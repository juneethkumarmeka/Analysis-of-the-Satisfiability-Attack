module basic_5000_50000_5000_200_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_209,In_4064);
nor U1 (N_1,In_3416,In_2806);
nor U2 (N_2,In_1955,In_4370);
nand U3 (N_3,In_710,In_4524);
xor U4 (N_4,In_1908,In_2531);
and U5 (N_5,In_4500,In_1269);
or U6 (N_6,In_4217,In_4065);
or U7 (N_7,In_3564,In_2818);
nor U8 (N_8,In_3344,In_1656);
nand U9 (N_9,In_2668,In_4730);
nor U10 (N_10,In_223,In_4246);
and U11 (N_11,In_1432,In_1037);
and U12 (N_12,In_3842,In_2400);
and U13 (N_13,In_3233,In_1011);
nor U14 (N_14,In_1521,In_2550);
xor U15 (N_15,In_4425,In_795);
xor U16 (N_16,In_3619,In_3058);
nand U17 (N_17,In_236,In_2948);
or U18 (N_18,In_3482,In_932);
xor U19 (N_19,In_1958,In_1401);
or U20 (N_20,In_128,In_1622);
nor U21 (N_21,In_3737,In_578);
nor U22 (N_22,In_2248,In_4617);
xnor U23 (N_23,In_100,In_4728);
nor U24 (N_24,In_4743,In_4794);
and U25 (N_25,In_2520,In_2383);
nand U26 (N_26,In_2378,In_2076);
xnor U27 (N_27,In_2064,In_3869);
nand U28 (N_28,In_1888,In_3661);
and U29 (N_29,In_1988,In_1490);
and U30 (N_30,In_3726,In_2697);
nand U31 (N_31,In_3751,In_3041);
xnor U32 (N_32,In_1885,In_2290);
and U33 (N_33,In_2964,In_676);
or U34 (N_34,In_4287,In_2757);
nor U35 (N_35,In_3969,In_78);
or U36 (N_36,In_904,In_120);
xnor U37 (N_37,In_3871,In_9);
nor U38 (N_38,In_3920,In_825);
and U39 (N_39,In_4045,In_277);
nand U40 (N_40,In_4355,In_2967);
nor U41 (N_41,In_1774,In_1479);
nand U42 (N_42,In_1067,In_4279);
xor U43 (N_43,In_2240,In_2274);
nand U44 (N_44,In_1499,In_989);
or U45 (N_45,In_351,In_3377);
and U46 (N_46,In_738,In_81);
or U47 (N_47,In_4595,In_2606);
xnor U48 (N_48,In_621,In_3068);
nand U49 (N_49,In_960,In_388);
nor U50 (N_50,In_2188,In_4536);
nand U51 (N_51,In_3879,In_560);
and U52 (N_52,In_3099,In_503);
nor U53 (N_53,In_1404,In_3831);
xor U54 (N_54,In_4593,In_2228);
xnor U55 (N_55,In_3629,In_1664);
and U56 (N_56,In_4791,In_1305);
nor U57 (N_57,In_1041,In_1472);
and U58 (N_58,In_1733,In_2437);
and U59 (N_59,In_4960,In_4163);
and U60 (N_60,In_766,In_4472);
xor U61 (N_61,In_2354,In_2051);
and U62 (N_62,In_838,In_3929);
nand U63 (N_63,In_776,In_792);
or U64 (N_64,In_268,In_1460);
nand U65 (N_65,In_1071,In_3115);
or U66 (N_66,In_2316,In_4106);
xnor U67 (N_67,In_2397,In_266);
xnor U68 (N_68,In_1098,In_4686);
and U69 (N_69,In_4248,In_4481);
xor U70 (N_70,In_453,In_1693);
nor U71 (N_71,In_1168,In_4720);
and U72 (N_72,In_2779,In_1250);
nand U73 (N_73,In_466,In_4012);
nor U74 (N_74,In_1073,In_481);
nor U75 (N_75,In_2505,In_3297);
or U76 (N_76,In_92,In_429);
nand U77 (N_77,In_3269,In_1862);
nor U78 (N_78,In_3353,In_1387);
nand U79 (N_79,In_1423,In_1678);
or U80 (N_80,In_1983,In_452);
or U81 (N_81,In_1528,In_3000);
and U82 (N_82,In_1261,In_927);
nand U83 (N_83,In_1308,In_2984);
and U84 (N_84,In_2225,In_3412);
xor U85 (N_85,In_4624,In_3317);
xnor U86 (N_86,In_4392,In_2702);
and U87 (N_87,In_4590,In_2280);
nand U88 (N_88,In_435,In_1430);
nor U89 (N_89,In_4809,In_3280);
nand U90 (N_90,In_3500,In_3817);
and U91 (N_91,In_3898,In_3565);
xnor U92 (N_92,In_1543,In_569);
nand U93 (N_93,In_2145,In_3473);
or U94 (N_94,In_2692,In_3571);
nand U95 (N_95,In_4373,In_3609);
nand U96 (N_96,In_4690,In_1502);
nor U97 (N_97,In_1378,In_106);
nor U98 (N_98,In_4316,In_422);
or U99 (N_99,In_1417,In_2582);
and U100 (N_100,In_1416,In_931);
xnor U101 (N_101,In_4171,In_2824);
nor U102 (N_102,In_1652,In_802);
or U103 (N_103,In_4134,In_4085);
xor U104 (N_104,In_1800,In_2499);
and U105 (N_105,In_3821,In_4519);
xor U106 (N_106,In_3931,In_4480);
xnor U107 (N_107,In_4840,In_4927);
or U108 (N_108,In_4745,In_3237);
nand U109 (N_109,In_4154,In_2935);
xnor U110 (N_110,In_1745,In_3947);
and U111 (N_111,In_4,In_2184);
or U112 (N_112,In_4311,In_817);
nand U113 (N_113,In_1277,In_3345);
nor U114 (N_114,In_3132,In_4240);
and U115 (N_115,In_2879,In_4748);
nand U116 (N_116,In_3531,In_2410);
and U117 (N_117,In_1796,In_4363);
nand U118 (N_118,In_2933,In_4994);
or U119 (N_119,In_2991,In_4409);
and U120 (N_120,In_2580,In_2099);
and U121 (N_121,In_1090,In_3277);
nor U122 (N_122,In_2937,In_1902);
nand U123 (N_123,In_2200,In_1253);
and U124 (N_124,In_1589,In_4461);
nor U125 (N_125,In_3962,In_2838);
and U126 (N_126,In_2601,In_3484);
nor U127 (N_127,In_2256,In_2516);
or U128 (N_128,In_896,In_3036);
or U129 (N_129,In_3550,In_1497);
or U130 (N_130,In_2124,In_2513);
xor U131 (N_131,In_2053,In_228);
nor U132 (N_132,In_4178,In_2976);
xor U133 (N_133,In_1730,In_2756);
and U134 (N_134,In_708,In_1706);
nand U135 (N_135,In_844,In_1035);
xnor U136 (N_136,In_918,In_4968);
nor U137 (N_137,In_4114,In_4605);
and U138 (N_138,In_3975,In_494);
xnor U139 (N_139,In_1957,In_3253);
or U140 (N_140,In_3949,In_3211);
and U141 (N_141,In_2556,In_4639);
nand U142 (N_142,In_478,In_1206);
nand U143 (N_143,In_2527,In_1389);
nand U144 (N_144,In_3305,In_1836);
xnor U145 (N_145,In_4868,In_1669);
xor U146 (N_146,In_4095,In_3026);
and U147 (N_147,In_2704,In_901);
and U148 (N_148,In_1402,In_1525);
nor U149 (N_149,In_3953,In_4371);
or U150 (N_150,In_255,In_3727);
or U151 (N_151,In_827,In_1886);
or U152 (N_152,In_2203,In_2627);
nor U153 (N_153,In_4061,In_2323);
or U154 (N_154,In_432,In_940);
xor U155 (N_155,In_1029,In_2363);
nor U156 (N_156,In_1360,In_859);
and U157 (N_157,In_2558,In_2685);
nor U158 (N_158,In_889,In_96);
nor U159 (N_159,In_3075,In_3187);
and U160 (N_160,In_1530,In_659);
nand U161 (N_161,In_1960,In_48);
and U162 (N_162,In_1439,In_1156);
nand U163 (N_163,In_1309,In_1150);
xor U164 (N_164,In_4517,In_4939);
or U165 (N_165,In_751,In_3653);
nand U166 (N_166,In_3426,In_1245);
or U167 (N_167,In_1200,In_4263);
nand U168 (N_168,In_1344,In_2707);
and U169 (N_169,In_2899,In_2968);
xor U170 (N_170,In_2444,In_303);
xor U171 (N_171,In_2414,In_3171);
or U172 (N_172,In_1271,In_3244);
and U173 (N_173,In_216,In_345);
xor U174 (N_174,In_2317,In_1461);
or U175 (N_175,In_4521,In_1992);
and U176 (N_176,In_448,In_715);
or U177 (N_177,In_3238,In_3232);
nor U178 (N_178,In_747,In_2713);
or U179 (N_179,In_788,In_1840);
and U180 (N_180,In_7,In_2574);
xor U181 (N_181,In_3159,In_2512);
or U182 (N_182,In_1816,In_2595);
or U183 (N_183,In_2063,In_3862);
nor U184 (N_184,In_1788,In_2628);
or U185 (N_185,In_3409,In_1809);
nand U186 (N_186,In_635,In_1354);
nand U187 (N_187,In_443,In_2086);
and U188 (N_188,In_3847,In_4169);
and U189 (N_189,In_4221,In_35);
nor U190 (N_190,In_2730,In_3538);
nor U191 (N_191,In_897,In_1446);
nand U192 (N_192,In_837,In_4261);
or U193 (N_193,In_4010,In_3596);
xnor U194 (N_194,In_3384,In_2615);
nand U195 (N_195,In_4274,In_2111);
and U196 (N_196,In_4360,In_794);
nand U197 (N_197,In_4553,In_1017);
or U198 (N_198,In_767,In_357);
or U199 (N_199,In_4842,In_3883);
xnor U200 (N_200,In_4199,In_1786);
nand U201 (N_201,In_1252,In_4667);
nand U202 (N_202,In_4244,In_3646);
and U203 (N_203,In_4034,In_4057);
and U204 (N_204,In_1743,In_436);
and U205 (N_205,In_4807,In_3177);
nor U206 (N_206,In_2850,In_3769);
and U207 (N_207,In_3508,In_4844);
nand U208 (N_208,In_4918,In_903);
nand U209 (N_209,In_2191,In_4328);
and U210 (N_210,In_1054,In_4225);
or U211 (N_211,In_2902,In_1143);
or U212 (N_212,In_1657,In_864);
nand U213 (N_213,In_3381,In_1667);
nand U214 (N_214,In_1165,In_2536);
or U215 (N_215,In_3833,In_4405);
or U216 (N_216,In_437,In_3865);
and U217 (N_217,In_2877,In_4945);
nand U218 (N_218,In_4419,In_1129);
or U219 (N_219,In_4305,In_2650);
xor U220 (N_220,In_3524,In_2896);
xnor U221 (N_221,In_224,In_275);
xor U222 (N_222,In_1567,In_958);
nand U223 (N_223,In_4789,In_4156);
and U224 (N_224,In_1692,In_95);
and U225 (N_225,In_3778,In_1659);
nand U226 (N_226,In_1620,In_3124);
xor U227 (N_227,In_1414,In_2958);
xor U228 (N_228,In_1611,In_4003);
nor U229 (N_229,In_4573,In_3835);
and U230 (N_230,In_2945,In_4857);
or U231 (N_231,In_4043,In_4951);
or U232 (N_232,In_302,In_2673);
nor U233 (N_233,In_3096,In_2570);
xor U234 (N_234,In_4346,In_4320);
nand U235 (N_235,In_1588,In_2277);
or U236 (N_236,In_3485,In_3723);
nand U237 (N_237,In_537,In_136);
xnor U238 (N_238,In_464,In_3888);
xor U239 (N_239,In_3364,In_4626);
xnor U240 (N_240,In_1734,In_641);
xnor U241 (N_241,In_1297,In_217);
or U242 (N_242,In_2807,In_1646);
and U243 (N_243,In_4837,In_4887);
xnor U244 (N_244,In_2551,In_575);
nor U245 (N_245,In_610,In_1122);
nor U246 (N_246,In_4008,In_3690);
xnor U247 (N_247,In_3383,In_227);
and U248 (N_248,In_1070,In_19);
and U249 (N_249,In_4737,In_482);
xnor U250 (N_250,In_4976,In_87);
or U251 (N_251,In_3884,In_4204);
nand U252 (N_252,In_3243,In_1428);
or U253 (N_253,In_2755,In_637);
and U254 (N_254,In_4428,In_948);
xnor U255 (N_255,In_2996,In_4841);
xnor U256 (N_256,In_16,In_2929);
nand U257 (N_257,N_145,In_3752);
nor U258 (N_258,In_4893,In_3556);
nor U259 (N_259,N_71,In_4139);
nor U260 (N_260,In_744,In_4660);
and U261 (N_261,In_3094,In_108);
nand U262 (N_262,In_1556,In_3189);
and U263 (N_263,In_2738,In_3521);
xor U264 (N_264,In_1393,In_3441);
xor U265 (N_265,In_699,In_3714);
nand U266 (N_266,In_2117,In_4440);
and U267 (N_267,In_3415,In_1107);
xnor U268 (N_268,In_3807,In_381);
nand U269 (N_269,In_4591,In_2503);
xor U270 (N_270,In_4990,In_4804);
nor U271 (N_271,In_4533,In_389);
nor U272 (N_272,In_1237,N_24);
or U273 (N_273,In_129,In_14);
nand U274 (N_274,In_4056,In_4909);
and U275 (N_275,In_427,In_850);
and U276 (N_276,In_1986,In_3776);
nand U277 (N_277,In_1368,In_815);
xor U278 (N_278,In_3991,In_3860);
or U279 (N_279,In_2408,In_204);
or U280 (N_280,In_2584,In_4736);
xnor U281 (N_281,In_2997,In_401);
xor U282 (N_282,In_2176,In_1384);
or U283 (N_283,In_2889,In_1984);
nor U284 (N_284,In_2081,In_2645);
and U285 (N_285,In_3555,In_3301);
xnor U286 (N_286,In_3056,In_2908);
nand U287 (N_287,In_1766,In_470);
or U288 (N_288,In_492,In_632);
and U289 (N_289,N_98,N_111);
xor U290 (N_290,N_110,In_4278);
nor U291 (N_291,In_1415,In_2067);
nand U292 (N_292,In_1487,In_3527);
xnor U293 (N_293,In_505,In_461);
or U294 (N_294,In_994,In_1959);
nor U295 (N_295,In_2494,In_1382);
nor U296 (N_296,In_1927,In_3464);
xnor U297 (N_297,In_4635,In_3985);
or U298 (N_298,In_619,In_4268);
nor U299 (N_299,In_3276,In_4167);
xor U300 (N_300,In_556,In_1560);
xnor U301 (N_301,In_2583,In_2987);
nand U302 (N_302,In_1887,In_2796);
nor U303 (N_303,In_3598,In_3558);
and U304 (N_304,In_2093,In_2624);
xor U305 (N_305,In_2537,In_1023);
and U306 (N_306,In_2275,In_2508);
xnor U307 (N_307,In_2544,In_1449);
and U308 (N_308,In_1194,In_2241);
nand U309 (N_309,In_3761,In_4972);
or U310 (N_310,In_3729,In_174);
nor U311 (N_311,In_772,In_2440);
or U312 (N_312,In_2123,In_4486);
nor U313 (N_313,In_664,In_431);
xor U314 (N_314,In_2001,N_109);
and U315 (N_315,In_1863,In_3293);
or U316 (N_316,In_4779,In_1127);
and U317 (N_317,In_4997,In_4172);
xnor U318 (N_318,In_3667,In_4788);
xnor U319 (N_319,In_3624,In_3675);
nand U320 (N_320,In_424,In_72);
nor U321 (N_321,In_4019,In_891);
or U322 (N_322,In_2263,In_1913);
xor U323 (N_323,In_949,In_4487);
or U324 (N_324,In_3070,In_4739);
nor U325 (N_325,In_3337,In_373);
nor U326 (N_326,In_1830,In_159);
and U327 (N_327,In_2898,In_2151);
xor U328 (N_328,In_2517,In_2119);
xor U329 (N_329,In_4120,In_2449);
xor U330 (N_330,In_3091,In_2847);
xnor U331 (N_331,In_2082,In_4304);
xnor U332 (N_332,In_806,In_391);
nor U333 (N_333,In_4787,In_1105);
and U334 (N_334,In_1495,In_3081);
nor U335 (N_335,In_4820,In_3210);
or U336 (N_336,In_440,In_4026);
nor U337 (N_337,In_4477,In_2614);
nand U338 (N_338,In_663,In_310);
or U339 (N_339,In_3637,In_1142);
nand U340 (N_340,In_1114,In_1741);
xor U341 (N_341,In_3939,In_3150);
nand U342 (N_342,In_2459,In_4239);
xnor U343 (N_343,In_4529,In_867);
and U344 (N_344,In_3891,In_2425);
xnor U345 (N_345,In_3529,In_273);
or U346 (N_346,In_3168,In_2046);
xnor U347 (N_347,In_4883,N_155);
or U348 (N_348,In_3162,In_1680);
nand U349 (N_349,In_3618,In_3432);
or U350 (N_350,In_4954,In_2072);
nand U351 (N_351,In_1333,In_314);
nand U352 (N_352,In_4333,In_1034);
xor U353 (N_353,In_608,In_2174);
or U354 (N_354,In_1493,In_856);
or U355 (N_355,In_2320,In_2735);
nor U356 (N_356,In_2025,In_982);
and U357 (N_357,In_4522,In_3288);
and U358 (N_358,In_667,In_1334);
nand U359 (N_359,In_1221,In_3530);
nor U360 (N_360,In_2457,In_3850);
or U361 (N_361,N_72,In_4413);
and U362 (N_362,In_2532,In_442);
and U363 (N_363,In_2170,In_2742);
and U364 (N_364,In_2985,In_4141);
nor U365 (N_365,In_4295,In_4862);
xor U366 (N_366,In_4738,In_316);
nand U367 (N_367,In_2166,In_934);
or U368 (N_368,In_4859,In_113);
nand U369 (N_369,In_1128,N_176);
and U370 (N_370,In_3837,In_4438);
or U371 (N_371,In_3016,In_4116);
xor U372 (N_372,In_616,In_3010);
nor U373 (N_373,In_4614,N_75);
or U374 (N_374,N_28,In_2179);
nand U375 (N_375,In_4429,In_2456);
nor U376 (N_376,In_1909,In_2514);
and U377 (N_377,In_1329,N_125);
or U378 (N_378,In_2481,In_1636);
xnor U379 (N_379,In_1939,In_1813);
nand U380 (N_380,In_3780,In_2815);
nor U381 (N_381,In_4389,In_3321);
or U382 (N_382,In_730,In_3589);
and U383 (N_383,In_3622,In_4931);
and U384 (N_384,In_1640,In_2788);
or U385 (N_385,In_1281,In_1290);
nand U386 (N_386,In_318,In_4645);
and U387 (N_387,In_648,In_2792);
or U388 (N_388,In_3736,In_4619);
and U389 (N_389,In_1244,In_2522);
or U390 (N_390,In_3701,In_4161);
xor U391 (N_391,In_1954,In_2428);
nor U392 (N_392,In_2011,In_4797);
xor U393 (N_393,In_3586,In_1369);
and U394 (N_394,In_942,In_961);
xor U395 (N_395,In_1028,In_4588);
xnor U396 (N_396,In_409,In_915);
or U397 (N_397,In_4391,In_149);
or U398 (N_398,In_3648,In_1973);
nor U399 (N_399,In_2862,In_842);
or U400 (N_400,In_46,In_4688);
nand U401 (N_401,In_2905,In_4946);
nor U402 (N_402,In_1058,In_3015);
nor U403 (N_403,In_1690,In_3332);
nor U404 (N_404,In_706,In_3421);
and U405 (N_405,In_1106,In_2100);
or U406 (N_406,In_4041,In_1650);
xnor U407 (N_407,In_4266,In_1896);
xor U408 (N_408,N_172,N_19);
nor U409 (N_409,In_40,In_4290);
nand U410 (N_410,N_102,In_990);
nor U411 (N_411,In_967,In_116);
or U412 (N_412,In_2127,In_2804);
xnor U413 (N_413,In_2292,In_2342);
nand U414 (N_414,N_216,In_2836);
nand U415 (N_415,In_589,In_2830);
nor U416 (N_416,In_1010,In_1931);
nor U417 (N_417,In_564,In_4707);
and U418 (N_418,In_3104,In_4498);
and U419 (N_419,In_964,In_3513);
nor U420 (N_420,N_201,In_2473);
nor U421 (N_421,In_1578,In_4042);
or U422 (N_422,In_4582,In_2092);
nand U423 (N_423,In_3102,In_1781);
or U424 (N_424,In_2484,In_613);
nor U425 (N_425,In_1408,In_438);
nand U426 (N_426,In_4881,In_2351);
nand U427 (N_427,In_2839,N_164);
and U428 (N_428,In_1398,In_847);
or U429 (N_429,In_146,In_4032);
or U430 (N_430,In_3234,In_4080);
nand U431 (N_431,In_530,In_3823);
nand U432 (N_432,In_1634,In_654);
and U433 (N_433,In_1022,In_4740);
or U434 (N_434,In_2500,In_3764);
nor U435 (N_435,In_3781,In_2825);
nand U436 (N_436,In_4592,In_4082);
nor U437 (N_437,In_3106,N_185);
xor U438 (N_438,N_165,In_528);
nor U439 (N_439,In_3362,In_3155);
or U440 (N_440,In_2284,In_3628);
nor U441 (N_441,In_4983,In_2315);
nor U442 (N_442,In_3385,In_2222);
nor U443 (N_443,In_1649,In_184);
xnor U444 (N_444,In_454,In_4917);
nor U445 (N_445,In_4022,In_3536);
nand U446 (N_446,In_235,In_2333);
xnor U447 (N_447,In_3007,In_3797);
nor U448 (N_448,In_2157,In_274);
xor U449 (N_449,N_161,In_3148);
nor U450 (N_450,In_3625,In_3945);
nor U451 (N_451,In_294,In_4603);
nand U452 (N_452,In_3760,In_2926);
nand U453 (N_453,In_1085,In_1306);
xor U454 (N_454,In_1944,N_48);
xnor U455 (N_455,In_2758,N_235);
nor U456 (N_456,In_3291,In_951);
and U457 (N_457,In_1714,N_33);
nor U458 (N_458,In_4712,In_3899);
and U459 (N_459,In_3181,In_1431);
nand U460 (N_460,In_4280,In_1923);
nor U461 (N_461,In_1370,In_1895);
or U462 (N_462,In_143,In_2693);
nand U463 (N_463,In_740,In_4648);
xor U464 (N_464,In_45,In_4212);
and U465 (N_465,N_205,In_3188);
nand U466 (N_466,In_3396,In_2547);
xnor U467 (N_467,In_313,In_1691);
and U468 (N_468,In_3614,In_1440);
nor U469 (N_469,In_286,In_2015);
nor U470 (N_470,In_4299,In_3496);
and U471 (N_471,In_1376,In_1219);
xor U472 (N_472,In_2963,In_4494);
xor U473 (N_473,In_2657,In_4604);
and U474 (N_474,In_1814,In_1110);
or U475 (N_475,In_529,In_4924);
nor U476 (N_476,In_3656,In_688);
nor U477 (N_477,In_4766,In_1198);
xor U478 (N_478,In_2366,In_4991);
nor U479 (N_479,In_3204,In_1558);
and U480 (N_480,In_2364,In_3959);
nor U481 (N_481,In_4811,In_1783);
xor U482 (N_482,In_3501,In_292);
or U483 (N_483,In_3429,In_3551);
or U484 (N_484,In_4324,In_628);
or U485 (N_485,In_2922,In_1409);
nand U486 (N_486,In_4051,In_3987);
xor U487 (N_487,In_2856,In_2700);
and U488 (N_488,In_853,In_4399);
xor U489 (N_489,In_1183,In_3014);
or U490 (N_490,In_3052,N_38);
nand U491 (N_491,In_720,In_1551);
nand U492 (N_492,In_317,In_2307);
xnor U493 (N_493,N_232,In_4164);
nor U494 (N_494,In_119,In_179);
nand U495 (N_495,In_970,In_1832);
nor U496 (N_496,In_1314,In_2762);
nor U497 (N_497,In_4272,In_4584);
xnor U498 (N_498,In_4833,In_2533);
or U499 (N_499,N_26,In_1249);
and U500 (N_500,In_3072,In_2541);
nand U501 (N_501,In_2143,In_3679);
xnor U502 (N_502,In_2680,In_2266);
nor U503 (N_503,In_1116,In_3897);
nor U504 (N_504,In_4416,In_68);
nand U505 (N_505,In_1214,In_1737);
or U506 (N_506,In_781,In_4928);
xnor U507 (N_507,In_1554,In_3575);
xnor U508 (N_508,In_4180,In_3996);
xor U509 (N_509,In_649,In_97);
or U510 (N_510,In_894,In_4724);
xnor U511 (N_511,N_319,In_1676);
or U512 (N_512,In_4979,In_1710);
nor U513 (N_513,In_2927,N_35);
xnor U514 (N_514,In_4150,In_3105);
xor U515 (N_515,In_3095,In_919);
nand U516 (N_516,N_285,In_4159);
xnor U517 (N_517,In_3065,In_109);
or U518 (N_518,N_277,In_681);
nand U519 (N_519,In_3319,In_3370);
nor U520 (N_520,In_826,In_3687);
nor U521 (N_521,In_3922,In_3854);
xnor U522 (N_522,N_340,In_1280);
or U523 (N_523,In_1831,In_647);
nor U524 (N_524,In_1454,In_1727);
nand U525 (N_525,In_156,In_13);
nand U526 (N_526,In_1731,In_1317);
xor U527 (N_527,N_225,In_1891);
xnor U528 (N_528,In_752,In_711);
or U529 (N_529,In_3918,In_2640);
or U530 (N_530,In_2813,In_4652);
and U531 (N_531,In_2108,In_598);
or U532 (N_532,N_179,In_3641);
or U533 (N_533,In_3405,In_1803);
xnor U534 (N_534,In_2552,In_4067);
and U535 (N_535,N_93,In_2027);
nor U536 (N_536,In_3912,In_1291);
nand U537 (N_537,N_105,In_4744);
nor U538 (N_538,In_4356,In_4950);
and U539 (N_539,In_816,In_1374);
nand U540 (N_540,In_3858,In_4108);
xor U541 (N_541,In_3404,In_1117);
or U542 (N_542,In_1477,In_3433);
or U543 (N_543,N_312,In_4113);
or U544 (N_544,In_2095,In_2014);
and U545 (N_545,In_4802,In_1043);
nand U546 (N_546,In_2309,In_714);
nor U547 (N_547,In_3042,In_3844);
nand U548 (N_548,In_127,In_2385);
and U549 (N_549,N_303,In_3263);
and U550 (N_550,In_150,In_469);
nor U551 (N_551,In_2587,In_3469);
and U552 (N_552,In_2369,In_4236);
nor U553 (N_553,In_1205,In_692);
xnor U554 (N_554,N_301,In_4670);
nand U555 (N_555,In_732,In_44);
and U556 (N_556,In_3284,N_188);
or U557 (N_557,In_1753,In_1789);
xnor U558 (N_558,In_3895,In_4235);
nand U559 (N_559,N_84,In_1982);
nor U560 (N_560,In_1671,In_1538);
nor U561 (N_561,In_3549,N_446);
nand U562 (N_562,In_477,In_3515);
and U563 (N_563,In_4258,In_705);
xor U564 (N_564,N_375,In_349);
or U565 (N_565,In_3574,In_3427);
or U566 (N_566,N_450,In_539);
nor U567 (N_567,In_1381,In_3503);
and U568 (N_568,In_565,In_1158);
or U569 (N_569,In_1050,In_219);
or U570 (N_570,In_3061,In_1695);
xor U571 (N_571,In_3805,In_2764);
nand U572 (N_572,In_1042,In_4891);
and U573 (N_573,In_4062,In_1841);
nand U574 (N_574,In_629,In_3110);
nand U575 (N_575,In_3604,In_3399);
xnor U576 (N_576,In_300,In_1759);
xnor U577 (N_577,In_4735,In_3180);
nor U578 (N_578,In_836,In_1777);
nor U579 (N_579,N_306,In_1049);
or U580 (N_580,In_1192,In_3649);
nand U581 (N_581,In_3479,In_2895);
nor U582 (N_582,In_15,In_3859);
or U583 (N_583,In_1413,In_4096);
and U584 (N_584,In_3191,In_1492);
nor U585 (N_585,N_354,In_1104);
nand U586 (N_586,In_226,In_3818);
and U587 (N_587,In_793,N_401);
or U588 (N_588,In_1264,In_3779);
and U589 (N_589,In_66,In_848);
nor U590 (N_590,N_66,In_3672);
nor U591 (N_591,In_4310,In_3999);
xnor U592 (N_592,In_4622,In_3491);
nand U593 (N_593,In_3149,In_1696);
nor U594 (N_594,N_376,In_4332);
or U595 (N_595,In_499,In_4072);
xnor U596 (N_596,In_258,In_293);
xor U597 (N_597,In_1508,In_3126);
nor U598 (N_598,In_2431,In_3800);
nand U599 (N_599,In_1820,In_1977);
xor U600 (N_600,In_2163,In_1421);
nor U601 (N_601,In_1824,N_283);
and U602 (N_602,In_3223,In_37);
xor U603 (N_603,In_1467,In_3033);
xnor U604 (N_604,In_3299,In_3815);
xor U605 (N_605,N_332,N_260);
xor U606 (N_606,In_3356,In_765);
or U607 (N_607,In_2142,In_1003);
nand U608 (N_608,In_4339,In_1853);
nand U609 (N_609,In_346,In_1044);
and U610 (N_610,N_103,In_2182);
nor U611 (N_611,In_2297,In_625);
or U612 (N_612,In_355,In_4663);
nand U613 (N_613,In_2303,In_818);
and U614 (N_614,In_4723,In_702);
and U615 (N_615,In_1687,In_1570);
or U616 (N_616,In_1856,In_2686);
or U617 (N_617,In_2107,In_2080);
xnor U618 (N_618,In_3542,In_2827);
xnor U619 (N_619,In_2068,In_3376);
and U620 (N_620,In_4117,N_57);
nor U621 (N_621,In_3227,In_220);
or U622 (N_622,In_2597,In_2507);
xnor U623 (N_623,In_457,In_3788);
xor U624 (N_624,In_3363,In_2348);
xnor U625 (N_625,In_3795,In_337);
nand U626 (N_626,In_4434,In_4759);
nand U627 (N_627,In_1412,In_2585);
or U628 (N_628,In_368,In_3594);
nand U629 (N_629,In_3452,In_2132);
nand U630 (N_630,N_5,N_482);
xnor U631 (N_631,N_112,In_3430);
xor U632 (N_632,In_187,In_1956);
xnor U633 (N_633,In_1924,In_4218);
or U634 (N_634,N_108,In_2299);
or U635 (N_635,In_4121,In_4650);
or U636 (N_636,In_4701,In_3450);
and U637 (N_637,In_2038,In_4623);
or U638 (N_638,In_543,In_1286);
or U639 (N_639,In_1683,In_4646);
xnor U640 (N_640,In_4183,In_779);
nand U641 (N_641,In_2442,In_3744);
or U642 (N_642,In_4685,In_3419);
and U643 (N_643,In_4515,In_3792);
xor U644 (N_644,In_2740,In_1482);
or U645 (N_645,In_2474,In_4301);
nand U646 (N_646,In_922,In_4550);
xor U647 (N_647,In_3179,In_2468);
or U648 (N_648,In_4963,In_4559);
nand U649 (N_649,In_585,In_3047);
or U650 (N_650,In_2511,N_209);
and U651 (N_651,In_4048,In_2344);
nand U652 (N_652,In_2268,In_11);
xnor U653 (N_653,N_76,In_1320);
xnor U654 (N_654,N_180,In_2821);
or U655 (N_655,In_3057,In_2773);
and U656 (N_656,In_2175,In_1364);
nand U657 (N_657,In_397,In_3765);
and U658 (N_658,In_504,In_661);
nor U659 (N_659,In_3514,In_3930);
nor U660 (N_660,In_58,In_3497);
xnor U661 (N_661,In_3108,In_500);
or U662 (N_662,In_1858,In_4763);
nor U663 (N_663,In_1780,In_1749);
or U664 (N_664,In_1903,In_3205);
xor U665 (N_665,In_4826,In_4027);
xor U666 (N_666,In_2956,In_197);
nor U667 (N_667,N_380,In_607);
nor U668 (N_668,In_4307,In_4255);
nor U669 (N_669,N_392,In_2765);
and U670 (N_670,In_4147,In_3853);
nor U671 (N_671,N_341,In_1509);
nor U672 (N_672,In_2881,In_3437);
or U673 (N_673,In_1263,In_416);
nand U674 (N_674,In_396,In_4849);
nand U675 (N_675,In_4975,In_2489);
or U676 (N_676,In_232,N_449);
xnor U677 (N_677,In_1920,In_2720);
nand U678 (N_678,In_1694,In_536);
nand U679 (N_679,In_3798,In_4656);
xnor U680 (N_680,In_2975,In_4467);
nor U681 (N_681,In_3086,In_2102);
xnor U682 (N_682,In_1585,In_1137);
nor U683 (N_683,In_624,In_304);
and U684 (N_684,In_916,In_1052);
and U685 (N_685,In_4662,In_3163);
nor U686 (N_686,In_4230,In_2699);
nand U687 (N_687,In_4913,In_332);
and U688 (N_688,In_3134,In_4375);
and U689 (N_689,In_2805,In_4796);
xnor U690 (N_690,In_1770,In_3613);
or U691 (N_691,In_2868,In_1091);
or U692 (N_692,In_2273,In_563);
nor U693 (N_693,In_2696,In_2147);
or U694 (N_694,In_614,In_521);
or U695 (N_695,In_2387,In_1867);
or U696 (N_696,In_572,In_1631);
or U697 (N_697,In_3926,In_1025);
nor U698 (N_698,In_3490,N_339);
or U699 (N_699,In_2078,In_4607);
or U700 (N_700,N_477,In_3864);
nor U701 (N_701,In_1846,In_3201);
or U702 (N_702,In_155,In_4490);
nand U703 (N_703,In_2793,In_3591);
xor U704 (N_704,N_409,In_390);
nand U705 (N_705,In_4189,In_463);
nor U706 (N_706,In_3995,In_4110);
or U707 (N_707,In_1583,In_3826);
and U708 (N_708,In_2594,In_2942);
xnor U709 (N_709,N_274,In_3060);
nor U710 (N_710,In_2656,In_2204);
nand U711 (N_711,In_2155,In_1892);
xnor U712 (N_712,In_4866,In_4651);
xor U713 (N_713,N_0,In_876);
xor U714 (N_714,N_237,In_2834);
nor U715 (N_715,In_3846,In_2024);
nand U716 (N_716,N_271,In_4644);
or U717 (N_717,In_4502,N_146);
nand U718 (N_718,In_1310,In_3287);
xnor U719 (N_719,In_4308,In_4297);
nand U720 (N_720,In_1875,N_284);
xnor U721 (N_721,In_3983,In_1148);
or U722 (N_722,In_4111,In_1469);
nand U723 (N_723,N_472,In_1187);
or U724 (N_724,In_2258,In_3537);
nand U725 (N_725,In_1964,In_2392);
nand U726 (N_726,In_2045,In_25);
or U727 (N_727,In_1438,In_2719);
and U728 (N_728,In_3,In_1377);
or U729 (N_729,In_47,In_3829);
nor U730 (N_730,In_176,In_2158);
nor U731 (N_731,In_3819,In_4300);
and U732 (N_732,In_4282,In_580);
nor U733 (N_733,In_507,In_428);
xor U734 (N_734,In_4873,In_4511);
xnor U735 (N_735,In_943,In_21);
xnor U736 (N_736,N_259,In_4403);
and U737 (N_737,In_4845,In_4875);
xnor U738 (N_738,In_2436,In_3323);
xnor U739 (N_739,In_1778,In_430);
nand U740 (N_740,In_973,In_944);
or U741 (N_741,In_803,In_561);
nor U742 (N_742,In_1870,In_1522);
nand U743 (N_743,In_203,In_3137);
xor U744 (N_744,N_9,In_4450);
or U745 (N_745,In_1178,In_3794);
and U746 (N_746,In_4816,In_4534);
xor U747 (N_747,In_1092,In_4288);
and U748 (N_748,In_712,In_2608);
and U749 (N_749,N_183,In_387);
nor U750 (N_750,In_1260,In_2831);
xnor U751 (N_751,N_157,N_25);
xor U752 (N_752,In_105,N_100);
or U753 (N_753,In_4475,In_1099);
or U754 (N_754,In_1392,In_4241);
and U755 (N_755,In_2289,In_3241);
or U756 (N_756,In_170,In_4458);
xnor U757 (N_757,In_1450,In_4703);
or U758 (N_758,In_1582,In_1204);
nand U759 (N_759,In_2033,N_126);
and U760 (N_760,In_832,In_1352);
and U761 (N_761,In_324,N_115);
xnor U762 (N_762,In_3247,In_952);
nor U763 (N_763,In_177,In_2869);
or U764 (N_764,In_1940,In_3138);
or U765 (N_765,In_2169,In_1532);
and U766 (N_766,N_293,In_579);
xnor U767 (N_767,In_4423,N_489);
and U768 (N_768,In_4633,In_2007);
xor U769 (N_769,In_1436,In_3013);
and U770 (N_770,In_421,In_3109);
nor U771 (N_771,In_3216,In_2778);
nor U772 (N_772,In_3318,In_898);
xnor U773 (N_773,N_97,In_2485);
nand U774 (N_774,In_3342,In_1765);
nand U775 (N_775,In_4503,N_445);
or U776 (N_776,In_4036,In_3877);
or U777 (N_777,In_2048,In_2106);
or U778 (N_778,In_3526,In_2801);
and U779 (N_779,In_2446,In_3382);
nor U780 (N_780,In_953,In_4585);
or U781 (N_781,In_2578,In_4586);
and U782 (N_782,In_1096,In_3250);
xor U783 (N_783,In_2849,In_2662);
xnor U784 (N_784,In_3902,In_633);
nor U785 (N_785,In_4974,N_357);
nor U786 (N_786,In_2465,In_2853);
or U787 (N_787,In_3278,N_367);
or U788 (N_788,In_2949,In_4471);
or U789 (N_789,In_2098,In_1324);
xor U790 (N_790,N_484,In_1705);
and U791 (N_791,In_379,In_4693);
nand U792 (N_792,In_2802,In_142);
nand U793 (N_793,In_1849,In_282);
nor U794 (N_794,In_1597,In_3784);
and U795 (N_795,In_713,In_1945);
and U796 (N_796,In_1575,In_4944);
and U797 (N_797,In_1894,In_2034);
xnor U798 (N_798,N_243,In_4247);
nor U799 (N_799,In_1174,In_3226);
nor U800 (N_800,In_131,In_1321);
nor U801 (N_801,In_189,N_169);
nor U802 (N_802,In_4099,N_671);
or U803 (N_803,N_512,In_3669);
xor U804 (N_804,In_3261,In_4277);
nand U805 (N_805,N_178,In_4906);
xor U806 (N_806,In_153,N_667);
xor U807 (N_807,In_995,In_399);
or U808 (N_808,In_4675,In_330);
xnor U809 (N_809,In_798,N_17);
nand U810 (N_810,N_657,N_44);
nand U811 (N_811,N_523,In_1235);
and U812 (N_812,In_2790,In_4805);
or U813 (N_813,In_4131,In_3135);
and U814 (N_814,In_190,In_270);
nor U815 (N_815,In_3657,In_2377);
or U816 (N_816,In_555,In_103);
nor U817 (N_817,In_2005,In_2291);
nand U818 (N_818,In_2978,In_2832);
or U819 (N_819,In_2314,N_190);
and U820 (N_820,In_3934,N_252);
and U821 (N_821,N_287,N_456);
nor U822 (N_822,N_692,N_563);
or U823 (N_823,In_1861,In_473);
nor U824 (N_824,In_2682,In_3742);
or U825 (N_825,In_2950,In_3249);
and U826 (N_826,In_1750,In_2596);
xor U827 (N_827,In_1303,In_2331);
or U828 (N_828,In_557,In_3114);
and U829 (N_829,N_162,In_2321);
nor U830 (N_830,In_4023,In_2739);
and U831 (N_831,N_461,In_4599);
and U832 (N_832,In_1203,In_2523);
and U833 (N_833,In_1462,In_4388);
or U834 (N_834,N_415,In_3209);
nand U835 (N_835,In_3878,N_470);
nor U836 (N_836,In_650,In_3569);
or U837 (N_837,In_2710,In_1553);
nor U838 (N_838,In_1076,In_2282);
and U839 (N_839,In_2144,In_2412);
xnor U840 (N_840,In_3043,In_2096);
xor U841 (N_841,In_4283,N_273);
xnor U842 (N_842,In_376,In_3360);
xnor U843 (N_843,N_447,N_649);
or U844 (N_844,N_278,In_3502);
or U845 (N_845,In_719,In_2477);
and U846 (N_846,In_487,In_3271);
or U847 (N_847,In_3044,In_1039);
nor U848 (N_848,In_1818,In_4075);
nor U849 (N_849,N_628,N_604);
nand U850 (N_850,In_4101,In_2355);
xnor U851 (N_851,In_1080,In_508);
and U852 (N_852,In_4160,In_288);
or U853 (N_853,In_1637,In_3395);
nand U854 (N_854,N_352,In_414);
nand U855 (N_855,N_292,In_985);
nand U856 (N_856,In_3700,N_618);
and U857 (N_857,N_742,N_624);
and U858 (N_858,In_1523,In_1976);
nand U859 (N_859,In_353,In_2122);
or U860 (N_860,In_1593,In_760);
or U861 (N_861,N_707,N_732);
and U862 (N_862,In_364,In_4385);
nor U863 (N_863,In_2610,In_1292);
and U864 (N_864,In_3129,N_730);
or U865 (N_865,In_3825,N_137);
and U866 (N_866,In_601,In_1708);
and U867 (N_867,In_137,N_212);
or U868 (N_868,In_2690,N_497);
nor U869 (N_869,In_1391,N_699);
nand U870 (N_870,N_602,In_4143);
nand U871 (N_871,In_3467,In_4476);
nand U872 (N_872,In_384,In_3265);
or U873 (N_873,In_4709,In_60);
xnor U874 (N_874,N_454,In_3488);
nand U875 (N_875,In_3198,In_2006);
xnor U876 (N_876,In_814,In_479);
xnor U877 (N_877,In_1934,N_211);
or U878 (N_878,In_3466,In_3196);
nor U879 (N_879,In_4412,In_4700);
and U880 (N_880,N_52,N_174);
xor U881 (N_881,In_4215,In_1488);
or U882 (N_882,In_3686,N_379);
xor U883 (N_883,In_2934,In_2525);
nand U884 (N_884,In_2218,In_551);
and U885 (N_885,In_3706,In_1);
and U886 (N_886,In_4665,In_61);
nand U887 (N_887,In_1890,In_4013);
nand U888 (N_888,N_316,In_359);
xor U889 (N_889,In_4465,In_3548);
and U890 (N_890,In_3358,In_3932);
nor U891 (N_891,In_3937,N_427);
nor U892 (N_892,In_88,In_999);
nand U893 (N_893,In_917,In_683);
nor U894 (N_894,In_2510,In_761);
or U895 (N_895,In_1160,In_2890);
nand U896 (N_896,In_3562,In_568);
and U897 (N_897,In_2833,In_3621);
or U898 (N_898,In_340,In_4806);
or U899 (N_899,In_1776,In_2837);
nor U900 (N_900,In_4882,In_1397);
nor U901 (N_901,In_4396,In_3992);
and U902 (N_902,N_451,In_4758);
nor U903 (N_903,In_1967,In_3777);
xnor U904 (N_904,In_1529,In_2193);
and U905 (N_905,In_3103,N_214);
nor U906 (N_906,In_3031,In_3650);
nor U907 (N_907,In_3365,In_1215);
xor U908 (N_908,In_3012,In_1876);
or U909 (N_909,In_2185,In_4947);
xnor U910 (N_910,In_3248,N_87);
xnor U911 (N_911,In_4188,In_4819);
nand U912 (N_912,In_4902,In_1715);
or U913 (N_913,In_2115,N_432);
nand U914 (N_914,N_331,In_3127);
nor U915 (N_915,In_801,In_3228);
nand U916 (N_916,In_344,In_3647);
nor U917 (N_917,In_1139,N_573);
nor U918 (N_918,In_1760,In_1661);
nor U919 (N_919,In_4233,In_725);
xnor U920 (N_920,N_503,In_1184);
nand U921 (N_921,In_4361,In_2665);
and U922 (N_922,In_311,In_1141);
or U923 (N_923,In_1170,In_407);
and U924 (N_924,In_2036,In_2725);
and U925 (N_925,N_711,In_4190);
or U926 (N_926,In_1751,In_3214);
and U927 (N_927,In_4336,In_1806);
nand U928 (N_928,In_3768,In_2017);
nand U929 (N_929,In_2463,In_3772);
xor U930 (N_930,In_1238,In_4822);
and U931 (N_931,In_2953,In_778);
or U932 (N_932,In_2162,In_888);
nor U933 (N_933,In_789,N_74);
or U934 (N_934,In_3541,In_3944);
xor U935 (N_935,In_1212,N_683);
nand U936 (N_936,N_498,N_625);
or U937 (N_937,N_159,In_495);
nor U938 (N_938,In_3112,In_2518);
xnor U939 (N_939,In_2808,N_589);
or U940 (N_940,In_3528,N_324);
nor U941 (N_941,In_3525,In_1026);
nor U942 (N_942,N_641,N_517);
xor U943 (N_943,In_858,In_2567);
and U944 (N_944,In_2037,In_233);
nor U945 (N_945,In_12,In_3048);
nand U946 (N_946,N_203,In_2864);
nor U947 (N_947,N_32,N_55);
or U948 (N_948,In_4291,In_4460);
nand U949 (N_949,In_1182,In_4276);
or U950 (N_950,In_3139,In_3793);
or U951 (N_951,In_1325,In_402);
nor U952 (N_952,In_1100,In_532);
nor U953 (N_953,In_3583,In_2221);
or U954 (N_954,N_239,In_1282);
nor U955 (N_955,In_2763,N_236);
xor U956 (N_956,In_4334,In_3329);
and U957 (N_957,In_2391,In_4808);
or U958 (N_958,In_2695,In_2466);
nand U959 (N_959,In_83,In_4629);
nand U960 (N_960,N_719,In_2694);
nor U961 (N_961,In_2324,In_4015);
nor U962 (N_962,In_1494,In_1994);
xor U963 (N_963,In_4774,In_2646);
xnor U964 (N_964,In_205,In_1524);
nand U965 (N_965,In_380,In_2125);
nand U966 (N_966,In_1399,In_1501);
or U967 (N_967,In_2009,In_4920);
and U968 (N_968,In_1990,In_2794);
or U969 (N_969,N_364,In_1763);
nor U970 (N_970,In_206,N_429);
xnor U971 (N_971,In_4242,N_231);
or U972 (N_972,N_654,In_604);
nor U973 (N_973,In_2564,In_1612);
or U974 (N_974,In_3231,In_2407);
nor U975 (N_975,In_4400,In_4044);
or U976 (N_976,In_1843,In_1180);
nand U977 (N_977,N_34,In_4801);
and U978 (N_978,In_2302,In_1700);
xor U979 (N_979,In_2283,In_4961);
xor U980 (N_980,In_3140,In_1859);
or U981 (N_981,N_666,In_3292);
xor U982 (N_982,In_2070,In_1302);
nor U983 (N_983,In_3388,N_234);
and U984 (N_984,In_465,N_601);
nand U985 (N_985,N_575,N_88);
or U986 (N_986,N_463,In_2878);
or U987 (N_987,In_3296,In_4817);
xor U988 (N_988,In_3767,In_1388);
and U989 (N_989,N_485,In_4296);
nor U990 (N_990,In_1752,In_2939);
nor U991 (N_991,N_525,In_41);
or U992 (N_992,In_1557,In_2245);
xor U993 (N_993,In_3724,In_2938);
or U994 (N_994,In_2236,In_1845);
or U995 (N_995,In_3523,In_231);
nand U996 (N_996,N_264,N_356);
xor U997 (N_997,In_4322,In_4831);
nor U998 (N_998,In_2897,N_734);
or U999 (N_999,In_2893,In_2008);
nor U1000 (N_1000,N_101,In_1294);
xor U1001 (N_1001,N_3,In_2050);
nand U1002 (N_1002,N_223,In_200);
nor U1003 (N_1003,In_4436,In_3511);
nand U1004 (N_1004,In_2913,In_913);
and U1005 (N_1005,In_2654,In_2661);
nand U1006 (N_1006,N_394,In_1190);
nor U1007 (N_1007,N_514,In_736);
and U1008 (N_1008,In_2988,In_840);
nor U1009 (N_1009,In_10,In_2672);
xor U1010 (N_1010,N_531,In_2851);
nor U1011 (N_1011,N_917,In_2811);
and U1012 (N_1012,In_1978,In_2664);
nor U1013 (N_1013,N_973,In_1713);
nand U1014 (N_1014,In_20,N_128);
xor U1015 (N_1015,N_743,In_3197);
nor U1016 (N_1016,In_3916,In_39);
xor U1017 (N_1017,In_1063,In_4719);
and U1018 (N_1018,In_2264,In_3039);
xnor U1019 (N_1019,In_975,In_2546);
nor U1020 (N_1020,In_3285,In_3021);
and U1021 (N_1021,In_3544,In_4834);
nand U1022 (N_1022,In_534,In_53);
nand U1023 (N_1023,In_4860,In_43);
and U1024 (N_1024,In_4338,In_4418);
and U1025 (N_1025,In_1056,In_139);
nor U1026 (N_1026,In_723,In_618);
and U1027 (N_1027,In_290,In_3410);
xnor U1028 (N_1028,In_1102,In_4815);
xor U1029 (N_1029,In_2154,In_3476);
nor U1030 (N_1030,In_3534,In_3820);
nand U1031 (N_1031,In_1804,In_787);
nor U1032 (N_1032,In_4516,In_2172);
nand U1033 (N_1033,In_3771,In_4764);
nand U1034 (N_1034,N_985,N_448);
or U1035 (N_1035,N_167,In_328);
nand U1036 (N_1036,In_936,In_1045);
and U1037 (N_1037,N_991,In_4907);
nor U1038 (N_1038,In_1601,N_579);
or U1039 (N_1039,In_797,N_979);
xnor U1040 (N_1040,In_1346,In_2390);
xor U1041 (N_1041,N_47,In_2430);
nor U1042 (N_1042,In_1635,N_272);
or U1043 (N_1043,In_4732,In_26);
nor U1044 (N_1044,In_1185,N_297);
or U1045 (N_1045,In_3446,In_3951);
or U1046 (N_1046,N_858,In_875);
xnor U1047 (N_1047,In_1241,In_4407);
nor U1048 (N_1048,In_739,In_239);
and U1049 (N_1049,N_992,N_663);
nand U1050 (N_1050,In_3457,N_932);
and U1051 (N_1051,In_194,In_1549);
xnor U1052 (N_1052,In_1224,In_1605);
xnor U1053 (N_1053,N_492,In_2678);
xor U1054 (N_1054,In_1162,In_2957);
nand U1055 (N_1055,In_2288,N_705);
or U1056 (N_1056,In_320,In_1808);
nor U1057 (N_1057,In_2932,In_2341);
xnor U1058 (N_1058,In_2278,In_3309);
xnor U1059 (N_1059,In_4135,In_4773);
nand U1060 (N_1060,In_2687,In_1481);
nor U1061 (N_1061,In_3841,In_2705);
xnor U1062 (N_1062,In_2304,In_3352);
nand U1063 (N_1063,In_2894,In_3389);
xnor U1064 (N_1064,In_271,N_689);
or U1065 (N_1065,In_309,N_210);
or U1066 (N_1066,N_717,In_1108);
nand U1067 (N_1067,In_2962,In_4612);
xor U1068 (N_1068,In_852,N_334);
or U1069 (N_1069,In_597,N_20);
and U1070 (N_1070,In_4271,N_767);
and U1071 (N_1071,N_729,In_4948);
xor U1072 (N_1072,In_693,In_821);
xnor U1073 (N_1073,In_762,In_2367);
nor U1074 (N_1074,In_1866,In_4149);
nor U1075 (N_1075,In_2622,In_4047);
nor U1076 (N_1076,In_2198,In_756);
nand U1077 (N_1077,In_3122,In_3952);
nand U1078 (N_1078,N_171,In_4762);
xnor U1079 (N_1079,In_3133,In_759);
nand U1080 (N_1080,In_1897,N_653);
and U1081 (N_1081,In_4539,In_377);
xnor U1082 (N_1082,In_3483,In_3694);
and U1083 (N_1083,In_2150,In_2094);
xnor U1084 (N_1084,In_3477,In_3568);
nand U1085 (N_1085,N_804,In_1120);
xor U1086 (N_1086,N_6,In_1254);
and U1087 (N_1087,In_2791,In_1546);
nand U1088 (N_1088,In_3855,In_3146);
nor U1089 (N_1089,In_458,In_352);
xor U1090 (N_1090,N_266,In_2438);
nor U1091 (N_1091,In_3390,In_2983);
nand U1092 (N_1092,In_4934,In_1517);
nor U1093 (N_1093,N_275,In_3236);
and U1094 (N_1094,In_4046,In_1304);
xor U1095 (N_1095,In_1386,In_411);
xor U1096 (N_1096,In_4557,In_4545);
nor U1097 (N_1097,N_987,N_924);
xor U1098 (N_1098,In_2534,In_1223);
xor U1099 (N_1099,In_957,In_363);
nor U1100 (N_1100,In_42,In_2620);
xnor U1101 (N_1101,N_530,N_542);
nand U1102 (N_1102,In_4077,In_4021);
or U1103 (N_1103,N_311,N_826);
xnor U1104 (N_1104,In_4200,In_4598);
xor U1105 (N_1105,In_2197,In_4641);
nor U1106 (N_1106,N_288,In_154);
nand U1107 (N_1107,N_422,In_4209);
xnor U1108 (N_1108,In_334,In_4501);
or U1109 (N_1109,In_2901,In_3252);
or U1110 (N_1110,N_913,In_914);
xor U1111 (N_1111,In_1761,In_1005);
nor U1112 (N_1112,N_322,N_669);
xnor U1113 (N_1113,In_2345,In_4993);
nor U1114 (N_1114,In_1654,In_2346);
or U1115 (N_1115,In_4289,In_2469);
nand U1116 (N_1116,In_171,In_1658);
and U1117 (N_1117,In_3192,In_4203);
nand U1118 (N_1118,N_834,In_1764);
xor U1119 (N_1119,N_562,N_258);
nand U1120 (N_1120,In_3172,In_1662);
and U1121 (N_1121,In_2812,In_941);
nor U1122 (N_1122,N_864,In_2924);
and U1123 (N_1123,In_65,In_253);
or U1124 (N_1124,In_1163,In_3941);
nand U1125 (N_1125,In_4657,In_4342);
nor U1126 (N_1126,N_491,In_1802);
xor U1127 (N_1127,In_134,In_51);
nor U1128 (N_1128,In_3073,In_4079);
nor U1129 (N_1129,In_3354,In_2716);
and U1130 (N_1130,In_2379,In_1512);
and U1131 (N_1131,In_4129,In_2239);
or U1132 (N_1132,In_4838,In_82);
and U1133 (N_1133,In_1651,In_1699);
xor U1134 (N_1134,In_3141,In_553);
nand U1135 (N_1135,In_3164,N_722);
nor U1136 (N_1136,In_1618,In_4897);
or U1137 (N_1137,N_898,In_285);
xor U1138 (N_1138,In_3509,In_4259);
or U1139 (N_1139,In_2885,In_4996);
and U1140 (N_1140,In_933,In_509);
and U1141 (N_1141,In_1550,In_2854);
nand U1142 (N_1142,N_935,In_3710);
xnor U1143 (N_1143,In_2875,In_3166);
nor U1144 (N_1144,In_1704,In_3008);
xor U1145 (N_1145,In_2482,In_4437);
xor U1146 (N_1146,In_166,In_4710);
and U1147 (N_1147,N_142,In_3560);
xnor U1148 (N_1148,In_413,In_1917);
nand U1149 (N_1149,In_1884,In_2652);
nand U1150 (N_1150,In_4107,In_812);
or U1151 (N_1151,In_1134,In_4631);
or U1152 (N_1152,In_777,N_733);
xnor U1153 (N_1153,In_4177,In_2281);
or U1154 (N_1154,In_3326,In_3957);
xor U1155 (N_1155,In_2884,In_3747);
nor U1156 (N_1156,N_377,In_3119);
xor U1157 (N_1157,In_935,In_2305);
and U1158 (N_1158,In_3972,In_3563);
and U1159 (N_1159,In_1981,In_4133);
nand U1160 (N_1160,In_439,In_1476);
and U1161 (N_1161,In_930,In_2010);
xor U1162 (N_1162,In_191,N_850);
xor U1163 (N_1163,In_4506,In_1267);
nor U1164 (N_1164,In_4094,In_2999);
or U1165 (N_1165,In_2723,In_2943);
and U1166 (N_1166,In_4874,In_3220);
nor U1167 (N_1167,In_4485,In_3128);
and U1168 (N_1168,N_83,In_4102);
xnor U1169 (N_1169,In_2365,N_849);
or U1170 (N_1170,In_4195,In_3167);
and U1171 (N_1171,In_141,In_1555);
or U1172 (N_1172,In_2069,In_4505);
nand U1173 (N_1173,In_1810,N_500);
or U1174 (N_1174,N_765,In_459);
nor U1175 (N_1175,N_965,N_890);
and U1176 (N_1176,In_3195,In_4366);
nor U1177 (N_1177,In_811,N_853);
or U1178 (N_1178,N_335,In_514);
nand U1179 (N_1179,In_3750,In_2226);
and U1180 (N_1180,In_4880,In_2800);
nor U1181 (N_1181,N_964,In_2271);
nand U1182 (N_1182,In_4926,In_29);
nor U1183 (N_1183,In_1343,In_1255);
xnor U1184 (N_1184,In_3051,In_283);
nor U1185 (N_1185,N_630,In_1288);
nor U1186 (N_1186,In_107,N_396);
nor U1187 (N_1187,N_468,In_1707);
xnor U1188 (N_1188,In_1904,In_566);
nor U1189 (N_1189,In_4313,In_581);
and U1190 (N_1190,N_242,In_3756);
nand U1191 (N_1191,In_1468,In_450);
and U1192 (N_1192,In_2334,In_1580);
xnor U1193 (N_1193,In_1779,In_4965);
nand U1194 (N_1194,In_2480,N_773);
xor U1195 (N_1195,In_1616,In_656);
or U1196 (N_1196,In_573,In_1535);
nor U1197 (N_1197,In_3442,In_4661);
and U1198 (N_1198,In_4925,In_3170);
xor U1199 (N_1199,In_4569,In_1748);
nand U1200 (N_1200,In_1257,In_2146);
nand U1201 (N_1201,In_2761,In_3597);
xor U1202 (N_1202,In_1385,In_829);
and U1203 (N_1203,N_474,N_952);
xnor U1204 (N_1204,In_3702,In_4453);
and U1205 (N_1205,In_4778,In_2429);
xor U1206 (N_1206,In_2422,N_715);
and U1207 (N_1207,In_257,In_456);
nor U1208 (N_1208,In_2084,In_1193);
nand U1209 (N_1209,In_84,N_672);
xnor U1210 (N_1210,N_434,N_988);
nand U1211 (N_1211,N_222,In_3587);
nor U1212 (N_1212,In_4871,N_433);
xor U1213 (N_1213,In_4464,N_943);
or U1214 (N_1214,In_2571,In_3660);
and U1215 (N_1215,In_1447,In_622);
xnor U1216 (N_1216,In_2767,In_240);
and U1217 (N_1217,In_2649,In_486);
and U1218 (N_1218,In_1547,In_1922);
xor U1219 (N_1219,In_748,In_2114);
and U1220 (N_1220,In_1548,In_3567);
nand U1221 (N_1221,In_3470,In_59);
xnor U1222 (N_1222,N_156,N_637);
and U1223 (N_1223,N_11,In_2882);
or U1224 (N_1224,In_360,In_3942);
nand U1225 (N_1225,In_2961,In_3207);
nor U1226 (N_1226,In_3006,N_437);
xnor U1227 (N_1227,N_844,N_8);
nand U1228 (N_1228,In_1598,In_1379);
xnor U1229 (N_1229,In_2301,In_1262);
or U1230 (N_1230,In_1997,N_10);
nor U1231 (N_1231,In_1935,In_215);
nand U1232 (N_1232,In_2566,N_68);
xnor U1233 (N_1233,In_4401,In_4832);
and U1234 (N_1234,In_152,In_1838);
nor U1235 (N_1235,N_501,In_4953);
xor U1236 (N_1236,N_771,N_384);
xor U1237 (N_1237,In_2133,In_2629);
or U1238 (N_1238,In_1087,N_803);
xor U1239 (N_1239,In_3593,In_36);
nor U1240 (N_1240,In_1062,N_993);
xor U1241 (N_1241,N_62,In_4474);
and U1242 (N_1242,In_1653,In_4186);
or U1243 (N_1243,In_172,In_3174);
or U1244 (N_1244,N_424,In_2493);
and U1245 (N_1245,In_1337,In_2306);
nand U1246 (N_1246,In_3546,In_69);
and U1247 (N_1247,In_2328,In_1159);
and U1248 (N_1248,In_3703,In_4264);
nor U1249 (N_1249,N_839,In_3435);
and U1250 (N_1250,In_2322,In_3539);
xnor U1251 (N_1251,In_1332,N_1091);
and U1252 (N_1252,In_4145,In_4406);
or U1253 (N_1253,In_3713,N_355);
and U1254 (N_1254,In_4577,In_3734);
xor U1255 (N_1255,N_788,In_2285);
and U1256 (N_1256,In_1879,In_2651);
and U1257 (N_1257,N_761,In_341);
nand U1258 (N_1258,In_2325,In_3281);
nor U1259 (N_1259,In_645,In_576);
xor U1260 (N_1260,In_1628,In_180);
nand U1261 (N_1261,N_1155,In_3906);
nor U1262 (N_1262,N_1012,In_4828);
nand U1263 (N_1263,In_1189,In_3603);
nand U1264 (N_1264,N_960,In_515);
and U1265 (N_1265,In_540,In_33);
or U1266 (N_1266,N_877,N_1045);
nor U1267 (N_1267,In_2439,In_3666);
nand U1268 (N_1268,In_2058,In_2617);
and U1269 (N_1269,In_1864,In_2848);
nand U1270 (N_1270,In_1932,In_3553);
nand U1271 (N_1271,N_1229,In_1239);
nand U1272 (N_1272,In_902,In_483);
xnor U1273 (N_1273,N_805,In_2644);
and U1274 (N_1274,In_524,In_329);
nand U1275 (N_1275,In_2972,In_157);
xnor U1276 (N_1276,N_1190,In_62);
nor U1277 (N_1277,In_690,In_299);
nor U1278 (N_1278,In_3867,In_3474);
nor U1279 (N_1279,In_3691,In_3783);
nand U1280 (N_1280,In_1081,In_671);
and U1281 (N_1281,In_3422,In_3933);
nand U1282 (N_1282,In_1188,In_854);
nor U1283 (N_1283,In_168,In_17);
nand U1284 (N_1284,N_900,In_4468);
or U1285 (N_1285,N_215,In_276);
nor U1286 (N_1286,In_4544,In_3034);
nor U1287 (N_1287,In_4964,In_1268);
and U1288 (N_1288,In_2003,In_2399);
or U1289 (N_1289,N_565,N_1079);
and U1290 (N_1290,N_1230,In_91);
and U1291 (N_1291,N_471,In_2420);
or U1292 (N_1292,N_751,N_723);
or U1293 (N_1293,N_1008,N_21);
nand U1294 (N_1294,In_4329,In_2398);
or U1295 (N_1295,N_1126,N_166);
nand U1296 (N_1296,In_322,In_3320);
and U1297 (N_1297,In_709,N_969);
nor U1298 (N_1298,In_1172,In_2159);
nor U1299 (N_1299,In_2568,N_90);
or U1300 (N_1300,N_921,N_887);
nor U1301 (N_1301,N_610,In_2487);
and U1302 (N_1302,In_4176,In_112);
or U1303 (N_1303,In_4456,In_3239);
nand U1304 (N_1304,In_2104,N_1047);
nand U1305 (N_1305,N_802,In_4770);
or U1306 (N_1306,In_851,In_2729);
and U1307 (N_1307,In_991,N_1169);
or U1308 (N_1308,In_2402,N_132);
nand U1309 (N_1309,In_3974,In_4220);
and U1310 (N_1310,N_230,N_696);
and U1311 (N_1311,N_1015,In_1411);
nand U1312 (N_1312,In_3960,N_902);
xor U1313 (N_1313,In_4512,In_1441);
or U1314 (N_1314,In_3753,In_4952);
nand U1315 (N_1315,In_2137,N_740);
or U1316 (N_1316,In_484,In_3938);
nand U1317 (N_1317,In_873,N_597);
xor U1318 (N_1318,In_4549,In_3993);
and U1319 (N_1319,N_300,N_270);
nand U1320 (N_1320,In_3721,In_831);
nand U1321 (N_1321,In_1503,In_809);
nor U1322 (N_1322,In_1093,In_4752);
nor U1323 (N_1323,N_69,In_2928);
or U1324 (N_1324,In_2495,In_4618);
xor U1325 (N_1325,In_4583,In_2613);
or U1326 (N_1326,In_1596,In_2413);
nand U1327 (N_1327,In_1910,In_4562);
nor U1328 (N_1328,N_823,In_2065);
xor U1329 (N_1329,N_226,In_3852);
nor U1330 (N_1330,In_70,In_2129);
and U1331 (N_1331,In_3144,In_2);
xor U1332 (N_1332,In_735,In_1991);
nor U1333 (N_1333,In_250,In_305);
and U1334 (N_1334,In_3872,N_374);
or U1335 (N_1335,N_435,N_571);
and U1336 (N_1336,In_600,In_704);
or U1337 (N_1337,In_342,In_843);
xnor U1338 (N_1338,In_2911,In_4286);
nor U1339 (N_1339,In_3520,N_23);
nand U1340 (N_1340,In_3507,N_1221);
nor U1341 (N_1341,In_3408,In_4166);
nor U1342 (N_1342,In_2189,N_368);
or U1343 (N_1343,N_152,In_643);
nand U1344 (N_1344,In_2453,N_681);
and U1345 (N_1345,N_1180,N_405);
or U1346 (N_1346,In_2047,In_3324);
nand U1347 (N_1347,In_126,In_4017);
nor U1348 (N_1348,In_1729,N_923);
xnor U1349 (N_1349,N_1065,In_758);
xor U1350 (N_1350,In_3282,N_1);
and U1351 (N_1351,In_57,In_3425);
nor U1352 (N_1352,N_1189,In_3455);
nand U1353 (N_1353,In_185,In_4971);
or U1354 (N_1354,In_3030,In_4410);
nand U1355 (N_1355,In_4330,N_1130);
nand U1356 (N_1356,In_1443,In_1356);
or U1357 (N_1357,N_810,N_1080);
nand U1358 (N_1358,In_4527,N_1205);
xnor U1359 (N_1359,In_1136,N_738);
nor U1360 (N_1360,N_1175,In_4181);
nor U1361 (N_1361,In_4357,N_67);
and U1362 (N_1362,In_1515,In_312);
and U1363 (N_1363,In_3158,N_457);
and U1364 (N_1364,N_587,In_1083);
nand U1365 (N_1365,In_2476,N_1236);
nand U1366 (N_1366,In_2272,In_1872);
nor U1367 (N_1367,In_265,N_414);
or U1368 (N_1368,N_1170,In_371);
or U1369 (N_1369,In_3581,In_333);
or U1370 (N_1370,In_877,In_4243);
and U1371 (N_1371,In_4352,In_1298);
or U1372 (N_1372,In_2982,In_1470);
nor U1373 (N_1373,In_2389,N_218);
xnor U1374 (N_1374,N_1123,N_238);
xor U1375 (N_1375,In_298,In_1514);
or U1376 (N_1376,In_1826,N_327);
xnor U1377 (N_1377,In_214,In_3313);
nor U1378 (N_1378,N_1004,In_1046);
or U1379 (N_1379,In_4790,In_4454);
nand U1380 (N_1380,In_1540,In_3749);
or U1381 (N_1381,In_3307,In_3704);
or U1382 (N_1382,N_698,In_2049);
xnor U1383 (N_1383,In_1946,In_2822);
or U1384 (N_1384,In_734,N_1244);
and U1385 (N_1385,In_3510,In_2423);
or U1386 (N_1386,In_841,In_4068);
or U1387 (N_1387,N_574,In_1625);
nor U1388 (N_1388,N_333,N_1002);
nor U1389 (N_1389,N_1203,In_512);
nand U1390 (N_1390,In_446,In_1966);
or U1391 (N_1391,In_415,In_2237);
xor U1392 (N_1392,In_4933,In_3272);
xor U1393 (N_1393,In_3755,In_3984);
or U1394 (N_1394,In_3498,N_1083);
nor U1395 (N_1395,N_63,In_3590);
xor U1396 (N_1396,In_2177,In_4402);
or U1397 (N_1397,In_4725,In_1688);
xnor U1398 (N_1398,In_1322,In_2880);
nand U1399 (N_1399,In_1738,In_306);
nor U1400 (N_1400,N_739,In_2841);
nor U1401 (N_1401,In_3806,In_1584);
nor U1402 (N_1402,N_665,In_3632);
or U1403 (N_1403,In_3400,In_4492);
or U1404 (N_1404,In_1251,N_736);
and U1405 (N_1405,N_248,In_2863);
and U1406 (N_1406,In_2441,In_2521);
and U1407 (N_1407,In_696,N_970);
nor U1408 (N_1408,In_920,N_247);
nor U1409 (N_1409,In_2156,In_4941);
and U1410 (N_1410,N_1089,N_329);
or U1411 (N_1411,In_1103,N_1024);
or U1412 (N_1412,In_4014,N_1210);
and U1413 (N_1413,In_718,In_3423);
or U1414 (N_1414,In_3890,In_386);
nand U1415 (N_1415,In_4430,In_3346);
and U1416 (N_1416,In_3640,In_3489);
or U1417 (N_1417,N_194,In_2019);
and U1418 (N_1418,In_2752,In_4600);
xnor U1419 (N_1419,In_800,In_4937);
and U1420 (N_1420,In_151,In_542);
nand U1421 (N_1421,In_2677,In_4792);
nor U1422 (N_1422,N_59,N_1149);
and U1423 (N_1423,N_1095,In_977);
nor U1424 (N_1424,In_887,In_3964);
or U1425 (N_1425,In_2260,In_3224);
nor U1426 (N_1426,In_4273,In_4344);
and U1427 (N_1427,N_957,In_3763);
nor U1428 (N_1428,In_3361,In_1834);
xor U1429 (N_1429,N_54,In_3392);
nor U1430 (N_1430,In_1819,In_677);
and U1431 (N_1431,In_2073,In_3958);
xor U1432 (N_1432,In_4580,In_1742);
nor U1433 (N_1433,In_3678,In_1606);
or U1434 (N_1434,N_550,In_144);
xor U1435 (N_1435,In_3071,In_2454);
nor U1436 (N_1436,N_661,In_4999);
nand U1437 (N_1437,In_2451,In_3966);
or U1438 (N_1438,In_2820,In_2085);
nand U1439 (N_1439,In_1949,In_1566);
nor U1440 (N_1440,In_2989,In_839);
nand U1441 (N_1441,In_805,In_2602);
xor U1442 (N_1442,In_3274,In_4753);
or U1443 (N_1443,In_4314,N_1103);
nor U1444 (N_1444,N_980,N_848);
nor U1445 (N_1445,N_510,N_833);
nor U1446 (N_1446,In_3559,N_1020);
xnor U1447 (N_1447,In_4666,In_4331);
nand U1448 (N_1448,In_4001,In_3157);
nand U1449 (N_1449,In_3350,In_4466);
xor U1450 (N_1450,In_4415,In_3242);
nor U1451 (N_1451,In_471,In_3875);
nor U1452 (N_1452,N_1238,In_4053);
or U1453 (N_1453,In_1407,In_3378);
and U1454 (N_1454,In_3064,In_3741);
nor U1455 (N_1455,In_4780,In_4267);
or U1456 (N_1456,In_210,In_1065);
nor U1457 (N_1457,N_596,In_3024);
xnor U1458 (N_1458,In_2840,In_1246);
and U1459 (N_1459,In_4742,In_2426);
nor U1460 (N_1460,In_3275,In_2319);
and U1461 (N_1461,N_547,In_1698);
nand U1462 (N_1462,In_2760,In_147);
or U1463 (N_1463,In_3333,N_642);
nor U1464 (N_1464,In_3738,In_3386);
xnor U1465 (N_1465,In_1827,In_4208);
xnor U1466 (N_1466,In_3019,In_2388);
and U1467 (N_1467,In_1287,In_2642);
xor U1468 (N_1468,In_4867,In_2669);
xor U1469 (N_1469,In_4814,In_4853);
xnor U1470 (N_1470,In_1725,In_1520);
or U1471 (N_1471,N_27,N_1062);
and U1472 (N_1472,In_3635,In_1647);
xor U1473 (N_1473,In_3267,In_8);
and U1474 (N_1474,In_2004,In_3462);
nor U1475 (N_1475,In_1315,N_315);
xnor U1476 (N_1476,In_24,In_1507);
nand U1477 (N_1477,In_3004,In_3919);
nor U1478 (N_1478,In_3634,N_1053);
nor U1479 (N_1479,In_3373,In_1726);
and U1480 (N_1480,In_1568,In_1424);
xnor U1481 (N_1481,In_746,In_2639);
and U1482 (N_1482,In_652,N_801);
nor U1483 (N_1483,In_2748,In_2232);
or U1484 (N_1484,In_4877,In_4033);
or U1485 (N_1485,N_382,N_927);
and U1486 (N_1486,N_198,In_2223);
nor U1487 (N_1487,In_1595,In_327);
and U1488 (N_1488,In_4682,In_383);
nand U1489 (N_1489,In_2918,In_1961);
and U1490 (N_1490,In_755,N_1016);
and U1491 (N_1491,In_2676,In_3873);
xor U1492 (N_1492,In_1455,N_560);
xnor U1493 (N_1493,In_1123,In_2786);
or U1494 (N_1494,In_863,In_3118);
nor U1495 (N_1495,In_2828,N_1014);
and U1496 (N_1496,In_3910,In_3347);
or U1497 (N_1497,N_1140,N_1066);
nor U1498 (N_1498,In_279,In_1059);
xnor U1499 (N_1499,In_3475,In_4348);
and U1500 (N_1500,N_651,In_3306);
and U1501 (N_1501,In_3804,N_1419);
xnor U1502 (N_1502,N_325,In_1316);
or U1503 (N_1503,In_4509,In_1617);
nand U1504 (N_1504,In_2658,In_4349);
nor U1505 (N_1505,N_139,In_491);
xnor U1506 (N_1506,In_3896,In_1452);
nand U1507 (N_1507,In_3676,In_3454);
nand U1508 (N_1508,In_2152,N_1165);
or U1509 (N_1509,N_1447,In_3903);
nand U1510 (N_1510,In_3968,N_1057);
and U1511 (N_1511,N_726,In_4628);
or U1512 (N_1512,In_2888,In_4998);
nand U1513 (N_1513,N_861,In_98);
or U1514 (N_1514,N_1334,In_2404);
nor U1515 (N_1515,In_963,N_241);
xor U1516 (N_1516,In_4127,In_3682);
nand U1517 (N_1517,In_2254,In_684);
or U1518 (N_1518,In_3049,In_2075);
nor U1519 (N_1519,In_1723,In_4445);
nor U1520 (N_1520,In_4555,In_1513);
nor U1521 (N_1521,N_1078,In_1668);
nor U1522 (N_1522,In_1390,N_1036);
xor U1523 (N_1523,N_221,In_4448);
and U1524 (N_1524,In_1972,In_3328);
nor U1525 (N_1525,In_4004,In_4625);
or U1526 (N_1526,N_670,N_1255);
and U1527 (N_1527,N_878,N_191);
nor U1528 (N_1528,In_757,N_752);
nand U1529 (N_1529,In_1119,N_977);
nor U1530 (N_1530,In_2279,In_1860);
nor U1531 (N_1531,N_1382,In_3602);
and U1532 (N_1532,In_4768,In_2771);
nand U1533 (N_1533,In_3848,N_421);
or U1534 (N_1534,In_1115,In_4182);
or U1535 (N_1535,N_944,In_4252);
or U1536 (N_1536,In_1311,In_3147);
or U1537 (N_1537,In_4489,In_955);
and U1538 (N_1538,In_3670,In_3493);
or U1539 (N_1539,N_220,N_344);
or U1540 (N_1540,N_1461,In_2557);
nand U1541 (N_1541,In_3074,N_107);
nor U1542 (N_1542,In_2131,In_1717);
or U1543 (N_1543,In_1373,N_89);
and U1544 (N_1544,N_785,N_182);
or U1545 (N_1545,In_2138,In_2843);
or U1546 (N_1546,N_527,In_2670);
xnor U1547 (N_1547,In_1030,In_3839);
nor U1548 (N_1548,In_4694,In_1769);
and U1549 (N_1549,In_405,In_1576);
or U1550 (N_1550,In_3936,N_1195);
nand U1551 (N_1551,In_1684,N_832);
or U1552 (N_1552,In_2433,In_2140);
nor U1553 (N_1553,In_3518,In_2993);
and U1554 (N_1554,In_1006,In_4579);
or U1555 (N_1555,In_4684,In_978);
or U1556 (N_1556,In_4850,N_307);
xnor U1557 (N_1557,In_2504,In_527);
nor U1558 (N_1558,N_1116,In_3314);
or U1559 (N_1559,In_121,In_3471);
nand U1560 (N_1560,In_900,In_1675);
or U1561 (N_1561,In_2971,In_1336);
nor U1562 (N_1562,N_359,In_4335);
nor U1563 (N_1563,In_4006,In_3447);
or U1564 (N_1564,In_246,In_2638);
or U1565 (N_1565,In_2648,In_945);
xnor U1566 (N_1566,In_2016,In_343);
nand U1567 (N_1567,In_2242,In_4823);
xor U1568 (N_1568,In_4910,In_3623);
nand U1569 (N_1569,N_1499,In_3182);
nand U1570 (N_1570,In_549,N_1496);
nand U1571 (N_1571,In_1002,In_4157);
and U1572 (N_1572,In_3225,In_3017);
and U1573 (N_1573,N_549,In_2641);
or U1574 (N_1574,In_1230,N_1157);
nand U1575 (N_1575,In_4587,In_1928);
nor U1576 (N_1576,In_3348,N_1411);
nor U1577 (N_1577,N_896,N_1154);
nor U1578 (N_1578,In_2675,In_2121);
and U1579 (N_1579,In_4275,In_1283);
xor U1580 (N_1580,N_1456,In_1191);
nand U1581 (N_1581,N_954,N_606);
nand U1582 (N_1582,In_212,N_1403);
nand U1583 (N_1583,N_1405,In_1793);
nor U1584 (N_1584,N_600,In_1638);
nor U1585 (N_1585,In_1197,In_4038);
and U1586 (N_1586,N_1119,N_118);
nor U1587 (N_1587,N_1213,In_4532);
and U1588 (N_1588,N_691,In_685);
nand U1589 (N_1589,In_4118,In_3218);
xor U1590 (N_1590,In_1526,In_879);
xor U1591 (N_1591,In_339,N_504);
or U1592 (N_1592,In_4442,N_404);
nand U1593 (N_1593,N_862,In_1055);
xnor U1594 (N_1594,In_2149,In_2207);
nor U1595 (N_1595,In_3674,N_40);
xnor U1596 (N_1596,In_3221,In_269);
nand U1597 (N_1597,In_1771,In_1296);
nor U1598 (N_1598,N_1445,N_431);
or U1599 (N_1599,In_3255,In_4404);
nand U1600 (N_1600,In_2635,N_487);
nor U1601 (N_1601,In_2688,In_188);
nor U1602 (N_1602,In_2816,In_3642);
or U1603 (N_1603,In_4059,In_567);
nor U1604 (N_1604,N_999,In_4915);
nor U1605 (N_1605,In_4196,In_417);
nand U1606 (N_1606,In_1795,N_918);
and U1607 (N_1607,N_1168,N_1058);
or U1608 (N_1608,N_257,In_3801);
xnor U1609 (N_1609,In_1475,N_830);
xnor U1610 (N_1610,In_2066,In_3169);
nand U1611 (N_1611,In_799,N_85);
and U1612 (N_1612,In_2603,N_113);
xnor U1613 (N_1613,N_817,N_1090);
and U1614 (N_1614,N_1311,In_1276);
and U1615 (N_1615,In_263,In_4173);
or U1616 (N_1616,In_2944,N_1162);
nand U1617 (N_1617,In_2674,In_909);
nand U1618 (N_1618,In_145,N_43);
or U1619 (N_1619,In_2021,N_1263);
nor U1620 (N_1620,In_38,In_2373);
nor U1621 (N_1621,In_3340,In_130);
xor U1622 (N_1622,In_4447,N_253);
and U1623 (N_1623,N_706,N_1148);
nor U1624 (N_1624,In_3986,In_4146);
xnor U1625 (N_1625,In_2684,In_1355);
nand U1626 (N_1626,In_1367,In_791);
nor U1627 (N_1627,In_3283,N_626);
or U1628 (N_1628,N_1344,N_1067);
and U1629 (N_1629,In_3230,In_1433);
nand U1630 (N_1630,In_32,N_455);
nand U1631 (N_1631,In_4069,N_966);
nand U1632 (N_1632,In_3662,N_388);
or U1633 (N_1633,In_782,N_1144);
nand U1634 (N_1634,In_289,In_1847);
xnor U1635 (N_1635,N_1425,In_2088);
nand U1636 (N_1636,N_1495,In_1933);
and U1637 (N_1637,In_3973,In_2359);
nor U1638 (N_1638,In_4427,In_2372);
xnor U1639 (N_1639,In_3486,In_1829);
and U1640 (N_1640,In_3183,In_1167);
nor U1641 (N_1641,N_1034,N_685);
and U1642 (N_1642,In_2462,In_4970);
or U1643 (N_1643,In_4507,In_2703);
nand U1644 (N_1644,In_4966,In_2326);
and U1645 (N_1645,In_3411,In_4632);
xnor U1646 (N_1646,In_4306,In_3813);
xnor U1647 (N_1647,In_2871,In_3380);
and U1648 (N_1648,In_101,N_989);
nand U1649 (N_1649,N_1237,N_1044);
or U1650 (N_1650,In_2356,In_1942);
xnor U1651 (N_1651,N_631,In_3961);
and U1652 (N_1652,In_3406,In_2411);
nand U1653 (N_1653,In_4734,In_1426);
and U1654 (N_1654,N_1356,N_1454);
xnor U1655 (N_1655,In_2734,N_423);
nor U1656 (N_1656,N_323,In_4708);
xnor U1657 (N_1657,N_1262,N_508);
nand U1658 (N_1658,N_950,N_1026);
and U1659 (N_1659,In_1210,In_2194);
or U1660 (N_1660,In_1014,In_1552);
or U1661 (N_1661,In_4165,In_3184);
xor U1662 (N_1662,In_1464,In_1541);
nor U1663 (N_1663,In_3087,In_4830);
or U1664 (N_1664,In_4659,In_3327);
and U1665 (N_1665,N_1005,N_779);
and U1666 (N_1666,N_912,In_202);
xor U1667 (N_1667,In_1645,In_4422);
xnor U1668 (N_1668,N_121,In_4315);
or U1669 (N_1669,In_2519,In_4362);
or U1670 (N_1670,In_2542,In_2711);
or U1671 (N_1671,N_1436,In_1817);
nor U1672 (N_1672,In_4514,N_1231);
nand U1673 (N_1673,In_3254,N_1192);
and U1674 (N_1674,In_3746,In_4443);
and U1675 (N_1675,N_737,In_4795);
nor U1676 (N_1676,In_408,N_1291);
xor U1677 (N_1677,In_1274,In_3037);
nor U1678 (N_1678,N_1097,In_1768);
xor U1679 (N_1679,In_675,N_941);
xor U1680 (N_1680,In_2842,In_272);
nor U1681 (N_1681,N_614,In_186);
and U1682 (N_1682,In_1273,In_2312);
or U1683 (N_1683,In_3213,N_741);
nand U1684 (N_1684,In_2265,In_1921);
or U1685 (N_1685,In_4184,In_3175);
or U1686 (N_1686,In_3665,N_1471);
or U1687 (N_1687,In_1674,In_2581);
nor U1688 (N_1688,N_1212,In_117);
nand U1689 (N_1689,In_4749,In_822);
nand U1690 (N_1690,In_3712,In_1573);
nand U1691 (N_1691,In_4119,In_666);
xor U1692 (N_1692,N_1353,In_2349);
nand U1693 (N_1693,N_1077,In_2415);
xnor U1694 (N_1694,N_281,In_3200);
nor U1695 (N_1695,In_698,In_3069);
nor U1696 (N_1696,N_584,N_541);
or U1697 (N_1697,N_1117,N_1393);
nand U1698 (N_1698,N_1040,In_2450);
nand U1699 (N_1699,N_478,In_3088);
or U1700 (N_1700,N_22,In_4678);
nand U1701 (N_1701,In_1489,In_4908);
or U1702 (N_1702,In_3830,In_3866);
or U1703 (N_1703,In_50,In_1019);
or U1704 (N_1704,In_771,N_1396);
nor U1705 (N_1705,In_1874,In_3402);
xor U1706 (N_1706,In_3886,N_951);
or U1707 (N_1707,N_330,In_3802);
xnor U1708 (N_1708,In_3294,In_3773);
and U1709 (N_1709,N_197,In_2432);
nand U1710 (N_1710,In_2781,In_1218);
or U1711 (N_1711,In_2736,In_750);
or U1712 (N_1712,In_3894,In_4781);
or U1713 (N_1713,N_595,In_4892);
or U1714 (N_1714,In_3311,In_423);
nor U1715 (N_1715,In_2337,In_2160);
xnor U1716 (N_1716,In_2077,In_1248);
xnor U1717 (N_1717,N_1215,In_2586);
and U1718 (N_1718,In_892,In_4191);
xor U1719 (N_1719,N_910,N_639);
or U1720 (N_1720,In_1728,N_809);
nand U1721 (N_1721,In_2973,In_3011);
and U1722 (N_1722,In_3708,In_4777);
or U1723 (N_1723,N_240,In_1679);
xnor U1724 (N_1724,In_4729,In_4767);
and U1725 (N_1725,N_36,In_2565);
and U1726 (N_1726,In_1569,In_1097);
nor U1727 (N_1727,In_691,N_1030);
nand U1728 (N_1728,In_301,In_4613);
nor U1729 (N_1729,N_254,In_55);
nand U1730 (N_1730,In_2374,In_3917);
nor U1731 (N_1731,In_4193,N_612);
or U1732 (N_1732,In_780,N_1071);
nor U1733 (N_1733,In_426,N_872);
and U1734 (N_1734,In_2981,N_1374);
nand U1735 (N_1735,In_921,N_1093);
and U1736 (N_1736,In_2726,In_2823);
nor U1737 (N_1737,In_4621,N_1171);
nor U1738 (N_1738,In_4548,In_2589);
and U1739 (N_1739,In_4683,N_851);
xnor U1740 (N_1740,In_2769,In_1285);
xor U1741 (N_1741,N_1270,N_1105);
or U1742 (N_1742,In_687,N_608);
or U1743 (N_1743,N_1272,In_1590);
or U1744 (N_1744,N_1328,In_2261);
nand U1745 (N_1745,N_1308,In_3684);
and U1746 (N_1746,N_1049,In_4198);
nand U1747 (N_1747,In_979,In_1995);
xor U1748 (N_1748,In_3654,N_1414);
or U1749 (N_1749,In_1445,N_974);
or U1750 (N_1750,In_4390,N_1223);
nor U1751 (N_1751,In_1660,In_4219);
xor U1752 (N_1752,In_3980,In_3716);
xor U1753 (N_1753,In_133,N_981);
nor U1754 (N_1754,In_4761,In_910);
and U1755 (N_1755,In_3645,In_3154);
nand U1756 (N_1756,N_1439,N_903);
or U1757 (N_1757,In_544,In_2467);
or U1758 (N_1758,N_1545,In_774);
and U1759 (N_1759,In_1610,In_287);
xnor U1760 (N_1760,N_889,N_1299);
nor U1761 (N_1761,In_2553,N_1665);
and U1762 (N_1762,In_2384,In_749);
or U1763 (N_1763,In_3606,N_1675);
xor U1764 (N_1764,In_3611,In_3082);
and U1765 (N_1765,N_1068,N_1387);
xnor U1766 (N_1766,In_2912,In_3977);
or U1767 (N_1767,N_381,In_3599);
and U1768 (N_1768,In_1722,In_195);
nand U1769 (N_1769,In_1971,N_690);
or U1770 (N_1770,In_4518,In_4197);
nor U1771 (N_1771,In_2196,In_4959);
nor U1772 (N_1772,In_1217,In_538);
nor U1773 (N_1773,N_1410,N_794);
or U1774 (N_1774,N_971,N_1562);
and U1775 (N_1775,N_1584,In_2995);
nor U1776 (N_1776,In_4066,N_1709);
nand U1777 (N_1777,In_2659,N_1715);
nor U1778 (N_1778,N_578,In_1359);
and U1779 (N_1779,N_1585,N_886);
nand U1780 (N_1780,N_1194,In_594);
or U1781 (N_1781,N_267,In_3151);
xnor U1782 (N_1782,In_4772,N_1197);
nor U1783 (N_1783,In_4384,In_1074);
nand U1784 (N_1784,N_959,In_243);
nor U1785 (N_1785,N_1300,In_4123);
nand U1786 (N_1786,In_2358,N_648);
nand U1787 (N_1787,In_686,In_460);
xnor U1788 (N_1788,In_4513,In_3838);
or U1789 (N_1789,In_2921,N_1616);
xnor U1790 (N_1790,In_541,In_1644);
nand U1791 (N_1791,In_90,N_1399);
nand U1792 (N_1792,N_793,In_1425);
xnor U1793 (N_1793,In_4091,N_708);
and U1794 (N_1794,In_3517,N_526);
nand U1795 (N_1795,In_4885,N_680);
nand U1796 (N_1796,N_576,In_3203);
xor U1797 (N_1797,In_1429,In_2579);
nor U1798 (N_1798,N_1293,N_486);
xnor U1799 (N_1799,N_1697,N_1572);
nand U1800 (N_1800,In_4546,In_2101);
nor U1801 (N_1801,In_3367,N_1503);
xnor U1802 (N_1802,N_515,In_2930);
nor U1803 (N_1803,In_4039,N_1422);
or U1804 (N_1804,N_1246,N_1397);
or U1805 (N_1805,In_2577,In_4696);
xor U1806 (N_1806,In_2083,In_4444);
nand U1807 (N_1807,In_3393,In_4706);
nor U1808 (N_1808,N_819,In_3982);
nand U1809 (N_1809,In_2031,In_4327);
xnor U1810 (N_1810,In_3260,In_1673);
nor U1811 (N_1811,N_524,In_1594);
xnor U1812 (N_1812,In_3020,N_1133);
or U1813 (N_1813,In_3849,In_1275);
xnor U1814 (N_1814,In_4089,N_905);
or U1815 (N_1815,In_4643,N_106);
xor U1816 (N_1816,In_1794,In_4341);
and U1817 (N_1817,In_3028,In_670);
nand U1818 (N_1818,N_204,In_1395);
nand U1819 (N_1819,In_1036,N_569);
nand U1820 (N_1820,In_3160,In_165);
nor U1821 (N_1821,In_3816,N_1482);
xnor U1822 (N_1822,In_3472,In_4229);
nand U1823 (N_1823,N_1658,In_4504);
nand U1824 (N_1824,In_2858,N_763);
nand U1825 (N_1825,In_4318,In_3371);
xnor U1826 (N_1826,In_2252,In_1868);
nand U1827 (N_1827,In_3343,In_1811);
and U1828 (N_1828,N_265,N_545);
nand U1829 (N_1829,In_3460,In_3098);
nand U1830 (N_1830,N_444,N_528);
and U1831 (N_1831,In_3880,In_2270);
nor U1832 (N_1832,In_3251,In_4029);
xor U1833 (N_1833,N_789,In_4757);
and U1834 (N_1834,In_4050,In_2168);
nor U1835 (N_1835,N_473,In_1016);
xnor U1836 (N_1836,N_522,N_386);
nand U1837 (N_1837,In_2528,In_474);
or U1838 (N_1838,In_653,In_4340);
or U1839 (N_1839,In_3461,In_2103);
xor U1840 (N_1840,In_2780,In_1232);
or U1841 (N_1841,In_4483,In_2623);
nor U1842 (N_1842,In_1880,In_726);
and U1843 (N_1843,In_768,In_1009);
nor U1844 (N_1844,In_2803,In_878);
xor U1845 (N_1845,In_2262,In_1486);
nand U1846 (N_1846,In_4421,In_522);
or U1847 (N_1847,In_4520,In_369);
or U1848 (N_1848,In_4705,N_911);
nor U1849 (N_1849,In_4398,N_1181);
nand U1850 (N_1850,In_4856,In_2588);
and U1851 (N_1851,In_2845,In_1672);
and U1852 (N_1852,In_1131,In_2141);
nand U1853 (N_1853,N_1383,In_412);
nand U1854 (N_1854,In_3444,N_1570);
or U1855 (N_1855,In_1848,N_1009);
nor U1856 (N_1856,In_1905,In_2667);
and U1857 (N_1857,In_420,N_556);
nand U1858 (N_1858,In_489,N_268);
or U1859 (N_1859,In_4904,In_4126);
and U1860 (N_1860,In_546,In_1842);
and U1861 (N_1861,In_954,N_1398);
or U1862 (N_1862,In_4847,N_1085);
xnor U1863 (N_1863,In_1394,N_1714);
or U1864 (N_1864,In_2599,In_75);
and U1865 (N_1865,N_713,In_4722);
nand U1866 (N_1866,In_2970,In_946);
nand U1867 (N_1867,N_1476,In_4852);
and U1868 (N_1868,N_582,N_1727);
or U1869 (N_1869,In_1295,In_3579);
nand U1870 (N_1870,N_936,In_2042);
and U1871 (N_1871,N_1618,In_3304);
nand U1872 (N_1872,In_3557,In_3077);
or U1873 (N_1873,N_1199,In_2721);
nor U1874 (N_1874,N_914,N_990);
nand U1875 (N_1875,In_586,In_865);
nand U1876 (N_1876,In_2491,N_49);
nand U1877 (N_1877,In_899,N_1266);
and U1878 (N_1878,In_1639,In_3994);
xnor U1879 (N_1879,In_2744,In_4949);
nand U1880 (N_1880,In_3789,N_1276);
nor U1881 (N_1881,N_1274,N_1651);
nor U1882 (N_1882,In_2475,In_241);
and U1883 (N_1883,In_1950,In_3976);
nand U1884 (N_1884,N_469,N_1687);
nor U1885 (N_1885,N_1707,N_1265);
nor U1886 (N_1886,N_638,N_1031);
or U1887 (N_1887,N_1725,In_4086);
xor U1888 (N_1888,In_1451,In_4496);
nor U1889 (N_1889,In_1563,N_1186);
or U1890 (N_1890,In_3810,N_502);
or U1891 (N_1891,N_939,In_4081);
nor U1892 (N_1892,In_2215,In_3463);
xor U1893 (N_1893,N_784,N_347);
xnor U1894 (N_1894,N_813,In_4462);
or U1895 (N_1895,In_3120,N_758);
nor U1896 (N_1896,In_4981,N_402);
and U1897 (N_1897,In_4281,N_728);
or U1898 (N_1898,In_2540,In_2486);
and U1899 (N_1899,In_2611,N_676);
xor U1900 (N_1900,In_366,In_3308);
and U1901 (N_1901,In_1504,N_829);
and U1902 (N_1902,N_369,N_46);
xnor U1903 (N_1903,N_778,N_800);
and U1904 (N_1904,In_4005,In_4351);
nand U1905 (N_1905,In_4865,In_3190);
xnor U1906 (N_1906,In_849,In_4775);
nor U1907 (N_1907,In_857,In_2370);
and U1908 (N_1908,In_1720,N_1370);
nand U1909 (N_1909,In_3908,In_925);
xor U1910 (N_1910,In_4640,In_3911);
nand U1911 (N_1911,N_1094,In_4253);
xor U1912 (N_1912,In_67,N_1098);
xnor U1913 (N_1913,In_510,N_1735);
nand U1914 (N_1914,N_1525,In_552);
and U1915 (N_1915,In_3540,N_1217);
or U1916 (N_1916,N_79,In_2210);
xnor U1917 (N_1917,N_60,N_1591);
nand U1918 (N_1918,In_3882,In_162);
nor U1919 (N_1919,N_843,N_899);
nor U1920 (N_1920,N_1376,In_1146);
or U1921 (N_1921,N_1690,N_1558);
nand U1922 (N_1922,In_2600,N_1463);
xnor U1923 (N_1923,N_1710,N_1354);
nand U1924 (N_1924,In_2992,N_1599);
xor U1925 (N_1925,In_2994,In_3372);
xor U1926 (N_1926,In_3707,In_4459);
xnor U1927 (N_1927,N_1460,N_1373);
xnor U1928 (N_1928,In_3901,N_189);
nor U1929 (N_1929,In_1996,N_299);
xor U1930 (N_1930,N_534,N_148);
or U1931 (N_1931,N_1379,N_296);
nand U1932 (N_1932,In_3636,N_1109);
xnor U1933 (N_1933,In_721,In_1701);
nor U1934 (N_1934,In_2030,N_1081);
and U1935 (N_1935,In_4431,In_4397);
nor U1936 (N_1936,N_82,In_3136);
and U1937 (N_1937,In_3438,N_1590);
and U1938 (N_1938,In_2052,N_1375);
nor U1939 (N_1939,N_1135,In_4368);
xor U1940 (N_1940,In_4699,N_1717);
xor U1941 (N_1941,In_3827,In_3403);
nand U1942 (N_1942,In_965,In_3258);
and U1943 (N_1943,N_1084,In_3018);
nor U1944 (N_1944,In_3436,In_1157);
nor U1945 (N_1945,N_249,In_393);
nor U1946 (N_1946,In_419,N_412);
xor U1947 (N_1947,In_1821,N_1337);
and U1948 (N_1948,In_4192,N_1347);
and U1949 (N_1949,N_217,In_4843);
or U1950 (N_1950,In_80,In_754);
xor U1951 (N_1951,N_1209,In_2022);
nand U1952 (N_1952,In_2886,N_370);
nor U1953 (N_1953,In_1222,In_1587);
nand U1954 (N_1954,N_92,N_1575);
or U1955 (N_1955,N_1358,In_1623);
and U1956 (N_1956,In_498,N_1193);
and U1957 (N_1957,In_2712,In_1366);
and U1958 (N_1958,N_1256,N_1106);
xnor U1959 (N_1959,N_42,In_3626);
xnor U1960 (N_1960,In_4417,N_787);
nand U1961 (N_1961,In_4097,In_2940);
nor U1962 (N_1962,In_1435,In_1358);
or U1963 (N_1963,In_3199,In_1607);
or U1964 (N_1964,N_411,In_1208);
nor U1965 (N_1965,In_4337,N_543);
xnor U1966 (N_1966,In_3341,N_926);
nand U1967 (N_1967,N_1164,N_827);
or U1968 (N_1968,N_1019,In_418);
xor U1969 (N_1969,N_187,N_143);
and U1970 (N_1970,In_1718,N_346);
xnor U1971 (N_1971,In_4018,In_2701);
nand U1972 (N_1972,In_3316,In_4658);
and U1973 (N_1973,N_797,In_2091);
xor U1974 (N_1974,In_1629,In_3533);
or U1975 (N_1975,N_1747,In_2859);
xor U1976 (N_1976,In_4201,In_1686);
or U1977 (N_1977,N_1200,In_1604);
nor U1978 (N_1978,N_282,In_30);
or U1979 (N_1979,In_2619,In_2980);
or U1980 (N_1980,In_4238,In_3458);
nand U1981 (N_1981,In_4093,In_2231);
nor U1982 (N_1982,In_3111,N_1407);
or U1983 (N_1983,N_206,In_2417);
xnor U1984 (N_1984,In_1109,In_4714);
xnor U1985 (N_1985,In_4226,In_4168);
nor U1986 (N_1986,N_1671,In_3420);
xnor U1987 (N_1987,N_466,In_828);
nor U1988 (N_1988,N_1208,N_592);
xnor U1989 (N_1989,In_2250,N_53);
nand U1990 (N_1990,In_52,In_3576);
xor U1991 (N_1991,N_1153,In_593);
or U1992 (N_1992,In_2634,N_1151);
xor U1993 (N_1993,In_4142,In_3059);
nor U1994 (N_1994,N_192,In_2452);
and U1995 (N_1995,N_1338,In_548);
xnor U1996 (N_1996,In_1448,N_1533);
xor U1997 (N_1997,N_1325,In_3355);
nor U1998 (N_1998,N_506,In_1207);
xor U1999 (N_1999,In_1228,In_3002);
and U2000 (N_2000,N_1556,In_444);
nand U2001 (N_2001,In_280,N_1657);
and U2002 (N_2002,In_861,In_4224);
xnor U2003 (N_2003,N_757,In_1670);
and U2004 (N_2004,N_291,In_4609);
and U2005 (N_2005,N_1784,N_385);
nor U2006 (N_2006,In_1348,In_4839);
xnor U2007 (N_2007,N_869,In_4020);
nor U2008 (N_2008,N_1909,N_1513);
and U2009 (N_2009,N_460,In_1427);
nand U2010 (N_2010,N_1537,In_4140);
xnor U2011 (N_2011,In_3290,N_702);
and U2012 (N_2012,In_2754,In_4234);
xnor U2013 (N_2013,N_138,N_1510);
xor U2014 (N_2014,N_536,N_721);
or U2015 (N_2015,N_336,In_4128);
xor U2016 (N_2016,N_593,In_3315);
nand U2017 (N_2017,In_1457,N_821);
and U2018 (N_2018,N_1978,N_1142);
and U2019 (N_2019,In_4369,N_1369);
xnor U2020 (N_2020,N_1452,N_679);
and U2021 (N_2021,In_2234,In_609);
nor U2022 (N_2022,In_2904,In_4936);
and U2023 (N_2023,N_1435,N_1225);
nor U2024 (N_2024,N_1803,In_4343);
xor U2025 (N_2025,N_1933,N_1490);
or U2026 (N_2026,In_937,In_4138);
xor U2027 (N_2027,N_1638,N_1640);
xnor U2028 (N_2028,In_1225,N_1486);
or U2029 (N_2029,N_1625,In_4387);
or U2030 (N_2030,In_1289,N_1125);
xnor U2031 (N_2031,In_885,In_237);
or U2032 (N_2032,In_2621,N_1879);
nor U2033 (N_2033,In_485,N_1839);
nor U2034 (N_2034,In_4672,N_856);
and U2035 (N_2035,In_4319,N_1881);
xor U2036 (N_2036,N_1206,In_630);
or U2037 (N_2037,In_2318,In_2708);
or U2038 (N_2038,N_383,N_831);
and U2039 (N_2039,In_1323,In_3431);
nor U2040 (N_2040,N_1010,In_4071);
and U2041 (N_2041,In_4912,N_1131);
nand U2042 (N_2042,N_678,In_1126);
nor U2043 (N_2043,N_1674,In_4435);
or U2044 (N_2044,In_2353,In_3445);
or U2045 (N_2045,In_3748,In_694);
nor U2046 (N_2046,In_4232,N_727);
xor U2047 (N_2047,In_2128,In_4451);
nor U2048 (N_2048,N_774,In_1463);
nand U2049 (N_2049,In_992,In_1498);
xor U2050 (N_2050,N_1035,N_1548);
xnor U2051 (N_2051,In_2257,N_688);
nand U2052 (N_2052,N_475,N_1767);
and U2053 (N_2053,In_2018,In_1797);
or U2054 (N_2054,In_1301,In_3680);
and U2055 (N_2055,In_947,In_588);
xnor U2056 (N_2056,In_587,N_1327);
or U2057 (N_2057,In_4298,In_2447);
and U2058 (N_2058,N_1457,In_1666);
xnor U2059 (N_2059,In_4076,N_1348);
xnor U2060 (N_2060,N_358,In_4671);
or U2061 (N_2061,In_2435,In_1782);
xor U2062 (N_2062,N_1477,In_4358);
xnor U2063 (N_2063,In_1434,N_1874);
and U2064 (N_2064,In_4711,In_3302);
or U2065 (N_2065,In_3066,In_4124);
xnor U2066 (N_2066,In_763,In_3808);
nand U2067 (N_2067,In_1330,In_626);
or U2068 (N_2068,In_1458,In_810);
nand U2069 (N_2069,In_737,In_4350);
nand U2070 (N_2070,In_1001,In_1033);
and U2071 (N_2071,N_1267,N_643);
or U2072 (N_2072,N_1574,N_513);
nand U2073 (N_2073,In_3732,In_2852);
xnor U2074 (N_2074,N_897,In_717);
xnor U2075 (N_2075,In_1641,In_2909);
nor U2076 (N_2076,In_3266,In_533);
nor U2077 (N_2077,In_872,In_5);
nand U2078 (N_2078,N_1588,In_3273);
or U2079 (N_2079,In_4499,N_1003);
nor U2080 (N_2080,N_1386,In_3845);
and U2081 (N_2081,N_1566,In_520);
nor U2082 (N_2082,N_1807,In_4174);
or U2083 (N_2083,In_1124,In_1318);
or U2084 (N_2084,In_4395,In_3003);
xor U2085 (N_2085,In_1307,N_1770);
nand U2086 (N_2086,In_3428,N_419);
xor U2087 (N_2087,N_764,N_1762);
and U2088 (N_2088,In_3222,N_1688);
nor U2089 (N_2089,N_867,In_4231);
or U2090 (N_2090,N_623,In_2561);
nor U2091 (N_2091,N_629,N_1517);
xor U2092 (N_2092,In_4756,N_931);
nand U2093 (N_2093,In_571,N_1972);
and U2094 (N_2094,In_4813,In_3289);
nand U2095 (N_2095,In_1020,In_1021);
xnor U2096 (N_2096,N_1777,In_2607);
or U2097 (N_2097,In_1948,N_462);
nor U2098 (N_2098,In_2977,N_1516);
and U2099 (N_2099,N_196,In_1799);
and U2100 (N_2100,In_2109,N_1760);
nor U2101 (N_2101,N_1772,In_627);
and U2102 (N_2102,In_1837,N_1870);
xnor U2103 (N_2103,N_1876,In_1353);
xnor U2104 (N_2104,N_769,N_1254);
xor U2105 (N_2105,N_746,N_1795);
and U2106 (N_2106,In_4898,N_1685);
or U2107 (N_2107,In_1175,In_2733);
and U2108 (N_2108,In_679,N_894);
xor U2109 (N_2109,N_1840,In_3259);
nor U2110 (N_2110,N_391,In_1335);
and U2111 (N_2111,In_3516,N_173);
xnor U2112 (N_2112,N_1160,In_104);
xor U2113 (N_2113,In_4216,In_1544);
xor U2114 (N_2114,In_2165,In_4982);
nor U2115 (N_2115,In_4488,In_871);
nand U2116 (N_2116,N_929,In_3080);
nor U2117 (N_2117,N_687,In_1564);
and U2118 (N_2118,N_1916,N_1796);
and U2119 (N_2119,In_102,N_1547);
nor U2120 (N_2120,N_1544,N_1987);
nand U2121 (N_2121,In_3633,In_3698);
xnor U2122 (N_2122,In_3887,In_2056);
or U2123 (N_2123,In_1328,N_664);
nand U2124 (N_2124,In_1919,In_596);
or U2125 (N_2125,In_2393,In_85);
or U2126 (N_2126,N_1667,In_3580);
nor U2127 (N_2127,In_835,In_251);
xor U2128 (N_2128,N_1438,N_2);
xor U2129 (N_2129,N_1880,In_4469);
and U2130 (N_2130,In_2217,N_1224);
and U2131 (N_2131,N_1966,N_1782);
nand U2132 (N_2132,In_2798,In_3718);
and U2133 (N_2133,In_2515,N_1121);
or U2134 (N_2134,In_3009,In_2233);
and U2135 (N_2135,In_1240,In_3570);
nand U2136 (N_2136,N_1453,N_818);
nor U2137 (N_2137,In_196,N_882);
nor U2138 (N_2138,N_1975,N_1699);
or U2139 (N_2139,In_4144,In_367);
xor U2140 (N_2140,In_1716,In_2136);
xnor U2141 (N_2141,In_1510,In_2947);
nor U2142 (N_2142,N_1521,N_1895);
nor U2143 (N_2143,In_3268,In_1484);
or U2144 (N_2144,In_2498,N_538);
nor U2145 (N_2145,N_1505,In_1881);
and U2146 (N_2146,N_620,In_868);
nor U2147 (N_2147,In_3963,N_56);
xnor U2148 (N_2148,N_1491,In_1152);
nor U2149 (N_2149,In_3279,N_888);
or U2150 (N_2150,In_1882,In_3904);
nand U2151 (N_2151,N_1621,N_1742);
xnor U2152 (N_2152,In_4636,N_99);
or U2153 (N_2153,In_64,In_1516);
nor U2154 (N_2154,N_1855,N_1041);
nand U2155 (N_2155,In_606,In_3851);
xnor U2156 (N_2156,N_775,N_1297);
nand U2157 (N_2157,N_1351,N_686);
and U2158 (N_2158,In_2313,N_1763);
xor U2159 (N_2159,In_2060,N_633);
and U2160 (N_2160,In_1169,In_4030);
and U2161 (N_2161,N_1163,N_1156);
nor U2162 (N_2162,N_615,In_3639);
nand U2163 (N_2163,N_1324,In_4783);
xnor U2164 (N_2164,N_163,N_1466);
nor U2165 (N_2165,In_1491,N_747);
or U2166 (N_2166,In_2747,N_1993);
nor U2167 (N_2167,N_1974,In_1980);
nor U2168 (N_2168,N_1166,N_947);
or U2169 (N_2169,N_632,In_655);
nand U2170 (N_2170,N_1596,N_1442);
xnor U2171 (N_2171,In_595,In_2206);
nor U2172 (N_2172,In_1599,N_1541);
nand U2173 (N_2173,N_1576,In_3397);
nand U2174 (N_2174,In_531,N_901);
and U2175 (N_2175,N_1159,In_4132);
or U2176 (N_2176,In_2267,N_1371);
nor U2177 (N_2177,In_1112,In_3874);
nand U2178 (N_2178,In_2087,In_1681);
or U2179 (N_2179,N_227,N_1780);
or U2180 (N_2180,In_4988,In_1419);
xor U2181 (N_2181,In_3506,N_972);
xnor U2182 (N_2182,In_3668,In_2590);
nor U2183 (N_2183,N_1228,In_722);
nor U2184 (N_2184,N_1943,N_1415);
xnor U2185 (N_2185,In_4009,In_993);
or U2186 (N_2186,In_657,In_1229);
nor U2187 (N_2187,In_3246,In_969);
or U2188 (N_2188,N_1485,N_1634);
xor U2189 (N_2189,N_417,In_3889);
nor U2190 (N_2190,In_4060,N_1312);
xor U2191 (N_2191,In_1075,N_1986);
nor U2192 (N_2192,N_836,N_1046);
nand U2193 (N_2193,N_1394,In_3535);
or U2194 (N_2194,N_1985,In_1893);
nand U2195 (N_2195,In_2887,In_4821);
xor U2196 (N_2196,In_4827,In_1807);
or U2197 (N_2197,In_1331,In_2855);
or U2198 (N_2198,N_652,N_1025);
xnor U2199 (N_2199,N_1112,N_1342);
and U2200 (N_2200,N_389,N_756);
nand U2201 (N_2201,N_1441,N_1800);
or U2202 (N_2202,In_2238,In_2560);
nor U2203 (N_2203,In_1833,N_1261);
nand U2204 (N_2204,In_2421,In_4292);
nor U2205 (N_2205,In_4674,N_1819);
nand U2206 (N_2206,N_1622,N_1701);
or U2207 (N_2207,In_4372,N_1911);
nor U2208 (N_2208,In_4878,N_586);
xnor U2209 (N_2209,N_714,In_1926);
nor U2210 (N_2210,N_104,N_1852);
nand U2211 (N_2211,In_1024,N_656);
nor U2212 (N_2212,In_1113,N_186);
nand U2213 (N_2213,In_2135,N_1955);
and U2214 (N_2214,In_1970,In_584);
nand U2215 (N_2215,In_790,In_2612);
nand U2216 (N_2216,In_3552,N_1653);
or U2217 (N_2217,In_1724,In_4052);
nand U2218 (N_2218,In_2809,In_615);
and U2219 (N_2219,N_1150,In_4836);
nor U2220 (N_2220,In_2026,In_984);
nor U2221 (N_2221,In_3979,N_1845);
xor U2222 (N_2222,N_418,In_4493);
nand U2223 (N_2223,In_4620,In_4202);
nand U2224 (N_2224,In_2061,N_1404);
xnor U2225 (N_2225,In_3608,In_1785);
xor U2226 (N_2226,N_1749,In_2598);
or U2227 (N_2227,N_704,N_12);
nand U2228 (N_2228,N_1834,N_1684);
nand U2229 (N_2229,N_509,In_2562);
nor U2230 (N_2230,N_529,In_3050);
xnor U2231 (N_2231,In_1478,In_1873);
xnor U2232 (N_2232,N_1939,N_1793);
or U2233 (N_2233,In_2055,N_1799);
and U2234 (N_2234,In_680,N_1607);
nor U2235 (N_2235,In_701,N_4);
nor U2236 (N_2236,In_2294,In_2784);
nand U2237 (N_2237,In_1363,N_1022);
nand U2238 (N_2238,N_1814,In_1815);
nor U2239 (N_2239,N_812,In_4677);
xnor U2240 (N_2240,N_1595,In_2201);
xor U2241 (N_2241,N_776,In_307);
xor U2242 (N_2242,In_4608,In_4379);
nand U2243 (N_2243,In_783,N_1940);
or U2244 (N_2244,N_1524,N_1761);
xor U2245 (N_2245,In_3607,In_4153);
nand U2246 (N_2246,In_211,In_4668);
and U2247 (N_2247,N_1345,N_1417);
nand U2248 (N_2248,In_2872,N_403);
nor U2249 (N_2249,In_1975,N_1317);
or U2250 (N_2250,In_4957,N_1860);
xor U2251 (N_2251,N_682,N_2205);
and U2252 (N_2252,In_4616,N_2192);
xor U2253 (N_2253,In_4087,N_1730);
xnor U2254 (N_2254,In_4152,N_2166);
or U2255 (N_2255,In_535,In_880);
xor U2256 (N_2256,N_1172,N_2077);
xnor U2257 (N_2257,In_3651,In_4919);
or U2258 (N_2258,In_2381,N_1930);
or U2259 (N_2259,N_1377,In_336);
nor U2260 (N_2260,In_3303,In_1213);
nor U2261 (N_2261,In_2776,N_1678);
xor U2262 (N_2262,In_986,In_4721);
or U2263 (N_2263,In_3754,N_1138);
nand U2264 (N_2264,N_219,In_599);
nand U2265 (N_2265,N_1821,N_1235);
and U2266 (N_2266,N_1818,N_703);
and U2267 (N_2267,In_2243,In_3206);
xor U2268 (N_2268,N_199,N_2222);
or U2269 (N_2269,N_1811,In_3582);
and U2270 (N_2270,N_1459,In_3785);
nor U2271 (N_2271,In_2308,In_1912);
nor U2272 (N_2272,In_3310,In_27);
nor U2273 (N_2273,N_644,In_4383);
or U2274 (N_2274,In_3643,In_1365);
nor U2275 (N_2275,In_3123,In_3063);
and U2276 (N_2276,N_251,In_2035);
nor U2277 (N_2277,N_1641,In_1327);
or U2278 (N_2278,In_99,In_3262);
or U2279 (N_2279,N_2230,N_673);
or U2280 (N_2280,In_3025,In_4063);
nor U2281 (N_2281,In_4323,In_4377);
nand U2282 (N_2282,N_1889,N_2064);
xor U2283 (N_2283,N_496,In_2759);
and U2284 (N_2284,N_1054,In_2782);
and U2285 (N_2285,N_2085,N_2231);
nand U2286 (N_2286,N_1989,In_2906);
nand U2287 (N_2287,N_1809,N_2038);
xor U2288 (N_2288,N_65,In_4989);
xnor U2289 (N_2289,N_2136,In_3413);
nand U2290 (N_2290,N_820,In_475);
and U2291 (N_2291,N_2220,N_1969);
and U2292 (N_2292,N_548,N_2140);
or U2293 (N_2293,In_2023,In_2403);
and U2294 (N_2294,N_1992,In_278);
nand U2295 (N_2295,In_1372,N_2152);
nand U2296 (N_2296,In_1068,In_2296);
nor U2297 (N_2297,N_1960,In_6);
nor U2298 (N_2298,In_4894,In_2029);
and U2299 (N_2299,N_1648,In_2492);
and U2300 (N_2300,In_3893,N_799);
and U2301 (N_2301,In_4386,In_4810);
xor U2302 (N_2302,In_2770,In_2208);
nand U2303 (N_2303,In_4367,In_3683);
and U2304 (N_2304,N_697,In_2249);
xnor U2305 (N_2305,N_968,In_1850);
xnor U2306 (N_2306,In_1711,N_1773);
nor U2307 (N_2307,N_1111,In_3693);
and U2308 (N_2308,N_1284,In_1985);
nand U2309 (N_2309,N_1861,In_4726);
or U2310 (N_2310,N_1938,In_2259);
xnor U2311 (N_2311,In_519,N_1392);
nand U2312 (N_2312,In_1697,N_677);
or U2313 (N_2313,In_1258,N_1075);
or U2314 (N_2314,In_247,In_4610);
xnor U2315 (N_2315,In_1086,N_1529);
xnor U2316 (N_2316,N_1871,In_4863);
and U2317 (N_2317,N_748,N_1635);
xnor U2318 (N_2318,N_655,N_81);
xor U2319 (N_2319,N_1887,N_1990);
nor U2320 (N_2320,In_1278,In_1313);
nand U2321 (N_2321,In_3950,N_1137);
nor U2322 (N_2322,N_1136,In_4364);
nand U2323 (N_2323,In_3125,N_627);
xnor U2324 (N_2324,N_313,In_4647);
and U2325 (N_2325,In_94,In_2173);
and U2326 (N_2326,In_1787,In_2835);
or U2327 (N_2327,N_815,In_356);
or U2328 (N_2328,N_942,In_2548);
and U2329 (N_2329,In_261,N_583);
nor U2330 (N_2330,In_4750,N_1724);
xor U2331 (N_2331,In_3312,N_1147);
nor U2332 (N_2332,In_1216,N_731);
nor U2333 (N_2333,In_2002,In_2952);
and U2334 (N_2334,N_1579,N_594);
nand U2335 (N_2335,N_1528,N_2142);
or U2336 (N_2336,In_1665,In_769);
or U2337 (N_2337,N_1813,N_1613);
and U2338 (N_2338,N_1526,N_1628);
xor U2339 (N_2339,In_2276,In_4940);
nor U2340 (N_2340,N_1363,N_2042);
or U2341 (N_2341,N_622,In_1839);
and U2342 (N_2342,In_3728,N_909);
xor U2343 (N_2343,In_2224,N_1820);
nor U2344 (N_2344,N_2208,In_3022);
or U2345 (N_2345,In_2951,N_136);
nor U2346 (N_2346,In_323,In_2955);
xnor U2347 (N_2347,N_1826,N_975);
xnor U2348 (N_2348,In_4921,N_1514);
and U2349 (N_2349,In_93,In_2330);
or U2350 (N_2350,N_1873,N_1679);
and U2351 (N_2351,In_54,In_716);
nor U2352 (N_2352,In_745,In_3368);
nor U2353 (N_2353,In_1032,In_558);
nor U2354 (N_2354,In_3178,N_2133);
xnor U2355 (N_2355,In_1256,In_4491);
nor U2356 (N_2356,In_4552,In_2917);
nand U2357 (N_2357,In_3572,In_2655);
nor U2358 (N_2358,In_3786,N_1443);
or U2359 (N_2359,N_1329,In_441);
and U2360 (N_2360,In_1405,N_2082);
xor U2361 (N_2361,In_1437,In_893);
nand U2362 (N_2362,In_4560,N_934);
and U2363 (N_2363,In_3605,In_4025);
xnor U2364 (N_2364,In_2925,N_2187);
and U2365 (N_2365,In_4007,N_1429);
xor U2366 (N_2366,In_1130,N_495);
xnor U2367 (N_2367,N_790,In_3351);
nand U2368 (N_2368,N_781,In_4495);
or U2369 (N_2369,In_2954,N_1586);
nor U2370 (N_2370,N_1804,N_1950);
or U2371 (N_2371,N_1636,N_520);
or U2372 (N_2372,In_3719,In_1901);
or U2373 (N_2373,In_3857,N_1683);
nor U2374 (N_2374,In_1602,In_4473);
xnor U2375 (N_2375,N_1891,In_3107);
nand U2376 (N_2376,In_4223,N_2171);
nand U2377 (N_2377,N_1483,N_1448);
and U2378 (N_2378,In_4566,N_2035);
xor U2379 (N_2379,In_2714,In_135);
nor U2380 (N_2380,In_3245,In_1914);
nand U2381 (N_2381,In_1968,N_1841);
nand U2382 (N_2382,In_2743,N_1903);
nor U2383 (N_2383,N_229,In_2497);
and U2384 (N_2384,N_2021,In_3868);
nor U2385 (N_2385,In_182,In_1453);
nor U2386 (N_2386,In_2892,N_1732);
nor U2387 (N_2387,N_701,In_2471);
and U2388 (N_2388,In_395,In_284);
nor U2389 (N_2389,N_2176,In_4869);
and U2390 (N_2390,In_3459,N_1649);
xnor U2391 (N_2391,In_1166,In_2209);
nand U2392 (N_2392,N_2138,N_1816);
or U2393 (N_2393,In_2000,N_884);
or U2394 (N_2394,N_1728,N_572);
and U2395 (N_2395,In_3658,N_2121);
nor U2396 (N_2396,In_375,N_1831);
nor U2397 (N_2397,In_2153,In_3113);
and U2398 (N_2398,N_160,N_2119);
xnor U2399 (N_2399,In_1444,In_3480);
or U2400 (N_2400,In_1201,N_1315);
or U2401 (N_2401,N_2207,N_1868);
nor U2402 (N_2402,N_1268,N_320);
nand U2403 (N_2403,In_2916,N_1615);
and U2404 (N_2404,In_242,In_1133);
or U2405 (N_2405,N_2204,In_3176);
or U2406 (N_2406,N_2079,In_1164);
and U2407 (N_2407,N_770,In_4935);
nand U2408 (N_2408,In_158,In_4185);
xor U2409 (N_2409,N_1250,N_2108);
nor U2410 (N_2410,In_1852,In_1627);
and U2411 (N_2411,In_2394,N_2013);
nand U2412 (N_2412,In_2336,N_958);
xnor U2413 (N_2413,In_1712,N_2054);
or U2414 (N_2414,N_440,N_310);
and U2415 (N_2415,In_2774,In_2461);
nor U2416 (N_2416,In_1279,N_443);
nand U2417 (N_2417,In_1018,N_1543);
xor U2418 (N_2418,In_4747,In_3770);
and U2419 (N_2419,In_3257,N_1389);
and U2420 (N_2420,In_2139,N_2084);
and U2421 (N_2421,In_1735,In_3997);
xor U2422 (N_2422,N_873,In_406);
and U2423 (N_2423,In_3909,In_3495);
xnor U2424 (N_2424,In_2768,N_807);
nand U2425 (N_2425,In_4581,In_3577);
nand U2426 (N_2426,In_2679,In_2418);
xor U2427 (N_2427,N_1734,N_1070);
or U2428 (N_2428,N_77,N_91);
nand U2429 (N_2429,In_855,N_847);
and U2430 (N_2430,In_1941,N_1294);
nand U2431 (N_2431,N_646,In_3566);
nand U2432 (N_2432,N_2000,N_1326);
nand U2433 (N_2433,In_870,In_56);
or U2434 (N_2434,N_1201,In_4537);
nand U2435 (N_2435,N_413,N_1251);
nor U2436 (N_2436,In_3161,In_3117);
xnor U2437 (N_2437,N_1113,N_1542);
nand U2438 (N_2438,N_2094,In_4923);
or U2439 (N_2439,N_1827,In_1060);
xnor U2440 (N_2440,In_1925,N_1064);
and U2441 (N_2441,In_2360,N_1339);
nor U2442 (N_2442,N_1017,In_2717);
nor U2443 (N_2443,N_1918,In_860);
xor U2444 (N_2444,N_1219,N_1998);
or U2445 (N_2445,In_3398,N_1538);
xor U2446 (N_2446,In_3053,In_4000);
nand U2447 (N_2447,N_518,N_406);
xnor U2448 (N_2448,In_1877,N_1355);
and U2449 (N_2449,In_2079,In_4175);
nor U2450 (N_2450,N_1331,In_2338);
and U2451 (N_2451,N_1802,N_1645);
xnor U2452 (N_2452,N_1937,N_1559);
or U2453 (N_2453,N_37,N_2080);
xor U2454 (N_2454,In_2062,In_296);
and U2455 (N_2455,N_2107,N_1561);
nor U2456 (N_2456,N_617,In_623);
nor U2457 (N_2457,In_4818,N_1905);
nand U2458 (N_2458,In_577,N_1922);
xnor U2459 (N_2459,In_77,In_2817);
nor U2460 (N_2460,N_1712,N_2189);
nand U2461 (N_2461,N_151,In_1565);
and U2462 (N_2462,N_2052,In_1410);
xnor U2463 (N_2463,In_796,In_3775);
xor U2464 (N_2464,In_3739,N_1713);
or U2465 (N_2465,N_452,N_1218);
or U2466 (N_2466,In_1615,In_4090);
or U2467 (N_2467,In_2012,In_2861);
and U2468 (N_2468,In_1577,N_2194);
or U2469 (N_2469,N_1018,In_3401);
and U2470 (N_2470,N_2015,In_1805);
and U2471 (N_2471,In_4741,In_3100);
xor U2472 (N_2472,N_2093,In_3843);
nand U2473 (N_2473,N_1629,In_1600);
or U2474 (N_2474,In_385,In_3758);
xnor U2475 (N_2475,In_2946,In_1703);
nand U2476 (N_2476,In_4800,In_3032);
and U2477 (N_2477,N_2105,In_4088);
and U2478 (N_2478,N_837,In_175);
xnor U2479 (N_2479,In_467,In_974);
nor U2480 (N_2480,N_828,N_2069);
xor U2481 (N_2481,In_1993,In_350);
nand U2482 (N_2482,In_3692,N_2165);
and U2483 (N_2483,In_4589,N_1455);
nor U2484 (N_2484,In_1078,N_1610);
xnor U2485 (N_2485,In_1871,N_824);
and U2486 (N_2486,N_1847,N_1872);
nor U2487 (N_2487,In_3561,N_1245);
or U2488 (N_2488,N_407,N_1765);
nor U2489 (N_2489,N_1021,In_3131);
or U2490 (N_2490,N_2153,N_1661);
nand U2491 (N_2491,N_1924,In_4228);
nand U2492 (N_2492,N_2144,N_494);
and U2493 (N_2493,In_1051,N_1273);
xnor U2494 (N_2494,N_1952,N_2247);
nand U2495 (N_2495,N_337,N_1214);
xnor U2496 (N_2496,N_1973,N_410);
and U2497 (N_2497,In_4122,N_428);
or U2498 (N_2498,N_1995,N_1931);
xnor U2499 (N_2499,In_361,In_3638);
nor U2500 (N_2500,N_2177,In_1747);
and U2501 (N_2501,N_546,N_1812);
or U2502 (N_2502,N_1539,N_2028);
xor U2503 (N_2503,In_71,N_1352);
and U2504 (N_2504,N_2216,In_983);
and U2505 (N_2505,In_1177,N_2041);
xnor U2506 (N_2506,In_1989,N_1614);
and U2507 (N_2507,N_80,In_883);
nand U2508 (N_2508,N_759,N_1307);
nand U2509 (N_2509,N_2203,In_488);
xnor U2510 (N_2510,N_1705,N_1605);
nand U2511 (N_2511,N_1851,N_1152);
xor U2512 (N_2512,In_808,In_3374);
xnor U2513 (N_2513,In_4439,N_2332);
or U2514 (N_2514,In_1418,In_2013);
nand U2515 (N_2515,In_4962,In_636);
or U2516 (N_2516,N_1167,N_2299);
or U2517 (N_2517,In_1537,In_733);
nand U2518 (N_2518,In_2753,N_2408);
and U2519 (N_2519,N_2201,N_2265);
xnor U2520 (N_2520,In_591,N_2483);
and U2521 (N_2521,In_2545,N_2103);
and U2522 (N_2522,N_1964,In_2192);
nor U2523 (N_2523,N_2461,In_662);
nor U2524 (N_2524,N_2293,In_1527);
xor U2525 (N_2525,N_2477,In_764);
and U2526 (N_2526,N_780,N_811);
xor U2527 (N_2527,N_1704,N_2442);
nand U2528 (N_2528,In_4642,N_2090);
and U2529 (N_2529,N_2072,N_1141);
nand U2530 (N_2530,N_2097,In_1272);
nor U2531 (N_2531,In_4207,N_228);
or U2532 (N_2532,In_2814,N_591);
xor U2533 (N_2533,In_3062,In_1938);
nand U2534 (N_2534,N_2320,N_1581);
or U2535 (N_2535,N_2481,N_2313);
and U2536 (N_2536,N_2322,In_1132);
nand U2537 (N_2537,In_4554,In_1420);
xnor U2538 (N_2538,In_2931,N_2292);
and U2539 (N_2539,N_2278,N_73);
and U2540 (N_2540,In_3924,In_673);
nor U2541 (N_2541,N_2061,In_1643);
xor U2542 (N_2542,In_2666,N_2223);
nand U2543 (N_2543,In_2698,In_672);
xnor U2544 (N_2544,N_961,N_946);
or U2545 (N_2545,N_2363,N_675);
and U2546 (N_2546,In_4104,In_447);
xor U2547 (N_2547,In_319,N_684);
or U2548 (N_2548,In_3612,N_2274);
xor U2549 (N_2549,N_1104,N_1906);
xor U2550 (N_2550,In_2539,In_3989);
or U2551 (N_2551,In_245,In_4864);
and U2552 (N_2552,In_823,In_4571);
and U2553 (N_2553,N_1259,N_2424);
xor U2554 (N_2554,N_2115,In_4978);
and U2555 (N_2555,N_925,In_1865);
nor U2556 (N_2556,N_1520,N_1604);
and U2557 (N_2557,In_2637,In_4002);
nand U2558 (N_2558,In_3914,N_1962);
nor U2559 (N_2559,N_2348,In_2706);
nand U2560 (N_2560,In_1064,N_1464);
nand U2561 (N_2561,In_2032,In_1349);
xnor U2562 (N_2562,In_3046,In_3375);
nand U2563 (N_2563,N_2047,In_3664);
or U2564 (N_2564,In_2846,N_360);
or U2565 (N_2565,N_1055,In_4691);
nand U2566 (N_2566,In_611,In_1511);
nand U2567 (N_2567,N_1568,In_252);
or U2568 (N_2568,N_1502,In_3130);
nand U2569 (N_2569,In_4872,N_2065);
and U2570 (N_2570,In_2819,In_2470);
or U2571 (N_2571,In_3743,In_570);
and U2572 (N_2572,N_1706,N_1801);
and U2573 (N_2573,In_4786,In_3519);
and U2574 (N_2574,N_2214,In_695);
nor U2575 (N_2575,N_2284,In_4992);
nor U2576 (N_2576,N_1673,N_2100);
or U2577 (N_2577,N_1032,In_1118);
nand U2578 (N_2578,In_4269,In_358);
nor U2579 (N_2579,In_173,N_2074);
xor U2580 (N_2580,N_1222,In_291);
nor U2581 (N_2581,N_2301,In_4105);
and U2582 (N_2582,In_2220,N_2316);
xnor U2583 (N_2583,N_15,N_1431);
or U2584 (N_2584,In_1138,N_1716);
or U2585 (N_2585,N_1956,N_660);
nand U2586 (N_2586,In_201,N_2025);
nand U2587 (N_2587,N_2347,N_892);
or U2588 (N_2588,N_1609,N_1798);
nand U2589 (N_2589,In_2826,In_2310);
xnor U2590 (N_2590,N_1296,N_1593);
xnor U2591 (N_2591,N_2454,N_2295);
nand U2592 (N_2592,In_425,In_4653);
nand U2593 (N_2593,In_2919,In_3588);
nand U2594 (N_2594,In_370,In_267);
xnor U2595 (N_2595,In_4222,N_2050);
nand U2596 (N_2596,N_1680,N_2306);
nand U2597 (N_2597,In_1591,In_4870);
xor U2598 (N_2598,N_557,N_2470);
or U2599 (N_2599,In_3504,N_2209);
nand U2600 (N_2600,N_2305,In_1154);
nor U2601 (N_2601,In_1561,In_392);
nand U2602 (N_2602,N_1523,N_2418);
nand U2603 (N_2603,In_3652,In_2625);
nand U2604 (N_2604,In_4825,In_3240);
and U2605 (N_2605,N_1907,N_2492);
nand U2606 (N_2606,N_885,N_116);
xor U2607 (N_2607,N_1480,In_4260);
and U2608 (N_2608,N_1423,N_387);
or U2609 (N_2609,In_4359,In_2105);
nor U2610 (N_2610,N_2149,N_1557);
xor U2611 (N_2611,In_741,In_2883);
xor U2612 (N_2612,N_1449,In_3359);
and U2613 (N_2613,N_1947,In_1586);
nand U2614 (N_2614,N_700,N_1275);
xnor U2615 (N_2615,In_2424,In_2339);
or U2616 (N_2616,N_2132,N_1063);
xnor U2617 (N_2617,N_1869,In_2749);
xor U2618 (N_2618,N_521,In_1790);
nand U2619 (N_2619,N_2441,N_1319);
xor U2620 (N_2620,In_4565,N_1954);
xnor U2621 (N_2621,N_1825,N_2428);
and U2622 (N_2622,In_4568,N_2388);
nor U2623 (N_2623,In_4484,N_2087);
xor U2624 (N_2624,N_1602,N_1242);
xnor U2625 (N_2625,In_4716,In_2609);
nor U2626 (N_2626,In_118,In_74);
and U2627 (N_2627,In_547,In_1798);
and U2628 (N_2628,In_3796,N_351);
or U2629 (N_2629,In_181,In_3955);
nand U2630 (N_2630,In_1624,In_400);
and U2631 (N_2631,N_2211,N_1518);
or U2632 (N_2632,In_2715,In_980);
or U2633 (N_2633,N_177,N_1569);
xnor U2634 (N_2634,N_725,In_1736);
or U2635 (N_2635,N_1994,N_2400);
or U2636 (N_2636,N_568,In_2097);
nor U2637 (N_2637,N_1875,In_132);
nor U2638 (N_2638,N_1963,In_1347);
nor U2639 (N_2639,In_403,N_154);
xor U2640 (N_2640,In_3143,N_1849);
or U2641 (N_2641,N_1508,In_2458);
nand U2642 (N_2642,N_2340,In_79);
and U2643 (N_2643,In_3757,N_1384);
and U2644 (N_2644,In_4130,N_1832);
or U2645 (N_2645,In_1801,N_2395);
nand U2646 (N_2646,N_1437,N_2030);
and U2647 (N_2647,N_1785,N_1927);
or U2648 (N_2648,N_1867,N_1549);
nand U2649 (N_2649,N_1346,In_4824);
xor U2650 (N_2650,In_4835,N_2385);
xor U2651 (N_2651,In_1756,In_3595);
or U2652 (N_2652,N_846,N_1676);
nand U2653 (N_2653,In_1300,In_962);
nor U2654 (N_2654,N_200,N_1234);
and U2655 (N_2655,N_1612,In_2455);
or U2656 (N_2656,In_2386,In_1293);
and U2657 (N_2657,N_1708,N_930);
xnor U2658 (N_2658,N_1122,In_1069);
nand U2659 (N_2659,N_1850,In_2183);
or U2660 (N_2660,In_1171,In_3217);
nand U2661 (N_2661,In_4986,N_2401);
xnor U2662 (N_2662,In_3027,N_1846);
nand U2663 (N_2663,In_1380,N_2168);
nor U2664 (N_2664,In_2797,In_3023);
and U2665 (N_2665,In_1151,In_998);
nor U2666 (N_2666,N_709,In_221);
nor U2667 (N_2667,In_583,N_1330);
and U2668 (N_2668,In_3970,In_728);
or U2669 (N_2669,N_1368,N_263);
xnor U2670 (N_2670,N_2200,In_4073);
xor U2671 (N_2671,In_1211,N_516);
nand U2672 (N_2672,In_3079,N_906);
and U2673 (N_2673,N_78,N_1478);
nand U2674 (N_2674,In_3731,N_1434);
nand U2675 (N_2675,In_229,In_3705);
or U2676 (N_2676,N_710,In_89);
and U2677 (N_2677,In_518,In_939);
and U2678 (N_2678,N_2456,In_846);
xnor U2679 (N_2679,In_4455,N_30);
xor U2680 (N_2680,In_545,N_2233);
or U2681 (N_2681,N_1185,N_279);
and U2682 (N_2682,N_1372,In_2543);
nor U2683 (N_2683,In_2120,In_4564);
nor U2684 (N_2684,In_956,In_4424);
nand U2685 (N_2685,In_114,In_4148);
or U2686 (N_2686,In_161,In_506);
nor U2687 (N_2687,N_598,N_29);
nand U2688 (N_2688,In_2737,N_436);
nand U2689 (N_2689,N_1771,In_259);
nand U2690 (N_2690,In_2891,In_4697);
nor U2691 (N_2691,In_1226,In_2380);
nand U2692 (N_2692,N_2242,N_2279);
or U2693 (N_2693,In_2750,N_1082);
nand U2694 (N_2694,In_3336,In_1342);
xnor U2695 (N_2695,N_342,N_1145);
and U2696 (N_2696,In_4932,In_2247);
nor U2697 (N_2697,In_4162,In_3212);
nor U2698 (N_2698,In_3417,In_2860);
nand U2699 (N_2699,In_2605,N_1967);
or U2700 (N_2700,N_2023,N_636);
and U2701 (N_2701,N_619,N_2236);
nand U2702 (N_2702,In_4210,N_1571);
nor U2703 (N_2703,N_1751,N_2235);
or U2704 (N_2704,N_195,In_4347);
xnor U2705 (N_2705,In_493,In_511);
xor U2706 (N_2706,In_1406,In_4482);
xnor U2707 (N_2707,N_1468,N_255);
xor U2708 (N_2708,N_735,N_2303);
nor U2709 (N_2709,N_95,In_3927);
and U2710 (N_2710,N_1890,N_1833);
and U2711 (N_2711,In_2059,N_863);
xnor U2712 (N_2712,In_2178,N_2158);
nand U2713 (N_2713,N_1754,N_2004);
nand U2714 (N_2714,In_4930,In_1000);
nor U2715 (N_2715,In_1937,In_2920);
xnor U2716 (N_2716,In_2113,N_1920);
and U2717 (N_2717,In_4249,N_2113);
nor U2718 (N_2718,In_3092,N_893);
nand U2719 (N_2719,N_621,N_1074);
or U2720 (N_2720,In_1341,In_1828);
nand U2721 (N_2721,In_160,N_1980);
xor U2722 (N_2722,In_2538,N_825);
nand U2723 (N_2723,N_2249,In_1007);
and U2724 (N_2724,N_2116,N_1531);
nor U2725 (N_2725,N_544,In_1161);
nand U2726 (N_2726,In_4572,N_922);
nor U2727 (N_2727,N_1096,N_2261);
or U2728 (N_2728,In_1754,N_1965);
nand U2729 (N_2729,N_140,In_3215);
nand U2730 (N_2730,N_2078,N_1378);
nand U2731 (N_2731,In_434,In_4855);
nand U2732 (N_2732,N_1774,In_3967);
nor U2733 (N_2733,N_982,N_295);
nor U2734 (N_2734,In_582,N_798);
or U2735 (N_2735,N_976,In_786);
nand U2736 (N_2736,N_2493,N_2392);
nand U2737 (N_2737,In_4031,In_820);
nand U2738 (N_2738,N_2359,N_1864);
nor U2739 (N_2739,N_2276,N_1501);
nand U2740 (N_2740,In_374,N_1893);
nand U2741 (N_2741,N_1737,N_1689);
xor U2742 (N_2742,N_1740,N_933);
nor U2743 (N_2743,In_2028,N_1416);
and U2744 (N_2744,N_613,In_4293);
and U2745 (N_2745,In_2287,In_1878);
nand U2746 (N_2746,N_1694,In_3264);
nor U2747 (N_2747,In_1383,In_4213);
or U2748 (N_2748,In_785,N_131);
nand U2749 (N_2749,In_1456,N_1340);
or U2750 (N_2750,In_4911,In_525);
and U2751 (N_2751,In_1057,N_1332);
xnor U2752 (N_2752,In_1739,N_567);
xor U2753 (N_2753,In_929,N_2338);
nand U2754 (N_2754,N_2039,In_1084);
and U2755 (N_2755,N_1589,N_2651);
nand U2756 (N_2756,N_2386,N_1290);
xnor U2757 (N_2757,In_476,In_926);
xnor U2758 (N_2758,In_2350,N_2479);
xor U2759 (N_2759,In_4525,N_712);
or U2760 (N_2760,N_1440,N_493);
and U2761 (N_2761,N_605,N_1598);
nor U2762 (N_2762,N_2071,N_874);
nand U2763 (N_2763,In_2199,N_1546);
and U2764 (N_2764,In_2941,N_662);
xor U2765 (N_2765,N_1631,N_425);
xnor U2766 (N_2766,In_244,N_2537);
xnor U2767 (N_2767,N_2707,N_2583);
nor U2768 (N_2768,In_1259,In_501);
and U2769 (N_2769,In_4058,N_564);
xnor U2770 (N_2770,N_2725,N_904);
xnor U2771 (N_2771,N_1726,In_2506);
nor U2772 (N_2772,In_1196,N_2059);
nor U2773 (N_2773,N_2031,In_4680);
xor U2774 (N_2774,In_665,In_4601);
and U2775 (N_2775,N_2405,N_2180);
nand U2776 (N_2776,N_2611,N_2129);
and U2777 (N_2777,N_294,In_199);
and U2778 (N_2778,N_603,N_1433);
nand U2779 (N_2779,In_213,In_4441);
xnor U2780 (N_2780,In_1350,In_1357);
and U2781 (N_2781,In_881,N_1925);
xnor U2782 (N_2782,In_4905,N_2264);
nand U2783 (N_2783,N_519,In_4638);
nor U2784 (N_2784,In_724,N_2569);
xnor U2785 (N_2785,In_707,N_133);
or U2786 (N_2786,In_3005,N_559);
nor U2787 (N_2787,N_1320,N_1522);
and U2788 (N_2788,N_321,In_3892);
xnor U2789 (N_2789,N_1654,N_1866);
or U2790 (N_2790,N_792,In_1974);
or U2791 (N_2791,N_2542,N_1913);
nor U2792 (N_2792,N_2719,In_4303);
and U2793 (N_2793,N_1322,N_2036);
and U2794 (N_2794,In_394,N_2749);
nand U2795 (N_2795,In_4955,N_2110);
and U2796 (N_2796,In_2118,In_3229);
xnor U2797 (N_2797,In_3856,In_1186);
nand U2798 (N_2798,N_1806,In_4479);
xor U2799 (N_2799,In_2915,N_2239);
nor U2800 (N_2800,N_2297,N_2574);
xor U2801 (N_2801,N_2687,N_2335);
xnor U2802 (N_2802,N_1949,In_4664);
nor U2803 (N_2803,N_585,In_2332);
nor U2804 (N_2804,N_1808,In_308);
and U2805 (N_2805,N_1479,N_1489);
and U2806 (N_2806,N_2268,In_950);
nor U2807 (N_2807,N_1817,N_2742);
xor U2808 (N_2808,In_2352,In_4888);
nor U2809 (N_2809,N_535,In_2636);
nand U2810 (N_2810,N_2536,In_3861);
and U2811 (N_2811,In_2293,N_1976);
xor U2812 (N_2812,In_3685,N_2309);
and U2813 (N_2813,In_4251,In_1930);
and U2814 (N_2814,N_1739,In_4848);
xor U2815 (N_2815,N_2304,N_2548);
nor U2816 (N_2816,N_2664,In_4262);
nor U2817 (N_2817,N_1288,N_2383);
and U2818 (N_2818,In_3121,N_2259);
xor U2819 (N_2819,N_2244,N_1775);
or U2820 (N_2820,N_286,N_2262);
or U2821 (N_2821,N_1421,N_2411);
nor U2822 (N_2822,In_1677,In_3418);
nor U2823 (N_2823,In_3828,In_225);
or U2824 (N_2824,N_1146,N_2019);
and U2825 (N_2825,N_2691,N_2101);
nand U2826 (N_2826,In_4634,N_2377);
nand U2827 (N_2827,In_2044,N_2426);
or U2828 (N_2828,N_305,N_551);
or U2829 (N_2829,N_919,N_895);
or U2830 (N_2830,In_4321,In_2405);
nor U2831 (N_2831,In_2496,N_1627);
and U2832 (N_2832,In_4103,In_2689);
and U2833 (N_2833,In_2631,N_561);
nand U2834 (N_2834,In_4900,N_2354);
xor U2835 (N_2835,In_3863,N_2497);
xor U2836 (N_2836,In_4886,N_2022);
and U2837 (N_2837,N_170,N_2436);
and U2838 (N_2838,N_2638,N_716);
xnor U2839 (N_2839,N_650,In_1784);
and U2840 (N_2840,In_111,N_963);
xnor U2841 (N_2841,In_3101,In_2376);
nand U2842 (N_2842,N_2689,In_1053);
or U2843 (N_2843,N_2314,In_3456);
or U2844 (N_2844,N_1857,In_3443);
nor U2845 (N_2845,In_1047,In_1719);
or U2846 (N_2846,In_1505,N_2727);
and U2847 (N_2847,N_2724,N_2450);
or U2848 (N_2848,In_297,In_3369);
or U2849 (N_2849,N_2040,N_1878);
xor U2850 (N_2850,In_2396,N_1946);
or U2851 (N_2851,In_2180,N_1469);
nor U2852 (N_2852,In_3907,In_3832);
xor U2853 (N_2853,N_1692,N_749);
and U2854 (N_2854,In_4558,N_426);
and U2855 (N_2855,N_1932,N_920);
xnor U2856 (N_2856,In_1792,N_1983);
and U2857 (N_2857,In_3414,N_1848);
xor U2858 (N_2858,N_2487,N_1042);
nor U2859 (N_2859,N_2625,In_4596);
nor U2860 (N_2860,In_3812,N_2679);
or U2861 (N_2861,In_3787,In_1094);
xnor U2862 (N_2862,In_2630,In_1345);
xnor U2863 (N_2863,N_2151,N_995);
nor U2864 (N_2864,N_1720,N_479);
or U2865 (N_2865,N_755,N_378);
or U2866 (N_2866,N_2352,N_2520);
or U2867 (N_2867,N_2653,N_2033);
xor U2868 (N_2868,N_2500,N_480);
or U2869 (N_2869,In_1101,N_2494);
or U2870 (N_2870,N_754,N_555);
nand U2871 (N_2871,N_1139,N_1056);
and U2872 (N_2872,N_2126,N_2665);
and U2873 (N_2873,In_230,In_3334);
nand U2874 (N_2874,In_1648,N_540);
nand U2875 (N_2875,In_3881,N_2485);
or U2876 (N_2876,In_2479,In_1371);
xnor U2877 (N_2877,N_2632,In_4414);
nor U2878 (N_2878,N_2291,N_1824);
xnor U2879 (N_2879,N_1390,In_4879);
and U2880 (N_2880,In_3001,N_2228);
nor U2881 (N_2881,N_96,In_2914);
xor U2882 (N_2882,In_1663,In_3545);
and U2883 (N_2883,N_2125,N_2604);
xor U2884 (N_2884,In_4151,In_658);
xor U2885 (N_2885,In_1812,N_2051);
nor U2886 (N_2886,In_1614,In_4078);
or U2887 (N_2887,N_2182,N_233);
xor U2888 (N_2888,In_3145,N_2349);
and U2889 (N_2889,N_2367,N_149);
nand U2890 (N_2890,In_1906,In_1767);
and U2891 (N_2891,In_1176,N_1555);
xnor U2892 (N_2892,N_2601,N_2056);
or U2893 (N_2893,In_3935,N_2195);
nand U2894 (N_2894,In_462,In_1242);
or U2895 (N_2895,In_325,In_1632);
xnor U2896 (N_2896,In_4542,N_213);
xnor U2897 (N_2897,In_1519,In_2427);
or U2898 (N_2898,N_1318,In_2039);
xor U2899 (N_2899,N_1001,N_141);
nand U2900 (N_2900,In_912,In_4411);
or U2901 (N_2901,N_122,In_1339);
or U2902 (N_2902,In_4083,N_18);
xnor U2903 (N_2903,N_2190,N_1666);
nor U2904 (N_2904,In_2246,N_1498);
nand U2905 (N_2905,In_3300,N_1258);
and U2906 (N_2906,N_806,N_1626);
nor U2907 (N_2907,In_3673,N_2333);
or U2908 (N_2908,N_2407,N_2218);
xnor U2909 (N_2909,N_1999,N_2057);
xor U2910 (N_2910,N_768,In_1147);
nand U2911 (N_2911,N_41,N_2315);
nand U2912 (N_2912,In_1609,In_2214);
and U2913 (N_2913,N_1746,N_2731);
and U2914 (N_2914,N_1580,In_3946);
xor U2915 (N_2915,In_4574,N_2114);
xnor U2916 (N_2916,N_2421,N_854);
or U2917 (N_2917,N_1052,In_4615);
nand U2918 (N_2918,In_4943,N_2296);
nor U2919 (N_2919,In_3468,In_605);
and U2920 (N_2920,In_1038,In_1963);
xnor U2921 (N_2921,In_3449,In_2502);
nor U2922 (N_2922,In_4284,N_1279);
xnor U2923 (N_2923,N_1472,N_398);
nor U2924 (N_2924,N_362,N_1577);
and U2925 (N_2925,N_2647,N_2646);
nor U2926 (N_2926,N_2453,In_4345);
nand U2927 (N_2927,N_1174,N_2083);
or U2928 (N_2928,N_2538,N_2394);
or U2929 (N_2929,In_4541,N_1587);
nand U2930 (N_2930,N_2661,N_783);
and U2931 (N_2931,In_167,In_638);
or U2932 (N_2932,N_1277,In_2974);
and U2933 (N_2933,N_1738,N_2008);
or U2934 (N_2934,In_3083,In_192);
and U2935 (N_2935,N_262,N_2438);
nand U2936 (N_2936,N_2368,In_3745);
nand U2937 (N_2937,N_2682,N_1247);
nor U2938 (N_2938,N_2525,In_3689);
or U2939 (N_2939,In_1506,N_86);
xnor U2940 (N_2940,N_2444,N_2396);
xnor U2941 (N_2941,N_2232,N_2370);
nand U2942 (N_2942,N_2413,In_3978);
nand U2943 (N_2943,In_4754,In_207);
nor U2944 (N_2944,N_2219,N_1776);
nand U2945 (N_2945,In_968,N_1600);
and U2946 (N_2946,N_891,N_2167);
nand U2947 (N_2947,N_2513,N_2582);
or U2948 (N_2948,N_2435,N_2716);
nor U2949 (N_2949,In_1539,N_2578);
xnor U2950 (N_2950,N_2570,In_3067);
or U2951 (N_2951,In_4576,N_611);
nor U2952 (N_2952,In_4312,N_1182);
and U2953 (N_2953,N_1711,N_2663);
xor U2954 (N_2954,N_1029,In_3256);
xor U2955 (N_2955,N_537,N_1910);
xnor U2956 (N_2956,N_2594,In_4669);
nor U2957 (N_2957,N_2654,In_1082);
xor U2958 (N_2958,N_1718,N_1642);
nand U2959 (N_2959,In_451,In_148);
nand U2960 (N_2960,In_2572,In_18);
nor U2961 (N_2961,N_2043,N_2726);
xor U2962 (N_2962,N_1567,N_2254);
and U2963 (N_2963,In_2990,N_2575);
xnor U2964 (N_2964,In_480,N_363);
and U2965 (N_2965,N_114,N_2154);
nor U2966 (N_2966,N_1086,In_2576);
nor U2967 (N_2967,In_3434,In_2616);
and U2968 (N_2968,In_4760,N_2480);
xor U2969 (N_2969,In_2483,N_144);
xnor U2970 (N_2970,N_481,N_1582);
and U2971 (N_2971,N_845,N_1011);
nand U2972 (N_2972,N_1039,N_2141);
and U2973 (N_2973,N_1815,In_4977);
nor U2974 (N_2974,In_222,In_3644);
nor U2975 (N_2975,In_2130,In_4317);
nand U2976 (N_2976,N_1853,In_4890);
and U2977 (N_2977,In_2357,N_1865);
nor U2978 (N_2978,N_1494,In_2799);
nand U2979 (N_2979,In_2653,In_4884);
xnor U2980 (N_2980,N_2088,N_124);
nor U2981 (N_2981,In_2416,N_2243);
nand U2982 (N_2982,N_1335,In_2211);
nor U2983 (N_2983,N_14,N_2312);
or U2984 (N_2984,N_1693,In_1762);
and U2985 (N_2985,N_1791,N_2344);
or U2986 (N_2986,In_4049,In_981);
nand U2987 (N_2987,N_1948,In_2592);
and U2988 (N_2988,N_430,In_988);
nand U2989 (N_2989,N_2252,In_0);
or U2990 (N_2990,In_1145,N_2577);
and U2991 (N_2991,N_2657,In_1326);
xor U2992 (N_2992,N_256,N_1467);
nand U2993 (N_2993,N_2416,N_1072);
nand U2994 (N_2994,In_2116,N_1278);
and U2995 (N_2995,N_2572,N_852);
nor U2996 (N_2996,In_3339,N_1227);
nor U2997 (N_2997,In_2235,In_3928);
or U2998 (N_2998,N_1698,In_3699);
nand U2999 (N_2999,In_4914,N_250);
xor U3000 (N_3000,N_2584,N_1271);
or U3001 (N_3001,In_455,N_2449);
nand U3002 (N_3002,In_4531,N_2286);
xor U3003 (N_3003,In_2298,N_1617);
nor U3004 (N_3004,N_2860,N_2760);
and U3005 (N_3005,N_1991,N_2747);
or U3006 (N_3006,N_1451,N_2649);
and U3007 (N_3007,N_2770,N_2202);
nand U3008 (N_3008,In_3322,N_1280);
xor U3009 (N_3009,In_3630,N_2835);
nor U3010 (N_3010,In_1613,N_2884);
and U3011 (N_3011,In_3499,In_372);
nand U3012 (N_3012,In_4547,N_2193);
xor U3013 (N_3013,In_3790,In_523);
xnor U3014 (N_3014,N_1412,N_1722);
nor U3015 (N_3015,N_1601,In_1851);
nor U3016 (N_3016,In_1883,In_526);
and U3017 (N_3017,N_883,N_1700);
and U3018 (N_3018,N_2155,In_1088);
or U3019 (N_3019,N_2592,N_2973);
or U3020 (N_3020,In_234,N_577);
nand U3021 (N_3021,In_410,N_2362);
xnor U3022 (N_3022,N_1630,N_2784);
and U3023 (N_3023,In_1473,In_1299);
xnor U3024 (N_3024,N_1239,N_1110);
xnor U3025 (N_3025,In_1466,In_4654);
nor U3026 (N_3026,N_2459,N_1606);
or U3027 (N_3027,N_1409,In_4353);
xor U3028 (N_3028,In_1362,N_2373);
and U3029 (N_3029,In_2789,N_2277);
or U3030 (N_3030,N_1458,In_634);
xor U3031 (N_3031,N_1532,N_2955);
nand U3032 (N_3032,In_2575,In_2900);
nor U3033 (N_3033,In_1480,N_1552);
xnor U3034 (N_3034,N_2834,N_2406);
or U3035 (N_3035,N_1560,In_1340);
and U3036 (N_3036,N_2892,In_2229);
nor U3037 (N_3037,In_2728,In_3054);
nor U3038 (N_3038,N_2793,N_1470);
and U3039 (N_3039,N_2853,N_1888);
xnor U3040 (N_3040,N_2710,N_490);
nand U3041 (N_3041,N_2139,In_3076);
xor U3042 (N_3042,In_1015,In_2255);
or U3043 (N_3043,N_2732,In_4028);
and U3044 (N_3044,In_996,N_1198);
or U3045 (N_3045,N_2325,In_4769);
xor U3046 (N_3046,N_1573,N_193);
or U3047 (N_3047,N_2641,N_772);
nor U3048 (N_3048,N_2250,In_2134);
and U3049 (N_3049,N_2330,In_2161);
and U3050 (N_3050,N_580,In_3338);
nor U3051 (N_3051,N_1647,In_3505);
or U3052 (N_3052,N_1178,In_3078);
xor U3053 (N_3053,N_390,N_439);
and U3054 (N_3054,N_1493,In_4903);
nand U3055 (N_3055,In_3615,In_4510);
nor U3056 (N_3056,In_238,N_2334);
xor U3057 (N_3057,N_1446,N_2875);
nor U3058 (N_3058,In_3688,N_1736);
xnor U3059 (N_3059,N_127,In_2526);
xnor U3060 (N_3060,N_1188,N_366);
or U3061 (N_3061,In_2478,N_2945);
nand U3062 (N_3062,N_2567,N_208);
xor U3063 (N_3063,In_2998,N_2501);
xor U3064 (N_3064,In_4497,N_2432);
and U3065 (N_3065,N_1908,N_2005);
xnor U3066 (N_3066,N_2389,In_4125);
nand U3067 (N_3067,N_2210,N_1768);
xnor U3068 (N_3068,In_4637,In_1969);
nor U3069 (N_3069,N_2841,N_2169);
nand U3070 (N_3070,N_2566,N_2960);
xnor U3071 (N_3071,In_3610,In_218);
nand U3072 (N_3072,N_245,In_4170);
nand U3073 (N_3073,In_882,In_4100);
nor U3074 (N_3074,N_1357,In_1442);
nor U3075 (N_3075,In_1947,In_1061);
nand U3076 (N_3076,N_2159,N_2624);
and U3077 (N_3077,N_302,In_3286);
nor U3078 (N_3078,In_1361,In_1545);
nor U3079 (N_3079,N_2378,N_1759);
and U3080 (N_3080,N_373,N_2106);
xor U3081 (N_3081,N_1942,In_4597);
nand U3082 (N_3082,N_2614,In_4294);
nor U3083 (N_3083,N_2458,N_2832);
nor U3084 (N_3084,N_2678,In_2731);
or U3085 (N_3085,In_1987,In_1642);
and U3086 (N_3086,N_1896,In_727);
or U3087 (N_3087,N_2164,N_2539);
nor U3088 (N_3088,N_123,In_2632);
xnor U3089 (N_3089,In_2593,N_2986);
nor U3090 (N_3090,In_3655,In_678);
and U3091 (N_3091,In_1247,In_1962);
nor U3092 (N_3092,N_2534,N_269);
or U3093 (N_3093,N_1743,N_1432);
or U3094 (N_3094,In_2591,In_2219);
xnor U3095 (N_3095,In_3836,In_3085);
nand U3096 (N_3096,N_13,N_558);
and U3097 (N_3097,N_1669,In_2202);
and U3098 (N_3098,N_940,In_697);
nand U3099 (N_3099,N_1359,N_2854);
xor U3100 (N_3100,N_2911,N_1914);
xor U3101 (N_3101,N_865,N_2746);
or U3102 (N_3102,In_1633,N_397);
or U3103 (N_3103,N_2901,N_2027);
and U3104 (N_3104,N_1401,N_1764);
nor U3105 (N_3105,N_1336,N_39);
xor U3106 (N_3106,N_2016,N_1289);
and U3107 (N_3107,N_2803,N_2852);
nor U3108 (N_3108,In_4713,In_1496);
xor U3109 (N_3109,N_2931,In_315);
nand U3110 (N_3110,N_1321,In_1471);
and U3111 (N_3111,N_2098,N_2788);
and U3112 (N_3112,N_2921,N_2422);
nand U3113 (N_3113,In_4556,N_2648);
xor U3114 (N_3114,N_2387,In_4563);
and U3115 (N_3115,N_51,N_393);
xor U3116 (N_3116,In_3185,N_956);
nand U3117 (N_3117,N_2655,In_2509);
xor U3118 (N_3118,N_2179,In_178);
nand U3119 (N_3119,N_2636,N_875);
nand U3120 (N_3120,N_2965,N_2452);
nor U3121 (N_3121,In_2501,N_2812);
and U3122 (N_3122,N_2382,N_2868);
or U3123 (N_3123,N_1788,N_1858);
nand U3124 (N_3124,N_2666,N_1102);
and U3125 (N_3125,N_2738,N_2430);
nand U3126 (N_3126,In_362,N_2894);
nand U3127 (N_3127,In_2691,In_4530);
xnor U3128 (N_3128,N_2709,In_3696);
or U3129 (N_3129,N_1388,N_2768);
and U3130 (N_3130,In_2563,N_777);
and U3131 (N_3131,In_3954,In_4889);
nand U3132 (N_3132,N_2994,N_2823);
and U3133 (N_3133,N_94,In_122);
xnor U3134 (N_3134,In_3097,N_345);
nor U3135 (N_3135,N_1886,In_4858);
nand U3136 (N_3136,In_3331,N_2507);
or U3137 (N_3137,N_2014,N_2468);
nand U3138 (N_3138,In_4254,In_1772);
xor U3139 (N_3139,N_2186,In_73);
nand U3140 (N_3140,N_2473,N_2032);
nor U3141 (N_3141,N_1862,N_1509);
nand U3142 (N_3142,N_2905,In_639);
and U3143 (N_3143,N_1118,In_2727);
xnor U3144 (N_3144,In_862,In_3915);
nor U3145 (N_3145,N_2130,N_1672);
xnor U3146 (N_3146,N_1968,N_2398);
or U3147 (N_3147,In_1685,N_2608);
xnor U3148 (N_3148,In_1125,N_2763);
nand U3149 (N_3149,In_468,In_4702);
or U3150 (N_3150,N_2978,N_2521);
and U3151 (N_3151,N_2796,N_2765);
or U3152 (N_3152,N_2226,N_2623);
and U3153 (N_3153,N_1750,In_3811);
or U3154 (N_3154,N_2640,N_2693);
xnor U3155 (N_3155,N_1620,N_871);
or U3156 (N_3156,In_1195,N_1349);
xor U3157 (N_3157,N_2409,In_4084);
and U3158 (N_3158,N_1935,N_1183);
nand U3159 (N_3159,N_2476,N_2393);
nand U3160 (N_3160,N_2837,In_2227);
or U3161 (N_3161,N_2729,In_3791);
xnor U3162 (N_3162,N_2807,In_804);
and U3163 (N_3163,In_2979,N_750);
xnor U3164 (N_3164,N_181,In_4689);
and U3165 (N_3165,N_2415,N_2886);
nor U3166 (N_3166,N_7,In_784);
xnor U3167 (N_3167,N_2010,In_4257);
nand U3168 (N_3168,N_2163,In_4285);
or U3169 (N_3169,In_2844,N_2616);
nor U3170 (N_3170,N_408,In_1936);
and U3171 (N_3171,N_2962,In_348);
nand U3172 (N_3172,N_507,N_2321);
or U3173 (N_3173,N_1006,N_2029);
xnor U3174 (N_3174,N_2946,N_1462);
and U3175 (N_3175,N_2627,N_2547);
nor U3176 (N_3176,In_3709,N_1741);
or U3177 (N_3177,In_3142,In_3038);
nor U3178 (N_3178,In_2960,N_2374);
nor U3179 (N_3179,In_4679,N_2474);
xor U3180 (N_3180,N_2541,N_2433);
xnor U3181 (N_3181,N_2599,In_1757);
or U3182 (N_3182,N_1837,N_2692);
nand U3183 (N_3183,N_2867,N_361);
xnor U3184 (N_3184,N_2772,In_3663);
or U3185 (N_3185,N_1719,In_2732);
nor U3186 (N_3186,In_398,In_4829);
nor U3187 (N_3187,N_2075,N_647);
nand U3188 (N_3188,N_2350,N_2981);
nor U3189 (N_3189,N_2675,N_2705);
xor U3190 (N_3190,In_4016,In_2959);
and U3191 (N_3191,N_1497,N_2869);
xor U3192 (N_3192,N_1779,N_2024);
or U3193 (N_3193,In_1630,In_1040);
xor U3194 (N_3194,N_2778,N_2791);
nor U3195 (N_3195,In_4765,N_2127);
or U3196 (N_3196,N_2753,In_4109);
or U3197 (N_3197,N_720,N_1395);
or U3198 (N_3198,In_28,N_2443);
nor U3199 (N_3199,N_1013,N_2878);
and U3200 (N_3200,N_2445,N_2733);
xnor U3201 (N_3201,N_2067,N_2120);
nand U3202 (N_3202,In_262,In_2874);
nor U3203 (N_3203,In_2718,N_1506);
xnor U3204 (N_3204,In_3492,In_4378);
nor U3205 (N_3205,In_3585,N_2672);
xnor U3206 (N_3206,In_4408,N_2308);
nor U3207 (N_3207,N_2237,N_2882);
and U3208 (N_3208,N_816,In_3717);
and U3209 (N_3209,N_2957,N_2346);
or U3210 (N_3210,N_2972,N_1564);
xnor U3211 (N_3211,In_4899,N_2754);
or U3212 (N_3212,In_2775,N_1652);
xnor U3213 (N_3213,N_1316,In_689);
nand U3214 (N_3214,In_2724,N_467);
xor U3215 (N_3215,In_3578,N_2870);
nor U3216 (N_3216,N_2698,N_1240);
xnor U3217 (N_3217,N_1668,N_2918);
and U3218 (N_3218,N_2034,N_2579);
nor U3219 (N_3219,N_1894,N_2669);
nand U3220 (N_3220,N_2620,N_2684);
nor U3221 (N_3221,N_1360,In_4561);
and U3222 (N_3222,In_4958,N_317);
or U3223 (N_3223,In_3620,N_2076);
or U3224 (N_3224,N_1128,N_1639);
or U3225 (N_3225,N_1069,N_2104);
and U3226 (N_3226,In_1135,N_2799);
and U3227 (N_3227,In_2382,N_2410);
and U3228 (N_3228,N_2708,In_1998);
xnor U3229 (N_3229,N_2591,N_1859);
nor U3230 (N_3230,In_2903,N_1787);
and U3231 (N_3231,In_1755,N_2518);
or U3232 (N_3232,N_2364,In_2329);
and U3233 (N_3233,In_164,In_2966);
and U3234 (N_3234,In_3840,In_1483);
nor U3235 (N_3235,N_2118,N_2950);
nand U3236 (N_3236,N_1000,N_1563);
or U3237 (N_3237,N_1264,N_420);
or U3238 (N_3238,In_4967,In_2171);
xnor U3239 (N_3239,N_693,N_2722);
xor U3240 (N_3240,N_1958,N_2457);
nor U3241 (N_3241,In_3735,N_945);
nand U3242 (N_3242,N_855,In_3971);
nor U3243 (N_3243,In_1791,In_4158);
xor U3244 (N_3244,N_2275,N_2535);
xnor U3245 (N_3245,N_1778,In_2434);
or U3246 (N_3246,N_868,N_207);
nor U3247 (N_3247,In_445,N_2685);
xor U3248 (N_3248,N_2257,N_2699);
and U3249 (N_3249,N_1302,N_2055);
xor U3250 (N_3250,In_4956,N_1124);
or U3251 (N_3251,N_2809,N_3228);
xor U3252 (N_3252,N_2915,N_3032);
nand U3253 (N_3253,N_3212,N_3152);
xor U3254 (N_3254,N_3106,In_4649);
nand U3255 (N_3255,N_2511,N_399);
or U3256 (N_3256,In_603,N_2551);
nand U3257 (N_3257,N_2089,N_2437);
or U3258 (N_3258,N_566,In_874);
and U3259 (N_3259,N_1882,N_1099);
xnor U3260 (N_3260,N_2528,N_3223);
nor U3261 (N_3261,N_3036,In_966);
or U3262 (N_3262,N_3008,N_2563);
nor U3263 (N_3263,N_2366,In_1031);
nand U3264 (N_3264,In_2362,N_3177);
nor U3265 (N_3265,In_4206,N_2414);
nor U3266 (N_3266,N_2776,In_1869);
nand U3267 (N_3267,In_3055,In_193);
or U3268 (N_3268,In_845,In_2643);
nand U3269 (N_3269,In_365,N_2440);
or U3270 (N_3270,In_1351,N_1753);
and U3271 (N_3271,N_2643,N_1592);
nor U3272 (N_3272,N_760,In_3627);
nand U3273 (N_3273,N_3037,N_3035);
or U3274 (N_3274,In_254,In_382);
or U3275 (N_3275,N_2559,N_3017);
or U3276 (N_3276,In_4155,N_1884);
and U3277 (N_3277,N_3163,In_1682);
nor U3278 (N_3278,N_3161,N_2598);
and U3279 (N_3279,In_4037,N_2526);
and U3280 (N_3280,In_620,In_1758);
xnor U3281 (N_3281,N_1915,N_58);
or U3282 (N_3282,N_2674,N_3188);
xnor U3283 (N_3283,N_1381,N_2302);
and U3284 (N_3284,In_4755,N_997);
and U3285 (N_3285,In_4237,In_2647);
nand U3286 (N_3286,N_3085,N_2956);
nand U3287 (N_3287,N_1341,N_2712);
or U3288 (N_3288,N_2260,N_2690);
and U3289 (N_3289,N_2995,N_2795);
nand U3290 (N_3290,N_2977,In_2777);
xor U3291 (N_3291,In_4929,N_3022);
xnor U3292 (N_3292,In_640,N_1367);
nor U3293 (N_3293,N_2922,In_4602);
nor U3294 (N_3294,N_2472,N_2263);
nor U3295 (N_3295,N_70,N_3069);
or U3296 (N_3296,N_3060,N_1733);
and U3297 (N_3297,In_4115,N_2673);
nor U3298 (N_3298,N_2343,N_1187);
nor U3299 (N_3299,N_1450,In_1854);
nand U3300 (N_3300,N_1530,N_2802);
xnor U3301 (N_3301,In_2746,In_1536);
nor U3302 (N_3302,N_2593,In_3554);
or U3303 (N_3303,N_2630,In_4478);
or U3304 (N_3304,In_3040,N_2197);
and U3305 (N_3305,In_3814,N_2213);
nor U3306 (N_3306,N_3142,In_1732);
nand U3307 (N_3307,N_928,In_1284);
nand U3308 (N_3308,N_2199,N_2419);
nand U3309 (N_3309,N_3204,N_2565);
nand U3310 (N_3310,N_3102,In_1465);
nor U3311 (N_3311,N_3211,N_2941);
xnor U3312 (N_3312,In_3601,N_2081);
nor U3313 (N_3313,N_1143,N_2439);
xnor U3314 (N_3314,N_350,N_2128);
and U3315 (N_3315,N_3233,N_2966);
and U3316 (N_3316,In_4854,N_1269);
nor U3317 (N_3317,In_742,N_261);
nand U3318 (N_3318,N_1830,In_3481);
or U3319 (N_3319,N_2843,In_4751);
nand U3320 (N_3320,N_3135,N_1643);
nor U3321 (N_3321,N_1204,N_2423);
or U3322 (N_3322,In_4354,N_3061);
nor U3323 (N_3323,N_1364,N_3227);
nand U3324 (N_3324,In_3715,N_3182);
nand U3325 (N_3325,N_3159,N_962);
nor U3326 (N_3326,In_2343,N_2736);
nor U3327 (N_3327,N_2755,In_63);
nor U3328 (N_3328,N_3206,In_2071);
or U3329 (N_3329,N_1474,N_2811);
xnor U3330 (N_3330,In_1144,N_2060);
nor U3331 (N_3331,In_972,N_1134);
and U3332 (N_3332,In_3349,N_1565);
and U3333 (N_3333,N_2997,In_4365);
xor U3334 (N_3334,In_123,N_1207);
xnor U3335 (N_3335,N_2002,N_2863);
or U3336 (N_3336,N_1997,N_915);
or U3337 (N_3337,N_953,N_3108);
and U3338 (N_3338,N_1794,N_2544);
nand U3339 (N_3339,N_3075,In_4092);
or U3340 (N_3340,In_1825,N_2974);
xnor U3341 (N_3341,In_4876,N_2522);
and U3342 (N_3342,N_1076,N_2855);
xnor U3343 (N_3343,N_3104,N_3098);
nand U3344 (N_3344,In_830,N_3202);
xor U3345 (N_3345,N_3158,N_2819);
or U3346 (N_3346,N_499,In_1542);
and U3347 (N_3347,N_3004,In_2212);
nand U3348 (N_3348,In_4302,N_2622);
and U3349 (N_3349,N_2888,N_3082);
nand U3350 (N_3350,N_3057,N_1844);
nor U3351 (N_3351,N_3055,In_2361);
and U3352 (N_3352,N_3229,In_4463);
nand U3353 (N_3353,N_2919,In_3834);
nand U3354 (N_3354,In_559,In_2216);
and U3355 (N_3355,N_2948,N_2451);
or U3356 (N_3356,N_2975,N_2642);
or U3357 (N_3357,In_3045,In_404);
or U3358 (N_3358,N_1281,N_2810);
nand U3359 (N_3359,N_2466,N_2215);
or U3360 (N_3360,N_2717,N_2225);
xnor U3361 (N_3361,In_3782,In_1626);
nand U3362 (N_3362,N_1758,N_2906);
and U3363 (N_3363,N_134,N_2606);
or U3364 (N_3364,N_881,N_3180);
xnor U3365 (N_3365,N_3215,N_1232);
nand U3366 (N_3366,In_4394,N_3208);
nor U3367 (N_3367,N_2720,N_609);
xor U3368 (N_3368,In_3487,N_1902);
nor U3369 (N_3369,N_2323,In_140);
and U3370 (N_3370,N_2967,N_2943);
nand U3371 (N_3371,In_3677,N_3056);
and U3372 (N_3372,N_2361,In_4098);
and U3373 (N_3373,N_442,In_2745);
and U3374 (N_3374,N_158,N_3101);
xor U3375 (N_3375,N_2848,N_3183);
or U3376 (N_3376,N_2181,In_4381);
nand U3377 (N_3377,N_2644,N_2688);
or U3378 (N_3378,In_3440,N_3007);
and U3379 (N_3379,N_1430,N_2813);
nor U3380 (N_3380,In_1153,N_2756);
nor U3381 (N_3381,In_729,N_2046);
nand U3382 (N_3382,In_1571,N_3155);
xnor U3383 (N_3383,N_2198,N_2897);
or U3384 (N_3384,N_2147,In_2251);
nand U3385 (N_3385,N_2961,N_766);
xnor U3386 (N_3386,N_3238,In_1823);
nand U3387 (N_3387,N_3006,N_1900);
nand U3388 (N_3388,N_289,N_570);
xor U3389 (N_3389,N_1241,In_338);
nor U3390 (N_3390,N_483,In_4687);
nand U3391 (N_3391,N_2801,In_574);
nor U3392 (N_3392,N_3178,In_3697);
nand U3393 (N_3393,N_2979,N_1953);
nor U3394 (N_3394,In_3156,N_2238);
xor U3395 (N_3395,N_2049,In_807);
nand U3396 (N_3396,N_2829,In_1835);
xor U3397 (N_3397,N_2949,N_2980);
and U3398 (N_3398,N_3132,In_4270);
xnor U3399 (N_3399,N_3067,In_3659);
nor U3400 (N_3400,N_3021,N_2564);
xnor U3401 (N_3401,N_3078,In_2783);
and U3402 (N_3402,In_2529,N_668);
nor U3403 (N_3403,In_3965,N_2904);
nor U3404 (N_3404,N_1885,In_3186);
or U3405 (N_3405,N_2221,N_3138);
nand U3406 (N_3406,N_1702,N_2714);
and U3407 (N_3407,N_458,In_3235);
xnor U3408 (N_3408,In_86,N_1176);
nand U3409 (N_3409,N_1623,N_2849);
or U3410 (N_3410,N_1656,N_353);
and U3411 (N_3411,In_1855,In_4508);
and U3412 (N_3412,In_4543,N_2174);
nor U3413 (N_3413,In_660,N_2637);
nand U3414 (N_3414,In_249,N_2984);
nand U3415 (N_3415,In_1004,In_2741);
nand U3416 (N_3416,In_1066,In_2530);
or U3417 (N_3417,N_2706,N_1904);
or U3418 (N_3418,In_592,In_753);
and U3419 (N_3419,N_2447,N_2764);
nor U3420 (N_3420,In_1744,N_2618);
xor U3421 (N_3421,N_2771,N_2490);
xor U3422 (N_3422,N_2844,N_795);
or U3423 (N_3423,In_1689,N_3115);
nor U3424 (N_3424,N_3094,N_1691);
xor U3425 (N_3425,N_994,N_3071);
or U3426 (N_3426,N_3149,N_599);
and U3427 (N_3427,N_658,N_3139);
or U3428 (N_3428,N_553,N_1305);
or U3429 (N_3429,N_1838,N_1843);
xor U3430 (N_3430,N_1723,N_3028);
nand U3431 (N_3431,In_612,N_2893);
xnor U3432 (N_3432,N_2372,In_3394);
nor U3433 (N_3433,In_2040,N_2576);
and U3434 (N_3434,N_1310,N_2814);
xor U3435 (N_3435,N_3168,N_1945);
and U3436 (N_3436,In_1140,In_819);
or U3437 (N_3437,N_2224,N_464);
xnor U3438 (N_3438,N_1248,In_2057);
or U3439 (N_3439,N_718,N_2329);
or U3440 (N_3440,N_866,In_4449);
nor U3441 (N_3441,In_2213,N_1786);
and U3442 (N_3442,N_2944,In_4540);
nand U3443 (N_3443,N_2741,In_1746);
and U3444 (N_3444,N_2066,N_117);
xor U3445 (N_3445,N_2879,N_2319);
and U3446 (N_3446,In_644,In_264);
and U3447 (N_3447,In_2810,N_2917);
or U3448 (N_3448,N_879,In_517);
or U3449 (N_3449,In_2965,N_2968);
or U3450 (N_3450,In_884,N_2947);
and U3451 (N_3451,In_22,N_1536);
nor U3452 (N_3452,In_4681,N_2403);
and U3453 (N_3453,N_3247,N_588);
nand U3454 (N_3454,N_2086,N_3195);
nand U3455 (N_3455,N_2465,N_2998);
and U3456 (N_3456,N_3112,N_1073);
or U3457 (N_3457,In_4136,N_314);
nand U3458 (N_3458,N_1898,N_2073);
nand U3459 (N_3459,In_4538,N_1257);
nor U3460 (N_3460,In_869,In_115);
or U3461 (N_3461,N_2369,N_3058);
nand U3462 (N_3462,In_281,In_4446);
nand U3463 (N_3463,N_3026,N_3077);
nand U3464 (N_3464,N_3073,N_2283);
nand U3465 (N_3465,N_3018,N_1361);
xor U3466 (N_3466,N_2448,In_938);
nor U3467 (N_3467,N_2298,N_3114);
xor U3468 (N_3468,In_3803,N_3024);
nand U3469 (N_3469,In_554,N_2585);
and U3470 (N_3470,N_2484,In_4040);
and U3471 (N_3471,In_4187,N_3092);
and U3472 (N_3472,N_2696,In_4214);
nand U3473 (N_3473,N_1061,In_668);
nand U3474 (N_3474,N_2543,N_1043);
xor U3475 (N_3475,In_1179,N_3173);
nor U3476 (N_3476,N_2486,N_2820);
nor U3477 (N_3477,N_2850,In_4024);
nor U3478 (N_3478,N_2694,N_2580);
and U3479 (N_3479,N_2514,In_928);
and U3480 (N_3480,In_1209,N_1380);
nand U3481 (N_3481,N_2112,N_2881);
xor U3482 (N_3482,N_2652,N_1527);
and U3483 (N_3483,N_607,N_1929);
nor U3484 (N_3484,N_2864,In_4309);
and U3485 (N_3485,In_1844,N_3125);
nor U3486 (N_3486,N_1979,N_1624);
and U3487 (N_3487,N_3096,In_1474);
xor U3488 (N_3488,N_978,N_2281);
nand U3489 (N_3489,N_2327,In_2986);
and U3490 (N_3490,N_2767,N_1823);
xor U3491 (N_3491,In_4535,N_3136);
nand U3492 (N_3492,In_4325,In_1500);
nor U3493 (N_3493,N_1912,N_2099);
nand U3494 (N_3494,In_3295,N_2851);
nor U3495 (N_3495,N_2816,N_1427);
or U3496 (N_3496,In_2269,N_2818);
or U3497 (N_3497,N_3087,N_2248);
nor U3498 (N_3498,N_1400,N_2134);
or U3499 (N_3499,In_1396,In_3876);
or U3500 (N_3500,N_908,In_2923);
xnor U3501 (N_3501,N_3351,N_3249);
nor U3502 (N_3502,In_3298,In_3093);
xnor U3503 (N_3503,N_2607,N_3174);
and U3504 (N_3504,N_2045,N_2018);
or U3505 (N_3505,N_3072,In_4074);
xor U3506 (N_3506,N_3398,N_2455);
and U3507 (N_3507,In_3439,N_2256);
or U3508 (N_3508,N_3042,N_3214);
nand U3509 (N_3509,N_2131,N_3151);
and U3510 (N_3510,N_2148,In_4980);
xor U3511 (N_3511,N_3219,In_2829);
and U3512 (N_3512,In_651,In_4715);
and U3513 (N_3513,N_2273,In_4179);
or U3514 (N_3514,N_2929,In_4205);
and U3515 (N_3515,N_1554,N_1402);
nand U3516 (N_3516,N_64,N_808);
xor U3517 (N_3517,In_2190,N_3235);
nand U3518 (N_3518,N_3435,In_4432);
nor U3519 (N_3519,N_2982,N_3466);
nor U3520 (N_3520,N_796,N_2122);
or U3521 (N_3521,In_890,In_1822);
xnor U3522 (N_3522,N_880,N_2425);
nand U3523 (N_3523,N_2938,In_110);
nand U3524 (N_3524,N_1027,N_2838);
and U3525 (N_3525,N_2650,N_1088);
or U3526 (N_3526,N_2676,N_3209);
xnor U3527 (N_3527,N_2890,N_916);
nor U3528 (N_3528,In_833,N_1115);
nand U3529 (N_3529,In_3084,N_1362);
or U3530 (N_3530,N_2914,N_2068);
nor U3531 (N_3531,N_3424,N_2375);
nand U3532 (N_3532,In_2460,N_3426);
or U3533 (N_3533,N_3105,In_3671);
nor U3534 (N_3534,N_3123,N_3361);
and U3535 (N_3535,N_937,N_3124);
xor U3536 (N_3536,N_3369,N_3310);
and U3537 (N_3537,N_3279,N_1731);
nor U3538 (N_3538,N_3048,N_1977);
or U3539 (N_3539,N_3412,N_2339);
xnor U3540 (N_3540,In_2559,N_3148);
nor U3541 (N_3541,In_2335,N_2681);
nand U3542 (N_3542,N_2822,N_3464);
nor U3543 (N_3543,N_2560,N_1295);
or U3544 (N_3544,N_3416,N_2510);
nand U3545 (N_3545,N_1132,In_886);
xnor U3546 (N_3546,N_2769,N_1033);
xor U3547 (N_3547,N_2600,N_3415);
nand U3548 (N_3548,N_1655,In_1236);
nor U3549 (N_3549,N_3318,In_3988);
or U3550 (N_3550,In_4692,N_2091);
xnor U3551 (N_3551,N_3390,N_3244);
nand U3552 (N_3552,In_4470,In_2936);
and U3553 (N_3553,N_3300,In_4551);
or U3554 (N_3554,N_2610,N_168);
nor U3555 (N_3555,In_472,N_3396);
nand U3556 (N_3556,N_2269,N_814);
xnor U3557 (N_3557,N_2160,N_2156);
nor U3558 (N_3558,N_2185,N_1633);
nand U3559 (N_3559,N_3045,N_1473);
nand U3560 (N_3560,N_1504,In_169);
xnor U3561 (N_3561,N_3270,N_2744);
or U3562 (N_3562,N_2390,N_2462);
nor U3563 (N_3563,In_646,N_2862);
and U3564 (N_3564,In_2554,N_2828);
or U3565 (N_3565,In_4717,N_3425);
xor U3566 (N_3566,In_987,N_3355);
or U3567 (N_3567,In_2751,In_3730);
nor U3568 (N_3568,In_1857,N_3315);
nand U3569 (N_3569,N_1391,N_2773);
nand U3570 (N_3570,N_2524,N_1608);
nand U3571 (N_3571,N_3273,N_2463);
and U3572 (N_3572,In_2205,In_4256);
nor U3573 (N_3573,N_184,In_3981);
or U3574 (N_3574,N_1173,N_2757);
nand U3575 (N_3575,In_2167,N_2554);
or U3576 (N_3576,In_1608,N_328);
and U3577 (N_3577,In_4995,In_513);
or U3578 (N_3578,N_2615,N_2617);
nand U3579 (N_3579,N_2953,N_659);
and U3580 (N_3580,N_1790,N_3401);
and U3581 (N_3581,N_224,N_3483);
or U3582 (N_3582,In_4380,N_3253);
and U3583 (N_3583,N_1127,N_3263);
and U3584 (N_3584,In_1943,In_2663);
and U3585 (N_3585,N_1981,N_2782);
or U3586 (N_3586,N_3378,N_2621);
xor U3587 (N_3587,N_2161,N_2798);
and U3588 (N_3588,N_3288,N_2003);
nand U3589 (N_3589,N_3099,N_3471);
nand U3590 (N_3590,N_3342,In_4457);
or U3591 (N_3591,In_2187,N_2797);
or U3592 (N_3592,In_2295,N_2889);
and U3593 (N_3593,N_2775,N_1934);
nor U3594 (N_3594,N_3472,N_841);
and U3595 (N_3595,N_753,N_1304);
xor U3596 (N_3596,In_4942,N_581);
or U3597 (N_3597,N_276,In_3733);
nand U3598 (N_3598,N_3302,N_2954);
xor U3599 (N_3599,N_2934,N_246);
nor U3600 (N_3600,N_2804,In_2555);
xnor U3601 (N_3601,In_1579,N_120);
nand U3602 (N_3602,N_870,N_3406);
nor U3603 (N_3603,N_1792,N_371);
nor U3604 (N_3604,N_1048,In_824);
nand U3605 (N_3605,N_2983,N_1789);
nor U3606 (N_3606,In_321,In_3219);
nor U3607 (N_3607,N_2891,In_2787);
or U3608 (N_3608,In_449,In_2368);
or U3609 (N_3609,N_441,N_1769);
or U3610 (N_3610,N_2469,In_1900);
or U3611 (N_3611,N_744,N_1921);
xnor U3612 (N_3612,N_3312,N_2172);
or U3613 (N_3613,In_4137,In_1266);
or U3614 (N_3614,N_3344,N_3084);
nor U3615 (N_3615,N_949,N_2603);
nor U3616 (N_3616,In_1089,N_1632);
nor U3617 (N_3617,N_3360,N_3210);
xnor U3618 (N_3618,N_3299,N_1007);
and U3619 (N_3619,N_1301,N_840);
and U3620 (N_3620,N_3399,In_3822);
nand U3621 (N_3621,N_2907,N_2588);
and U3622 (N_3622,N_3493,N_1426);
or U3623 (N_3623,N_3455,N_3276);
xor U3624 (N_3624,N_1216,N_3394);
and U3625 (N_3625,N_3034,N_1051);
or U3626 (N_3626,N_3193,In_631);
nand U3627 (N_3627,N_3167,N_309);
xnor U3628 (N_3628,N_2529,N_2446);
nor U3629 (N_3629,In_23,N_2280);
xor U3630 (N_3630,N_3091,N_2629);
nand U3631 (N_3631,N_2331,N_2958);
and U3632 (N_3632,N_1957,In_3089);
nand U3633 (N_3633,N_3258,N_3070);
nand U3634 (N_3634,N_2845,N_3404);
nand U3635 (N_3635,N_3224,In_703);
xnor U3636 (N_3636,N_3062,In_2785);
nand U3637 (N_3637,In_3766,In_4746);
xnor U3638 (N_3638,N_1578,N_2876);
nand U3639 (N_3639,N_1842,N_590);
nor U3640 (N_3640,N_3012,N_1926);
xor U3641 (N_3641,N_2895,N_3266);
and U3642 (N_3642,N_3086,N_998);
nor U3643 (N_3643,N_3262,In_4771);
xnor U3644 (N_3644,N_2070,In_4916);
and U3645 (N_3645,In_2286,In_1952);
nor U3646 (N_3646,N_31,In_2873);
nand U3647 (N_3647,N_1892,N_3450);
or U3648 (N_3648,In_3194,N_2887);
and U3649 (N_3649,N_1092,N_1828);
or U3650 (N_3650,N_1923,N_3400);
nor U3651 (N_3651,N_1594,N_3475);
nor U3652 (N_3652,N_2976,N_2683);
nand U3653 (N_3653,N_3065,N_1611);
xnor U3654 (N_3654,N_3257,N_130);
and U3655 (N_3655,N_3089,N_2009);
nand U3656 (N_3656,N_1695,N_3088);
nand U3657 (N_3657,N_3278,N_1282);
nand U3658 (N_3658,N_3307,In_3547);
nand U3659 (N_3659,N_2631,N_2925);
and U3660 (N_3660,In_959,N_2146);
nor U3661 (N_3661,N_3079,N_3146);
xor U3662 (N_3662,N_2839,In_4245);
xnor U3663 (N_3663,N_3434,In_1916);
xnor U3664 (N_3664,N_3131,In_433);
or U3665 (N_3665,In_3774,In_4523);
nand U3666 (N_3666,In_1518,N_2391);
or U3667 (N_3667,N_2124,N_1050);
nor U3668 (N_3668,N_3325,In_1531);
nor U3669 (N_3669,N_2503,N_2857);
or U3670 (N_3670,N_3203,N_3050);
xnor U3671 (N_3671,N_1664,N_3457);
and U3672 (N_3672,In_248,N_2750);
nor U3673 (N_3673,N_1507,In_3424);
or U3674 (N_3674,N_3119,In_1702);
nand U3675 (N_3675,N_3081,In_2709);
xor U3676 (N_3676,N_372,N_3009);
and U3677 (N_3677,N_1037,In_2340);
and U3678 (N_3678,N_3063,In_3905);
nand U3679 (N_3679,N_147,In_163);
xnor U3680 (N_3680,N_3109,N_3372);
and U3681 (N_3681,N_1350,In_347);
xor U3682 (N_3682,N_2515,In_3600);
xnor U3683 (N_3683,N_3480,N_2991);
nor U3684 (N_3684,N_1202,N_3144);
or U3685 (N_3685,N_1406,N_3341);
xnor U3686 (N_3686,N_326,In_2857);
nor U3687 (N_3687,In_3573,N_2628);
nand U3688 (N_3688,In_4782,N_2899);
xnor U3689 (N_3689,In_502,N_2815);
or U3690 (N_3690,N_3120,N_3349);
nand U3691 (N_3691,In_770,In_2110);
nor U3692 (N_3692,N_308,N_2117);
xnor U3693 (N_3693,N_3237,N_3156);
or U3694 (N_3694,N_1249,N_2240);
and U3695 (N_3695,N_3165,N_3001);
xor U3696 (N_3696,N_3126,N_2735);
nor U3697 (N_3697,In_669,N_2959);
nor U3698 (N_3698,N_1971,N_1108);
xnor U3699 (N_3699,In_2633,N_3040);
and U3700 (N_3700,N_2670,N_3377);
and U3701 (N_3701,N_453,N_505);
xor U3702 (N_3702,N_2504,N_2318);
or U3703 (N_3703,N_2910,N_3494);
and U3704 (N_3704,N_2660,N_2865);
or U3705 (N_3705,N_2096,N_1101);
xnor U3706 (N_3706,In_923,N_1936);
xnor U3707 (N_3707,N_3268,N_3166);
xor U3708 (N_3708,N_2695,N_3417);
nand U3709 (N_3709,N_2053,N_2499);
or U3710 (N_3710,In_731,N_2531);
and U3711 (N_3711,In_1999,N_3334);
and U3712 (N_3712,N_2786,In_490);
nand U3713 (N_3713,N_1286,In_4812);
xnor U3714 (N_3714,N_3287,In_3809);
nand U3715 (N_3715,N_1897,N_1196);
or U3716 (N_3716,N_2840,N_3470);
xnor U3717 (N_3717,In_924,N_2989);
xor U3718 (N_3718,In_2347,N_2058);
and U3719 (N_3719,N_2111,N_2992);
nand U3720 (N_3720,In_4731,N_2779);
xor U3721 (N_3721,N_16,N_2902);
and U3722 (N_3722,In_3695,N_2376);
and U3723 (N_3723,N_2766,In_3759);
nand U3724 (N_3724,N_2063,In_4630);
xor U3725 (N_3725,N_2745,In_1422);
or U3726 (N_3726,N_2491,N_3442);
or U3727 (N_3727,In_4211,N_1745);
and U3728 (N_3728,In_260,N_2703);
xor U3729 (N_3729,N_1408,N_2777);
xnor U3730 (N_3730,In_4420,In_4528);
nand U3731 (N_3731,N_3191,In_4846);
nor U3732 (N_3732,N_2609,N_1781);
xor U3733 (N_3733,N_3169,N_3052);
nand U3734 (N_3734,In_2683,N_2562);
and U3735 (N_3735,N_2384,N_2612);
xor U3736 (N_3736,N_2903,N_2940);
xor U3737 (N_3737,N_2935,N_2734);
nand U3738 (N_3738,N_786,N_2752);
nor U3739 (N_3739,In_3913,In_335);
and U3740 (N_3740,N_2371,In_2253);
or U3741 (N_3741,N_3345,N_2353);
xnor U3742 (N_3742,N_2336,N_2781);
nand U3743 (N_3743,N_2532,N_3137);
xor U3744 (N_3744,N_3083,N_3130);
or U3745 (N_3745,N_2721,N_3025);
nand U3746 (N_3746,N_3236,N_3389);
and U3747 (N_3747,In_3330,N_3486);
or U3748 (N_3748,N_3051,N_2328);
xor U3749 (N_3749,N_3469,N_1670);
or U3750 (N_3750,N_2831,N_3566);
and U3751 (N_3751,In_2870,N_2429);
or U3752 (N_3752,In_4698,N_3582);
nand U3753 (N_3753,N_3648,N_3205);
nand U3754 (N_3754,N_2885,In_997);
and U3755 (N_3755,N_2271,N_1253);
nor U3756 (N_3756,In_1027,N_1662);
xnor U3757 (N_3757,N_2552,N_1179);
nand U3758 (N_3758,In_1889,N_2740);
or U3759 (N_3759,N_554,N_2794);
and U3760 (N_3760,N_3175,N_3500);
or U3761 (N_3761,N_3107,In_4776);
and U3762 (N_3762,In_2660,N_1583);
and U3763 (N_3763,N_1797,In_1048);
xor U3764 (N_3764,N_3461,N_2402);
nand U3765 (N_3765,N_175,In_3543);
nand U3766 (N_3766,In_1202,N_3327);
and U3767 (N_3767,N_3368,In_1400);
nand U3768 (N_3768,N_3199,N_3141);
and U3769 (N_3769,N_3277,In_2671);
nand U3770 (N_3770,In_3720,N_3735);
and U3771 (N_3771,N_2355,N_1951);
nand U3772 (N_3772,In_4112,In_1899);
xor U3773 (N_3773,N_3029,N_3283);
xor U3774 (N_3774,In_2443,N_3340);
nor U3775 (N_3775,N_1487,N_3516);
xnor U3776 (N_3776,In_4896,N_724);
and U3777 (N_3777,In_2230,N_3452);
and U3778 (N_3778,N_1744,N_3644);
nand U3779 (N_3779,In_911,N_3023);
nor U3780 (N_3780,N_3696,N_3561);
nand U3781 (N_3781,N_2556,N_3314);
nor U3782 (N_3782,N_3328,In_1740);
xnor U3783 (N_3783,N_2817,N_2506);
xnor U3784 (N_3784,N_2266,N_2300);
nor U3785 (N_3785,N_3709,In_76);
or U3786 (N_3786,N_3700,In_1574);
xnor U3787 (N_3787,N_2952,N_2639);
and U3788 (N_3788,N_2987,N_1681);
xnor U3789 (N_3789,N_3690,N_1534);
and U3790 (N_3790,In_3391,N_318);
nor U3791 (N_3791,N_2920,N_3076);
or U3792 (N_3792,N_2898,In_4376);
xnor U3793 (N_3793,In_4526,N_1982);
nor U3794 (N_3794,N_3440,In_208);
and U3795 (N_3795,N_2324,N_3100);
xnor U3796 (N_3796,N_616,N_3405);
xor U3797 (N_3797,N_3620,N_3323);
or U3798 (N_3798,N_3733,N_2700);
nor U3799 (N_3799,N_3259,N_3190);
nand U3800 (N_3800,N_3544,In_1709);
nor U3801 (N_3801,N_3720,N_2496);
nor U3802 (N_3802,N_1766,In_2488);
and U3803 (N_3803,N_2397,N_3393);
nor U3804 (N_3804,In_1533,In_4973);
nor U3805 (N_3805,N_3683,N_1220);
or U3806 (N_3806,N_2662,N_2846);
xnor U3807 (N_3807,N_2680,N_3090);
or U3808 (N_3808,N_2488,N_3617);
xnor U3809 (N_3809,N_3316,N_3632);
and U3810 (N_3810,N_2806,N_3386);
nand U3811 (N_3811,N_2290,N_2939);
nor U3812 (N_3812,N_3702,In_125);
nand U3813 (N_3813,N_3664,N_1822);
xor U3814 (N_3814,N_3520,In_3923);
xor U3815 (N_3815,In_2375,In_2186);
or U3816 (N_3816,N_1292,N_150);
xor U3817 (N_3817,N_3011,N_3489);
and U3818 (N_3818,In_1592,N_1492);
and U3819 (N_3819,N_3395,N_3511);
and U3820 (N_3820,N_3605,N_3311);
nor U3821 (N_3821,N_3482,N_1805);
or U3822 (N_3822,N_3103,N_3463);
nand U3823 (N_3823,N_3038,N_1829);
xor U3824 (N_3824,N_3459,N_3286);
xor U3825 (N_3825,N_2590,In_1655);
or U3826 (N_3826,N_2288,In_971);
nor U3827 (N_3827,In_3940,In_4011);
and U3828 (N_3828,In_3532,N_3557);
or U3829 (N_3829,N_3451,N_3588);
nand U3830 (N_3830,In_4611,N_3294);
nor U3831 (N_3831,N_1418,N_3290);
or U3832 (N_3832,In_4673,N_3539);
nor U3833 (N_3833,In_2464,N_1810);
nor U3834 (N_3834,N_3226,N_1211);
nor U3835 (N_3835,N_3655,N_1475);
or U3836 (N_3836,N_1752,N_3491);
or U3837 (N_3837,In_4695,N_3422);
and U3838 (N_3838,In_2907,N_2007);
xor U3839 (N_3839,N_3473,In_2074);
nand U3840 (N_3840,N_1129,N_842);
and U3841 (N_3841,N_2739,N_1984);
nand U3842 (N_3842,In_183,N_3651);
nor U3843 (N_3843,N_2272,N_3337);
or U3844 (N_3844,N_3250,N_3242);
or U3845 (N_3845,In_2311,N_2659);
nor U3846 (N_3846,N_3677,N_3689);
or U3847 (N_3847,In_3202,In_354);
nand U3848 (N_3848,N_2789,In_4985);
xnor U3849 (N_3849,N_1535,N_1696);
or U3850 (N_3850,N_1177,In_602);
nor U3851 (N_3851,N_3506,N_2478);
xnor U3852 (N_3852,N_2527,N_280);
and U3853 (N_3853,N_3589,In_1121);
nor U3854 (N_3854,In_1220,N_2517);
and U3855 (N_3855,N_3343,N_3591);
nand U3856 (N_3856,N_3667,N_2558);
or U3857 (N_3857,N_1682,N_2988);
nand U3858 (N_3858,N_3725,N_1444);
or U3859 (N_3859,N_2317,N_3111);
and U3860 (N_3860,N_2549,In_2148);
and U3861 (N_3861,N_3728,In_3029);
nor U3862 (N_3862,N_3066,N_3255);
and U3863 (N_3863,N_2253,N_3718);
or U3864 (N_3864,N_3681,N_1659);
xor U3865 (N_3865,In_2401,N_3746);
or U3866 (N_3866,In_3740,In_3165);
or U3867 (N_3867,N_938,N_3338);
nor U3868 (N_3868,N_3552,N_3678);
xor U3869 (N_3869,N_3306,N_3738);
nand U3870 (N_3870,In_617,N_3584);
and U3871 (N_3871,In_4861,In_4901);
or U3872 (N_3872,N_3317,N_3367);
or U3873 (N_3873,N_3635,N_3420);
xor U3874 (N_3874,N_3624,In_1907);
and U3875 (N_3875,N_2702,In_2772);
nand U3876 (N_3876,N_2006,In_3921);
xor U3877 (N_3877,N_3484,N_3503);
nor U3878 (N_3878,N_2704,N_1919);
nand U3879 (N_3879,N_3385,N_2866);
and U3880 (N_3880,N_476,N_3737);
nand U3881 (N_3881,N_3613,N_3411);
xnor U3882 (N_3882,N_135,N_1677);
or U3883 (N_3883,N_2596,N_3336);
nand U3884 (N_3884,N_3623,N_3269);
and U3885 (N_3885,In_496,N_2759);
and U3886 (N_3886,N_2399,N_3356);
or U3887 (N_3887,In_4606,N_3636);
and U3888 (N_3888,In_1898,N_2379);
xor U3889 (N_3889,N_2912,N_3402);
and U3890 (N_3890,N_3134,N_2482);
xnor U3891 (N_3891,N_3658,In_3631);
nor U3892 (N_3892,N_3380,N_3660);
nand U3893 (N_3893,N_1686,N_907);
and U3894 (N_3894,N_3694,N_2586);
xnor U3895 (N_3895,N_3333,N_3267);
nor U3896 (N_3896,N_3548,N_3682);
nor U3897 (N_3897,N_3668,N_1856);
nand U3898 (N_3898,N_2619,N_3736);
nand U3899 (N_3899,N_2431,N_3616);
xnor U3900 (N_3900,N_3436,N_2937);
and U3901 (N_3901,N_3409,N_3705);
xor U3902 (N_3902,N_3630,N_745);
nor U3903 (N_3903,N_3672,In_2181);
nand U3904 (N_3904,N_3245,In_1243);
xor U3905 (N_3905,N_2877,N_129);
nor U3906 (N_3906,N_3467,N_2217);
and U3907 (N_3907,N_3514,N_3734);
and U3908 (N_3908,In_3681,N_3614);
nor U3909 (N_3909,N_3397,N_3731);
nand U3910 (N_3910,N_2555,N_2743);
xnor U3911 (N_3911,N_2985,In_1012);
nor U3912 (N_3912,In_1403,N_2587);
or U3913 (N_3913,N_3441,N_2930);
nand U3914 (N_3914,N_2012,N_3282);
nor U3915 (N_3915,N_3241,N_3421);
or U3916 (N_3916,N_634,In_1095);
nor U3917 (N_3917,N_3575,In_2490);
and U3918 (N_3918,N_3453,N_2102);
xor U3919 (N_3919,N_1059,N_3408);
and U3920 (N_3920,N_3507,N_3715);
xnor U3921 (N_3921,N_3454,In_1562);
and U3922 (N_3922,In_4054,N_2170);
and U3923 (N_3923,In_3512,N_2827);
or U3924 (N_3924,N_533,N_1191);
and U3925 (N_3925,N_695,N_1863);
xnor U3926 (N_3926,N_3438,N_1941);
or U3927 (N_3927,N_2783,N_3528);
nand U3928 (N_3928,N_3639,N_1721);
nand U3929 (N_3929,N_3534,N_2206);
and U3930 (N_3930,In_2448,In_4895);
xnor U3931 (N_3931,N_3362,N_2909);
nand U3932 (N_3932,In_2090,N_3540);
xor U3933 (N_3933,N_3221,In_3366);
or U3934 (N_3934,N_3626,N_2360);
or U3935 (N_3935,N_3329,In_895);
nand U3936 (N_3936,In_4799,N_3261);
xnor U3937 (N_3937,N_3304,N_3350);
and U3938 (N_3938,In_3448,In_3451);
or U3939 (N_3939,In_256,In_1929);
or U3940 (N_3940,N_3631,N_1306);
and U3941 (N_3941,In_4055,N_2916);
nand U3942 (N_3942,N_3216,N_3357);
and U3943 (N_3943,In_2041,In_2371);
or U3944 (N_3944,In_976,N_3599);
nand U3945 (N_3945,N_3381,In_2876);
or U3946 (N_3946,N_762,N_3301);
or U3947 (N_3947,N_3176,N_3496);
xor U3948 (N_3948,In_3522,N_2188);
and U3949 (N_3949,N_2602,N_2626);
nor U3950 (N_3950,N_3522,N_3376);
nor U3951 (N_3951,In_906,N_3596);
xnor U3952 (N_3952,In_4452,N_2595);
xnor U3953 (N_3953,In_4984,N_3546);
xor U3954 (N_3954,In_31,N_3370);
and U3955 (N_3955,N_3320,N_1038);
or U3956 (N_3956,N_2926,N_3392);
and U3957 (N_3957,N_2728,N_3117);
and U3958 (N_3958,N_2017,N_1233);
xnor U3959 (N_3959,N_3558,N_1783);
nand U3960 (N_3960,In_2406,N_3456);
nand U3961 (N_3961,In_908,N_3629);
xor U3962 (N_3962,N_1511,N_2475);
xor U3963 (N_3963,N_2993,N_3140);
xnor U3964 (N_3964,N_3147,N_3704);
nand U3965 (N_3965,N_2701,N_3384);
nor U3966 (N_3966,N_3688,In_2327);
nor U3967 (N_3967,In_3152,N_2246);
xnor U3968 (N_3968,N_2900,N_3730);
nand U3969 (N_3969,N_3128,N_3207);
xor U3970 (N_3970,N_3578,N_3192);
or U3971 (N_3971,N_2671,N_2351);
nor U3972 (N_3972,N_2883,N_2191);
and U3973 (N_3973,N_3527,N_3674);
or U3974 (N_3974,In_4326,N_3563);
xnor U3975 (N_3975,N_3429,N_1428);
nand U3976 (N_3976,N_2686,N_2923);
xnor U3977 (N_3977,In_2524,N_2420);
nand U3978 (N_3978,N_3324,N_3280);
and U3979 (N_3979,N_3181,N_3252);
and U3980 (N_3980,N_3427,In_1008);
or U3981 (N_3981,N_2942,N_3594);
or U3982 (N_3982,N_2356,N_3121);
and U3983 (N_3983,N_2667,N_3059);
or U3984 (N_3984,N_2365,N_2212);
nand U3985 (N_3985,In_905,In_4627);
nand U3986 (N_3986,N_1488,N_1854);
nor U3987 (N_3987,In_4922,N_1996);
nand U3988 (N_3988,N_3621,N_2718);
and U3989 (N_3989,N_2326,N_2825);
nand U3990 (N_3990,In_1619,N_2123);
and U3991 (N_3991,N_3271,N_1959);
nor U3992 (N_3992,N_3010,N_3413);
or U3993 (N_3993,N_3364,N_3382);
xnor U3994 (N_3994,N_3033,In_3116);
or U3995 (N_3995,N_3519,In_4655);
xor U3996 (N_3996,N_3447,In_4798);
nor U3997 (N_3997,N_3749,N_1114);
nor U3998 (N_3998,N_3495,In_3925);
and U3999 (N_3999,N_3662,N_3653);
nor U4000 (N_4000,N_3951,N_3964);
nand U4001 (N_4001,N_2668,N_365);
xor U4002 (N_4002,N_2173,N_1343);
or U4003 (N_4003,N_61,In_3153);
nand U4004 (N_4004,N_1285,N_3764);
or U4005 (N_4005,N_3220,N_3110);
nand U4006 (N_4006,N_2533,N_3281);
and U4007 (N_4007,N_3650,N_3526);
or U4008 (N_4008,N_3902,N_3721);
or U4009 (N_4009,In_3325,N_3864);
nand U4010 (N_4010,N_3592,N_3637);
or U4011 (N_4011,N_3217,N_2761);
nand U4012 (N_4012,N_3887,N_3497);
and U4013 (N_4013,N_3999,In_2969);
xor U4014 (N_4014,N_2658,N_2697);
or U4015 (N_4015,N_3722,N_3837);
nand U4016 (N_4016,N_2495,N_3371);
or U4017 (N_4017,N_3153,In_1951);
or U4018 (N_4018,N_3988,N_1413);
nand U4019 (N_4019,N_3877,N_3982);
or U4020 (N_4020,N_3905,N_3602);
nor U4021 (N_4021,N_3788,In_326);
and U4022 (N_4022,N_3305,In_2573);
xnor U4023 (N_4023,N_290,N_2001);
nand U4024 (N_4024,N_2557,N_1646);
xnor U4025 (N_4025,In_3335,N_3583);
and U4026 (N_4026,N_2150,N_3914);
xnor U4027 (N_4027,N_3828,N_3858);
nand U4028 (N_4028,N_1944,N_3911);
or U4029 (N_4029,In_2910,N_3809);
or U4030 (N_4030,N_3831,N_3418);
nor U4031 (N_4031,In_2626,N_1650);
or U4032 (N_4032,N_3595,N_1252);
or U4033 (N_4033,N_3150,N_3231);
or U4034 (N_4034,In_700,N_3816);
xor U4035 (N_4035,N_3953,In_3725);
nand U4036 (N_4036,N_2872,N_2489);
nor U4037 (N_4037,In_4250,N_3889);
nor U4038 (N_4038,N_3388,N_3600);
nor U4039 (N_4039,N_3555,N_3846);
nor U4040 (N_4040,N_3541,N_2546);
xor U4041 (N_4041,In_550,N_694);
nor U4042 (N_4042,N_3691,N_3882);
xor U4043 (N_4043,N_2836,N_3937);
and U4044 (N_4044,N_791,N_3646);
nand U4045 (N_4045,N_3625,In_3465);
nand U4046 (N_4046,N_3912,N_3423);
xnor U4047 (N_4047,N_3847,N_2711);
nand U4048 (N_4048,N_3884,In_1312);
or U4049 (N_4049,N_3995,N_3363);
and U4050 (N_4050,N_3145,N_2026);
or U4051 (N_4051,N_3900,N_3710);
and U4052 (N_4052,N_2969,N_2404);
xor U4053 (N_4053,N_3003,In_2604);
xnor U4054 (N_4054,N_3488,N_3732);
or U4055 (N_4055,In_2089,N_2635);
and U4056 (N_4056,N_3755,N_3777);
nand U4057 (N_4057,N_3821,N_2062);
nor U4058 (N_4058,N_3989,N_3127);
nor U4059 (N_4059,In_4194,N_400);
xnor U4060 (N_4060,N_3654,N_2824);
and U4061 (N_4061,N_2145,In_4727);
or U4062 (N_4062,N_3043,N_967);
nand U4063 (N_4063,In_1603,N_3761);
nor U4064 (N_4064,N_2780,N_3538);
nor U4065 (N_4065,N_3941,N_3551);
nand U4066 (N_4066,In_1485,N_3232);
nor U4067 (N_4067,N_3936,N_3610);
xor U4068 (N_4068,In_4785,N_3509);
nand U4069 (N_4069,N_2502,In_4851);
or U4070 (N_4070,N_3772,N_3529);
nor U4071 (N_4071,N_3387,In_2126);
and U4072 (N_4072,N_3666,N_1287);
or U4073 (N_4073,N_3194,N_876);
xor U4074 (N_4074,N_3000,N_3049);
nand U4075 (N_4075,N_3874,N_3502);
nand U4076 (N_4076,N_3792,N_1835);
xnor U4077 (N_4077,N_3535,N_3765);
nand U4078 (N_4078,N_3771,In_1199);
xor U4079 (N_4079,In_3870,In_1181);
nor U4080 (N_4080,In_1149,N_3627);
and U4081 (N_4081,N_1184,N_3292);
and U4082 (N_4082,N_3955,N_3414);
nand U4083 (N_4083,N_3603,In_674);
xnor U4084 (N_4084,In_3494,N_3570);
and U4085 (N_4085,In_4070,N_3814);
or U4086 (N_4086,N_3685,N_1550);
xor U4087 (N_4087,N_2856,N_3196);
nand U4088 (N_4088,N_3501,N_2833);
and U4089 (N_4089,In_1918,N_3850);
nand U4090 (N_4090,N_2289,N_635);
nor U4091 (N_4091,N_3553,N_2135);
or U4092 (N_4092,N_1420,N_3322);
and U4093 (N_4093,N_3498,N_838);
nand U4094 (N_4094,N_1303,N_1663);
xor U4095 (N_4095,N_3713,N_3604);
or U4096 (N_4096,N_3876,N_395);
nor U4097 (N_4097,N_3524,N_3918);
or U4098 (N_4098,In_2549,N_3687);
xor U4099 (N_4099,N_3712,N_2581);
and U4100 (N_4100,In_4938,In_4987);
nand U4101 (N_4101,N_1703,N_1298);
nor U4102 (N_4102,N_3867,N_3606);
nand U4103 (N_4103,In_1234,In_1621);
nor U4104 (N_4104,N_3113,N_416);
nor U4105 (N_4105,N_3444,In_1572);
nor U4106 (N_4106,N_3778,N_3985);
and U4107 (N_4107,N_2826,N_3836);
or U4108 (N_4108,N_2358,N_3767);
nor U4109 (N_4109,In_49,N_3807);
nor U4110 (N_4110,N_3848,N_2748);
xnor U4111 (N_4111,N_1757,N_2342);
nor U4112 (N_4112,N_3934,N_859);
nand U4113 (N_4113,N_3295,N_3948);
xor U4114 (N_4114,In_497,N_3275);
or U4115 (N_4115,N_2913,N_3796);
nor U4116 (N_4116,N_2792,N_3726);
nor U4117 (N_4117,N_3762,N_3642);
nand U4118 (N_4118,N_3893,N_3946);
xnor U4119 (N_4119,N_3886,N_3485);
xor U4120 (N_4120,N_3643,In_1965);
and U4121 (N_4121,N_3201,N_3118);
and U4122 (N_4122,N_3272,N_857);
nor U4123 (N_4123,N_2337,N_3987);
and U4124 (N_4124,N_3359,In_834);
and U4125 (N_4125,N_1755,N_3309);
xnor U4126 (N_4126,In_3407,N_3407);
xor U4127 (N_4127,In_2569,N_2178);
nand U4128 (N_4128,N_2109,In_1581);
and U4129 (N_4129,N_2758,N_3213);
nor U4130 (N_4130,N_3699,In_4570);
nand U4131 (N_4131,N_3554,N_3716);
and U4132 (N_4132,N_2871,N_3326);
nand U4133 (N_4133,N_3790,N_2381);
and U4134 (N_4134,N_1424,N_3590);
and U4135 (N_4135,N_3031,In_1375);
xnor U4136 (N_4136,N_3053,N_3160);
and U4137 (N_4137,N_3419,N_1500);
and U4138 (N_4138,N_3717,N_3824);
nor U4139 (N_4139,N_3701,N_3907);
nand U4140 (N_4140,N_2858,N_2183);
nand U4141 (N_4141,N_3296,N_1515);
nand U4142 (N_4142,N_3564,N_2990);
xor U4143 (N_4143,N_3339,N_3931);
nor U4144 (N_4144,N_3559,N_2936);
xor U4145 (N_4145,N_3791,N_1309);
xor U4146 (N_4146,N_2656,N_3775);
xor U4147 (N_4147,N_3901,N_3675);
xnor U4148 (N_4148,N_2345,N_3898);
xnor U4149 (N_4149,N_2589,In_34);
nand U4150 (N_4150,N_3517,N_3248);
or U4151 (N_4151,N_3913,N_3983);
or U4152 (N_4152,In_3357,N_3358);
xnor U4153 (N_4153,In_1953,N_3994);
nor U4154 (N_4154,N_2251,N_3823);
xor U4155 (N_4155,N_2785,In_4594);
xnor U4156 (N_4156,N_3243,N_3291);
xor U4157 (N_4157,N_539,N_3162);
nor U4158 (N_4158,N_3403,N_3975);
or U4159 (N_4159,In_2535,In_2300);
nor U4160 (N_4160,In_2164,In_3173);
or U4161 (N_4161,N_3862,N_3064);
or U4162 (N_4162,N_3543,N_459);
nor U4163 (N_4163,N_1161,N_3921);
nand U4164 (N_4164,N_3303,N_3477);
nand U4165 (N_4165,N_3189,N_244);
nand U4166 (N_4166,N_2229,In_2195);
xor U4167 (N_4167,N_3465,N_2634);
xnor U4168 (N_4168,N_3759,N_2933);
xor U4169 (N_4169,N_3963,N_349);
or U4170 (N_4170,N_2808,N_3133);
nand U4171 (N_4171,N_3926,N_3871);
xor U4172 (N_4172,In_1338,N_3751);
nand U4173 (N_4173,N_1553,In_3617);
or U4174 (N_4174,N_3899,N_3569);
xor U4175 (N_4175,N_3944,N_3225);
and U4176 (N_4176,N_2505,N_3973);
or U4177 (N_4177,In_198,N_3885);
and U4178 (N_4178,N_822,N_3872);
nand U4179 (N_4179,N_1087,N_3910);
and U4180 (N_4180,N_3873,In_3711);
xnor U4181 (N_4181,N_1961,N_2467);
or U4182 (N_4182,N_3962,In_2766);
and U4183 (N_4183,In_1079,N_511);
and U4184 (N_4184,N_3817,N_3492);
or U4185 (N_4185,N_3861,N_3164);
xnor U4186 (N_4186,N_3352,N_3852);
nor U4187 (N_4187,In_4793,N_3976);
nor U4188 (N_4188,N_3757,N_3256);
or U4189 (N_4189,N_2460,N_1484);
nor U4190 (N_4190,N_3825,N_3428);
and U4191 (N_4191,N_3187,N_3014);
nor U4192 (N_4192,N_3532,In_743);
and U4193 (N_4193,N_3857,N_3330);
xor U4194 (N_4194,N_3609,N_2540);
nor U4195 (N_4195,N_3686,In_138);
and U4196 (N_4196,N_3573,N_2605);
or U4197 (N_4197,N_348,N_3891);
nor U4198 (N_4198,N_2464,In_3990);
or U4199 (N_4199,N_3835,N_3537);
or U4200 (N_4200,N_3968,N_3947);
nor U4201 (N_4201,N_3766,In_2867);
nor U4202 (N_4202,N_3916,N_298);
or U4203 (N_4203,N_3978,N_3285);
or U4204 (N_4204,In_3824,N_3806);
nand U4205 (N_4205,N_3875,In_3956);
nand U4206 (N_4206,N_3608,N_3793);
xor U4207 (N_4207,N_3601,N_3919);
xor U4208 (N_4208,In_3948,In_1319);
or U4209 (N_4209,In_3193,N_3618);
nor U4210 (N_4210,N_674,N_3826);
xnor U4211 (N_4211,N_338,N_3179);
nand U4212 (N_4212,In_1233,N_1756);
xnor U4213 (N_4213,N_3980,N_202);
nor U4214 (N_4214,N_3996,N_3745);
nor U4215 (N_4215,N_3549,N_3878);
nand U4216 (N_4216,N_3839,In_4704);
nand U4217 (N_4217,In_3592,N_438);
and U4218 (N_4218,N_3044,N_3903);
and U4219 (N_4219,N_645,N_2963);
nand U4220 (N_4220,N_3365,N_3840);
nor U4221 (N_4221,N_3849,N_3641);
nand U4222 (N_4222,In_866,N_3016);
nand U4223 (N_4223,In_2054,N_3958);
and U4224 (N_4224,N_3783,N_3562);
nor U4225 (N_4225,In_2244,N_3523);
and U4226 (N_4226,N_3347,N_3246);
and U4227 (N_4227,N_3866,N_1366);
xor U4228 (N_4228,In_1013,N_996);
nor U4229 (N_4229,In_4676,N_153);
nor U4230 (N_4230,N_1644,N_3822);
or U4231 (N_4231,In_2618,N_2307);
xor U4232 (N_4232,N_3449,N_3593);
nor U4233 (N_4233,N_3753,N_1323);
nor U4234 (N_4234,N_2095,N_782);
nor U4235 (N_4235,N_1519,N_3954);
nand U4236 (N_4236,N_3046,In_295);
and U4237 (N_4237,N_3993,N_3986);
nand U4238 (N_4238,N_3068,N_3615);
nor U4239 (N_4239,N_3530,N_3254);
or U4240 (N_4240,N_1660,N_3634);
nor U4241 (N_4241,In_4803,N_3928);
nor U4242 (N_4242,N_3758,N_3927);
nand U4243 (N_4243,N_488,N_3820);
nor U4244 (N_4244,N_3446,N_2234);
or U4245 (N_4245,In_3387,In_3035);
nor U4246 (N_4246,N_2519,N_3391);
nor U4247 (N_4247,N_3284,N_3740);
nor U4248 (N_4248,N_3027,N_3794);
xor U4249 (N_4249,N_3935,N_3499);
xor U4250 (N_4250,N_2471,N_4033);
xnor U4251 (N_4251,N_3054,In_4374);
xnor U4252 (N_4252,N_2048,N_3895);
or U4253 (N_4253,N_3448,N_2908);
xnor U4254 (N_4254,N_4066,N_1928);
or U4255 (N_4255,N_4048,N_4051);
and U4256 (N_4256,N_4050,N_4177);
nand U4257 (N_4257,N_1243,N_3780);
nor U4258 (N_4258,N_4070,N_3774);
or U4259 (N_4259,N_4133,N_4170);
nand U4260 (N_4260,N_2285,N_4014);
and U4261 (N_4261,In_1227,N_835);
and U4262 (N_4262,N_3956,N_3917);
xnor U4263 (N_4263,N_2553,In_4969);
and U4264 (N_4264,N_3545,N_3513);
nand U4265 (N_4265,In_378,N_4139);
and U4266 (N_4266,In_4433,N_3800);
xnor U4267 (N_4267,N_2762,N_4166);
nor U4268 (N_4268,N_3829,In_1173);
xor U4269 (N_4269,N_3714,N_4049);
nand U4270 (N_4270,N_3586,N_3727);
xor U4271 (N_4271,N_4245,N_3550);
xnor U4272 (N_4272,N_4192,N_3708);
nand U4273 (N_4273,N_3776,N_4005);
and U4274 (N_4274,N_4195,N_1028);
nand U4275 (N_4275,N_3143,N_3533);
nand U4276 (N_4276,N_4025,N_4161);
and U4277 (N_4277,N_3542,N_3904);
nand U4278 (N_4278,N_4090,N_3628);
xnor U4279 (N_4279,N_4168,In_2445);
and U4280 (N_4280,N_3510,N_3801);
nor U4281 (N_4281,N_4078,N_4234);
xnor U4282 (N_4282,N_3784,N_4167);
nand U4283 (N_4283,In_1534,N_4221);
xor U4284 (N_4284,N_4147,In_4718);
or U4285 (N_4285,N_4043,N_3515);
and U4286 (N_4286,N_4185,In_4578);
xnor U4287 (N_4287,N_3692,N_1226);
or U4288 (N_4288,N_1603,N_3965);
xnor U4289 (N_4289,N_3585,In_3998);
or U4290 (N_4290,N_3789,N_4179);
xnor U4291 (N_4291,N_3785,N_4013);
xnor U4292 (N_4292,In_1231,N_1060);
nor U4293 (N_4293,N_3567,N_4240);
and U4294 (N_4294,N_3929,N_4227);
or U4295 (N_4295,N_4223,N_4112);
nand U4296 (N_4296,N_4243,N_4083);
or U4297 (N_4297,In_4393,N_4239);
or U4298 (N_4298,N_2427,In_1072);
nor U4299 (N_4299,N_4231,N_3770);
or U4300 (N_4300,In_1265,N_640);
and U4301 (N_4301,N_4073,N_3744);
or U4302 (N_4302,N_4021,N_4099);
xor U4303 (N_4303,N_3005,N_4157);
xnor U4304 (N_4304,N_4208,N_4110);
or U4305 (N_4305,N_4122,N_2842);
and U4306 (N_4306,In_4265,N_4190);
nand U4307 (N_4307,N_2568,N_3750);
nand U4308 (N_4308,N_3669,In_331);
nor U4309 (N_4309,N_4035,N_4145);
or U4310 (N_4310,N_4186,N_3556);
nor U4311 (N_4311,N_3607,N_4017);
and U4312 (N_4312,N_3490,N_3970);
xnor U4313 (N_4313,N_4052,N_3431);
nand U4314 (N_4314,N_3240,N_3719);
xor U4315 (N_4315,N_4130,N_3645);
xnor U4316 (N_4316,N_4019,N_983);
and U4317 (N_4317,N_4241,N_3458);
nor U4318 (N_4318,N_4207,N_3915);
xor U4319 (N_4319,N_4137,N_3859);
and U4320 (N_4320,N_3445,N_3218);
or U4321 (N_4321,N_3938,N_2530);
nand U4322 (N_4322,N_1970,N_4086);
xor U4323 (N_4323,N_1877,N_4054);
nor U4324 (N_4324,N_3373,In_1911);
nand U4325 (N_4325,N_4209,N_2294);
nor U4326 (N_4326,N_4092,N_4031);
or U4327 (N_4327,N_3652,N_45);
nand U4328 (N_4328,N_4180,N_3984);
nor U4329 (N_4329,N_4134,In_1773);
xor U4330 (N_4330,N_4129,N_2162);
nand U4331 (N_4331,N_4213,N_3525);
and U4332 (N_4332,N_2774,N_3443);
nor U4333 (N_4333,N_4159,In_4784);
nand U4334 (N_4334,In_3616,N_3531);
nor U4335 (N_4335,N_4045,N_1901);
xnor U4336 (N_4336,In_2865,N_4059);
nor U4337 (N_4337,N_3185,N_3560);
or U4338 (N_4338,N_2184,N_4136);
and U4339 (N_4339,N_3093,N_4238);
and U4340 (N_4340,N_3883,N_3930);
nor U4341 (N_4341,N_3640,N_4146);
or U4342 (N_4342,N_4120,N_1465);
xor U4343 (N_4343,N_4210,N_3487);
nand U4344 (N_4344,N_3920,N_3002);
xnor U4345 (N_4345,N_3030,N_3074);
and U4346 (N_4346,N_1313,N_4188);
xnor U4347 (N_4347,N_3844,In_775);
nand U4348 (N_4348,N_3805,N_1729);
or U4349 (N_4349,N_3869,N_1023);
and U4350 (N_4350,N_2873,N_4094);
nor U4351 (N_4351,In_2395,In_773);
xnor U4352 (N_4352,N_4026,N_4176);
nand U4353 (N_4353,N_4058,N_3769);
nand U4354 (N_4354,N_3799,N_3830);
and U4355 (N_4355,N_4230,N_4229);
xnor U4356 (N_4356,N_2996,In_2419);
and U4357 (N_4357,N_3289,N_4063);
and U4358 (N_4358,N_3649,N_4012);
nor U4359 (N_4359,N_3433,N_4084);
and U4360 (N_4360,N_3855,N_4202);
or U4361 (N_4361,N_2677,N_3773);
and U4362 (N_4362,N_2241,N_2357);
and U4363 (N_4363,N_3587,N_3812);
nor U4364 (N_4364,N_3819,N_4141);
nand U4365 (N_4365,N_3879,N_3942);
nand U4366 (N_4366,N_2516,N_4156);
nand U4367 (N_4367,N_3379,N_3576);
and U4368 (N_4368,N_4091,N_3892);
nand U4369 (N_4369,N_3366,N_3665);
xor U4370 (N_4370,N_2512,N_4040);
or U4371 (N_4371,N_3853,N_1883);
nor U4372 (N_4372,N_4062,N_3992);
nor U4373 (N_4373,N_2037,In_813);
or U4374 (N_4374,N_4047,N_3673);
nand U4375 (N_4375,N_3579,N_3571);
or U4376 (N_4376,N_3949,N_4232);
or U4377 (N_4377,N_4107,N_3991);
nand U4378 (N_4378,N_4125,N_4219);
and U4379 (N_4379,N_2508,N_3854);
xor U4380 (N_4380,N_3536,N_4193);
or U4381 (N_4381,N_2412,In_2472);
nand U4382 (N_4382,N_955,N_4164);
nand U4383 (N_4383,N_3939,N_4191);
xnor U4384 (N_4384,N_4165,In_2043);
nor U4385 (N_4385,In_3270,N_2847);
xor U4386 (N_4386,N_4143,N_3741);
xnor U4387 (N_4387,In_4733,N_3810);
nor U4388 (N_4388,N_3990,N_3581);
nand U4389 (N_4389,N_3264,N_3781);
or U4390 (N_4390,N_3047,N_3754);
or U4391 (N_4391,N_2861,N_2380);
xor U4392 (N_4392,N_2137,N_3577);
nand U4393 (N_4393,N_4199,N_4088);
or U4394 (N_4394,In_907,N_4169);
nand U4395 (N_4395,N_4142,N_4095);
xor U4396 (N_4396,N_3230,In_3478);
xor U4397 (N_4397,N_3981,N_3957);
or U4398 (N_4398,N_3265,N_4016);
xor U4399 (N_4399,N_3908,In_590);
or U4400 (N_4400,N_1314,N_4150);
nor U4401 (N_4401,N_4153,N_3838);
and U4402 (N_4402,N_3786,N_3697);
nand U4403 (N_4403,N_3657,N_2550);
xor U4404 (N_4404,N_2044,N_4102);
xnor U4405 (N_4405,N_1333,N_3661);
and U4406 (N_4406,N_3313,In_1155);
nand U4407 (N_4407,N_2175,N_1988);
or U4408 (N_4408,N_3239,N_984);
nor U4409 (N_4409,N_4057,N_2730);
xor U4410 (N_4410,N_4071,N_2311);
or U4411 (N_4411,In_1979,N_4126);
or U4412 (N_4412,N_3950,N_4113);
xnor U4413 (N_4413,N_4233,N_3880);
and U4414 (N_4414,N_2751,N_1481);
or U4415 (N_4415,N_3748,N_3197);
xor U4416 (N_4416,N_3680,N_4160);
nand U4417 (N_4417,N_3743,N_2821);
xnor U4418 (N_4418,N_3476,N_4100);
nand U4419 (N_4419,N_3795,N_1512);
or U4420 (N_4420,N_3374,N_4149);
xnor U4421 (N_4421,N_1917,N_532);
xnor U4422 (N_4422,N_552,N_3695);
nor U4423 (N_4423,N_3693,N_4224);
nor U4424 (N_4424,N_4148,N_3802);
and U4425 (N_4425,N_2971,N_3679);
or U4426 (N_4426,N_2417,In_1775);
and U4427 (N_4427,N_3945,N_2613);
xor U4428 (N_4428,N_3572,N_3332);
or U4429 (N_4429,N_4039,In_4426);
nor U4430 (N_4430,N_4079,N_4068);
nand U4431 (N_4431,N_2267,N_4218);
xnor U4432 (N_4432,N_3154,N_3375);
or U4433 (N_4433,N_3122,N_3308);
or U4434 (N_4434,N_2287,N_3186);
nor U4435 (N_4435,N_4173,N_4155);
and U4436 (N_4436,N_3703,N_3818);
nor U4437 (N_4437,N_3080,N_4087);
nand U4438 (N_4438,N_4064,N_2928);
xnor U4439 (N_4439,N_3808,N_3940);
or U4440 (N_4440,N_2715,N_3612);
nor U4441 (N_4441,N_3698,N_3383);
nor U4442 (N_4442,In_4035,N_2561);
nor U4443 (N_4443,N_3670,N_2341);
xor U4444 (N_4444,N_3568,N_3508);
nor U4445 (N_4445,N_4010,N_3580);
nor U4446 (N_4446,N_4036,N_3565);
nand U4447 (N_4447,N_3171,N_3518);
or U4448 (N_4448,N_1107,N_3676);
nor U4449 (N_4449,N_3979,N_4121);
xor U4450 (N_4450,In_4567,N_4203);
nor U4451 (N_4451,N_2830,N_4204);
or U4452 (N_4452,N_2227,N_3198);
nor U4453 (N_4453,N_4075,N_4123);
nor U4454 (N_4454,N_3959,N_4022);
nand U4455 (N_4455,In_2681,N_3811);
nand U4456 (N_4456,N_3798,N_4237);
or U4457 (N_4457,N_4029,N_3097);
nor U4458 (N_4458,N_3684,N_3184);
and U4459 (N_4459,N_4246,In_2795);
and U4460 (N_4460,N_1100,N_4000);
or U4461 (N_4461,N_4116,N_3998);
nor U4462 (N_4462,N_4115,N_3095);
nor U4463 (N_4463,N_4096,N_2787);
nand U4464 (N_4464,N_3763,N_3462);
or U4465 (N_4465,N_4065,N_3321);
xnor U4466 (N_4466,N_2092,N_4056);
or U4467 (N_4467,N_3742,N_3019);
and U4468 (N_4468,N_4131,N_4080);
and U4469 (N_4469,N_4015,In_3900);
nor U4470 (N_4470,N_3923,N_3933);
xnor U4471 (N_4471,N_4104,N_2282);
nand U4472 (N_4472,N_3845,N_3832);
nand U4473 (N_4473,N_4011,N_1619);
nor U4474 (N_4474,N_3346,N_3768);
xor U4475 (N_4475,N_2880,N_4119);
nand U4476 (N_4476,N_4132,N_3020);
nand U4477 (N_4477,N_3671,N_4163);
or U4478 (N_4478,N_3971,In_4227);
or U4479 (N_4479,In_1915,N_4069);
or U4480 (N_4480,N_4002,N_3234);
nand U4481 (N_4481,N_2723,N_3460);
nand U4482 (N_4482,N_4222,N_4151);
nand U4483 (N_4483,N_4097,In_124);
or U4484 (N_4484,In_562,N_2713);
nor U4485 (N_4485,N_3787,N_4034);
and U4486 (N_4486,N_3479,N_4144);
and U4487 (N_4487,N_4171,N_3711);
and U4488 (N_4488,N_3960,N_2790);
or U4489 (N_4489,In_2020,In_3943);
and U4490 (N_4490,N_3354,N_4127);
nor U4491 (N_4491,N_4211,N_4124);
nor U4492 (N_4492,N_3547,N_4236);
nor U4493 (N_4493,N_2545,N_4037);
and U4494 (N_4494,N_343,N_3925);
xnor U4495 (N_4495,In_3885,N_4006);
xor U4496 (N_4496,N_3922,N_4200);
xnor U4497 (N_4497,N_4152,N_4175);
or U4498 (N_4498,N_4215,N_3860);
nor U4499 (N_4499,N_3638,N_3619);
nor U4500 (N_4500,N_4296,N_3521);
nand U4501 (N_4501,N_2245,N_4381);
xnor U4502 (N_4502,N_4497,N_3633);
nor U4503 (N_4503,N_3967,N_4085);
nor U4504 (N_4504,N_4268,N_4007);
xnor U4505 (N_4505,N_4162,N_4418);
and U4506 (N_4506,N_4436,N_4491);
nand U4507 (N_4507,N_4074,N_4263);
xor U4508 (N_4508,N_4346,N_4341);
and U4509 (N_4509,N_2932,N_4284);
and U4510 (N_4510,N_4340,N_4350);
or U4511 (N_4511,N_2573,N_4439);
xnor U4512 (N_4512,N_3274,N_3894);
and U4513 (N_4513,N_4394,N_2143);
nand U4514 (N_4514,N_4365,N_4421);
or U4515 (N_4515,N_4442,N_4435);
nor U4516 (N_4516,N_4479,N_860);
and U4517 (N_4517,N_4024,N_4333);
nor U4518 (N_4518,N_1260,N_304);
and U4519 (N_4519,N_3015,N_4271);
or U4520 (N_4520,N_4348,N_3813);
and U4521 (N_4521,N_4277,N_4406);
nand U4522 (N_4522,N_3729,N_4323);
xor U4523 (N_4523,N_3747,N_3906);
xnor U4524 (N_4524,N_4462,N_4488);
or U4525 (N_4525,N_4269,N_3611);
xor U4526 (N_4526,N_4461,N_4293);
and U4527 (N_4527,N_4279,N_4308);
nand U4528 (N_4528,N_3932,N_3888);
and U4529 (N_4529,N_4449,N_3909);
nand U4530 (N_4530,N_4128,N_4369);
and U4531 (N_4531,N_4228,N_4041);
nor U4532 (N_4532,N_4255,N_4286);
nor U4533 (N_4533,N_4481,N_3622);
and U4534 (N_4534,N_4189,N_2196);
and U4535 (N_4535,N_3170,N_4212);
nor U4536 (N_4536,N_1597,In_1111);
or U4537 (N_4537,N_4414,N_2509);
xnor U4538 (N_4538,N_4306,N_4198);
nor U4539 (N_4539,N_4468,N_4448);
xor U4540 (N_4540,N_4138,N_4055);
or U4541 (N_4541,N_4247,N_4032);
xnor U4542 (N_4542,N_4476,N_1899);
xnor U4543 (N_4543,N_4261,N_4225);
or U4544 (N_4544,N_4242,N_4334);
nand U4545 (N_4545,N_4318,N_4419);
xnor U4546 (N_4546,N_4376,N_3863);
nand U4547 (N_4547,N_2523,N_2597);
nand U4548 (N_4548,N_4259,N_4423);
nor U4549 (N_4549,N_4492,N_4264);
nor U4550 (N_4550,N_3512,N_4226);
and U4551 (N_4551,N_3760,N_4388);
and U4552 (N_4552,N_4289,N_3129);
or U4553 (N_4553,N_4273,N_4413);
or U4554 (N_4554,N_4408,In_3379);
or U4555 (N_4555,N_3293,N_4415);
and U4556 (N_4556,N_3478,In_3584);
and U4557 (N_4557,N_4427,N_4103);
nand U4558 (N_4558,N_4290,N_4432);
or U4559 (N_4559,N_4313,N_3013);
nor U4560 (N_4560,N_4266,N_4285);
nor U4561 (N_4561,N_4446,N_3842);
and U4562 (N_4562,N_4440,N_4252);
and U4563 (N_4563,N_4257,N_2258);
and U4564 (N_4564,In_1459,N_4329);
nor U4565 (N_4565,In_1721,N_4402);
or U4566 (N_4566,N_4383,N_4336);
or U4567 (N_4567,N_3756,N_4477);
xnor U4568 (N_4568,N_3504,N_4499);
nand U4569 (N_4569,N_3969,N_4003);
or U4570 (N_4570,N_3157,N_4475);
nand U4571 (N_4571,N_4473,N_4298);
or U4572 (N_4572,N_4373,N_4322);
nor U4573 (N_4573,N_4486,N_4372);
and U4574 (N_4574,N_4028,N_4244);
or U4575 (N_4575,N_4400,N_3222);
or U4576 (N_4576,N_3952,N_4352);
or U4577 (N_4577,N_2498,N_3172);
nor U4578 (N_4578,N_4314,N_4326);
and U4579 (N_4579,N_3647,N_4471);
and U4580 (N_4580,N_4201,N_4248);
xnor U4581 (N_4581,N_4454,N_4288);
xnor U4582 (N_4582,N_4281,N_4455);
and U4583 (N_4583,N_3335,In_2112);
nand U4584 (N_4584,N_3331,N_4349);
or U4585 (N_4585,N_4392,N_4008);
and U4586 (N_4586,N_4437,N_3260);
and U4587 (N_4587,N_4386,N_3468);
and U4588 (N_4588,N_4379,N_986);
nor U4589 (N_4589,N_4262,N_3041);
and U4590 (N_4590,N_4297,N_3439);
or U4591 (N_4591,In_642,N_4370);
nand U4592 (N_4592,N_3298,N_4451);
nor U4593 (N_4593,N_4044,N_4354);
or U4594 (N_4594,N_4001,N_4342);
and U4595 (N_4595,N_4182,N_3797);
or U4596 (N_4596,N_4391,N_3972);
nand U4597 (N_4597,N_4101,N_4411);
nor U4598 (N_4598,N_4390,N_2020);
or U4599 (N_4599,N_4339,N_4483);
or U4600 (N_4600,N_4158,N_3656);
nor U4601 (N_4601,N_3881,N_4109);
xnor U4602 (N_4602,N_2800,N_4382);
nand U4603 (N_4603,N_2964,N_4428);
xnor U4604 (N_4604,N_4278,N_4367);
or U4605 (N_4605,N_1283,N_4407);
or U4606 (N_4606,In_3208,N_3815);
or U4607 (N_4607,N_4396,In_1270);
xor U4608 (N_4608,N_3997,N_4467);
or U4609 (N_4609,N_4114,N_2874);
xor U4610 (N_4610,N_3706,N_4434);
xnor U4611 (N_4611,N_3896,N_3890);
nor U4612 (N_4612,N_119,N_4315);
nand U4613 (N_4613,N_4393,N_2157);
and U4614 (N_4614,N_4307,N_4174);
and U4615 (N_4615,N_4345,N_4378);
xor U4616 (N_4616,N_465,N_4321);
or U4617 (N_4617,N_4178,N_1836);
nand U4618 (N_4618,N_4270,N_4325);
and U4619 (N_4619,N_4401,N_3437);
nor U4620 (N_4620,N_3803,N_4357);
and U4621 (N_4621,N_4305,N_4154);
xor U4622 (N_4622,N_3474,N_3966);
and U4623 (N_4623,N_3804,N_3410);
or U4624 (N_4624,In_2722,N_4292);
and U4625 (N_4625,N_3251,N_4291);
or U4626 (N_4626,N_4356,N_3319);
and U4627 (N_4627,N_4495,N_2270);
nor U4628 (N_4628,N_2927,N_4250);
or U4629 (N_4629,N_4140,N_1385);
nand U4630 (N_4630,N_3870,N_2255);
xor U4631 (N_4631,N_4430,N_2999);
and U4632 (N_4632,N_3200,N_4403);
or U4633 (N_4633,N_4441,In_3722);
or U4634 (N_4634,N_4445,N_4267);
and U4635 (N_4635,N_4361,In_3762);
or U4636 (N_4636,N_4181,N_1120);
xnor U4637 (N_4637,N_4009,N_4425);
and U4638 (N_4638,N_4332,N_4276);
nor U4639 (N_4639,N_4496,N_4433);
xor U4640 (N_4640,N_4494,N_3297);
nand U4641 (N_4641,In_4575,N_4482);
or U4642 (N_4642,N_4108,N_2951);
xor U4643 (N_4643,N_4384,N_4217);
nor U4644 (N_4644,N_4076,N_3659);
nor U4645 (N_4645,N_3598,N_4251);
or U4646 (N_4646,N_4380,N_3723);
xnor U4647 (N_4647,N_4387,In_3090);
xnor U4648 (N_4648,N_4106,N_1637);
xor U4649 (N_4649,N_4474,N_4300);
nand U4650 (N_4650,N_4135,N_4030);
nor U4651 (N_4651,N_3897,N_3724);
or U4652 (N_4652,N_4463,N_1551);
or U4653 (N_4653,N_4282,N_4042);
nand U4654 (N_4654,N_4265,N_3833);
or U4655 (N_4655,N_4429,N_4295);
xor U4656 (N_4656,N_2011,N_3943);
xor U4657 (N_4657,N_4490,N_4424);
xor U4658 (N_4658,N_4275,N_4320);
xor U4659 (N_4659,N_4487,N_4412);
and U4660 (N_4660,In_2409,N_4420);
nor U4661 (N_4661,N_3868,N_4489);
and U4662 (N_4662,N_4197,N_4235);
and U4663 (N_4663,In_3453,N_3739);
nor U4664 (N_4664,N_4457,N_3827);
nor U4665 (N_4665,N_3782,N_4067);
nand U4666 (N_4666,N_50,N_4389);
nor U4667 (N_4667,N_3974,N_4194);
and U4668 (N_4668,N_3977,N_3851);
nand U4669 (N_4669,N_2859,N_4077);
nand U4670 (N_4670,N_4472,N_4453);
nand U4671 (N_4671,N_4310,N_4371);
and U4672 (N_4672,N_4478,N_4480);
xnor U4673 (N_4673,N_4355,N_4395);
nor U4674 (N_4674,N_4366,N_4324);
or U4675 (N_4675,N_4466,N_4431);
nand U4676 (N_4676,N_4364,N_4312);
or U4677 (N_4677,N_4469,N_3663);
nand U4678 (N_4678,N_2737,N_4464);
nor U4679 (N_4679,N_4330,N_4206);
nand U4680 (N_4680,N_3841,N_4256);
and U4681 (N_4681,N_2924,N_4023);
nor U4682 (N_4682,N_4303,N_4493);
xnor U4683 (N_4683,N_4410,N_4452);
nand U4684 (N_4684,N_4111,N_4343);
nor U4685 (N_4685,N_4294,N_4299);
xor U4686 (N_4686,N_2633,N_4374);
or U4687 (N_4687,N_4098,N_4443);
nor U4688 (N_4688,N_4027,N_4331);
xnor U4689 (N_4689,N_3707,N_4117);
nand U4690 (N_4690,N_4220,N_4072);
and U4691 (N_4691,N_2896,N_4283);
or U4692 (N_4692,N_4484,N_4301);
nor U4693 (N_4693,N_4196,N_4358);
xor U4694 (N_4694,N_4498,N_4405);
and U4695 (N_4695,N_4205,N_3961);
and U4696 (N_4696,N_4485,N_4184);
nor U4697 (N_4697,N_1158,N_4093);
or U4698 (N_4698,N_2645,N_3039);
xor U4699 (N_4699,N_4338,N_4327);
nor U4700 (N_4700,N_2571,N_4458);
xor U4701 (N_4701,N_4368,N_4311);
nor U4702 (N_4702,N_4335,N_3865);
and U4703 (N_4703,N_4385,N_4258);
and U4704 (N_4704,N_4280,N_4444);
nand U4705 (N_4705,N_4053,N_4399);
xor U4706 (N_4706,N_3779,N_4187);
and U4707 (N_4707,N_4081,N_948);
nor U4708 (N_4708,N_4018,N_4172);
or U4709 (N_4709,N_3843,N_3481);
and U4710 (N_4710,N_1748,N_4118);
nor U4711 (N_4711,N_4351,N_4046);
or U4712 (N_4712,N_4020,N_4214);
or U4713 (N_4713,N_4316,N_4447);
xnor U4714 (N_4714,N_4319,N_4470);
and U4715 (N_4715,N_4353,N_4409);
nand U4716 (N_4716,N_4426,N_4061);
and U4717 (N_4717,N_4460,N_4362);
or U4718 (N_4718,In_2866,N_1540);
or U4719 (N_4719,N_4317,N_4274);
xnor U4720 (N_4720,N_4249,N_3348);
xnor U4721 (N_4721,N_3505,N_4422);
and U4722 (N_4722,N_4404,N_4359);
and U4723 (N_4723,N_4416,N_3924);
nand U4724 (N_4724,In_1559,N_4260);
or U4725 (N_4725,N_4456,N_4253);
nand U4726 (N_4726,N_4363,N_2310);
or U4727 (N_4727,N_4360,N_4060);
or U4728 (N_4728,N_4465,N_4004);
nor U4729 (N_4729,N_4397,N_4082);
xor U4730 (N_4730,N_3856,N_3834);
xor U4731 (N_4731,N_2805,In_4382);
nand U4732 (N_4732,N_4089,N_4183);
xor U4733 (N_4733,N_3597,N_4398);
nand U4734 (N_4734,N_4344,N_2434);
and U4735 (N_4735,N_4302,N_4438);
and U4736 (N_4736,N_4304,N_4377);
xnor U4737 (N_4737,N_3116,N_4417);
and U4738 (N_4738,In_3799,N_4216);
nor U4739 (N_4739,N_3752,N_4105);
and U4740 (N_4740,N_4287,N_3432);
or U4741 (N_4741,In_1077,N_3353);
xnor U4742 (N_4742,N_4450,N_1365);
nor U4743 (N_4743,N_4375,N_3430);
nor U4744 (N_4744,N_4309,N_2970);
nand U4745 (N_4745,N_4347,N_4459);
and U4746 (N_4746,N_4272,N_4038);
nand U4747 (N_4747,N_4254,In_516);
xor U4748 (N_4748,N_4328,In_682);
nand U4749 (N_4749,N_3574,N_4337);
xor U4750 (N_4750,N_4644,N_4589);
nor U4751 (N_4751,N_4696,N_4564);
nand U4752 (N_4752,N_4583,N_4604);
and U4753 (N_4753,N_4731,N_4542);
or U4754 (N_4754,N_4570,N_4651);
and U4755 (N_4755,N_4592,N_4551);
xnor U4756 (N_4756,N_4671,N_4668);
xnor U4757 (N_4757,N_4584,N_4580);
or U4758 (N_4758,N_4700,N_4693);
or U4759 (N_4759,N_4521,N_4523);
or U4760 (N_4760,N_4555,N_4682);
and U4761 (N_4761,N_4742,N_4710);
xor U4762 (N_4762,N_4686,N_4591);
nor U4763 (N_4763,N_4738,N_4608);
or U4764 (N_4764,N_4505,N_4728);
nand U4765 (N_4765,N_4552,N_4640);
or U4766 (N_4766,N_4639,N_4629);
nand U4767 (N_4767,N_4743,N_4709);
nand U4768 (N_4768,N_4548,N_4574);
and U4769 (N_4769,N_4507,N_4582);
nand U4770 (N_4770,N_4503,N_4605);
and U4771 (N_4771,N_4661,N_4735);
xor U4772 (N_4772,N_4539,N_4610);
xor U4773 (N_4773,N_4697,N_4732);
nor U4774 (N_4774,N_4606,N_4681);
and U4775 (N_4775,N_4745,N_4520);
xor U4776 (N_4776,N_4729,N_4624);
nand U4777 (N_4777,N_4657,N_4588);
nand U4778 (N_4778,N_4741,N_4641);
and U4779 (N_4779,N_4667,N_4734);
nand U4780 (N_4780,N_4566,N_4692);
nand U4781 (N_4781,N_4663,N_4561);
nand U4782 (N_4782,N_4655,N_4642);
or U4783 (N_4783,N_4670,N_4634);
and U4784 (N_4784,N_4510,N_4748);
nand U4785 (N_4785,N_4649,N_4553);
or U4786 (N_4786,N_4637,N_4685);
xnor U4787 (N_4787,N_4724,N_4719);
nand U4788 (N_4788,N_4660,N_4509);
nand U4789 (N_4789,N_4699,N_4549);
nor U4790 (N_4790,N_4704,N_4576);
or U4791 (N_4791,N_4543,N_4617);
nor U4792 (N_4792,N_4623,N_4601);
xnor U4793 (N_4793,N_4609,N_4594);
or U4794 (N_4794,N_4712,N_4658);
and U4795 (N_4795,N_4744,N_4645);
or U4796 (N_4796,N_4602,N_4577);
or U4797 (N_4797,N_4679,N_4746);
nand U4798 (N_4798,N_4636,N_4695);
and U4799 (N_4799,N_4526,N_4654);
or U4800 (N_4800,N_4500,N_4721);
xnor U4801 (N_4801,N_4530,N_4627);
or U4802 (N_4802,N_4519,N_4727);
nor U4803 (N_4803,N_4718,N_4586);
nand U4804 (N_4804,N_4508,N_4717);
nand U4805 (N_4805,N_4702,N_4567);
or U4806 (N_4806,N_4534,N_4689);
nor U4807 (N_4807,N_4665,N_4632);
and U4808 (N_4808,N_4714,N_4533);
xnor U4809 (N_4809,N_4678,N_4653);
xnor U4810 (N_4810,N_4677,N_4573);
nor U4811 (N_4811,N_4711,N_4687);
and U4812 (N_4812,N_4706,N_4547);
nand U4813 (N_4813,N_4554,N_4688);
or U4814 (N_4814,N_4513,N_4648);
nor U4815 (N_4815,N_4698,N_4733);
nand U4816 (N_4816,N_4633,N_4585);
or U4817 (N_4817,N_4662,N_4647);
and U4818 (N_4818,N_4638,N_4611);
xnor U4819 (N_4819,N_4643,N_4664);
nor U4820 (N_4820,N_4707,N_4532);
nor U4821 (N_4821,N_4650,N_4720);
nor U4822 (N_4822,N_4544,N_4504);
or U4823 (N_4823,N_4502,N_4587);
xor U4824 (N_4824,N_4622,N_4691);
or U4825 (N_4825,N_4626,N_4625);
nor U4826 (N_4826,N_4619,N_4597);
nand U4827 (N_4827,N_4512,N_4527);
xor U4828 (N_4828,N_4716,N_4723);
nand U4829 (N_4829,N_4524,N_4736);
or U4830 (N_4830,N_4579,N_4615);
or U4831 (N_4831,N_4581,N_4518);
nor U4832 (N_4832,N_4614,N_4631);
and U4833 (N_4833,N_4703,N_4747);
or U4834 (N_4834,N_4646,N_4529);
nor U4835 (N_4835,N_4531,N_4511);
nand U4836 (N_4836,N_4621,N_4517);
and U4837 (N_4837,N_4514,N_4708);
or U4838 (N_4838,N_4669,N_4536);
nor U4839 (N_4839,N_4550,N_4538);
or U4840 (N_4840,N_4676,N_4565);
and U4841 (N_4841,N_4557,N_4558);
or U4842 (N_4842,N_4572,N_4730);
nand U4843 (N_4843,N_4659,N_4590);
xor U4844 (N_4844,N_4569,N_4607);
and U4845 (N_4845,N_4684,N_4635);
nand U4846 (N_4846,N_4596,N_4603);
nor U4847 (N_4847,N_4683,N_4578);
and U4848 (N_4848,N_4749,N_4535);
nor U4849 (N_4849,N_4722,N_4705);
nand U4850 (N_4850,N_4726,N_4715);
and U4851 (N_4851,N_4620,N_4739);
nor U4852 (N_4852,N_4690,N_4501);
and U4853 (N_4853,N_4598,N_4674);
or U4854 (N_4854,N_4652,N_4701);
nor U4855 (N_4855,N_4575,N_4568);
nor U4856 (N_4856,N_4562,N_4628);
or U4857 (N_4857,N_4559,N_4656);
xnor U4858 (N_4858,N_4593,N_4616);
nand U4859 (N_4859,N_4680,N_4541);
or U4860 (N_4860,N_4666,N_4694);
xor U4861 (N_4861,N_4713,N_4630);
and U4862 (N_4862,N_4599,N_4506);
and U4863 (N_4863,N_4545,N_4537);
or U4864 (N_4864,N_4595,N_4618);
nand U4865 (N_4865,N_4556,N_4540);
nand U4866 (N_4866,N_4673,N_4522);
nor U4867 (N_4867,N_4600,N_4675);
nor U4868 (N_4868,N_4546,N_4571);
and U4869 (N_4869,N_4525,N_4725);
nand U4870 (N_4870,N_4528,N_4563);
and U4871 (N_4871,N_4515,N_4560);
nor U4872 (N_4872,N_4516,N_4672);
xor U4873 (N_4873,N_4740,N_4612);
nor U4874 (N_4874,N_4737,N_4613);
and U4875 (N_4875,N_4705,N_4536);
nand U4876 (N_4876,N_4520,N_4715);
nor U4877 (N_4877,N_4691,N_4648);
xnor U4878 (N_4878,N_4638,N_4532);
xnor U4879 (N_4879,N_4504,N_4660);
nand U4880 (N_4880,N_4571,N_4690);
xnor U4881 (N_4881,N_4530,N_4698);
or U4882 (N_4882,N_4685,N_4698);
or U4883 (N_4883,N_4573,N_4712);
nand U4884 (N_4884,N_4733,N_4552);
and U4885 (N_4885,N_4697,N_4552);
xor U4886 (N_4886,N_4610,N_4646);
nand U4887 (N_4887,N_4621,N_4569);
nor U4888 (N_4888,N_4642,N_4741);
and U4889 (N_4889,N_4670,N_4702);
and U4890 (N_4890,N_4570,N_4610);
or U4891 (N_4891,N_4549,N_4577);
or U4892 (N_4892,N_4725,N_4500);
nand U4893 (N_4893,N_4611,N_4506);
and U4894 (N_4894,N_4554,N_4634);
and U4895 (N_4895,N_4645,N_4650);
nand U4896 (N_4896,N_4726,N_4686);
xnor U4897 (N_4897,N_4512,N_4603);
nor U4898 (N_4898,N_4669,N_4578);
and U4899 (N_4899,N_4684,N_4570);
nand U4900 (N_4900,N_4666,N_4618);
nor U4901 (N_4901,N_4673,N_4724);
xor U4902 (N_4902,N_4518,N_4633);
xnor U4903 (N_4903,N_4694,N_4637);
or U4904 (N_4904,N_4588,N_4717);
xnor U4905 (N_4905,N_4654,N_4594);
nand U4906 (N_4906,N_4723,N_4680);
nand U4907 (N_4907,N_4637,N_4636);
or U4908 (N_4908,N_4590,N_4503);
nor U4909 (N_4909,N_4679,N_4542);
or U4910 (N_4910,N_4704,N_4559);
nor U4911 (N_4911,N_4643,N_4719);
xor U4912 (N_4912,N_4641,N_4595);
and U4913 (N_4913,N_4617,N_4713);
nand U4914 (N_4914,N_4615,N_4635);
nor U4915 (N_4915,N_4674,N_4518);
and U4916 (N_4916,N_4550,N_4681);
xnor U4917 (N_4917,N_4544,N_4672);
nand U4918 (N_4918,N_4725,N_4537);
nor U4919 (N_4919,N_4690,N_4660);
and U4920 (N_4920,N_4513,N_4548);
xor U4921 (N_4921,N_4670,N_4635);
nand U4922 (N_4922,N_4644,N_4687);
nor U4923 (N_4923,N_4743,N_4673);
xor U4924 (N_4924,N_4560,N_4711);
nor U4925 (N_4925,N_4706,N_4670);
nor U4926 (N_4926,N_4515,N_4613);
or U4927 (N_4927,N_4571,N_4548);
or U4928 (N_4928,N_4524,N_4531);
or U4929 (N_4929,N_4603,N_4641);
nand U4930 (N_4930,N_4606,N_4503);
nand U4931 (N_4931,N_4544,N_4520);
and U4932 (N_4932,N_4521,N_4658);
or U4933 (N_4933,N_4688,N_4626);
nand U4934 (N_4934,N_4556,N_4696);
xor U4935 (N_4935,N_4711,N_4541);
nand U4936 (N_4936,N_4688,N_4598);
or U4937 (N_4937,N_4601,N_4652);
or U4938 (N_4938,N_4588,N_4667);
and U4939 (N_4939,N_4619,N_4605);
and U4940 (N_4940,N_4645,N_4656);
and U4941 (N_4941,N_4549,N_4568);
and U4942 (N_4942,N_4544,N_4587);
or U4943 (N_4943,N_4718,N_4623);
xor U4944 (N_4944,N_4610,N_4593);
nand U4945 (N_4945,N_4738,N_4566);
nand U4946 (N_4946,N_4733,N_4688);
or U4947 (N_4947,N_4639,N_4549);
nor U4948 (N_4948,N_4565,N_4609);
and U4949 (N_4949,N_4577,N_4698);
or U4950 (N_4950,N_4520,N_4610);
nand U4951 (N_4951,N_4664,N_4636);
and U4952 (N_4952,N_4566,N_4706);
nand U4953 (N_4953,N_4547,N_4712);
xnor U4954 (N_4954,N_4654,N_4529);
or U4955 (N_4955,N_4691,N_4747);
or U4956 (N_4956,N_4685,N_4622);
xnor U4957 (N_4957,N_4726,N_4645);
xnor U4958 (N_4958,N_4604,N_4597);
and U4959 (N_4959,N_4539,N_4682);
nand U4960 (N_4960,N_4538,N_4702);
nand U4961 (N_4961,N_4651,N_4537);
nor U4962 (N_4962,N_4687,N_4731);
and U4963 (N_4963,N_4627,N_4670);
and U4964 (N_4964,N_4700,N_4545);
xor U4965 (N_4965,N_4649,N_4604);
nand U4966 (N_4966,N_4548,N_4527);
and U4967 (N_4967,N_4674,N_4675);
xnor U4968 (N_4968,N_4663,N_4630);
nand U4969 (N_4969,N_4593,N_4687);
or U4970 (N_4970,N_4745,N_4631);
nand U4971 (N_4971,N_4698,N_4641);
xnor U4972 (N_4972,N_4636,N_4503);
xor U4973 (N_4973,N_4520,N_4542);
and U4974 (N_4974,N_4581,N_4631);
xnor U4975 (N_4975,N_4730,N_4567);
or U4976 (N_4976,N_4657,N_4656);
nand U4977 (N_4977,N_4582,N_4702);
nor U4978 (N_4978,N_4631,N_4543);
or U4979 (N_4979,N_4689,N_4522);
xor U4980 (N_4980,N_4580,N_4653);
or U4981 (N_4981,N_4503,N_4577);
nor U4982 (N_4982,N_4702,N_4513);
nor U4983 (N_4983,N_4571,N_4580);
and U4984 (N_4984,N_4544,N_4725);
xnor U4985 (N_4985,N_4684,N_4523);
or U4986 (N_4986,N_4649,N_4650);
xnor U4987 (N_4987,N_4694,N_4673);
and U4988 (N_4988,N_4681,N_4608);
nor U4989 (N_4989,N_4668,N_4552);
or U4990 (N_4990,N_4652,N_4602);
nor U4991 (N_4991,N_4576,N_4748);
and U4992 (N_4992,N_4625,N_4739);
nand U4993 (N_4993,N_4709,N_4669);
xnor U4994 (N_4994,N_4665,N_4508);
xor U4995 (N_4995,N_4710,N_4632);
nand U4996 (N_4996,N_4682,N_4505);
xor U4997 (N_4997,N_4622,N_4602);
or U4998 (N_4998,N_4746,N_4539);
and U4999 (N_4999,N_4711,N_4542);
xor U5000 (N_5000,N_4862,N_4866);
nor U5001 (N_5001,N_4774,N_4771);
xnor U5002 (N_5002,N_4910,N_4947);
or U5003 (N_5003,N_4904,N_4926);
xor U5004 (N_5004,N_4785,N_4888);
nor U5005 (N_5005,N_4822,N_4795);
xnor U5006 (N_5006,N_4818,N_4808);
or U5007 (N_5007,N_4952,N_4870);
or U5008 (N_5008,N_4970,N_4913);
xnor U5009 (N_5009,N_4900,N_4813);
or U5010 (N_5010,N_4833,N_4846);
nand U5011 (N_5011,N_4765,N_4816);
nand U5012 (N_5012,N_4809,N_4908);
and U5013 (N_5013,N_4950,N_4769);
xnor U5014 (N_5014,N_4814,N_4890);
nor U5015 (N_5015,N_4750,N_4954);
or U5016 (N_5016,N_4907,N_4906);
or U5017 (N_5017,N_4828,N_4827);
nor U5018 (N_5018,N_4902,N_4789);
nand U5019 (N_5019,N_4930,N_4983);
and U5020 (N_5020,N_4892,N_4791);
and U5021 (N_5021,N_4971,N_4759);
or U5022 (N_5022,N_4770,N_4756);
nor U5023 (N_5023,N_4886,N_4937);
nor U5024 (N_5024,N_4920,N_4855);
and U5025 (N_5025,N_4847,N_4875);
nand U5026 (N_5026,N_4777,N_4802);
nand U5027 (N_5027,N_4979,N_4896);
or U5028 (N_5028,N_4836,N_4831);
or U5029 (N_5029,N_4850,N_4996);
xnor U5030 (N_5030,N_4845,N_4824);
nor U5031 (N_5031,N_4905,N_4819);
xnor U5032 (N_5032,N_4849,N_4931);
nand U5033 (N_5033,N_4976,N_4865);
or U5034 (N_5034,N_4891,N_4767);
nand U5035 (N_5035,N_4974,N_4864);
or U5036 (N_5036,N_4988,N_4805);
xnor U5037 (N_5037,N_4782,N_4923);
xor U5038 (N_5038,N_4914,N_4867);
xnor U5039 (N_5039,N_4945,N_4953);
nor U5040 (N_5040,N_4977,N_4811);
or U5041 (N_5041,N_4925,N_4984);
nor U5042 (N_5042,N_4879,N_4852);
nor U5043 (N_5043,N_4962,N_4779);
or U5044 (N_5044,N_4911,N_4963);
and U5045 (N_5045,N_4972,N_4843);
xor U5046 (N_5046,N_4844,N_4885);
nor U5047 (N_5047,N_4815,N_4820);
and U5048 (N_5048,N_4882,N_4994);
xnor U5049 (N_5049,N_4948,N_4960);
and U5050 (N_5050,N_4793,N_4932);
xnor U5051 (N_5051,N_4853,N_4830);
and U5052 (N_5052,N_4758,N_4941);
xnor U5053 (N_5053,N_4764,N_4924);
nand U5054 (N_5054,N_4939,N_4776);
and U5055 (N_5055,N_4762,N_4861);
or U5056 (N_5056,N_4978,N_4942);
xnor U5057 (N_5057,N_4835,N_4944);
and U5058 (N_5058,N_4753,N_4991);
or U5059 (N_5059,N_4949,N_4946);
and U5060 (N_5060,N_4992,N_4797);
xor U5061 (N_5061,N_4995,N_4881);
nand U5062 (N_5062,N_4751,N_4982);
or U5063 (N_5063,N_4778,N_4783);
and U5064 (N_5064,N_4859,N_4993);
nor U5065 (N_5065,N_4938,N_4887);
nor U5066 (N_5066,N_4915,N_4817);
nor U5067 (N_5067,N_4966,N_4754);
and U5068 (N_5068,N_4755,N_4784);
or U5069 (N_5069,N_4825,N_4958);
or U5070 (N_5070,N_4981,N_4940);
nor U5071 (N_5071,N_4842,N_4772);
and U5072 (N_5072,N_4922,N_4893);
and U5073 (N_5073,N_4957,N_4799);
xor U5074 (N_5074,N_4903,N_4796);
nor U5075 (N_5075,N_4928,N_4921);
and U5076 (N_5076,N_4841,N_4874);
and U5077 (N_5077,N_4969,N_4975);
xnor U5078 (N_5078,N_4840,N_4810);
nor U5079 (N_5079,N_4832,N_4951);
and U5080 (N_5080,N_4858,N_4956);
xnor U5081 (N_5081,N_4829,N_4851);
xnor U5082 (N_5082,N_4880,N_4883);
and U5083 (N_5083,N_4794,N_4826);
nand U5084 (N_5084,N_4894,N_4919);
nand U5085 (N_5085,N_4868,N_4790);
nor U5086 (N_5086,N_4934,N_4760);
xnor U5087 (N_5087,N_4834,N_4857);
or U5088 (N_5088,N_4801,N_4786);
nand U5089 (N_5089,N_4871,N_4973);
or U5090 (N_5090,N_4916,N_4927);
or U5091 (N_5091,N_4763,N_4838);
or U5092 (N_5092,N_4837,N_4967);
nand U5093 (N_5093,N_4901,N_4897);
nand U5094 (N_5094,N_4860,N_4773);
nor U5095 (N_5095,N_4986,N_4757);
xor U5096 (N_5096,N_4935,N_4895);
nand U5097 (N_5097,N_4839,N_4899);
nor U5098 (N_5098,N_4876,N_4990);
xor U5099 (N_5099,N_4807,N_4997);
or U5100 (N_5100,N_4812,N_4987);
and U5101 (N_5101,N_4936,N_4943);
and U5102 (N_5102,N_4792,N_4806);
nand U5103 (N_5103,N_4889,N_4980);
and U5104 (N_5104,N_4863,N_4909);
or U5105 (N_5105,N_4856,N_4854);
and U5106 (N_5106,N_4787,N_4884);
and U5107 (N_5107,N_4804,N_4998);
and U5108 (N_5108,N_4965,N_4929);
xor U5109 (N_5109,N_4873,N_4917);
or U5110 (N_5110,N_4964,N_4912);
xor U5111 (N_5111,N_4821,N_4800);
or U5112 (N_5112,N_4959,N_4985);
or U5113 (N_5113,N_4877,N_4869);
nand U5114 (N_5114,N_4766,N_4999);
nand U5115 (N_5115,N_4878,N_4823);
nor U5116 (N_5116,N_4989,N_4798);
or U5117 (N_5117,N_4780,N_4933);
and U5118 (N_5118,N_4803,N_4768);
and U5119 (N_5119,N_4752,N_4788);
nor U5120 (N_5120,N_4898,N_4781);
nand U5121 (N_5121,N_4968,N_4775);
xor U5122 (N_5122,N_4848,N_4918);
and U5123 (N_5123,N_4961,N_4872);
xor U5124 (N_5124,N_4955,N_4761);
nand U5125 (N_5125,N_4983,N_4948);
xor U5126 (N_5126,N_4825,N_4932);
or U5127 (N_5127,N_4896,N_4790);
nor U5128 (N_5128,N_4977,N_4949);
or U5129 (N_5129,N_4928,N_4936);
xor U5130 (N_5130,N_4823,N_4872);
nand U5131 (N_5131,N_4934,N_4863);
and U5132 (N_5132,N_4881,N_4923);
nor U5133 (N_5133,N_4788,N_4830);
nor U5134 (N_5134,N_4989,N_4992);
or U5135 (N_5135,N_4951,N_4753);
or U5136 (N_5136,N_4785,N_4809);
nor U5137 (N_5137,N_4822,N_4825);
nand U5138 (N_5138,N_4980,N_4971);
and U5139 (N_5139,N_4803,N_4970);
nor U5140 (N_5140,N_4936,N_4975);
xor U5141 (N_5141,N_4986,N_4853);
and U5142 (N_5142,N_4803,N_4860);
nand U5143 (N_5143,N_4935,N_4867);
and U5144 (N_5144,N_4851,N_4844);
nor U5145 (N_5145,N_4824,N_4783);
xnor U5146 (N_5146,N_4988,N_4761);
and U5147 (N_5147,N_4854,N_4875);
or U5148 (N_5148,N_4754,N_4785);
and U5149 (N_5149,N_4925,N_4987);
or U5150 (N_5150,N_4956,N_4840);
nor U5151 (N_5151,N_4769,N_4867);
or U5152 (N_5152,N_4925,N_4883);
or U5153 (N_5153,N_4752,N_4803);
or U5154 (N_5154,N_4943,N_4890);
xnor U5155 (N_5155,N_4895,N_4765);
nand U5156 (N_5156,N_4753,N_4805);
xnor U5157 (N_5157,N_4955,N_4777);
xor U5158 (N_5158,N_4956,N_4760);
nor U5159 (N_5159,N_4920,N_4854);
nand U5160 (N_5160,N_4789,N_4943);
or U5161 (N_5161,N_4907,N_4876);
or U5162 (N_5162,N_4978,N_4947);
and U5163 (N_5163,N_4841,N_4973);
xor U5164 (N_5164,N_4906,N_4966);
xor U5165 (N_5165,N_4817,N_4811);
or U5166 (N_5166,N_4931,N_4858);
or U5167 (N_5167,N_4757,N_4865);
and U5168 (N_5168,N_4837,N_4797);
nand U5169 (N_5169,N_4866,N_4815);
nand U5170 (N_5170,N_4960,N_4864);
and U5171 (N_5171,N_4828,N_4823);
and U5172 (N_5172,N_4760,N_4850);
or U5173 (N_5173,N_4785,N_4825);
nor U5174 (N_5174,N_4918,N_4900);
xnor U5175 (N_5175,N_4805,N_4763);
and U5176 (N_5176,N_4784,N_4799);
nor U5177 (N_5177,N_4867,N_4827);
nor U5178 (N_5178,N_4802,N_4984);
or U5179 (N_5179,N_4796,N_4936);
nand U5180 (N_5180,N_4854,N_4842);
nand U5181 (N_5181,N_4794,N_4789);
xor U5182 (N_5182,N_4863,N_4995);
or U5183 (N_5183,N_4972,N_4788);
nor U5184 (N_5184,N_4843,N_4857);
xnor U5185 (N_5185,N_4855,N_4846);
nand U5186 (N_5186,N_4938,N_4802);
nor U5187 (N_5187,N_4799,N_4833);
nand U5188 (N_5188,N_4776,N_4999);
xnor U5189 (N_5189,N_4839,N_4784);
nand U5190 (N_5190,N_4803,N_4967);
nand U5191 (N_5191,N_4944,N_4986);
or U5192 (N_5192,N_4989,N_4979);
xor U5193 (N_5193,N_4916,N_4913);
or U5194 (N_5194,N_4807,N_4967);
xnor U5195 (N_5195,N_4840,N_4892);
or U5196 (N_5196,N_4970,N_4773);
nor U5197 (N_5197,N_4800,N_4774);
nor U5198 (N_5198,N_4976,N_4795);
nand U5199 (N_5199,N_4953,N_4957);
xnor U5200 (N_5200,N_4940,N_4867);
xor U5201 (N_5201,N_4782,N_4938);
nand U5202 (N_5202,N_4912,N_4918);
or U5203 (N_5203,N_4984,N_4771);
and U5204 (N_5204,N_4807,N_4974);
or U5205 (N_5205,N_4770,N_4790);
or U5206 (N_5206,N_4761,N_4821);
xor U5207 (N_5207,N_4910,N_4767);
nor U5208 (N_5208,N_4768,N_4802);
or U5209 (N_5209,N_4769,N_4887);
or U5210 (N_5210,N_4786,N_4763);
xor U5211 (N_5211,N_4752,N_4791);
nor U5212 (N_5212,N_4850,N_4863);
and U5213 (N_5213,N_4788,N_4902);
nor U5214 (N_5214,N_4824,N_4890);
and U5215 (N_5215,N_4789,N_4762);
and U5216 (N_5216,N_4919,N_4880);
and U5217 (N_5217,N_4976,N_4855);
nand U5218 (N_5218,N_4944,N_4931);
nor U5219 (N_5219,N_4970,N_4809);
and U5220 (N_5220,N_4767,N_4998);
nor U5221 (N_5221,N_4929,N_4857);
xnor U5222 (N_5222,N_4864,N_4795);
nand U5223 (N_5223,N_4823,N_4838);
xnor U5224 (N_5224,N_4993,N_4999);
and U5225 (N_5225,N_4986,N_4915);
nand U5226 (N_5226,N_4856,N_4808);
or U5227 (N_5227,N_4937,N_4823);
or U5228 (N_5228,N_4753,N_4752);
nor U5229 (N_5229,N_4771,N_4838);
nand U5230 (N_5230,N_4799,N_4919);
nor U5231 (N_5231,N_4884,N_4943);
xnor U5232 (N_5232,N_4967,N_4808);
xnor U5233 (N_5233,N_4783,N_4912);
xor U5234 (N_5234,N_4808,N_4817);
or U5235 (N_5235,N_4903,N_4789);
nand U5236 (N_5236,N_4862,N_4795);
xnor U5237 (N_5237,N_4867,N_4998);
xor U5238 (N_5238,N_4955,N_4952);
nand U5239 (N_5239,N_4918,N_4780);
and U5240 (N_5240,N_4754,N_4758);
and U5241 (N_5241,N_4939,N_4972);
nor U5242 (N_5242,N_4988,N_4973);
or U5243 (N_5243,N_4772,N_4806);
nor U5244 (N_5244,N_4844,N_4953);
and U5245 (N_5245,N_4887,N_4907);
and U5246 (N_5246,N_4818,N_4886);
xnor U5247 (N_5247,N_4786,N_4751);
and U5248 (N_5248,N_4759,N_4870);
xnor U5249 (N_5249,N_4910,N_4901);
nor U5250 (N_5250,N_5098,N_5206);
nand U5251 (N_5251,N_5009,N_5111);
and U5252 (N_5252,N_5107,N_5246);
nor U5253 (N_5253,N_5083,N_5093);
or U5254 (N_5254,N_5062,N_5142);
nor U5255 (N_5255,N_5140,N_5001);
xor U5256 (N_5256,N_5053,N_5036);
and U5257 (N_5257,N_5190,N_5041);
and U5258 (N_5258,N_5088,N_5248);
nand U5259 (N_5259,N_5004,N_5167);
or U5260 (N_5260,N_5050,N_5149);
and U5261 (N_5261,N_5236,N_5226);
nor U5262 (N_5262,N_5225,N_5085);
xnor U5263 (N_5263,N_5202,N_5034);
xor U5264 (N_5264,N_5019,N_5229);
xor U5265 (N_5265,N_5220,N_5101);
nor U5266 (N_5266,N_5227,N_5079);
xor U5267 (N_5267,N_5040,N_5201);
and U5268 (N_5268,N_5194,N_5123);
xor U5269 (N_5269,N_5104,N_5161);
and U5270 (N_5270,N_5165,N_5135);
nor U5271 (N_5271,N_5131,N_5143);
nor U5272 (N_5272,N_5221,N_5021);
nand U5273 (N_5273,N_5000,N_5211);
nand U5274 (N_5274,N_5162,N_5129);
and U5275 (N_5275,N_5081,N_5169);
or U5276 (N_5276,N_5058,N_5046);
and U5277 (N_5277,N_5109,N_5240);
xnor U5278 (N_5278,N_5061,N_5144);
nor U5279 (N_5279,N_5146,N_5137);
or U5280 (N_5280,N_5033,N_5159);
nand U5281 (N_5281,N_5056,N_5234);
xnor U5282 (N_5282,N_5178,N_5026);
and U5283 (N_5283,N_5064,N_5055);
or U5284 (N_5284,N_5097,N_5181);
or U5285 (N_5285,N_5022,N_5183);
and U5286 (N_5286,N_5207,N_5116);
nor U5287 (N_5287,N_5200,N_5139);
or U5288 (N_5288,N_5249,N_5080);
or U5289 (N_5289,N_5099,N_5007);
nand U5290 (N_5290,N_5071,N_5106);
or U5291 (N_5291,N_5032,N_5230);
nand U5292 (N_5292,N_5152,N_5044);
xor U5293 (N_5293,N_5084,N_5175);
or U5294 (N_5294,N_5112,N_5243);
and U5295 (N_5295,N_5160,N_5090);
nor U5296 (N_5296,N_5029,N_5209);
nand U5297 (N_5297,N_5065,N_5244);
nor U5298 (N_5298,N_5204,N_5070);
nor U5299 (N_5299,N_5002,N_5122);
nor U5300 (N_5300,N_5205,N_5128);
or U5301 (N_5301,N_5233,N_5072);
or U5302 (N_5302,N_5067,N_5196);
nand U5303 (N_5303,N_5133,N_5091);
nor U5304 (N_5304,N_5024,N_5006);
nor U5305 (N_5305,N_5018,N_5130);
nor U5306 (N_5306,N_5037,N_5245);
nand U5307 (N_5307,N_5223,N_5087);
or U5308 (N_5308,N_5115,N_5114);
xnor U5309 (N_5309,N_5075,N_5103);
nand U5310 (N_5310,N_5158,N_5108);
or U5311 (N_5311,N_5198,N_5125);
nor U5312 (N_5312,N_5185,N_5008);
or U5313 (N_5313,N_5020,N_5145);
nand U5314 (N_5314,N_5073,N_5012);
nor U5315 (N_5315,N_5141,N_5154);
xor U5316 (N_5316,N_5184,N_5192);
and U5317 (N_5317,N_5096,N_5164);
nand U5318 (N_5318,N_5110,N_5186);
or U5319 (N_5319,N_5124,N_5118);
nand U5320 (N_5320,N_5076,N_5082);
and U5321 (N_5321,N_5126,N_5176);
nor U5322 (N_5322,N_5031,N_5005);
and U5323 (N_5323,N_5014,N_5214);
nor U5324 (N_5324,N_5078,N_5238);
xor U5325 (N_5325,N_5188,N_5028);
and U5326 (N_5326,N_5048,N_5172);
xnor U5327 (N_5327,N_5195,N_5113);
nor U5328 (N_5328,N_5210,N_5136);
nor U5329 (N_5329,N_5049,N_5069);
or U5330 (N_5330,N_5003,N_5212);
or U5331 (N_5331,N_5177,N_5077);
and U5332 (N_5332,N_5057,N_5013);
nor U5333 (N_5333,N_5100,N_5222);
nor U5334 (N_5334,N_5016,N_5239);
xnor U5335 (N_5335,N_5120,N_5089);
nor U5336 (N_5336,N_5132,N_5231);
or U5337 (N_5337,N_5241,N_5155);
nor U5338 (N_5338,N_5199,N_5052);
nor U5339 (N_5339,N_5156,N_5213);
and U5340 (N_5340,N_5045,N_5237);
nand U5341 (N_5341,N_5102,N_5127);
xnor U5342 (N_5342,N_5074,N_5148);
nand U5343 (N_5343,N_5059,N_5039);
nand U5344 (N_5344,N_5066,N_5147);
xor U5345 (N_5345,N_5119,N_5151);
nand U5346 (N_5346,N_5197,N_5208);
nand U5347 (N_5347,N_5170,N_5010);
nor U5348 (N_5348,N_5138,N_5191);
and U5349 (N_5349,N_5173,N_5054);
xor U5350 (N_5350,N_5179,N_5011);
and U5351 (N_5351,N_5094,N_5166);
xor U5352 (N_5352,N_5015,N_5218);
and U5353 (N_5353,N_5051,N_5219);
nand U5354 (N_5354,N_5171,N_5117);
xor U5355 (N_5355,N_5086,N_5043);
or U5356 (N_5356,N_5157,N_5224);
or U5357 (N_5357,N_5105,N_5095);
and U5358 (N_5358,N_5121,N_5180);
and U5359 (N_5359,N_5232,N_5038);
or U5360 (N_5360,N_5092,N_5242);
nor U5361 (N_5361,N_5060,N_5134);
nor U5362 (N_5362,N_5182,N_5017);
or U5363 (N_5363,N_5153,N_5187);
and U5364 (N_5364,N_5025,N_5193);
or U5365 (N_5365,N_5163,N_5217);
or U5366 (N_5366,N_5215,N_5235);
and U5367 (N_5367,N_5203,N_5168);
nor U5368 (N_5368,N_5042,N_5068);
nor U5369 (N_5369,N_5228,N_5174);
and U5370 (N_5370,N_5027,N_5247);
nand U5371 (N_5371,N_5035,N_5030);
xor U5372 (N_5372,N_5023,N_5189);
xor U5373 (N_5373,N_5063,N_5216);
and U5374 (N_5374,N_5150,N_5047);
xor U5375 (N_5375,N_5123,N_5175);
nor U5376 (N_5376,N_5111,N_5022);
and U5377 (N_5377,N_5227,N_5202);
or U5378 (N_5378,N_5066,N_5182);
nand U5379 (N_5379,N_5195,N_5120);
nand U5380 (N_5380,N_5048,N_5044);
nor U5381 (N_5381,N_5045,N_5182);
nand U5382 (N_5382,N_5133,N_5018);
nor U5383 (N_5383,N_5229,N_5216);
xnor U5384 (N_5384,N_5204,N_5200);
nor U5385 (N_5385,N_5248,N_5126);
nand U5386 (N_5386,N_5083,N_5136);
nand U5387 (N_5387,N_5164,N_5217);
nor U5388 (N_5388,N_5134,N_5131);
nand U5389 (N_5389,N_5113,N_5075);
or U5390 (N_5390,N_5150,N_5221);
and U5391 (N_5391,N_5208,N_5194);
or U5392 (N_5392,N_5014,N_5211);
nor U5393 (N_5393,N_5230,N_5020);
xnor U5394 (N_5394,N_5173,N_5163);
and U5395 (N_5395,N_5119,N_5044);
nand U5396 (N_5396,N_5003,N_5198);
nand U5397 (N_5397,N_5139,N_5007);
nand U5398 (N_5398,N_5038,N_5017);
nor U5399 (N_5399,N_5064,N_5233);
or U5400 (N_5400,N_5162,N_5144);
nand U5401 (N_5401,N_5094,N_5225);
xnor U5402 (N_5402,N_5105,N_5150);
and U5403 (N_5403,N_5171,N_5204);
or U5404 (N_5404,N_5031,N_5148);
or U5405 (N_5405,N_5023,N_5087);
nand U5406 (N_5406,N_5106,N_5060);
or U5407 (N_5407,N_5068,N_5113);
xor U5408 (N_5408,N_5056,N_5094);
or U5409 (N_5409,N_5087,N_5115);
nor U5410 (N_5410,N_5222,N_5192);
nor U5411 (N_5411,N_5095,N_5164);
nor U5412 (N_5412,N_5212,N_5029);
nand U5413 (N_5413,N_5192,N_5051);
nand U5414 (N_5414,N_5002,N_5021);
nor U5415 (N_5415,N_5111,N_5032);
xor U5416 (N_5416,N_5053,N_5182);
nor U5417 (N_5417,N_5136,N_5094);
nor U5418 (N_5418,N_5217,N_5107);
and U5419 (N_5419,N_5029,N_5099);
nor U5420 (N_5420,N_5170,N_5062);
nor U5421 (N_5421,N_5126,N_5199);
nand U5422 (N_5422,N_5082,N_5043);
nor U5423 (N_5423,N_5199,N_5023);
and U5424 (N_5424,N_5114,N_5245);
xor U5425 (N_5425,N_5225,N_5109);
nor U5426 (N_5426,N_5247,N_5188);
and U5427 (N_5427,N_5075,N_5193);
or U5428 (N_5428,N_5038,N_5013);
nor U5429 (N_5429,N_5160,N_5174);
nand U5430 (N_5430,N_5224,N_5019);
xor U5431 (N_5431,N_5192,N_5151);
nor U5432 (N_5432,N_5178,N_5051);
or U5433 (N_5433,N_5192,N_5216);
xnor U5434 (N_5434,N_5112,N_5219);
and U5435 (N_5435,N_5098,N_5045);
nand U5436 (N_5436,N_5179,N_5153);
nor U5437 (N_5437,N_5077,N_5240);
xnor U5438 (N_5438,N_5097,N_5171);
nor U5439 (N_5439,N_5014,N_5072);
nand U5440 (N_5440,N_5180,N_5048);
nand U5441 (N_5441,N_5205,N_5061);
and U5442 (N_5442,N_5012,N_5211);
or U5443 (N_5443,N_5218,N_5038);
and U5444 (N_5444,N_5244,N_5164);
nor U5445 (N_5445,N_5150,N_5177);
xnor U5446 (N_5446,N_5212,N_5247);
nand U5447 (N_5447,N_5037,N_5110);
xnor U5448 (N_5448,N_5005,N_5243);
xor U5449 (N_5449,N_5204,N_5037);
or U5450 (N_5450,N_5176,N_5242);
nor U5451 (N_5451,N_5144,N_5088);
nor U5452 (N_5452,N_5227,N_5136);
xnor U5453 (N_5453,N_5192,N_5066);
nand U5454 (N_5454,N_5227,N_5167);
nand U5455 (N_5455,N_5103,N_5102);
nor U5456 (N_5456,N_5179,N_5087);
nand U5457 (N_5457,N_5156,N_5082);
or U5458 (N_5458,N_5129,N_5245);
or U5459 (N_5459,N_5203,N_5064);
and U5460 (N_5460,N_5170,N_5015);
xnor U5461 (N_5461,N_5245,N_5108);
nand U5462 (N_5462,N_5040,N_5245);
xor U5463 (N_5463,N_5129,N_5112);
nand U5464 (N_5464,N_5045,N_5189);
or U5465 (N_5465,N_5242,N_5002);
xnor U5466 (N_5466,N_5180,N_5087);
and U5467 (N_5467,N_5148,N_5172);
and U5468 (N_5468,N_5036,N_5052);
nand U5469 (N_5469,N_5231,N_5083);
or U5470 (N_5470,N_5070,N_5194);
nor U5471 (N_5471,N_5016,N_5142);
xor U5472 (N_5472,N_5099,N_5136);
nor U5473 (N_5473,N_5044,N_5144);
and U5474 (N_5474,N_5121,N_5186);
and U5475 (N_5475,N_5017,N_5161);
and U5476 (N_5476,N_5073,N_5140);
and U5477 (N_5477,N_5192,N_5016);
and U5478 (N_5478,N_5138,N_5030);
nor U5479 (N_5479,N_5012,N_5008);
xnor U5480 (N_5480,N_5027,N_5055);
and U5481 (N_5481,N_5139,N_5224);
xnor U5482 (N_5482,N_5055,N_5089);
nor U5483 (N_5483,N_5117,N_5192);
or U5484 (N_5484,N_5077,N_5159);
nor U5485 (N_5485,N_5096,N_5011);
and U5486 (N_5486,N_5019,N_5045);
and U5487 (N_5487,N_5195,N_5119);
or U5488 (N_5488,N_5240,N_5168);
or U5489 (N_5489,N_5214,N_5146);
nand U5490 (N_5490,N_5214,N_5077);
nor U5491 (N_5491,N_5081,N_5053);
and U5492 (N_5492,N_5117,N_5106);
nand U5493 (N_5493,N_5191,N_5148);
and U5494 (N_5494,N_5157,N_5196);
nor U5495 (N_5495,N_5032,N_5069);
nand U5496 (N_5496,N_5018,N_5106);
nand U5497 (N_5497,N_5174,N_5242);
xnor U5498 (N_5498,N_5039,N_5198);
or U5499 (N_5499,N_5107,N_5236);
and U5500 (N_5500,N_5288,N_5454);
or U5501 (N_5501,N_5415,N_5400);
and U5502 (N_5502,N_5303,N_5362);
nor U5503 (N_5503,N_5447,N_5422);
and U5504 (N_5504,N_5485,N_5356);
nor U5505 (N_5505,N_5265,N_5274);
or U5506 (N_5506,N_5459,N_5340);
or U5507 (N_5507,N_5461,N_5359);
and U5508 (N_5508,N_5466,N_5438);
and U5509 (N_5509,N_5278,N_5441);
nand U5510 (N_5510,N_5373,N_5478);
xor U5511 (N_5511,N_5457,N_5368);
and U5512 (N_5512,N_5488,N_5260);
or U5513 (N_5513,N_5403,N_5435);
nand U5514 (N_5514,N_5264,N_5431);
or U5515 (N_5515,N_5463,N_5483);
and U5516 (N_5516,N_5292,N_5452);
nor U5517 (N_5517,N_5273,N_5487);
xnor U5518 (N_5518,N_5439,N_5381);
xor U5519 (N_5519,N_5370,N_5277);
and U5520 (N_5520,N_5257,N_5304);
or U5521 (N_5521,N_5331,N_5378);
and U5522 (N_5522,N_5396,N_5448);
and U5523 (N_5523,N_5460,N_5271);
nand U5524 (N_5524,N_5491,N_5261);
and U5525 (N_5525,N_5468,N_5456);
xor U5526 (N_5526,N_5464,N_5253);
nand U5527 (N_5527,N_5315,N_5290);
nand U5528 (N_5528,N_5345,N_5424);
nor U5529 (N_5529,N_5286,N_5436);
nor U5530 (N_5530,N_5280,N_5379);
and U5531 (N_5531,N_5302,N_5285);
nand U5532 (N_5532,N_5332,N_5446);
and U5533 (N_5533,N_5371,N_5372);
or U5534 (N_5534,N_5440,N_5406);
or U5535 (N_5535,N_5481,N_5350);
nor U5536 (N_5536,N_5430,N_5275);
xor U5537 (N_5537,N_5327,N_5484);
xnor U5538 (N_5538,N_5364,N_5429);
nand U5539 (N_5539,N_5495,N_5357);
nor U5540 (N_5540,N_5311,N_5320);
xor U5541 (N_5541,N_5269,N_5348);
or U5542 (N_5542,N_5480,N_5252);
xor U5543 (N_5543,N_5449,N_5308);
or U5544 (N_5544,N_5262,N_5462);
nand U5545 (N_5545,N_5313,N_5266);
nor U5546 (N_5546,N_5316,N_5344);
nor U5547 (N_5547,N_5453,N_5374);
nand U5548 (N_5548,N_5305,N_5420);
or U5549 (N_5549,N_5391,N_5337);
and U5550 (N_5550,N_5319,N_5479);
and U5551 (N_5551,N_5296,N_5499);
xor U5552 (N_5552,N_5476,N_5455);
nand U5553 (N_5553,N_5390,N_5465);
xnor U5554 (N_5554,N_5318,N_5301);
nor U5555 (N_5555,N_5492,N_5380);
or U5556 (N_5556,N_5343,N_5346);
nand U5557 (N_5557,N_5494,N_5404);
xor U5558 (N_5558,N_5423,N_5467);
or U5559 (N_5559,N_5409,N_5291);
or U5560 (N_5560,N_5333,N_5433);
and U5561 (N_5561,N_5298,N_5360);
xnor U5562 (N_5562,N_5411,N_5402);
xor U5563 (N_5563,N_5375,N_5407);
nand U5564 (N_5564,N_5419,N_5351);
xnor U5565 (N_5565,N_5472,N_5369);
nor U5566 (N_5566,N_5498,N_5255);
or U5567 (N_5567,N_5425,N_5386);
nor U5568 (N_5568,N_5270,N_5489);
or U5569 (N_5569,N_5477,N_5437);
and U5570 (N_5570,N_5383,N_5287);
or U5571 (N_5571,N_5254,N_5324);
xor U5572 (N_5572,N_5470,N_5282);
nor U5573 (N_5573,N_5307,N_5401);
and U5574 (N_5574,N_5317,N_5377);
xnor U5575 (N_5575,N_5334,N_5445);
nand U5576 (N_5576,N_5289,N_5300);
and U5577 (N_5577,N_5363,N_5493);
nor U5578 (N_5578,N_5496,N_5325);
xnor U5579 (N_5579,N_5358,N_5310);
nand U5580 (N_5580,N_5392,N_5418);
xor U5581 (N_5581,N_5354,N_5284);
xnor U5582 (N_5582,N_5427,N_5323);
nor U5583 (N_5583,N_5469,N_5294);
and U5584 (N_5584,N_5421,N_5394);
and U5585 (N_5585,N_5426,N_5342);
or U5586 (N_5586,N_5432,N_5434);
xnor U5587 (N_5587,N_5376,N_5443);
xnor U5588 (N_5588,N_5338,N_5471);
and U5589 (N_5589,N_5329,N_5251);
nand U5590 (N_5590,N_5295,N_5328);
nand U5591 (N_5591,N_5416,N_5412);
xnor U5592 (N_5592,N_5417,N_5428);
nor U5593 (N_5593,N_5475,N_5474);
and U5594 (N_5594,N_5250,N_5450);
nor U5595 (N_5595,N_5388,N_5312);
or U5596 (N_5596,N_5408,N_5321);
and U5597 (N_5597,N_5293,N_5281);
nand U5598 (N_5598,N_5355,N_5347);
and U5599 (N_5599,N_5393,N_5263);
nor U5600 (N_5600,N_5444,N_5410);
and U5601 (N_5601,N_5384,N_5339);
nor U5602 (N_5602,N_5387,N_5361);
or U5603 (N_5603,N_5276,N_5397);
or U5604 (N_5604,N_5330,N_5299);
nand U5605 (N_5605,N_5365,N_5399);
nand U5606 (N_5606,N_5314,N_5322);
xnor U5607 (N_5607,N_5395,N_5336);
and U5608 (N_5608,N_5306,N_5497);
xor U5609 (N_5609,N_5473,N_5482);
nor U5610 (N_5610,N_5458,N_5353);
nand U5611 (N_5611,N_5405,N_5258);
xor U5612 (N_5612,N_5366,N_5382);
or U5613 (N_5613,N_5385,N_5442);
nor U5614 (N_5614,N_5341,N_5451);
nand U5615 (N_5615,N_5413,N_5267);
xor U5616 (N_5616,N_5283,N_5279);
nand U5617 (N_5617,N_5309,N_5367);
xnor U5618 (N_5618,N_5259,N_5272);
xor U5619 (N_5619,N_5326,N_5414);
nor U5620 (N_5620,N_5268,N_5352);
and U5621 (N_5621,N_5349,N_5335);
and U5622 (N_5622,N_5398,N_5389);
and U5623 (N_5623,N_5256,N_5486);
or U5624 (N_5624,N_5297,N_5490);
and U5625 (N_5625,N_5403,N_5490);
or U5626 (N_5626,N_5411,N_5347);
xnor U5627 (N_5627,N_5388,N_5436);
xnor U5628 (N_5628,N_5450,N_5354);
nor U5629 (N_5629,N_5397,N_5452);
nand U5630 (N_5630,N_5388,N_5351);
xor U5631 (N_5631,N_5372,N_5461);
nor U5632 (N_5632,N_5430,N_5470);
or U5633 (N_5633,N_5298,N_5374);
or U5634 (N_5634,N_5461,N_5424);
nor U5635 (N_5635,N_5278,N_5422);
nand U5636 (N_5636,N_5252,N_5386);
nand U5637 (N_5637,N_5429,N_5424);
and U5638 (N_5638,N_5399,N_5267);
xor U5639 (N_5639,N_5271,N_5259);
nor U5640 (N_5640,N_5301,N_5492);
or U5641 (N_5641,N_5307,N_5473);
or U5642 (N_5642,N_5485,N_5361);
and U5643 (N_5643,N_5349,N_5359);
xor U5644 (N_5644,N_5438,N_5250);
or U5645 (N_5645,N_5251,N_5346);
nand U5646 (N_5646,N_5311,N_5499);
and U5647 (N_5647,N_5452,N_5297);
or U5648 (N_5648,N_5356,N_5447);
nor U5649 (N_5649,N_5434,N_5447);
or U5650 (N_5650,N_5389,N_5309);
and U5651 (N_5651,N_5311,N_5263);
or U5652 (N_5652,N_5471,N_5424);
and U5653 (N_5653,N_5266,N_5435);
nand U5654 (N_5654,N_5255,N_5293);
nand U5655 (N_5655,N_5326,N_5446);
and U5656 (N_5656,N_5296,N_5363);
or U5657 (N_5657,N_5489,N_5259);
and U5658 (N_5658,N_5327,N_5309);
nor U5659 (N_5659,N_5404,N_5484);
nand U5660 (N_5660,N_5270,N_5394);
nand U5661 (N_5661,N_5281,N_5294);
xnor U5662 (N_5662,N_5444,N_5428);
nand U5663 (N_5663,N_5319,N_5387);
xor U5664 (N_5664,N_5325,N_5395);
or U5665 (N_5665,N_5317,N_5458);
nor U5666 (N_5666,N_5278,N_5373);
or U5667 (N_5667,N_5312,N_5250);
xnor U5668 (N_5668,N_5440,N_5306);
and U5669 (N_5669,N_5351,N_5473);
nand U5670 (N_5670,N_5415,N_5333);
nor U5671 (N_5671,N_5476,N_5261);
xor U5672 (N_5672,N_5412,N_5438);
nor U5673 (N_5673,N_5285,N_5291);
nand U5674 (N_5674,N_5427,N_5333);
or U5675 (N_5675,N_5351,N_5492);
xnor U5676 (N_5676,N_5254,N_5445);
and U5677 (N_5677,N_5316,N_5466);
xor U5678 (N_5678,N_5438,N_5480);
and U5679 (N_5679,N_5290,N_5267);
xor U5680 (N_5680,N_5411,N_5447);
nor U5681 (N_5681,N_5297,N_5270);
nand U5682 (N_5682,N_5460,N_5399);
or U5683 (N_5683,N_5448,N_5274);
xor U5684 (N_5684,N_5257,N_5252);
or U5685 (N_5685,N_5417,N_5379);
or U5686 (N_5686,N_5416,N_5362);
and U5687 (N_5687,N_5255,N_5451);
or U5688 (N_5688,N_5364,N_5448);
nor U5689 (N_5689,N_5260,N_5313);
and U5690 (N_5690,N_5327,N_5315);
xnor U5691 (N_5691,N_5417,N_5434);
nand U5692 (N_5692,N_5477,N_5272);
nor U5693 (N_5693,N_5370,N_5468);
xor U5694 (N_5694,N_5451,N_5365);
nor U5695 (N_5695,N_5288,N_5298);
and U5696 (N_5696,N_5490,N_5357);
nor U5697 (N_5697,N_5284,N_5297);
nand U5698 (N_5698,N_5320,N_5393);
nor U5699 (N_5699,N_5297,N_5341);
nor U5700 (N_5700,N_5255,N_5364);
or U5701 (N_5701,N_5372,N_5291);
xor U5702 (N_5702,N_5258,N_5254);
nor U5703 (N_5703,N_5316,N_5349);
or U5704 (N_5704,N_5447,N_5297);
nand U5705 (N_5705,N_5413,N_5462);
nor U5706 (N_5706,N_5390,N_5300);
and U5707 (N_5707,N_5284,N_5401);
nand U5708 (N_5708,N_5412,N_5495);
or U5709 (N_5709,N_5458,N_5436);
or U5710 (N_5710,N_5300,N_5407);
nor U5711 (N_5711,N_5299,N_5483);
or U5712 (N_5712,N_5296,N_5435);
and U5713 (N_5713,N_5454,N_5264);
xor U5714 (N_5714,N_5301,N_5250);
nand U5715 (N_5715,N_5340,N_5288);
xnor U5716 (N_5716,N_5436,N_5330);
xor U5717 (N_5717,N_5429,N_5320);
or U5718 (N_5718,N_5477,N_5326);
nor U5719 (N_5719,N_5347,N_5337);
nand U5720 (N_5720,N_5442,N_5271);
nor U5721 (N_5721,N_5299,N_5485);
nor U5722 (N_5722,N_5446,N_5408);
or U5723 (N_5723,N_5325,N_5427);
or U5724 (N_5724,N_5396,N_5416);
or U5725 (N_5725,N_5266,N_5321);
nor U5726 (N_5726,N_5432,N_5362);
nor U5727 (N_5727,N_5281,N_5317);
nand U5728 (N_5728,N_5444,N_5344);
and U5729 (N_5729,N_5272,N_5311);
or U5730 (N_5730,N_5474,N_5275);
and U5731 (N_5731,N_5374,N_5312);
nor U5732 (N_5732,N_5356,N_5263);
or U5733 (N_5733,N_5354,N_5499);
nor U5734 (N_5734,N_5474,N_5311);
and U5735 (N_5735,N_5477,N_5430);
nor U5736 (N_5736,N_5313,N_5448);
and U5737 (N_5737,N_5495,N_5405);
and U5738 (N_5738,N_5384,N_5459);
xor U5739 (N_5739,N_5333,N_5455);
and U5740 (N_5740,N_5275,N_5350);
nand U5741 (N_5741,N_5340,N_5296);
or U5742 (N_5742,N_5336,N_5309);
nand U5743 (N_5743,N_5293,N_5282);
or U5744 (N_5744,N_5307,N_5315);
nor U5745 (N_5745,N_5430,N_5414);
or U5746 (N_5746,N_5368,N_5382);
xor U5747 (N_5747,N_5290,N_5364);
nand U5748 (N_5748,N_5313,N_5470);
or U5749 (N_5749,N_5498,N_5290);
xor U5750 (N_5750,N_5529,N_5694);
nand U5751 (N_5751,N_5567,N_5548);
and U5752 (N_5752,N_5738,N_5592);
and U5753 (N_5753,N_5615,N_5576);
and U5754 (N_5754,N_5616,N_5698);
and U5755 (N_5755,N_5561,N_5525);
nor U5756 (N_5756,N_5749,N_5530);
nor U5757 (N_5757,N_5507,N_5685);
nor U5758 (N_5758,N_5634,N_5500);
xnor U5759 (N_5759,N_5640,N_5716);
nor U5760 (N_5760,N_5725,N_5612);
nor U5761 (N_5761,N_5723,N_5601);
and U5762 (N_5762,N_5538,N_5627);
nor U5763 (N_5763,N_5652,N_5546);
nand U5764 (N_5764,N_5644,N_5720);
xnor U5765 (N_5765,N_5669,N_5633);
and U5766 (N_5766,N_5599,N_5721);
and U5767 (N_5767,N_5635,N_5605);
and U5768 (N_5768,N_5728,N_5501);
and U5769 (N_5769,N_5580,N_5586);
or U5770 (N_5770,N_5717,N_5512);
and U5771 (N_5771,N_5731,N_5682);
nand U5772 (N_5772,N_5547,N_5691);
or U5773 (N_5773,N_5664,N_5674);
nor U5774 (N_5774,N_5671,N_5637);
and U5775 (N_5775,N_5630,N_5670);
nand U5776 (N_5776,N_5541,N_5587);
or U5777 (N_5777,N_5503,N_5724);
nor U5778 (N_5778,N_5729,N_5710);
nor U5779 (N_5779,N_5647,N_5735);
and U5780 (N_5780,N_5636,N_5504);
nor U5781 (N_5781,N_5509,N_5539);
nor U5782 (N_5782,N_5524,N_5549);
xnor U5783 (N_5783,N_5632,N_5642);
or U5784 (N_5784,N_5563,N_5643);
xnor U5785 (N_5785,N_5718,N_5703);
nand U5786 (N_5786,N_5641,N_5534);
nand U5787 (N_5787,N_5619,N_5590);
or U5788 (N_5788,N_5528,N_5745);
nand U5789 (N_5789,N_5543,N_5727);
and U5790 (N_5790,N_5571,N_5626);
xor U5791 (N_5791,N_5617,N_5657);
nor U5792 (N_5792,N_5741,N_5689);
or U5793 (N_5793,N_5579,N_5715);
nor U5794 (N_5794,N_5589,N_5654);
or U5795 (N_5795,N_5701,N_5552);
or U5796 (N_5796,N_5740,N_5709);
nor U5797 (N_5797,N_5742,N_5712);
nand U5798 (N_5798,N_5692,N_5648);
nand U5799 (N_5799,N_5734,N_5609);
and U5800 (N_5800,N_5747,N_5575);
or U5801 (N_5801,N_5722,N_5744);
nor U5802 (N_5802,N_5620,N_5660);
xnor U5803 (N_5803,N_5551,N_5677);
nand U5804 (N_5804,N_5678,N_5676);
nor U5805 (N_5805,N_5555,N_5679);
xor U5806 (N_5806,N_5667,N_5697);
nand U5807 (N_5807,N_5683,N_5553);
or U5808 (N_5808,N_5600,N_5520);
and U5809 (N_5809,N_5540,N_5628);
or U5810 (N_5810,N_5655,N_5699);
and U5811 (N_5811,N_5514,N_5577);
and U5812 (N_5812,N_5550,N_5638);
nor U5813 (N_5813,N_5613,N_5610);
and U5814 (N_5814,N_5526,N_5663);
nor U5815 (N_5815,N_5560,N_5690);
and U5816 (N_5816,N_5523,N_5746);
nor U5817 (N_5817,N_5522,N_5649);
nand U5818 (N_5818,N_5595,N_5516);
and U5819 (N_5819,N_5673,N_5608);
nand U5820 (N_5820,N_5726,N_5533);
and U5821 (N_5821,N_5645,N_5506);
or U5822 (N_5822,N_5656,N_5598);
or U5823 (N_5823,N_5545,N_5582);
nor U5824 (N_5824,N_5733,N_5536);
nand U5825 (N_5825,N_5719,N_5659);
and U5826 (N_5826,N_5508,N_5650);
and U5827 (N_5827,N_5743,N_5565);
xor U5828 (N_5828,N_5624,N_5537);
nand U5829 (N_5829,N_5531,N_5702);
or U5830 (N_5830,N_5518,N_5629);
and U5831 (N_5831,N_5578,N_5597);
nor U5832 (N_5832,N_5625,N_5708);
or U5833 (N_5833,N_5510,N_5519);
or U5834 (N_5834,N_5662,N_5700);
nand U5835 (N_5835,N_5696,N_5631);
nand U5836 (N_5836,N_5713,N_5603);
or U5837 (N_5837,N_5588,N_5535);
or U5838 (N_5838,N_5688,N_5739);
xor U5839 (N_5839,N_5730,N_5604);
or U5840 (N_5840,N_5668,N_5618);
nand U5841 (N_5841,N_5748,N_5693);
and U5842 (N_5842,N_5570,N_5594);
nor U5843 (N_5843,N_5711,N_5707);
nand U5844 (N_5844,N_5658,N_5513);
or U5845 (N_5845,N_5665,N_5542);
nor U5846 (N_5846,N_5593,N_5651);
nand U5847 (N_5847,N_5675,N_5661);
or U5848 (N_5848,N_5602,N_5544);
and U5849 (N_5849,N_5585,N_5705);
xnor U5850 (N_5850,N_5532,N_5607);
and U5851 (N_5851,N_5622,N_5515);
nand U5852 (N_5852,N_5606,N_5505);
nor U5853 (N_5853,N_5687,N_5556);
and U5854 (N_5854,N_5564,N_5517);
nand U5855 (N_5855,N_5574,N_5584);
or U5856 (N_5856,N_5695,N_5557);
nand U5857 (N_5857,N_5639,N_5573);
nor U5858 (N_5858,N_5732,N_5572);
nand U5859 (N_5859,N_5591,N_5653);
or U5860 (N_5860,N_5502,N_5623);
nor U5861 (N_5861,N_5511,N_5704);
or U5862 (N_5862,N_5737,N_5568);
nand U5863 (N_5863,N_5566,N_5672);
nor U5864 (N_5864,N_5569,N_5521);
nand U5865 (N_5865,N_5611,N_5559);
xnor U5866 (N_5866,N_5583,N_5558);
and U5867 (N_5867,N_5714,N_5614);
nor U5868 (N_5868,N_5562,N_5646);
xor U5869 (N_5869,N_5686,N_5666);
and U5870 (N_5870,N_5680,N_5621);
and U5871 (N_5871,N_5554,N_5681);
nor U5872 (N_5872,N_5596,N_5527);
or U5873 (N_5873,N_5684,N_5581);
nand U5874 (N_5874,N_5736,N_5706);
and U5875 (N_5875,N_5587,N_5686);
or U5876 (N_5876,N_5508,N_5616);
nor U5877 (N_5877,N_5626,N_5688);
or U5878 (N_5878,N_5595,N_5610);
nand U5879 (N_5879,N_5605,N_5530);
or U5880 (N_5880,N_5683,N_5501);
or U5881 (N_5881,N_5667,N_5665);
and U5882 (N_5882,N_5702,N_5602);
and U5883 (N_5883,N_5682,N_5506);
nor U5884 (N_5884,N_5726,N_5724);
xnor U5885 (N_5885,N_5582,N_5577);
nor U5886 (N_5886,N_5723,N_5531);
and U5887 (N_5887,N_5680,N_5707);
nand U5888 (N_5888,N_5515,N_5513);
and U5889 (N_5889,N_5724,N_5599);
or U5890 (N_5890,N_5649,N_5628);
nand U5891 (N_5891,N_5526,N_5642);
and U5892 (N_5892,N_5540,N_5726);
nor U5893 (N_5893,N_5688,N_5645);
or U5894 (N_5894,N_5706,N_5559);
nand U5895 (N_5895,N_5664,N_5587);
nand U5896 (N_5896,N_5660,N_5696);
nand U5897 (N_5897,N_5642,N_5672);
nand U5898 (N_5898,N_5736,N_5546);
nor U5899 (N_5899,N_5723,N_5618);
and U5900 (N_5900,N_5656,N_5672);
and U5901 (N_5901,N_5528,N_5601);
nand U5902 (N_5902,N_5712,N_5599);
xor U5903 (N_5903,N_5708,N_5623);
or U5904 (N_5904,N_5707,N_5572);
xnor U5905 (N_5905,N_5641,N_5740);
nor U5906 (N_5906,N_5540,N_5644);
and U5907 (N_5907,N_5700,N_5555);
and U5908 (N_5908,N_5591,N_5616);
and U5909 (N_5909,N_5584,N_5569);
and U5910 (N_5910,N_5507,N_5632);
or U5911 (N_5911,N_5746,N_5514);
and U5912 (N_5912,N_5661,N_5608);
nor U5913 (N_5913,N_5657,N_5699);
nor U5914 (N_5914,N_5530,N_5659);
and U5915 (N_5915,N_5535,N_5691);
and U5916 (N_5916,N_5537,N_5661);
nor U5917 (N_5917,N_5731,N_5508);
nor U5918 (N_5918,N_5622,N_5532);
or U5919 (N_5919,N_5639,N_5510);
nand U5920 (N_5920,N_5571,N_5588);
xnor U5921 (N_5921,N_5714,N_5652);
nand U5922 (N_5922,N_5600,N_5566);
nor U5923 (N_5923,N_5566,N_5742);
nand U5924 (N_5924,N_5568,N_5567);
xor U5925 (N_5925,N_5745,N_5640);
nor U5926 (N_5926,N_5672,N_5673);
and U5927 (N_5927,N_5565,N_5721);
nor U5928 (N_5928,N_5696,N_5622);
or U5929 (N_5929,N_5743,N_5571);
nand U5930 (N_5930,N_5604,N_5653);
or U5931 (N_5931,N_5613,N_5666);
or U5932 (N_5932,N_5502,N_5688);
xor U5933 (N_5933,N_5531,N_5537);
nand U5934 (N_5934,N_5712,N_5540);
or U5935 (N_5935,N_5697,N_5592);
nor U5936 (N_5936,N_5642,N_5537);
nand U5937 (N_5937,N_5708,N_5657);
xor U5938 (N_5938,N_5651,N_5523);
nand U5939 (N_5939,N_5623,N_5597);
nand U5940 (N_5940,N_5659,N_5633);
and U5941 (N_5941,N_5530,N_5692);
and U5942 (N_5942,N_5612,N_5742);
or U5943 (N_5943,N_5571,N_5670);
nand U5944 (N_5944,N_5622,N_5602);
and U5945 (N_5945,N_5642,N_5728);
and U5946 (N_5946,N_5718,N_5729);
or U5947 (N_5947,N_5720,N_5521);
xor U5948 (N_5948,N_5671,N_5532);
nand U5949 (N_5949,N_5524,N_5721);
and U5950 (N_5950,N_5631,N_5695);
nand U5951 (N_5951,N_5686,N_5650);
or U5952 (N_5952,N_5710,N_5657);
xnor U5953 (N_5953,N_5673,N_5526);
or U5954 (N_5954,N_5587,N_5621);
or U5955 (N_5955,N_5522,N_5717);
or U5956 (N_5956,N_5630,N_5676);
nand U5957 (N_5957,N_5524,N_5540);
xor U5958 (N_5958,N_5595,N_5512);
and U5959 (N_5959,N_5560,N_5692);
and U5960 (N_5960,N_5671,N_5549);
nand U5961 (N_5961,N_5669,N_5716);
xor U5962 (N_5962,N_5637,N_5718);
nand U5963 (N_5963,N_5551,N_5614);
xor U5964 (N_5964,N_5650,N_5536);
nor U5965 (N_5965,N_5574,N_5577);
nor U5966 (N_5966,N_5533,N_5505);
and U5967 (N_5967,N_5716,N_5703);
nand U5968 (N_5968,N_5548,N_5716);
and U5969 (N_5969,N_5533,N_5619);
or U5970 (N_5970,N_5520,N_5725);
xor U5971 (N_5971,N_5640,N_5648);
nor U5972 (N_5972,N_5529,N_5678);
nor U5973 (N_5973,N_5709,N_5538);
nand U5974 (N_5974,N_5634,N_5568);
nand U5975 (N_5975,N_5520,N_5581);
and U5976 (N_5976,N_5690,N_5611);
or U5977 (N_5977,N_5678,N_5628);
or U5978 (N_5978,N_5548,N_5544);
xor U5979 (N_5979,N_5663,N_5551);
xor U5980 (N_5980,N_5717,N_5530);
nand U5981 (N_5981,N_5616,N_5542);
nand U5982 (N_5982,N_5532,N_5678);
or U5983 (N_5983,N_5731,N_5669);
xnor U5984 (N_5984,N_5654,N_5681);
nand U5985 (N_5985,N_5730,N_5571);
nor U5986 (N_5986,N_5634,N_5722);
xor U5987 (N_5987,N_5544,N_5572);
and U5988 (N_5988,N_5716,N_5577);
nor U5989 (N_5989,N_5726,N_5522);
xnor U5990 (N_5990,N_5519,N_5568);
nor U5991 (N_5991,N_5671,N_5552);
or U5992 (N_5992,N_5635,N_5510);
or U5993 (N_5993,N_5604,N_5520);
nand U5994 (N_5994,N_5540,N_5589);
and U5995 (N_5995,N_5591,N_5544);
and U5996 (N_5996,N_5553,N_5685);
nor U5997 (N_5997,N_5572,N_5727);
xor U5998 (N_5998,N_5665,N_5611);
nand U5999 (N_5999,N_5501,N_5588);
xor U6000 (N_6000,N_5975,N_5764);
nand U6001 (N_6001,N_5838,N_5790);
nor U6002 (N_6002,N_5769,N_5841);
nand U6003 (N_6003,N_5781,N_5852);
nand U6004 (N_6004,N_5960,N_5759);
nor U6005 (N_6005,N_5878,N_5779);
xnor U6006 (N_6006,N_5798,N_5983);
xor U6007 (N_6007,N_5865,N_5892);
and U6008 (N_6008,N_5846,N_5965);
and U6009 (N_6009,N_5847,N_5949);
nor U6010 (N_6010,N_5929,N_5782);
and U6011 (N_6011,N_5791,N_5848);
or U6012 (N_6012,N_5986,N_5925);
nor U6013 (N_6013,N_5922,N_5807);
and U6014 (N_6014,N_5944,N_5997);
nand U6015 (N_6015,N_5817,N_5858);
nor U6016 (N_6016,N_5973,N_5873);
nor U6017 (N_6017,N_5753,N_5953);
xnor U6018 (N_6018,N_5832,N_5978);
nor U6019 (N_6019,N_5976,N_5824);
and U6020 (N_6020,N_5950,N_5926);
or U6021 (N_6021,N_5979,N_5971);
or U6022 (N_6022,N_5884,N_5876);
or U6023 (N_6023,N_5947,N_5801);
nand U6024 (N_6024,N_5886,N_5906);
xnor U6025 (N_6025,N_5845,N_5933);
or U6026 (N_6026,N_5877,N_5943);
xor U6027 (N_6027,N_5834,N_5895);
nand U6028 (N_6028,N_5859,N_5797);
nand U6029 (N_6029,N_5889,N_5890);
or U6030 (N_6030,N_5962,N_5868);
nor U6031 (N_6031,N_5785,N_5830);
and U6032 (N_6032,N_5980,N_5989);
or U6033 (N_6033,N_5816,N_5970);
nand U6034 (N_6034,N_5789,N_5918);
nor U6035 (N_6035,N_5800,N_5901);
nor U6036 (N_6036,N_5957,N_5823);
and U6037 (N_6037,N_5840,N_5869);
or U6038 (N_6038,N_5945,N_5977);
nand U6039 (N_6039,N_5972,N_5793);
and U6040 (N_6040,N_5760,N_5930);
xnor U6041 (N_6041,N_5818,N_5828);
and U6042 (N_6042,N_5750,N_5754);
xor U6043 (N_6043,N_5941,N_5870);
xor U6044 (N_6044,N_5780,N_5829);
xor U6045 (N_6045,N_5827,N_5912);
xor U6046 (N_6046,N_5855,N_5826);
nor U6047 (N_6047,N_5887,N_5773);
nor U6048 (N_6048,N_5784,N_5851);
nand U6049 (N_6049,N_5821,N_5996);
nand U6050 (N_6050,N_5844,N_5920);
xnor U6051 (N_6051,N_5936,N_5776);
nand U6052 (N_6052,N_5905,N_5874);
xnor U6053 (N_6053,N_5835,N_5880);
xnor U6054 (N_6054,N_5908,N_5778);
nor U6055 (N_6055,N_5861,N_5775);
xnor U6056 (N_6056,N_5963,N_5893);
or U6057 (N_6057,N_5871,N_5898);
nand U6058 (N_6058,N_5899,N_5909);
or U6059 (N_6059,N_5966,N_5819);
nor U6060 (N_6060,N_5808,N_5991);
nand U6061 (N_6061,N_5872,N_5921);
xor U6062 (N_6062,N_5867,N_5853);
or U6063 (N_6063,N_5928,N_5923);
nor U6064 (N_6064,N_5836,N_5924);
and U6065 (N_6065,N_5783,N_5932);
xor U6066 (N_6066,N_5894,N_5856);
and U6067 (N_6067,N_5752,N_5854);
nand U6068 (N_6068,N_5927,N_5935);
or U6069 (N_6069,N_5849,N_5958);
nand U6070 (N_6070,N_5990,N_5879);
and U6071 (N_6071,N_5796,N_5761);
nand U6072 (N_6072,N_5910,N_5952);
xnor U6073 (N_6073,N_5770,N_5758);
nor U6074 (N_6074,N_5897,N_5951);
xnor U6075 (N_6075,N_5799,N_5967);
or U6076 (N_6076,N_5820,N_5917);
nand U6077 (N_6077,N_5964,N_5862);
nor U6078 (N_6078,N_5911,N_5974);
xor U6079 (N_6079,N_5757,N_5888);
xnor U6080 (N_6080,N_5777,N_5988);
xnor U6081 (N_6081,N_5810,N_5839);
nor U6082 (N_6082,N_5806,N_5857);
nor U6083 (N_6083,N_5866,N_5787);
xor U6084 (N_6084,N_5805,N_5771);
nand U6085 (N_6085,N_5956,N_5763);
and U6086 (N_6086,N_5984,N_5786);
nand U6087 (N_6087,N_5993,N_5885);
or U6088 (N_6088,N_5755,N_5969);
nor U6089 (N_6089,N_5995,N_5825);
nand U6090 (N_6090,N_5915,N_5794);
or U6091 (N_6091,N_5998,N_5772);
nor U6092 (N_6092,N_5768,N_5968);
nand U6093 (N_6093,N_5954,N_5914);
nand U6094 (N_6094,N_5904,N_5931);
and U6095 (N_6095,N_5774,N_5802);
or U6096 (N_6096,N_5756,N_5937);
nor U6097 (N_6097,N_5809,N_5987);
and U6098 (N_6098,N_5948,N_5902);
nor U6099 (N_6099,N_5882,N_5815);
nand U6100 (N_6100,N_5831,N_5961);
xor U6101 (N_6101,N_5795,N_5999);
nor U6102 (N_6102,N_5833,N_5788);
xnor U6103 (N_6103,N_5822,N_5994);
xor U6104 (N_6104,N_5837,N_5959);
nor U6105 (N_6105,N_5940,N_5811);
and U6106 (N_6106,N_5913,N_5992);
nand U6107 (N_6107,N_5946,N_5843);
nand U6108 (N_6108,N_5981,N_5792);
or U6109 (N_6109,N_5842,N_5850);
nor U6110 (N_6110,N_5938,N_5900);
xor U6111 (N_6111,N_5907,N_5803);
nand U6112 (N_6112,N_5939,N_5919);
or U6113 (N_6113,N_5875,N_5903);
or U6114 (N_6114,N_5751,N_5896);
xnor U6115 (N_6115,N_5982,N_5916);
xnor U6116 (N_6116,N_5804,N_5955);
and U6117 (N_6117,N_5812,N_5766);
xnor U6118 (N_6118,N_5765,N_5863);
nor U6119 (N_6119,N_5814,N_5864);
and U6120 (N_6120,N_5985,N_5762);
and U6121 (N_6121,N_5891,N_5813);
or U6122 (N_6122,N_5883,N_5881);
xor U6123 (N_6123,N_5767,N_5934);
nor U6124 (N_6124,N_5942,N_5860);
and U6125 (N_6125,N_5980,N_5905);
xor U6126 (N_6126,N_5771,N_5945);
nand U6127 (N_6127,N_5855,N_5850);
nand U6128 (N_6128,N_5840,N_5778);
nand U6129 (N_6129,N_5928,N_5906);
nor U6130 (N_6130,N_5968,N_5892);
or U6131 (N_6131,N_5882,N_5923);
xor U6132 (N_6132,N_5987,N_5879);
nand U6133 (N_6133,N_5765,N_5903);
and U6134 (N_6134,N_5789,N_5903);
or U6135 (N_6135,N_5969,N_5914);
nand U6136 (N_6136,N_5845,N_5919);
nor U6137 (N_6137,N_5977,N_5877);
nor U6138 (N_6138,N_5909,N_5937);
or U6139 (N_6139,N_5792,N_5797);
nor U6140 (N_6140,N_5806,N_5784);
xnor U6141 (N_6141,N_5864,N_5978);
and U6142 (N_6142,N_5903,N_5785);
nor U6143 (N_6143,N_5868,N_5835);
nand U6144 (N_6144,N_5920,N_5977);
xor U6145 (N_6145,N_5910,N_5834);
nand U6146 (N_6146,N_5927,N_5877);
nand U6147 (N_6147,N_5911,N_5788);
nor U6148 (N_6148,N_5883,N_5943);
nand U6149 (N_6149,N_5832,N_5986);
and U6150 (N_6150,N_5837,N_5897);
nor U6151 (N_6151,N_5789,N_5892);
and U6152 (N_6152,N_5836,N_5820);
or U6153 (N_6153,N_5966,N_5826);
and U6154 (N_6154,N_5799,N_5985);
and U6155 (N_6155,N_5762,N_5913);
and U6156 (N_6156,N_5920,N_5911);
nand U6157 (N_6157,N_5753,N_5948);
xnor U6158 (N_6158,N_5862,N_5914);
nand U6159 (N_6159,N_5760,N_5820);
or U6160 (N_6160,N_5824,N_5778);
and U6161 (N_6161,N_5831,N_5839);
nand U6162 (N_6162,N_5913,N_5845);
nor U6163 (N_6163,N_5775,N_5804);
and U6164 (N_6164,N_5774,N_5922);
or U6165 (N_6165,N_5952,N_5828);
nand U6166 (N_6166,N_5763,N_5845);
nand U6167 (N_6167,N_5987,N_5786);
nand U6168 (N_6168,N_5760,N_5801);
nor U6169 (N_6169,N_5975,N_5866);
and U6170 (N_6170,N_5784,N_5872);
xnor U6171 (N_6171,N_5879,N_5873);
xnor U6172 (N_6172,N_5886,N_5892);
nor U6173 (N_6173,N_5760,N_5880);
nor U6174 (N_6174,N_5936,N_5869);
nor U6175 (N_6175,N_5752,N_5918);
xor U6176 (N_6176,N_5862,N_5974);
or U6177 (N_6177,N_5867,N_5864);
and U6178 (N_6178,N_5926,N_5877);
or U6179 (N_6179,N_5925,N_5798);
and U6180 (N_6180,N_5864,N_5905);
or U6181 (N_6181,N_5921,N_5933);
and U6182 (N_6182,N_5795,N_5982);
and U6183 (N_6183,N_5985,N_5910);
nand U6184 (N_6184,N_5873,N_5802);
and U6185 (N_6185,N_5866,N_5924);
or U6186 (N_6186,N_5779,N_5995);
and U6187 (N_6187,N_5863,N_5869);
and U6188 (N_6188,N_5798,N_5957);
xor U6189 (N_6189,N_5966,N_5992);
or U6190 (N_6190,N_5755,N_5766);
nor U6191 (N_6191,N_5878,N_5788);
nor U6192 (N_6192,N_5764,N_5812);
xnor U6193 (N_6193,N_5868,N_5895);
and U6194 (N_6194,N_5993,N_5948);
xnor U6195 (N_6195,N_5877,N_5970);
and U6196 (N_6196,N_5936,N_5854);
or U6197 (N_6197,N_5874,N_5957);
or U6198 (N_6198,N_5924,N_5775);
or U6199 (N_6199,N_5831,N_5808);
and U6200 (N_6200,N_5756,N_5890);
xor U6201 (N_6201,N_5931,N_5851);
nor U6202 (N_6202,N_5991,N_5823);
xnor U6203 (N_6203,N_5950,N_5981);
nand U6204 (N_6204,N_5814,N_5972);
nand U6205 (N_6205,N_5904,N_5778);
nor U6206 (N_6206,N_5944,N_5817);
xor U6207 (N_6207,N_5958,N_5793);
nand U6208 (N_6208,N_5824,N_5794);
xnor U6209 (N_6209,N_5992,N_5858);
xnor U6210 (N_6210,N_5849,N_5927);
or U6211 (N_6211,N_5894,N_5817);
xor U6212 (N_6212,N_5768,N_5830);
and U6213 (N_6213,N_5935,N_5798);
xor U6214 (N_6214,N_5859,N_5793);
or U6215 (N_6215,N_5967,N_5764);
and U6216 (N_6216,N_5949,N_5767);
nand U6217 (N_6217,N_5774,N_5825);
xnor U6218 (N_6218,N_5918,N_5848);
xor U6219 (N_6219,N_5843,N_5838);
xor U6220 (N_6220,N_5832,N_5979);
nor U6221 (N_6221,N_5829,N_5955);
and U6222 (N_6222,N_5942,N_5791);
xor U6223 (N_6223,N_5798,N_5963);
nand U6224 (N_6224,N_5763,N_5870);
or U6225 (N_6225,N_5812,N_5753);
or U6226 (N_6226,N_5773,N_5942);
xor U6227 (N_6227,N_5955,N_5757);
nand U6228 (N_6228,N_5969,N_5908);
xnor U6229 (N_6229,N_5863,N_5888);
nor U6230 (N_6230,N_5879,N_5889);
nand U6231 (N_6231,N_5978,N_5902);
or U6232 (N_6232,N_5755,N_5837);
xnor U6233 (N_6233,N_5966,N_5874);
nand U6234 (N_6234,N_5915,N_5897);
or U6235 (N_6235,N_5782,N_5886);
nor U6236 (N_6236,N_5766,N_5780);
nor U6237 (N_6237,N_5938,N_5912);
nand U6238 (N_6238,N_5788,N_5829);
nand U6239 (N_6239,N_5812,N_5980);
nor U6240 (N_6240,N_5810,N_5765);
nand U6241 (N_6241,N_5760,N_5895);
and U6242 (N_6242,N_5865,N_5956);
nor U6243 (N_6243,N_5861,N_5935);
and U6244 (N_6244,N_5819,N_5812);
xnor U6245 (N_6245,N_5762,N_5798);
nand U6246 (N_6246,N_5997,N_5872);
nor U6247 (N_6247,N_5904,N_5888);
or U6248 (N_6248,N_5756,N_5935);
and U6249 (N_6249,N_5825,N_5978);
nand U6250 (N_6250,N_6132,N_6169);
or U6251 (N_6251,N_6141,N_6220);
xor U6252 (N_6252,N_6113,N_6033);
nor U6253 (N_6253,N_6210,N_6093);
or U6254 (N_6254,N_6233,N_6140);
nor U6255 (N_6255,N_6034,N_6230);
or U6256 (N_6256,N_6173,N_6245);
or U6257 (N_6257,N_6189,N_6242);
nand U6258 (N_6258,N_6087,N_6082);
or U6259 (N_6259,N_6192,N_6160);
or U6260 (N_6260,N_6066,N_6117);
xor U6261 (N_6261,N_6244,N_6213);
nor U6262 (N_6262,N_6020,N_6203);
nand U6263 (N_6263,N_6126,N_6199);
nor U6264 (N_6264,N_6143,N_6144);
xor U6265 (N_6265,N_6238,N_6237);
and U6266 (N_6266,N_6156,N_6080);
xnor U6267 (N_6267,N_6150,N_6016);
xor U6268 (N_6268,N_6154,N_6130);
xor U6269 (N_6269,N_6198,N_6178);
nor U6270 (N_6270,N_6099,N_6114);
nor U6271 (N_6271,N_6124,N_6094);
nor U6272 (N_6272,N_6201,N_6078);
xor U6273 (N_6273,N_6157,N_6159);
nand U6274 (N_6274,N_6176,N_6004);
nand U6275 (N_6275,N_6221,N_6069);
nor U6276 (N_6276,N_6215,N_6030);
nand U6277 (N_6277,N_6088,N_6089);
nand U6278 (N_6278,N_6142,N_6064);
xnor U6279 (N_6279,N_6101,N_6223);
and U6280 (N_6280,N_6059,N_6038);
nor U6281 (N_6281,N_6183,N_6228);
xor U6282 (N_6282,N_6180,N_6118);
nand U6283 (N_6283,N_6047,N_6191);
and U6284 (N_6284,N_6218,N_6027);
nand U6285 (N_6285,N_6205,N_6096);
xnor U6286 (N_6286,N_6010,N_6011);
xnor U6287 (N_6287,N_6207,N_6107);
xnor U6288 (N_6288,N_6163,N_6013);
and U6289 (N_6289,N_6104,N_6017);
or U6290 (N_6290,N_6060,N_6138);
xnor U6291 (N_6291,N_6184,N_6023);
or U6292 (N_6292,N_6090,N_6200);
and U6293 (N_6293,N_6211,N_6097);
or U6294 (N_6294,N_6236,N_6056);
and U6295 (N_6295,N_6036,N_6052);
nor U6296 (N_6296,N_6042,N_6084);
xor U6297 (N_6297,N_6147,N_6021);
nand U6298 (N_6298,N_6098,N_6070);
or U6299 (N_6299,N_6015,N_6081);
or U6300 (N_6300,N_6162,N_6137);
and U6301 (N_6301,N_6077,N_6185);
or U6302 (N_6302,N_6106,N_6136);
or U6303 (N_6303,N_6134,N_6073);
or U6304 (N_6304,N_6045,N_6240);
nand U6305 (N_6305,N_6234,N_6014);
or U6306 (N_6306,N_6125,N_6071);
nand U6307 (N_6307,N_6048,N_6123);
or U6308 (N_6308,N_6241,N_6131);
or U6309 (N_6309,N_6041,N_6006);
nor U6310 (N_6310,N_6044,N_6243);
and U6311 (N_6311,N_6146,N_6002);
xnor U6312 (N_6312,N_6012,N_6110);
and U6313 (N_6313,N_6095,N_6005);
xnor U6314 (N_6314,N_6151,N_6153);
or U6315 (N_6315,N_6170,N_6072);
nand U6316 (N_6316,N_6206,N_6092);
nand U6317 (N_6317,N_6196,N_6067);
xor U6318 (N_6318,N_6083,N_6202);
or U6319 (N_6319,N_6039,N_6239);
nor U6320 (N_6320,N_6164,N_6024);
nand U6321 (N_6321,N_6018,N_6128);
nand U6322 (N_6322,N_6171,N_6108);
and U6323 (N_6323,N_6186,N_6148);
nand U6324 (N_6324,N_6166,N_6219);
or U6325 (N_6325,N_6122,N_6001);
or U6326 (N_6326,N_6031,N_6019);
or U6327 (N_6327,N_6195,N_6079);
or U6328 (N_6328,N_6226,N_6103);
nor U6329 (N_6329,N_6187,N_6248);
nand U6330 (N_6330,N_6247,N_6100);
nor U6331 (N_6331,N_6053,N_6172);
and U6332 (N_6332,N_6161,N_6050);
or U6333 (N_6333,N_6065,N_6058);
nor U6334 (N_6334,N_6111,N_6208);
nor U6335 (N_6335,N_6217,N_6158);
or U6336 (N_6336,N_6179,N_6209);
or U6337 (N_6337,N_6116,N_6076);
or U6338 (N_6338,N_6035,N_6091);
xor U6339 (N_6339,N_6229,N_6177);
or U6340 (N_6340,N_6249,N_6168);
nand U6341 (N_6341,N_6037,N_6175);
nor U6342 (N_6342,N_6102,N_6000);
xnor U6343 (N_6343,N_6212,N_6246);
or U6344 (N_6344,N_6190,N_6227);
nor U6345 (N_6345,N_6174,N_6121);
or U6346 (N_6346,N_6197,N_6231);
and U6347 (N_6347,N_6007,N_6167);
xor U6348 (N_6348,N_6105,N_6120);
xnor U6349 (N_6349,N_6222,N_6055);
xor U6350 (N_6350,N_6152,N_6155);
or U6351 (N_6351,N_6235,N_6182);
and U6352 (N_6352,N_6165,N_6149);
nor U6353 (N_6353,N_6086,N_6135);
xor U6354 (N_6354,N_6194,N_6028);
and U6355 (N_6355,N_6009,N_6188);
xor U6356 (N_6356,N_6181,N_6043);
nor U6357 (N_6357,N_6112,N_6216);
or U6358 (N_6358,N_6224,N_6204);
xor U6359 (N_6359,N_6061,N_6032);
nand U6360 (N_6360,N_6003,N_6029);
or U6361 (N_6361,N_6049,N_6225);
and U6362 (N_6362,N_6068,N_6046);
xor U6363 (N_6363,N_6115,N_6109);
nand U6364 (N_6364,N_6232,N_6075);
xor U6365 (N_6365,N_6008,N_6040);
or U6366 (N_6366,N_6129,N_6062);
xnor U6367 (N_6367,N_6133,N_6051);
nand U6368 (N_6368,N_6139,N_6022);
nand U6369 (N_6369,N_6025,N_6119);
xnor U6370 (N_6370,N_6026,N_6085);
and U6371 (N_6371,N_6145,N_6063);
xnor U6372 (N_6372,N_6057,N_6054);
nor U6373 (N_6373,N_6127,N_6214);
nor U6374 (N_6374,N_6074,N_6193);
or U6375 (N_6375,N_6186,N_6112);
xor U6376 (N_6376,N_6166,N_6173);
nor U6377 (N_6377,N_6074,N_6096);
or U6378 (N_6378,N_6181,N_6115);
and U6379 (N_6379,N_6085,N_6195);
and U6380 (N_6380,N_6153,N_6148);
xnor U6381 (N_6381,N_6007,N_6136);
or U6382 (N_6382,N_6007,N_6216);
xor U6383 (N_6383,N_6207,N_6069);
xnor U6384 (N_6384,N_6041,N_6049);
nor U6385 (N_6385,N_6145,N_6154);
xnor U6386 (N_6386,N_6124,N_6123);
or U6387 (N_6387,N_6063,N_6013);
nor U6388 (N_6388,N_6245,N_6231);
nand U6389 (N_6389,N_6224,N_6032);
and U6390 (N_6390,N_6056,N_6190);
or U6391 (N_6391,N_6035,N_6149);
xnor U6392 (N_6392,N_6225,N_6206);
or U6393 (N_6393,N_6188,N_6083);
nand U6394 (N_6394,N_6052,N_6147);
nand U6395 (N_6395,N_6176,N_6056);
nand U6396 (N_6396,N_6206,N_6023);
nand U6397 (N_6397,N_6135,N_6199);
nand U6398 (N_6398,N_6229,N_6081);
and U6399 (N_6399,N_6066,N_6108);
nor U6400 (N_6400,N_6106,N_6015);
nand U6401 (N_6401,N_6152,N_6056);
nor U6402 (N_6402,N_6077,N_6120);
nand U6403 (N_6403,N_6061,N_6002);
xnor U6404 (N_6404,N_6235,N_6140);
xor U6405 (N_6405,N_6044,N_6114);
nand U6406 (N_6406,N_6248,N_6019);
xor U6407 (N_6407,N_6135,N_6091);
nor U6408 (N_6408,N_6047,N_6236);
nor U6409 (N_6409,N_6190,N_6014);
nand U6410 (N_6410,N_6187,N_6092);
xor U6411 (N_6411,N_6093,N_6220);
or U6412 (N_6412,N_6191,N_6077);
nand U6413 (N_6413,N_6219,N_6188);
nand U6414 (N_6414,N_6175,N_6119);
or U6415 (N_6415,N_6089,N_6211);
xor U6416 (N_6416,N_6243,N_6056);
nand U6417 (N_6417,N_6230,N_6088);
nor U6418 (N_6418,N_6249,N_6237);
xor U6419 (N_6419,N_6182,N_6055);
and U6420 (N_6420,N_6217,N_6151);
nand U6421 (N_6421,N_6008,N_6135);
nor U6422 (N_6422,N_6059,N_6237);
and U6423 (N_6423,N_6228,N_6022);
and U6424 (N_6424,N_6075,N_6027);
and U6425 (N_6425,N_6033,N_6090);
or U6426 (N_6426,N_6182,N_6234);
and U6427 (N_6427,N_6133,N_6136);
and U6428 (N_6428,N_6007,N_6135);
and U6429 (N_6429,N_6050,N_6054);
nor U6430 (N_6430,N_6218,N_6215);
or U6431 (N_6431,N_6087,N_6073);
nand U6432 (N_6432,N_6033,N_6085);
or U6433 (N_6433,N_6000,N_6226);
nand U6434 (N_6434,N_6109,N_6175);
nand U6435 (N_6435,N_6024,N_6038);
nand U6436 (N_6436,N_6147,N_6120);
nor U6437 (N_6437,N_6049,N_6213);
nand U6438 (N_6438,N_6006,N_6204);
or U6439 (N_6439,N_6053,N_6086);
and U6440 (N_6440,N_6225,N_6035);
nor U6441 (N_6441,N_6105,N_6104);
or U6442 (N_6442,N_6029,N_6119);
and U6443 (N_6443,N_6070,N_6205);
and U6444 (N_6444,N_6065,N_6240);
nor U6445 (N_6445,N_6137,N_6017);
nand U6446 (N_6446,N_6174,N_6157);
nor U6447 (N_6447,N_6104,N_6060);
or U6448 (N_6448,N_6223,N_6229);
or U6449 (N_6449,N_6221,N_6194);
and U6450 (N_6450,N_6086,N_6163);
nor U6451 (N_6451,N_6079,N_6041);
and U6452 (N_6452,N_6187,N_6145);
xor U6453 (N_6453,N_6149,N_6243);
nor U6454 (N_6454,N_6088,N_6215);
and U6455 (N_6455,N_6124,N_6046);
nand U6456 (N_6456,N_6034,N_6025);
xnor U6457 (N_6457,N_6027,N_6158);
nor U6458 (N_6458,N_6058,N_6075);
nand U6459 (N_6459,N_6236,N_6096);
and U6460 (N_6460,N_6225,N_6123);
nand U6461 (N_6461,N_6243,N_6006);
or U6462 (N_6462,N_6209,N_6194);
or U6463 (N_6463,N_6010,N_6189);
and U6464 (N_6464,N_6248,N_6059);
nor U6465 (N_6465,N_6168,N_6009);
xnor U6466 (N_6466,N_6053,N_6227);
nor U6467 (N_6467,N_6194,N_6192);
nand U6468 (N_6468,N_6038,N_6055);
nand U6469 (N_6469,N_6237,N_6065);
nor U6470 (N_6470,N_6124,N_6154);
nand U6471 (N_6471,N_6067,N_6108);
or U6472 (N_6472,N_6248,N_6011);
nand U6473 (N_6473,N_6237,N_6221);
xnor U6474 (N_6474,N_6112,N_6172);
nand U6475 (N_6475,N_6128,N_6166);
nand U6476 (N_6476,N_6196,N_6177);
or U6477 (N_6477,N_6023,N_6059);
and U6478 (N_6478,N_6020,N_6180);
xnor U6479 (N_6479,N_6202,N_6012);
and U6480 (N_6480,N_6150,N_6010);
or U6481 (N_6481,N_6004,N_6239);
and U6482 (N_6482,N_6005,N_6093);
nor U6483 (N_6483,N_6127,N_6131);
or U6484 (N_6484,N_6108,N_6179);
nor U6485 (N_6485,N_6069,N_6097);
nand U6486 (N_6486,N_6046,N_6238);
nor U6487 (N_6487,N_6183,N_6087);
nand U6488 (N_6488,N_6174,N_6187);
nor U6489 (N_6489,N_6054,N_6023);
nand U6490 (N_6490,N_6077,N_6145);
nor U6491 (N_6491,N_6050,N_6073);
nand U6492 (N_6492,N_6212,N_6113);
or U6493 (N_6493,N_6046,N_6216);
xnor U6494 (N_6494,N_6249,N_6032);
xnor U6495 (N_6495,N_6248,N_6039);
nand U6496 (N_6496,N_6198,N_6121);
or U6497 (N_6497,N_6104,N_6209);
or U6498 (N_6498,N_6059,N_6131);
or U6499 (N_6499,N_6209,N_6204);
and U6500 (N_6500,N_6387,N_6453);
or U6501 (N_6501,N_6407,N_6308);
and U6502 (N_6502,N_6428,N_6339);
and U6503 (N_6503,N_6426,N_6286);
or U6504 (N_6504,N_6309,N_6476);
nand U6505 (N_6505,N_6266,N_6349);
nor U6506 (N_6506,N_6402,N_6258);
nor U6507 (N_6507,N_6285,N_6287);
nand U6508 (N_6508,N_6317,N_6382);
nor U6509 (N_6509,N_6434,N_6293);
xnor U6510 (N_6510,N_6283,N_6303);
or U6511 (N_6511,N_6272,N_6263);
or U6512 (N_6512,N_6424,N_6381);
nand U6513 (N_6513,N_6401,N_6416);
xor U6514 (N_6514,N_6444,N_6466);
xor U6515 (N_6515,N_6473,N_6371);
nand U6516 (N_6516,N_6415,N_6411);
and U6517 (N_6517,N_6331,N_6423);
or U6518 (N_6518,N_6327,N_6481);
nand U6519 (N_6519,N_6267,N_6374);
nor U6520 (N_6520,N_6467,N_6408);
nand U6521 (N_6521,N_6457,N_6398);
and U6522 (N_6522,N_6346,N_6383);
nand U6523 (N_6523,N_6372,N_6456);
xor U6524 (N_6524,N_6284,N_6274);
nand U6525 (N_6525,N_6412,N_6436);
nand U6526 (N_6526,N_6449,N_6482);
nor U6527 (N_6527,N_6432,N_6437);
xor U6528 (N_6528,N_6433,N_6280);
or U6529 (N_6529,N_6319,N_6363);
nand U6530 (N_6530,N_6450,N_6356);
nor U6531 (N_6531,N_6307,N_6311);
and U6532 (N_6532,N_6262,N_6257);
xor U6533 (N_6533,N_6275,N_6276);
nand U6534 (N_6534,N_6343,N_6323);
nand U6535 (N_6535,N_6312,N_6400);
or U6536 (N_6536,N_6337,N_6299);
or U6537 (N_6537,N_6345,N_6338);
and U6538 (N_6538,N_6479,N_6393);
xor U6539 (N_6539,N_6461,N_6290);
nand U6540 (N_6540,N_6314,N_6354);
and U6541 (N_6541,N_6471,N_6347);
or U6542 (N_6542,N_6326,N_6348);
or U6543 (N_6543,N_6336,N_6421);
xnor U6544 (N_6544,N_6252,N_6264);
xnor U6545 (N_6545,N_6364,N_6498);
xnor U6546 (N_6546,N_6333,N_6489);
and U6547 (N_6547,N_6413,N_6458);
or U6548 (N_6548,N_6459,N_6306);
and U6549 (N_6549,N_6296,N_6268);
nand U6550 (N_6550,N_6497,N_6386);
xnor U6551 (N_6551,N_6321,N_6366);
or U6552 (N_6552,N_6451,N_6391);
nor U6553 (N_6553,N_6344,N_6406);
nand U6554 (N_6554,N_6404,N_6465);
nand U6555 (N_6555,N_6472,N_6397);
nand U6556 (N_6556,N_6385,N_6279);
nor U6557 (N_6557,N_6439,N_6255);
and U6558 (N_6558,N_6419,N_6452);
or U6559 (N_6559,N_6379,N_6492);
nand U6560 (N_6560,N_6313,N_6484);
xor U6561 (N_6561,N_6496,N_6341);
or U6562 (N_6562,N_6475,N_6427);
xor U6563 (N_6563,N_6361,N_6487);
nand U6564 (N_6564,N_6414,N_6455);
or U6565 (N_6565,N_6445,N_6277);
nand U6566 (N_6566,N_6384,N_6295);
xor U6567 (N_6567,N_6294,N_6320);
xor U6568 (N_6568,N_6297,N_6259);
xnor U6569 (N_6569,N_6369,N_6420);
nand U6570 (N_6570,N_6352,N_6495);
xnor U6571 (N_6571,N_6447,N_6301);
and U6572 (N_6572,N_6380,N_6477);
and U6573 (N_6573,N_6330,N_6362);
nand U6574 (N_6574,N_6394,N_6329);
xnor U6575 (N_6575,N_6431,N_6494);
and U6576 (N_6576,N_6324,N_6360);
nor U6577 (N_6577,N_6340,N_6390);
nor U6578 (N_6578,N_6392,N_6388);
nand U6579 (N_6579,N_6334,N_6488);
nand U6580 (N_6580,N_6468,N_6464);
nand U6581 (N_6581,N_6469,N_6367);
or U6582 (N_6582,N_6395,N_6396);
or U6583 (N_6583,N_6425,N_6378);
and U6584 (N_6584,N_6357,N_6422);
nor U6585 (N_6585,N_6438,N_6460);
xnor U6586 (N_6586,N_6478,N_6288);
or U6587 (N_6587,N_6271,N_6376);
nand U6588 (N_6588,N_6250,N_6332);
xnor U6589 (N_6589,N_6305,N_6485);
nor U6590 (N_6590,N_6373,N_6322);
or U6591 (N_6591,N_6265,N_6298);
and U6592 (N_6592,N_6429,N_6273);
and U6593 (N_6593,N_6328,N_6463);
or U6594 (N_6594,N_6491,N_6375);
nor U6595 (N_6595,N_6399,N_6410);
and U6596 (N_6596,N_6454,N_6300);
nor U6597 (N_6597,N_6289,N_6358);
or U6598 (N_6598,N_6405,N_6417);
and U6599 (N_6599,N_6318,N_6409);
xnor U6600 (N_6600,N_6270,N_6278);
xnor U6601 (N_6601,N_6281,N_6370);
xnor U6602 (N_6602,N_6282,N_6315);
and U6603 (N_6603,N_6304,N_6474);
nor U6604 (N_6604,N_6483,N_6443);
xor U6605 (N_6605,N_6389,N_6325);
or U6606 (N_6606,N_6261,N_6440);
nor U6607 (N_6607,N_6442,N_6377);
or U6608 (N_6608,N_6441,N_6462);
nor U6609 (N_6609,N_6359,N_6269);
nand U6610 (N_6610,N_6490,N_6256);
or U6611 (N_6611,N_6253,N_6292);
nor U6612 (N_6612,N_6302,N_6430);
or U6613 (N_6613,N_6310,N_6486);
xnor U6614 (N_6614,N_6260,N_6418);
xor U6615 (N_6615,N_6470,N_6351);
nor U6616 (N_6616,N_6254,N_6480);
or U6617 (N_6617,N_6350,N_6316);
nand U6618 (N_6618,N_6291,N_6499);
nand U6619 (N_6619,N_6368,N_6448);
nor U6620 (N_6620,N_6335,N_6435);
xor U6621 (N_6621,N_6251,N_6353);
nor U6622 (N_6622,N_6446,N_6355);
and U6623 (N_6623,N_6403,N_6365);
or U6624 (N_6624,N_6342,N_6493);
xnor U6625 (N_6625,N_6450,N_6417);
nand U6626 (N_6626,N_6425,N_6400);
xnor U6627 (N_6627,N_6391,N_6445);
nor U6628 (N_6628,N_6404,N_6378);
nor U6629 (N_6629,N_6366,N_6309);
xnor U6630 (N_6630,N_6252,N_6278);
and U6631 (N_6631,N_6498,N_6383);
or U6632 (N_6632,N_6323,N_6288);
xor U6633 (N_6633,N_6270,N_6372);
xor U6634 (N_6634,N_6441,N_6392);
or U6635 (N_6635,N_6349,N_6252);
xnor U6636 (N_6636,N_6456,N_6367);
nor U6637 (N_6637,N_6362,N_6483);
or U6638 (N_6638,N_6365,N_6495);
xnor U6639 (N_6639,N_6295,N_6336);
nor U6640 (N_6640,N_6294,N_6307);
or U6641 (N_6641,N_6468,N_6354);
xnor U6642 (N_6642,N_6335,N_6485);
xor U6643 (N_6643,N_6436,N_6340);
nor U6644 (N_6644,N_6269,N_6354);
nor U6645 (N_6645,N_6365,N_6457);
or U6646 (N_6646,N_6333,N_6468);
and U6647 (N_6647,N_6270,N_6293);
or U6648 (N_6648,N_6290,N_6430);
xnor U6649 (N_6649,N_6389,N_6426);
and U6650 (N_6650,N_6274,N_6496);
nor U6651 (N_6651,N_6357,N_6277);
nor U6652 (N_6652,N_6299,N_6320);
xor U6653 (N_6653,N_6465,N_6436);
nor U6654 (N_6654,N_6498,N_6410);
nand U6655 (N_6655,N_6492,N_6281);
or U6656 (N_6656,N_6355,N_6272);
and U6657 (N_6657,N_6299,N_6463);
and U6658 (N_6658,N_6429,N_6409);
xor U6659 (N_6659,N_6295,N_6472);
nand U6660 (N_6660,N_6422,N_6445);
xnor U6661 (N_6661,N_6313,N_6464);
or U6662 (N_6662,N_6305,N_6357);
nor U6663 (N_6663,N_6276,N_6328);
nand U6664 (N_6664,N_6450,N_6324);
xor U6665 (N_6665,N_6316,N_6446);
nand U6666 (N_6666,N_6341,N_6276);
nand U6667 (N_6667,N_6399,N_6404);
nor U6668 (N_6668,N_6371,N_6287);
nand U6669 (N_6669,N_6361,N_6393);
and U6670 (N_6670,N_6303,N_6369);
xor U6671 (N_6671,N_6360,N_6290);
and U6672 (N_6672,N_6378,N_6319);
xor U6673 (N_6673,N_6260,N_6319);
and U6674 (N_6674,N_6479,N_6272);
or U6675 (N_6675,N_6289,N_6440);
and U6676 (N_6676,N_6404,N_6496);
and U6677 (N_6677,N_6430,N_6336);
or U6678 (N_6678,N_6394,N_6462);
nor U6679 (N_6679,N_6270,N_6331);
nand U6680 (N_6680,N_6429,N_6354);
or U6681 (N_6681,N_6415,N_6394);
and U6682 (N_6682,N_6310,N_6453);
xor U6683 (N_6683,N_6309,N_6426);
nor U6684 (N_6684,N_6332,N_6255);
xnor U6685 (N_6685,N_6412,N_6463);
and U6686 (N_6686,N_6381,N_6470);
nor U6687 (N_6687,N_6454,N_6405);
or U6688 (N_6688,N_6447,N_6375);
nand U6689 (N_6689,N_6270,N_6315);
or U6690 (N_6690,N_6384,N_6324);
or U6691 (N_6691,N_6274,N_6429);
or U6692 (N_6692,N_6278,N_6365);
nor U6693 (N_6693,N_6471,N_6452);
nor U6694 (N_6694,N_6494,N_6423);
or U6695 (N_6695,N_6268,N_6498);
nand U6696 (N_6696,N_6476,N_6379);
xor U6697 (N_6697,N_6464,N_6306);
nand U6698 (N_6698,N_6322,N_6419);
and U6699 (N_6699,N_6398,N_6484);
xnor U6700 (N_6700,N_6294,N_6438);
nor U6701 (N_6701,N_6403,N_6498);
nand U6702 (N_6702,N_6474,N_6344);
or U6703 (N_6703,N_6397,N_6375);
or U6704 (N_6704,N_6329,N_6272);
xnor U6705 (N_6705,N_6288,N_6379);
nor U6706 (N_6706,N_6433,N_6449);
nor U6707 (N_6707,N_6484,N_6478);
xnor U6708 (N_6708,N_6486,N_6326);
nand U6709 (N_6709,N_6324,N_6341);
or U6710 (N_6710,N_6486,N_6390);
or U6711 (N_6711,N_6425,N_6385);
nand U6712 (N_6712,N_6277,N_6250);
xnor U6713 (N_6713,N_6440,N_6385);
nand U6714 (N_6714,N_6290,N_6469);
nor U6715 (N_6715,N_6409,N_6368);
or U6716 (N_6716,N_6337,N_6375);
xor U6717 (N_6717,N_6253,N_6346);
nand U6718 (N_6718,N_6369,N_6399);
xnor U6719 (N_6719,N_6491,N_6442);
or U6720 (N_6720,N_6321,N_6446);
and U6721 (N_6721,N_6275,N_6498);
nor U6722 (N_6722,N_6320,N_6317);
nand U6723 (N_6723,N_6392,N_6283);
and U6724 (N_6724,N_6426,N_6436);
nor U6725 (N_6725,N_6338,N_6324);
and U6726 (N_6726,N_6426,N_6262);
nor U6727 (N_6727,N_6254,N_6402);
or U6728 (N_6728,N_6302,N_6329);
nor U6729 (N_6729,N_6360,N_6272);
nor U6730 (N_6730,N_6350,N_6335);
and U6731 (N_6731,N_6267,N_6446);
nand U6732 (N_6732,N_6450,N_6326);
nand U6733 (N_6733,N_6466,N_6310);
or U6734 (N_6734,N_6258,N_6446);
or U6735 (N_6735,N_6485,N_6353);
or U6736 (N_6736,N_6267,N_6432);
nor U6737 (N_6737,N_6424,N_6251);
and U6738 (N_6738,N_6311,N_6467);
nand U6739 (N_6739,N_6365,N_6332);
nor U6740 (N_6740,N_6492,N_6308);
and U6741 (N_6741,N_6466,N_6391);
xnor U6742 (N_6742,N_6407,N_6402);
nand U6743 (N_6743,N_6471,N_6437);
nand U6744 (N_6744,N_6494,N_6479);
xor U6745 (N_6745,N_6423,N_6354);
and U6746 (N_6746,N_6329,N_6369);
xnor U6747 (N_6747,N_6304,N_6398);
xnor U6748 (N_6748,N_6307,N_6356);
or U6749 (N_6749,N_6429,N_6276);
nor U6750 (N_6750,N_6638,N_6666);
or U6751 (N_6751,N_6624,N_6569);
xnor U6752 (N_6752,N_6529,N_6513);
and U6753 (N_6753,N_6640,N_6580);
xor U6754 (N_6754,N_6522,N_6507);
xor U6755 (N_6755,N_6504,N_6581);
xnor U6756 (N_6756,N_6706,N_6599);
nor U6757 (N_6757,N_6668,N_6744);
or U6758 (N_6758,N_6653,N_6607);
xor U6759 (N_6759,N_6722,N_6739);
nand U6760 (N_6760,N_6628,N_6589);
and U6761 (N_6761,N_6642,N_6691);
or U6762 (N_6762,N_6710,N_6736);
and U6763 (N_6763,N_6594,N_6585);
nor U6764 (N_6764,N_6728,N_6662);
nand U6765 (N_6765,N_6692,N_6541);
and U6766 (N_6766,N_6561,N_6696);
nor U6767 (N_6767,N_6742,N_6530);
xnor U6768 (N_6768,N_6588,N_6553);
and U6769 (N_6769,N_6574,N_6697);
or U6770 (N_6770,N_6512,N_6577);
nor U6771 (N_6771,N_6702,N_6715);
and U6772 (N_6772,N_6674,N_6737);
and U6773 (N_6773,N_6731,N_6546);
xor U6774 (N_6774,N_6559,N_6694);
nor U6775 (N_6775,N_6595,N_6545);
and U6776 (N_6776,N_6667,N_6564);
or U6777 (N_6777,N_6604,N_6709);
nor U6778 (N_6778,N_6665,N_6724);
xor U6779 (N_6779,N_6505,N_6535);
nand U6780 (N_6780,N_6705,N_6718);
nand U6781 (N_6781,N_6747,N_6575);
and U6782 (N_6782,N_6528,N_6536);
xnor U6783 (N_6783,N_6621,N_6679);
nor U6784 (N_6784,N_6717,N_6684);
xor U6785 (N_6785,N_6551,N_6556);
nand U6786 (N_6786,N_6740,N_6741);
xor U6787 (N_6787,N_6675,N_6548);
or U6788 (N_6788,N_6681,N_6669);
or U6789 (N_6789,N_6590,N_6544);
nand U6790 (N_6790,N_6622,N_6605);
xnor U6791 (N_6791,N_6656,N_6555);
or U6792 (N_6792,N_6519,N_6620);
or U6793 (N_6793,N_6576,N_6664);
nor U6794 (N_6794,N_6516,N_6699);
or U6795 (N_6795,N_6734,N_6560);
nor U6796 (N_6796,N_6749,N_6523);
and U6797 (N_6797,N_6501,N_6597);
xor U6798 (N_6798,N_6524,N_6641);
and U6799 (N_6799,N_6554,N_6713);
xor U6800 (N_6800,N_6704,N_6693);
nor U6801 (N_6801,N_6543,N_6683);
and U6802 (N_6802,N_6626,N_6707);
nor U6803 (N_6803,N_6647,N_6526);
xor U6804 (N_6804,N_6745,N_6644);
xor U6805 (N_6805,N_6629,N_6730);
or U6806 (N_6806,N_6592,N_6733);
or U6807 (N_6807,N_6708,N_6547);
nand U6808 (N_6808,N_6518,N_6578);
xnor U6809 (N_6809,N_6601,N_6610);
or U6810 (N_6810,N_6630,N_6502);
and U6811 (N_6811,N_6615,N_6623);
and U6812 (N_6812,N_6506,N_6671);
xnor U6813 (N_6813,N_6635,N_6698);
xor U6814 (N_6814,N_6567,N_6658);
and U6815 (N_6815,N_6582,N_6688);
nand U6816 (N_6816,N_6539,N_6652);
or U6817 (N_6817,N_6570,N_6533);
or U6818 (N_6818,N_6631,N_6643);
xnor U6819 (N_6819,N_6525,N_6746);
xnor U6820 (N_6820,N_6735,N_6657);
or U6821 (N_6821,N_6617,N_6720);
nor U6822 (N_6822,N_6682,N_6534);
or U6823 (N_6823,N_6686,N_6609);
nor U6824 (N_6824,N_6579,N_6723);
nor U6825 (N_6825,N_6727,N_6510);
xnor U6826 (N_6826,N_6711,N_6689);
xnor U6827 (N_6827,N_6616,N_6673);
xor U6828 (N_6828,N_6532,N_6612);
or U6829 (N_6829,N_6562,N_6508);
xnor U6830 (N_6830,N_6586,N_6583);
xor U6831 (N_6831,N_6695,N_6558);
nor U6832 (N_6832,N_6654,N_6587);
nand U6833 (N_6833,N_6650,N_6625);
and U6834 (N_6834,N_6627,N_6633);
xor U6835 (N_6835,N_6677,N_6568);
and U6836 (N_6836,N_6634,N_6619);
or U6837 (N_6837,N_6596,N_6703);
xnor U6838 (N_6838,N_6690,N_6611);
nor U6839 (N_6839,N_6712,N_6542);
or U6840 (N_6840,N_6632,N_6738);
or U6841 (N_6841,N_6655,N_6670);
and U6842 (N_6842,N_6593,N_6520);
xor U6843 (N_6843,N_6608,N_6637);
and U6844 (N_6844,N_6552,N_6663);
nor U6845 (N_6845,N_6613,N_6729);
xor U6846 (N_6846,N_6719,N_6748);
xor U6847 (N_6847,N_6639,N_6531);
nand U6848 (N_6848,N_6700,N_6661);
or U6849 (N_6849,N_6680,N_6509);
nor U6850 (N_6850,N_6726,N_6687);
nor U6851 (N_6851,N_6618,N_6725);
nand U6852 (N_6852,N_6565,N_6573);
or U6853 (N_6853,N_6571,N_6716);
and U6854 (N_6854,N_6598,N_6743);
and U6855 (N_6855,N_6514,N_6646);
nor U6856 (N_6856,N_6721,N_6549);
xnor U6857 (N_6857,N_6500,N_6659);
nor U6858 (N_6858,N_6649,N_6732);
xor U6859 (N_6859,N_6563,N_6511);
xor U6860 (N_6860,N_6550,N_6645);
nor U6861 (N_6861,N_6685,N_6660);
nor U6862 (N_6862,N_6606,N_6527);
xor U6863 (N_6863,N_6603,N_6600);
or U6864 (N_6864,N_6572,N_6591);
xor U6865 (N_6865,N_6517,N_6701);
xor U6866 (N_6866,N_6503,N_6614);
nand U6867 (N_6867,N_6678,N_6540);
or U6868 (N_6868,N_6515,N_6566);
and U6869 (N_6869,N_6651,N_6648);
and U6870 (N_6870,N_6584,N_6537);
nor U6871 (N_6871,N_6557,N_6672);
nor U6872 (N_6872,N_6636,N_6538);
or U6873 (N_6873,N_6714,N_6602);
nand U6874 (N_6874,N_6521,N_6676);
and U6875 (N_6875,N_6577,N_6709);
xor U6876 (N_6876,N_6697,N_6526);
and U6877 (N_6877,N_6633,N_6741);
nor U6878 (N_6878,N_6689,N_6588);
xor U6879 (N_6879,N_6542,N_6657);
nor U6880 (N_6880,N_6701,N_6602);
and U6881 (N_6881,N_6615,N_6687);
xor U6882 (N_6882,N_6566,N_6705);
or U6883 (N_6883,N_6519,N_6548);
xor U6884 (N_6884,N_6567,N_6598);
or U6885 (N_6885,N_6584,N_6721);
and U6886 (N_6886,N_6546,N_6653);
and U6887 (N_6887,N_6739,N_6703);
xor U6888 (N_6888,N_6549,N_6543);
xnor U6889 (N_6889,N_6600,N_6661);
nor U6890 (N_6890,N_6598,N_6724);
nand U6891 (N_6891,N_6651,N_6749);
nor U6892 (N_6892,N_6581,N_6595);
xor U6893 (N_6893,N_6502,N_6661);
nand U6894 (N_6894,N_6663,N_6719);
or U6895 (N_6895,N_6501,N_6611);
nor U6896 (N_6896,N_6684,N_6588);
and U6897 (N_6897,N_6704,N_6660);
or U6898 (N_6898,N_6569,N_6697);
and U6899 (N_6899,N_6653,N_6692);
or U6900 (N_6900,N_6572,N_6716);
nor U6901 (N_6901,N_6747,N_6566);
xor U6902 (N_6902,N_6606,N_6727);
or U6903 (N_6903,N_6747,N_6548);
or U6904 (N_6904,N_6745,N_6668);
nor U6905 (N_6905,N_6537,N_6639);
nor U6906 (N_6906,N_6563,N_6699);
nand U6907 (N_6907,N_6533,N_6736);
xor U6908 (N_6908,N_6710,N_6553);
nor U6909 (N_6909,N_6583,N_6730);
nor U6910 (N_6910,N_6506,N_6514);
and U6911 (N_6911,N_6517,N_6573);
xnor U6912 (N_6912,N_6671,N_6630);
nor U6913 (N_6913,N_6678,N_6677);
nand U6914 (N_6914,N_6637,N_6631);
or U6915 (N_6915,N_6676,N_6612);
xor U6916 (N_6916,N_6652,N_6577);
xnor U6917 (N_6917,N_6654,N_6670);
xor U6918 (N_6918,N_6691,N_6509);
nor U6919 (N_6919,N_6593,N_6542);
and U6920 (N_6920,N_6652,N_6542);
nor U6921 (N_6921,N_6534,N_6702);
xnor U6922 (N_6922,N_6687,N_6538);
xnor U6923 (N_6923,N_6651,N_6644);
xnor U6924 (N_6924,N_6509,N_6592);
or U6925 (N_6925,N_6616,N_6665);
nor U6926 (N_6926,N_6731,N_6527);
nor U6927 (N_6927,N_6628,N_6564);
xor U6928 (N_6928,N_6739,N_6533);
nor U6929 (N_6929,N_6627,N_6648);
and U6930 (N_6930,N_6603,N_6573);
or U6931 (N_6931,N_6638,N_6687);
and U6932 (N_6932,N_6638,N_6678);
xnor U6933 (N_6933,N_6645,N_6731);
or U6934 (N_6934,N_6617,N_6537);
xnor U6935 (N_6935,N_6635,N_6614);
nor U6936 (N_6936,N_6724,N_6600);
and U6937 (N_6937,N_6691,N_6625);
xnor U6938 (N_6938,N_6503,N_6723);
xor U6939 (N_6939,N_6702,N_6725);
nor U6940 (N_6940,N_6619,N_6673);
or U6941 (N_6941,N_6749,N_6542);
and U6942 (N_6942,N_6611,N_6658);
and U6943 (N_6943,N_6646,N_6531);
xnor U6944 (N_6944,N_6733,N_6628);
nand U6945 (N_6945,N_6568,N_6613);
and U6946 (N_6946,N_6718,N_6559);
and U6947 (N_6947,N_6597,N_6677);
and U6948 (N_6948,N_6722,N_6665);
nand U6949 (N_6949,N_6673,N_6708);
and U6950 (N_6950,N_6559,N_6721);
xor U6951 (N_6951,N_6515,N_6748);
nand U6952 (N_6952,N_6650,N_6594);
nand U6953 (N_6953,N_6719,N_6689);
and U6954 (N_6954,N_6659,N_6749);
nand U6955 (N_6955,N_6623,N_6719);
xnor U6956 (N_6956,N_6588,N_6565);
or U6957 (N_6957,N_6696,N_6533);
xnor U6958 (N_6958,N_6650,N_6633);
and U6959 (N_6959,N_6503,N_6591);
nor U6960 (N_6960,N_6687,N_6525);
nand U6961 (N_6961,N_6585,N_6662);
nor U6962 (N_6962,N_6601,N_6705);
xor U6963 (N_6963,N_6595,N_6541);
nor U6964 (N_6964,N_6688,N_6731);
nand U6965 (N_6965,N_6585,N_6660);
or U6966 (N_6966,N_6612,N_6645);
or U6967 (N_6967,N_6571,N_6742);
or U6968 (N_6968,N_6724,N_6648);
nand U6969 (N_6969,N_6702,N_6517);
and U6970 (N_6970,N_6722,N_6602);
xnor U6971 (N_6971,N_6672,N_6713);
xor U6972 (N_6972,N_6665,N_6537);
nor U6973 (N_6973,N_6632,N_6697);
xor U6974 (N_6974,N_6505,N_6536);
or U6975 (N_6975,N_6517,N_6681);
xor U6976 (N_6976,N_6707,N_6570);
or U6977 (N_6977,N_6620,N_6647);
nand U6978 (N_6978,N_6508,N_6612);
nor U6979 (N_6979,N_6601,N_6712);
nor U6980 (N_6980,N_6582,N_6699);
xnor U6981 (N_6981,N_6541,N_6699);
nor U6982 (N_6982,N_6748,N_6632);
nor U6983 (N_6983,N_6519,N_6621);
nand U6984 (N_6984,N_6518,N_6638);
nand U6985 (N_6985,N_6554,N_6502);
nor U6986 (N_6986,N_6704,N_6574);
nand U6987 (N_6987,N_6548,N_6595);
or U6988 (N_6988,N_6595,N_6621);
nand U6989 (N_6989,N_6745,N_6734);
xnor U6990 (N_6990,N_6698,N_6553);
or U6991 (N_6991,N_6556,N_6533);
nand U6992 (N_6992,N_6514,N_6591);
nand U6993 (N_6993,N_6638,N_6684);
nand U6994 (N_6994,N_6612,N_6540);
nor U6995 (N_6995,N_6506,N_6596);
or U6996 (N_6996,N_6569,N_6629);
and U6997 (N_6997,N_6534,N_6735);
nand U6998 (N_6998,N_6635,N_6733);
nor U6999 (N_6999,N_6679,N_6513);
or U7000 (N_7000,N_6795,N_6981);
nor U7001 (N_7001,N_6871,N_6986);
nand U7002 (N_7002,N_6844,N_6923);
nor U7003 (N_7003,N_6814,N_6967);
and U7004 (N_7004,N_6954,N_6810);
xor U7005 (N_7005,N_6957,N_6983);
or U7006 (N_7006,N_6935,N_6834);
xor U7007 (N_7007,N_6945,N_6947);
nor U7008 (N_7008,N_6802,N_6968);
xnor U7009 (N_7009,N_6752,N_6888);
nand U7010 (N_7010,N_6780,N_6946);
and U7011 (N_7011,N_6851,N_6782);
nand U7012 (N_7012,N_6926,N_6969);
nand U7013 (N_7013,N_6950,N_6924);
xor U7014 (N_7014,N_6987,N_6766);
xnor U7015 (N_7015,N_6966,N_6833);
or U7016 (N_7016,N_6750,N_6886);
xnor U7017 (N_7017,N_6789,N_6919);
xor U7018 (N_7018,N_6872,N_6955);
and U7019 (N_7019,N_6857,N_6865);
and U7020 (N_7020,N_6774,N_6912);
and U7021 (N_7021,N_6881,N_6991);
nor U7022 (N_7022,N_6993,N_6849);
and U7023 (N_7023,N_6831,N_6760);
nor U7024 (N_7024,N_6917,N_6862);
nand U7025 (N_7025,N_6835,N_6895);
nand U7026 (N_7026,N_6822,N_6842);
or U7027 (N_7027,N_6816,N_6909);
xor U7028 (N_7028,N_6798,N_6885);
xnor U7029 (N_7029,N_6804,N_6762);
and U7030 (N_7030,N_6818,N_6904);
xnor U7031 (N_7031,N_6972,N_6860);
nor U7032 (N_7032,N_6803,N_6942);
nand U7033 (N_7033,N_6850,N_6910);
xor U7034 (N_7034,N_6847,N_6866);
nand U7035 (N_7035,N_6769,N_6894);
nor U7036 (N_7036,N_6922,N_6824);
and U7037 (N_7037,N_6876,N_6979);
and U7038 (N_7038,N_6773,N_6751);
or U7039 (N_7039,N_6775,N_6870);
nand U7040 (N_7040,N_6905,N_6877);
nor U7041 (N_7041,N_6827,N_6953);
and U7042 (N_7042,N_6845,N_6920);
xor U7043 (N_7043,N_6765,N_6777);
xor U7044 (N_7044,N_6826,N_6973);
nand U7045 (N_7045,N_6755,N_6929);
nor U7046 (N_7046,N_6989,N_6927);
nor U7047 (N_7047,N_6875,N_6999);
xnor U7048 (N_7048,N_6813,N_6829);
nand U7049 (N_7049,N_6936,N_6965);
xnor U7050 (N_7050,N_6868,N_6990);
nand U7051 (N_7051,N_6943,N_6776);
xnor U7052 (N_7052,N_6930,N_6960);
and U7053 (N_7053,N_6959,N_6889);
and U7054 (N_7054,N_6772,N_6840);
and U7055 (N_7055,N_6825,N_6938);
nor U7056 (N_7056,N_6839,N_6820);
or U7057 (N_7057,N_6792,N_6884);
or U7058 (N_7058,N_6819,N_6757);
or U7059 (N_7059,N_6956,N_6996);
nand U7060 (N_7060,N_6784,N_6809);
nor U7061 (N_7061,N_6997,N_6754);
nor U7062 (N_7062,N_6763,N_6913);
nor U7063 (N_7063,N_6908,N_6984);
nand U7064 (N_7064,N_6882,N_6998);
nand U7065 (N_7065,N_6787,N_6994);
nand U7066 (N_7066,N_6793,N_6800);
nor U7067 (N_7067,N_6974,N_6873);
or U7068 (N_7068,N_6932,N_6828);
or U7069 (N_7069,N_6768,N_6977);
nor U7070 (N_7070,N_6867,N_6846);
nand U7071 (N_7071,N_6783,N_6896);
nor U7072 (N_7072,N_6964,N_6911);
and U7073 (N_7073,N_6864,N_6801);
nand U7074 (N_7074,N_6985,N_6958);
and U7075 (N_7075,N_6883,N_6797);
xor U7076 (N_7076,N_6916,N_6806);
nor U7077 (N_7077,N_6940,N_6962);
nor U7078 (N_7078,N_6856,N_6941);
and U7079 (N_7079,N_6821,N_6812);
nand U7080 (N_7080,N_6805,N_6855);
and U7081 (N_7081,N_6925,N_6971);
nor U7082 (N_7082,N_6837,N_6900);
or U7083 (N_7083,N_6907,N_6970);
xor U7084 (N_7084,N_6758,N_6817);
nand U7085 (N_7085,N_6949,N_6933);
nand U7086 (N_7086,N_6854,N_6879);
and U7087 (N_7087,N_6790,N_6753);
xnor U7088 (N_7088,N_6788,N_6902);
and U7089 (N_7089,N_6939,N_6952);
or U7090 (N_7090,N_6975,N_6890);
or U7091 (N_7091,N_6869,N_6963);
nand U7092 (N_7092,N_6841,N_6898);
nand U7093 (N_7093,N_6764,N_6811);
or U7094 (N_7094,N_6861,N_6799);
nand U7095 (N_7095,N_6761,N_6948);
nor U7096 (N_7096,N_6901,N_6830);
nor U7097 (N_7097,N_6770,N_6899);
xor U7098 (N_7098,N_6903,N_6931);
or U7099 (N_7099,N_6836,N_6921);
or U7100 (N_7100,N_6944,N_6992);
nor U7101 (N_7101,N_6778,N_6978);
xnor U7102 (N_7102,N_6848,N_6756);
and U7103 (N_7103,N_6863,N_6893);
nand U7104 (N_7104,N_6980,N_6823);
xnor U7105 (N_7105,N_6853,N_6937);
xnor U7106 (N_7106,N_6928,N_6918);
xor U7107 (N_7107,N_6815,N_6976);
xor U7108 (N_7108,N_6785,N_6759);
or U7109 (N_7109,N_6852,N_6767);
xnor U7110 (N_7110,N_6859,N_6891);
xor U7111 (N_7111,N_6874,N_6961);
xor U7112 (N_7112,N_6838,N_6843);
xor U7113 (N_7113,N_6988,N_6779);
and U7114 (N_7114,N_6880,N_6951);
or U7115 (N_7115,N_6796,N_6915);
nand U7116 (N_7116,N_6906,N_6858);
nor U7117 (N_7117,N_6832,N_6791);
and U7118 (N_7118,N_6878,N_6914);
and U7119 (N_7119,N_6892,N_6786);
xor U7120 (N_7120,N_6934,N_6995);
and U7121 (N_7121,N_6781,N_6897);
or U7122 (N_7122,N_6771,N_6982);
and U7123 (N_7123,N_6808,N_6794);
or U7124 (N_7124,N_6807,N_6887);
or U7125 (N_7125,N_6959,N_6826);
nand U7126 (N_7126,N_6762,N_6861);
nand U7127 (N_7127,N_6924,N_6898);
nor U7128 (N_7128,N_6770,N_6877);
or U7129 (N_7129,N_6814,N_6996);
nand U7130 (N_7130,N_6843,N_6811);
nand U7131 (N_7131,N_6977,N_6802);
nand U7132 (N_7132,N_6859,N_6838);
nor U7133 (N_7133,N_6753,N_6809);
xnor U7134 (N_7134,N_6937,N_6843);
or U7135 (N_7135,N_6933,N_6833);
or U7136 (N_7136,N_6935,N_6778);
xor U7137 (N_7137,N_6851,N_6955);
or U7138 (N_7138,N_6835,N_6901);
or U7139 (N_7139,N_6900,N_6938);
xor U7140 (N_7140,N_6790,N_6966);
nand U7141 (N_7141,N_6939,N_6840);
xnor U7142 (N_7142,N_6808,N_6949);
or U7143 (N_7143,N_6981,N_6769);
nand U7144 (N_7144,N_6787,N_6954);
xor U7145 (N_7145,N_6750,N_6951);
nor U7146 (N_7146,N_6889,N_6917);
nor U7147 (N_7147,N_6760,N_6948);
nand U7148 (N_7148,N_6830,N_6954);
nor U7149 (N_7149,N_6769,N_6947);
nand U7150 (N_7150,N_6822,N_6829);
xor U7151 (N_7151,N_6908,N_6845);
xor U7152 (N_7152,N_6838,N_6942);
nand U7153 (N_7153,N_6871,N_6824);
or U7154 (N_7154,N_6877,N_6959);
xor U7155 (N_7155,N_6808,N_6909);
or U7156 (N_7156,N_6762,N_6894);
and U7157 (N_7157,N_6764,N_6971);
and U7158 (N_7158,N_6943,N_6807);
nand U7159 (N_7159,N_6962,N_6815);
nor U7160 (N_7160,N_6902,N_6939);
or U7161 (N_7161,N_6758,N_6906);
nand U7162 (N_7162,N_6970,N_6971);
and U7163 (N_7163,N_6845,N_6768);
and U7164 (N_7164,N_6946,N_6861);
nor U7165 (N_7165,N_6760,N_6801);
and U7166 (N_7166,N_6780,N_6871);
xor U7167 (N_7167,N_6917,N_6914);
or U7168 (N_7168,N_6831,N_6942);
xor U7169 (N_7169,N_6947,N_6927);
xnor U7170 (N_7170,N_6789,N_6969);
nand U7171 (N_7171,N_6963,N_6942);
or U7172 (N_7172,N_6870,N_6838);
nor U7173 (N_7173,N_6896,N_6892);
or U7174 (N_7174,N_6951,N_6995);
xnor U7175 (N_7175,N_6937,N_6968);
nand U7176 (N_7176,N_6776,N_6872);
or U7177 (N_7177,N_6768,N_6890);
nor U7178 (N_7178,N_6914,N_6929);
and U7179 (N_7179,N_6922,N_6802);
and U7180 (N_7180,N_6945,N_6977);
xnor U7181 (N_7181,N_6923,N_6819);
and U7182 (N_7182,N_6794,N_6878);
nand U7183 (N_7183,N_6927,N_6778);
nor U7184 (N_7184,N_6895,N_6932);
nand U7185 (N_7185,N_6785,N_6842);
and U7186 (N_7186,N_6823,N_6833);
xor U7187 (N_7187,N_6929,N_6984);
nor U7188 (N_7188,N_6785,N_6906);
nor U7189 (N_7189,N_6900,N_6777);
xor U7190 (N_7190,N_6807,N_6895);
xor U7191 (N_7191,N_6934,N_6999);
nor U7192 (N_7192,N_6760,N_6789);
nor U7193 (N_7193,N_6926,N_6766);
nor U7194 (N_7194,N_6987,N_6896);
nor U7195 (N_7195,N_6890,N_6876);
nor U7196 (N_7196,N_6804,N_6755);
nand U7197 (N_7197,N_6985,N_6788);
xor U7198 (N_7198,N_6799,N_6837);
nor U7199 (N_7199,N_6996,N_6934);
xor U7200 (N_7200,N_6833,N_6974);
nand U7201 (N_7201,N_6898,N_6976);
and U7202 (N_7202,N_6835,N_6956);
nand U7203 (N_7203,N_6806,N_6816);
nor U7204 (N_7204,N_6835,N_6853);
nor U7205 (N_7205,N_6869,N_6834);
nor U7206 (N_7206,N_6799,N_6848);
nand U7207 (N_7207,N_6956,N_6995);
nand U7208 (N_7208,N_6952,N_6972);
xnor U7209 (N_7209,N_6992,N_6793);
or U7210 (N_7210,N_6776,N_6922);
nor U7211 (N_7211,N_6905,N_6835);
xor U7212 (N_7212,N_6990,N_6886);
nand U7213 (N_7213,N_6887,N_6926);
nand U7214 (N_7214,N_6954,N_6985);
xnor U7215 (N_7215,N_6924,N_6989);
or U7216 (N_7216,N_6831,N_6934);
and U7217 (N_7217,N_6765,N_6774);
nand U7218 (N_7218,N_6901,N_6841);
and U7219 (N_7219,N_6927,N_6922);
nand U7220 (N_7220,N_6754,N_6821);
and U7221 (N_7221,N_6755,N_6831);
and U7222 (N_7222,N_6768,N_6894);
and U7223 (N_7223,N_6956,N_6772);
nor U7224 (N_7224,N_6885,N_6818);
nor U7225 (N_7225,N_6814,N_6845);
nor U7226 (N_7226,N_6962,N_6912);
nand U7227 (N_7227,N_6936,N_6903);
nand U7228 (N_7228,N_6803,N_6882);
or U7229 (N_7229,N_6780,N_6799);
or U7230 (N_7230,N_6893,N_6948);
nand U7231 (N_7231,N_6822,N_6819);
nor U7232 (N_7232,N_6906,N_6804);
nand U7233 (N_7233,N_6811,N_6776);
or U7234 (N_7234,N_6959,N_6885);
nor U7235 (N_7235,N_6864,N_6817);
nand U7236 (N_7236,N_6875,N_6848);
or U7237 (N_7237,N_6771,N_6858);
nand U7238 (N_7238,N_6761,N_6762);
xor U7239 (N_7239,N_6922,N_6923);
and U7240 (N_7240,N_6873,N_6825);
nor U7241 (N_7241,N_6872,N_6891);
and U7242 (N_7242,N_6775,N_6857);
nor U7243 (N_7243,N_6994,N_6991);
and U7244 (N_7244,N_6926,N_6856);
nor U7245 (N_7245,N_6752,N_6845);
nand U7246 (N_7246,N_6805,N_6889);
xnor U7247 (N_7247,N_6800,N_6918);
or U7248 (N_7248,N_6846,N_6892);
xor U7249 (N_7249,N_6977,N_6830);
nor U7250 (N_7250,N_7076,N_7012);
nor U7251 (N_7251,N_7046,N_7157);
or U7252 (N_7252,N_7183,N_7019);
nand U7253 (N_7253,N_7205,N_7196);
and U7254 (N_7254,N_7179,N_7083);
and U7255 (N_7255,N_7241,N_7146);
xor U7256 (N_7256,N_7182,N_7118);
or U7257 (N_7257,N_7188,N_7151);
xnor U7258 (N_7258,N_7111,N_7153);
and U7259 (N_7259,N_7159,N_7036);
xnor U7260 (N_7260,N_7098,N_7197);
nand U7261 (N_7261,N_7053,N_7014);
xor U7262 (N_7262,N_7231,N_7123);
and U7263 (N_7263,N_7068,N_7247);
nand U7264 (N_7264,N_7212,N_7015);
xor U7265 (N_7265,N_7177,N_7035);
and U7266 (N_7266,N_7180,N_7218);
xnor U7267 (N_7267,N_7028,N_7104);
nor U7268 (N_7268,N_7087,N_7204);
nor U7269 (N_7269,N_7114,N_7061);
or U7270 (N_7270,N_7129,N_7049);
xnor U7271 (N_7271,N_7165,N_7216);
or U7272 (N_7272,N_7088,N_7007);
nand U7273 (N_7273,N_7060,N_7236);
and U7274 (N_7274,N_7033,N_7004);
and U7275 (N_7275,N_7184,N_7194);
nand U7276 (N_7276,N_7172,N_7121);
nor U7277 (N_7277,N_7213,N_7117);
and U7278 (N_7278,N_7168,N_7136);
xnor U7279 (N_7279,N_7243,N_7190);
nand U7280 (N_7280,N_7214,N_7025);
nand U7281 (N_7281,N_7181,N_7219);
and U7282 (N_7282,N_7145,N_7070);
xnor U7283 (N_7283,N_7020,N_7207);
xnor U7284 (N_7284,N_7072,N_7137);
xnor U7285 (N_7285,N_7127,N_7110);
nand U7286 (N_7286,N_7115,N_7154);
xor U7287 (N_7287,N_7034,N_7021);
and U7288 (N_7288,N_7043,N_7103);
or U7289 (N_7289,N_7189,N_7038);
and U7290 (N_7290,N_7006,N_7139);
or U7291 (N_7291,N_7191,N_7178);
or U7292 (N_7292,N_7078,N_7011);
or U7293 (N_7293,N_7002,N_7032);
xor U7294 (N_7294,N_7080,N_7091);
or U7295 (N_7295,N_7162,N_7031);
and U7296 (N_7296,N_7044,N_7164);
or U7297 (N_7297,N_7202,N_7167);
and U7298 (N_7298,N_7005,N_7186);
and U7299 (N_7299,N_7084,N_7106);
or U7300 (N_7300,N_7242,N_7239);
nor U7301 (N_7301,N_7171,N_7233);
nor U7302 (N_7302,N_7234,N_7039);
or U7303 (N_7303,N_7105,N_7187);
xor U7304 (N_7304,N_7126,N_7228);
xor U7305 (N_7305,N_7174,N_7211);
or U7306 (N_7306,N_7071,N_7100);
and U7307 (N_7307,N_7130,N_7238);
and U7308 (N_7308,N_7090,N_7010);
nor U7309 (N_7309,N_7166,N_7063);
or U7310 (N_7310,N_7237,N_7099);
nor U7311 (N_7311,N_7016,N_7023);
or U7312 (N_7312,N_7097,N_7086);
or U7313 (N_7313,N_7037,N_7064);
or U7314 (N_7314,N_7235,N_7081);
xor U7315 (N_7315,N_7108,N_7244);
nor U7316 (N_7316,N_7042,N_7109);
and U7317 (N_7317,N_7203,N_7215);
nor U7318 (N_7318,N_7200,N_7027);
and U7319 (N_7319,N_7067,N_7112);
nor U7320 (N_7320,N_7065,N_7169);
nand U7321 (N_7321,N_7226,N_7227);
xor U7322 (N_7322,N_7026,N_7249);
and U7323 (N_7323,N_7040,N_7024);
xor U7324 (N_7324,N_7000,N_7057);
or U7325 (N_7325,N_7066,N_7206);
nand U7326 (N_7326,N_7092,N_7147);
nand U7327 (N_7327,N_7142,N_7210);
nand U7328 (N_7328,N_7096,N_7009);
nor U7329 (N_7329,N_7119,N_7141);
xnor U7330 (N_7330,N_7245,N_7085);
nor U7331 (N_7331,N_7101,N_7116);
nand U7332 (N_7332,N_7017,N_7201);
and U7333 (N_7333,N_7133,N_7055);
nand U7334 (N_7334,N_7221,N_7192);
and U7335 (N_7335,N_7232,N_7173);
nand U7336 (N_7336,N_7124,N_7082);
and U7337 (N_7337,N_7229,N_7220);
nor U7338 (N_7338,N_7029,N_7059);
nand U7339 (N_7339,N_7048,N_7095);
nand U7340 (N_7340,N_7030,N_7208);
nand U7341 (N_7341,N_7125,N_7077);
xnor U7342 (N_7342,N_7193,N_7062);
and U7343 (N_7343,N_7158,N_7075);
nor U7344 (N_7344,N_7122,N_7069);
nand U7345 (N_7345,N_7209,N_7094);
nand U7346 (N_7346,N_7056,N_7051);
or U7347 (N_7347,N_7018,N_7003);
and U7348 (N_7348,N_7013,N_7223);
nor U7349 (N_7349,N_7170,N_7155);
and U7350 (N_7350,N_7185,N_7152);
or U7351 (N_7351,N_7176,N_7022);
or U7352 (N_7352,N_7161,N_7225);
and U7353 (N_7353,N_7131,N_7248);
or U7354 (N_7354,N_7001,N_7073);
xnor U7355 (N_7355,N_7198,N_7150);
xor U7356 (N_7356,N_7120,N_7041);
xnor U7357 (N_7357,N_7113,N_7102);
nor U7358 (N_7358,N_7240,N_7107);
or U7359 (N_7359,N_7160,N_7132);
xor U7360 (N_7360,N_7156,N_7093);
nor U7361 (N_7361,N_7230,N_7045);
xnor U7362 (N_7362,N_7222,N_7074);
and U7363 (N_7363,N_7199,N_7050);
nor U7364 (N_7364,N_7195,N_7163);
and U7365 (N_7365,N_7143,N_7079);
and U7366 (N_7366,N_7135,N_7138);
xnor U7367 (N_7367,N_7144,N_7058);
or U7368 (N_7368,N_7089,N_7047);
xor U7369 (N_7369,N_7008,N_7149);
xor U7370 (N_7370,N_7217,N_7054);
or U7371 (N_7371,N_7175,N_7052);
nand U7372 (N_7372,N_7224,N_7148);
nor U7373 (N_7373,N_7140,N_7128);
nand U7374 (N_7374,N_7134,N_7246);
xor U7375 (N_7375,N_7108,N_7242);
and U7376 (N_7376,N_7214,N_7053);
nand U7377 (N_7377,N_7177,N_7111);
nor U7378 (N_7378,N_7104,N_7029);
and U7379 (N_7379,N_7188,N_7186);
nor U7380 (N_7380,N_7149,N_7158);
or U7381 (N_7381,N_7179,N_7090);
and U7382 (N_7382,N_7088,N_7206);
and U7383 (N_7383,N_7249,N_7160);
nand U7384 (N_7384,N_7002,N_7188);
xor U7385 (N_7385,N_7035,N_7062);
or U7386 (N_7386,N_7121,N_7161);
xor U7387 (N_7387,N_7106,N_7186);
nand U7388 (N_7388,N_7166,N_7049);
nor U7389 (N_7389,N_7177,N_7076);
or U7390 (N_7390,N_7078,N_7162);
or U7391 (N_7391,N_7108,N_7101);
nand U7392 (N_7392,N_7066,N_7009);
nor U7393 (N_7393,N_7163,N_7062);
nor U7394 (N_7394,N_7127,N_7062);
nand U7395 (N_7395,N_7003,N_7095);
or U7396 (N_7396,N_7007,N_7076);
or U7397 (N_7397,N_7210,N_7108);
or U7398 (N_7398,N_7006,N_7223);
xnor U7399 (N_7399,N_7112,N_7019);
or U7400 (N_7400,N_7156,N_7104);
and U7401 (N_7401,N_7108,N_7193);
nor U7402 (N_7402,N_7148,N_7111);
or U7403 (N_7403,N_7088,N_7204);
and U7404 (N_7404,N_7145,N_7101);
nand U7405 (N_7405,N_7132,N_7049);
nand U7406 (N_7406,N_7068,N_7185);
xnor U7407 (N_7407,N_7126,N_7066);
nor U7408 (N_7408,N_7128,N_7157);
or U7409 (N_7409,N_7044,N_7236);
or U7410 (N_7410,N_7058,N_7106);
nand U7411 (N_7411,N_7096,N_7218);
xnor U7412 (N_7412,N_7102,N_7081);
or U7413 (N_7413,N_7139,N_7231);
nand U7414 (N_7414,N_7136,N_7235);
nor U7415 (N_7415,N_7054,N_7067);
xor U7416 (N_7416,N_7020,N_7083);
nor U7417 (N_7417,N_7044,N_7110);
or U7418 (N_7418,N_7147,N_7060);
xnor U7419 (N_7419,N_7173,N_7152);
and U7420 (N_7420,N_7160,N_7226);
or U7421 (N_7421,N_7222,N_7108);
xnor U7422 (N_7422,N_7224,N_7037);
nand U7423 (N_7423,N_7248,N_7163);
xnor U7424 (N_7424,N_7036,N_7120);
and U7425 (N_7425,N_7103,N_7126);
nand U7426 (N_7426,N_7072,N_7188);
and U7427 (N_7427,N_7178,N_7023);
nand U7428 (N_7428,N_7223,N_7135);
or U7429 (N_7429,N_7024,N_7038);
nand U7430 (N_7430,N_7150,N_7069);
nor U7431 (N_7431,N_7104,N_7215);
xor U7432 (N_7432,N_7047,N_7223);
nor U7433 (N_7433,N_7212,N_7060);
xnor U7434 (N_7434,N_7074,N_7034);
nand U7435 (N_7435,N_7039,N_7154);
and U7436 (N_7436,N_7228,N_7152);
xnor U7437 (N_7437,N_7030,N_7179);
nor U7438 (N_7438,N_7183,N_7199);
xnor U7439 (N_7439,N_7225,N_7019);
or U7440 (N_7440,N_7184,N_7200);
nor U7441 (N_7441,N_7172,N_7038);
nor U7442 (N_7442,N_7120,N_7060);
and U7443 (N_7443,N_7055,N_7035);
nor U7444 (N_7444,N_7015,N_7191);
and U7445 (N_7445,N_7063,N_7038);
or U7446 (N_7446,N_7000,N_7183);
or U7447 (N_7447,N_7196,N_7097);
xnor U7448 (N_7448,N_7106,N_7147);
and U7449 (N_7449,N_7145,N_7130);
nor U7450 (N_7450,N_7203,N_7168);
nor U7451 (N_7451,N_7108,N_7042);
and U7452 (N_7452,N_7118,N_7031);
nor U7453 (N_7453,N_7004,N_7061);
and U7454 (N_7454,N_7185,N_7229);
or U7455 (N_7455,N_7080,N_7127);
and U7456 (N_7456,N_7044,N_7171);
or U7457 (N_7457,N_7243,N_7149);
xnor U7458 (N_7458,N_7189,N_7153);
or U7459 (N_7459,N_7247,N_7085);
nand U7460 (N_7460,N_7189,N_7101);
nor U7461 (N_7461,N_7072,N_7116);
xnor U7462 (N_7462,N_7109,N_7113);
nor U7463 (N_7463,N_7087,N_7031);
nand U7464 (N_7464,N_7237,N_7002);
or U7465 (N_7465,N_7044,N_7090);
and U7466 (N_7466,N_7013,N_7235);
nand U7467 (N_7467,N_7037,N_7187);
nand U7468 (N_7468,N_7123,N_7078);
nor U7469 (N_7469,N_7078,N_7216);
nor U7470 (N_7470,N_7206,N_7197);
nand U7471 (N_7471,N_7036,N_7075);
and U7472 (N_7472,N_7150,N_7025);
nand U7473 (N_7473,N_7021,N_7008);
and U7474 (N_7474,N_7083,N_7011);
and U7475 (N_7475,N_7098,N_7147);
or U7476 (N_7476,N_7023,N_7073);
xnor U7477 (N_7477,N_7171,N_7165);
and U7478 (N_7478,N_7244,N_7173);
and U7479 (N_7479,N_7126,N_7039);
or U7480 (N_7480,N_7238,N_7020);
nand U7481 (N_7481,N_7167,N_7126);
and U7482 (N_7482,N_7088,N_7139);
xor U7483 (N_7483,N_7175,N_7207);
xor U7484 (N_7484,N_7087,N_7111);
or U7485 (N_7485,N_7047,N_7171);
nor U7486 (N_7486,N_7238,N_7243);
or U7487 (N_7487,N_7055,N_7200);
or U7488 (N_7488,N_7035,N_7026);
nor U7489 (N_7489,N_7166,N_7096);
and U7490 (N_7490,N_7180,N_7042);
or U7491 (N_7491,N_7157,N_7229);
and U7492 (N_7492,N_7168,N_7223);
nor U7493 (N_7493,N_7237,N_7138);
xnor U7494 (N_7494,N_7026,N_7070);
nor U7495 (N_7495,N_7077,N_7160);
or U7496 (N_7496,N_7046,N_7214);
nand U7497 (N_7497,N_7082,N_7194);
xor U7498 (N_7498,N_7042,N_7016);
xor U7499 (N_7499,N_7134,N_7052);
or U7500 (N_7500,N_7364,N_7410);
or U7501 (N_7501,N_7391,N_7283);
nand U7502 (N_7502,N_7279,N_7417);
or U7503 (N_7503,N_7304,N_7382);
or U7504 (N_7504,N_7483,N_7258);
nand U7505 (N_7505,N_7250,N_7374);
or U7506 (N_7506,N_7274,N_7386);
nor U7507 (N_7507,N_7438,N_7300);
or U7508 (N_7508,N_7497,N_7331);
nand U7509 (N_7509,N_7440,N_7394);
and U7510 (N_7510,N_7351,N_7339);
or U7511 (N_7511,N_7381,N_7439);
xnor U7512 (N_7512,N_7491,N_7421);
xor U7513 (N_7513,N_7401,N_7356);
nor U7514 (N_7514,N_7414,N_7366);
and U7515 (N_7515,N_7253,N_7294);
and U7516 (N_7516,N_7388,N_7392);
or U7517 (N_7517,N_7474,N_7475);
nor U7518 (N_7518,N_7457,N_7435);
xnor U7519 (N_7519,N_7499,N_7349);
or U7520 (N_7520,N_7313,N_7334);
or U7521 (N_7521,N_7390,N_7275);
nand U7522 (N_7522,N_7252,N_7357);
xor U7523 (N_7523,N_7473,N_7362);
nand U7524 (N_7524,N_7321,N_7345);
and U7525 (N_7525,N_7376,N_7324);
xnor U7526 (N_7526,N_7299,N_7288);
and U7527 (N_7527,N_7437,N_7365);
and U7528 (N_7528,N_7347,N_7477);
xor U7529 (N_7529,N_7260,N_7416);
xnor U7530 (N_7530,N_7389,N_7293);
or U7531 (N_7531,N_7261,N_7450);
nand U7532 (N_7532,N_7480,N_7444);
xnor U7533 (N_7533,N_7269,N_7367);
xnor U7534 (N_7534,N_7340,N_7485);
and U7535 (N_7535,N_7470,N_7441);
or U7536 (N_7536,N_7354,N_7335);
nor U7537 (N_7537,N_7436,N_7447);
nor U7538 (N_7538,N_7251,N_7433);
or U7539 (N_7539,N_7396,N_7449);
xor U7540 (N_7540,N_7492,N_7412);
nand U7541 (N_7541,N_7307,N_7332);
or U7542 (N_7542,N_7338,N_7282);
or U7543 (N_7543,N_7264,N_7445);
nor U7544 (N_7544,N_7478,N_7325);
xor U7545 (N_7545,N_7272,N_7333);
nor U7546 (N_7546,N_7378,N_7284);
xnor U7547 (N_7547,N_7400,N_7326);
or U7548 (N_7548,N_7327,N_7434);
xnor U7549 (N_7549,N_7476,N_7271);
nand U7550 (N_7550,N_7432,N_7280);
xor U7551 (N_7551,N_7496,N_7442);
and U7552 (N_7552,N_7419,N_7346);
and U7553 (N_7553,N_7263,N_7256);
nor U7554 (N_7554,N_7430,N_7418);
or U7555 (N_7555,N_7296,N_7454);
or U7556 (N_7556,N_7486,N_7393);
and U7557 (N_7557,N_7451,N_7377);
or U7558 (N_7558,N_7494,N_7289);
xnor U7559 (N_7559,N_7472,N_7471);
xnor U7560 (N_7560,N_7341,N_7452);
nor U7561 (N_7561,N_7318,N_7427);
and U7562 (N_7562,N_7411,N_7460);
nand U7563 (N_7563,N_7461,N_7479);
or U7564 (N_7564,N_7459,N_7311);
or U7565 (N_7565,N_7397,N_7404);
or U7566 (N_7566,N_7387,N_7265);
and U7567 (N_7567,N_7384,N_7355);
xor U7568 (N_7568,N_7266,N_7484);
and U7569 (N_7569,N_7425,N_7488);
nand U7570 (N_7570,N_7462,N_7295);
or U7571 (N_7571,N_7270,N_7358);
nor U7572 (N_7572,N_7276,N_7398);
and U7573 (N_7573,N_7361,N_7422);
nand U7574 (N_7574,N_7286,N_7466);
or U7575 (N_7575,N_7257,N_7302);
or U7576 (N_7576,N_7278,N_7353);
and U7577 (N_7577,N_7385,N_7262);
nand U7578 (N_7578,N_7343,N_7373);
and U7579 (N_7579,N_7429,N_7352);
nand U7580 (N_7580,N_7489,N_7424);
or U7581 (N_7581,N_7330,N_7281);
or U7582 (N_7582,N_7490,N_7464);
nor U7583 (N_7583,N_7453,N_7426);
xnor U7584 (N_7584,N_7405,N_7254);
xor U7585 (N_7585,N_7255,N_7312);
or U7586 (N_7586,N_7370,N_7360);
xor U7587 (N_7587,N_7322,N_7431);
nor U7588 (N_7588,N_7369,N_7399);
nand U7589 (N_7589,N_7359,N_7290);
nand U7590 (N_7590,N_7305,N_7423);
nand U7591 (N_7591,N_7277,N_7337);
nor U7592 (N_7592,N_7380,N_7498);
nand U7593 (N_7593,N_7409,N_7446);
nand U7594 (N_7594,N_7487,N_7448);
or U7595 (N_7595,N_7482,N_7292);
nor U7596 (N_7596,N_7316,N_7420);
nand U7597 (N_7597,N_7303,N_7465);
nand U7598 (N_7598,N_7315,N_7363);
nand U7599 (N_7599,N_7402,N_7308);
and U7600 (N_7600,N_7371,N_7481);
or U7601 (N_7601,N_7350,N_7291);
or U7602 (N_7602,N_7467,N_7495);
nand U7603 (N_7603,N_7259,N_7317);
xor U7604 (N_7604,N_7395,N_7415);
nor U7605 (N_7605,N_7458,N_7320);
nor U7606 (N_7606,N_7379,N_7323);
nand U7607 (N_7607,N_7328,N_7463);
nor U7608 (N_7608,N_7336,N_7314);
and U7609 (N_7609,N_7267,N_7443);
nand U7610 (N_7610,N_7297,N_7301);
and U7611 (N_7611,N_7403,N_7348);
nand U7612 (N_7612,N_7408,N_7287);
xor U7613 (N_7613,N_7319,N_7428);
and U7614 (N_7614,N_7306,N_7329);
nand U7615 (N_7615,N_7375,N_7298);
xor U7616 (N_7616,N_7383,N_7469);
and U7617 (N_7617,N_7285,N_7268);
or U7618 (N_7618,N_7372,N_7455);
nor U7619 (N_7619,N_7406,N_7407);
nor U7620 (N_7620,N_7273,N_7309);
or U7621 (N_7621,N_7342,N_7413);
nor U7622 (N_7622,N_7344,N_7368);
nor U7623 (N_7623,N_7468,N_7456);
and U7624 (N_7624,N_7310,N_7493);
or U7625 (N_7625,N_7496,N_7418);
nand U7626 (N_7626,N_7366,N_7470);
nand U7627 (N_7627,N_7404,N_7367);
nand U7628 (N_7628,N_7278,N_7372);
nand U7629 (N_7629,N_7375,N_7301);
or U7630 (N_7630,N_7384,N_7257);
or U7631 (N_7631,N_7269,N_7289);
nor U7632 (N_7632,N_7398,N_7466);
or U7633 (N_7633,N_7377,N_7351);
and U7634 (N_7634,N_7306,N_7494);
nor U7635 (N_7635,N_7493,N_7490);
xnor U7636 (N_7636,N_7457,N_7307);
xnor U7637 (N_7637,N_7393,N_7398);
and U7638 (N_7638,N_7461,N_7368);
nor U7639 (N_7639,N_7373,N_7267);
and U7640 (N_7640,N_7493,N_7374);
or U7641 (N_7641,N_7252,N_7404);
and U7642 (N_7642,N_7267,N_7491);
nand U7643 (N_7643,N_7414,N_7423);
nand U7644 (N_7644,N_7389,N_7351);
nor U7645 (N_7645,N_7452,N_7295);
xnor U7646 (N_7646,N_7291,N_7311);
nor U7647 (N_7647,N_7459,N_7384);
xor U7648 (N_7648,N_7472,N_7446);
nor U7649 (N_7649,N_7470,N_7264);
nor U7650 (N_7650,N_7427,N_7433);
xnor U7651 (N_7651,N_7379,N_7278);
xnor U7652 (N_7652,N_7418,N_7342);
and U7653 (N_7653,N_7301,N_7419);
nor U7654 (N_7654,N_7374,N_7469);
xnor U7655 (N_7655,N_7400,N_7263);
xor U7656 (N_7656,N_7480,N_7326);
or U7657 (N_7657,N_7280,N_7456);
or U7658 (N_7658,N_7260,N_7375);
nand U7659 (N_7659,N_7347,N_7376);
nor U7660 (N_7660,N_7283,N_7306);
or U7661 (N_7661,N_7439,N_7480);
nand U7662 (N_7662,N_7321,N_7376);
nor U7663 (N_7663,N_7497,N_7460);
xnor U7664 (N_7664,N_7423,N_7382);
nor U7665 (N_7665,N_7277,N_7288);
and U7666 (N_7666,N_7352,N_7395);
or U7667 (N_7667,N_7308,N_7278);
and U7668 (N_7668,N_7471,N_7349);
xnor U7669 (N_7669,N_7278,N_7403);
or U7670 (N_7670,N_7451,N_7397);
and U7671 (N_7671,N_7425,N_7332);
xor U7672 (N_7672,N_7479,N_7434);
xor U7673 (N_7673,N_7260,N_7328);
and U7674 (N_7674,N_7299,N_7359);
or U7675 (N_7675,N_7460,N_7393);
or U7676 (N_7676,N_7499,N_7274);
xor U7677 (N_7677,N_7346,N_7307);
nor U7678 (N_7678,N_7304,N_7330);
nor U7679 (N_7679,N_7346,N_7283);
nor U7680 (N_7680,N_7445,N_7492);
and U7681 (N_7681,N_7481,N_7269);
nor U7682 (N_7682,N_7269,N_7447);
or U7683 (N_7683,N_7290,N_7307);
nand U7684 (N_7684,N_7471,N_7362);
and U7685 (N_7685,N_7332,N_7293);
or U7686 (N_7686,N_7309,N_7355);
nand U7687 (N_7687,N_7499,N_7350);
nor U7688 (N_7688,N_7383,N_7322);
or U7689 (N_7689,N_7491,N_7294);
nand U7690 (N_7690,N_7357,N_7460);
or U7691 (N_7691,N_7259,N_7292);
nor U7692 (N_7692,N_7359,N_7477);
xor U7693 (N_7693,N_7430,N_7362);
xor U7694 (N_7694,N_7493,N_7487);
nor U7695 (N_7695,N_7387,N_7492);
and U7696 (N_7696,N_7251,N_7469);
or U7697 (N_7697,N_7485,N_7298);
and U7698 (N_7698,N_7463,N_7281);
xnor U7699 (N_7699,N_7352,N_7499);
or U7700 (N_7700,N_7486,N_7333);
nor U7701 (N_7701,N_7406,N_7328);
nor U7702 (N_7702,N_7251,N_7254);
or U7703 (N_7703,N_7254,N_7425);
or U7704 (N_7704,N_7484,N_7443);
nor U7705 (N_7705,N_7430,N_7376);
nand U7706 (N_7706,N_7354,N_7253);
and U7707 (N_7707,N_7497,N_7277);
or U7708 (N_7708,N_7282,N_7336);
or U7709 (N_7709,N_7432,N_7411);
and U7710 (N_7710,N_7350,N_7267);
or U7711 (N_7711,N_7287,N_7399);
xor U7712 (N_7712,N_7358,N_7410);
and U7713 (N_7713,N_7311,N_7379);
and U7714 (N_7714,N_7364,N_7369);
nor U7715 (N_7715,N_7415,N_7354);
nand U7716 (N_7716,N_7257,N_7435);
and U7717 (N_7717,N_7287,N_7286);
or U7718 (N_7718,N_7393,N_7440);
and U7719 (N_7719,N_7433,N_7261);
or U7720 (N_7720,N_7343,N_7418);
and U7721 (N_7721,N_7453,N_7275);
and U7722 (N_7722,N_7426,N_7263);
and U7723 (N_7723,N_7339,N_7270);
or U7724 (N_7724,N_7253,N_7319);
and U7725 (N_7725,N_7256,N_7251);
and U7726 (N_7726,N_7378,N_7494);
xor U7727 (N_7727,N_7335,N_7290);
and U7728 (N_7728,N_7438,N_7338);
and U7729 (N_7729,N_7331,N_7309);
xor U7730 (N_7730,N_7279,N_7466);
or U7731 (N_7731,N_7436,N_7499);
xor U7732 (N_7732,N_7332,N_7336);
nand U7733 (N_7733,N_7294,N_7320);
xnor U7734 (N_7734,N_7371,N_7449);
nor U7735 (N_7735,N_7267,N_7445);
or U7736 (N_7736,N_7338,N_7325);
or U7737 (N_7737,N_7422,N_7478);
and U7738 (N_7738,N_7342,N_7457);
nor U7739 (N_7739,N_7315,N_7422);
xor U7740 (N_7740,N_7316,N_7434);
nor U7741 (N_7741,N_7273,N_7331);
nand U7742 (N_7742,N_7347,N_7372);
and U7743 (N_7743,N_7345,N_7412);
and U7744 (N_7744,N_7437,N_7408);
or U7745 (N_7745,N_7406,N_7466);
or U7746 (N_7746,N_7273,N_7356);
nor U7747 (N_7747,N_7251,N_7429);
and U7748 (N_7748,N_7376,N_7459);
and U7749 (N_7749,N_7402,N_7459);
and U7750 (N_7750,N_7501,N_7706);
nor U7751 (N_7751,N_7574,N_7687);
nor U7752 (N_7752,N_7597,N_7600);
or U7753 (N_7753,N_7726,N_7683);
and U7754 (N_7754,N_7567,N_7700);
nand U7755 (N_7755,N_7662,N_7565);
or U7756 (N_7756,N_7697,N_7592);
and U7757 (N_7757,N_7663,N_7715);
nand U7758 (N_7758,N_7576,N_7545);
nand U7759 (N_7759,N_7743,N_7618);
nor U7760 (N_7760,N_7611,N_7729);
and U7761 (N_7761,N_7733,N_7735);
xnor U7762 (N_7762,N_7710,N_7608);
xnor U7763 (N_7763,N_7723,N_7630);
and U7764 (N_7764,N_7605,N_7676);
and U7765 (N_7765,N_7519,N_7581);
xor U7766 (N_7766,N_7626,N_7711);
and U7767 (N_7767,N_7577,N_7691);
xnor U7768 (N_7768,N_7699,N_7705);
and U7769 (N_7769,N_7725,N_7516);
and U7770 (N_7770,N_7526,N_7507);
or U7771 (N_7771,N_7696,N_7669);
xnor U7772 (N_7772,N_7732,N_7503);
xnor U7773 (N_7773,N_7606,N_7547);
and U7774 (N_7774,N_7544,N_7745);
xnor U7775 (N_7775,N_7601,N_7553);
and U7776 (N_7776,N_7742,N_7744);
nor U7777 (N_7777,N_7656,N_7555);
nor U7778 (N_7778,N_7677,N_7635);
nor U7779 (N_7779,N_7511,N_7746);
xor U7780 (N_7780,N_7655,N_7649);
xor U7781 (N_7781,N_7632,N_7653);
xor U7782 (N_7782,N_7564,N_7651);
or U7783 (N_7783,N_7747,N_7595);
nor U7784 (N_7784,N_7578,N_7690);
and U7785 (N_7785,N_7563,N_7532);
or U7786 (N_7786,N_7510,N_7612);
and U7787 (N_7787,N_7659,N_7521);
xnor U7788 (N_7788,N_7522,N_7708);
or U7789 (N_7789,N_7739,N_7622);
xnor U7790 (N_7790,N_7625,N_7624);
and U7791 (N_7791,N_7554,N_7568);
xor U7792 (N_7792,N_7712,N_7589);
and U7793 (N_7793,N_7566,N_7702);
and U7794 (N_7794,N_7513,N_7551);
xor U7795 (N_7795,N_7598,N_7720);
or U7796 (N_7796,N_7514,N_7685);
and U7797 (N_7797,N_7546,N_7628);
nor U7798 (N_7798,N_7562,N_7693);
nand U7799 (N_7799,N_7692,N_7665);
nand U7800 (N_7800,N_7714,N_7643);
nand U7801 (N_7801,N_7550,N_7536);
nand U7802 (N_7802,N_7637,N_7585);
nor U7803 (N_7803,N_7530,N_7583);
and U7804 (N_7804,N_7542,N_7572);
xnor U7805 (N_7805,N_7541,N_7640);
and U7806 (N_7806,N_7737,N_7638);
and U7807 (N_7807,N_7686,N_7664);
and U7808 (N_7808,N_7703,N_7641);
nor U7809 (N_7809,N_7548,N_7504);
nand U7810 (N_7810,N_7525,N_7500);
xor U7811 (N_7811,N_7650,N_7661);
xor U7812 (N_7812,N_7681,N_7556);
xor U7813 (N_7813,N_7694,N_7730);
nor U7814 (N_7814,N_7623,N_7678);
nand U7815 (N_7815,N_7658,N_7538);
and U7816 (N_7816,N_7552,N_7736);
xnor U7817 (N_7817,N_7561,N_7518);
or U7818 (N_7818,N_7543,N_7588);
nand U7819 (N_7819,N_7717,N_7593);
nand U7820 (N_7820,N_7602,N_7594);
nand U7821 (N_7821,N_7657,N_7528);
nand U7822 (N_7822,N_7679,N_7629);
or U7823 (N_7823,N_7724,N_7698);
and U7824 (N_7824,N_7573,N_7533);
and U7825 (N_7825,N_7741,N_7614);
and U7826 (N_7826,N_7560,N_7660);
nor U7827 (N_7827,N_7520,N_7738);
nand U7828 (N_7828,N_7701,N_7529);
nand U7829 (N_7829,N_7722,N_7680);
nor U7830 (N_7830,N_7673,N_7689);
nand U7831 (N_7831,N_7627,N_7579);
nand U7832 (N_7832,N_7666,N_7534);
nor U7833 (N_7833,N_7642,N_7636);
xor U7834 (N_7834,N_7549,N_7539);
and U7835 (N_7835,N_7684,N_7506);
xor U7836 (N_7836,N_7675,N_7639);
nor U7837 (N_7837,N_7569,N_7604);
xnor U7838 (N_7838,N_7652,N_7575);
or U7839 (N_7839,N_7648,N_7617);
nand U7840 (N_7840,N_7587,N_7570);
or U7841 (N_7841,N_7671,N_7704);
nand U7842 (N_7842,N_7670,N_7749);
and U7843 (N_7843,N_7505,N_7557);
xnor U7844 (N_7844,N_7633,N_7709);
xnor U7845 (N_7845,N_7695,N_7674);
nand U7846 (N_7846,N_7740,N_7668);
nor U7847 (N_7847,N_7716,N_7609);
or U7848 (N_7848,N_7582,N_7527);
and U7849 (N_7849,N_7512,N_7728);
and U7850 (N_7850,N_7707,N_7508);
and U7851 (N_7851,N_7616,N_7631);
xor U7852 (N_7852,N_7644,N_7731);
and U7853 (N_7853,N_7603,N_7517);
xor U7854 (N_7854,N_7531,N_7615);
xnor U7855 (N_7855,N_7502,N_7591);
nand U7856 (N_7856,N_7721,N_7596);
and U7857 (N_7857,N_7584,N_7509);
xor U7858 (N_7858,N_7580,N_7537);
nor U7859 (N_7859,N_7515,N_7734);
and U7860 (N_7860,N_7559,N_7634);
and U7861 (N_7861,N_7610,N_7647);
nor U7862 (N_7862,N_7672,N_7571);
xor U7863 (N_7863,N_7727,N_7599);
nor U7864 (N_7864,N_7682,N_7558);
or U7865 (N_7865,N_7535,N_7523);
or U7866 (N_7866,N_7667,N_7718);
nor U7867 (N_7867,N_7613,N_7719);
nand U7868 (N_7868,N_7524,N_7586);
nor U7869 (N_7869,N_7713,N_7619);
or U7870 (N_7870,N_7654,N_7590);
nor U7871 (N_7871,N_7645,N_7688);
nand U7872 (N_7872,N_7621,N_7607);
nor U7873 (N_7873,N_7540,N_7646);
and U7874 (N_7874,N_7748,N_7620);
nand U7875 (N_7875,N_7700,N_7599);
nand U7876 (N_7876,N_7715,N_7684);
and U7877 (N_7877,N_7570,N_7642);
and U7878 (N_7878,N_7563,N_7615);
xnor U7879 (N_7879,N_7618,N_7549);
nor U7880 (N_7880,N_7680,N_7636);
xnor U7881 (N_7881,N_7575,N_7748);
or U7882 (N_7882,N_7584,N_7578);
nor U7883 (N_7883,N_7749,N_7727);
nand U7884 (N_7884,N_7649,N_7513);
or U7885 (N_7885,N_7612,N_7722);
xor U7886 (N_7886,N_7654,N_7655);
and U7887 (N_7887,N_7517,N_7669);
or U7888 (N_7888,N_7513,N_7564);
and U7889 (N_7889,N_7700,N_7514);
and U7890 (N_7890,N_7577,N_7684);
xor U7891 (N_7891,N_7564,N_7588);
nand U7892 (N_7892,N_7528,N_7701);
nor U7893 (N_7893,N_7669,N_7682);
and U7894 (N_7894,N_7661,N_7730);
nor U7895 (N_7895,N_7673,N_7745);
nand U7896 (N_7896,N_7521,N_7742);
and U7897 (N_7897,N_7727,N_7510);
and U7898 (N_7898,N_7683,N_7637);
nand U7899 (N_7899,N_7591,N_7667);
nand U7900 (N_7900,N_7582,N_7562);
and U7901 (N_7901,N_7690,N_7731);
or U7902 (N_7902,N_7594,N_7515);
nand U7903 (N_7903,N_7542,N_7595);
and U7904 (N_7904,N_7731,N_7563);
nand U7905 (N_7905,N_7724,N_7661);
and U7906 (N_7906,N_7690,N_7516);
nor U7907 (N_7907,N_7703,N_7633);
or U7908 (N_7908,N_7512,N_7735);
nand U7909 (N_7909,N_7623,N_7538);
nor U7910 (N_7910,N_7692,N_7636);
nor U7911 (N_7911,N_7629,N_7724);
xor U7912 (N_7912,N_7651,N_7558);
nor U7913 (N_7913,N_7578,N_7683);
and U7914 (N_7914,N_7734,N_7631);
nand U7915 (N_7915,N_7709,N_7664);
or U7916 (N_7916,N_7664,N_7502);
nor U7917 (N_7917,N_7531,N_7665);
and U7918 (N_7918,N_7556,N_7522);
or U7919 (N_7919,N_7736,N_7679);
or U7920 (N_7920,N_7647,N_7620);
nand U7921 (N_7921,N_7725,N_7551);
xor U7922 (N_7922,N_7610,N_7633);
and U7923 (N_7923,N_7556,N_7748);
or U7924 (N_7924,N_7560,N_7680);
nand U7925 (N_7925,N_7571,N_7557);
xnor U7926 (N_7926,N_7729,N_7628);
or U7927 (N_7927,N_7649,N_7536);
and U7928 (N_7928,N_7585,N_7697);
or U7929 (N_7929,N_7615,N_7519);
and U7930 (N_7930,N_7581,N_7598);
and U7931 (N_7931,N_7530,N_7608);
nor U7932 (N_7932,N_7581,N_7670);
nand U7933 (N_7933,N_7734,N_7532);
nor U7934 (N_7934,N_7550,N_7618);
xnor U7935 (N_7935,N_7634,N_7566);
xor U7936 (N_7936,N_7746,N_7616);
nand U7937 (N_7937,N_7632,N_7520);
or U7938 (N_7938,N_7726,N_7737);
xnor U7939 (N_7939,N_7556,N_7534);
or U7940 (N_7940,N_7598,N_7516);
xor U7941 (N_7941,N_7531,N_7631);
nor U7942 (N_7942,N_7533,N_7709);
and U7943 (N_7943,N_7528,N_7564);
nor U7944 (N_7944,N_7627,N_7694);
or U7945 (N_7945,N_7543,N_7709);
or U7946 (N_7946,N_7504,N_7560);
nand U7947 (N_7947,N_7525,N_7588);
and U7948 (N_7948,N_7627,N_7558);
xnor U7949 (N_7949,N_7636,N_7645);
and U7950 (N_7950,N_7741,N_7552);
nand U7951 (N_7951,N_7726,N_7510);
and U7952 (N_7952,N_7698,N_7590);
xor U7953 (N_7953,N_7593,N_7680);
and U7954 (N_7954,N_7671,N_7560);
xor U7955 (N_7955,N_7556,N_7532);
and U7956 (N_7956,N_7672,N_7595);
xor U7957 (N_7957,N_7600,N_7502);
nand U7958 (N_7958,N_7640,N_7542);
and U7959 (N_7959,N_7594,N_7741);
and U7960 (N_7960,N_7536,N_7510);
xor U7961 (N_7961,N_7645,N_7623);
xor U7962 (N_7962,N_7721,N_7585);
nand U7963 (N_7963,N_7588,N_7701);
or U7964 (N_7964,N_7714,N_7646);
and U7965 (N_7965,N_7529,N_7607);
nand U7966 (N_7966,N_7638,N_7659);
nor U7967 (N_7967,N_7553,N_7743);
xor U7968 (N_7968,N_7722,N_7535);
xor U7969 (N_7969,N_7607,N_7691);
or U7970 (N_7970,N_7649,N_7681);
or U7971 (N_7971,N_7676,N_7656);
nand U7972 (N_7972,N_7671,N_7722);
nand U7973 (N_7973,N_7628,N_7555);
nand U7974 (N_7974,N_7675,N_7717);
xnor U7975 (N_7975,N_7588,N_7609);
nor U7976 (N_7976,N_7670,N_7713);
or U7977 (N_7977,N_7532,N_7652);
nand U7978 (N_7978,N_7584,N_7616);
and U7979 (N_7979,N_7721,N_7602);
xnor U7980 (N_7980,N_7633,N_7533);
or U7981 (N_7981,N_7601,N_7690);
nand U7982 (N_7982,N_7558,N_7700);
xnor U7983 (N_7983,N_7564,N_7566);
and U7984 (N_7984,N_7627,N_7705);
nor U7985 (N_7985,N_7587,N_7535);
and U7986 (N_7986,N_7572,N_7619);
nand U7987 (N_7987,N_7618,N_7572);
and U7988 (N_7988,N_7639,N_7553);
nor U7989 (N_7989,N_7581,N_7524);
nor U7990 (N_7990,N_7569,N_7714);
xor U7991 (N_7991,N_7737,N_7528);
and U7992 (N_7992,N_7717,N_7545);
nand U7993 (N_7993,N_7536,N_7670);
nor U7994 (N_7994,N_7598,N_7544);
or U7995 (N_7995,N_7583,N_7618);
or U7996 (N_7996,N_7632,N_7597);
xor U7997 (N_7997,N_7591,N_7603);
and U7998 (N_7998,N_7616,N_7619);
and U7999 (N_7999,N_7548,N_7588);
and U8000 (N_8000,N_7764,N_7844);
xor U8001 (N_8001,N_7952,N_7885);
and U8002 (N_8002,N_7767,N_7772);
and U8003 (N_8003,N_7963,N_7752);
nand U8004 (N_8004,N_7912,N_7909);
xor U8005 (N_8005,N_7869,N_7804);
or U8006 (N_8006,N_7968,N_7888);
nand U8007 (N_8007,N_7874,N_7945);
or U8008 (N_8008,N_7791,N_7876);
nand U8009 (N_8009,N_7796,N_7965);
nor U8010 (N_8010,N_7838,N_7935);
nor U8011 (N_8011,N_7982,N_7851);
nor U8012 (N_8012,N_7793,N_7998);
or U8013 (N_8013,N_7760,N_7921);
xor U8014 (N_8014,N_7959,N_7900);
and U8015 (N_8015,N_7755,N_7992);
or U8016 (N_8016,N_7815,N_7894);
and U8017 (N_8017,N_7865,N_7908);
or U8018 (N_8018,N_7957,N_7800);
or U8019 (N_8019,N_7941,N_7899);
nand U8020 (N_8020,N_7821,N_7848);
xor U8021 (N_8021,N_7973,N_7811);
and U8022 (N_8022,N_7829,N_7843);
nor U8023 (N_8023,N_7798,N_7886);
nor U8024 (N_8024,N_7757,N_7814);
nand U8025 (N_8025,N_7940,N_7769);
or U8026 (N_8026,N_7771,N_7847);
and U8027 (N_8027,N_7871,N_7987);
xnor U8028 (N_8028,N_7766,N_7839);
xnor U8029 (N_8029,N_7884,N_7823);
nor U8030 (N_8030,N_7993,N_7972);
and U8031 (N_8031,N_7974,N_7975);
xnor U8032 (N_8032,N_7939,N_7873);
and U8033 (N_8033,N_7761,N_7901);
or U8034 (N_8034,N_7954,N_7787);
or U8035 (N_8035,N_7898,N_7933);
nor U8036 (N_8036,N_7961,N_7845);
nor U8037 (N_8037,N_7846,N_7902);
xnor U8038 (N_8038,N_7820,N_7768);
nor U8039 (N_8039,N_7880,N_7758);
nand U8040 (N_8040,N_7863,N_7976);
or U8041 (N_8041,N_7895,N_7930);
and U8042 (N_8042,N_7926,N_7770);
xor U8043 (N_8043,N_7818,N_7842);
nand U8044 (N_8044,N_7805,N_7942);
nand U8045 (N_8045,N_7803,N_7924);
nor U8046 (N_8046,N_7824,N_7951);
nand U8047 (N_8047,N_7953,N_7775);
and U8048 (N_8048,N_7970,N_7754);
nor U8049 (N_8049,N_7934,N_7799);
or U8050 (N_8050,N_7789,N_7750);
nor U8051 (N_8051,N_7907,N_7860);
and U8052 (N_8052,N_7986,N_7994);
and U8053 (N_8053,N_7990,N_7792);
or U8054 (N_8054,N_7925,N_7762);
nor U8055 (N_8055,N_7849,N_7920);
nor U8056 (N_8056,N_7753,N_7922);
or U8057 (N_8057,N_7831,N_7773);
or U8058 (N_8058,N_7944,N_7810);
or U8059 (N_8059,N_7866,N_7856);
xnor U8060 (N_8060,N_7779,N_7837);
or U8061 (N_8061,N_7802,N_7840);
and U8062 (N_8062,N_7949,N_7872);
and U8063 (N_8063,N_7988,N_7911);
nor U8064 (N_8064,N_7892,N_7777);
nand U8065 (N_8065,N_7997,N_7841);
and U8066 (N_8066,N_7958,N_7910);
xor U8067 (N_8067,N_7862,N_7967);
nor U8068 (N_8068,N_7966,N_7859);
nand U8069 (N_8069,N_7828,N_7776);
and U8070 (N_8070,N_7960,N_7875);
nand U8071 (N_8071,N_7917,N_7931);
nand U8072 (N_8072,N_7947,N_7905);
nand U8073 (N_8073,N_7903,N_7879);
nand U8074 (N_8074,N_7897,N_7937);
nand U8075 (N_8075,N_7932,N_7890);
or U8076 (N_8076,N_7778,N_7807);
nor U8077 (N_8077,N_7834,N_7817);
or U8078 (N_8078,N_7836,N_7977);
and U8079 (N_8079,N_7785,N_7882);
nor U8080 (N_8080,N_7801,N_7833);
xor U8081 (N_8081,N_7864,N_7825);
xnor U8082 (N_8082,N_7889,N_7855);
and U8083 (N_8083,N_7780,N_7782);
or U8084 (N_8084,N_7996,N_7948);
nor U8085 (N_8085,N_7781,N_7826);
and U8086 (N_8086,N_7822,N_7896);
nor U8087 (N_8087,N_7835,N_7985);
nor U8088 (N_8088,N_7906,N_7914);
and U8089 (N_8089,N_7819,N_7795);
nor U8090 (N_8090,N_7788,N_7946);
or U8091 (N_8091,N_7858,N_7893);
nand U8092 (N_8092,N_7916,N_7956);
nand U8093 (N_8093,N_7786,N_7816);
or U8094 (N_8094,N_7984,N_7929);
xnor U8095 (N_8095,N_7980,N_7854);
nand U8096 (N_8096,N_7850,N_7923);
xor U8097 (N_8097,N_7794,N_7765);
nand U8098 (N_8098,N_7983,N_7878);
or U8099 (N_8099,N_7928,N_7867);
nor U8100 (N_8100,N_7904,N_7861);
or U8101 (N_8101,N_7756,N_7852);
and U8102 (N_8102,N_7827,N_7927);
xor U8103 (N_8103,N_7962,N_7809);
and U8104 (N_8104,N_7919,N_7981);
or U8105 (N_8105,N_7783,N_7857);
nor U8106 (N_8106,N_7806,N_7808);
and U8107 (N_8107,N_7870,N_7991);
or U8108 (N_8108,N_7881,N_7797);
xor U8109 (N_8109,N_7759,N_7868);
nand U8110 (N_8110,N_7751,N_7812);
or U8111 (N_8111,N_7943,N_7999);
nand U8112 (N_8112,N_7883,N_7918);
xnor U8113 (N_8113,N_7830,N_7915);
and U8114 (N_8114,N_7774,N_7790);
nand U8115 (N_8115,N_7887,N_7950);
or U8116 (N_8116,N_7936,N_7955);
nor U8117 (N_8117,N_7853,N_7938);
or U8118 (N_8118,N_7784,N_7989);
and U8119 (N_8119,N_7913,N_7979);
nand U8120 (N_8120,N_7969,N_7877);
or U8121 (N_8121,N_7832,N_7813);
nor U8122 (N_8122,N_7763,N_7891);
and U8123 (N_8123,N_7995,N_7971);
or U8124 (N_8124,N_7978,N_7964);
or U8125 (N_8125,N_7765,N_7788);
and U8126 (N_8126,N_7989,N_7778);
and U8127 (N_8127,N_7902,N_7816);
xor U8128 (N_8128,N_7960,N_7809);
nor U8129 (N_8129,N_7829,N_7810);
xnor U8130 (N_8130,N_7914,N_7780);
nand U8131 (N_8131,N_7797,N_7851);
xnor U8132 (N_8132,N_7956,N_7810);
nand U8133 (N_8133,N_7804,N_7780);
and U8134 (N_8134,N_7847,N_7958);
and U8135 (N_8135,N_7929,N_7811);
nand U8136 (N_8136,N_7823,N_7795);
or U8137 (N_8137,N_7915,N_7814);
xor U8138 (N_8138,N_7948,N_7902);
nand U8139 (N_8139,N_7820,N_7798);
nor U8140 (N_8140,N_7850,N_7977);
and U8141 (N_8141,N_7996,N_7994);
xnor U8142 (N_8142,N_7934,N_7936);
and U8143 (N_8143,N_7810,N_7754);
nand U8144 (N_8144,N_7827,N_7823);
nand U8145 (N_8145,N_7780,N_7763);
xnor U8146 (N_8146,N_7936,N_7769);
nand U8147 (N_8147,N_7927,N_7892);
nand U8148 (N_8148,N_7864,N_7986);
or U8149 (N_8149,N_7773,N_7842);
and U8150 (N_8150,N_7828,N_7829);
xor U8151 (N_8151,N_7982,N_7780);
nand U8152 (N_8152,N_7896,N_7866);
xnor U8153 (N_8153,N_7889,N_7856);
or U8154 (N_8154,N_7764,N_7945);
nor U8155 (N_8155,N_7753,N_7791);
or U8156 (N_8156,N_7980,N_7888);
xnor U8157 (N_8157,N_7979,N_7999);
and U8158 (N_8158,N_7886,N_7910);
nand U8159 (N_8159,N_7969,N_7902);
xnor U8160 (N_8160,N_7900,N_7775);
xnor U8161 (N_8161,N_7838,N_7886);
xor U8162 (N_8162,N_7915,N_7993);
and U8163 (N_8163,N_7927,N_7877);
xnor U8164 (N_8164,N_7847,N_7903);
nand U8165 (N_8165,N_7828,N_7944);
nand U8166 (N_8166,N_7940,N_7983);
xnor U8167 (N_8167,N_7793,N_7751);
nor U8168 (N_8168,N_7781,N_7854);
and U8169 (N_8169,N_7810,N_7974);
nor U8170 (N_8170,N_7861,N_7984);
nor U8171 (N_8171,N_7924,N_7940);
nand U8172 (N_8172,N_7794,N_7879);
nand U8173 (N_8173,N_7903,N_7819);
xor U8174 (N_8174,N_7776,N_7762);
or U8175 (N_8175,N_7833,N_7962);
or U8176 (N_8176,N_7799,N_7760);
nand U8177 (N_8177,N_7786,N_7858);
xnor U8178 (N_8178,N_7966,N_7980);
or U8179 (N_8179,N_7785,N_7918);
nor U8180 (N_8180,N_7952,N_7891);
or U8181 (N_8181,N_7793,N_7755);
and U8182 (N_8182,N_7921,N_7766);
or U8183 (N_8183,N_7842,N_7925);
xnor U8184 (N_8184,N_7832,N_7779);
xnor U8185 (N_8185,N_7892,N_7907);
nand U8186 (N_8186,N_7867,N_7812);
nand U8187 (N_8187,N_7865,N_7789);
xnor U8188 (N_8188,N_7808,N_7789);
xnor U8189 (N_8189,N_7905,N_7798);
nand U8190 (N_8190,N_7855,N_7944);
and U8191 (N_8191,N_7800,N_7935);
and U8192 (N_8192,N_7891,N_7947);
nor U8193 (N_8193,N_7931,N_7921);
xor U8194 (N_8194,N_7760,N_7781);
or U8195 (N_8195,N_7849,N_7798);
and U8196 (N_8196,N_7906,N_7842);
xnor U8197 (N_8197,N_7842,N_7935);
or U8198 (N_8198,N_7765,N_7978);
nand U8199 (N_8199,N_7814,N_7868);
nor U8200 (N_8200,N_7792,N_7970);
or U8201 (N_8201,N_7802,N_7896);
nand U8202 (N_8202,N_7889,N_7849);
and U8203 (N_8203,N_7774,N_7870);
nor U8204 (N_8204,N_7909,N_7750);
and U8205 (N_8205,N_7904,N_7930);
xor U8206 (N_8206,N_7888,N_7929);
nor U8207 (N_8207,N_7783,N_7822);
nor U8208 (N_8208,N_7751,N_7754);
xor U8209 (N_8209,N_7921,N_7882);
or U8210 (N_8210,N_7813,N_7857);
xor U8211 (N_8211,N_7937,N_7875);
xor U8212 (N_8212,N_7946,N_7813);
and U8213 (N_8213,N_7979,N_7965);
or U8214 (N_8214,N_7877,N_7865);
nor U8215 (N_8215,N_7830,N_7798);
and U8216 (N_8216,N_7794,N_7833);
or U8217 (N_8217,N_7853,N_7842);
or U8218 (N_8218,N_7841,N_7943);
xor U8219 (N_8219,N_7787,N_7767);
or U8220 (N_8220,N_7804,N_7875);
or U8221 (N_8221,N_7769,N_7792);
xor U8222 (N_8222,N_7938,N_7888);
nor U8223 (N_8223,N_7911,N_7792);
nor U8224 (N_8224,N_7864,N_7835);
and U8225 (N_8225,N_7995,N_7939);
or U8226 (N_8226,N_7887,N_7866);
and U8227 (N_8227,N_7772,N_7975);
nor U8228 (N_8228,N_7795,N_7836);
nand U8229 (N_8229,N_7915,N_7935);
and U8230 (N_8230,N_7896,N_7849);
and U8231 (N_8231,N_7892,N_7870);
nor U8232 (N_8232,N_7751,N_7957);
or U8233 (N_8233,N_7977,N_7901);
nor U8234 (N_8234,N_7997,N_7759);
nand U8235 (N_8235,N_7904,N_7889);
or U8236 (N_8236,N_7977,N_7796);
or U8237 (N_8237,N_7887,N_7932);
or U8238 (N_8238,N_7938,N_7816);
nor U8239 (N_8239,N_7897,N_7752);
or U8240 (N_8240,N_7937,N_7826);
nand U8241 (N_8241,N_7955,N_7987);
xor U8242 (N_8242,N_7766,N_7822);
and U8243 (N_8243,N_7860,N_7763);
nor U8244 (N_8244,N_7761,N_7827);
nand U8245 (N_8245,N_7863,N_7908);
nand U8246 (N_8246,N_7942,N_7956);
xor U8247 (N_8247,N_7948,N_7832);
nor U8248 (N_8248,N_7877,N_7777);
nand U8249 (N_8249,N_7903,N_7887);
nor U8250 (N_8250,N_8017,N_8098);
nand U8251 (N_8251,N_8195,N_8021);
nand U8252 (N_8252,N_8114,N_8176);
nand U8253 (N_8253,N_8192,N_8145);
xor U8254 (N_8254,N_8088,N_8008);
and U8255 (N_8255,N_8031,N_8148);
and U8256 (N_8256,N_8188,N_8082);
and U8257 (N_8257,N_8045,N_8181);
or U8258 (N_8258,N_8220,N_8249);
nand U8259 (N_8259,N_8240,N_8113);
nand U8260 (N_8260,N_8222,N_8172);
nand U8261 (N_8261,N_8058,N_8047);
and U8262 (N_8262,N_8175,N_8206);
or U8263 (N_8263,N_8140,N_8080);
nor U8264 (N_8264,N_8146,N_8104);
xnor U8265 (N_8265,N_8030,N_8081);
xor U8266 (N_8266,N_8018,N_8120);
nor U8267 (N_8267,N_8089,N_8214);
and U8268 (N_8268,N_8090,N_8044);
nor U8269 (N_8269,N_8035,N_8116);
nand U8270 (N_8270,N_8213,N_8194);
nand U8271 (N_8271,N_8007,N_8121);
nor U8272 (N_8272,N_8155,N_8205);
xor U8273 (N_8273,N_8247,N_8037);
and U8274 (N_8274,N_8233,N_8078);
xnor U8275 (N_8275,N_8009,N_8006);
and U8276 (N_8276,N_8052,N_8144);
xnor U8277 (N_8277,N_8199,N_8135);
nor U8278 (N_8278,N_8087,N_8010);
nand U8279 (N_8279,N_8042,N_8019);
and U8280 (N_8280,N_8190,N_8202);
or U8281 (N_8281,N_8132,N_8131);
nand U8282 (N_8282,N_8151,N_8211);
or U8283 (N_8283,N_8083,N_8150);
nor U8284 (N_8284,N_8112,N_8138);
nor U8285 (N_8285,N_8160,N_8126);
xnor U8286 (N_8286,N_8022,N_8029);
nand U8287 (N_8287,N_8062,N_8077);
and U8288 (N_8288,N_8165,N_8033);
nand U8289 (N_8289,N_8095,N_8034);
nand U8290 (N_8290,N_8170,N_8149);
or U8291 (N_8291,N_8073,N_8003);
nor U8292 (N_8292,N_8106,N_8187);
and U8293 (N_8293,N_8005,N_8036);
and U8294 (N_8294,N_8056,N_8166);
xor U8295 (N_8295,N_8232,N_8183);
and U8296 (N_8296,N_8248,N_8065);
or U8297 (N_8297,N_8173,N_8158);
xnor U8298 (N_8298,N_8063,N_8096);
or U8299 (N_8299,N_8200,N_8171);
or U8300 (N_8300,N_8244,N_8004);
or U8301 (N_8301,N_8105,N_8099);
nor U8302 (N_8302,N_8204,N_8013);
or U8303 (N_8303,N_8178,N_8002);
and U8304 (N_8304,N_8152,N_8084);
or U8305 (N_8305,N_8075,N_8050);
nand U8306 (N_8306,N_8147,N_8108);
nand U8307 (N_8307,N_8234,N_8027);
nand U8308 (N_8308,N_8012,N_8246);
xor U8309 (N_8309,N_8111,N_8209);
nor U8310 (N_8310,N_8119,N_8127);
nor U8311 (N_8311,N_8094,N_8102);
xor U8312 (N_8312,N_8226,N_8086);
nand U8313 (N_8313,N_8103,N_8016);
and U8314 (N_8314,N_8215,N_8227);
nand U8315 (N_8315,N_8186,N_8193);
nor U8316 (N_8316,N_8101,N_8011);
and U8317 (N_8317,N_8085,N_8000);
nand U8318 (N_8318,N_8168,N_8137);
nand U8319 (N_8319,N_8129,N_8225);
nor U8320 (N_8320,N_8242,N_8141);
and U8321 (N_8321,N_8185,N_8048);
and U8322 (N_8322,N_8040,N_8230);
or U8323 (N_8323,N_8218,N_8208);
or U8324 (N_8324,N_8219,N_8071);
xor U8325 (N_8325,N_8241,N_8072);
nor U8326 (N_8326,N_8142,N_8097);
nand U8327 (N_8327,N_8217,N_8153);
and U8328 (N_8328,N_8053,N_8051);
and U8329 (N_8329,N_8196,N_8212);
nor U8330 (N_8330,N_8117,N_8032);
nor U8331 (N_8331,N_8161,N_8107);
nor U8332 (N_8332,N_8068,N_8091);
xor U8333 (N_8333,N_8189,N_8059);
xnor U8334 (N_8334,N_8046,N_8038);
and U8335 (N_8335,N_8197,N_8136);
and U8336 (N_8336,N_8159,N_8224);
or U8337 (N_8337,N_8025,N_8066);
nand U8338 (N_8338,N_8154,N_8015);
or U8339 (N_8339,N_8239,N_8169);
nor U8340 (N_8340,N_8014,N_8115);
nor U8341 (N_8341,N_8236,N_8133);
nor U8342 (N_8342,N_8054,N_8203);
xnor U8343 (N_8343,N_8180,N_8070);
or U8344 (N_8344,N_8049,N_8143);
or U8345 (N_8345,N_8243,N_8079);
or U8346 (N_8346,N_8238,N_8067);
or U8347 (N_8347,N_8060,N_8057);
xor U8348 (N_8348,N_8164,N_8020);
nor U8349 (N_8349,N_8061,N_8109);
or U8350 (N_8350,N_8100,N_8064);
nor U8351 (N_8351,N_8229,N_8167);
or U8352 (N_8352,N_8039,N_8231);
or U8353 (N_8353,N_8125,N_8179);
xor U8354 (N_8354,N_8069,N_8162);
nand U8355 (N_8355,N_8023,N_8174);
xor U8356 (N_8356,N_8139,N_8184);
nand U8357 (N_8357,N_8055,N_8182);
nor U8358 (N_8358,N_8092,N_8123);
nor U8359 (N_8359,N_8216,N_8245);
or U8360 (N_8360,N_8041,N_8093);
xnor U8361 (N_8361,N_8026,N_8130);
nor U8362 (N_8362,N_8076,N_8177);
nor U8363 (N_8363,N_8118,N_8028);
nand U8364 (N_8364,N_8198,N_8201);
or U8365 (N_8365,N_8221,N_8228);
and U8366 (N_8366,N_8163,N_8001);
nand U8367 (N_8367,N_8134,N_8191);
and U8368 (N_8368,N_8157,N_8235);
and U8369 (N_8369,N_8110,N_8207);
and U8370 (N_8370,N_8156,N_8210);
or U8371 (N_8371,N_8124,N_8024);
nor U8372 (N_8372,N_8074,N_8122);
nand U8373 (N_8373,N_8128,N_8237);
nor U8374 (N_8374,N_8223,N_8043);
xor U8375 (N_8375,N_8128,N_8110);
nand U8376 (N_8376,N_8197,N_8031);
and U8377 (N_8377,N_8033,N_8197);
or U8378 (N_8378,N_8184,N_8040);
or U8379 (N_8379,N_8082,N_8143);
nand U8380 (N_8380,N_8208,N_8071);
xor U8381 (N_8381,N_8131,N_8015);
xnor U8382 (N_8382,N_8218,N_8146);
xor U8383 (N_8383,N_8203,N_8248);
or U8384 (N_8384,N_8168,N_8077);
or U8385 (N_8385,N_8063,N_8205);
and U8386 (N_8386,N_8177,N_8228);
xor U8387 (N_8387,N_8199,N_8224);
or U8388 (N_8388,N_8027,N_8204);
nor U8389 (N_8389,N_8123,N_8094);
nand U8390 (N_8390,N_8228,N_8042);
nand U8391 (N_8391,N_8140,N_8095);
or U8392 (N_8392,N_8228,N_8038);
xor U8393 (N_8393,N_8007,N_8112);
xnor U8394 (N_8394,N_8047,N_8097);
and U8395 (N_8395,N_8170,N_8039);
or U8396 (N_8396,N_8095,N_8209);
xnor U8397 (N_8397,N_8155,N_8249);
nor U8398 (N_8398,N_8100,N_8197);
nand U8399 (N_8399,N_8099,N_8147);
and U8400 (N_8400,N_8190,N_8088);
and U8401 (N_8401,N_8200,N_8022);
or U8402 (N_8402,N_8129,N_8034);
nor U8403 (N_8403,N_8121,N_8192);
nor U8404 (N_8404,N_8128,N_8191);
nor U8405 (N_8405,N_8111,N_8104);
nand U8406 (N_8406,N_8093,N_8117);
and U8407 (N_8407,N_8229,N_8060);
or U8408 (N_8408,N_8093,N_8243);
and U8409 (N_8409,N_8061,N_8131);
nand U8410 (N_8410,N_8124,N_8201);
nor U8411 (N_8411,N_8238,N_8181);
nand U8412 (N_8412,N_8239,N_8182);
and U8413 (N_8413,N_8243,N_8130);
and U8414 (N_8414,N_8141,N_8004);
and U8415 (N_8415,N_8056,N_8004);
nor U8416 (N_8416,N_8061,N_8091);
and U8417 (N_8417,N_8112,N_8175);
nand U8418 (N_8418,N_8122,N_8061);
nand U8419 (N_8419,N_8143,N_8117);
and U8420 (N_8420,N_8246,N_8143);
xnor U8421 (N_8421,N_8029,N_8202);
or U8422 (N_8422,N_8054,N_8223);
nor U8423 (N_8423,N_8091,N_8234);
nand U8424 (N_8424,N_8201,N_8244);
and U8425 (N_8425,N_8126,N_8120);
xnor U8426 (N_8426,N_8128,N_8095);
or U8427 (N_8427,N_8189,N_8090);
xor U8428 (N_8428,N_8005,N_8201);
or U8429 (N_8429,N_8088,N_8191);
and U8430 (N_8430,N_8035,N_8090);
nor U8431 (N_8431,N_8174,N_8147);
xnor U8432 (N_8432,N_8229,N_8105);
xor U8433 (N_8433,N_8092,N_8186);
nor U8434 (N_8434,N_8229,N_8074);
nor U8435 (N_8435,N_8123,N_8041);
nor U8436 (N_8436,N_8177,N_8097);
nor U8437 (N_8437,N_8075,N_8240);
nand U8438 (N_8438,N_8153,N_8209);
xnor U8439 (N_8439,N_8005,N_8177);
xor U8440 (N_8440,N_8248,N_8185);
or U8441 (N_8441,N_8139,N_8193);
or U8442 (N_8442,N_8050,N_8096);
and U8443 (N_8443,N_8151,N_8214);
and U8444 (N_8444,N_8147,N_8123);
nor U8445 (N_8445,N_8091,N_8064);
and U8446 (N_8446,N_8088,N_8206);
nand U8447 (N_8447,N_8189,N_8220);
nand U8448 (N_8448,N_8210,N_8058);
nand U8449 (N_8449,N_8137,N_8013);
or U8450 (N_8450,N_8095,N_8196);
xnor U8451 (N_8451,N_8190,N_8011);
nand U8452 (N_8452,N_8246,N_8112);
nand U8453 (N_8453,N_8008,N_8133);
and U8454 (N_8454,N_8000,N_8240);
nand U8455 (N_8455,N_8047,N_8223);
xnor U8456 (N_8456,N_8237,N_8170);
nor U8457 (N_8457,N_8094,N_8168);
and U8458 (N_8458,N_8069,N_8075);
or U8459 (N_8459,N_8231,N_8155);
and U8460 (N_8460,N_8065,N_8140);
nand U8461 (N_8461,N_8166,N_8184);
and U8462 (N_8462,N_8051,N_8093);
nor U8463 (N_8463,N_8166,N_8010);
nor U8464 (N_8464,N_8235,N_8082);
and U8465 (N_8465,N_8170,N_8183);
xnor U8466 (N_8466,N_8158,N_8243);
and U8467 (N_8467,N_8035,N_8061);
nor U8468 (N_8468,N_8173,N_8196);
nor U8469 (N_8469,N_8224,N_8193);
or U8470 (N_8470,N_8232,N_8090);
xor U8471 (N_8471,N_8009,N_8200);
xor U8472 (N_8472,N_8009,N_8120);
nor U8473 (N_8473,N_8190,N_8182);
nand U8474 (N_8474,N_8090,N_8101);
nor U8475 (N_8475,N_8019,N_8183);
or U8476 (N_8476,N_8237,N_8038);
and U8477 (N_8477,N_8050,N_8015);
nand U8478 (N_8478,N_8139,N_8099);
nor U8479 (N_8479,N_8064,N_8202);
or U8480 (N_8480,N_8111,N_8210);
xnor U8481 (N_8481,N_8114,N_8038);
xor U8482 (N_8482,N_8150,N_8140);
nor U8483 (N_8483,N_8248,N_8115);
nor U8484 (N_8484,N_8218,N_8187);
or U8485 (N_8485,N_8072,N_8249);
or U8486 (N_8486,N_8232,N_8010);
xnor U8487 (N_8487,N_8050,N_8049);
and U8488 (N_8488,N_8082,N_8228);
xnor U8489 (N_8489,N_8152,N_8112);
xor U8490 (N_8490,N_8130,N_8197);
and U8491 (N_8491,N_8247,N_8079);
and U8492 (N_8492,N_8236,N_8178);
and U8493 (N_8493,N_8009,N_8077);
nor U8494 (N_8494,N_8006,N_8054);
xor U8495 (N_8495,N_8088,N_8201);
xor U8496 (N_8496,N_8076,N_8225);
nand U8497 (N_8497,N_8233,N_8186);
nor U8498 (N_8498,N_8092,N_8034);
or U8499 (N_8499,N_8044,N_8119);
nand U8500 (N_8500,N_8425,N_8431);
xnor U8501 (N_8501,N_8477,N_8411);
nand U8502 (N_8502,N_8288,N_8344);
or U8503 (N_8503,N_8394,N_8383);
and U8504 (N_8504,N_8480,N_8490);
or U8505 (N_8505,N_8389,N_8290);
or U8506 (N_8506,N_8282,N_8315);
and U8507 (N_8507,N_8427,N_8261);
nor U8508 (N_8508,N_8271,N_8355);
xor U8509 (N_8509,N_8348,N_8436);
nor U8510 (N_8510,N_8316,N_8292);
and U8511 (N_8511,N_8255,N_8435);
nand U8512 (N_8512,N_8281,N_8373);
and U8513 (N_8513,N_8350,N_8371);
xnor U8514 (N_8514,N_8446,N_8467);
or U8515 (N_8515,N_8317,N_8474);
xor U8516 (N_8516,N_8415,N_8481);
and U8517 (N_8517,N_8289,N_8485);
nand U8518 (N_8518,N_8302,N_8341);
and U8519 (N_8519,N_8252,N_8268);
xnor U8520 (N_8520,N_8295,N_8449);
nor U8521 (N_8521,N_8484,N_8280);
or U8522 (N_8522,N_8378,N_8346);
and U8523 (N_8523,N_8418,N_8419);
or U8524 (N_8524,N_8463,N_8479);
and U8525 (N_8525,N_8256,N_8420);
or U8526 (N_8526,N_8486,N_8366);
nor U8527 (N_8527,N_8382,N_8258);
and U8528 (N_8528,N_8438,N_8307);
or U8529 (N_8529,N_8487,N_8364);
xnor U8530 (N_8530,N_8254,N_8381);
or U8531 (N_8531,N_8426,N_8262);
and U8532 (N_8532,N_8417,N_8314);
nor U8533 (N_8533,N_8319,N_8454);
and U8534 (N_8534,N_8489,N_8329);
xnor U8535 (N_8535,N_8343,N_8468);
nand U8536 (N_8536,N_8345,N_8422);
xor U8537 (N_8537,N_8321,N_8465);
or U8538 (N_8538,N_8392,N_8395);
xnor U8539 (N_8539,N_8380,N_8396);
or U8540 (N_8540,N_8325,N_8328);
nand U8541 (N_8541,N_8372,N_8340);
xor U8542 (N_8542,N_8305,N_8297);
nand U8543 (N_8543,N_8267,N_8464);
nand U8544 (N_8544,N_8452,N_8284);
nor U8545 (N_8545,N_8461,N_8301);
or U8546 (N_8546,N_8483,N_8457);
nor U8547 (N_8547,N_8401,N_8351);
and U8548 (N_8548,N_8407,N_8400);
nor U8549 (N_8549,N_8403,N_8264);
and U8550 (N_8550,N_8434,N_8398);
or U8551 (N_8551,N_8270,N_8306);
and U8552 (N_8552,N_8499,N_8361);
or U8553 (N_8553,N_8349,N_8478);
xor U8554 (N_8554,N_8260,N_8354);
nor U8555 (N_8555,N_8429,N_8326);
nand U8556 (N_8556,N_8450,N_8253);
nand U8557 (N_8557,N_8387,N_8285);
nor U8558 (N_8558,N_8496,N_8250);
xnor U8559 (N_8559,N_8384,N_8416);
nand U8560 (N_8560,N_8304,N_8405);
nand U8561 (N_8561,N_8488,N_8455);
and U8562 (N_8562,N_8421,N_8441);
nor U8563 (N_8563,N_8330,N_8327);
xor U8564 (N_8564,N_8347,N_8462);
nand U8565 (N_8565,N_8363,N_8437);
nand U8566 (N_8566,N_8296,N_8473);
xor U8567 (N_8567,N_8283,N_8494);
nand U8568 (N_8568,N_8265,N_8375);
and U8569 (N_8569,N_8369,N_8412);
nor U8570 (N_8570,N_8370,N_8287);
and U8571 (N_8571,N_8495,N_8424);
nor U8572 (N_8572,N_8311,N_8413);
nand U8573 (N_8573,N_8498,N_8472);
or U8574 (N_8574,N_8274,N_8353);
and U8575 (N_8575,N_8277,N_8456);
and U8576 (N_8576,N_8377,N_8460);
nand U8577 (N_8577,N_8337,N_8263);
and U8578 (N_8578,N_8493,N_8322);
xnor U8579 (N_8579,N_8294,N_8433);
or U8580 (N_8580,N_8356,N_8333);
nand U8581 (N_8581,N_8410,N_8313);
nand U8582 (N_8582,N_8497,N_8393);
or U8583 (N_8583,N_8338,N_8273);
xor U8584 (N_8584,N_8357,N_8443);
xnor U8585 (N_8585,N_8445,N_8299);
or U8586 (N_8586,N_8332,N_8358);
nor U8587 (N_8587,N_8459,N_8342);
and U8588 (N_8588,N_8323,N_8439);
xnor U8589 (N_8589,N_8453,N_8286);
and U8590 (N_8590,N_8430,N_8428);
xnor U8591 (N_8591,N_8298,N_8276);
nor U8592 (N_8592,N_8444,N_8404);
and U8593 (N_8593,N_8336,N_8269);
xnor U8594 (N_8594,N_8259,N_8408);
xor U8595 (N_8595,N_8476,N_8324);
and U8596 (N_8596,N_8492,N_8335);
or U8597 (N_8597,N_8339,N_8471);
or U8598 (N_8598,N_8458,N_8385);
nor U8599 (N_8599,N_8308,N_8448);
xor U8600 (N_8600,N_8368,N_8352);
or U8601 (N_8601,N_8409,N_8379);
nand U8602 (N_8602,N_8318,N_8251);
and U8603 (N_8603,N_8334,N_8278);
xnor U8604 (N_8604,N_8482,N_8470);
xnor U8605 (N_8605,N_8275,N_8367);
and U8606 (N_8606,N_8440,N_8442);
nor U8607 (N_8607,N_8399,N_8257);
or U8608 (N_8608,N_8320,N_8272);
nor U8609 (N_8609,N_8376,N_8447);
nor U8610 (N_8610,N_8397,N_8374);
or U8611 (N_8611,N_8475,N_8365);
nand U8612 (N_8612,N_8359,N_8266);
and U8613 (N_8613,N_8390,N_8331);
and U8614 (N_8614,N_8310,N_8391);
and U8615 (N_8615,N_8279,N_8300);
and U8616 (N_8616,N_8388,N_8312);
nor U8617 (N_8617,N_8303,N_8466);
xor U8618 (N_8618,N_8491,N_8386);
nor U8619 (N_8619,N_8423,N_8360);
or U8620 (N_8620,N_8291,N_8309);
nor U8621 (N_8621,N_8469,N_8293);
xnor U8622 (N_8622,N_8362,N_8402);
nand U8623 (N_8623,N_8414,N_8432);
or U8624 (N_8624,N_8406,N_8451);
xnor U8625 (N_8625,N_8426,N_8357);
and U8626 (N_8626,N_8421,N_8454);
or U8627 (N_8627,N_8485,N_8446);
nand U8628 (N_8628,N_8366,N_8376);
nand U8629 (N_8629,N_8384,N_8394);
nor U8630 (N_8630,N_8405,N_8443);
nor U8631 (N_8631,N_8355,N_8454);
and U8632 (N_8632,N_8367,N_8475);
nand U8633 (N_8633,N_8421,N_8273);
or U8634 (N_8634,N_8487,N_8415);
and U8635 (N_8635,N_8321,N_8337);
or U8636 (N_8636,N_8352,N_8433);
and U8637 (N_8637,N_8321,N_8258);
and U8638 (N_8638,N_8282,N_8294);
and U8639 (N_8639,N_8427,N_8295);
or U8640 (N_8640,N_8406,N_8301);
nor U8641 (N_8641,N_8310,N_8497);
and U8642 (N_8642,N_8432,N_8451);
and U8643 (N_8643,N_8487,N_8485);
nand U8644 (N_8644,N_8399,N_8458);
or U8645 (N_8645,N_8321,N_8429);
xnor U8646 (N_8646,N_8283,N_8464);
nor U8647 (N_8647,N_8411,N_8442);
nor U8648 (N_8648,N_8367,N_8428);
or U8649 (N_8649,N_8356,N_8290);
nor U8650 (N_8650,N_8327,N_8412);
and U8651 (N_8651,N_8424,N_8260);
and U8652 (N_8652,N_8325,N_8395);
nand U8653 (N_8653,N_8279,N_8369);
and U8654 (N_8654,N_8391,N_8404);
nand U8655 (N_8655,N_8348,N_8320);
or U8656 (N_8656,N_8311,N_8380);
and U8657 (N_8657,N_8449,N_8338);
nand U8658 (N_8658,N_8484,N_8325);
nor U8659 (N_8659,N_8344,N_8306);
or U8660 (N_8660,N_8292,N_8471);
nor U8661 (N_8661,N_8418,N_8399);
xor U8662 (N_8662,N_8294,N_8471);
nor U8663 (N_8663,N_8385,N_8287);
nor U8664 (N_8664,N_8324,N_8266);
nand U8665 (N_8665,N_8480,N_8422);
and U8666 (N_8666,N_8282,N_8384);
nor U8667 (N_8667,N_8478,N_8326);
nor U8668 (N_8668,N_8359,N_8284);
and U8669 (N_8669,N_8318,N_8314);
or U8670 (N_8670,N_8265,N_8430);
nor U8671 (N_8671,N_8435,N_8286);
nor U8672 (N_8672,N_8370,N_8454);
nor U8673 (N_8673,N_8384,N_8420);
or U8674 (N_8674,N_8451,N_8314);
xnor U8675 (N_8675,N_8388,N_8255);
or U8676 (N_8676,N_8363,N_8398);
nand U8677 (N_8677,N_8409,N_8328);
xor U8678 (N_8678,N_8422,N_8275);
xnor U8679 (N_8679,N_8344,N_8285);
nor U8680 (N_8680,N_8299,N_8319);
nor U8681 (N_8681,N_8339,N_8448);
xor U8682 (N_8682,N_8344,N_8293);
nand U8683 (N_8683,N_8452,N_8411);
or U8684 (N_8684,N_8449,N_8329);
xor U8685 (N_8685,N_8337,N_8376);
nor U8686 (N_8686,N_8267,N_8381);
nor U8687 (N_8687,N_8499,N_8283);
nand U8688 (N_8688,N_8462,N_8468);
and U8689 (N_8689,N_8428,N_8301);
or U8690 (N_8690,N_8257,N_8276);
xor U8691 (N_8691,N_8457,N_8356);
and U8692 (N_8692,N_8390,N_8275);
nand U8693 (N_8693,N_8384,N_8342);
and U8694 (N_8694,N_8254,N_8469);
nor U8695 (N_8695,N_8275,N_8451);
and U8696 (N_8696,N_8397,N_8492);
xor U8697 (N_8697,N_8422,N_8321);
nor U8698 (N_8698,N_8377,N_8367);
and U8699 (N_8699,N_8280,N_8276);
xnor U8700 (N_8700,N_8262,N_8381);
nand U8701 (N_8701,N_8312,N_8349);
nand U8702 (N_8702,N_8494,N_8326);
and U8703 (N_8703,N_8490,N_8383);
and U8704 (N_8704,N_8274,N_8415);
nand U8705 (N_8705,N_8308,N_8354);
or U8706 (N_8706,N_8347,N_8374);
and U8707 (N_8707,N_8290,N_8336);
xnor U8708 (N_8708,N_8310,N_8415);
xor U8709 (N_8709,N_8313,N_8390);
and U8710 (N_8710,N_8491,N_8364);
nor U8711 (N_8711,N_8382,N_8368);
nand U8712 (N_8712,N_8394,N_8321);
xor U8713 (N_8713,N_8482,N_8313);
or U8714 (N_8714,N_8357,N_8250);
xor U8715 (N_8715,N_8304,N_8296);
nor U8716 (N_8716,N_8416,N_8423);
and U8717 (N_8717,N_8333,N_8341);
nand U8718 (N_8718,N_8268,N_8449);
or U8719 (N_8719,N_8487,N_8351);
and U8720 (N_8720,N_8317,N_8258);
nand U8721 (N_8721,N_8289,N_8407);
nor U8722 (N_8722,N_8354,N_8346);
nand U8723 (N_8723,N_8447,N_8387);
and U8724 (N_8724,N_8300,N_8362);
and U8725 (N_8725,N_8338,N_8355);
or U8726 (N_8726,N_8252,N_8395);
nand U8727 (N_8727,N_8265,N_8318);
nand U8728 (N_8728,N_8353,N_8332);
xor U8729 (N_8729,N_8302,N_8434);
or U8730 (N_8730,N_8319,N_8406);
and U8731 (N_8731,N_8460,N_8311);
and U8732 (N_8732,N_8445,N_8439);
xnor U8733 (N_8733,N_8409,N_8422);
nor U8734 (N_8734,N_8482,N_8368);
nor U8735 (N_8735,N_8309,N_8348);
and U8736 (N_8736,N_8322,N_8286);
and U8737 (N_8737,N_8360,N_8291);
or U8738 (N_8738,N_8303,N_8492);
xor U8739 (N_8739,N_8266,N_8447);
nor U8740 (N_8740,N_8268,N_8313);
nand U8741 (N_8741,N_8268,N_8461);
nand U8742 (N_8742,N_8337,N_8348);
nor U8743 (N_8743,N_8410,N_8435);
nand U8744 (N_8744,N_8436,N_8350);
and U8745 (N_8745,N_8262,N_8306);
or U8746 (N_8746,N_8449,N_8481);
and U8747 (N_8747,N_8468,N_8395);
or U8748 (N_8748,N_8329,N_8472);
nor U8749 (N_8749,N_8371,N_8388);
or U8750 (N_8750,N_8508,N_8695);
xnor U8751 (N_8751,N_8727,N_8506);
xnor U8752 (N_8752,N_8604,N_8540);
nor U8753 (N_8753,N_8574,N_8564);
xnor U8754 (N_8754,N_8669,N_8636);
nand U8755 (N_8755,N_8552,N_8624);
nand U8756 (N_8756,N_8593,N_8514);
and U8757 (N_8757,N_8516,N_8535);
nand U8758 (N_8758,N_8573,N_8545);
and U8759 (N_8759,N_8654,N_8656);
xor U8760 (N_8760,N_8575,N_8583);
nand U8761 (N_8761,N_8700,N_8725);
or U8762 (N_8762,N_8529,N_8606);
xnor U8763 (N_8763,N_8536,N_8584);
nand U8764 (N_8764,N_8722,N_8732);
xor U8765 (N_8765,N_8647,N_8663);
nand U8766 (N_8766,N_8625,N_8607);
and U8767 (N_8767,N_8561,N_8547);
or U8768 (N_8768,N_8659,N_8702);
xor U8769 (N_8769,N_8661,N_8621);
and U8770 (N_8770,N_8524,N_8719);
and U8771 (N_8771,N_8605,N_8541);
and U8772 (N_8772,N_8671,N_8664);
nor U8773 (N_8773,N_8518,N_8530);
xor U8774 (N_8774,N_8739,N_8646);
and U8775 (N_8775,N_8592,N_8628);
xnor U8776 (N_8776,N_8579,N_8511);
nand U8777 (N_8777,N_8568,N_8572);
nand U8778 (N_8778,N_8505,N_8691);
nor U8779 (N_8779,N_8692,N_8714);
nand U8780 (N_8780,N_8715,N_8509);
or U8781 (N_8781,N_8716,N_8635);
and U8782 (N_8782,N_8705,N_8675);
or U8783 (N_8783,N_8610,N_8587);
or U8784 (N_8784,N_8611,N_8595);
nand U8785 (N_8785,N_8682,N_8566);
nor U8786 (N_8786,N_8602,N_8502);
nand U8787 (N_8787,N_8737,N_8665);
nand U8788 (N_8788,N_8658,N_8687);
nand U8789 (N_8789,N_8570,N_8527);
xnor U8790 (N_8790,N_8676,N_8588);
xnor U8791 (N_8791,N_8679,N_8551);
or U8792 (N_8792,N_8614,N_8730);
or U8793 (N_8793,N_8504,N_8550);
and U8794 (N_8794,N_8603,N_8720);
xor U8795 (N_8795,N_8598,N_8642);
nor U8796 (N_8796,N_8539,N_8711);
and U8797 (N_8797,N_8630,N_8553);
nand U8798 (N_8798,N_8660,N_8620);
xnor U8799 (N_8799,N_8723,N_8688);
or U8800 (N_8800,N_8637,N_8651);
or U8801 (N_8801,N_8668,N_8670);
nand U8802 (N_8802,N_8734,N_8726);
nand U8803 (N_8803,N_8576,N_8662);
nand U8804 (N_8804,N_8645,N_8742);
nand U8805 (N_8805,N_8554,N_8699);
and U8806 (N_8806,N_8537,N_8736);
or U8807 (N_8807,N_8741,N_8608);
or U8808 (N_8808,N_8600,N_8613);
xnor U8809 (N_8809,N_8643,N_8672);
nor U8810 (N_8810,N_8743,N_8707);
or U8811 (N_8811,N_8728,N_8559);
or U8812 (N_8812,N_8589,N_8685);
xnor U8813 (N_8813,N_8717,N_8657);
xor U8814 (N_8814,N_8683,N_8693);
nor U8815 (N_8815,N_8582,N_8631);
nor U8816 (N_8816,N_8738,N_8565);
and U8817 (N_8817,N_8562,N_8681);
and U8818 (N_8818,N_8684,N_8627);
or U8819 (N_8819,N_8713,N_8617);
nor U8820 (N_8820,N_8513,N_8534);
nand U8821 (N_8821,N_8612,N_8650);
and U8822 (N_8822,N_8718,N_8525);
xor U8823 (N_8823,N_8640,N_8500);
xnor U8824 (N_8824,N_8615,N_8526);
or U8825 (N_8825,N_8735,N_8749);
or U8826 (N_8826,N_8649,N_8667);
xor U8827 (N_8827,N_8619,N_8698);
xor U8828 (N_8828,N_8706,N_8558);
and U8829 (N_8829,N_8744,N_8708);
or U8830 (N_8830,N_8548,N_8597);
or U8831 (N_8831,N_8515,N_8577);
or U8832 (N_8832,N_8510,N_8528);
and U8833 (N_8833,N_8648,N_8653);
nor U8834 (N_8834,N_8644,N_8521);
nand U8835 (N_8835,N_8520,N_8517);
or U8836 (N_8836,N_8544,N_8599);
nor U8837 (N_8837,N_8609,N_8501);
nor U8838 (N_8838,N_8542,N_8678);
xor U8839 (N_8839,N_8578,N_8622);
nand U8840 (N_8840,N_8721,N_8616);
or U8841 (N_8841,N_8686,N_8694);
and U8842 (N_8842,N_8532,N_8712);
or U8843 (N_8843,N_8503,N_8507);
nor U8844 (N_8844,N_8567,N_8632);
nand U8845 (N_8845,N_8690,N_8512);
xnor U8846 (N_8846,N_8747,N_8709);
nand U8847 (N_8847,N_8733,N_8560);
and U8848 (N_8848,N_8557,N_8666);
or U8849 (N_8849,N_8522,N_8543);
nor U8850 (N_8850,N_8549,N_8652);
xor U8851 (N_8851,N_8673,N_8563);
and U8852 (N_8852,N_8533,N_8569);
nor U8853 (N_8853,N_8586,N_8638);
nand U8854 (N_8854,N_8639,N_8519);
or U8855 (N_8855,N_8689,N_8740);
or U8856 (N_8856,N_8531,N_8680);
xor U8857 (N_8857,N_8696,N_8729);
nand U8858 (N_8858,N_8555,N_8731);
nor U8859 (N_8859,N_8591,N_8601);
or U8860 (N_8860,N_8748,N_8641);
and U8861 (N_8861,N_8745,N_8703);
and U8862 (N_8862,N_8697,N_8594);
nor U8863 (N_8863,N_8538,N_8556);
xnor U8864 (N_8864,N_8590,N_8704);
and U8865 (N_8865,N_8655,N_8623);
and U8866 (N_8866,N_8546,N_8701);
or U8867 (N_8867,N_8523,N_8585);
or U8868 (N_8868,N_8724,N_8634);
or U8869 (N_8869,N_8596,N_8626);
or U8870 (N_8870,N_8571,N_8633);
xor U8871 (N_8871,N_8677,N_8581);
or U8872 (N_8872,N_8746,N_8618);
and U8873 (N_8873,N_8580,N_8674);
nor U8874 (N_8874,N_8710,N_8629);
nand U8875 (N_8875,N_8738,N_8541);
or U8876 (N_8876,N_8716,N_8741);
and U8877 (N_8877,N_8597,N_8627);
or U8878 (N_8878,N_8668,N_8596);
nand U8879 (N_8879,N_8501,N_8544);
xnor U8880 (N_8880,N_8632,N_8578);
nor U8881 (N_8881,N_8732,N_8739);
nand U8882 (N_8882,N_8634,N_8568);
nor U8883 (N_8883,N_8625,N_8619);
nor U8884 (N_8884,N_8737,N_8515);
nor U8885 (N_8885,N_8537,N_8701);
and U8886 (N_8886,N_8629,N_8686);
nor U8887 (N_8887,N_8581,N_8708);
nand U8888 (N_8888,N_8524,N_8746);
xor U8889 (N_8889,N_8645,N_8739);
and U8890 (N_8890,N_8575,N_8636);
nor U8891 (N_8891,N_8676,N_8737);
and U8892 (N_8892,N_8582,N_8617);
and U8893 (N_8893,N_8603,N_8723);
or U8894 (N_8894,N_8601,N_8689);
xor U8895 (N_8895,N_8538,N_8688);
xnor U8896 (N_8896,N_8518,N_8607);
xnor U8897 (N_8897,N_8716,N_8699);
xnor U8898 (N_8898,N_8613,N_8557);
or U8899 (N_8899,N_8500,N_8662);
nor U8900 (N_8900,N_8549,N_8736);
nand U8901 (N_8901,N_8659,N_8612);
nand U8902 (N_8902,N_8719,N_8701);
xor U8903 (N_8903,N_8600,N_8671);
xor U8904 (N_8904,N_8650,N_8574);
nand U8905 (N_8905,N_8644,N_8690);
or U8906 (N_8906,N_8688,N_8747);
and U8907 (N_8907,N_8520,N_8656);
or U8908 (N_8908,N_8514,N_8594);
and U8909 (N_8909,N_8583,N_8733);
nand U8910 (N_8910,N_8642,N_8588);
nor U8911 (N_8911,N_8539,N_8603);
and U8912 (N_8912,N_8512,N_8544);
nand U8913 (N_8913,N_8606,N_8614);
or U8914 (N_8914,N_8506,N_8535);
xnor U8915 (N_8915,N_8690,N_8546);
nand U8916 (N_8916,N_8534,N_8599);
xor U8917 (N_8917,N_8574,N_8600);
and U8918 (N_8918,N_8523,N_8746);
nand U8919 (N_8919,N_8678,N_8596);
xnor U8920 (N_8920,N_8620,N_8736);
nand U8921 (N_8921,N_8553,N_8693);
and U8922 (N_8922,N_8674,N_8507);
and U8923 (N_8923,N_8595,N_8543);
nand U8924 (N_8924,N_8742,N_8677);
nor U8925 (N_8925,N_8601,N_8664);
xnor U8926 (N_8926,N_8675,N_8537);
nor U8927 (N_8927,N_8587,N_8692);
nor U8928 (N_8928,N_8536,N_8546);
or U8929 (N_8929,N_8655,N_8615);
nor U8930 (N_8930,N_8728,N_8651);
nand U8931 (N_8931,N_8533,N_8586);
or U8932 (N_8932,N_8732,N_8557);
and U8933 (N_8933,N_8629,N_8742);
xor U8934 (N_8934,N_8675,N_8658);
nand U8935 (N_8935,N_8662,N_8695);
or U8936 (N_8936,N_8683,N_8565);
nand U8937 (N_8937,N_8561,N_8658);
or U8938 (N_8938,N_8723,N_8671);
nand U8939 (N_8939,N_8689,N_8636);
nand U8940 (N_8940,N_8591,N_8613);
nor U8941 (N_8941,N_8588,N_8547);
and U8942 (N_8942,N_8622,N_8572);
nand U8943 (N_8943,N_8626,N_8591);
nor U8944 (N_8944,N_8568,N_8553);
nand U8945 (N_8945,N_8697,N_8694);
or U8946 (N_8946,N_8573,N_8539);
nor U8947 (N_8947,N_8657,N_8539);
xnor U8948 (N_8948,N_8580,N_8607);
nor U8949 (N_8949,N_8710,N_8501);
nand U8950 (N_8950,N_8701,N_8641);
nand U8951 (N_8951,N_8704,N_8672);
or U8952 (N_8952,N_8654,N_8718);
or U8953 (N_8953,N_8510,N_8693);
xor U8954 (N_8954,N_8659,N_8742);
nand U8955 (N_8955,N_8518,N_8608);
or U8956 (N_8956,N_8535,N_8672);
nor U8957 (N_8957,N_8505,N_8729);
nor U8958 (N_8958,N_8613,N_8744);
nor U8959 (N_8959,N_8593,N_8539);
nor U8960 (N_8960,N_8714,N_8560);
and U8961 (N_8961,N_8557,N_8700);
and U8962 (N_8962,N_8519,N_8505);
xor U8963 (N_8963,N_8505,N_8534);
and U8964 (N_8964,N_8673,N_8686);
or U8965 (N_8965,N_8500,N_8618);
and U8966 (N_8966,N_8562,N_8612);
nand U8967 (N_8967,N_8633,N_8707);
and U8968 (N_8968,N_8556,N_8549);
xor U8969 (N_8969,N_8617,N_8630);
or U8970 (N_8970,N_8748,N_8716);
and U8971 (N_8971,N_8510,N_8635);
and U8972 (N_8972,N_8683,N_8619);
nand U8973 (N_8973,N_8601,N_8535);
nor U8974 (N_8974,N_8714,N_8598);
and U8975 (N_8975,N_8556,N_8663);
nand U8976 (N_8976,N_8546,N_8741);
nand U8977 (N_8977,N_8732,N_8655);
xnor U8978 (N_8978,N_8597,N_8668);
nor U8979 (N_8979,N_8647,N_8542);
nand U8980 (N_8980,N_8719,N_8663);
or U8981 (N_8981,N_8681,N_8563);
nand U8982 (N_8982,N_8684,N_8578);
and U8983 (N_8983,N_8614,N_8595);
and U8984 (N_8984,N_8665,N_8671);
nand U8985 (N_8985,N_8513,N_8655);
nand U8986 (N_8986,N_8639,N_8512);
nand U8987 (N_8987,N_8670,N_8625);
or U8988 (N_8988,N_8593,N_8541);
nor U8989 (N_8989,N_8662,N_8632);
and U8990 (N_8990,N_8599,N_8683);
nand U8991 (N_8991,N_8738,N_8667);
nand U8992 (N_8992,N_8664,N_8579);
or U8993 (N_8993,N_8689,N_8688);
xor U8994 (N_8994,N_8572,N_8718);
nor U8995 (N_8995,N_8594,N_8668);
xor U8996 (N_8996,N_8674,N_8592);
xnor U8997 (N_8997,N_8706,N_8531);
or U8998 (N_8998,N_8627,N_8517);
or U8999 (N_8999,N_8692,N_8748);
nor U9000 (N_9000,N_8817,N_8957);
and U9001 (N_9001,N_8949,N_8778);
xor U9002 (N_9002,N_8855,N_8991);
nand U9003 (N_9003,N_8816,N_8809);
nand U9004 (N_9004,N_8948,N_8942);
and U9005 (N_9005,N_8850,N_8854);
and U9006 (N_9006,N_8937,N_8763);
or U9007 (N_9007,N_8988,N_8874);
nor U9008 (N_9008,N_8878,N_8846);
nand U9009 (N_9009,N_8917,N_8784);
nor U9010 (N_9010,N_8896,N_8931);
xor U9011 (N_9011,N_8925,N_8836);
xor U9012 (N_9012,N_8813,N_8773);
nor U9013 (N_9013,N_8819,N_8835);
xnor U9014 (N_9014,N_8873,N_8939);
nor U9015 (N_9015,N_8914,N_8760);
nor U9016 (N_9016,N_8822,N_8840);
and U9017 (N_9017,N_8843,N_8879);
xnor U9018 (N_9018,N_8791,N_8828);
nor U9019 (N_9019,N_8811,N_8834);
nor U9020 (N_9020,N_8865,N_8987);
xnor U9021 (N_9021,N_8792,N_8989);
or U9022 (N_9022,N_8969,N_8812);
and U9023 (N_9023,N_8802,N_8797);
or U9024 (N_9024,N_8909,N_8882);
xnor U9025 (N_9025,N_8783,N_8839);
and U9026 (N_9026,N_8990,N_8848);
nand U9027 (N_9027,N_8963,N_8830);
or U9028 (N_9028,N_8867,N_8768);
nand U9029 (N_9029,N_8968,N_8757);
nor U9030 (N_9030,N_8751,N_8858);
and U9031 (N_9031,N_8984,N_8789);
and U9032 (N_9032,N_8982,N_8892);
or U9033 (N_9033,N_8871,N_8851);
nand U9034 (N_9034,N_8952,N_8947);
xnor U9035 (N_9035,N_8894,N_8814);
or U9036 (N_9036,N_8861,N_8767);
nand U9037 (N_9037,N_8924,N_8979);
nand U9038 (N_9038,N_8774,N_8771);
or U9039 (N_9039,N_8859,N_8862);
and U9040 (N_9040,N_8764,N_8903);
nand U9041 (N_9041,N_8964,N_8908);
nor U9042 (N_9042,N_8772,N_8777);
nor U9043 (N_9043,N_8825,N_8842);
or U9044 (N_9044,N_8953,N_8833);
nor U9045 (N_9045,N_8911,N_8943);
and U9046 (N_9046,N_8936,N_8945);
nor U9047 (N_9047,N_8794,N_8927);
nand U9048 (N_9048,N_8818,N_8923);
nor U9049 (N_9049,N_8913,N_8820);
nand U9050 (N_9050,N_8847,N_8750);
or U9051 (N_9051,N_8844,N_8761);
nor U9052 (N_9052,N_8907,N_8829);
or U9053 (N_9053,N_8920,N_8826);
nor U9054 (N_9054,N_8916,N_8869);
or U9055 (N_9055,N_8889,N_8800);
xnor U9056 (N_9056,N_8770,N_8863);
nor U9057 (N_9057,N_8785,N_8769);
nand U9058 (N_9058,N_8827,N_8995);
or U9059 (N_9059,N_8870,N_8912);
xnor U9060 (N_9060,N_8806,N_8919);
nand U9061 (N_9061,N_8838,N_8926);
nand U9062 (N_9062,N_8753,N_8849);
and U9063 (N_9063,N_8886,N_8877);
xor U9064 (N_9064,N_8985,N_8910);
or U9065 (N_9065,N_8853,N_8993);
or U9066 (N_9066,N_8810,N_8994);
or U9067 (N_9067,N_8966,N_8956);
or U9068 (N_9068,N_8946,N_8845);
nor U9069 (N_9069,N_8796,N_8805);
xor U9070 (N_9070,N_8958,N_8932);
nand U9071 (N_9071,N_8997,N_8996);
and U9072 (N_9072,N_8951,N_8961);
xnor U9073 (N_9073,N_8999,N_8795);
nor U9074 (N_9074,N_8790,N_8980);
nand U9075 (N_9075,N_8758,N_8856);
nor U9076 (N_9076,N_8974,N_8897);
nor U9077 (N_9077,N_8793,N_8918);
and U9078 (N_9078,N_8821,N_8883);
xor U9079 (N_9079,N_8954,N_8905);
nor U9080 (N_9080,N_8782,N_8803);
xnor U9081 (N_9081,N_8754,N_8787);
nor U9082 (N_9082,N_8752,N_8786);
nor U9083 (N_9083,N_8807,N_8959);
nor U9084 (N_9084,N_8832,N_8938);
or U9085 (N_9085,N_8895,N_8798);
xor U9086 (N_9086,N_8866,N_8935);
xor U9087 (N_9087,N_8900,N_8823);
nor U9088 (N_9088,N_8899,N_8981);
or U9089 (N_9089,N_8940,N_8950);
or U9090 (N_9090,N_8887,N_8781);
nor U9091 (N_9091,N_8901,N_8902);
or U9092 (N_9092,N_8766,N_8978);
or U9093 (N_9093,N_8967,N_8801);
or U9094 (N_9094,N_8880,N_8824);
and U9095 (N_9095,N_8804,N_8998);
or U9096 (N_9096,N_8884,N_8972);
nor U9097 (N_9097,N_8759,N_8992);
or U9098 (N_9098,N_8872,N_8970);
or U9099 (N_9099,N_8971,N_8775);
nand U9100 (N_9100,N_8906,N_8831);
and U9101 (N_9101,N_8976,N_8780);
and U9102 (N_9102,N_8929,N_8930);
and U9103 (N_9103,N_8941,N_8915);
xnor U9104 (N_9104,N_8944,N_8841);
or U9105 (N_9105,N_8922,N_8779);
xor U9106 (N_9106,N_8788,N_8977);
and U9107 (N_9107,N_8815,N_8864);
nor U9108 (N_9108,N_8852,N_8885);
or U9109 (N_9109,N_8868,N_8756);
nand U9110 (N_9110,N_8762,N_8921);
xor U9111 (N_9111,N_8875,N_8860);
or U9112 (N_9112,N_8857,N_8973);
or U9113 (N_9113,N_8808,N_8965);
nand U9114 (N_9114,N_8983,N_8876);
and U9115 (N_9115,N_8934,N_8888);
nand U9116 (N_9116,N_8890,N_8891);
nor U9117 (N_9117,N_8765,N_8837);
or U9118 (N_9118,N_8960,N_8799);
nand U9119 (N_9119,N_8986,N_8904);
xor U9120 (N_9120,N_8962,N_8933);
or U9121 (N_9121,N_8955,N_8893);
and U9122 (N_9122,N_8776,N_8898);
and U9123 (N_9123,N_8755,N_8881);
and U9124 (N_9124,N_8975,N_8928);
xnor U9125 (N_9125,N_8803,N_8962);
nand U9126 (N_9126,N_8828,N_8820);
or U9127 (N_9127,N_8982,N_8808);
nand U9128 (N_9128,N_8913,N_8764);
and U9129 (N_9129,N_8926,N_8854);
xor U9130 (N_9130,N_8917,N_8793);
or U9131 (N_9131,N_8837,N_8867);
and U9132 (N_9132,N_8887,N_8897);
and U9133 (N_9133,N_8897,N_8862);
xor U9134 (N_9134,N_8902,N_8759);
and U9135 (N_9135,N_8750,N_8761);
nor U9136 (N_9136,N_8969,N_8834);
nand U9137 (N_9137,N_8997,N_8953);
and U9138 (N_9138,N_8918,N_8825);
nor U9139 (N_9139,N_8884,N_8910);
or U9140 (N_9140,N_8774,N_8881);
or U9141 (N_9141,N_8752,N_8918);
and U9142 (N_9142,N_8801,N_8877);
nand U9143 (N_9143,N_8755,N_8821);
or U9144 (N_9144,N_8763,N_8826);
or U9145 (N_9145,N_8927,N_8751);
xnor U9146 (N_9146,N_8973,N_8879);
xnor U9147 (N_9147,N_8896,N_8966);
and U9148 (N_9148,N_8751,N_8806);
xor U9149 (N_9149,N_8969,N_8779);
nand U9150 (N_9150,N_8904,N_8974);
nor U9151 (N_9151,N_8851,N_8816);
or U9152 (N_9152,N_8986,N_8979);
nand U9153 (N_9153,N_8762,N_8924);
xor U9154 (N_9154,N_8814,N_8789);
nand U9155 (N_9155,N_8987,N_8868);
nor U9156 (N_9156,N_8803,N_8783);
nand U9157 (N_9157,N_8789,N_8983);
nor U9158 (N_9158,N_8878,N_8803);
or U9159 (N_9159,N_8824,N_8994);
xor U9160 (N_9160,N_8911,N_8874);
and U9161 (N_9161,N_8896,N_8898);
and U9162 (N_9162,N_8786,N_8814);
and U9163 (N_9163,N_8826,N_8765);
or U9164 (N_9164,N_8968,N_8816);
and U9165 (N_9165,N_8796,N_8852);
nor U9166 (N_9166,N_8919,N_8974);
nand U9167 (N_9167,N_8943,N_8849);
or U9168 (N_9168,N_8964,N_8954);
xor U9169 (N_9169,N_8985,N_8979);
and U9170 (N_9170,N_8763,N_8797);
nand U9171 (N_9171,N_8921,N_8937);
nor U9172 (N_9172,N_8849,N_8938);
and U9173 (N_9173,N_8752,N_8758);
xnor U9174 (N_9174,N_8946,N_8884);
and U9175 (N_9175,N_8885,N_8821);
and U9176 (N_9176,N_8760,N_8840);
nand U9177 (N_9177,N_8853,N_8999);
nand U9178 (N_9178,N_8923,N_8893);
and U9179 (N_9179,N_8781,N_8791);
and U9180 (N_9180,N_8887,N_8951);
xor U9181 (N_9181,N_8794,N_8841);
xnor U9182 (N_9182,N_8998,N_8920);
nor U9183 (N_9183,N_8820,N_8942);
nor U9184 (N_9184,N_8973,N_8914);
and U9185 (N_9185,N_8833,N_8857);
nor U9186 (N_9186,N_8877,N_8943);
or U9187 (N_9187,N_8863,N_8867);
or U9188 (N_9188,N_8941,N_8958);
and U9189 (N_9189,N_8791,N_8940);
nor U9190 (N_9190,N_8921,N_8782);
nand U9191 (N_9191,N_8753,N_8918);
nor U9192 (N_9192,N_8829,N_8959);
nand U9193 (N_9193,N_8944,N_8983);
nand U9194 (N_9194,N_8993,N_8918);
or U9195 (N_9195,N_8888,N_8913);
or U9196 (N_9196,N_8808,N_8860);
or U9197 (N_9197,N_8860,N_8945);
nand U9198 (N_9198,N_8798,N_8986);
and U9199 (N_9199,N_8942,N_8937);
and U9200 (N_9200,N_8798,N_8898);
and U9201 (N_9201,N_8787,N_8872);
nand U9202 (N_9202,N_8775,N_8975);
nor U9203 (N_9203,N_8992,N_8764);
or U9204 (N_9204,N_8828,N_8997);
xor U9205 (N_9205,N_8757,N_8924);
or U9206 (N_9206,N_8757,N_8917);
or U9207 (N_9207,N_8821,N_8878);
nand U9208 (N_9208,N_8830,N_8886);
nor U9209 (N_9209,N_8845,N_8979);
xor U9210 (N_9210,N_8909,N_8768);
nor U9211 (N_9211,N_8837,N_8943);
or U9212 (N_9212,N_8820,N_8994);
or U9213 (N_9213,N_8767,N_8888);
nand U9214 (N_9214,N_8751,N_8788);
and U9215 (N_9215,N_8763,N_8954);
or U9216 (N_9216,N_8762,N_8825);
xor U9217 (N_9217,N_8966,N_8843);
nor U9218 (N_9218,N_8805,N_8878);
nor U9219 (N_9219,N_8959,N_8955);
xor U9220 (N_9220,N_8921,N_8802);
xor U9221 (N_9221,N_8963,N_8752);
nor U9222 (N_9222,N_8823,N_8860);
xnor U9223 (N_9223,N_8940,N_8944);
nor U9224 (N_9224,N_8999,N_8777);
or U9225 (N_9225,N_8757,N_8881);
or U9226 (N_9226,N_8928,N_8996);
xor U9227 (N_9227,N_8801,N_8890);
or U9228 (N_9228,N_8769,N_8963);
xnor U9229 (N_9229,N_8904,N_8758);
nor U9230 (N_9230,N_8907,N_8859);
and U9231 (N_9231,N_8792,N_8981);
and U9232 (N_9232,N_8841,N_8793);
and U9233 (N_9233,N_8832,N_8860);
nand U9234 (N_9234,N_8961,N_8856);
nand U9235 (N_9235,N_8815,N_8840);
or U9236 (N_9236,N_8914,N_8953);
or U9237 (N_9237,N_8918,N_8818);
and U9238 (N_9238,N_8904,N_8814);
xnor U9239 (N_9239,N_8814,N_8806);
xnor U9240 (N_9240,N_8849,N_8752);
nor U9241 (N_9241,N_8930,N_8853);
xor U9242 (N_9242,N_8916,N_8828);
and U9243 (N_9243,N_8873,N_8776);
nor U9244 (N_9244,N_8919,N_8978);
nand U9245 (N_9245,N_8887,N_8852);
nor U9246 (N_9246,N_8780,N_8951);
and U9247 (N_9247,N_8894,N_8890);
nand U9248 (N_9248,N_8972,N_8784);
xor U9249 (N_9249,N_8911,N_8871);
and U9250 (N_9250,N_9180,N_9186);
and U9251 (N_9251,N_9000,N_9051);
nor U9252 (N_9252,N_9028,N_9063);
and U9253 (N_9253,N_9197,N_9171);
xor U9254 (N_9254,N_9007,N_9016);
nand U9255 (N_9255,N_9229,N_9239);
xor U9256 (N_9256,N_9097,N_9209);
or U9257 (N_9257,N_9027,N_9108);
nor U9258 (N_9258,N_9191,N_9029);
nand U9259 (N_9259,N_9129,N_9151);
nor U9260 (N_9260,N_9124,N_9144);
or U9261 (N_9261,N_9162,N_9178);
or U9262 (N_9262,N_9048,N_9181);
or U9263 (N_9263,N_9207,N_9226);
xor U9264 (N_9264,N_9185,N_9070);
xnor U9265 (N_9265,N_9231,N_9135);
nand U9266 (N_9266,N_9174,N_9216);
and U9267 (N_9267,N_9009,N_9023);
and U9268 (N_9268,N_9213,N_9044);
xor U9269 (N_9269,N_9082,N_9179);
and U9270 (N_9270,N_9134,N_9106);
xnor U9271 (N_9271,N_9177,N_9221);
xnor U9272 (N_9272,N_9212,N_9034);
and U9273 (N_9273,N_9224,N_9208);
nor U9274 (N_9274,N_9033,N_9030);
or U9275 (N_9275,N_9159,N_9107);
xor U9276 (N_9276,N_9073,N_9215);
and U9277 (N_9277,N_9094,N_9093);
nor U9278 (N_9278,N_9117,N_9182);
or U9279 (N_9279,N_9080,N_9133);
nor U9280 (N_9280,N_9014,N_9214);
nor U9281 (N_9281,N_9205,N_9166);
xnor U9282 (N_9282,N_9172,N_9223);
nor U9283 (N_9283,N_9052,N_9195);
or U9284 (N_9284,N_9010,N_9150);
nand U9285 (N_9285,N_9025,N_9217);
nand U9286 (N_9286,N_9118,N_9188);
or U9287 (N_9287,N_9086,N_9131);
or U9288 (N_9288,N_9031,N_9170);
or U9289 (N_9289,N_9098,N_9194);
nand U9290 (N_9290,N_9243,N_9038);
nand U9291 (N_9291,N_9112,N_9109);
nand U9292 (N_9292,N_9020,N_9167);
or U9293 (N_9293,N_9163,N_9200);
nand U9294 (N_9294,N_9183,N_9228);
xnor U9295 (N_9295,N_9203,N_9176);
nor U9296 (N_9296,N_9077,N_9138);
or U9297 (N_9297,N_9004,N_9045);
xor U9298 (N_9298,N_9210,N_9237);
or U9299 (N_9299,N_9060,N_9152);
xnor U9300 (N_9300,N_9041,N_9100);
xnor U9301 (N_9301,N_9090,N_9068);
xnor U9302 (N_9302,N_9246,N_9196);
nand U9303 (N_9303,N_9003,N_9130);
nor U9304 (N_9304,N_9184,N_9132);
xnor U9305 (N_9305,N_9247,N_9111);
nor U9306 (N_9306,N_9227,N_9046);
nand U9307 (N_9307,N_9099,N_9039);
and U9308 (N_9308,N_9116,N_9206);
and U9309 (N_9309,N_9232,N_9062);
or U9310 (N_9310,N_9083,N_9235);
or U9311 (N_9311,N_9049,N_9218);
xnor U9312 (N_9312,N_9160,N_9050);
and U9313 (N_9313,N_9120,N_9015);
xor U9314 (N_9314,N_9055,N_9140);
nand U9315 (N_9315,N_9219,N_9149);
nor U9316 (N_9316,N_9242,N_9156);
and U9317 (N_9317,N_9084,N_9145);
nand U9318 (N_9318,N_9040,N_9095);
nand U9319 (N_9319,N_9187,N_9240);
nand U9320 (N_9320,N_9190,N_9026);
or U9321 (N_9321,N_9008,N_9067);
and U9322 (N_9322,N_9079,N_9220);
xor U9323 (N_9323,N_9173,N_9076);
nand U9324 (N_9324,N_9043,N_9126);
and U9325 (N_9325,N_9245,N_9192);
nand U9326 (N_9326,N_9136,N_9175);
and U9327 (N_9327,N_9137,N_9085);
and U9328 (N_9328,N_9072,N_9081);
nand U9329 (N_9329,N_9092,N_9164);
xnor U9330 (N_9330,N_9248,N_9204);
xnor U9331 (N_9331,N_9249,N_9065);
nand U9332 (N_9332,N_9211,N_9168);
xnor U9333 (N_9333,N_9054,N_9238);
nor U9334 (N_9334,N_9103,N_9121);
or U9335 (N_9335,N_9096,N_9113);
and U9336 (N_9336,N_9193,N_9110);
or U9337 (N_9337,N_9021,N_9234);
and U9338 (N_9338,N_9061,N_9078);
nand U9339 (N_9339,N_9037,N_9169);
and U9340 (N_9340,N_9053,N_9241);
or U9341 (N_9341,N_9042,N_9056);
and U9342 (N_9342,N_9089,N_9146);
nand U9343 (N_9343,N_9155,N_9142);
or U9344 (N_9344,N_9153,N_9017);
or U9345 (N_9345,N_9001,N_9036);
nor U9346 (N_9346,N_9011,N_9087);
xnor U9347 (N_9347,N_9022,N_9075);
or U9348 (N_9348,N_9147,N_9202);
or U9349 (N_9349,N_9225,N_9161);
nand U9350 (N_9350,N_9157,N_9102);
or U9351 (N_9351,N_9141,N_9066);
xor U9352 (N_9352,N_9158,N_9064);
and U9353 (N_9353,N_9013,N_9018);
or U9354 (N_9354,N_9198,N_9127);
nor U9355 (N_9355,N_9104,N_9101);
and U9356 (N_9356,N_9057,N_9123);
xnor U9357 (N_9357,N_9201,N_9125);
and U9358 (N_9358,N_9091,N_9244);
or U9359 (N_9359,N_9058,N_9222);
and U9360 (N_9360,N_9154,N_9189);
and U9361 (N_9361,N_9115,N_9059);
xnor U9362 (N_9362,N_9128,N_9088);
xnor U9363 (N_9363,N_9006,N_9071);
or U9364 (N_9364,N_9114,N_9236);
nand U9365 (N_9365,N_9119,N_9230);
xor U9366 (N_9366,N_9035,N_9005);
or U9367 (N_9367,N_9032,N_9165);
nand U9368 (N_9368,N_9199,N_9002);
xor U9369 (N_9369,N_9047,N_9233);
nand U9370 (N_9370,N_9069,N_9024);
xnor U9371 (N_9371,N_9148,N_9122);
and U9372 (N_9372,N_9074,N_9105);
nor U9373 (N_9373,N_9139,N_9019);
nor U9374 (N_9374,N_9012,N_9143);
xor U9375 (N_9375,N_9034,N_9115);
nor U9376 (N_9376,N_9232,N_9193);
or U9377 (N_9377,N_9133,N_9017);
nor U9378 (N_9378,N_9205,N_9219);
and U9379 (N_9379,N_9179,N_9022);
and U9380 (N_9380,N_9071,N_9170);
and U9381 (N_9381,N_9167,N_9184);
or U9382 (N_9382,N_9232,N_9242);
xor U9383 (N_9383,N_9239,N_9246);
or U9384 (N_9384,N_9084,N_9177);
and U9385 (N_9385,N_9031,N_9116);
nor U9386 (N_9386,N_9085,N_9218);
and U9387 (N_9387,N_9204,N_9198);
xnor U9388 (N_9388,N_9123,N_9083);
nand U9389 (N_9389,N_9132,N_9095);
xnor U9390 (N_9390,N_9073,N_9244);
and U9391 (N_9391,N_9174,N_9119);
nor U9392 (N_9392,N_9022,N_9119);
nor U9393 (N_9393,N_9234,N_9140);
nor U9394 (N_9394,N_9142,N_9006);
nand U9395 (N_9395,N_9126,N_9125);
and U9396 (N_9396,N_9133,N_9208);
or U9397 (N_9397,N_9232,N_9142);
nand U9398 (N_9398,N_9220,N_9031);
xor U9399 (N_9399,N_9099,N_9171);
or U9400 (N_9400,N_9121,N_9187);
and U9401 (N_9401,N_9066,N_9005);
or U9402 (N_9402,N_9241,N_9248);
nand U9403 (N_9403,N_9107,N_9236);
nand U9404 (N_9404,N_9083,N_9110);
xnor U9405 (N_9405,N_9245,N_9220);
nor U9406 (N_9406,N_9163,N_9032);
and U9407 (N_9407,N_9218,N_9141);
or U9408 (N_9408,N_9043,N_9050);
nand U9409 (N_9409,N_9176,N_9003);
nand U9410 (N_9410,N_9094,N_9004);
nand U9411 (N_9411,N_9140,N_9201);
nor U9412 (N_9412,N_9094,N_9096);
nand U9413 (N_9413,N_9181,N_9091);
and U9414 (N_9414,N_9022,N_9205);
nor U9415 (N_9415,N_9049,N_9059);
xor U9416 (N_9416,N_9196,N_9068);
and U9417 (N_9417,N_9057,N_9181);
nor U9418 (N_9418,N_9036,N_9222);
nand U9419 (N_9419,N_9160,N_9066);
and U9420 (N_9420,N_9117,N_9193);
and U9421 (N_9421,N_9001,N_9086);
and U9422 (N_9422,N_9108,N_9160);
xnor U9423 (N_9423,N_9139,N_9086);
xnor U9424 (N_9424,N_9142,N_9223);
nand U9425 (N_9425,N_9164,N_9121);
nor U9426 (N_9426,N_9248,N_9228);
or U9427 (N_9427,N_9029,N_9193);
and U9428 (N_9428,N_9179,N_9107);
nor U9429 (N_9429,N_9070,N_9091);
xor U9430 (N_9430,N_9100,N_9193);
nor U9431 (N_9431,N_9194,N_9112);
and U9432 (N_9432,N_9197,N_9056);
or U9433 (N_9433,N_9249,N_9044);
nand U9434 (N_9434,N_9227,N_9074);
and U9435 (N_9435,N_9058,N_9052);
nand U9436 (N_9436,N_9127,N_9191);
nand U9437 (N_9437,N_9144,N_9115);
xor U9438 (N_9438,N_9156,N_9143);
or U9439 (N_9439,N_9028,N_9241);
xnor U9440 (N_9440,N_9159,N_9095);
xnor U9441 (N_9441,N_9028,N_9057);
nand U9442 (N_9442,N_9027,N_9003);
or U9443 (N_9443,N_9015,N_9148);
nand U9444 (N_9444,N_9182,N_9071);
nand U9445 (N_9445,N_9000,N_9236);
and U9446 (N_9446,N_9094,N_9047);
and U9447 (N_9447,N_9037,N_9163);
or U9448 (N_9448,N_9243,N_9034);
nand U9449 (N_9449,N_9133,N_9177);
and U9450 (N_9450,N_9080,N_9209);
or U9451 (N_9451,N_9018,N_9096);
and U9452 (N_9452,N_9162,N_9061);
or U9453 (N_9453,N_9186,N_9026);
nor U9454 (N_9454,N_9143,N_9175);
or U9455 (N_9455,N_9153,N_9024);
or U9456 (N_9456,N_9193,N_9217);
and U9457 (N_9457,N_9029,N_9225);
and U9458 (N_9458,N_9221,N_9178);
or U9459 (N_9459,N_9154,N_9222);
nand U9460 (N_9460,N_9089,N_9184);
or U9461 (N_9461,N_9015,N_9228);
xor U9462 (N_9462,N_9151,N_9186);
nand U9463 (N_9463,N_9033,N_9112);
or U9464 (N_9464,N_9096,N_9023);
nor U9465 (N_9465,N_9160,N_9022);
nor U9466 (N_9466,N_9056,N_9121);
and U9467 (N_9467,N_9085,N_9091);
nand U9468 (N_9468,N_9197,N_9063);
nor U9469 (N_9469,N_9022,N_9028);
or U9470 (N_9470,N_9161,N_9121);
xor U9471 (N_9471,N_9083,N_9093);
nor U9472 (N_9472,N_9238,N_9189);
nand U9473 (N_9473,N_9114,N_9145);
nor U9474 (N_9474,N_9141,N_9063);
xor U9475 (N_9475,N_9216,N_9043);
xnor U9476 (N_9476,N_9001,N_9103);
nand U9477 (N_9477,N_9137,N_9108);
or U9478 (N_9478,N_9093,N_9159);
xnor U9479 (N_9479,N_9128,N_9049);
nand U9480 (N_9480,N_9235,N_9139);
nor U9481 (N_9481,N_9057,N_9103);
xor U9482 (N_9482,N_9055,N_9121);
and U9483 (N_9483,N_9089,N_9233);
nor U9484 (N_9484,N_9055,N_9096);
nor U9485 (N_9485,N_9075,N_9039);
and U9486 (N_9486,N_9241,N_9244);
nand U9487 (N_9487,N_9097,N_9186);
and U9488 (N_9488,N_9005,N_9133);
or U9489 (N_9489,N_9239,N_9141);
xnor U9490 (N_9490,N_9199,N_9107);
nor U9491 (N_9491,N_9018,N_9243);
nand U9492 (N_9492,N_9049,N_9077);
xnor U9493 (N_9493,N_9015,N_9058);
xnor U9494 (N_9494,N_9105,N_9168);
xor U9495 (N_9495,N_9138,N_9222);
nand U9496 (N_9496,N_9095,N_9208);
nand U9497 (N_9497,N_9243,N_9020);
or U9498 (N_9498,N_9151,N_9039);
nand U9499 (N_9499,N_9139,N_9047);
xor U9500 (N_9500,N_9306,N_9444);
nor U9501 (N_9501,N_9317,N_9481);
nand U9502 (N_9502,N_9373,N_9251);
and U9503 (N_9503,N_9318,N_9483);
or U9504 (N_9504,N_9439,N_9377);
nand U9505 (N_9505,N_9300,N_9312);
xnor U9506 (N_9506,N_9342,N_9428);
or U9507 (N_9507,N_9299,N_9424);
or U9508 (N_9508,N_9388,N_9260);
or U9509 (N_9509,N_9253,N_9265);
nor U9510 (N_9510,N_9485,N_9297);
nand U9511 (N_9511,N_9291,N_9325);
or U9512 (N_9512,N_9418,N_9262);
nor U9513 (N_9513,N_9304,N_9358);
nor U9514 (N_9514,N_9316,N_9264);
xnor U9515 (N_9515,N_9386,N_9448);
xor U9516 (N_9516,N_9463,N_9307);
or U9517 (N_9517,N_9349,N_9412);
nand U9518 (N_9518,N_9414,N_9496);
xnor U9519 (N_9519,N_9427,N_9362);
nand U9520 (N_9520,N_9438,N_9492);
xnor U9521 (N_9521,N_9403,N_9399);
nor U9522 (N_9522,N_9415,N_9437);
or U9523 (N_9523,N_9322,N_9259);
nor U9524 (N_9524,N_9335,N_9445);
nand U9525 (N_9525,N_9310,N_9390);
nand U9526 (N_9526,N_9442,N_9446);
and U9527 (N_9527,N_9371,N_9423);
xnor U9528 (N_9528,N_9408,N_9268);
xnor U9529 (N_9529,N_9337,N_9287);
or U9530 (N_9530,N_9263,N_9473);
nor U9531 (N_9531,N_9256,N_9350);
or U9532 (N_9532,N_9394,N_9449);
nor U9533 (N_9533,N_9383,N_9491);
xor U9534 (N_9534,N_9339,N_9488);
or U9535 (N_9535,N_9401,N_9393);
nor U9536 (N_9536,N_9450,N_9289);
nand U9537 (N_9537,N_9426,N_9254);
nor U9538 (N_9538,N_9486,N_9462);
and U9539 (N_9539,N_9459,N_9348);
and U9540 (N_9540,N_9308,N_9368);
and U9541 (N_9541,N_9315,N_9277);
nor U9542 (N_9542,N_9319,N_9425);
or U9543 (N_9543,N_9366,N_9255);
or U9544 (N_9544,N_9406,N_9364);
nand U9545 (N_9545,N_9476,N_9497);
nand U9546 (N_9546,N_9484,N_9435);
nor U9547 (N_9547,N_9326,N_9471);
or U9548 (N_9548,N_9278,N_9392);
xor U9549 (N_9549,N_9271,N_9498);
xor U9550 (N_9550,N_9290,N_9402);
nor U9551 (N_9551,N_9344,N_9280);
nor U9552 (N_9552,N_9381,N_9279);
xor U9553 (N_9553,N_9327,N_9283);
xnor U9554 (N_9554,N_9396,N_9420);
or U9555 (N_9555,N_9343,N_9477);
and U9556 (N_9556,N_9365,N_9455);
and U9557 (N_9557,N_9313,N_9285);
nor U9558 (N_9558,N_9417,N_9338);
and U9559 (N_9559,N_9398,N_9469);
xor U9560 (N_9560,N_9372,N_9434);
and U9561 (N_9561,N_9303,N_9369);
nor U9562 (N_9562,N_9457,N_9487);
nand U9563 (N_9563,N_9341,N_9475);
xor U9564 (N_9564,N_9452,N_9458);
and U9565 (N_9565,N_9353,N_9433);
xor U9566 (N_9566,N_9490,N_9361);
and U9567 (N_9567,N_9269,N_9272);
xor U9568 (N_9568,N_9465,N_9384);
or U9569 (N_9569,N_9472,N_9385);
and U9570 (N_9570,N_9461,N_9382);
nand U9571 (N_9571,N_9411,N_9466);
xnor U9572 (N_9572,N_9321,N_9389);
nand U9573 (N_9573,N_9478,N_9309);
and U9574 (N_9574,N_9295,N_9354);
xor U9575 (N_9575,N_9422,N_9324);
or U9576 (N_9576,N_9467,N_9429);
nand U9577 (N_9577,N_9347,N_9495);
or U9578 (N_9578,N_9419,N_9404);
nor U9579 (N_9579,N_9410,N_9331);
nor U9580 (N_9580,N_9293,N_9274);
or U9581 (N_9581,N_9376,N_9480);
nor U9582 (N_9582,N_9298,N_9250);
xor U9583 (N_9583,N_9284,N_9387);
nor U9584 (N_9584,N_9356,N_9286);
nor U9585 (N_9585,N_9447,N_9405);
nand U9586 (N_9586,N_9430,N_9267);
nand U9587 (N_9587,N_9440,N_9380);
nand U9588 (N_9588,N_9421,N_9351);
or U9589 (N_9589,N_9258,N_9363);
or U9590 (N_9590,N_9332,N_9266);
or U9591 (N_9591,N_9370,N_9328);
nand U9592 (N_9592,N_9296,N_9416);
xnor U9593 (N_9593,N_9311,N_9275);
xnor U9594 (N_9594,N_9499,N_9357);
or U9595 (N_9595,N_9340,N_9454);
or U9596 (N_9596,N_9456,N_9441);
or U9597 (N_9597,N_9333,N_9288);
nand U9598 (N_9598,N_9379,N_9468);
and U9599 (N_9599,N_9474,N_9346);
nand U9600 (N_9600,N_9443,N_9367);
xnor U9601 (N_9601,N_9323,N_9436);
or U9602 (N_9602,N_9432,N_9352);
xor U9603 (N_9603,N_9294,N_9329);
or U9604 (N_9604,N_9282,N_9378);
and U9605 (N_9605,N_9453,N_9345);
and U9606 (N_9606,N_9270,N_9395);
nor U9607 (N_9607,N_9334,N_9409);
and U9608 (N_9608,N_9273,N_9407);
or U9609 (N_9609,N_9451,N_9470);
or U9610 (N_9610,N_9482,N_9391);
nor U9611 (N_9611,N_9413,N_9301);
nor U9612 (N_9612,N_9359,N_9360);
xor U9613 (N_9613,N_9320,N_9397);
xnor U9614 (N_9614,N_9336,N_9355);
or U9615 (N_9615,N_9292,N_9400);
nor U9616 (N_9616,N_9494,N_9493);
or U9617 (N_9617,N_9261,N_9464);
and U9618 (N_9618,N_9314,N_9257);
or U9619 (N_9619,N_9330,N_9375);
xor U9620 (N_9620,N_9431,N_9276);
or U9621 (N_9621,N_9479,N_9252);
xor U9622 (N_9622,N_9374,N_9281);
nor U9623 (N_9623,N_9460,N_9489);
and U9624 (N_9624,N_9305,N_9302);
nor U9625 (N_9625,N_9439,N_9255);
nor U9626 (N_9626,N_9367,N_9300);
and U9627 (N_9627,N_9421,N_9329);
nand U9628 (N_9628,N_9347,N_9306);
or U9629 (N_9629,N_9457,N_9393);
xor U9630 (N_9630,N_9295,N_9292);
nor U9631 (N_9631,N_9300,N_9253);
or U9632 (N_9632,N_9396,N_9455);
nor U9633 (N_9633,N_9344,N_9495);
or U9634 (N_9634,N_9435,N_9390);
or U9635 (N_9635,N_9376,N_9263);
xor U9636 (N_9636,N_9497,N_9290);
or U9637 (N_9637,N_9421,N_9288);
and U9638 (N_9638,N_9398,N_9295);
and U9639 (N_9639,N_9383,N_9490);
nor U9640 (N_9640,N_9447,N_9438);
xnor U9641 (N_9641,N_9377,N_9357);
nand U9642 (N_9642,N_9354,N_9435);
nand U9643 (N_9643,N_9298,N_9287);
nand U9644 (N_9644,N_9348,N_9493);
nor U9645 (N_9645,N_9337,N_9474);
or U9646 (N_9646,N_9365,N_9258);
xnor U9647 (N_9647,N_9289,N_9351);
and U9648 (N_9648,N_9425,N_9290);
xor U9649 (N_9649,N_9270,N_9497);
xnor U9650 (N_9650,N_9407,N_9258);
and U9651 (N_9651,N_9411,N_9322);
and U9652 (N_9652,N_9292,N_9489);
nor U9653 (N_9653,N_9465,N_9333);
xor U9654 (N_9654,N_9396,N_9378);
nand U9655 (N_9655,N_9367,N_9333);
nor U9656 (N_9656,N_9344,N_9309);
xnor U9657 (N_9657,N_9298,N_9393);
nor U9658 (N_9658,N_9363,N_9375);
nor U9659 (N_9659,N_9399,N_9354);
and U9660 (N_9660,N_9266,N_9272);
nand U9661 (N_9661,N_9420,N_9284);
and U9662 (N_9662,N_9444,N_9416);
nand U9663 (N_9663,N_9341,N_9270);
nand U9664 (N_9664,N_9468,N_9283);
xnor U9665 (N_9665,N_9384,N_9486);
or U9666 (N_9666,N_9465,N_9320);
nor U9667 (N_9667,N_9286,N_9476);
nand U9668 (N_9668,N_9269,N_9461);
xor U9669 (N_9669,N_9324,N_9496);
or U9670 (N_9670,N_9381,N_9436);
or U9671 (N_9671,N_9370,N_9431);
xnor U9672 (N_9672,N_9493,N_9277);
nand U9673 (N_9673,N_9490,N_9379);
and U9674 (N_9674,N_9447,N_9341);
nor U9675 (N_9675,N_9280,N_9339);
or U9676 (N_9676,N_9441,N_9371);
xor U9677 (N_9677,N_9282,N_9287);
nor U9678 (N_9678,N_9386,N_9457);
and U9679 (N_9679,N_9374,N_9465);
and U9680 (N_9680,N_9438,N_9445);
nand U9681 (N_9681,N_9285,N_9452);
xor U9682 (N_9682,N_9267,N_9311);
xnor U9683 (N_9683,N_9469,N_9386);
or U9684 (N_9684,N_9432,N_9372);
nand U9685 (N_9685,N_9486,N_9317);
nor U9686 (N_9686,N_9333,N_9408);
xor U9687 (N_9687,N_9267,N_9305);
nor U9688 (N_9688,N_9350,N_9329);
xnor U9689 (N_9689,N_9276,N_9397);
nor U9690 (N_9690,N_9283,N_9489);
or U9691 (N_9691,N_9262,N_9495);
nand U9692 (N_9692,N_9299,N_9477);
nor U9693 (N_9693,N_9306,N_9451);
and U9694 (N_9694,N_9347,N_9440);
or U9695 (N_9695,N_9284,N_9428);
nor U9696 (N_9696,N_9417,N_9255);
xor U9697 (N_9697,N_9354,N_9434);
nor U9698 (N_9698,N_9345,N_9330);
nand U9699 (N_9699,N_9497,N_9431);
and U9700 (N_9700,N_9463,N_9453);
nand U9701 (N_9701,N_9493,N_9314);
xor U9702 (N_9702,N_9265,N_9294);
and U9703 (N_9703,N_9327,N_9326);
xnor U9704 (N_9704,N_9434,N_9379);
and U9705 (N_9705,N_9407,N_9305);
xnor U9706 (N_9706,N_9259,N_9499);
nand U9707 (N_9707,N_9280,N_9405);
nand U9708 (N_9708,N_9420,N_9288);
nor U9709 (N_9709,N_9410,N_9496);
and U9710 (N_9710,N_9492,N_9464);
xor U9711 (N_9711,N_9422,N_9429);
nand U9712 (N_9712,N_9328,N_9434);
nand U9713 (N_9713,N_9488,N_9490);
xor U9714 (N_9714,N_9451,N_9348);
xnor U9715 (N_9715,N_9435,N_9275);
and U9716 (N_9716,N_9333,N_9416);
nand U9717 (N_9717,N_9450,N_9466);
nand U9718 (N_9718,N_9255,N_9476);
or U9719 (N_9719,N_9467,N_9446);
nor U9720 (N_9720,N_9430,N_9408);
and U9721 (N_9721,N_9376,N_9439);
xnor U9722 (N_9722,N_9440,N_9296);
nor U9723 (N_9723,N_9414,N_9442);
nor U9724 (N_9724,N_9334,N_9491);
nand U9725 (N_9725,N_9397,N_9437);
and U9726 (N_9726,N_9348,N_9265);
nand U9727 (N_9727,N_9452,N_9282);
nor U9728 (N_9728,N_9250,N_9414);
xor U9729 (N_9729,N_9349,N_9435);
xor U9730 (N_9730,N_9392,N_9448);
or U9731 (N_9731,N_9444,N_9369);
or U9732 (N_9732,N_9457,N_9451);
or U9733 (N_9733,N_9386,N_9429);
nand U9734 (N_9734,N_9434,N_9458);
xnor U9735 (N_9735,N_9411,N_9268);
or U9736 (N_9736,N_9356,N_9496);
xnor U9737 (N_9737,N_9377,N_9425);
or U9738 (N_9738,N_9257,N_9468);
xor U9739 (N_9739,N_9320,N_9463);
nor U9740 (N_9740,N_9472,N_9318);
xor U9741 (N_9741,N_9265,N_9316);
and U9742 (N_9742,N_9250,N_9365);
and U9743 (N_9743,N_9487,N_9262);
xor U9744 (N_9744,N_9441,N_9277);
nand U9745 (N_9745,N_9364,N_9332);
nor U9746 (N_9746,N_9443,N_9404);
nor U9747 (N_9747,N_9270,N_9454);
nor U9748 (N_9748,N_9468,N_9323);
or U9749 (N_9749,N_9383,N_9350);
and U9750 (N_9750,N_9543,N_9611);
and U9751 (N_9751,N_9707,N_9538);
and U9752 (N_9752,N_9731,N_9725);
xor U9753 (N_9753,N_9522,N_9510);
nand U9754 (N_9754,N_9667,N_9527);
nor U9755 (N_9755,N_9741,N_9629);
xnor U9756 (N_9756,N_9672,N_9593);
or U9757 (N_9757,N_9519,N_9564);
or U9758 (N_9758,N_9625,N_9682);
or U9759 (N_9759,N_9563,N_9653);
nor U9760 (N_9760,N_9681,N_9709);
xnor U9761 (N_9761,N_9525,N_9701);
nand U9762 (N_9762,N_9665,N_9640);
or U9763 (N_9763,N_9670,N_9738);
and U9764 (N_9764,N_9680,N_9536);
nand U9765 (N_9765,N_9506,N_9679);
or U9766 (N_9766,N_9746,N_9717);
nor U9767 (N_9767,N_9696,N_9704);
and U9768 (N_9768,N_9555,N_9643);
nor U9769 (N_9769,N_9561,N_9677);
and U9770 (N_9770,N_9617,N_9609);
xor U9771 (N_9771,N_9657,N_9652);
nor U9772 (N_9772,N_9509,N_9719);
nand U9773 (N_9773,N_9548,N_9631);
nand U9774 (N_9774,N_9579,N_9708);
nor U9775 (N_9775,N_9650,N_9624);
nor U9776 (N_9776,N_9596,N_9539);
and U9777 (N_9777,N_9688,N_9637);
xnor U9778 (N_9778,N_9645,N_9549);
nand U9779 (N_9779,N_9711,N_9571);
and U9780 (N_9780,N_9545,N_9520);
and U9781 (N_9781,N_9675,N_9605);
xnor U9782 (N_9782,N_9556,N_9621);
and U9783 (N_9783,N_9595,N_9697);
and U9784 (N_9784,N_9695,N_9619);
and U9785 (N_9785,N_9546,N_9511);
nor U9786 (N_9786,N_9505,N_9674);
nand U9787 (N_9787,N_9602,N_9534);
nor U9788 (N_9788,N_9736,N_9633);
xor U9789 (N_9789,N_9531,N_9698);
and U9790 (N_9790,N_9582,N_9636);
and U9791 (N_9791,N_9713,N_9504);
or U9792 (N_9792,N_9668,N_9634);
or U9793 (N_9793,N_9692,N_9607);
nand U9794 (N_9794,N_9568,N_9591);
xnor U9795 (N_9795,N_9739,N_9723);
nor U9796 (N_9796,N_9676,N_9661);
or U9797 (N_9797,N_9612,N_9554);
xnor U9798 (N_9798,N_9603,N_9550);
nor U9799 (N_9799,N_9533,N_9663);
xor U9800 (N_9800,N_9716,N_9649);
nor U9801 (N_9801,N_9671,N_9655);
nand U9802 (N_9802,N_9678,N_9669);
nor U9803 (N_9803,N_9647,N_9518);
xnor U9804 (N_9804,N_9574,N_9687);
and U9805 (N_9805,N_9508,N_9702);
nor U9806 (N_9806,N_9620,N_9608);
nand U9807 (N_9807,N_9748,N_9628);
and U9808 (N_9808,N_9515,N_9623);
xnor U9809 (N_9809,N_9552,N_9714);
or U9810 (N_9810,N_9632,N_9584);
and U9811 (N_9811,N_9642,N_9635);
or U9812 (N_9812,N_9566,N_9613);
nand U9813 (N_9813,N_9513,N_9659);
nand U9814 (N_9814,N_9706,N_9565);
nand U9815 (N_9815,N_9700,N_9598);
nand U9816 (N_9816,N_9516,N_9727);
nand U9817 (N_9817,N_9654,N_9673);
xnor U9818 (N_9818,N_9614,N_9502);
nor U9819 (N_9819,N_9604,N_9600);
xor U9820 (N_9820,N_9537,N_9583);
xnor U9821 (N_9821,N_9587,N_9630);
nor U9822 (N_9822,N_9588,N_9572);
nand U9823 (N_9823,N_9622,N_9526);
xor U9824 (N_9824,N_9733,N_9724);
and U9825 (N_9825,N_9589,N_9599);
and U9826 (N_9826,N_9562,N_9710);
or U9827 (N_9827,N_9734,N_9745);
and U9828 (N_9828,N_9573,N_9646);
or U9829 (N_9829,N_9524,N_9729);
nor U9830 (N_9830,N_9627,N_9742);
or U9831 (N_9831,N_9581,N_9744);
xnor U9832 (N_9832,N_9594,N_9683);
nand U9833 (N_9833,N_9641,N_9703);
or U9834 (N_9834,N_9610,N_9666);
or U9835 (N_9835,N_9658,N_9530);
xnor U9836 (N_9836,N_9521,N_9626);
nor U9837 (N_9837,N_9644,N_9656);
nor U9838 (N_9838,N_9523,N_9535);
nand U9839 (N_9839,N_9732,N_9540);
xor U9840 (N_9840,N_9586,N_9615);
or U9841 (N_9841,N_9567,N_9560);
nand U9842 (N_9842,N_9576,N_9722);
xor U9843 (N_9843,N_9662,N_9551);
and U9844 (N_9844,N_9693,N_9570);
xor U9845 (N_9845,N_9514,N_9749);
nor U9846 (N_9846,N_9684,N_9639);
and U9847 (N_9847,N_9721,N_9686);
nand U9848 (N_9848,N_9712,N_9720);
nand U9849 (N_9849,N_9705,N_9507);
nand U9850 (N_9850,N_9694,N_9569);
nand U9851 (N_9851,N_9606,N_9726);
xnor U9852 (N_9852,N_9638,N_9578);
xnor U9853 (N_9853,N_9580,N_9699);
nand U9854 (N_9854,N_9528,N_9648);
nor U9855 (N_9855,N_9553,N_9715);
and U9856 (N_9856,N_9743,N_9740);
and U9857 (N_9857,N_9737,N_9660);
nand U9858 (N_9858,N_9532,N_9590);
and U9859 (N_9859,N_9689,N_9577);
or U9860 (N_9860,N_9547,N_9651);
xor U9861 (N_9861,N_9690,N_9541);
nand U9862 (N_9862,N_9585,N_9747);
and U9863 (N_9863,N_9575,N_9735);
nand U9864 (N_9864,N_9542,N_9529);
or U9865 (N_9865,N_9558,N_9685);
xor U9866 (N_9866,N_9601,N_9616);
nor U9867 (N_9867,N_9544,N_9503);
xor U9868 (N_9868,N_9618,N_9559);
and U9869 (N_9869,N_9592,N_9501);
xnor U9870 (N_9870,N_9728,N_9500);
or U9871 (N_9871,N_9691,N_9730);
nand U9872 (N_9872,N_9718,N_9597);
xnor U9873 (N_9873,N_9517,N_9557);
nor U9874 (N_9874,N_9664,N_9512);
and U9875 (N_9875,N_9526,N_9671);
and U9876 (N_9876,N_9664,N_9570);
or U9877 (N_9877,N_9713,N_9727);
or U9878 (N_9878,N_9564,N_9609);
nand U9879 (N_9879,N_9600,N_9677);
xor U9880 (N_9880,N_9678,N_9521);
xor U9881 (N_9881,N_9700,N_9654);
or U9882 (N_9882,N_9538,N_9522);
nand U9883 (N_9883,N_9708,N_9569);
and U9884 (N_9884,N_9746,N_9599);
nor U9885 (N_9885,N_9731,N_9647);
xnor U9886 (N_9886,N_9671,N_9511);
or U9887 (N_9887,N_9723,N_9720);
xor U9888 (N_9888,N_9531,N_9657);
xnor U9889 (N_9889,N_9640,N_9634);
xor U9890 (N_9890,N_9675,N_9742);
xnor U9891 (N_9891,N_9596,N_9512);
nor U9892 (N_9892,N_9510,N_9616);
xor U9893 (N_9893,N_9545,N_9631);
nand U9894 (N_9894,N_9530,N_9583);
nor U9895 (N_9895,N_9662,N_9533);
nor U9896 (N_9896,N_9609,N_9654);
and U9897 (N_9897,N_9568,N_9631);
nand U9898 (N_9898,N_9736,N_9536);
xor U9899 (N_9899,N_9639,N_9611);
nor U9900 (N_9900,N_9593,N_9666);
nand U9901 (N_9901,N_9648,N_9577);
nor U9902 (N_9902,N_9532,N_9630);
xor U9903 (N_9903,N_9612,N_9671);
nor U9904 (N_9904,N_9576,N_9686);
or U9905 (N_9905,N_9621,N_9720);
or U9906 (N_9906,N_9557,N_9631);
nor U9907 (N_9907,N_9631,N_9694);
xor U9908 (N_9908,N_9688,N_9568);
and U9909 (N_9909,N_9696,N_9568);
or U9910 (N_9910,N_9645,N_9686);
and U9911 (N_9911,N_9607,N_9558);
or U9912 (N_9912,N_9503,N_9513);
nor U9913 (N_9913,N_9612,N_9512);
xnor U9914 (N_9914,N_9733,N_9721);
nand U9915 (N_9915,N_9712,N_9730);
and U9916 (N_9916,N_9512,N_9600);
xor U9917 (N_9917,N_9592,N_9587);
and U9918 (N_9918,N_9736,N_9618);
nand U9919 (N_9919,N_9572,N_9540);
or U9920 (N_9920,N_9599,N_9549);
and U9921 (N_9921,N_9699,N_9513);
xnor U9922 (N_9922,N_9671,N_9708);
nand U9923 (N_9923,N_9567,N_9540);
and U9924 (N_9924,N_9605,N_9635);
or U9925 (N_9925,N_9556,N_9733);
xnor U9926 (N_9926,N_9620,N_9693);
xnor U9927 (N_9927,N_9520,N_9732);
or U9928 (N_9928,N_9501,N_9558);
nand U9929 (N_9929,N_9680,N_9700);
or U9930 (N_9930,N_9729,N_9731);
or U9931 (N_9931,N_9712,N_9704);
nand U9932 (N_9932,N_9566,N_9678);
nand U9933 (N_9933,N_9723,N_9707);
nand U9934 (N_9934,N_9677,N_9688);
nor U9935 (N_9935,N_9662,N_9588);
or U9936 (N_9936,N_9518,N_9625);
nor U9937 (N_9937,N_9599,N_9722);
nor U9938 (N_9938,N_9672,N_9642);
nor U9939 (N_9939,N_9667,N_9748);
xor U9940 (N_9940,N_9585,N_9693);
or U9941 (N_9941,N_9566,N_9747);
or U9942 (N_9942,N_9524,N_9603);
and U9943 (N_9943,N_9613,N_9546);
or U9944 (N_9944,N_9618,N_9543);
nand U9945 (N_9945,N_9613,N_9518);
nor U9946 (N_9946,N_9512,N_9695);
nand U9947 (N_9947,N_9571,N_9594);
xnor U9948 (N_9948,N_9724,N_9571);
or U9949 (N_9949,N_9672,N_9572);
nand U9950 (N_9950,N_9740,N_9523);
or U9951 (N_9951,N_9568,N_9531);
or U9952 (N_9952,N_9563,N_9716);
xor U9953 (N_9953,N_9670,N_9584);
xor U9954 (N_9954,N_9643,N_9557);
and U9955 (N_9955,N_9558,N_9667);
and U9956 (N_9956,N_9739,N_9551);
nand U9957 (N_9957,N_9610,N_9572);
and U9958 (N_9958,N_9679,N_9674);
xnor U9959 (N_9959,N_9501,N_9694);
xor U9960 (N_9960,N_9707,N_9617);
and U9961 (N_9961,N_9504,N_9620);
or U9962 (N_9962,N_9680,N_9734);
or U9963 (N_9963,N_9542,N_9512);
and U9964 (N_9964,N_9627,N_9544);
nand U9965 (N_9965,N_9744,N_9517);
nor U9966 (N_9966,N_9692,N_9687);
nor U9967 (N_9967,N_9702,N_9631);
xor U9968 (N_9968,N_9521,N_9614);
or U9969 (N_9969,N_9595,N_9530);
nor U9970 (N_9970,N_9530,N_9522);
nand U9971 (N_9971,N_9504,N_9506);
or U9972 (N_9972,N_9551,N_9532);
nand U9973 (N_9973,N_9705,N_9740);
or U9974 (N_9974,N_9536,N_9748);
and U9975 (N_9975,N_9569,N_9653);
or U9976 (N_9976,N_9666,N_9526);
and U9977 (N_9977,N_9506,N_9619);
or U9978 (N_9978,N_9679,N_9655);
nor U9979 (N_9979,N_9562,N_9614);
nor U9980 (N_9980,N_9606,N_9719);
nand U9981 (N_9981,N_9650,N_9677);
or U9982 (N_9982,N_9683,N_9739);
nand U9983 (N_9983,N_9625,N_9545);
nor U9984 (N_9984,N_9605,N_9734);
or U9985 (N_9985,N_9533,N_9670);
or U9986 (N_9986,N_9575,N_9729);
nand U9987 (N_9987,N_9584,N_9669);
nand U9988 (N_9988,N_9648,N_9711);
nor U9989 (N_9989,N_9712,N_9710);
and U9990 (N_9990,N_9631,N_9671);
and U9991 (N_9991,N_9527,N_9511);
xor U9992 (N_9992,N_9506,N_9590);
and U9993 (N_9993,N_9657,N_9625);
and U9994 (N_9994,N_9524,N_9670);
xnor U9995 (N_9995,N_9561,N_9678);
and U9996 (N_9996,N_9637,N_9723);
nand U9997 (N_9997,N_9704,N_9509);
nand U9998 (N_9998,N_9707,N_9721);
nor U9999 (N_9999,N_9633,N_9560);
nand U10000 (N_10000,N_9957,N_9823);
nor U10001 (N_10001,N_9894,N_9886);
nand U10002 (N_10002,N_9786,N_9842);
and U10003 (N_10003,N_9963,N_9775);
nor U10004 (N_10004,N_9929,N_9960);
or U10005 (N_10005,N_9897,N_9954);
and U10006 (N_10006,N_9759,N_9757);
nor U10007 (N_10007,N_9896,N_9989);
or U10008 (N_10008,N_9812,N_9750);
nor U10009 (N_10009,N_9755,N_9903);
nand U10010 (N_10010,N_9943,N_9876);
or U10011 (N_10011,N_9922,N_9843);
or U10012 (N_10012,N_9888,N_9931);
nand U10013 (N_10013,N_9904,N_9820);
xor U10014 (N_10014,N_9814,N_9821);
and U10015 (N_10015,N_9793,N_9999);
or U10016 (N_10016,N_9867,N_9794);
xnor U10017 (N_10017,N_9774,N_9981);
xor U10018 (N_10018,N_9968,N_9908);
nor U10019 (N_10019,N_9866,N_9836);
xor U10020 (N_10020,N_9780,N_9972);
or U10021 (N_10021,N_9785,N_9958);
or U10022 (N_10022,N_9875,N_9781);
or U10023 (N_10023,N_9884,N_9829);
nand U10024 (N_10024,N_9770,N_9984);
nand U10025 (N_10025,N_9782,N_9801);
nor U10026 (N_10026,N_9964,N_9760);
nand U10027 (N_10027,N_9863,N_9990);
nor U10028 (N_10028,N_9927,N_9764);
nor U10029 (N_10029,N_9913,N_9811);
nor U10030 (N_10030,N_9864,N_9763);
or U10031 (N_10031,N_9859,N_9877);
xnor U10032 (N_10032,N_9838,N_9965);
xor U10033 (N_10033,N_9840,N_9880);
xor U10034 (N_10034,N_9911,N_9878);
or U10035 (N_10035,N_9830,N_9998);
and U10036 (N_10036,N_9806,N_9895);
nand U10037 (N_10037,N_9887,N_9817);
xor U10038 (N_10038,N_9994,N_9848);
nor U10039 (N_10039,N_9892,N_9826);
nand U10040 (N_10040,N_9905,N_9874);
nand U10041 (N_10041,N_9756,N_9967);
xnor U10042 (N_10042,N_9799,N_9940);
nand U10043 (N_10043,N_9765,N_9945);
and U10044 (N_10044,N_9899,N_9844);
xor U10045 (N_10045,N_9815,N_9856);
and U10046 (N_10046,N_9810,N_9752);
xnor U10047 (N_10047,N_9991,N_9850);
nor U10048 (N_10048,N_9979,N_9930);
xnor U10049 (N_10049,N_9949,N_9795);
nor U10050 (N_10050,N_9798,N_9937);
nor U10051 (N_10051,N_9819,N_9831);
or U10052 (N_10052,N_9925,N_9946);
nand U10053 (N_10053,N_9805,N_9813);
nand U10054 (N_10054,N_9800,N_9824);
and U10055 (N_10055,N_9753,N_9973);
and U10056 (N_10056,N_9947,N_9993);
and U10057 (N_10057,N_9769,N_9906);
xnor U10058 (N_10058,N_9807,N_9825);
nor U10059 (N_10059,N_9898,N_9851);
nor U10060 (N_10060,N_9861,N_9822);
nor U10061 (N_10061,N_9766,N_9935);
nand U10062 (N_10062,N_9865,N_9910);
or U10063 (N_10063,N_9772,N_9862);
xnor U10064 (N_10064,N_9783,N_9996);
nand U10065 (N_10065,N_9939,N_9789);
and U10066 (N_10066,N_9995,N_9771);
and U10067 (N_10067,N_9849,N_9852);
nand U10068 (N_10068,N_9751,N_9902);
nand U10069 (N_10069,N_9966,N_9928);
xor U10070 (N_10070,N_9917,N_9776);
xor U10071 (N_10071,N_9941,N_9816);
xor U10072 (N_10072,N_9952,N_9882);
xor U10073 (N_10073,N_9959,N_9970);
and U10074 (N_10074,N_9983,N_9881);
or U10075 (N_10075,N_9953,N_9845);
xor U10076 (N_10076,N_9767,N_9942);
and U10077 (N_10077,N_9944,N_9901);
and U10078 (N_10078,N_9961,N_9857);
nor U10079 (N_10079,N_9969,N_9950);
or U10080 (N_10080,N_9841,N_9986);
nand U10081 (N_10081,N_9914,N_9985);
nor U10082 (N_10082,N_9883,N_9974);
xnor U10083 (N_10083,N_9915,N_9871);
nor U10084 (N_10084,N_9992,N_9853);
or U10085 (N_10085,N_9962,N_9846);
nor U10086 (N_10086,N_9988,N_9761);
nand U10087 (N_10087,N_9923,N_9936);
xor U10088 (N_10088,N_9938,N_9854);
nor U10089 (N_10089,N_9885,N_9919);
or U10090 (N_10090,N_9797,N_9920);
nor U10091 (N_10091,N_9997,N_9855);
or U10092 (N_10092,N_9933,N_9890);
or U10093 (N_10093,N_9790,N_9987);
nor U10094 (N_10094,N_9900,N_9879);
or U10095 (N_10095,N_9909,N_9872);
xnor U10096 (N_10096,N_9976,N_9833);
nand U10097 (N_10097,N_9934,N_9791);
and U10098 (N_10098,N_9768,N_9932);
nand U10099 (N_10099,N_9982,N_9924);
nor U10100 (N_10100,N_9828,N_9796);
and U10101 (N_10101,N_9977,N_9834);
xnor U10102 (N_10102,N_9773,N_9907);
nand U10103 (N_10103,N_9778,N_9948);
nor U10104 (N_10104,N_9870,N_9792);
nor U10105 (N_10105,N_9980,N_9847);
nand U10106 (N_10106,N_9978,N_9777);
xor U10107 (N_10107,N_9837,N_9912);
and U10108 (N_10108,N_9802,N_9832);
and U10109 (N_10109,N_9758,N_9762);
xor U10110 (N_10110,N_9893,N_9860);
and U10111 (N_10111,N_9889,N_9975);
or U10112 (N_10112,N_9779,N_9891);
and U10113 (N_10113,N_9808,N_9955);
or U10114 (N_10114,N_9754,N_9916);
nand U10115 (N_10115,N_9951,N_9827);
or U10116 (N_10116,N_9818,N_9809);
or U10117 (N_10117,N_9804,N_9956);
and U10118 (N_10118,N_9971,N_9926);
nand U10119 (N_10119,N_9788,N_9835);
nor U10120 (N_10120,N_9873,N_9918);
and U10121 (N_10121,N_9839,N_9858);
and U10122 (N_10122,N_9868,N_9784);
nor U10123 (N_10123,N_9921,N_9787);
nor U10124 (N_10124,N_9803,N_9869);
nand U10125 (N_10125,N_9923,N_9948);
nand U10126 (N_10126,N_9815,N_9783);
nor U10127 (N_10127,N_9767,N_9765);
or U10128 (N_10128,N_9782,N_9915);
nor U10129 (N_10129,N_9800,N_9825);
or U10130 (N_10130,N_9774,N_9937);
and U10131 (N_10131,N_9989,N_9980);
or U10132 (N_10132,N_9757,N_9887);
xnor U10133 (N_10133,N_9819,N_9938);
nand U10134 (N_10134,N_9888,N_9868);
and U10135 (N_10135,N_9845,N_9782);
or U10136 (N_10136,N_9933,N_9917);
xor U10137 (N_10137,N_9758,N_9797);
or U10138 (N_10138,N_9820,N_9795);
nand U10139 (N_10139,N_9817,N_9852);
or U10140 (N_10140,N_9991,N_9780);
and U10141 (N_10141,N_9842,N_9885);
nand U10142 (N_10142,N_9959,N_9861);
or U10143 (N_10143,N_9923,N_9905);
or U10144 (N_10144,N_9941,N_9783);
nand U10145 (N_10145,N_9986,N_9945);
nor U10146 (N_10146,N_9968,N_9762);
nand U10147 (N_10147,N_9803,N_9793);
nand U10148 (N_10148,N_9802,N_9781);
xor U10149 (N_10149,N_9890,N_9829);
xnor U10150 (N_10150,N_9854,N_9848);
nand U10151 (N_10151,N_9940,N_9771);
and U10152 (N_10152,N_9933,N_9756);
nor U10153 (N_10153,N_9847,N_9992);
xnor U10154 (N_10154,N_9988,N_9781);
nand U10155 (N_10155,N_9813,N_9822);
or U10156 (N_10156,N_9818,N_9771);
xor U10157 (N_10157,N_9920,N_9932);
or U10158 (N_10158,N_9839,N_9868);
or U10159 (N_10159,N_9870,N_9966);
or U10160 (N_10160,N_9915,N_9828);
or U10161 (N_10161,N_9941,N_9775);
and U10162 (N_10162,N_9941,N_9953);
nand U10163 (N_10163,N_9931,N_9764);
or U10164 (N_10164,N_9783,N_9864);
nor U10165 (N_10165,N_9987,N_9808);
or U10166 (N_10166,N_9947,N_9835);
nand U10167 (N_10167,N_9832,N_9902);
nand U10168 (N_10168,N_9814,N_9975);
nand U10169 (N_10169,N_9790,N_9972);
and U10170 (N_10170,N_9793,N_9868);
nor U10171 (N_10171,N_9860,N_9802);
xnor U10172 (N_10172,N_9878,N_9750);
nor U10173 (N_10173,N_9818,N_9950);
nand U10174 (N_10174,N_9805,N_9904);
or U10175 (N_10175,N_9781,N_9819);
nand U10176 (N_10176,N_9798,N_9942);
xor U10177 (N_10177,N_9788,N_9967);
and U10178 (N_10178,N_9889,N_9757);
and U10179 (N_10179,N_9981,N_9851);
and U10180 (N_10180,N_9794,N_9886);
and U10181 (N_10181,N_9990,N_9958);
nand U10182 (N_10182,N_9994,N_9976);
or U10183 (N_10183,N_9854,N_9835);
nand U10184 (N_10184,N_9842,N_9886);
or U10185 (N_10185,N_9785,N_9871);
and U10186 (N_10186,N_9870,N_9773);
and U10187 (N_10187,N_9881,N_9905);
or U10188 (N_10188,N_9964,N_9767);
or U10189 (N_10189,N_9761,N_9876);
or U10190 (N_10190,N_9962,N_9990);
nand U10191 (N_10191,N_9962,N_9958);
or U10192 (N_10192,N_9894,N_9881);
nand U10193 (N_10193,N_9911,N_9769);
or U10194 (N_10194,N_9867,N_9970);
or U10195 (N_10195,N_9807,N_9913);
or U10196 (N_10196,N_9910,N_9936);
nor U10197 (N_10197,N_9947,N_9898);
nor U10198 (N_10198,N_9953,N_9965);
xnor U10199 (N_10199,N_9895,N_9873);
or U10200 (N_10200,N_9924,N_9958);
xor U10201 (N_10201,N_9995,N_9846);
xor U10202 (N_10202,N_9823,N_9800);
or U10203 (N_10203,N_9893,N_9983);
or U10204 (N_10204,N_9878,N_9915);
or U10205 (N_10205,N_9851,N_9950);
nand U10206 (N_10206,N_9922,N_9982);
xor U10207 (N_10207,N_9875,N_9816);
or U10208 (N_10208,N_9848,N_9806);
nor U10209 (N_10209,N_9775,N_9872);
or U10210 (N_10210,N_9905,N_9909);
nand U10211 (N_10211,N_9963,N_9885);
nor U10212 (N_10212,N_9925,N_9818);
nand U10213 (N_10213,N_9871,N_9825);
and U10214 (N_10214,N_9773,N_9815);
nor U10215 (N_10215,N_9868,N_9918);
and U10216 (N_10216,N_9996,N_9867);
nand U10217 (N_10217,N_9870,N_9896);
and U10218 (N_10218,N_9753,N_9891);
nand U10219 (N_10219,N_9919,N_9985);
or U10220 (N_10220,N_9823,N_9903);
xor U10221 (N_10221,N_9809,N_9910);
xor U10222 (N_10222,N_9812,N_9937);
xnor U10223 (N_10223,N_9932,N_9890);
and U10224 (N_10224,N_9846,N_9851);
or U10225 (N_10225,N_9887,N_9752);
nand U10226 (N_10226,N_9815,N_9763);
nand U10227 (N_10227,N_9948,N_9821);
xnor U10228 (N_10228,N_9917,N_9894);
nor U10229 (N_10229,N_9845,N_9893);
xnor U10230 (N_10230,N_9811,N_9983);
nor U10231 (N_10231,N_9861,N_9855);
nand U10232 (N_10232,N_9971,N_9768);
nand U10233 (N_10233,N_9929,N_9950);
nand U10234 (N_10234,N_9997,N_9992);
nand U10235 (N_10235,N_9985,N_9955);
and U10236 (N_10236,N_9852,N_9844);
xor U10237 (N_10237,N_9767,N_9993);
and U10238 (N_10238,N_9932,N_9939);
or U10239 (N_10239,N_9928,N_9850);
xnor U10240 (N_10240,N_9895,N_9768);
xor U10241 (N_10241,N_9766,N_9902);
or U10242 (N_10242,N_9796,N_9773);
xnor U10243 (N_10243,N_9906,N_9863);
nor U10244 (N_10244,N_9889,N_9936);
nand U10245 (N_10245,N_9845,N_9938);
nor U10246 (N_10246,N_9906,N_9952);
xor U10247 (N_10247,N_9818,N_9912);
nand U10248 (N_10248,N_9870,N_9854);
nand U10249 (N_10249,N_9889,N_9927);
or U10250 (N_10250,N_10057,N_10248);
xor U10251 (N_10251,N_10209,N_10079);
nand U10252 (N_10252,N_10063,N_10151);
xnor U10253 (N_10253,N_10080,N_10033);
nor U10254 (N_10254,N_10246,N_10152);
or U10255 (N_10255,N_10093,N_10125);
xnor U10256 (N_10256,N_10201,N_10116);
or U10257 (N_10257,N_10249,N_10181);
and U10258 (N_10258,N_10010,N_10208);
or U10259 (N_10259,N_10081,N_10190);
nand U10260 (N_10260,N_10068,N_10122);
or U10261 (N_10261,N_10043,N_10003);
or U10262 (N_10262,N_10051,N_10013);
and U10263 (N_10263,N_10184,N_10217);
nor U10264 (N_10264,N_10180,N_10126);
or U10265 (N_10265,N_10089,N_10048);
and U10266 (N_10266,N_10117,N_10189);
xnor U10267 (N_10267,N_10045,N_10206);
xor U10268 (N_10268,N_10225,N_10019);
or U10269 (N_10269,N_10243,N_10215);
and U10270 (N_10270,N_10034,N_10064);
nor U10271 (N_10271,N_10077,N_10127);
xnor U10272 (N_10272,N_10224,N_10071);
and U10273 (N_10273,N_10046,N_10024);
or U10274 (N_10274,N_10195,N_10168);
nand U10275 (N_10275,N_10037,N_10247);
nand U10276 (N_10276,N_10076,N_10171);
and U10277 (N_10277,N_10192,N_10001);
xor U10278 (N_10278,N_10053,N_10166);
xor U10279 (N_10279,N_10022,N_10227);
xor U10280 (N_10280,N_10176,N_10005);
and U10281 (N_10281,N_10109,N_10169);
or U10282 (N_10282,N_10060,N_10017);
and U10283 (N_10283,N_10238,N_10000);
and U10284 (N_10284,N_10009,N_10092);
nand U10285 (N_10285,N_10244,N_10058);
xor U10286 (N_10286,N_10062,N_10015);
xor U10287 (N_10287,N_10229,N_10197);
nand U10288 (N_10288,N_10101,N_10183);
nand U10289 (N_10289,N_10200,N_10014);
and U10290 (N_10290,N_10030,N_10136);
nand U10291 (N_10291,N_10237,N_10012);
nand U10292 (N_10292,N_10090,N_10061);
nand U10293 (N_10293,N_10226,N_10102);
and U10294 (N_10294,N_10099,N_10194);
or U10295 (N_10295,N_10210,N_10055);
xor U10296 (N_10296,N_10170,N_10235);
or U10297 (N_10297,N_10230,N_10039);
nand U10298 (N_10298,N_10145,N_10065);
nor U10299 (N_10299,N_10028,N_10158);
nor U10300 (N_10300,N_10026,N_10214);
xor U10301 (N_10301,N_10198,N_10148);
or U10302 (N_10302,N_10044,N_10207);
nor U10303 (N_10303,N_10111,N_10199);
and U10304 (N_10304,N_10231,N_10123);
and U10305 (N_10305,N_10203,N_10149);
nand U10306 (N_10306,N_10016,N_10234);
xnor U10307 (N_10307,N_10031,N_10175);
and U10308 (N_10308,N_10173,N_10160);
or U10309 (N_10309,N_10054,N_10113);
nor U10310 (N_10310,N_10202,N_10134);
and U10311 (N_10311,N_10094,N_10107);
nor U10312 (N_10312,N_10032,N_10082);
and U10313 (N_10313,N_10172,N_10029);
or U10314 (N_10314,N_10002,N_10018);
and U10315 (N_10315,N_10241,N_10132);
nor U10316 (N_10316,N_10066,N_10050);
and U10317 (N_10317,N_10219,N_10072);
and U10318 (N_10318,N_10213,N_10073);
nor U10319 (N_10319,N_10228,N_10139);
or U10320 (N_10320,N_10130,N_10085);
nor U10321 (N_10321,N_10167,N_10159);
or U10322 (N_10322,N_10087,N_10097);
nor U10323 (N_10323,N_10008,N_10040);
nand U10324 (N_10324,N_10236,N_10163);
and U10325 (N_10325,N_10133,N_10147);
and U10326 (N_10326,N_10186,N_10174);
and U10327 (N_10327,N_10144,N_10021);
or U10328 (N_10328,N_10155,N_10075);
and U10329 (N_10329,N_10059,N_10154);
and U10330 (N_10330,N_10185,N_10041);
and U10331 (N_10331,N_10020,N_10129);
and U10332 (N_10332,N_10086,N_10100);
or U10333 (N_10333,N_10156,N_10232);
xnor U10334 (N_10334,N_10191,N_10162);
or U10335 (N_10335,N_10143,N_10178);
nor U10336 (N_10336,N_10083,N_10118);
nor U10337 (N_10337,N_10146,N_10193);
xor U10338 (N_10338,N_10011,N_10177);
and U10339 (N_10339,N_10096,N_10205);
nor U10340 (N_10340,N_10035,N_10153);
and U10341 (N_10341,N_10220,N_10131);
and U10342 (N_10342,N_10074,N_10098);
xnor U10343 (N_10343,N_10135,N_10188);
and U10344 (N_10344,N_10070,N_10218);
nand U10345 (N_10345,N_10137,N_10165);
nor U10346 (N_10346,N_10119,N_10142);
or U10347 (N_10347,N_10036,N_10006);
and U10348 (N_10348,N_10179,N_10222);
xor U10349 (N_10349,N_10182,N_10239);
or U10350 (N_10350,N_10157,N_10124);
or U10351 (N_10351,N_10106,N_10067);
xor U10352 (N_10352,N_10088,N_10120);
nand U10353 (N_10353,N_10084,N_10052);
or U10354 (N_10354,N_10161,N_10056);
nor U10355 (N_10355,N_10128,N_10027);
xor U10356 (N_10356,N_10138,N_10242);
xnor U10357 (N_10357,N_10115,N_10038);
or U10358 (N_10358,N_10187,N_10108);
or U10359 (N_10359,N_10141,N_10078);
nand U10360 (N_10360,N_10140,N_10114);
or U10361 (N_10361,N_10164,N_10221);
and U10362 (N_10362,N_10196,N_10204);
or U10363 (N_10363,N_10047,N_10240);
nor U10364 (N_10364,N_10007,N_10069);
or U10365 (N_10365,N_10212,N_10105);
and U10366 (N_10366,N_10004,N_10110);
nor U10367 (N_10367,N_10023,N_10233);
and U10368 (N_10368,N_10025,N_10245);
nand U10369 (N_10369,N_10049,N_10216);
nand U10370 (N_10370,N_10121,N_10091);
nor U10371 (N_10371,N_10042,N_10095);
nor U10372 (N_10372,N_10104,N_10211);
xnor U10373 (N_10373,N_10112,N_10103);
nor U10374 (N_10374,N_10150,N_10223);
and U10375 (N_10375,N_10142,N_10216);
or U10376 (N_10376,N_10145,N_10102);
nor U10377 (N_10377,N_10179,N_10076);
nand U10378 (N_10378,N_10179,N_10067);
nor U10379 (N_10379,N_10157,N_10237);
nor U10380 (N_10380,N_10202,N_10080);
xor U10381 (N_10381,N_10056,N_10037);
nor U10382 (N_10382,N_10056,N_10214);
or U10383 (N_10383,N_10007,N_10246);
nand U10384 (N_10384,N_10073,N_10191);
nand U10385 (N_10385,N_10092,N_10186);
nor U10386 (N_10386,N_10225,N_10233);
xor U10387 (N_10387,N_10042,N_10207);
and U10388 (N_10388,N_10147,N_10094);
nand U10389 (N_10389,N_10233,N_10135);
nor U10390 (N_10390,N_10008,N_10031);
nor U10391 (N_10391,N_10119,N_10019);
and U10392 (N_10392,N_10206,N_10115);
and U10393 (N_10393,N_10025,N_10032);
nand U10394 (N_10394,N_10204,N_10210);
xor U10395 (N_10395,N_10085,N_10001);
or U10396 (N_10396,N_10140,N_10166);
nor U10397 (N_10397,N_10081,N_10114);
nor U10398 (N_10398,N_10146,N_10215);
and U10399 (N_10399,N_10092,N_10073);
and U10400 (N_10400,N_10026,N_10119);
nand U10401 (N_10401,N_10066,N_10023);
xor U10402 (N_10402,N_10049,N_10050);
nor U10403 (N_10403,N_10194,N_10138);
nand U10404 (N_10404,N_10177,N_10150);
xnor U10405 (N_10405,N_10132,N_10175);
xnor U10406 (N_10406,N_10075,N_10148);
or U10407 (N_10407,N_10003,N_10202);
and U10408 (N_10408,N_10122,N_10019);
nand U10409 (N_10409,N_10157,N_10049);
nor U10410 (N_10410,N_10148,N_10040);
nand U10411 (N_10411,N_10042,N_10181);
xor U10412 (N_10412,N_10007,N_10107);
xnor U10413 (N_10413,N_10027,N_10000);
and U10414 (N_10414,N_10016,N_10118);
nor U10415 (N_10415,N_10124,N_10103);
nand U10416 (N_10416,N_10136,N_10231);
nand U10417 (N_10417,N_10248,N_10100);
and U10418 (N_10418,N_10015,N_10054);
and U10419 (N_10419,N_10149,N_10108);
or U10420 (N_10420,N_10222,N_10053);
nand U10421 (N_10421,N_10043,N_10012);
nand U10422 (N_10422,N_10011,N_10232);
xor U10423 (N_10423,N_10059,N_10094);
or U10424 (N_10424,N_10037,N_10185);
or U10425 (N_10425,N_10094,N_10125);
or U10426 (N_10426,N_10238,N_10202);
nand U10427 (N_10427,N_10052,N_10161);
and U10428 (N_10428,N_10097,N_10233);
nand U10429 (N_10429,N_10181,N_10199);
nor U10430 (N_10430,N_10098,N_10030);
xor U10431 (N_10431,N_10142,N_10097);
and U10432 (N_10432,N_10078,N_10133);
xnor U10433 (N_10433,N_10120,N_10196);
xnor U10434 (N_10434,N_10064,N_10161);
and U10435 (N_10435,N_10024,N_10154);
nor U10436 (N_10436,N_10237,N_10027);
nand U10437 (N_10437,N_10106,N_10240);
nor U10438 (N_10438,N_10221,N_10084);
or U10439 (N_10439,N_10229,N_10193);
nor U10440 (N_10440,N_10074,N_10217);
nor U10441 (N_10441,N_10193,N_10209);
or U10442 (N_10442,N_10090,N_10018);
nor U10443 (N_10443,N_10081,N_10206);
nand U10444 (N_10444,N_10056,N_10102);
and U10445 (N_10445,N_10070,N_10025);
and U10446 (N_10446,N_10239,N_10044);
nor U10447 (N_10447,N_10039,N_10241);
nand U10448 (N_10448,N_10119,N_10077);
nor U10449 (N_10449,N_10105,N_10113);
and U10450 (N_10450,N_10185,N_10197);
nor U10451 (N_10451,N_10006,N_10096);
and U10452 (N_10452,N_10085,N_10076);
xor U10453 (N_10453,N_10140,N_10025);
xnor U10454 (N_10454,N_10110,N_10234);
xor U10455 (N_10455,N_10059,N_10213);
nor U10456 (N_10456,N_10002,N_10009);
nor U10457 (N_10457,N_10039,N_10015);
and U10458 (N_10458,N_10025,N_10088);
and U10459 (N_10459,N_10200,N_10033);
or U10460 (N_10460,N_10047,N_10050);
nor U10461 (N_10461,N_10245,N_10219);
nand U10462 (N_10462,N_10129,N_10113);
nor U10463 (N_10463,N_10005,N_10218);
nand U10464 (N_10464,N_10116,N_10107);
xnor U10465 (N_10465,N_10128,N_10133);
nand U10466 (N_10466,N_10023,N_10089);
nand U10467 (N_10467,N_10185,N_10071);
or U10468 (N_10468,N_10011,N_10055);
nor U10469 (N_10469,N_10228,N_10016);
xnor U10470 (N_10470,N_10046,N_10217);
nor U10471 (N_10471,N_10054,N_10044);
nor U10472 (N_10472,N_10032,N_10040);
nand U10473 (N_10473,N_10040,N_10130);
and U10474 (N_10474,N_10070,N_10092);
or U10475 (N_10475,N_10119,N_10073);
nand U10476 (N_10476,N_10043,N_10194);
nand U10477 (N_10477,N_10244,N_10114);
and U10478 (N_10478,N_10187,N_10106);
or U10479 (N_10479,N_10216,N_10241);
xor U10480 (N_10480,N_10074,N_10134);
and U10481 (N_10481,N_10049,N_10042);
xor U10482 (N_10482,N_10197,N_10148);
nand U10483 (N_10483,N_10198,N_10107);
nor U10484 (N_10484,N_10204,N_10186);
nor U10485 (N_10485,N_10060,N_10171);
xnor U10486 (N_10486,N_10211,N_10173);
nand U10487 (N_10487,N_10191,N_10220);
or U10488 (N_10488,N_10184,N_10236);
nor U10489 (N_10489,N_10199,N_10035);
or U10490 (N_10490,N_10003,N_10248);
and U10491 (N_10491,N_10079,N_10094);
nor U10492 (N_10492,N_10169,N_10093);
xor U10493 (N_10493,N_10073,N_10176);
xor U10494 (N_10494,N_10139,N_10099);
xnor U10495 (N_10495,N_10068,N_10059);
and U10496 (N_10496,N_10022,N_10179);
or U10497 (N_10497,N_10154,N_10248);
and U10498 (N_10498,N_10021,N_10033);
nor U10499 (N_10499,N_10143,N_10187);
nor U10500 (N_10500,N_10298,N_10274);
or U10501 (N_10501,N_10339,N_10285);
nand U10502 (N_10502,N_10445,N_10322);
nand U10503 (N_10503,N_10379,N_10428);
or U10504 (N_10504,N_10453,N_10390);
nor U10505 (N_10505,N_10438,N_10296);
nand U10506 (N_10506,N_10257,N_10260);
nor U10507 (N_10507,N_10334,N_10469);
and U10508 (N_10508,N_10487,N_10336);
nand U10509 (N_10509,N_10278,N_10488);
nor U10510 (N_10510,N_10429,N_10407);
nor U10511 (N_10511,N_10493,N_10251);
nand U10512 (N_10512,N_10434,N_10343);
or U10513 (N_10513,N_10270,N_10495);
and U10514 (N_10514,N_10290,N_10464);
and U10515 (N_10515,N_10333,N_10399);
nand U10516 (N_10516,N_10395,N_10315);
xor U10517 (N_10517,N_10371,N_10338);
and U10518 (N_10518,N_10389,N_10484);
and U10519 (N_10519,N_10358,N_10344);
xnor U10520 (N_10520,N_10300,N_10346);
and U10521 (N_10521,N_10277,N_10430);
or U10522 (N_10522,N_10314,N_10326);
xor U10523 (N_10523,N_10268,N_10366);
or U10524 (N_10524,N_10446,N_10448);
nor U10525 (N_10525,N_10347,N_10293);
nor U10526 (N_10526,N_10377,N_10450);
nand U10527 (N_10527,N_10312,N_10266);
nand U10528 (N_10528,N_10352,N_10310);
nor U10529 (N_10529,N_10396,N_10265);
nor U10530 (N_10530,N_10282,N_10345);
or U10531 (N_10531,N_10421,N_10332);
xor U10532 (N_10532,N_10378,N_10455);
xor U10533 (N_10533,N_10404,N_10294);
or U10534 (N_10534,N_10423,N_10289);
nor U10535 (N_10535,N_10485,N_10409);
nor U10536 (N_10536,N_10305,N_10292);
or U10537 (N_10537,N_10427,N_10324);
or U10538 (N_10538,N_10309,N_10476);
xnor U10539 (N_10539,N_10380,N_10307);
nand U10540 (N_10540,N_10359,N_10436);
nor U10541 (N_10541,N_10462,N_10481);
or U10542 (N_10542,N_10330,N_10443);
nand U10543 (N_10543,N_10400,N_10325);
xnor U10544 (N_10544,N_10480,N_10454);
and U10545 (N_10545,N_10348,N_10317);
xor U10546 (N_10546,N_10386,N_10483);
nor U10547 (N_10547,N_10273,N_10272);
nor U10548 (N_10548,N_10468,N_10375);
xor U10549 (N_10549,N_10350,N_10320);
xnor U10550 (N_10550,N_10303,N_10362);
or U10551 (N_10551,N_10417,N_10431);
nand U10552 (N_10552,N_10406,N_10308);
nor U10553 (N_10553,N_10313,N_10280);
and U10554 (N_10554,N_10439,N_10490);
xnor U10555 (N_10555,N_10281,N_10318);
nor U10556 (N_10556,N_10424,N_10287);
nor U10557 (N_10557,N_10381,N_10460);
or U10558 (N_10558,N_10466,N_10369);
and U10559 (N_10559,N_10496,N_10271);
xor U10560 (N_10560,N_10323,N_10403);
and U10561 (N_10561,N_10269,N_10327);
or U10562 (N_10562,N_10349,N_10306);
xnor U10563 (N_10563,N_10385,N_10321);
xnor U10564 (N_10564,N_10444,N_10373);
xnor U10565 (N_10565,N_10367,N_10295);
and U10566 (N_10566,N_10452,N_10478);
and U10567 (N_10567,N_10405,N_10372);
nor U10568 (N_10568,N_10471,N_10420);
or U10569 (N_10569,N_10284,N_10252);
and U10570 (N_10570,N_10393,N_10254);
xnor U10571 (N_10571,N_10475,N_10384);
nor U10572 (N_10572,N_10456,N_10250);
nor U10573 (N_10573,N_10412,N_10276);
or U10574 (N_10574,N_10382,N_10337);
nand U10575 (N_10575,N_10474,N_10442);
nand U10576 (N_10576,N_10392,N_10357);
or U10577 (N_10577,N_10360,N_10457);
nor U10578 (N_10578,N_10401,N_10340);
and U10579 (N_10579,N_10451,N_10311);
and U10580 (N_10580,N_10368,N_10447);
or U10581 (N_10581,N_10433,N_10255);
or U10582 (N_10582,N_10408,N_10365);
and U10583 (N_10583,N_10440,N_10353);
or U10584 (N_10584,N_10477,N_10482);
nor U10585 (N_10585,N_10256,N_10473);
nor U10586 (N_10586,N_10414,N_10465);
and U10587 (N_10587,N_10370,N_10263);
xnor U10588 (N_10588,N_10275,N_10301);
nor U10589 (N_10589,N_10302,N_10398);
nor U10590 (N_10590,N_10264,N_10329);
and U10591 (N_10591,N_10472,N_10467);
nand U10592 (N_10592,N_10286,N_10288);
and U10593 (N_10593,N_10498,N_10459);
and U10594 (N_10594,N_10435,N_10383);
and U10595 (N_10595,N_10463,N_10486);
or U10596 (N_10596,N_10391,N_10397);
nand U10597 (N_10597,N_10432,N_10413);
or U10598 (N_10598,N_10253,N_10425);
xor U10599 (N_10599,N_10267,N_10497);
and U10600 (N_10600,N_10394,N_10388);
and U10601 (N_10601,N_10470,N_10416);
nand U10602 (N_10602,N_10262,N_10494);
nor U10603 (N_10603,N_10363,N_10328);
nor U10604 (N_10604,N_10341,N_10316);
xor U10605 (N_10605,N_10279,N_10355);
and U10606 (N_10606,N_10331,N_10335);
xnor U10607 (N_10607,N_10479,N_10491);
and U10608 (N_10608,N_10437,N_10492);
or U10609 (N_10609,N_10402,N_10356);
nand U10610 (N_10610,N_10304,N_10449);
and U10611 (N_10611,N_10259,N_10426);
xor U10612 (N_10612,N_10342,N_10376);
or U10613 (N_10613,N_10261,N_10411);
or U10614 (N_10614,N_10489,N_10364);
nand U10615 (N_10615,N_10351,N_10458);
and U10616 (N_10616,N_10410,N_10415);
and U10617 (N_10617,N_10387,N_10374);
or U10618 (N_10618,N_10361,N_10319);
nand U10619 (N_10619,N_10297,N_10419);
and U10620 (N_10620,N_10499,N_10283);
or U10621 (N_10621,N_10418,N_10422);
nand U10622 (N_10622,N_10354,N_10461);
nor U10623 (N_10623,N_10299,N_10291);
or U10624 (N_10624,N_10441,N_10258);
and U10625 (N_10625,N_10313,N_10375);
nand U10626 (N_10626,N_10407,N_10349);
xnor U10627 (N_10627,N_10471,N_10466);
and U10628 (N_10628,N_10263,N_10322);
xor U10629 (N_10629,N_10279,N_10367);
nor U10630 (N_10630,N_10268,N_10353);
and U10631 (N_10631,N_10472,N_10295);
nor U10632 (N_10632,N_10338,N_10274);
and U10633 (N_10633,N_10339,N_10275);
xor U10634 (N_10634,N_10361,N_10263);
and U10635 (N_10635,N_10452,N_10434);
nand U10636 (N_10636,N_10250,N_10259);
nor U10637 (N_10637,N_10466,N_10375);
nand U10638 (N_10638,N_10453,N_10291);
and U10639 (N_10639,N_10330,N_10259);
xnor U10640 (N_10640,N_10350,N_10296);
nor U10641 (N_10641,N_10313,N_10494);
xor U10642 (N_10642,N_10390,N_10385);
and U10643 (N_10643,N_10465,N_10380);
or U10644 (N_10644,N_10329,N_10303);
nor U10645 (N_10645,N_10448,N_10472);
nand U10646 (N_10646,N_10339,N_10327);
xnor U10647 (N_10647,N_10449,N_10400);
and U10648 (N_10648,N_10299,N_10418);
nand U10649 (N_10649,N_10297,N_10427);
nor U10650 (N_10650,N_10405,N_10335);
xor U10651 (N_10651,N_10281,N_10446);
xnor U10652 (N_10652,N_10328,N_10480);
and U10653 (N_10653,N_10265,N_10363);
nor U10654 (N_10654,N_10286,N_10457);
or U10655 (N_10655,N_10469,N_10438);
nand U10656 (N_10656,N_10352,N_10442);
nand U10657 (N_10657,N_10358,N_10479);
nand U10658 (N_10658,N_10484,N_10436);
and U10659 (N_10659,N_10453,N_10432);
and U10660 (N_10660,N_10473,N_10420);
or U10661 (N_10661,N_10288,N_10267);
or U10662 (N_10662,N_10389,N_10255);
or U10663 (N_10663,N_10276,N_10478);
and U10664 (N_10664,N_10379,N_10392);
and U10665 (N_10665,N_10407,N_10427);
xor U10666 (N_10666,N_10470,N_10289);
and U10667 (N_10667,N_10377,N_10415);
nor U10668 (N_10668,N_10425,N_10488);
and U10669 (N_10669,N_10291,N_10367);
or U10670 (N_10670,N_10287,N_10364);
and U10671 (N_10671,N_10423,N_10370);
xor U10672 (N_10672,N_10449,N_10450);
or U10673 (N_10673,N_10268,N_10365);
and U10674 (N_10674,N_10313,N_10351);
xnor U10675 (N_10675,N_10461,N_10284);
or U10676 (N_10676,N_10274,N_10325);
nor U10677 (N_10677,N_10462,N_10422);
nor U10678 (N_10678,N_10495,N_10257);
or U10679 (N_10679,N_10391,N_10291);
nand U10680 (N_10680,N_10434,N_10362);
xnor U10681 (N_10681,N_10361,N_10304);
or U10682 (N_10682,N_10361,N_10339);
or U10683 (N_10683,N_10388,N_10436);
nand U10684 (N_10684,N_10320,N_10308);
xnor U10685 (N_10685,N_10374,N_10436);
and U10686 (N_10686,N_10460,N_10345);
and U10687 (N_10687,N_10291,N_10290);
or U10688 (N_10688,N_10419,N_10381);
nand U10689 (N_10689,N_10475,N_10479);
or U10690 (N_10690,N_10259,N_10347);
xor U10691 (N_10691,N_10459,N_10257);
xnor U10692 (N_10692,N_10476,N_10380);
xor U10693 (N_10693,N_10310,N_10477);
and U10694 (N_10694,N_10474,N_10277);
xor U10695 (N_10695,N_10250,N_10404);
nand U10696 (N_10696,N_10352,N_10313);
nand U10697 (N_10697,N_10254,N_10302);
xor U10698 (N_10698,N_10434,N_10421);
or U10699 (N_10699,N_10458,N_10260);
xor U10700 (N_10700,N_10355,N_10291);
xor U10701 (N_10701,N_10323,N_10424);
and U10702 (N_10702,N_10295,N_10420);
xnor U10703 (N_10703,N_10307,N_10486);
xor U10704 (N_10704,N_10438,N_10431);
xor U10705 (N_10705,N_10449,N_10388);
nand U10706 (N_10706,N_10255,N_10328);
or U10707 (N_10707,N_10377,N_10407);
nor U10708 (N_10708,N_10314,N_10388);
nand U10709 (N_10709,N_10260,N_10407);
nand U10710 (N_10710,N_10445,N_10266);
and U10711 (N_10711,N_10294,N_10375);
nand U10712 (N_10712,N_10260,N_10310);
and U10713 (N_10713,N_10375,N_10401);
xnor U10714 (N_10714,N_10402,N_10482);
xor U10715 (N_10715,N_10372,N_10282);
and U10716 (N_10716,N_10353,N_10406);
xnor U10717 (N_10717,N_10436,N_10368);
or U10718 (N_10718,N_10256,N_10396);
and U10719 (N_10719,N_10329,N_10392);
xnor U10720 (N_10720,N_10271,N_10423);
xnor U10721 (N_10721,N_10375,N_10261);
nand U10722 (N_10722,N_10336,N_10497);
and U10723 (N_10723,N_10303,N_10308);
nand U10724 (N_10724,N_10461,N_10396);
nor U10725 (N_10725,N_10294,N_10252);
nor U10726 (N_10726,N_10305,N_10463);
xor U10727 (N_10727,N_10266,N_10355);
nor U10728 (N_10728,N_10332,N_10393);
or U10729 (N_10729,N_10393,N_10369);
nor U10730 (N_10730,N_10490,N_10467);
nor U10731 (N_10731,N_10427,N_10264);
and U10732 (N_10732,N_10398,N_10291);
xor U10733 (N_10733,N_10266,N_10444);
and U10734 (N_10734,N_10384,N_10430);
nand U10735 (N_10735,N_10360,N_10495);
xnor U10736 (N_10736,N_10463,N_10391);
and U10737 (N_10737,N_10274,N_10484);
nand U10738 (N_10738,N_10407,N_10461);
xnor U10739 (N_10739,N_10410,N_10253);
or U10740 (N_10740,N_10469,N_10278);
nor U10741 (N_10741,N_10290,N_10423);
or U10742 (N_10742,N_10308,N_10425);
or U10743 (N_10743,N_10370,N_10482);
xor U10744 (N_10744,N_10446,N_10428);
xnor U10745 (N_10745,N_10493,N_10495);
nand U10746 (N_10746,N_10329,N_10311);
or U10747 (N_10747,N_10312,N_10349);
nand U10748 (N_10748,N_10345,N_10495);
nor U10749 (N_10749,N_10396,N_10324);
and U10750 (N_10750,N_10630,N_10666);
and U10751 (N_10751,N_10622,N_10637);
xor U10752 (N_10752,N_10639,N_10620);
nand U10753 (N_10753,N_10506,N_10669);
nand U10754 (N_10754,N_10655,N_10540);
or U10755 (N_10755,N_10709,N_10707);
nand U10756 (N_10756,N_10665,N_10522);
xor U10757 (N_10757,N_10698,N_10582);
and U10758 (N_10758,N_10534,N_10573);
nor U10759 (N_10759,N_10725,N_10724);
or U10760 (N_10760,N_10696,N_10531);
nor U10761 (N_10761,N_10528,N_10502);
and U10762 (N_10762,N_10689,N_10570);
or U10763 (N_10763,N_10694,N_10626);
nand U10764 (N_10764,N_10608,N_10541);
or U10765 (N_10765,N_10663,N_10642);
or U10766 (N_10766,N_10635,N_10623);
or U10767 (N_10767,N_10564,N_10688);
nand U10768 (N_10768,N_10566,N_10735);
nand U10769 (N_10769,N_10731,N_10656);
xor U10770 (N_10770,N_10682,N_10511);
nor U10771 (N_10771,N_10543,N_10593);
xor U10772 (N_10772,N_10744,N_10599);
nor U10773 (N_10773,N_10662,N_10590);
or U10774 (N_10774,N_10537,N_10624);
nor U10775 (N_10775,N_10523,N_10684);
nand U10776 (N_10776,N_10733,N_10602);
xor U10777 (N_10777,N_10697,N_10551);
nand U10778 (N_10778,N_10548,N_10578);
nor U10779 (N_10779,N_10649,N_10546);
nor U10780 (N_10780,N_10644,N_10743);
nor U10781 (N_10781,N_10587,N_10618);
or U10782 (N_10782,N_10596,N_10518);
xnor U10783 (N_10783,N_10636,N_10706);
and U10784 (N_10784,N_10640,N_10520);
or U10785 (N_10785,N_10521,N_10585);
or U10786 (N_10786,N_10509,N_10650);
nor U10787 (N_10787,N_10519,N_10653);
or U10788 (N_10788,N_10609,N_10686);
or U10789 (N_10789,N_10503,N_10514);
nand U10790 (N_10790,N_10710,N_10500);
and U10791 (N_10791,N_10695,N_10621);
or U10792 (N_10792,N_10749,N_10678);
nand U10793 (N_10793,N_10536,N_10673);
and U10794 (N_10794,N_10579,N_10533);
or U10795 (N_10795,N_10571,N_10687);
nand U10796 (N_10796,N_10577,N_10638);
and U10797 (N_10797,N_10512,N_10614);
nand U10798 (N_10798,N_10646,N_10616);
and U10799 (N_10799,N_10713,N_10691);
nand U10800 (N_10800,N_10722,N_10595);
xor U10801 (N_10801,N_10535,N_10561);
xnor U10802 (N_10802,N_10584,N_10741);
nand U10803 (N_10803,N_10704,N_10544);
nand U10804 (N_10804,N_10591,N_10538);
or U10805 (N_10805,N_10726,N_10729);
and U10806 (N_10806,N_10658,N_10607);
nor U10807 (N_10807,N_10668,N_10586);
nand U10808 (N_10808,N_10738,N_10554);
or U10809 (N_10809,N_10734,N_10723);
xnor U10810 (N_10810,N_10661,N_10671);
nor U10811 (N_10811,N_10746,N_10574);
nand U10812 (N_10812,N_10603,N_10700);
nor U10813 (N_10813,N_10601,N_10712);
and U10814 (N_10814,N_10513,N_10632);
nor U10815 (N_10815,N_10575,N_10606);
or U10816 (N_10816,N_10641,N_10745);
nand U10817 (N_10817,N_10501,N_10627);
and U10818 (N_10818,N_10631,N_10702);
or U10819 (N_10819,N_10711,N_10556);
and U10820 (N_10820,N_10597,N_10679);
xor U10821 (N_10821,N_10718,N_10605);
xor U10822 (N_10822,N_10598,N_10742);
and U10823 (N_10823,N_10549,N_10716);
and U10824 (N_10824,N_10659,N_10550);
or U10825 (N_10825,N_10516,N_10558);
and U10826 (N_10826,N_10651,N_10563);
nor U10827 (N_10827,N_10730,N_10714);
or U10828 (N_10828,N_10553,N_10562);
nor U10829 (N_10829,N_10736,N_10545);
xor U10830 (N_10830,N_10611,N_10510);
nand U10831 (N_10831,N_10705,N_10505);
or U10832 (N_10832,N_10727,N_10654);
xor U10833 (N_10833,N_10555,N_10628);
nand U10834 (N_10834,N_10625,N_10542);
and U10835 (N_10835,N_10660,N_10748);
or U10836 (N_10836,N_10643,N_10667);
nor U10837 (N_10837,N_10615,N_10581);
and U10838 (N_10838,N_10670,N_10715);
nor U10839 (N_10839,N_10692,N_10634);
or U10840 (N_10840,N_10672,N_10674);
xnor U10841 (N_10841,N_10721,N_10708);
or U10842 (N_10842,N_10703,N_10530);
nor U10843 (N_10843,N_10675,N_10592);
and U10844 (N_10844,N_10645,N_10676);
nor U10845 (N_10845,N_10612,N_10588);
and U10846 (N_10846,N_10560,N_10629);
nor U10847 (N_10847,N_10677,N_10600);
xor U10848 (N_10848,N_10610,N_10525);
or U10849 (N_10849,N_10604,N_10685);
and U10850 (N_10850,N_10527,N_10580);
xor U10851 (N_10851,N_10594,N_10693);
nor U10852 (N_10852,N_10529,N_10683);
nand U10853 (N_10853,N_10717,N_10532);
nor U10854 (N_10854,N_10701,N_10664);
nand U10855 (N_10855,N_10583,N_10547);
or U10856 (N_10856,N_10613,N_10504);
nor U10857 (N_10857,N_10539,N_10567);
nor U10858 (N_10858,N_10747,N_10740);
nand U10859 (N_10859,N_10633,N_10576);
or U10860 (N_10860,N_10719,N_10732);
or U10861 (N_10861,N_10681,N_10559);
and U10862 (N_10862,N_10647,N_10552);
nor U10863 (N_10863,N_10508,N_10515);
nand U10864 (N_10864,N_10524,N_10680);
xor U10865 (N_10865,N_10565,N_10507);
and U10866 (N_10866,N_10728,N_10657);
xnor U10867 (N_10867,N_10617,N_10737);
nor U10868 (N_10868,N_10589,N_10568);
nor U10869 (N_10869,N_10648,N_10690);
xor U10870 (N_10870,N_10572,N_10619);
and U10871 (N_10871,N_10699,N_10526);
or U10872 (N_10872,N_10557,N_10569);
xor U10873 (N_10873,N_10739,N_10517);
xnor U10874 (N_10874,N_10720,N_10652);
or U10875 (N_10875,N_10734,N_10552);
or U10876 (N_10876,N_10531,N_10690);
nand U10877 (N_10877,N_10532,N_10538);
nand U10878 (N_10878,N_10749,N_10680);
nand U10879 (N_10879,N_10624,N_10649);
xnor U10880 (N_10880,N_10674,N_10694);
xor U10881 (N_10881,N_10677,N_10607);
nor U10882 (N_10882,N_10658,N_10695);
or U10883 (N_10883,N_10541,N_10701);
nand U10884 (N_10884,N_10630,N_10540);
nand U10885 (N_10885,N_10721,N_10687);
nand U10886 (N_10886,N_10600,N_10602);
nor U10887 (N_10887,N_10723,N_10712);
or U10888 (N_10888,N_10503,N_10502);
nor U10889 (N_10889,N_10720,N_10512);
nand U10890 (N_10890,N_10545,N_10653);
xor U10891 (N_10891,N_10589,N_10544);
or U10892 (N_10892,N_10539,N_10661);
and U10893 (N_10893,N_10525,N_10513);
or U10894 (N_10894,N_10650,N_10645);
and U10895 (N_10895,N_10671,N_10685);
or U10896 (N_10896,N_10706,N_10624);
or U10897 (N_10897,N_10587,N_10603);
nand U10898 (N_10898,N_10671,N_10520);
nor U10899 (N_10899,N_10730,N_10614);
or U10900 (N_10900,N_10689,N_10548);
or U10901 (N_10901,N_10553,N_10594);
or U10902 (N_10902,N_10596,N_10682);
xnor U10903 (N_10903,N_10504,N_10561);
xor U10904 (N_10904,N_10611,N_10514);
or U10905 (N_10905,N_10689,N_10635);
nor U10906 (N_10906,N_10560,N_10594);
nor U10907 (N_10907,N_10593,N_10599);
or U10908 (N_10908,N_10573,N_10667);
or U10909 (N_10909,N_10502,N_10642);
xor U10910 (N_10910,N_10569,N_10603);
xnor U10911 (N_10911,N_10510,N_10730);
nor U10912 (N_10912,N_10564,N_10580);
xor U10913 (N_10913,N_10504,N_10699);
or U10914 (N_10914,N_10501,N_10559);
nor U10915 (N_10915,N_10747,N_10688);
or U10916 (N_10916,N_10676,N_10691);
xor U10917 (N_10917,N_10685,N_10654);
and U10918 (N_10918,N_10631,N_10725);
and U10919 (N_10919,N_10573,N_10624);
or U10920 (N_10920,N_10717,N_10536);
and U10921 (N_10921,N_10509,N_10668);
and U10922 (N_10922,N_10621,N_10693);
nor U10923 (N_10923,N_10512,N_10677);
or U10924 (N_10924,N_10522,N_10588);
nor U10925 (N_10925,N_10623,N_10588);
nor U10926 (N_10926,N_10730,N_10557);
nand U10927 (N_10927,N_10668,N_10712);
xor U10928 (N_10928,N_10710,N_10637);
and U10929 (N_10929,N_10741,N_10643);
xnor U10930 (N_10930,N_10511,N_10501);
nor U10931 (N_10931,N_10562,N_10616);
or U10932 (N_10932,N_10668,N_10673);
or U10933 (N_10933,N_10622,N_10567);
xnor U10934 (N_10934,N_10569,N_10700);
nor U10935 (N_10935,N_10510,N_10579);
nand U10936 (N_10936,N_10659,N_10505);
xor U10937 (N_10937,N_10517,N_10552);
nor U10938 (N_10938,N_10593,N_10606);
nand U10939 (N_10939,N_10621,N_10734);
and U10940 (N_10940,N_10638,N_10519);
nand U10941 (N_10941,N_10708,N_10527);
and U10942 (N_10942,N_10523,N_10572);
xor U10943 (N_10943,N_10617,N_10647);
xor U10944 (N_10944,N_10695,N_10571);
nand U10945 (N_10945,N_10692,N_10501);
nand U10946 (N_10946,N_10662,N_10655);
nand U10947 (N_10947,N_10677,N_10626);
and U10948 (N_10948,N_10500,N_10743);
xnor U10949 (N_10949,N_10583,N_10630);
nor U10950 (N_10950,N_10701,N_10517);
nor U10951 (N_10951,N_10662,N_10570);
or U10952 (N_10952,N_10550,N_10613);
and U10953 (N_10953,N_10733,N_10533);
or U10954 (N_10954,N_10550,N_10512);
or U10955 (N_10955,N_10737,N_10681);
xor U10956 (N_10956,N_10653,N_10735);
nor U10957 (N_10957,N_10627,N_10663);
xnor U10958 (N_10958,N_10530,N_10524);
nand U10959 (N_10959,N_10587,N_10548);
nand U10960 (N_10960,N_10741,N_10629);
nor U10961 (N_10961,N_10710,N_10522);
xnor U10962 (N_10962,N_10551,N_10669);
and U10963 (N_10963,N_10746,N_10614);
xor U10964 (N_10964,N_10717,N_10732);
and U10965 (N_10965,N_10658,N_10533);
xor U10966 (N_10966,N_10716,N_10746);
or U10967 (N_10967,N_10578,N_10564);
or U10968 (N_10968,N_10638,N_10596);
nand U10969 (N_10969,N_10607,N_10558);
and U10970 (N_10970,N_10748,N_10652);
nand U10971 (N_10971,N_10539,N_10714);
nand U10972 (N_10972,N_10680,N_10734);
xor U10973 (N_10973,N_10741,N_10709);
xor U10974 (N_10974,N_10736,N_10601);
or U10975 (N_10975,N_10643,N_10720);
and U10976 (N_10976,N_10614,N_10710);
or U10977 (N_10977,N_10572,N_10719);
nand U10978 (N_10978,N_10735,N_10730);
nand U10979 (N_10979,N_10595,N_10606);
xnor U10980 (N_10980,N_10658,N_10717);
nor U10981 (N_10981,N_10607,N_10613);
and U10982 (N_10982,N_10727,N_10741);
or U10983 (N_10983,N_10632,N_10532);
nand U10984 (N_10984,N_10500,N_10529);
or U10985 (N_10985,N_10504,N_10559);
nand U10986 (N_10986,N_10651,N_10702);
nand U10987 (N_10987,N_10540,N_10620);
nor U10988 (N_10988,N_10650,N_10651);
nor U10989 (N_10989,N_10583,N_10565);
xnor U10990 (N_10990,N_10595,N_10625);
nand U10991 (N_10991,N_10551,N_10656);
nor U10992 (N_10992,N_10539,N_10612);
nand U10993 (N_10993,N_10639,N_10656);
and U10994 (N_10994,N_10730,N_10715);
or U10995 (N_10995,N_10537,N_10619);
nor U10996 (N_10996,N_10690,N_10533);
or U10997 (N_10997,N_10688,N_10578);
and U10998 (N_10998,N_10728,N_10684);
nand U10999 (N_10999,N_10660,N_10686);
or U11000 (N_11000,N_10889,N_10878);
and U11001 (N_11001,N_10897,N_10998);
nand U11002 (N_11002,N_10996,N_10942);
nand U11003 (N_11003,N_10980,N_10890);
or U11004 (N_11004,N_10817,N_10814);
nor U11005 (N_11005,N_10805,N_10789);
nor U11006 (N_11006,N_10757,N_10908);
and U11007 (N_11007,N_10779,N_10915);
and U11008 (N_11008,N_10975,N_10948);
nor U11009 (N_11009,N_10967,N_10857);
xor U11010 (N_11010,N_10919,N_10794);
xor U11011 (N_11011,N_10963,N_10910);
or U11012 (N_11012,N_10846,N_10811);
nand U11013 (N_11013,N_10753,N_10952);
xor U11014 (N_11014,N_10966,N_10933);
nor U11015 (N_11015,N_10944,N_10797);
nor U11016 (N_11016,N_10860,N_10982);
nor U11017 (N_11017,N_10911,N_10901);
nor U11018 (N_11018,N_10988,N_10843);
xor U11019 (N_11019,N_10859,N_10761);
nand U11020 (N_11020,N_10804,N_10820);
nand U11021 (N_11021,N_10877,N_10812);
nand U11022 (N_11022,N_10993,N_10872);
and U11023 (N_11023,N_10882,N_10887);
and U11024 (N_11024,N_10973,N_10929);
nor U11025 (N_11025,N_10949,N_10997);
nand U11026 (N_11026,N_10918,N_10821);
xor U11027 (N_11027,N_10879,N_10864);
and U11028 (N_11028,N_10808,N_10880);
xor U11029 (N_11029,N_10909,N_10869);
nor U11030 (N_11030,N_10947,N_10835);
nand U11031 (N_11031,N_10928,N_10924);
nor U11032 (N_11032,N_10920,N_10953);
nand U11033 (N_11033,N_10981,N_10840);
xnor U11034 (N_11034,N_10867,N_10945);
or U11035 (N_11035,N_10940,N_10774);
or U11036 (N_11036,N_10800,N_10813);
nor U11037 (N_11037,N_10913,N_10976);
xnor U11038 (N_11038,N_10806,N_10772);
and U11039 (N_11039,N_10763,N_10755);
and U11040 (N_11040,N_10934,N_10831);
and U11041 (N_11041,N_10954,N_10905);
nand U11042 (N_11042,N_10781,N_10939);
xnor U11043 (N_11043,N_10810,N_10902);
or U11044 (N_11044,N_10799,N_10984);
xor U11045 (N_11045,N_10758,N_10932);
and U11046 (N_11046,N_10855,N_10906);
nor U11047 (N_11047,N_10844,N_10793);
xnor U11048 (N_11048,N_10828,N_10790);
and U11049 (N_11049,N_10865,N_10815);
xnor U11050 (N_11050,N_10788,N_10839);
xnor U11051 (N_11051,N_10778,N_10863);
and U11052 (N_11052,N_10816,N_10912);
and U11053 (N_11053,N_10930,N_10951);
and U11054 (N_11054,N_10782,N_10836);
xnor U11055 (N_11055,N_10979,N_10925);
nor U11056 (N_11056,N_10922,N_10965);
xor U11057 (N_11057,N_10837,N_10861);
and U11058 (N_11058,N_10892,N_10853);
and U11059 (N_11059,N_10950,N_10914);
or U11060 (N_11060,N_10756,N_10931);
nand U11061 (N_11061,N_10978,N_10783);
xor U11062 (N_11062,N_10900,N_10927);
and U11063 (N_11063,N_10983,N_10895);
and U11064 (N_11064,N_10956,N_10830);
xnor U11065 (N_11065,N_10856,N_10786);
or U11066 (N_11066,N_10868,N_10769);
or U11067 (N_11067,N_10896,N_10866);
and U11068 (N_11068,N_10992,N_10958);
nor U11069 (N_11069,N_10776,N_10935);
xnor U11070 (N_11070,N_10768,N_10970);
nand U11071 (N_11071,N_10893,N_10759);
and U11072 (N_11072,N_10990,N_10943);
and U11073 (N_11073,N_10750,N_10838);
xor U11074 (N_11074,N_10847,N_10824);
xnor U11075 (N_11075,N_10796,N_10876);
xor U11076 (N_11076,N_10850,N_10827);
nand U11077 (N_11077,N_10775,N_10891);
xnor U11078 (N_11078,N_10762,N_10849);
xnor U11079 (N_11079,N_10851,N_10926);
and U11080 (N_11080,N_10916,N_10936);
nor U11081 (N_11081,N_10941,N_10792);
or U11082 (N_11082,N_10767,N_10995);
xnor U11083 (N_11083,N_10968,N_10765);
and U11084 (N_11084,N_10964,N_10903);
xor U11085 (N_11085,N_10899,N_10818);
nor U11086 (N_11086,N_10751,N_10801);
or U11087 (N_11087,N_10957,N_10985);
and U11088 (N_11088,N_10784,N_10871);
or U11089 (N_11089,N_10807,N_10885);
xnor U11090 (N_11090,N_10795,N_10754);
or U11091 (N_11091,N_10766,N_10923);
xor U11092 (N_11092,N_10994,N_10907);
nand U11093 (N_11093,N_10852,N_10848);
xor U11094 (N_11094,N_10991,N_10946);
and U11095 (N_11095,N_10826,N_10986);
xor U11096 (N_11096,N_10832,N_10822);
and U11097 (N_11097,N_10842,N_10841);
nor U11098 (N_11098,N_10937,N_10969);
nor U11099 (N_11099,N_10787,N_10825);
xnor U11100 (N_11100,N_10752,N_10955);
and U11101 (N_11101,N_10862,N_10875);
nand U11102 (N_11102,N_10833,N_10764);
nor U11103 (N_11103,N_10834,N_10881);
nand U11104 (N_11104,N_10770,N_10972);
or U11105 (N_11105,N_10829,N_10858);
and U11106 (N_11106,N_10974,N_10999);
or U11107 (N_11107,N_10898,N_10886);
and U11108 (N_11108,N_10962,N_10960);
nand U11109 (N_11109,N_10780,N_10771);
nor U11110 (N_11110,N_10959,N_10873);
xor U11111 (N_11111,N_10971,N_10938);
nor U11112 (N_11112,N_10894,N_10917);
xor U11113 (N_11113,N_10823,N_10760);
nor U11114 (N_11114,N_10785,N_10883);
nand U11115 (N_11115,N_10803,N_10884);
and U11116 (N_11116,N_10904,N_10989);
and U11117 (N_11117,N_10854,N_10802);
nor U11118 (N_11118,N_10777,N_10977);
nor U11119 (N_11119,N_10809,N_10845);
nand U11120 (N_11120,N_10870,N_10773);
nand U11121 (N_11121,N_10888,N_10819);
and U11122 (N_11122,N_10791,N_10961);
nand U11123 (N_11123,N_10987,N_10798);
or U11124 (N_11124,N_10874,N_10921);
nor U11125 (N_11125,N_10862,N_10907);
and U11126 (N_11126,N_10951,N_10791);
and U11127 (N_11127,N_10811,N_10768);
xnor U11128 (N_11128,N_10912,N_10881);
nor U11129 (N_11129,N_10945,N_10840);
xnor U11130 (N_11130,N_10977,N_10750);
xnor U11131 (N_11131,N_10959,N_10901);
or U11132 (N_11132,N_10932,N_10778);
xor U11133 (N_11133,N_10755,N_10890);
nand U11134 (N_11134,N_10957,N_10781);
xor U11135 (N_11135,N_10919,N_10868);
nand U11136 (N_11136,N_10846,N_10966);
nand U11137 (N_11137,N_10798,N_10981);
or U11138 (N_11138,N_10994,N_10910);
xor U11139 (N_11139,N_10872,N_10870);
nand U11140 (N_11140,N_10964,N_10913);
and U11141 (N_11141,N_10907,N_10757);
nand U11142 (N_11142,N_10942,N_10865);
nand U11143 (N_11143,N_10883,N_10798);
nand U11144 (N_11144,N_10807,N_10888);
nor U11145 (N_11145,N_10841,N_10886);
and U11146 (N_11146,N_10981,N_10834);
xor U11147 (N_11147,N_10991,N_10963);
nand U11148 (N_11148,N_10780,N_10935);
or U11149 (N_11149,N_10803,N_10958);
nor U11150 (N_11150,N_10835,N_10996);
or U11151 (N_11151,N_10897,N_10759);
nand U11152 (N_11152,N_10980,N_10835);
nor U11153 (N_11153,N_10927,N_10946);
nand U11154 (N_11154,N_10838,N_10754);
xor U11155 (N_11155,N_10982,N_10820);
and U11156 (N_11156,N_10934,N_10914);
or U11157 (N_11157,N_10803,N_10757);
or U11158 (N_11158,N_10980,N_10960);
nand U11159 (N_11159,N_10778,N_10954);
nor U11160 (N_11160,N_10886,N_10863);
nand U11161 (N_11161,N_10868,N_10876);
and U11162 (N_11162,N_10807,N_10814);
xor U11163 (N_11163,N_10967,N_10916);
nor U11164 (N_11164,N_10784,N_10781);
or U11165 (N_11165,N_10798,N_10947);
nor U11166 (N_11166,N_10908,N_10986);
and U11167 (N_11167,N_10894,N_10818);
nor U11168 (N_11168,N_10902,N_10861);
and U11169 (N_11169,N_10854,N_10963);
and U11170 (N_11170,N_10825,N_10820);
or U11171 (N_11171,N_10756,N_10975);
xnor U11172 (N_11172,N_10877,N_10750);
and U11173 (N_11173,N_10908,N_10885);
nor U11174 (N_11174,N_10986,N_10888);
and U11175 (N_11175,N_10854,N_10887);
or U11176 (N_11176,N_10957,N_10915);
and U11177 (N_11177,N_10878,N_10947);
nand U11178 (N_11178,N_10931,N_10928);
or U11179 (N_11179,N_10837,N_10947);
or U11180 (N_11180,N_10766,N_10836);
nor U11181 (N_11181,N_10972,N_10926);
xor U11182 (N_11182,N_10973,N_10832);
or U11183 (N_11183,N_10795,N_10808);
nand U11184 (N_11184,N_10864,N_10905);
nor U11185 (N_11185,N_10874,N_10918);
nand U11186 (N_11186,N_10790,N_10998);
nand U11187 (N_11187,N_10865,N_10847);
or U11188 (N_11188,N_10793,N_10924);
and U11189 (N_11189,N_10976,N_10874);
xor U11190 (N_11190,N_10762,N_10974);
nor U11191 (N_11191,N_10787,N_10881);
or U11192 (N_11192,N_10835,N_10948);
or U11193 (N_11193,N_10841,N_10787);
and U11194 (N_11194,N_10928,N_10945);
and U11195 (N_11195,N_10796,N_10848);
xor U11196 (N_11196,N_10886,N_10933);
nor U11197 (N_11197,N_10806,N_10812);
nand U11198 (N_11198,N_10956,N_10954);
xor U11199 (N_11199,N_10847,N_10849);
nand U11200 (N_11200,N_10994,N_10975);
nand U11201 (N_11201,N_10980,N_10929);
nand U11202 (N_11202,N_10925,N_10918);
or U11203 (N_11203,N_10808,N_10778);
and U11204 (N_11204,N_10999,N_10799);
and U11205 (N_11205,N_10978,N_10774);
nor U11206 (N_11206,N_10756,N_10948);
nor U11207 (N_11207,N_10761,N_10796);
xor U11208 (N_11208,N_10857,N_10896);
or U11209 (N_11209,N_10829,N_10797);
or U11210 (N_11210,N_10800,N_10887);
or U11211 (N_11211,N_10790,N_10819);
xor U11212 (N_11212,N_10931,N_10943);
nand U11213 (N_11213,N_10840,N_10762);
or U11214 (N_11214,N_10874,N_10866);
xor U11215 (N_11215,N_10859,N_10976);
xnor U11216 (N_11216,N_10811,N_10866);
nand U11217 (N_11217,N_10769,N_10958);
nand U11218 (N_11218,N_10875,N_10955);
xnor U11219 (N_11219,N_10932,N_10975);
xnor U11220 (N_11220,N_10873,N_10865);
or U11221 (N_11221,N_10981,N_10883);
and U11222 (N_11222,N_10858,N_10884);
and U11223 (N_11223,N_10839,N_10794);
nor U11224 (N_11224,N_10911,N_10881);
or U11225 (N_11225,N_10771,N_10877);
and U11226 (N_11226,N_10860,N_10983);
xor U11227 (N_11227,N_10752,N_10998);
nand U11228 (N_11228,N_10896,N_10814);
nand U11229 (N_11229,N_10901,N_10988);
nand U11230 (N_11230,N_10987,N_10983);
or U11231 (N_11231,N_10789,N_10756);
xnor U11232 (N_11232,N_10840,N_10764);
nor U11233 (N_11233,N_10937,N_10931);
nand U11234 (N_11234,N_10997,N_10955);
xor U11235 (N_11235,N_10905,N_10899);
and U11236 (N_11236,N_10970,N_10790);
xnor U11237 (N_11237,N_10869,N_10812);
xor U11238 (N_11238,N_10981,N_10923);
xor U11239 (N_11239,N_10808,N_10904);
nor U11240 (N_11240,N_10816,N_10916);
or U11241 (N_11241,N_10793,N_10808);
nor U11242 (N_11242,N_10779,N_10973);
or U11243 (N_11243,N_10824,N_10904);
nand U11244 (N_11244,N_10898,N_10938);
nand U11245 (N_11245,N_10962,N_10996);
nand U11246 (N_11246,N_10858,N_10820);
nor U11247 (N_11247,N_10868,N_10927);
or U11248 (N_11248,N_10942,N_10994);
or U11249 (N_11249,N_10752,N_10834);
nand U11250 (N_11250,N_11236,N_11243);
or U11251 (N_11251,N_11216,N_11195);
or U11252 (N_11252,N_11217,N_11068);
and U11253 (N_11253,N_11039,N_11003);
xnor U11254 (N_11254,N_11072,N_11156);
nor U11255 (N_11255,N_11166,N_11038);
nor U11256 (N_11256,N_11170,N_11214);
xnor U11257 (N_11257,N_11103,N_11018);
or U11258 (N_11258,N_11054,N_11107);
or U11259 (N_11259,N_11143,N_11240);
and U11260 (N_11260,N_11129,N_11164);
nor U11261 (N_11261,N_11190,N_11248);
or U11262 (N_11262,N_11015,N_11050);
and U11263 (N_11263,N_11042,N_11029);
and U11264 (N_11264,N_11076,N_11008);
nor U11265 (N_11265,N_11056,N_11223);
or U11266 (N_11266,N_11004,N_11235);
and U11267 (N_11267,N_11144,N_11071);
xnor U11268 (N_11268,N_11041,N_11099);
nor U11269 (N_11269,N_11069,N_11090);
and U11270 (N_11270,N_11181,N_11180);
nand U11271 (N_11271,N_11220,N_11052);
nand U11272 (N_11272,N_11022,N_11086);
nor U11273 (N_11273,N_11043,N_11098);
or U11274 (N_11274,N_11080,N_11177);
nand U11275 (N_11275,N_11161,N_11158);
nand U11276 (N_11276,N_11231,N_11013);
or U11277 (N_11277,N_11058,N_11197);
or U11278 (N_11278,N_11233,N_11193);
or U11279 (N_11279,N_11153,N_11055);
nor U11280 (N_11280,N_11135,N_11051);
xor U11281 (N_11281,N_11152,N_11094);
nand U11282 (N_11282,N_11210,N_11067);
nor U11283 (N_11283,N_11082,N_11186);
or U11284 (N_11284,N_11200,N_11101);
nor U11285 (N_11285,N_11085,N_11053);
xnor U11286 (N_11286,N_11245,N_11035);
and U11287 (N_11287,N_11145,N_11062);
or U11288 (N_11288,N_11064,N_11215);
or U11289 (N_11289,N_11226,N_11081);
and U11290 (N_11290,N_11237,N_11118);
and U11291 (N_11291,N_11128,N_11212);
or U11292 (N_11292,N_11100,N_11205);
or U11293 (N_11293,N_11092,N_11155);
nand U11294 (N_11294,N_11136,N_11079);
nand U11295 (N_11295,N_11061,N_11012);
nor U11296 (N_11296,N_11218,N_11150);
nand U11297 (N_11297,N_11117,N_11060);
nor U11298 (N_11298,N_11154,N_11213);
xor U11299 (N_11299,N_11134,N_11110);
or U11300 (N_11300,N_11227,N_11083);
nor U11301 (N_11301,N_11221,N_11207);
xnor U11302 (N_11302,N_11165,N_11014);
xor U11303 (N_11303,N_11095,N_11203);
nand U11304 (N_11304,N_11025,N_11239);
or U11305 (N_11305,N_11077,N_11201);
nor U11306 (N_11306,N_11202,N_11066);
and U11307 (N_11307,N_11157,N_11183);
or U11308 (N_11308,N_11059,N_11057);
and U11309 (N_11309,N_11148,N_11078);
nand U11310 (N_11310,N_11074,N_11234);
xnor U11311 (N_11311,N_11106,N_11142);
nor U11312 (N_11312,N_11151,N_11232);
nor U11313 (N_11313,N_11019,N_11131);
nor U11314 (N_11314,N_11209,N_11088);
or U11315 (N_11315,N_11189,N_11000);
nand U11316 (N_11316,N_11208,N_11097);
and U11317 (N_11317,N_11020,N_11172);
or U11318 (N_11318,N_11113,N_11141);
nor U11319 (N_11319,N_11119,N_11063);
and U11320 (N_11320,N_11191,N_11089);
and U11321 (N_11321,N_11044,N_11188);
or U11322 (N_11322,N_11198,N_11238);
or U11323 (N_11323,N_11030,N_11084);
or U11324 (N_11324,N_11031,N_11219);
xnor U11325 (N_11325,N_11046,N_11123);
xnor U11326 (N_11326,N_11026,N_11126);
nand U11327 (N_11327,N_11133,N_11109);
nand U11328 (N_11328,N_11230,N_11140);
xnor U11329 (N_11329,N_11127,N_11096);
and U11330 (N_11330,N_11138,N_11006);
nor U11331 (N_11331,N_11222,N_11045);
and U11332 (N_11332,N_11194,N_11173);
and U11333 (N_11333,N_11187,N_11047);
xnor U11334 (N_11334,N_11010,N_11249);
and U11335 (N_11335,N_11024,N_11225);
nor U11336 (N_11336,N_11105,N_11120);
or U11337 (N_11337,N_11159,N_11184);
nor U11338 (N_11338,N_11168,N_11174);
or U11339 (N_11339,N_11112,N_11073);
nand U11340 (N_11340,N_11048,N_11091);
or U11341 (N_11341,N_11196,N_11102);
and U11342 (N_11342,N_11229,N_11130);
nor U11343 (N_11343,N_11122,N_11028);
xnor U11344 (N_11344,N_11206,N_11002);
and U11345 (N_11345,N_11246,N_11027);
nor U11346 (N_11346,N_11001,N_11121);
nand U11347 (N_11347,N_11178,N_11146);
nand U11348 (N_11348,N_11149,N_11104);
xnor U11349 (N_11349,N_11037,N_11070);
or U11350 (N_11350,N_11242,N_11171);
or U11351 (N_11351,N_11033,N_11211);
or U11352 (N_11352,N_11007,N_11247);
or U11353 (N_11353,N_11204,N_11065);
xor U11354 (N_11354,N_11182,N_11192);
nand U11355 (N_11355,N_11108,N_11049);
nand U11356 (N_11356,N_11199,N_11032);
nand U11357 (N_11357,N_11163,N_11009);
or U11358 (N_11358,N_11115,N_11179);
and U11359 (N_11359,N_11241,N_11132);
and U11360 (N_11360,N_11116,N_11160);
nand U11361 (N_11361,N_11228,N_11111);
or U11362 (N_11362,N_11005,N_11167);
or U11363 (N_11363,N_11040,N_11169);
xnor U11364 (N_11364,N_11036,N_11185);
nor U11365 (N_11365,N_11137,N_11147);
nor U11366 (N_11366,N_11244,N_11016);
and U11367 (N_11367,N_11124,N_11087);
or U11368 (N_11368,N_11017,N_11175);
and U11369 (N_11369,N_11075,N_11011);
xnor U11370 (N_11370,N_11021,N_11139);
nand U11371 (N_11371,N_11093,N_11114);
xnor U11372 (N_11372,N_11023,N_11125);
or U11373 (N_11373,N_11176,N_11224);
xnor U11374 (N_11374,N_11162,N_11034);
and U11375 (N_11375,N_11144,N_11186);
or U11376 (N_11376,N_11240,N_11192);
or U11377 (N_11377,N_11210,N_11157);
nand U11378 (N_11378,N_11161,N_11036);
or U11379 (N_11379,N_11155,N_11247);
or U11380 (N_11380,N_11232,N_11026);
nor U11381 (N_11381,N_11051,N_11084);
nand U11382 (N_11382,N_11240,N_11236);
or U11383 (N_11383,N_11010,N_11179);
or U11384 (N_11384,N_11159,N_11241);
nand U11385 (N_11385,N_11241,N_11235);
nor U11386 (N_11386,N_11213,N_11099);
and U11387 (N_11387,N_11228,N_11003);
or U11388 (N_11388,N_11229,N_11107);
or U11389 (N_11389,N_11044,N_11019);
or U11390 (N_11390,N_11183,N_11208);
and U11391 (N_11391,N_11087,N_11211);
or U11392 (N_11392,N_11014,N_11085);
xor U11393 (N_11393,N_11228,N_11220);
nand U11394 (N_11394,N_11100,N_11097);
and U11395 (N_11395,N_11010,N_11110);
nor U11396 (N_11396,N_11247,N_11157);
xnor U11397 (N_11397,N_11099,N_11221);
or U11398 (N_11398,N_11033,N_11093);
nand U11399 (N_11399,N_11007,N_11169);
and U11400 (N_11400,N_11029,N_11121);
xor U11401 (N_11401,N_11061,N_11140);
nand U11402 (N_11402,N_11078,N_11086);
nor U11403 (N_11403,N_11194,N_11201);
nand U11404 (N_11404,N_11144,N_11139);
nand U11405 (N_11405,N_11011,N_11121);
or U11406 (N_11406,N_11012,N_11167);
nor U11407 (N_11407,N_11120,N_11182);
or U11408 (N_11408,N_11131,N_11071);
nor U11409 (N_11409,N_11231,N_11097);
xnor U11410 (N_11410,N_11054,N_11134);
or U11411 (N_11411,N_11018,N_11042);
nor U11412 (N_11412,N_11059,N_11208);
or U11413 (N_11413,N_11081,N_11202);
nand U11414 (N_11414,N_11247,N_11112);
nand U11415 (N_11415,N_11002,N_11152);
or U11416 (N_11416,N_11106,N_11229);
nor U11417 (N_11417,N_11228,N_11094);
nor U11418 (N_11418,N_11107,N_11030);
nor U11419 (N_11419,N_11108,N_11150);
nand U11420 (N_11420,N_11124,N_11024);
or U11421 (N_11421,N_11226,N_11163);
nor U11422 (N_11422,N_11159,N_11059);
xor U11423 (N_11423,N_11235,N_11100);
and U11424 (N_11424,N_11113,N_11068);
or U11425 (N_11425,N_11065,N_11000);
or U11426 (N_11426,N_11177,N_11216);
nand U11427 (N_11427,N_11233,N_11087);
xnor U11428 (N_11428,N_11170,N_11062);
nor U11429 (N_11429,N_11004,N_11140);
nor U11430 (N_11430,N_11233,N_11081);
nor U11431 (N_11431,N_11225,N_11004);
xor U11432 (N_11432,N_11210,N_11135);
and U11433 (N_11433,N_11169,N_11249);
xnor U11434 (N_11434,N_11137,N_11014);
nand U11435 (N_11435,N_11047,N_11032);
nand U11436 (N_11436,N_11002,N_11094);
or U11437 (N_11437,N_11187,N_11151);
or U11438 (N_11438,N_11012,N_11048);
nand U11439 (N_11439,N_11217,N_11048);
nor U11440 (N_11440,N_11215,N_11145);
or U11441 (N_11441,N_11085,N_11225);
nand U11442 (N_11442,N_11067,N_11110);
xor U11443 (N_11443,N_11180,N_11188);
xnor U11444 (N_11444,N_11173,N_11003);
nand U11445 (N_11445,N_11018,N_11077);
nand U11446 (N_11446,N_11116,N_11204);
and U11447 (N_11447,N_11127,N_11080);
and U11448 (N_11448,N_11009,N_11222);
nor U11449 (N_11449,N_11244,N_11001);
nor U11450 (N_11450,N_11133,N_11199);
nor U11451 (N_11451,N_11060,N_11057);
nand U11452 (N_11452,N_11140,N_11017);
nor U11453 (N_11453,N_11044,N_11229);
nand U11454 (N_11454,N_11009,N_11122);
or U11455 (N_11455,N_11200,N_11163);
nor U11456 (N_11456,N_11234,N_11229);
nand U11457 (N_11457,N_11168,N_11189);
and U11458 (N_11458,N_11228,N_11196);
nand U11459 (N_11459,N_11239,N_11038);
or U11460 (N_11460,N_11163,N_11064);
and U11461 (N_11461,N_11215,N_11138);
nor U11462 (N_11462,N_11030,N_11059);
nand U11463 (N_11463,N_11096,N_11026);
and U11464 (N_11464,N_11076,N_11026);
and U11465 (N_11465,N_11063,N_11199);
nor U11466 (N_11466,N_11157,N_11232);
xor U11467 (N_11467,N_11159,N_11185);
nor U11468 (N_11468,N_11249,N_11211);
and U11469 (N_11469,N_11005,N_11239);
nor U11470 (N_11470,N_11249,N_11085);
nor U11471 (N_11471,N_11132,N_11200);
nand U11472 (N_11472,N_11223,N_11027);
xor U11473 (N_11473,N_11010,N_11209);
nand U11474 (N_11474,N_11007,N_11153);
nand U11475 (N_11475,N_11129,N_11034);
nand U11476 (N_11476,N_11241,N_11213);
xnor U11477 (N_11477,N_11236,N_11203);
xor U11478 (N_11478,N_11201,N_11034);
or U11479 (N_11479,N_11226,N_11030);
nand U11480 (N_11480,N_11156,N_11201);
nand U11481 (N_11481,N_11069,N_11050);
xor U11482 (N_11482,N_11209,N_11186);
and U11483 (N_11483,N_11074,N_11100);
nand U11484 (N_11484,N_11004,N_11174);
nand U11485 (N_11485,N_11061,N_11094);
or U11486 (N_11486,N_11133,N_11029);
xnor U11487 (N_11487,N_11111,N_11193);
or U11488 (N_11488,N_11082,N_11163);
xor U11489 (N_11489,N_11000,N_11214);
or U11490 (N_11490,N_11173,N_11094);
or U11491 (N_11491,N_11127,N_11083);
xnor U11492 (N_11492,N_11035,N_11013);
nand U11493 (N_11493,N_11157,N_11075);
or U11494 (N_11494,N_11078,N_11125);
nand U11495 (N_11495,N_11114,N_11029);
or U11496 (N_11496,N_11033,N_11040);
xnor U11497 (N_11497,N_11170,N_11030);
nor U11498 (N_11498,N_11052,N_11010);
xor U11499 (N_11499,N_11201,N_11172);
nand U11500 (N_11500,N_11361,N_11485);
and U11501 (N_11501,N_11300,N_11293);
or U11502 (N_11502,N_11344,N_11388);
and U11503 (N_11503,N_11301,N_11367);
nand U11504 (N_11504,N_11402,N_11492);
xor U11505 (N_11505,N_11498,N_11470);
nand U11506 (N_11506,N_11345,N_11447);
xor U11507 (N_11507,N_11466,N_11264);
nand U11508 (N_11508,N_11291,N_11386);
nor U11509 (N_11509,N_11409,N_11333);
nand U11510 (N_11510,N_11355,N_11352);
or U11511 (N_11511,N_11396,N_11284);
or U11512 (N_11512,N_11406,N_11258);
and U11513 (N_11513,N_11268,N_11390);
nor U11514 (N_11514,N_11497,N_11286);
nor U11515 (N_11515,N_11395,N_11376);
xnor U11516 (N_11516,N_11330,N_11472);
or U11517 (N_11517,N_11360,N_11343);
and U11518 (N_11518,N_11374,N_11384);
and U11519 (N_11519,N_11477,N_11275);
nand U11520 (N_11520,N_11299,N_11281);
and U11521 (N_11521,N_11433,N_11454);
or U11522 (N_11522,N_11404,N_11254);
and U11523 (N_11523,N_11487,N_11480);
and U11524 (N_11524,N_11438,N_11279);
or U11525 (N_11525,N_11282,N_11385);
nand U11526 (N_11526,N_11484,N_11399);
xnor U11527 (N_11527,N_11434,N_11290);
xor U11528 (N_11528,N_11375,N_11354);
nor U11529 (N_11529,N_11474,N_11252);
nand U11530 (N_11530,N_11411,N_11415);
nor U11531 (N_11531,N_11295,N_11313);
nand U11532 (N_11532,N_11369,N_11283);
or U11533 (N_11533,N_11348,N_11260);
and U11534 (N_11534,N_11250,N_11469);
nor U11535 (N_11535,N_11257,N_11444);
xnor U11536 (N_11536,N_11347,N_11430);
nand U11537 (N_11537,N_11315,N_11332);
nor U11538 (N_11538,N_11473,N_11277);
nor U11539 (N_11539,N_11450,N_11364);
and U11540 (N_11540,N_11280,N_11471);
xor U11541 (N_11541,N_11381,N_11346);
or U11542 (N_11542,N_11297,N_11475);
and U11543 (N_11543,N_11314,N_11368);
nor U11544 (N_11544,N_11309,N_11426);
xnor U11545 (N_11545,N_11483,N_11445);
xor U11546 (N_11546,N_11493,N_11478);
or U11547 (N_11547,N_11420,N_11261);
nand U11548 (N_11548,N_11356,N_11294);
nand U11549 (N_11549,N_11432,N_11418);
nand U11550 (N_11550,N_11302,N_11378);
and U11551 (N_11551,N_11486,N_11453);
or U11552 (N_11552,N_11408,N_11351);
nand U11553 (N_11553,N_11391,N_11458);
nor U11554 (N_11554,N_11319,N_11272);
nand U11555 (N_11555,N_11461,N_11392);
nor U11556 (N_11556,N_11412,N_11379);
nor U11557 (N_11557,N_11489,N_11455);
nor U11558 (N_11558,N_11358,N_11339);
and U11559 (N_11559,N_11320,N_11436);
nand U11560 (N_11560,N_11407,N_11256);
nand U11561 (N_11561,N_11394,N_11441);
xnor U11562 (N_11562,N_11413,N_11273);
or U11563 (N_11563,N_11429,N_11366);
xnor U11564 (N_11564,N_11446,N_11298);
or U11565 (N_11565,N_11499,N_11398);
or U11566 (N_11566,N_11292,N_11372);
or U11567 (N_11567,N_11449,N_11359);
nand U11568 (N_11568,N_11382,N_11251);
nand U11569 (N_11569,N_11288,N_11479);
or U11570 (N_11570,N_11371,N_11327);
xnor U11571 (N_11571,N_11405,N_11465);
nand U11572 (N_11572,N_11324,N_11263);
nor U11573 (N_11573,N_11340,N_11306);
or U11574 (N_11574,N_11276,N_11427);
or U11575 (N_11575,N_11308,N_11439);
xor U11576 (N_11576,N_11421,N_11459);
or U11577 (N_11577,N_11370,N_11400);
or U11578 (N_11578,N_11323,N_11296);
or U11579 (N_11579,N_11329,N_11467);
xnor U11580 (N_11580,N_11266,N_11490);
nor U11581 (N_11581,N_11424,N_11322);
and U11582 (N_11582,N_11435,N_11336);
nor U11583 (N_11583,N_11317,N_11262);
nor U11584 (N_11584,N_11259,N_11387);
or U11585 (N_11585,N_11287,N_11349);
nand U11586 (N_11586,N_11274,N_11389);
or U11587 (N_11587,N_11419,N_11488);
nand U11588 (N_11588,N_11285,N_11383);
nand U11589 (N_11589,N_11422,N_11464);
and U11590 (N_11590,N_11321,N_11425);
or U11591 (N_11591,N_11442,N_11414);
or U11592 (N_11592,N_11440,N_11328);
and U11593 (N_11593,N_11494,N_11393);
nand U11594 (N_11594,N_11342,N_11311);
nand U11595 (N_11595,N_11403,N_11307);
nor U11596 (N_11596,N_11316,N_11495);
nand U11597 (N_11597,N_11431,N_11416);
xor U11598 (N_11598,N_11410,N_11463);
nor U11599 (N_11599,N_11357,N_11303);
nor U11600 (N_11600,N_11423,N_11460);
nor U11601 (N_11601,N_11341,N_11468);
or U11602 (N_11602,N_11448,N_11271);
nor U11603 (N_11603,N_11428,N_11325);
nor U11604 (N_11604,N_11310,N_11482);
xor U11605 (N_11605,N_11462,N_11278);
nand U11606 (N_11606,N_11270,N_11255);
nand U11607 (N_11607,N_11443,N_11269);
or U11608 (N_11608,N_11451,N_11362);
nand U11609 (N_11609,N_11365,N_11318);
xor U11610 (N_11610,N_11312,N_11481);
and U11611 (N_11611,N_11304,N_11326);
nand U11612 (N_11612,N_11335,N_11380);
and U11613 (N_11613,N_11373,N_11491);
and U11614 (N_11614,N_11457,N_11417);
nor U11615 (N_11615,N_11476,N_11377);
or U11616 (N_11616,N_11253,N_11496);
or U11617 (N_11617,N_11331,N_11452);
xor U11618 (N_11618,N_11456,N_11337);
or U11619 (N_11619,N_11397,N_11363);
nor U11620 (N_11620,N_11267,N_11401);
nand U11621 (N_11621,N_11437,N_11353);
or U11622 (N_11622,N_11265,N_11338);
nor U11623 (N_11623,N_11305,N_11334);
and U11624 (N_11624,N_11350,N_11289);
nand U11625 (N_11625,N_11308,N_11421);
xnor U11626 (N_11626,N_11326,N_11275);
and U11627 (N_11627,N_11325,N_11379);
nand U11628 (N_11628,N_11360,N_11351);
nand U11629 (N_11629,N_11286,N_11255);
nor U11630 (N_11630,N_11355,N_11306);
nor U11631 (N_11631,N_11382,N_11448);
nor U11632 (N_11632,N_11318,N_11378);
and U11633 (N_11633,N_11436,N_11426);
nand U11634 (N_11634,N_11445,N_11313);
and U11635 (N_11635,N_11408,N_11301);
and U11636 (N_11636,N_11393,N_11345);
nand U11637 (N_11637,N_11386,N_11363);
or U11638 (N_11638,N_11396,N_11417);
nor U11639 (N_11639,N_11322,N_11358);
and U11640 (N_11640,N_11390,N_11309);
nor U11641 (N_11641,N_11351,N_11275);
nor U11642 (N_11642,N_11330,N_11284);
xnor U11643 (N_11643,N_11340,N_11294);
nand U11644 (N_11644,N_11278,N_11429);
xor U11645 (N_11645,N_11387,N_11260);
and U11646 (N_11646,N_11460,N_11389);
nor U11647 (N_11647,N_11455,N_11267);
or U11648 (N_11648,N_11273,N_11458);
and U11649 (N_11649,N_11326,N_11378);
or U11650 (N_11650,N_11322,N_11324);
xor U11651 (N_11651,N_11406,N_11461);
and U11652 (N_11652,N_11339,N_11447);
nor U11653 (N_11653,N_11464,N_11345);
or U11654 (N_11654,N_11496,N_11341);
or U11655 (N_11655,N_11471,N_11252);
and U11656 (N_11656,N_11258,N_11313);
or U11657 (N_11657,N_11331,N_11370);
nand U11658 (N_11658,N_11471,N_11494);
nor U11659 (N_11659,N_11351,N_11310);
nand U11660 (N_11660,N_11454,N_11367);
or U11661 (N_11661,N_11290,N_11428);
nand U11662 (N_11662,N_11284,N_11266);
and U11663 (N_11663,N_11480,N_11255);
nor U11664 (N_11664,N_11493,N_11468);
xnor U11665 (N_11665,N_11410,N_11337);
and U11666 (N_11666,N_11367,N_11418);
nor U11667 (N_11667,N_11436,N_11455);
xor U11668 (N_11668,N_11361,N_11315);
nor U11669 (N_11669,N_11368,N_11410);
nor U11670 (N_11670,N_11346,N_11361);
nor U11671 (N_11671,N_11440,N_11489);
and U11672 (N_11672,N_11336,N_11408);
xor U11673 (N_11673,N_11380,N_11321);
or U11674 (N_11674,N_11357,N_11452);
and U11675 (N_11675,N_11449,N_11344);
xnor U11676 (N_11676,N_11485,N_11450);
or U11677 (N_11677,N_11473,N_11379);
nor U11678 (N_11678,N_11389,N_11300);
nand U11679 (N_11679,N_11264,N_11381);
xnor U11680 (N_11680,N_11379,N_11418);
and U11681 (N_11681,N_11357,N_11415);
nand U11682 (N_11682,N_11277,N_11286);
and U11683 (N_11683,N_11369,N_11316);
nor U11684 (N_11684,N_11362,N_11406);
nor U11685 (N_11685,N_11281,N_11318);
nand U11686 (N_11686,N_11499,N_11266);
and U11687 (N_11687,N_11312,N_11465);
xnor U11688 (N_11688,N_11259,N_11349);
nand U11689 (N_11689,N_11487,N_11374);
xnor U11690 (N_11690,N_11485,N_11381);
or U11691 (N_11691,N_11346,N_11387);
xor U11692 (N_11692,N_11470,N_11345);
and U11693 (N_11693,N_11370,N_11459);
nor U11694 (N_11694,N_11461,N_11437);
or U11695 (N_11695,N_11346,N_11420);
and U11696 (N_11696,N_11461,N_11370);
nand U11697 (N_11697,N_11499,N_11472);
and U11698 (N_11698,N_11381,N_11430);
or U11699 (N_11699,N_11263,N_11487);
xor U11700 (N_11700,N_11305,N_11417);
xor U11701 (N_11701,N_11428,N_11472);
and U11702 (N_11702,N_11261,N_11351);
nor U11703 (N_11703,N_11352,N_11309);
xnor U11704 (N_11704,N_11326,N_11398);
xor U11705 (N_11705,N_11267,N_11422);
nor U11706 (N_11706,N_11415,N_11268);
xor U11707 (N_11707,N_11370,N_11349);
and U11708 (N_11708,N_11483,N_11324);
xor U11709 (N_11709,N_11362,N_11470);
xor U11710 (N_11710,N_11458,N_11429);
or U11711 (N_11711,N_11297,N_11386);
nand U11712 (N_11712,N_11464,N_11300);
xor U11713 (N_11713,N_11329,N_11385);
nand U11714 (N_11714,N_11376,N_11258);
and U11715 (N_11715,N_11437,N_11422);
nor U11716 (N_11716,N_11391,N_11258);
nand U11717 (N_11717,N_11439,N_11306);
and U11718 (N_11718,N_11277,N_11378);
or U11719 (N_11719,N_11342,N_11445);
or U11720 (N_11720,N_11446,N_11363);
or U11721 (N_11721,N_11406,N_11255);
xnor U11722 (N_11722,N_11327,N_11267);
or U11723 (N_11723,N_11341,N_11401);
nand U11724 (N_11724,N_11341,N_11282);
nand U11725 (N_11725,N_11343,N_11479);
xnor U11726 (N_11726,N_11436,N_11310);
nand U11727 (N_11727,N_11337,N_11378);
nor U11728 (N_11728,N_11268,N_11407);
and U11729 (N_11729,N_11409,N_11352);
nor U11730 (N_11730,N_11349,N_11467);
nor U11731 (N_11731,N_11487,N_11258);
nand U11732 (N_11732,N_11407,N_11399);
xor U11733 (N_11733,N_11465,N_11400);
nand U11734 (N_11734,N_11322,N_11441);
xor U11735 (N_11735,N_11431,N_11407);
and U11736 (N_11736,N_11334,N_11364);
or U11737 (N_11737,N_11258,N_11430);
and U11738 (N_11738,N_11452,N_11354);
nor U11739 (N_11739,N_11332,N_11300);
or U11740 (N_11740,N_11343,N_11469);
or U11741 (N_11741,N_11294,N_11308);
xnor U11742 (N_11742,N_11351,N_11478);
nand U11743 (N_11743,N_11456,N_11273);
and U11744 (N_11744,N_11347,N_11326);
or U11745 (N_11745,N_11434,N_11385);
xnor U11746 (N_11746,N_11281,N_11274);
xor U11747 (N_11747,N_11488,N_11473);
nand U11748 (N_11748,N_11414,N_11367);
and U11749 (N_11749,N_11407,N_11285);
nor U11750 (N_11750,N_11692,N_11567);
nor U11751 (N_11751,N_11666,N_11621);
xnor U11752 (N_11752,N_11594,N_11586);
nand U11753 (N_11753,N_11605,N_11546);
and U11754 (N_11754,N_11609,N_11566);
nand U11755 (N_11755,N_11743,N_11510);
or U11756 (N_11756,N_11708,N_11695);
xnor U11757 (N_11757,N_11629,N_11678);
and U11758 (N_11758,N_11651,N_11710);
nand U11759 (N_11759,N_11725,N_11749);
nor U11760 (N_11760,N_11630,N_11559);
nor U11761 (N_11761,N_11745,N_11735);
and U11762 (N_11762,N_11671,N_11657);
nand U11763 (N_11763,N_11705,N_11730);
and U11764 (N_11764,N_11508,N_11739);
or U11765 (N_11765,N_11719,N_11602);
nor U11766 (N_11766,N_11561,N_11728);
and U11767 (N_11767,N_11744,N_11616);
xor U11768 (N_11768,N_11627,N_11556);
nand U11769 (N_11769,N_11670,N_11713);
nor U11770 (N_11770,N_11506,N_11531);
and U11771 (N_11771,N_11694,N_11523);
nor U11772 (N_11772,N_11702,N_11626);
and U11773 (N_11773,N_11722,N_11598);
and U11774 (N_11774,N_11664,N_11652);
xor U11775 (N_11775,N_11577,N_11623);
nand U11776 (N_11776,N_11599,N_11521);
nand U11777 (N_11777,N_11524,N_11672);
and U11778 (N_11778,N_11717,N_11679);
nor U11779 (N_11779,N_11654,N_11747);
xor U11780 (N_11780,N_11693,N_11742);
nor U11781 (N_11781,N_11607,N_11554);
xor U11782 (N_11782,N_11593,N_11587);
and U11783 (N_11783,N_11550,N_11689);
nor U11784 (N_11784,N_11700,N_11653);
nor U11785 (N_11785,N_11522,N_11535);
nand U11786 (N_11786,N_11649,N_11603);
xnor U11787 (N_11787,N_11646,N_11727);
nor U11788 (N_11788,N_11720,N_11676);
nor U11789 (N_11789,N_11677,N_11538);
or U11790 (N_11790,N_11513,N_11613);
and U11791 (N_11791,N_11548,N_11637);
nor U11792 (N_11792,N_11628,N_11686);
nor U11793 (N_11793,N_11588,N_11663);
nor U11794 (N_11794,N_11501,N_11589);
xnor U11795 (N_11795,N_11715,N_11711);
xor U11796 (N_11796,N_11631,N_11734);
or U11797 (N_11797,N_11574,N_11737);
nand U11798 (N_11798,N_11504,N_11580);
or U11799 (N_11799,N_11511,N_11576);
nand U11800 (N_11800,N_11684,N_11596);
or U11801 (N_11801,N_11517,N_11712);
or U11802 (N_11802,N_11509,N_11592);
or U11803 (N_11803,N_11633,N_11557);
or U11804 (N_11804,N_11721,N_11617);
xor U11805 (N_11805,N_11542,N_11748);
or U11806 (N_11806,N_11558,N_11595);
or U11807 (N_11807,N_11645,N_11632);
nor U11808 (N_11808,N_11563,N_11578);
and U11809 (N_11809,N_11555,N_11514);
and U11810 (N_11810,N_11610,N_11544);
nand U11811 (N_11811,N_11614,N_11724);
or U11812 (N_11812,N_11619,N_11667);
nor U11813 (N_11813,N_11519,N_11526);
and U11814 (N_11814,N_11530,N_11726);
xnor U11815 (N_11815,N_11641,N_11635);
xor U11816 (N_11816,N_11697,N_11634);
nor U11817 (N_11817,N_11618,N_11565);
and U11818 (N_11818,N_11655,N_11718);
nor U11819 (N_11819,N_11573,N_11738);
and U11820 (N_11820,N_11674,N_11650);
xnor U11821 (N_11821,N_11648,N_11690);
or U11822 (N_11822,N_11536,N_11662);
nand U11823 (N_11823,N_11591,N_11661);
or U11824 (N_11824,N_11703,N_11699);
nor U11825 (N_11825,N_11516,N_11740);
nor U11826 (N_11826,N_11644,N_11741);
xor U11827 (N_11827,N_11680,N_11560);
xor U11828 (N_11828,N_11601,N_11590);
nand U11829 (N_11829,N_11553,N_11547);
nor U11830 (N_11830,N_11543,N_11528);
xnor U11831 (N_11831,N_11608,N_11551);
and U11832 (N_11832,N_11515,N_11681);
and U11833 (N_11833,N_11668,N_11583);
or U11834 (N_11834,N_11723,N_11529);
xnor U11835 (N_11835,N_11691,N_11537);
and U11836 (N_11836,N_11642,N_11636);
nand U11837 (N_11837,N_11525,N_11600);
or U11838 (N_11838,N_11503,N_11647);
nand U11839 (N_11839,N_11582,N_11604);
and U11840 (N_11840,N_11643,N_11687);
nor U11841 (N_11841,N_11584,N_11597);
and U11842 (N_11842,N_11541,N_11532);
nor U11843 (N_11843,N_11545,N_11660);
nor U11844 (N_11844,N_11736,N_11624);
or U11845 (N_11845,N_11549,N_11714);
or U11846 (N_11846,N_11729,N_11696);
xor U11847 (N_11847,N_11716,N_11518);
and U11848 (N_11848,N_11611,N_11659);
or U11849 (N_11849,N_11606,N_11673);
or U11850 (N_11850,N_11658,N_11709);
nor U11851 (N_11851,N_11733,N_11688);
nor U11852 (N_11852,N_11746,N_11575);
nand U11853 (N_11853,N_11656,N_11675);
or U11854 (N_11854,N_11732,N_11639);
xor U11855 (N_11855,N_11620,N_11571);
nand U11856 (N_11856,N_11568,N_11638);
nor U11857 (N_11857,N_11507,N_11622);
nor U11858 (N_11858,N_11540,N_11625);
xnor U11859 (N_11859,N_11682,N_11698);
or U11860 (N_11860,N_11615,N_11539);
nor U11861 (N_11861,N_11731,N_11533);
nand U11862 (N_11862,N_11669,N_11612);
nand U11863 (N_11863,N_11640,N_11552);
or U11864 (N_11864,N_11502,N_11581);
or U11865 (N_11865,N_11512,N_11706);
nand U11866 (N_11866,N_11704,N_11570);
or U11867 (N_11867,N_11500,N_11520);
and U11868 (N_11868,N_11585,N_11564);
and U11869 (N_11869,N_11685,N_11579);
and U11870 (N_11870,N_11527,N_11707);
and U11871 (N_11871,N_11505,N_11683);
nor U11872 (N_11872,N_11572,N_11569);
nand U11873 (N_11873,N_11562,N_11665);
or U11874 (N_11874,N_11534,N_11701);
nand U11875 (N_11875,N_11697,N_11749);
xnor U11876 (N_11876,N_11610,N_11614);
xnor U11877 (N_11877,N_11687,N_11586);
nand U11878 (N_11878,N_11634,N_11572);
nand U11879 (N_11879,N_11683,N_11580);
or U11880 (N_11880,N_11682,N_11685);
xnor U11881 (N_11881,N_11572,N_11573);
or U11882 (N_11882,N_11698,N_11522);
nor U11883 (N_11883,N_11530,N_11687);
xnor U11884 (N_11884,N_11725,N_11584);
nor U11885 (N_11885,N_11703,N_11663);
or U11886 (N_11886,N_11601,N_11617);
and U11887 (N_11887,N_11573,N_11600);
and U11888 (N_11888,N_11717,N_11513);
nand U11889 (N_11889,N_11667,N_11695);
xor U11890 (N_11890,N_11535,N_11528);
nor U11891 (N_11891,N_11668,N_11536);
nand U11892 (N_11892,N_11563,N_11702);
nand U11893 (N_11893,N_11536,N_11747);
or U11894 (N_11894,N_11627,N_11639);
xor U11895 (N_11895,N_11579,N_11614);
nor U11896 (N_11896,N_11551,N_11515);
nor U11897 (N_11897,N_11595,N_11701);
and U11898 (N_11898,N_11720,N_11513);
nor U11899 (N_11899,N_11603,N_11670);
nand U11900 (N_11900,N_11660,N_11617);
nand U11901 (N_11901,N_11638,N_11631);
nor U11902 (N_11902,N_11592,N_11536);
or U11903 (N_11903,N_11717,N_11702);
or U11904 (N_11904,N_11621,N_11566);
xor U11905 (N_11905,N_11650,N_11566);
nand U11906 (N_11906,N_11728,N_11595);
and U11907 (N_11907,N_11651,N_11515);
xnor U11908 (N_11908,N_11631,N_11702);
nand U11909 (N_11909,N_11688,N_11702);
or U11910 (N_11910,N_11533,N_11749);
nor U11911 (N_11911,N_11565,N_11702);
nand U11912 (N_11912,N_11697,N_11536);
nor U11913 (N_11913,N_11606,N_11538);
nor U11914 (N_11914,N_11661,N_11659);
xnor U11915 (N_11915,N_11585,N_11713);
or U11916 (N_11916,N_11617,N_11589);
xnor U11917 (N_11917,N_11552,N_11520);
nand U11918 (N_11918,N_11691,N_11713);
or U11919 (N_11919,N_11595,N_11715);
xnor U11920 (N_11920,N_11666,N_11502);
xor U11921 (N_11921,N_11563,N_11622);
and U11922 (N_11922,N_11521,N_11597);
nand U11923 (N_11923,N_11689,N_11720);
and U11924 (N_11924,N_11500,N_11672);
and U11925 (N_11925,N_11506,N_11690);
nand U11926 (N_11926,N_11585,N_11621);
nor U11927 (N_11927,N_11720,N_11705);
or U11928 (N_11928,N_11626,N_11680);
and U11929 (N_11929,N_11684,N_11637);
nor U11930 (N_11930,N_11738,N_11663);
nor U11931 (N_11931,N_11503,N_11729);
nand U11932 (N_11932,N_11631,N_11622);
nor U11933 (N_11933,N_11565,N_11711);
or U11934 (N_11934,N_11567,N_11599);
xnor U11935 (N_11935,N_11567,N_11654);
or U11936 (N_11936,N_11730,N_11535);
xnor U11937 (N_11937,N_11600,N_11587);
and U11938 (N_11938,N_11638,N_11502);
and U11939 (N_11939,N_11555,N_11717);
nand U11940 (N_11940,N_11503,N_11562);
and U11941 (N_11941,N_11619,N_11624);
xor U11942 (N_11942,N_11593,N_11553);
xor U11943 (N_11943,N_11555,N_11515);
nor U11944 (N_11944,N_11569,N_11501);
or U11945 (N_11945,N_11745,N_11592);
nand U11946 (N_11946,N_11551,N_11543);
xor U11947 (N_11947,N_11696,N_11739);
or U11948 (N_11948,N_11739,N_11567);
nand U11949 (N_11949,N_11633,N_11530);
nor U11950 (N_11950,N_11705,N_11570);
nor U11951 (N_11951,N_11660,N_11747);
nand U11952 (N_11952,N_11732,N_11508);
and U11953 (N_11953,N_11662,N_11698);
or U11954 (N_11954,N_11674,N_11598);
xor U11955 (N_11955,N_11712,N_11520);
and U11956 (N_11956,N_11574,N_11733);
xnor U11957 (N_11957,N_11656,N_11728);
or U11958 (N_11958,N_11540,N_11612);
and U11959 (N_11959,N_11590,N_11661);
xnor U11960 (N_11960,N_11672,N_11749);
nand U11961 (N_11961,N_11584,N_11723);
nor U11962 (N_11962,N_11535,N_11628);
and U11963 (N_11963,N_11739,N_11510);
nand U11964 (N_11964,N_11672,N_11628);
xor U11965 (N_11965,N_11529,N_11631);
or U11966 (N_11966,N_11620,N_11521);
and U11967 (N_11967,N_11691,N_11543);
nor U11968 (N_11968,N_11613,N_11608);
nand U11969 (N_11969,N_11603,N_11697);
or U11970 (N_11970,N_11666,N_11501);
and U11971 (N_11971,N_11530,N_11585);
or U11972 (N_11972,N_11729,N_11571);
nor U11973 (N_11973,N_11736,N_11538);
xnor U11974 (N_11974,N_11515,N_11719);
and U11975 (N_11975,N_11524,N_11729);
or U11976 (N_11976,N_11661,N_11716);
nand U11977 (N_11977,N_11510,N_11711);
and U11978 (N_11978,N_11579,N_11629);
xor U11979 (N_11979,N_11562,N_11698);
nand U11980 (N_11980,N_11588,N_11545);
or U11981 (N_11981,N_11644,N_11592);
and U11982 (N_11982,N_11644,N_11589);
and U11983 (N_11983,N_11636,N_11683);
and U11984 (N_11984,N_11598,N_11745);
nor U11985 (N_11985,N_11597,N_11662);
nand U11986 (N_11986,N_11580,N_11663);
nand U11987 (N_11987,N_11548,N_11604);
or U11988 (N_11988,N_11707,N_11521);
nand U11989 (N_11989,N_11680,N_11712);
nand U11990 (N_11990,N_11599,N_11500);
xor U11991 (N_11991,N_11517,N_11749);
nor U11992 (N_11992,N_11748,N_11523);
or U11993 (N_11993,N_11711,N_11516);
xor U11994 (N_11994,N_11556,N_11619);
nand U11995 (N_11995,N_11629,N_11520);
nor U11996 (N_11996,N_11623,N_11640);
xor U11997 (N_11997,N_11706,N_11658);
or U11998 (N_11998,N_11725,N_11730);
nand U11999 (N_11999,N_11636,N_11627);
and U12000 (N_12000,N_11762,N_11940);
xor U12001 (N_12001,N_11981,N_11784);
nor U12002 (N_12002,N_11836,N_11787);
and U12003 (N_12003,N_11831,N_11898);
nor U12004 (N_12004,N_11982,N_11942);
nand U12005 (N_12005,N_11855,N_11755);
xor U12006 (N_12006,N_11969,N_11935);
nor U12007 (N_12007,N_11845,N_11890);
xnor U12008 (N_12008,N_11919,N_11824);
nor U12009 (N_12009,N_11875,N_11767);
and U12010 (N_12010,N_11992,N_11843);
nor U12011 (N_12011,N_11946,N_11889);
nor U12012 (N_12012,N_11886,N_11977);
nand U12013 (N_12013,N_11901,N_11926);
and U12014 (N_12014,N_11760,N_11863);
or U12015 (N_12015,N_11816,N_11996);
and U12016 (N_12016,N_11869,N_11954);
nor U12017 (N_12017,N_11949,N_11939);
nand U12018 (N_12018,N_11874,N_11789);
or U12019 (N_12019,N_11828,N_11833);
nand U12020 (N_12020,N_11983,N_11840);
nor U12021 (N_12021,N_11763,N_11930);
and U12022 (N_12022,N_11997,N_11795);
nor U12023 (N_12023,N_11776,N_11881);
nor U12024 (N_12024,N_11822,N_11777);
and U12025 (N_12025,N_11959,N_11927);
nand U12026 (N_12026,N_11974,N_11979);
or U12027 (N_12027,N_11908,N_11800);
xnor U12028 (N_12028,N_11827,N_11844);
xor U12029 (N_12029,N_11904,N_11923);
nor U12030 (N_12030,N_11765,N_11913);
or U12031 (N_12031,N_11798,N_11905);
and U12032 (N_12032,N_11814,N_11922);
nor U12033 (N_12033,N_11835,N_11810);
nor U12034 (N_12034,N_11903,N_11912);
nand U12035 (N_12035,N_11998,N_11803);
nand U12036 (N_12036,N_11860,N_11887);
or U12037 (N_12037,N_11915,N_11857);
nor U12038 (N_12038,N_11968,N_11955);
or U12039 (N_12039,N_11924,N_11988);
nand U12040 (N_12040,N_11995,N_11773);
nor U12041 (N_12041,N_11895,N_11779);
and U12042 (N_12042,N_11770,N_11782);
nand U12043 (N_12043,N_11952,N_11821);
xnor U12044 (N_12044,N_11984,N_11756);
nor U12045 (N_12045,N_11794,N_11853);
xnor U12046 (N_12046,N_11964,N_11873);
and U12047 (N_12047,N_11967,N_11790);
and U12048 (N_12048,N_11956,N_11953);
nor U12049 (N_12049,N_11879,N_11958);
nand U12050 (N_12050,N_11994,N_11754);
nor U12051 (N_12051,N_11902,N_11916);
xor U12052 (N_12052,N_11829,N_11896);
or U12053 (N_12053,N_11973,N_11808);
and U12054 (N_12054,N_11793,N_11847);
or U12055 (N_12055,N_11980,N_11972);
nand U12056 (N_12056,N_11870,N_11978);
and U12057 (N_12057,N_11757,N_11850);
or U12058 (N_12058,N_11768,N_11832);
nand U12059 (N_12059,N_11987,N_11830);
or U12060 (N_12060,N_11888,N_11841);
nor U12061 (N_12061,N_11778,N_11826);
nand U12062 (N_12062,N_11951,N_11788);
or U12063 (N_12063,N_11825,N_11945);
and U12064 (N_12064,N_11797,N_11911);
xor U12065 (N_12065,N_11976,N_11993);
nand U12066 (N_12066,N_11815,N_11918);
or U12067 (N_12067,N_11837,N_11943);
or U12068 (N_12068,N_11851,N_11868);
or U12069 (N_12069,N_11820,N_11750);
xor U12070 (N_12070,N_11891,N_11909);
xor U12071 (N_12071,N_11842,N_11906);
or U12072 (N_12072,N_11971,N_11878);
nor U12073 (N_12073,N_11948,N_11846);
xor U12074 (N_12074,N_11859,N_11771);
xnor U12075 (N_12075,N_11884,N_11766);
nand U12076 (N_12076,N_11986,N_11928);
and U12077 (N_12077,N_11933,N_11932);
or U12078 (N_12078,N_11806,N_11883);
nor U12079 (N_12079,N_11801,N_11944);
nand U12080 (N_12080,N_11819,N_11848);
nand U12081 (N_12081,N_11807,N_11805);
and U12082 (N_12082,N_11769,N_11900);
or U12083 (N_12083,N_11813,N_11882);
nand U12084 (N_12084,N_11936,N_11792);
nor U12085 (N_12085,N_11852,N_11907);
nand U12086 (N_12086,N_11961,N_11950);
xnor U12087 (N_12087,N_11897,N_11931);
or U12088 (N_12088,N_11812,N_11921);
and U12089 (N_12089,N_11938,N_11785);
and U12090 (N_12090,N_11751,N_11876);
or U12091 (N_12091,N_11910,N_11934);
nor U12092 (N_12092,N_11802,N_11772);
and U12093 (N_12093,N_11780,N_11817);
xor U12094 (N_12094,N_11929,N_11991);
xnor U12095 (N_12095,N_11796,N_11925);
xnor U12096 (N_12096,N_11894,N_11917);
or U12097 (N_12097,N_11963,N_11866);
xnor U12098 (N_12098,N_11809,N_11960);
xnor U12099 (N_12099,N_11914,N_11849);
nor U12100 (N_12100,N_11871,N_11864);
nor U12101 (N_12101,N_11858,N_11761);
nor U12102 (N_12102,N_11893,N_11786);
xnor U12103 (N_12103,N_11867,N_11872);
nor U12104 (N_12104,N_11783,N_11965);
xnor U12105 (N_12105,N_11989,N_11970);
xor U12106 (N_12106,N_11975,N_11764);
nand U12107 (N_12107,N_11999,N_11811);
nand U12108 (N_12108,N_11861,N_11839);
nand U12109 (N_12109,N_11804,N_11966);
and U12110 (N_12110,N_11892,N_11775);
nor U12111 (N_12111,N_11985,N_11799);
nand U12112 (N_12112,N_11838,N_11752);
or U12113 (N_12113,N_11818,N_11823);
or U12114 (N_12114,N_11990,N_11774);
nand U12115 (N_12115,N_11957,N_11856);
nand U12116 (N_12116,N_11854,N_11947);
xnor U12117 (N_12117,N_11791,N_11753);
or U12118 (N_12118,N_11862,N_11920);
nand U12119 (N_12119,N_11937,N_11834);
nand U12120 (N_12120,N_11885,N_11962);
and U12121 (N_12121,N_11899,N_11941);
and U12122 (N_12122,N_11781,N_11880);
nor U12123 (N_12123,N_11865,N_11877);
or U12124 (N_12124,N_11759,N_11758);
or U12125 (N_12125,N_11937,N_11920);
nand U12126 (N_12126,N_11869,N_11850);
nand U12127 (N_12127,N_11788,N_11994);
xor U12128 (N_12128,N_11804,N_11845);
nor U12129 (N_12129,N_11904,N_11793);
or U12130 (N_12130,N_11918,N_11757);
or U12131 (N_12131,N_11934,N_11965);
nand U12132 (N_12132,N_11806,N_11930);
xnor U12133 (N_12133,N_11861,N_11968);
nor U12134 (N_12134,N_11898,N_11861);
and U12135 (N_12135,N_11827,N_11783);
or U12136 (N_12136,N_11786,N_11854);
or U12137 (N_12137,N_11815,N_11919);
and U12138 (N_12138,N_11970,N_11964);
and U12139 (N_12139,N_11837,N_11968);
nand U12140 (N_12140,N_11822,N_11844);
and U12141 (N_12141,N_11773,N_11978);
xor U12142 (N_12142,N_11948,N_11854);
nand U12143 (N_12143,N_11948,N_11994);
or U12144 (N_12144,N_11967,N_11856);
and U12145 (N_12145,N_11962,N_11859);
nand U12146 (N_12146,N_11940,N_11804);
nand U12147 (N_12147,N_11996,N_11812);
or U12148 (N_12148,N_11927,N_11836);
nand U12149 (N_12149,N_11880,N_11914);
and U12150 (N_12150,N_11931,N_11909);
or U12151 (N_12151,N_11962,N_11765);
nand U12152 (N_12152,N_11954,N_11787);
nand U12153 (N_12153,N_11957,N_11927);
and U12154 (N_12154,N_11942,N_11956);
or U12155 (N_12155,N_11936,N_11818);
xor U12156 (N_12156,N_11876,N_11925);
or U12157 (N_12157,N_11853,N_11772);
nand U12158 (N_12158,N_11791,N_11815);
xnor U12159 (N_12159,N_11769,N_11983);
and U12160 (N_12160,N_11881,N_11920);
and U12161 (N_12161,N_11994,N_11964);
nand U12162 (N_12162,N_11930,N_11802);
nand U12163 (N_12163,N_11952,N_11879);
or U12164 (N_12164,N_11785,N_11830);
nand U12165 (N_12165,N_11831,N_11998);
nand U12166 (N_12166,N_11764,N_11921);
nand U12167 (N_12167,N_11868,N_11878);
xnor U12168 (N_12168,N_11942,N_11885);
xor U12169 (N_12169,N_11852,N_11768);
nand U12170 (N_12170,N_11995,N_11785);
nor U12171 (N_12171,N_11809,N_11860);
nand U12172 (N_12172,N_11763,N_11972);
and U12173 (N_12173,N_11924,N_11971);
or U12174 (N_12174,N_11906,N_11975);
or U12175 (N_12175,N_11919,N_11879);
nor U12176 (N_12176,N_11807,N_11990);
xnor U12177 (N_12177,N_11886,N_11873);
and U12178 (N_12178,N_11813,N_11878);
and U12179 (N_12179,N_11787,N_11969);
nor U12180 (N_12180,N_11996,N_11820);
and U12181 (N_12181,N_11948,N_11818);
nand U12182 (N_12182,N_11873,N_11785);
and U12183 (N_12183,N_11952,N_11766);
nand U12184 (N_12184,N_11845,N_11919);
xor U12185 (N_12185,N_11897,N_11987);
and U12186 (N_12186,N_11939,N_11760);
nor U12187 (N_12187,N_11965,N_11998);
and U12188 (N_12188,N_11943,N_11924);
xnor U12189 (N_12189,N_11841,N_11909);
nor U12190 (N_12190,N_11983,N_11978);
and U12191 (N_12191,N_11768,N_11972);
nand U12192 (N_12192,N_11825,N_11799);
and U12193 (N_12193,N_11778,N_11989);
nand U12194 (N_12194,N_11890,N_11996);
nor U12195 (N_12195,N_11991,N_11947);
and U12196 (N_12196,N_11896,N_11971);
xor U12197 (N_12197,N_11806,N_11852);
nand U12198 (N_12198,N_11904,N_11984);
nand U12199 (N_12199,N_11859,N_11849);
xor U12200 (N_12200,N_11837,N_11982);
and U12201 (N_12201,N_11809,N_11799);
nor U12202 (N_12202,N_11956,N_11901);
nand U12203 (N_12203,N_11920,N_11812);
nand U12204 (N_12204,N_11994,N_11912);
and U12205 (N_12205,N_11802,N_11968);
xnor U12206 (N_12206,N_11815,N_11979);
nor U12207 (N_12207,N_11815,N_11942);
or U12208 (N_12208,N_11757,N_11982);
xor U12209 (N_12209,N_11807,N_11901);
and U12210 (N_12210,N_11797,N_11803);
nor U12211 (N_12211,N_11928,N_11848);
and U12212 (N_12212,N_11778,N_11855);
nand U12213 (N_12213,N_11854,N_11894);
nand U12214 (N_12214,N_11800,N_11975);
xor U12215 (N_12215,N_11875,N_11832);
and U12216 (N_12216,N_11896,N_11992);
xnor U12217 (N_12217,N_11815,N_11884);
or U12218 (N_12218,N_11982,N_11909);
nor U12219 (N_12219,N_11774,N_11840);
nand U12220 (N_12220,N_11836,N_11876);
and U12221 (N_12221,N_11877,N_11786);
or U12222 (N_12222,N_11886,N_11769);
nor U12223 (N_12223,N_11919,N_11872);
nand U12224 (N_12224,N_11762,N_11825);
nor U12225 (N_12225,N_11852,N_11786);
and U12226 (N_12226,N_11948,N_11856);
nor U12227 (N_12227,N_11928,N_11850);
or U12228 (N_12228,N_11903,N_11780);
nand U12229 (N_12229,N_11941,N_11921);
nand U12230 (N_12230,N_11883,N_11807);
and U12231 (N_12231,N_11918,N_11996);
and U12232 (N_12232,N_11926,N_11864);
nand U12233 (N_12233,N_11830,N_11954);
and U12234 (N_12234,N_11984,N_11936);
xnor U12235 (N_12235,N_11913,N_11890);
nand U12236 (N_12236,N_11913,N_11861);
or U12237 (N_12237,N_11771,N_11861);
xnor U12238 (N_12238,N_11788,N_11798);
or U12239 (N_12239,N_11757,N_11813);
nor U12240 (N_12240,N_11898,N_11977);
nand U12241 (N_12241,N_11893,N_11824);
nor U12242 (N_12242,N_11984,N_11970);
nand U12243 (N_12243,N_11891,N_11887);
nand U12244 (N_12244,N_11895,N_11944);
or U12245 (N_12245,N_11894,N_11941);
or U12246 (N_12246,N_11859,N_11824);
and U12247 (N_12247,N_11982,N_11974);
and U12248 (N_12248,N_11943,N_11840);
and U12249 (N_12249,N_11875,N_11822);
nand U12250 (N_12250,N_12248,N_12023);
nor U12251 (N_12251,N_12028,N_12055);
and U12252 (N_12252,N_12136,N_12079);
xnor U12253 (N_12253,N_12194,N_12233);
or U12254 (N_12254,N_12169,N_12130);
and U12255 (N_12255,N_12060,N_12210);
nand U12256 (N_12256,N_12017,N_12190);
and U12257 (N_12257,N_12074,N_12120);
nand U12258 (N_12258,N_12051,N_12093);
nand U12259 (N_12259,N_12200,N_12228);
nand U12260 (N_12260,N_12087,N_12083);
nor U12261 (N_12261,N_12011,N_12167);
nor U12262 (N_12262,N_12149,N_12016);
xor U12263 (N_12263,N_12161,N_12242);
nor U12264 (N_12264,N_12088,N_12065);
and U12265 (N_12265,N_12125,N_12221);
and U12266 (N_12266,N_12072,N_12097);
xnor U12267 (N_12267,N_12177,N_12045);
nor U12268 (N_12268,N_12143,N_12212);
xnor U12269 (N_12269,N_12106,N_12195);
nor U12270 (N_12270,N_12135,N_12139);
or U12271 (N_12271,N_12246,N_12157);
xnor U12272 (N_12272,N_12064,N_12014);
or U12273 (N_12273,N_12176,N_12057);
or U12274 (N_12274,N_12213,N_12145);
nor U12275 (N_12275,N_12148,N_12008);
nor U12276 (N_12276,N_12129,N_12230);
nand U12277 (N_12277,N_12107,N_12225);
and U12278 (N_12278,N_12050,N_12199);
or U12279 (N_12279,N_12181,N_12010);
or U12280 (N_12280,N_12005,N_12049);
and U12281 (N_12281,N_12003,N_12207);
or U12282 (N_12282,N_12013,N_12142);
or U12283 (N_12283,N_12085,N_12175);
nor U12284 (N_12284,N_12162,N_12007);
and U12285 (N_12285,N_12193,N_12073);
xor U12286 (N_12286,N_12224,N_12096);
nand U12287 (N_12287,N_12211,N_12226);
or U12288 (N_12288,N_12025,N_12223);
nor U12289 (N_12289,N_12061,N_12119);
xor U12290 (N_12290,N_12189,N_12138);
nand U12291 (N_12291,N_12133,N_12184);
nor U12292 (N_12292,N_12070,N_12239);
and U12293 (N_12293,N_12063,N_12004);
and U12294 (N_12294,N_12044,N_12163);
xor U12295 (N_12295,N_12132,N_12171);
nor U12296 (N_12296,N_12056,N_12071);
and U12297 (N_12297,N_12147,N_12086);
nor U12298 (N_12298,N_12141,N_12066);
nand U12299 (N_12299,N_12216,N_12218);
nand U12300 (N_12300,N_12076,N_12240);
xnor U12301 (N_12301,N_12168,N_12227);
xnor U12302 (N_12302,N_12000,N_12179);
xnor U12303 (N_12303,N_12188,N_12117);
nand U12304 (N_12304,N_12234,N_12053);
and U12305 (N_12305,N_12123,N_12033);
nor U12306 (N_12306,N_12180,N_12155);
nand U12307 (N_12307,N_12182,N_12121);
and U12308 (N_12308,N_12206,N_12046);
xor U12309 (N_12309,N_12173,N_12116);
nand U12310 (N_12310,N_12222,N_12235);
nor U12311 (N_12311,N_12158,N_12219);
and U12312 (N_12312,N_12247,N_12144);
nand U12313 (N_12313,N_12178,N_12192);
and U12314 (N_12314,N_12040,N_12037);
and U12315 (N_12315,N_12203,N_12067);
nand U12316 (N_12316,N_12128,N_12112);
nor U12317 (N_12317,N_12183,N_12217);
nor U12318 (N_12318,N_12205,N_12196);
and U12319 (N_12319,N_12201,N_12156);
or U12320 (N_12320,N_12159,N_12202);
nor U12321 (N_12321,N_12100,N_12208);
nand U12322 (N_12322,N_12237,N_12024);
nand U12323 (N_12323,N_12187,N_12110);
and U12324 (N_12324,N_12164,N_12078);
nand U12325 (N_12325,N_12214,N_12172);
and U12326 (N_12326,N_12105,N_12036);
xnor U12327 (N_12327,N_12075,N_12041);
nor U12328 (N_12328,N_12101,N_12102);
and U12329 (N_12329,N_12027,N_12122);
and U12330 (N_12330,N_12244,N_12220);
or U12331 (N_12331,N_12094,N_12151);
xor U12332 (N_12332,N_12126,N_12099);
or U12333 (N_12333,N_12238,N_12204);
and U12334 (N_12334,N_12020,N_12131);
and U12335 (N_12335,N_12150,N_12080);
xnor U12336 (N_12336,N_12198,N_12029);
nor U12337 (N_12337,N_12209,N_12115);
nor U12338 (N_12338,N_12245,N_12006);
or U12339 (N_12339,N_12111,N_12215);
nand U12340 (N_12340,N_12113,N_12001);
nor U12341 (N_12341,N_12108,N_12054);
and U12342 (N_12342,N_12002,N_12134);
nand U12343 (N_12343,N_12160,N_12059);
xnor U12344 (N_12344,N_12166,N_12154);
xor U12345 (N_12345,N_12034,N_12229);
and U12346 (N_12346,N_12042,N_12243);
and U12347 (N_12347,N_12165,N_12035);
xnor U12348 (N_12348,N_12185,N_12236);
or U12349 (N_12349,N_12084,N_12058);
xor U12350 (N_12350,N_12174,N_12048);
xnor U12351 (N_12351,N_12038,N_12026);
xor U12352 (N_12352,N_12146,N_12077);
xnor U12353 (N_12353,N_12092,N_12047);
and U12354 (N_12354,N_12090,N_12015);
and U12355 (N_12355,N_12081,N_12140);
nor U12356 (N_12356,N_12104,N_12019);
nand U12357 (N_12357,N_12018,N_12091);
nor U12358 (N_12358,N_12127,N_12249);
xnor U12359 (N_12359,N_12232,N_12021);
xnor U12360 (N_12360,N_12191,N_12103);
and U12361 (N_12361,N_12114,N_12012);
and U12362 (N_12362,N_12062,N_12109);
nand U12363 (N_12363,N_12032,N_12186);
nand U12364 (N_12364,N_12241,N_12197);
xor U12365 (N_12365,N_12124,N_12068);
and U12366 (N_12366,N_12098,N_12089);
nor U12367 (N_12367,N_12043,N_12009);
nor U12368 (N_12368,N_12052,N_12153);
or U12369 (N_12369,N_12137,N_12030);
nand U12370 (N_12370,N_12031,N_12039);
nor U12371 (N_12371,N_12082,N_12118);
and U12372 (N_12372,N_12170,N_12069);
xnor U12373 (N_12373,N_12095,N_12152);
nand U12374 (N_12374,N_12022,N_12231);
and U12375 (N_12375,N_12231,N_12056);
nor U12376 (N_12376,N_12109,N_12162);
xor U12377 (N_12377,N_12154,N_12063);
nand U12378 (N_12378,N_12095,N_12242);
nor U12379 (N_12379,N_12238,N_12129);
nand U12380 (N_12380,N_12203,N_12189);
nor U12381 (N_12381,N_12092,N_12038);
nor U12382 (N_12382,N_12005,N_12219);
nor U12383 (N_12383,N_12009,N_12243);
nand U12384 (N_12384,N_12108,N_12049);
nand U12385 (N_12385,N_12102,N_12061);
nand U12386 (N_12386,N_12034,N_12187);
and U12387 (N_12387,N_12242,N_12142);
nand U12388 (N_12388,N_12195,N_12235);
xnor U12389 (N_12389,N_12113,N_12191);
xor U12390 (N_12390,N_12029,N_12244);
xnor U12391 (N_12391,N_12242,N_12127);
nor U12392 (N_12392,N_12058,N_12090);
and U12393 (N_12393,N_12174,N_12222);
or U12394 (N_12394,N_12073,N_12025);
nor U12395 (N_12395,N_12121,N_12034);
or U12396 (N_12396,N_12145,N_12036);
nor U12397 (N_12397,N_12031,N_12062);
nor U12398 (N_12398,N_12131,N_12133);
xnor U12399 (N_12399,N_12038,N_12132);
or U12400 (N_12400,N_12026,N_12201);
nand U12401 (N_12401,N_12046,N_12178);
xnor U12402 (N_12402,N_12019,N_12068);
xnor U12403 (N_12403,N_12165,N_12155);
and U12404 (N_12404,N_12194,N_12160);
or U12405 (N_12405,N_12098,N_12117);
xor U12406 (N_12406,N_12132,N_12175);
xnor U12407 (N_12407,N_12138,N_12020);
nand U12408 (N_12408,N_12158,N_12020);
nand U12409 (N_12409,N_12021,N_12240);
nand U12410 (N_12410,N_12164,N_12206);
and U12411 (N_12411,N_12003,N_12051);
nand U12412 (N_12412,N_12038,N_12195);
nor U12413 (N_12413,N_12051,N_12055);
nand U12414 (N_12414,N_12177,N_12111);
nor U12415 (N_12415,N_12112,N_12030);
or U12416 (N_12416,N_12103,N_12199);
xnor U12417 (N_12417,N_12054,N_12196);
nand U12418 (N_12418,N_12170,N_12203);
or U12419 (N_12419,N_12043,N_12108);
and U12420 (N_12420,N_12203,N_12044);
xnor U12421 (N_12421,N_12033,N_12095);
and U12422 (N_12422,N_12247,N_12118);
nand U12423 (N_12423,N_12178,N_12019);
or U12424 (N_12424,N_12153,N_12172);
nor U12425 (N_12425,N_12000,N_12149);
nor U12426 (N_12426,N_12206,N_12160);
nor U12427 (N_12427,N_12157,N_12033);
xor U12428 (N_12428,N_12173,N_12084);
or U12429 (N_12429,N_12138,N_12003);
nand U12430 (N_12430,N_12213,N_12219);
nor U12431 (N_12431,N_12078,N_12117);
xnor U12432 (N_12432,N_12214,N_12108);
xnor U12433 (N_12433,N_12186,N_12048);
and U12434 (N_12434,N_12001,N_12099);
nor U12435 (N_12435,N_12031,N_12023);
or U12436 (N_12436,N_12219,N_12249);
or U12437 (N_12437,N_12016,N_12039);
xnor U12438 (N_12438,N_12050,N_12041);
xnor U12439 (N_12439,N_12224,N_12245);
nand U12440 (N_12440,N_12230,N_12013);
or U12441 (N_12441,N_12202,N_12119);
xor U12442 (N_12442,N_12009,N_12127);
nor U12443 (N_12443,N_12211,N_12198);
or U12444 (N_12444,N_12064,N_12196);
nor U12445 (N_12445,N_12247,N_12189);
nand U12446 (N_12446,N_12196,N_12006);
nand U12447 (N_12447,N_12044,N_12154);
nor U12448 (N_12448,N_12148,N_12053);
or U12449 (N_12449,N_12222,N_12011);
xnor U12450 (N_12450,N_12143,N_12187);
and U12451 (N_12451,N_12208,N_12119);
and U12452 (N_12452,N_12123,N_12144);
or U12453 (N_12453,N_12084,N_12249);
nand U12454 (N_12454,N_12139,N_12218);
xor U12455 (N_12455,N_12160,N_12228);
xnor U12456 (N_12456,N_12035,N_12049);
nor U12457 (N_12457,N_12041,N_12109);
or U12458 (N_12458,N_12027,N_12045);
nor U12459 (N_12459,N_12193,N_12133);
and U12460 (N_12460,N_12118,N_12071);
and U12461 (N_12461,N_12147,N_12023);
xnor U12462 (N_12462,N_12033,N_12205);
xor U12463 (N_12463,N_12100,N_12216);
nor U12464 (N_12464,N_12188,N_12082);
nor U12465 (N_12465,N_12224,N_12225);
nand U12466 (N_12466,N_12136,N_12033);
and U12467 (N_12467,N_12088,N_12146);
nand U12468 (N_12468,N_12027,N_12200);
nand U12469 (N_12469,N_12243,N_12006);
xnor U12470 (N_12470,N_12170,N_12003);
xnor U12471 (N_12471,N_12073,N_12016);
and U12472 (N_12472,N_12175,N_12233);
nor U12473 (N_12473,N_12232,N_12198);
or U12474 (N_12474,N_12237,N_12010);
and U12475 (N_12475,N_12162,N_12244);
nor U12476 (N_12476,N_12204,N_12236);
nor U12477 (N_12477,N_12068,N_12010);
nor U12478 (N_12478,N_12000,N_12068);
nor U12479 (N_12479,N_12095,N_12093);
nor U12480 (N_12480,N_12114,N_12053);
nand U12481 (N_12481,N_12083,N_12221);
and U12482 (N_12482,N_12036,N_12127);
nand U12483 (N_12483,N_12122,N_12102);
xnor U12484 (N_12484,N_12224,N_12006);
or U12485 (N_12485,N_12133,N_12012);
nor U12486 (N_12486,N_12117,N_12069);
nand U12487 (N_12487,N_12145,N_12164);
and U12488 (N_12488,N_12246,N_12152);
and U12489 (N_12489,N_12019,N_12214);
nor U12490 (N_12490,N_12051,N_12045);
nor U12491 (N_12491,N_12088,N_12059);
and U12492 (N_12492,N_12138,N_12191);
and U12493 (N_12493,N_12019,N_12230);
and U12494 (N_12494,N_12032,N_12111);
nor U12495 (N_12495,N_12084,N_12055);
xnor U12496 (N_12496,N_12009,N_12197);
nand U12497 (N_12497,N_12165,N_12218);
or U12498 (N_12498,N_12002,N_12164);
nor U12499 (N_12499,N_12202,N_12151);
or U12500 (N_12500,N_12474,N_12276);
nor U12501 (N_12501,N_12371,N_12435);
or U12502 (N_12502,N_12291,N_12409);
nand U12503 (N_12503,N_12282,N_12317);
nand U12504 (N_12504,N_12436,N_12407);
or U12505 (N_12505,N_12412,N_12417);
nand U12506 (N_12506,N_12283,N_12419);
and U12507 (N_12507,N_12385,N_12482);
or U12508 (N_12508,N_12405,N_12457);
nor U12509 (N_12509,N_12493,N_12349);
xnor U12510 (N_12510,N_12354,N_12494);
and U12511 (N_12511,N_12321,N_12280);
nor U12512 (N_12512,N_12447,N_12341);
nor U12513 (N_12513,N_12431,N_12265);
or U12514 (N_12514,N_12414,N_12350);
and U12515 (N_12515,N_12468,N_12355);
nand U12516 (N_12516,N_12325,N_12364);
nor U12517 (N_12517,N_12342,N_12296);
or U12518 (N_12518,N_12346,N_12288);
and U12519 (N_12519,N_12281,N_12471);
or U12520 (N_12520,N_12467,N_12393);
and U12521 (N_12521,N_12279,N_12255);
xnor U12522 (N_12522,N_12290,N_12319);
nor U12523 (N_12523,N_12466,N_12392);
and U12524 (N_12524,N_12488,N_12318);
or U12525 (N_12525,N_12388,N_12332);
or U12526 (N_12526,N_12361,N_12453);
and U12527 (N_12527,N_12401,N_12335);
or U12528 (N_12528,N_12334,N_12433);
nor U12529 (N_12529,N_12261,N_12254);
nand U12530 (N_12530,N_12438,N_12399);
xor U12531 (N_12531,N_12495,N_12472);
xor U12532 (N_12532,N_12292,N_12287);
xor U12533 (N_12533,N_12340,N_12357);
or U12534 (N_12534,N_12397,N_12420);
nor U12535 (N_12535,N_12330,N_12286);
xor U12536 (N_12536,N_12404,N_12383);
and U12537 (N_12537,N_12490,N_12382);
or U12538 (N_12538,N_12285,N_12267);
xor U12539 (N_12539,N_12402,N_12400);
nand U12540 (N_12540,N_12273,N_12336);
nor U12541 (N_12541,N_12456,N_12415);
nand U12542 (N_12542,N_12394,N_12459);
nand U12543 (N_12543,N_12251,N_12499);
and U12544 (N_12544,N_12464,N_12268);
nand U12545 (N_12545,N_12485,N_12311);
nor U12546 (N_12546,N_12316,N_12338);
or U12547 (N_12547,N_12295,N_12387);
xnor U12548 (N_12548,N_12305,N_12367);
or U12549 (N_12549,N_12437,N_12439);
nor U12550 (N_12550,N_12374,N_12372);
nand U12551 (N_12551,N_12449,N_12398);
nor U12552 (N_12552,N_12284,N_12395);
nor U12553 (N_12553,N_12263,N_12358);
nand U12554 (N_12554,N_12379,N_12377);
or U12555 (N_12555,N_12496,N_12376);
nand U12556 (N_12556,N_12324,N_12454);
or U12557 (N_12557,N_12270,N_12298);
or U12558 (N_12558,N_12486,N_12362);
nand U12559 (N_12559,N_12356,N_12301);
nor U12560 (N_12560,N_12252,N_12473);
and U12561 (N_12561,N_12380,N_12333);
nor U12562 (N_12562,N_12422,N_12312);
and U12563 (N_12563,N_12443,N_12299);
xor U12564 (N_12564,N_12363,N_12329);
or U12565 (N_12565,N_12497,N_12462);
and U12566 (N_12566,N_12348,N_12479);
or U12567 (N_12567,N_12411,N_12476);
or U12568 (N_12568,N_12487,N_12257);
xnor U12569 (N_12569,N_12424,N_12300);
nor U12570 (N_12570,N_12271,N_12421);
and U12571 (N_12571,N_12322,N_12423);
or U12572 (N_12572,N_12430,N_12458);
nand U12573 (N_12573,N_12347,N_12306);
or U12574 (N_12574,N_12278,N_12396);
xor U12575 (N_12575,N_12337,N_12492);
or U12576 (N_12576,N_12410,N_12266);
nor U12577 (N_12577,N_12386,N_12277);
and U12578 (N_12578,N_12343,N_12352);
xnor U12579 (N_12579,N_12275,N_12432);
xor U12580 (N_12580,N_12408,N_12368);
nand U12581 (N_12581,N_12308,N_12480);
nand U12582 (N_12582,N_12470,N_12264);
nand U12583 (N_12583,N_12302,N_12307);
xor U12584 (N_12584,N_12429,N_12323);
or U12585 (N_12585,N_12272,N_12460);
nand U12586 (N_12586,N_12403,N_12451);
or U12587 (N_12587,N_12293,N_12446);
xnor U12588 (N_12588,N_12310,N_12259);
nor U12589 (N_12589,N_12445,N_12274);
nand U12590 (N_12590,N_12331,N_12304);
nand U12591 (N_12591,N_12384,N_12250);
and U12592 (N_12592,N_12389,N_12426);
or U12593 (N_12593,N_12294,N_12327);
and U12594 (N_12594,N_12303,N_12351);
nor U12595 (N_12595,N_12491,N_12469);
and U12596 (N_12596,N_12378,N_12434);
nor U12597 (N_12597,N_12258,N_12328);
xnor U12598 (N_12598,N_12381,N_12314);
and U12599 (N_12599,N_12326,N_12309);
nand U12600 (N_12600,N_12440,N_12484);
xor U12601 (N_12601,N_12289,N_12260);
and U12602 (N_12602,N_12253,N_12269);
or U12603 (N_12603,N_12418,N_12360);
and U12604 (N_12604,N_12413,N_12320);
nand U12605 (N_12605,N_12373,N_12465);
nand U12606 (N_12606,N_12416,N_12481);
nand U12607 (N_12607,N_12313,N_12444);
xnor U12608 (N_12608,N_12428,N_12461);
and U12609 (N_12609,N_12262,N_12297);
nor U12610 (N_12610,N_12498,N_12475);
xor U12611 (N_12611,N_12375,N_12448);
xnor U12612 (N_12612,N_12425,N_12463);
and U12613 (N_12613,N_12353,N_12406);
or U12614 (N_12614,N_12478,N_12366);
and U12615 (N_12615,N_12370,N_12427);
nor U12616 (N_12616,N_12359,N_12477);
nor U12617 (N_12617,N_12369,N_12442);
nor U12618 (N_12618,N_12489,N_12315);
nor U12619 (N_12619,N_12344,N_12390);
nor U12620 (N_12620,N_12455,N_12483);
and U12621 (N_12621,N_12441,N_12452);
nor U12622 (N_12622,N_12345,N_12339);
and U12623 (N_12623,N_12391,N_12365);
or U12624 (N_12624,N_12256,N_12450);
or U12625 (N_12625,N_12304,N_12484);
or U12626 (N_12626,N_12310,N_12398);
and U12627 (N_12627,N_12459,N_12432);
nor U12628 (N_12628,N_12423,N_12328);
xor U12629 (N_12629,N_12302,N_12484);
or U12630 (N_12630,N_12483,N_12381);
nor U12631 (N_12631,N_12421,N_12316);
or U12632 (N_12632,N_12493,N_12358);
nand U12633 (N_12633,N_12423,N_12418);
nand U12634 (N_12634,N_12289,N_12431);
and U12635 (N_12635,N_12480,N_12369);
nand U12636 (N_12636,N_12388,N_12457);
or U12637 (N_12637,N_12289,N_12297);
or U12638 (N_12638,N_12325,N_12499);
xnor U12639 (N_12639,N_12376,N_12400);
or U12640 (N_12640,N_12304,N_12483);
or U12641 (N_12641,N_12383,N_12352);
and U12642 (N_12642,N_12480,N_12327);
or U12643 (N_12643,N_12356,N_12331);
nor U12644 (N_12644,N_12348,N_12265);
and U12645 (N_12645,N_12391,N_12301);
or U12646 (N_12646,N_12452,N_12402);
nand U12647 (N_12647,N_12473,N_12387);
nor U12648 (N_12648,N_12442,N_12493);
xor U12649 (N_12649,N_12411,N_12250);
or U12650 (N_12650,N_12399,N_12387);
xnor U12651 (N_12651,N_12378,N_12383);
or U12652 (N_12652,N_12498,N_12427);
nor U12653 (N_12653,N_12364,N_12288);
nor U12654 (N_12654,N_12456,N_12485);
and U12655 (N_12655,N_12325,N_12274);
nor U12656 (N_12656,N_12452,N_12377);
and U12657 (N_12657,N_12498,N_12285);
and U12658 (N_12658,N_12306,N_12377);
xor U12659 (N_12659,N_12372,N_12319);
or U12660 (N_12660,N_12357,N_12415);
xor U12661 (N_12661,N_12331,N_12254);
nand U12662 (N_12662,N_12412,N_12487);
or U12663 (N_12663,N_12332,N_12294);
nand U12664 (N_12664,N_12297,N_12439);
nor U12665 (N_12665,N_12400,N_12385);
xnor U12666 (N_12666,N_12465,N_12442);
and U12667 (N_12667,N_12474,N_12343);
nand U12668 (N_12668,N_12255,N_12379);
xor U12669 (N_12669,N_12377,N_12260);
nor U12670 (N_12670,N_12366,N_12467);
xnor U12671 (N_12671,N_12493,N_12260);
xor U12672 (N_12672,N_12253,N_12400);
nor U12673 (N_12673,N_12472,N_12480);
and U12674 (N_12674,N_12360,N_12494);
nand U12675 (N_12675,N_12256,N_12422);
or U12676 (N_12676,N_12306,N_12490);
nor U12677 (N_12677,N_12365,N_12264);
nand U12678 (N_12678,N_12339,N_12272);
nand U12679 (N_12679,N_12475,N_12410);
nand U12680 (N_12680,N_12360,N_12479);
or U12681 (N_12681,N_12462,N_12391);
nor U12682 (N_12682,N_12468,N_12333);
and U12683 (N_12683,N_12433,N_12362);
nor U12684 (N_12684,N_12277,N_12446);
xor U12685 (N_12685,N_12422,N_12317);
xnor U12686 (N_12686,N_12404,N_12405);
or U12687 (N_12687,N_12268,N_12495);
nand U12688 (N_12688,N_12466,N_12296);
xor U12689 (N_12689,N_12330,N_12446);
and U12690 (N_12690,N_12315,N_12410);
nor U12691 (N_12691,N_12446,N_12360);
or U12692 (N_12692,N_12355,N_12410);
nand U12693 (N_12693,N_12437,N_12404);
xor U12694 (N_12694,N_12335,N_12353);
nand U12695 (N_12695,N_12480,N_12407);
or U12696 (N_12696,N_12449,N_12293);
and U12697 (N_12697,N_12384,N_12317);
xor U12698 (N_12698,N_12289,N_12377);
nor U12699 (N_12699,N_12370,N_12410);
nand U12700 (N_12700,N_12343,N_12359);
and U12701 (N_12701,N_12451,N_12261);
or U12702 (N_12702,N_12427,N_12257);
nand U12703 (N_12703,N_12288,N_12262);
or U12704 (N_12704,N_12265,N_12435);
nand U12705 (N_12705,N_12253,N_12282);
xor U12706 (N_12706,N_12376,N_12395);
or U12707 (N_12707,N_12276,N_12262);
xnor U12708 (N_12708,N_12374,N_12426);
and U12709 (N_12709,N_12290,N_12357);
or U12710 (N_12710,N_12301,N_12293);
nand U12711 (N_12711,N_12292,N_12334);
nand U12712 (N_12712,N_12351,N_12376);
xnor U12713 (N_12713,N_12469,N_12421);
nor U12714 (N_12714,N_12474,N_12394);
nor U12715 (N_12715,N_12368,N_12379);
nand U12716 (N_12716,N_12461,N_12466);
xnor U12717 (N_12717,N_12334,N_12333);
or U12718 (N_12718,N_12497,N_12411);
or U12719 (N_12719,N_12372,N_12359);
nor U12720 (N_12720,N_12293,N_12364);
or U12721 (N_12721,N_12369,N_12450);
nor U12722 (N_12722,N_12329,N_12287);
and U12723 (N_12723,N_12251,N_12344);
or U12724 (N_12724,N_12490,N_12360);
xnor U12725 (N_12725,N_12307,N_12361);
or U12726 (N_12726,N_12330,N_12378);
and U12727 (N_12727,N_12454,N_12372);
and U12728 (N_12728,N_12426,N_12456);
and U12729 (N_12729,N_12352,N_12472);
xnor U12730 (N_12730,N_12384,N_12466);
and U12731 (N_12731,N_12254,N_12324);
nor U12732 (N_12732,N_12479,N_12449);
nor U12733 (N_12733,N_12339,N_12353);
xnor U12734 (N_12734,N_12367,N_12470);
nor U12735 (N_12735,N_12361,N_12330);
xor U12736 (N_12736,N_12322,N_12356);
nand U12737 (N_12737,N_12360,N_12457);
and U12738 (N_12738,N_12267,N_12310);
xor U12739 (N_12739,N_12406,N_12447);
nand U12740 (N_12740,N_12389,N_12320);
xor U12741 (N_12741,N_12471,N_12455);
and U12742 (N_12742,N_12422,N_12340);
and U12743 (N_12743,N_12358,N_12391);
xnor U12744 (N_12744,N_12405,N_12353);
xnor U12745 (N_12745,N_12354,N_12460);
nor U12746 (N_12746,N_12318,N_12461);
and U12747 (N_12747,N_12409,N_12317);
nor U12748 (N_12748,N_12407,N_12401);
or U12749 (N_12749,N_12392,N_12292);
xor U12750 (N_12750,N_12654,N_12502);
xor U12751 (N_12751,N_12555,N_12665);
xor U12752 (N_12752,N_12634,N_12711);
or U12753 (N_12753,N_12676,N_12704);
or U12754 (N_12754,N_12726,N_12590);
nand U12755 (N_12755,N_12549,N_12699);
nand U12756 (N_12756,N_12743,N_12658);
xnor U12757 (N_12757,N_12526,N_12522);
and U12758 (N_12758,N_12523,N_12672);
xor U12759 (N_12759,N_12521,N_12524);
or U12760 (N_12760,N_12663,N_12749);
and U12761 (N_12761,N_12547,N_12705);
xor U12762 (N_12762,N_12735,N_12595);
nand U12763 (N_12763,N_12715,N_12566);
and U12764 (N_12764,N_12694,N_12732);
nand U12765 (N_12765,N_12510,N_12660);
and U12766 (N_12766,N_12557,N_12613);
or U12767 (N_12767,N_12575,N_12655);
nand U12768 (N_12768,N_12603,N_12721);
or U12769 (N_12769,N_12697,N_12629);
nand U12770 (N_12770,N_12625,N_12572);
or U12771 (N_12771,N_12618,N_12644);
nand U12772 (N_12772,N_12546,N_12611);
nand U12773 (N_12773,N_12543,N_12628);
or U12774 (N_12774,N_12552,N_12666);
nand U12775 (N_12775,N_12633,N_12545);
or U12776 (N_12776,N_12563,N_12738);
nand U12777 (N_12777,N_12703,N_12648);
xnor U12778 (N_12778,N_12667,N_12548);
or U12779 (N_12779,N_12560,N_12740);
xnor U12780 (N_12780,N_12737,N_12573);
xnor U12781 (N_12781,N_12541,N_12592);
nor U12782 (N_12782,N_12527,N_12559);
nor U12783 (N_12783,N_12723,N_12554);
nor U12784 (N_12784,N_12535,N_12561);
and U12785 (N_12785,N_12639,N_12649);
nor U12786 (N_12786,N_12605,N_12585);
or U12787 (N_12787,N_12696,N_12617);
and U12788 (N_12788,N_12578,N_12693);
nor U12789 (N_12789,N_12712,N_12651);
or U12790 (N_12790,N_12690,N_12642);
nor U12791 (N_12791,N_12565,N_12681);
xor U12792 (N_12792,N_12626,N_12708);
or U12793 (N_12793,N_12653,N_12632);
and U12794 (N_12794,N_12731,N_12505);
nand U12795 (N_12795,N_12587,N_12730);
nand U12796 (N_12796,N_12706,N_12677);
and U12797 (N_12797,N_12729,N_12602);
and U12798 (N_12798,N_12601,N_12727);
and U12799 (N_12799,N_12519,N_12586);
and U12800 (N_12800,N_12577,N_12668);
xnor U12801 (N_12801,N_12645,N_12584);
nand U12802 (N_12802,N_12513,N_12511);
nand U12803 (N_12803,N_12725,N_12722);
nor U12804 (N_12804,N_12536,N_12698);
xor U12805 (N_12805,N_12685,N_12701);
nand U12806 (N_12806,N_12564,N_12744);
nand U12807 (N_12807,N_12646,N_12673);
xor U12808 (N_12808,N_12678,N_12579);
xnor U12809 (N_12809,N_12692,N_12643);
nand U12810 (N_12810,N_12571,N_12717);
nor U12811 (N_12811,N_12518,N_12627);
xnor U12812 (N_12812,N_12707,N_12512);
nor U12813 (N_12813,N_12604,N_12500);
or U12814 (N_12814,N_12533,N_12616);
nor U12815 (N_12815,N_12550,N_12599);
nand U12816 (N_12816,N_12675,N_12635);
xor U12817 (N_12817,N_12733,N_12637);
or U12818 (N_12818,N_12719,N_12583);
xnor U12819 (N_12819,N_12624,N_12542);
nor U12820 (N_12820,N_12537,N_12539);
and U12821 (N_12821,N_12664,N_12695);
and U12822 (N_12822,N_12679,N_12640);
nor U12823 (N_12823,N_12680,N_12503);
and U12824 (N_12824,N_12615,N_12558);
nor U12825 (N_12825,N_12588,N_12638);
xnor U12826 (N_12826,N_12714,N_12623);
and U12827 (N_12827,N_12568,N_12538);
nor U12828 (N_12828,N_12607,N_12650);
and U12829 (N_12829,N_12534,N_12562);
nand U12830 (N_12830,N_12569,N_12508);
xnor U12831 (N_12831,N_12591,N_12532);
nor U12832 (N_12832,N_12619,N_12631);
nand U12833 (N_12833,N_12593,N_12504);
nand U12834 (N_12834,N_12580,N_12641);
xor U12835 (N_12835,N_12520,N_12606);
and U12836 (N_12836,N_12556,N_12509);
and U12837 (N_12837,N_12576,N_12530);
nor U12838 (N_12838,N_12745,N_12620);
nand U12839 (N_12839,N_12670,N_12516);
nand U12840 (N_12840,N_12669,N_12728);
nor U12841 (N_12841,N_12581,N_12621);
or U12842 (N_12842,N_12596,N_12736);
nand U12843 (N_12843,N_12531,N_12691);
or U12844 (N_12844,N_12540,N_12501);
or U12845 (N_12845,N_12724,N_12567);
or U12846 (N_12846,N_12684,N_12570);
and U12847 (N_12847,N_12529,N_12718);
and U12848 (N_12848,N_12742,N_12674);
nand U12849 (N_12849,N_12702,N_12528);
nor U12850 (N_12850,N_12506,N_12515);
and U12851 (N_12851,N_12636,N_12657);
nor U12852 (N_12852,N_12716,N_12746);
and U12853 (N_12853,N_12514,N_12507);
nor U12854 (N_12854,N_12747,N_12574);
nand U12855 (N_12855,N_12659,N_12748);
nand U12856 (N_12856,N_12734,N_12652);
nand U12857 (N_12857,N_12709,N_12525);
and U12858 (N_12858,N_12700,N_12689);
nand U12859 (N_12859,N_12594,N_12608);
nor U12860 (N_12860,N_12662,N_12622);
nand U12861 (N_12861,N_12582,N_12656);
and U12862 (N_12862,N_12741,N_12589);
xor U12863 (N_12863,N_12553,N_12686);
nand U12864 (N_12864,N_12710,N_12614);
nand U12865 (N_12865,N_12610,N_12661);
nor U12866 (N_12866,N_12671,N_12687);
and U12867 (N_12867,N_12551,N_12683);
nor U12868 (N_12868,N_12739,N_12600);
xnor U12869 (N_12869,N_12597,N_12647);
or U12870 (N_12870,N_12517,N_12688);
xor U12871 (N_12871,N_12720,N_12713);
nor U12872 (N_12872,N_12598,N_12682);
nand U12873 (N_12873,N_12612,N_12609);
nand U12874 (N_12874,N_12630,N_12544);
nor U12875 (N_12875,N_12615,N_12702);
xor U12876 (N_12876,N_12710,N_12560);
or U12877 (N_12877,N_12641,N_12706);
or U12878 (N_12878,N_12692,N_12602);
nand U12879 (N_12879,N_12584,N_12608);
or U12880 (N_12880,N_12543,N_12526);
xor U12881 (N_12881,N_12718,N_12621);
or U12882 (N_12882,N_12587,N_12652);
xnor U12883 (N_12883,N_12692,N_12703);
nand U12884 (N_12884,N_12715,N_12659);
or U12885 (N_12885,N_12732,N_12718);
nand U12886 (N_12886,N_12595,N_12524);
xnor U12887 (N_12887,N_12666,N_12557);
and U12888 (N_12888,N_12713,N_12562);
nor U12889 (N_12889,N_12560,N_12515);
nand U12890 (N_12890,N_12723,N_12570);
xor U12891 (N_12891,N_12639,N_12509);
xor U12892 (N_12892,N_12671,N_12697);
nor U12893 (N_12893,N_12570,N_12542);
nor U12894 (N_12894,N_12588,N_12537);
and U12895 (N_12895,N_12651,N_12505);
nor U12896 (N_12896,N_12703,N_12541);
nand U12897 (N_12897,N_12673,N_12548);
or U12898 (N_12898,N_12586,N_12582);
xnor U12899 (N_12899,N_12711,N_12534);
or U12900 (N_12900,N_12717,N_12583);
and U12901 (N_12901,N_12701,N_12510);
or U12902 (N_12902,N_12592,N_12550);
xnor U12903 (N_12903,N_12619,N_12731);
or U12904 (N_12904,N_12747,N_12675);
nand U12905 (N_12905,N_12712,N_12538);
nand U12906 (N_12906,N_12558,N_12629);
xnor U12907 (N_12907,N_12645,N_12637);
and U12908 (N_12908,N_12672,N_12508);
or U12909 (N_12909,N_12617,N_12701);
or U12910 (N_12910,N_12579,N_12654);
nor U12911 (N_12911,N_12502,N_12605);
xnor U12912 (N_12912,N_12712,N_12632);
nor U12913 (N_12913,N_12540,N_12705);
nand U12914 (N_12914,N_12679,N_12520);
xnor U12915 (N_12915,N_12567,N_12746);
and U12916 (N_12916,N_12584,N_12576);
nor U12917 (N_12917,N_12667,N_12513);
nor U12918 (N_12918,N_12596,N_12578);
and U12919 (N_12919,N_12591,N_12692);
nor U12920 (N_12920,N_12709,N_12500);
and U12921 (N_12921,N_12610,N_12552);
and U12922 (N_12922,N_12615,N_12710);
xnor U12923 (N_12923,N_12652,N_12677);
nor U12924 (N_12924,N_12685,N_12545);
or U12925 (N_12925,N_12522,N_12587);
nor U12926 (N_12926,N_12540,N_12586);
and U12927 (N_12927,N_12568,N_12506);
or U12928 (N_12928,N_12749,N_12569);
nand U12929 (N_12929,N_12597,N_12571);
nand U12930 (N_12930,N_12516,N_12567);
nand U12931 (N_12931,N_12714,N_12577);
or U12932 (N_12932,N_12628,N_12721);
nor U12933 (N_12933,N_12730,N_12612);
nor U12934 (N_12934,N_12511,N_12685);
nor U12935 (N_12935,N_12746,N_12516);
xor U12936 (N_12936,N_12739,N_12717);
nand U12937 (N_12937,N_12740,N_12554);
xnor U12938 (N_12938,N_12502,N_12626);
nand U12939 (N_12939,N_12612,N_12617);
nand U12940 (N_12940,N_12539,N_12511);
or U12941 (N_12941,N_12740,N_12645);
and U12942 (N_12942,N_12733,N_12707);
nand U12943 (N_12943,N_12582,N_12615);
and U12944 (N_12944,N_12658,N_12687);
nor U12945 (N_12945,N_12654,N_12657);
and U12946 (N_12946,N_12743,N_12746);
or U12947 (N_12947,N_12609,N_12549);
nor U12948 (N_12948,N_12520,N_12542);
or U12949 (N_12949,N_12652,N_12612);
or U12950 (N_12950,N_12741,N_12650);
xor U12951 (N_12951,N_12694,N_12661);
and U12952 (N_12952,N_12735,N_12699);
nand U12953 (N_12953,N_12649,N_12603);
xor U12954 (N_12954,N_12725,N_12583);
xor U12955 (N_12955,N_12715,N_12592);
nor U12956 (N_12956,N_12512,N_12633);
and U12957 (N_12957,N_12596,N_12558);
nor U12958 (N_12958,N_12584,N_12595);
nor U12959 (N_12959,N_12523,N_12602);
xnor U12960 (N_12960,N_12706,N_12704);
nor U12961 (N_12961,N_12554,N_12742);
and U12962 (N_12962,N_12597,N_12742);
or U12963 (N_12963,N_12619,N_12672);
or U12964 (N_12964,N_12673,N_12695);
xnor U12965 (N_12965,N_12719,N_12581);
and U12966 (N_12966,N_12747,N_12714);
nor U12967 (N_12967,N_12740,N_12697);
and U12968 (N_12968,N_12749,N_12697);
nor U12969 (N_12969,N_12686,N_12592);
nor U12970 (N_12970,N_12545,N_12566);
nand U12971 (N_12971,N_12526,N_12567);
nand U12972 (N_12972,N_12654,N_12676);
nor U12973 (N_12973,N_12654,N_12573);
or U12974 (N_12974,N_12509,N_12576);
xnor U12975 (N_12975,N_12590,N_12584);
or U12976 (N_12976,N_12681,N_12670);
and U12977 (N_12977,N_12612,N_12742);
and U12978 (N_12978,N_12699,N_12500);
nor U12979 (N_12979,N_12728,N_12722);
nand U12980 (N_12980,N_12729,N_12682);
nand U12981 (N_12981,N_12561,N_12522);
and U12982 (N_12982,N_12618,N_12514);
or U12983 (N_12983,N_12656,N_12654);
and U12984 (N_12984,N_12729,N_12592);
or U12985 (N_12985,N_12725,N_12614);
and U12986 (N_12986,N_12558,N_12716);
and U12987 (N_12987,N_12669,N_12642);
nand U12988 (N_12988,N_12606,N_12688);
nor U12989 (N_12989,N_12710,N_12598);
nor U12990 (N_12990,N_12636,N_12713);
or U12991 (N_12991,N_12608,N_12732);
xnor U12992 (N_12992,N_12745,N_12584);
xor U12993 (N_12993,N_12530,N_12594);
and U12994 (N_12994,N_12559,N_12586);
nand U12995 (N_12995,N_12737,N_12533);
and U12996 (N_12996,N_12597,N_12627);
xnor U12997 (N_12997,N_12714,N_12592);
nand U12998 (N_12998,N_12709,N_12570);
and U12999 (N_12999,N_12616,N_12658);
or U13000 (N_13000,N_12877,N_12995);
or U13001 (N_13001,N_12912,N_12874);
nor U13002 (N_13002,N_12892,N_12868);
and U13003 (N_13003,N_12969,N_12913);
or U13004 (N_13004,N_12769,N_12805);
and U13005 (N_13005,N_12800,N_12860);
nand U13006 (N_13006,N_12859,N_12854);
xnor U13007 (N_13007,N_12937,N_12793);
xor U13008 (N_13008,N_12974,N_12938);
nand U13009 (N_13009,N_12753,N_12960);
nand U13010 (N_13010,N_12849,N_12762);
nor U13011 (N_13011,N_12818,N_12889);
or U13012 (N_13012,N_12799,N_12878);
or U13013 (N_13013,N_12923,N_12829);
and U13014 (N_13014,N_12750,N_12816);
or U13015 (N_13015,N_12949,N_12803);
xnor U13016 (N_13016,N_12774,N_12837);
nor U13017 (N_13017,N_12756,N_12861);
nand U13018 (N_13018,N_12842,N_12789);
or U13019 (N_13019,N_12754,N_12939);
or U13020 (N_13020,N_12882,N_12914);
nor U13021 (N_13021,N_12944,N_12844);
nand U13022 (N_13022,N_12867,N_12802);
xnor U13023 (N_13023,N_12973,N_12951);
xor U13024 (N_13024,N_12831,N_12903);
or U13025 (N_13025,N_12898,N_12808);
or U13026 (N_13026,N_12847,N_12791);
nand U13027 (N_13027,N_12876,N_12872);
xor U13028 (N_13028,N_12947,N_12982);
nand U13029 (N_13029,N_12920,N_12921);
xnor U13030 (N_13030,N_12776,N_12865);
or U13031 (N_13031,N_12996,N_12993);
and U13032 (N_13032,N_12955,N_12991);
nand U13033 (N_13033,N_12824,N_12935);
nor U13034 (N_13034,N_12922,N_12948);
nand U13035 (N_13035,N_12907,N_12959);
or U13036 (N_13036,N_12839,N_12786);
and U13037 (N_13037,N_12883,N_12887);
nand U13038 (N_13038,N_12811,N_12886);
or U13039 (N_13039,N_12975,N_12813);
nor U13040 (N_13040,N_12751,N_12945);
or U13041 (N_13041,N_12843,N_12930);
nand U13042 (N_13042,N_12788,N_12804);
nor U13043 (N_13043,N_12881,N_12807);
and U13044 (N_13044,N_12798,N_12950);
nor U13045 (N_13045,N_12835,N_12984);
nand U13046 (N_13046,N_12992,N_12761);
xor U13047 (N_13047,N_12820,N_12927);
and U13048 (N_13048,N_12862,N_12891);
and U13049 (N_13049,N_12833,N_12760);
xor U13050 (N_13050,N_12954,N_12780);
nand U13051 (N_13051,N_12880,N_12787);
xnor U13052 (N_13052,N_12968,N_12775);
nand U13053 (N_13053,N_12896,N_12879);
nand U13054 (N_13054,N_12875,N_12997);
nand U13055 (N_13055,N_12953,N_12848);
and U13056 (N_13056,N_12925,N_12773);
xnor U13057 (N_13057,N_12758,N_12976);
xor U13058 (N_13058,N_12916,N_12797);
and U13059 (N_13059,N_12755,N_12885);
and U13060 (N_13060,N_12770,N_12785);
nand U13061 (N_13061,N_12765,N_12817);
nor U13062 (N_13062,N_12956,N_12772);
or U13063 (N_13063,N_12764,N_12928);
or U13064 (N_13064,N_12926,N_12863);
nand U13065 (N_13065,N_12917,N_12890);
and U13066 (N_13066,N_12819,N_12857);
or U13067 (N_13067,N_12792,N_12790);
and U13068 (N_13068,N_12958,N_12981);
xor U13069 (N_13069,N_12782,N_12894);
xor U13070 (N_13070,N_12919,N_12888);
nand U13071 (N_13071,N_12986,N_12961);
and U13072 (N_13072,N_12871,N_12910);
nand U13073 (N_13073,N_12994,N_12906);
xnor U13074 (N_13074,N_12943,N_12822);
xor U13075 (N_13075,N_12964,N_12941);
and U13076 (N_13076,N_12853,N_12884);
nor U13077 (N_13077,N_12856,N_12825);
nand U13078 (N_13078,N_12987,N_12971);
nand U13079 (N_13079,N_12779,N_12942);
xor U13080 (N_13080,N_12983,N_12827);
nand U13081 (N_13081,N_12936,N_12781);
nand U13082 (N_13082,N_12940,N_12977);
xor U13083 (N_13083,N_12757,N_12897);
nor U13084 (N_13084,N_12957,N_12900);
xnor U13085 (N_13085,N_12909,N_12929);
and U13086 (N_13086,N_12858,N_12759);
and U13087 (N_13087,N_12998,N_12836);
and U13088 (N_13088,N_12794,N_12767);
and U13089 (N_13089,N_12931,N_12989);
xnor U13090 (N_13090,N_12915,N_12852);
xor U13091 (N_13091,N_12873,N_12905);
nor U13092 (N_13092,N_12895,N_12933);
and U13093 (N_13093,N_12869,N_12768);
xor U13094 (N_13094,N_12864,N_12828);
xor U13095 (N_13095,N_12838,N_12766);
xnor U13096 (N_13096,N_12796,N_12870);
nand U13097 (N_13097,N_12990,N_12952);
nor U13098 (N_13098,N_12999,N_12963);
nand U13099 (N_13099,N_12855,N_12845);
nor U13100 (N_13100,N_12934,N_12771);
and U13101 (N_13101,N_12846,N_12752);
xnor U13102 (N_13102,N_12970,N_12866);
and U13103 (N_13103,N_12815,N_12826);
nor U13104 (N_13104,N_12962,N_12806);
and U13105 (N_13105,N_12830,N_12783);
xor U13106 (N_13106,N_12784,N_12932);
xor U13107 (N_13107,N_12823,N_12851);
xnor U13108 (N_13108,N_12778,N_12810);
or U13109 (N_13109,N_12946,N_12985);
or U13110 (N_13110,N_12978,N_12979);
nor U13111 (N_13111,N_12967,N_12904);
or U13112 (N_13112,N_12980,N_12801);
and U13113 (N_13113,N_12850,N_12840);
nor U13114 (N_13114,N_12899,N_12902);
and U13115 (N_13115,N_12812,N_12988);
xor U13116 (N_13116,N_12809,N_12777);
xor U13117 (N_13117,N_12841,N_12834);
xor U13118 (N_13118,N_12965,N_12911);
nand U13119 (N_13119,N_12972,N_12763);
xor U13120 (N_13120,N_12832,N_12814);
nand U13121 (N_13121,N_12966,N_12795);
and U13122 (N_13122,N_12901,N_12821);
nand U13123 (N_13123,N_12908,N_12893);
xor U13124 (N_13124,N_12918,N_12924);
nor U13125 (N_13125,N_12895,N_12845);
xnor U13126 (N_13126,N_12926,N_12897);
nand U13127 (N_13127,N_12942,N_12829);
nand U13128 (N_13128,N_12853,N_12881);
or U13129 (N_13129,N_12833,N_12791);
and U13130 (N_13130,N_12780,N_12978);
and U13131 (N_13131,N_12996,N_12895);
xnor U13132 (N_13132,N_12845,N_12964);
or U13133 (N_13133,N_12971,N_12904);
and U13134 (N_13134,N_12943,N_12972);
or U13135 (N_13135,N_12784,N_12775);
xnor U13136 (N_13136,N_12970,N_12762);
nor U13137 (N_13137,N_12914,N_12831);
nand U13138 (N_13138,N_12894,N_12902);
xor U13139 (N_13139,N_12873,N_12892);
and U13140 (N_13140,N_12839,N_12997);
nor U13141 (N_13141,N_12799,N_12978);
nand U13142 (N_13142,N_12998,N_12784);
or U13143 (N_13143,N_12782,N_12923);
nand U13144 (N_13144,N_12901,N_12813);
nor U13145 (N_13145,N_12942,N_12756);
nor U13146 (N_13146,N_12876,N_12950);
nor U13147 (N_13147,N_12887,N_12992);
xor U13148 (N_13148,N_12776,N_12878);
xor U13149 (N_13149,N_12769,N_12866);
or U13150 (N_13150,N_12751,N_12973);
or U13151 (N_13151,N_12970,N_12944);
xor U13152 (N_13152,N_12897,N_12963);
and U13153 (N_13153,N_12959,N_12897);
nand U13154 (N_13154,N_12765,N_12814);
or U13155 (N_13155,N_12919,N_12974);
or U13156 (N_13156,N_12861,N_12851);
nor U13157 (N_13157,N_12927,N_12966);
xor U13158 (N_13158,N_12932,N_12981);
or U13159 (N_13159,N_12996,N_12883);
and U13160 (N_13160,N_12856,N_12838);
nor U13161 (N_13161,N_12941,N_12830);
nor U13162 (N_13162,N_12802,N_12974);
xnor U13163 (N_13163,N_12819,N_12754);
or U13164 (N_13164,N_12925,N_12857);
nand U13165 (N_13165,N_12996,N_12872);
xor U13166 (N_13166,N_12791,N_12772);
and U13167 (N_13167,N_12777,N_12859);
nor U13168 (N_13168,N_12819,N_12897);
nor U13169 (N_13169,N_12828,N_12995);
and U13170 (N_13170,N_12763,N_12874);
nand U13171 (N_13171,N_12838,N_12942);
nor U13172 (N_13172,N_12852,N_12951);
nand U13173 (N_13173,N_12843,N_12754);
xnor U13174 (N_13174,N_12769,N_12903);
xor U13175 (N_13175,N_12882,N_12916);
nand U13176 (N_13176,N_12807,N_12759);
or U13177 (N_13177,N_12753,N_12868);
or U13178 (N_13178,N_12976,N_12995);
or U13179 (N_13179,N_12845,N_12954);
or U13180 (N_13180,N_12985,N_12856);
xor U13181 (N_13181,N_12994,N_12911);
xnor U13182 (N_13182,N_12881,N_12818);
and U13183 (N_13183,N_12911,N_12924);
nand U13184 (N_13184,N_12805,N_12864);
nor U13185 (N_13185,N_12795,N_12813);
nor U13186 (N_13186,N_12800,N_12871);
or U13187 (N_13187,N_12776,N_12913);
nand U13188 (N_13188,N_12979,N_12819);
and U13189 (N_13189,N_12799,N_12924);
and U13190 (N_13190,N_12991,N_12779);
nor U13191 (N_13191,N_12824,N_12831);
or U13192 (N_13192,N_12993,N_12859);
or U13193 (N_13193,N_12833,N_12977);
nand U13194 (N_13194,N_12791,N_12856);
nand U13195 (N_13195,N_12954,N_12767);
nor U13196 (N_13196,N_12786,N_12853);
nand U13197 (N_13197,N_12842,N_12824);
or U13198 (N_13198,N_12969,N_12861);
and U13199 (N_13199,N_12781,N_12986);
and U13200 (N_13200,N_12819,N_12856);
or U13201 (N_13201,N_12779,N_12785);
xnor U13202 (N_13202,N_12775,N_12875);
and U13203 (N_13203,N_12924,N_12773);
xnor U13204 (N_13204,N_12763,N_12976);
nor U13205 (N_13205,N_12862,N_12893);
xor U13206 (N_13206,N_12753,N_12930);
nor U13207 (N_13207,N_12966,N_12999);
or U13208 (N_13208,N_12965,N_12862);
and U13209 (N_13209,N_12934,N_12916);
nor U13210 (N_13210,N_12878,N_12824);
and U13211 (N_13211,N_12885,N_12855);
and U13212 (N_13212,N_12927,N_12991);
nor U13213 (N_13213,N_12895,N_12872);
nor U13214 (N_13214,N_12803,N_12815);
nor U13215 (N_13215,N_12754,N_12793);
and U13216 (N_13216,N_12850,N_12871);
nor U13217 (N_13217,N_12853,N_12910);
xor U13218 (N_13218,N_12938,N_12800);
and U13219 (N_13219,N_12995,N_12825);
or U13220 (N_13220,N_12834,N_12884);
nor U13221 (N_13221,N_12782,N_12965);
xnor U13222 (N_13222,N_12965,N_12934);
nand U13223 (N_13223,N_12950,N_12999);
or U13224 (N_13224,N_12986,N_12753);
or U13225 (N_13225,N_12813,N_12871);
or U13226 (N_13226,N_12913,N_12873);
or U13227 (N_13227,N_12908,N_12858);
nand U13228 (N_13228,N_12823,N_12898);
nor U13229 (N_13229,N_12857,N_12980);
nor U13230 (N_13230,N_12934,N_12822);
and U13231 (N_13231,N_12834,N_12981);
nor U13232 (N_13232,N_12934,N_12839);
nand U13233 (N_13233,N_12939,N_12952);
nand U13234 (N_13234,N_12866,N_12920);
or U13235 (N_13235,N_12950,N_12850);
nor U13236 (N_13236,N_12902,N_12896);
or U13237 (N_13237,N_12984,N_12847);
nor U13238 (N_13238,N_12939,N_12813);
nor U13239 (N_13239,N_12884,N_12985);
xor U13240 (N_13240,N_12982,N_12852);
nand U13241 (N_13241,N_12919,N_12910);
nand U13242 (N_13242,N_12988,N_12906);
or U13243 (N_13243,N_12883,N_12832);
and U13244 (N_13244,N_12887,N_12950);
or U13245 (N_13245,N_12871,N_12925);
and U13246 (N_13246,N_12870,N_12948);
nand U13247 (N_13247,N_12969,N_12991);
nor U13248 (N_13248,N_12843,N_12881);
nand U13249 (N_13249,N_12914,N_12948);
and U13250 (N_13250,N_13237,N_13068);
xor U13251 (N_13251,N_13135,N_13123);
nor U13252 (N_13252,N_13175,N_13097);
xnor U13253 (N_13253,N_13228,N_13002);
or U13254 (N_13254,N_13190,N_13227);
nor U13255 (N_13255,N_13127,N_13212);
xor U13256 (N_13256,N_13056,N_13049);
xor U13257 (N_13257,N_13025,N_13073);
nand U13258 (N_13258,N_13113,N_13075);
or U13259 (N_13259,N_13224,N_13236);
nor U13260 (N_13260,N_13194,N_13159);
and U13261 (N_13261,N_13089,N_13151);
or U13262 (N_13262,N_13196,N_13016);
xor U13263 (N_13263,N_13072,N_13100);
nor U13264 (N_13264,N_13112,N_13109);
or U13265 (N_13265,N_13206,N_13111);
nand U13266 (N_13266,N_13014,N_13182);
or U13267 (N_13267,N_13065,N_13091);
nand U13268 (N_13268,N_13116,N_13122);
and U13269 (N_13269,N_13012,N_13021);
xor U13270 (N_13270,N_13110,N_13219);
or U13271 (N_13271,N_13142,N_13061);
or U13272 (N_13272,N_13081,N_13235);
xor U13273 (N_13273,N_13031,N_13005);
or U13274 (N_13274,N_13169,N_13241);
xor U13275 (N_13275,N_13188,N_13119);
xor U13276 (N_13276,N_13043,N_13055);
nand U13277 (N_13277,N_13078,N_13167);
or U13278 (N_13278,N_13246,N_13150);
or U13279 (N_13279,N_13221,N_13059);
nand U13280 (N_13280,N_13071,N_13173);
xor U13281 (N_13281,N_13044,N_13028);
nand U13282 (N_13282,N_13018,N_13164);
and U13283 (N_13283,N_13132,N_13203);
nor U13284 (N_13284,N_13215,N_13128);
nor U13285 (N_13285,N_13160,N_13178);
nor U13286 (N_13286,N_13003,N_13226);
nand U13287 (N_13287,N_13153,N_13176);
and U13288 (N_13288,N_13172,N_13063);
nand U13289 (N_13289,N_13118,N_13138);
nand U13290 (N_13290,N_13171,N_13057);
xor U13291 (N_13291,N_13133,N_13248);
xnor U13292 (N_13292,N_13232,N_13201);
or U13293 (N_13293,N_13210,N_13168);
xor U13294 (N_13294,N_13101,N_13166);
or U13295 (N_13295,N_13230,N_13225);
or U13296 (N_13296,N_13129,N_13238);
nand U13297 (N_13297,N_13103,N_13036);
nor U13298 (N_13298,N_13008,N_13137);
xor U13299 (N_13299,N_13077,N_13050);
nor U13300 (N_13300,N_13195,N_13024);
nor U13301 (N_13301,N_13042,N_13156);
or U13302 (N_13302,N_13032,N_13147);
nor U13303 (N_13303,N_13192,N_13162);
nand U13304 (N_13304,N_13152,N_13035);
nand U13305 (N_13305,N_13247,N_13191);
nor U13306 (N_13306,N_13007,N_13045);
and U13307 (N_13307,N_13090,N_13180);
and U13308 (N_13308,N_13106,N_13058);
nand U13309 (N_13309,N_13023,N_13249);
or U13310 (N_13310,N_13177,N_13026);
xnor U13311 (N_13311,N_13205,N_13105);
nand U13312 (N_13312,N_13145,N_13202);
nor U13313 (N_13313,N_13189,N_13082);
nor U13314 (N_13314,N_13197,N_13011);
or U13315 (N_13315,N_13064,N_13170);
nand U13316 (N_13316,N_13074,N_13199);
or U13317 (N_13317,N_13141,N_13245);
and U13318 (N_13318,N_13051,N_13054);
nand U13319 (N_13319,N_13030,N_13087);
nor U13320 (N_13320,N_13001,N_13124);
nand U13321 (N_13321,N_13121,N_13213);
or U13322 (N_13322,N_13019,N_13200);
xnor U13323 (N_13323,N_13218,N_13174);
or U13324 (N_13324,N_13052,N_13066);
xor U13325 (N_13325,N_13130,N_13139);
nand U13326 (N_13326,N_13067,N_13234);
nand U13327 (N_13327,N_13204,N_13102);
or U13328 (N_13328,N_13086,N_13143);
xnor U13329 (N_13329,N_13069,N_13131);
nand U13330 (N_13330,N_13079,N_13239);
nor U13331 (N_13331,N_13107,N_13126);
or U13332 (N_13332,N_13181,N_13240);
nor U13333 (N_13333,N_13041,N_13125);
nand U13334 (N_13334,N_13038,N_13095);
or U13335 (N_13335,N_13193,N_13187);
xor U13336 (N_13336,N_13214,N_13163);
nor U13337 (N_13337,N_13149,N_13027);
xnor U13338 (N_13338,N_13062,N_13244);
nor U13339 (N_13339,N_13033,N_13155);
and U13340 (N_13340,N_13034,N_13093);
or U13341 (N_13341,N_13184,N_13220);
nand U13342 (N_13342,N_13208,N_13120);
nor U13343 (N_13343,N_13004,N_13243);
nand U13344 (N_13344,N_13104,N_13039);
nor U13345 (N_13345,N_13084,N_13136);
xnor U13346 (N_13346,N_13017,N_13006);
nor U13347 (N_13347,N_13165,N_13231);
or U13348 (N_13348,N_13134,N_13088);
nor U13349 (N_13349,N_13117,N_13216);
nand U13350 (N_13350,N_13185,N_13222);
and U13351 (N_13351,N_13048,N_13037);
xnor U13352 (N_13352,N_13096,N_13040);
xnor U13353 (N_13353,N_13053,N_13013);
and U13354 (N_13354,N_13211,N_13076);
and U13355 (N_13355,N_13094,N_13217);
and U13356 (N_13356,N_13207,N_13148);
nor U13357 (N_13357,N_13242,N_13198);
nand U13358 (N_13358,N_13209,N_13015);
nand U13359 (N_13359,N_13070,N_13154);
nor U13360 (N_13360,N_13083,N_13179);
nand U13361 (N_13361,N_13186,N_13020);
nand U13362 (N_13362,N_13140,N_13223);
xnor U13363 (N_13363,N_13092,N_13098);
or U13364 (N_13364,N_13085,N_13009);
and U13365 (N_13365,N_13046,N_13022);
or U13366 (N_13366,N_13047,N_13060);
nand U13367 (N_13367,N_13146,N_13144);
xnor U13368 (N_13368,N_13000,N_13183);
or U13369 (N_13369,N_13114,N_13115);
nor U13370 (N_13370,N_13080,N_13229);
or U13371 (N_13371,N_13108,N_13158);
and U13372 (N_13372,N_13161,N_13029);
nor U13373 (N_13373,N_13099,N_13233);
or U13374 (N_13374,N_13010,N_13157);
xnor U13375 (N_13375,N_13210,N_13141);
and U13376 (N_13376,N_13202,N_13028);
nand U13377 (N_13377,N_13159,N_13182);
or U13378 (N_13378,N_13067,N_13153);
nor U13379 (N_13379,N_13230,N_13087);
nor U13380 (N_13380,N_13181,N_13223);
nor U13381 (N_13381,N_13149,N_13050);
or U13382 (N_13382,N_13137,N_13088);
nor U13383 (N_13383,N_13100,N_13124);
and U13384 (N_13384,N_13070,N_13045);
or U13385 (N_13385,N_13157,N_13246);
and U13386 (N_13386,N_13062,N_13054);
xnor U13387 (N_13387,N_13182,N_13119);
and U13388 (N_13388,N_13065,N_13123);
xor U13389 (N_13389,N_13248,N_13132);
nor U13390 (N_13390,N_13235,N_13209);
and U13391 (N_13391,N_13110,N_13128);
nand U13392 (N_13392,N_13188,N_13120);
xnor U13393 (N_13393,N_13091,N_13070);
nand U13394 (N_13394,N_13131,N_13249);
nand U13395 (N_13395,N_13205,N_13125);
and U13396 (N_13396,N_13172,N_13088);
nor U13397 (N_13397,N_13065,N_13116);
or U13398 (N_13398,N_13180,N_13201);
and U13399 (N_13399,N_13011,N_13024);
or U13400 (N_13400,N_13221,N_13198);
and U13401 (N_13401,N_13066,N_13062);
and U13402 (N_13402,N_13088,N_13105);
nand U13403 (N_13403,N_13173,N_13103);
nor U13404 (N_13404,N_13074,N_13062);
xor U13405 (N_13405,N_13215,N_13141);
nor U13406 (N_13406,N_13139,N_13075);
nand U13407 (N_13407,N_13191,N_13119);
nand U13408 (N_13408,N_13088,N_13038);
nor U13409 (N_13409,N_13120,N_13147);
and U13410 (N_13410,N_13005,N_13079);
nor U13411 (N_13411,N_13172,N_13118);
and U13412 (N_13412,N_13220,N_13200);
and U13413 (N_13413,N_13187,N_13075);
and U13414 (N_13414,N_13054,N_13007);
nor U13415 (N_13415,N_13244,N_13133);
or U13416 (N_13416,N_13176,N_13235);
nor U13417 (N_13417,N_13102,N_13162);
or U13418 (N_13418,N_13200,N_13161);
and U13419 (N_13419,N_13236,N_13247);
or U13420 (N_13420,N_13094,N_13188);
and U13421 (N_13421,N_13236,N_13029);
or U13422 (N_13422,N_13071,N_13169);
nor U13423 (N_13423,N_13097,N_13148);
or U13424 (N_13424,N_13170,N_13074);
xor U13425 (N_13425,N_13220,N_13249);
xnor U13426 (N_13426,N_13241,N_13046);
nand U13427 (N_13427,N_13239,N_13226);
nor U13428 (N_13428,N_13181,N_13038);
xnor U13429 (N_13429,N_13105,N_13218);
nand U13430 (N_13430,N_13111,N_13204);
nor U13431 (N_13431,N_13177,N_13124);
and U13432 (N_13432,N_13029,N_13247);
nand U13433 (N_13433,N_13173,N_13131);
nand U13434 (N_13434,N_13125,N_13182);
nor U13435 (N_13435,N_13200,N_13238);
or U13436 (N_13436,N_13176,N_13079);
xor U13437 (N_13437,N_13235,N_13228);
and U13438 (N_13438,N_13023,N_13083);
nand U13439 (N_13439,N_13079,N_13204);
or U13440 (N_13440,N_13149,N_13165);
nor U13441 (N_13441,N_13079,N_13195);
nand U13442 (N_13442,N_13079,N_13081);
or U13443 (N_13443,N_13155,N_13131);
nor U13444 (N_13444,N_13236,N_13207);
nand U13445 (N_13445,N_13192,N_13064);
and U13446 (N_13446,N_13068,N_13072);
xnor U13447 (N_13447,N_13249,N_13033);
and U13448 (N_13448,N_13019,N_13240);
xnor U13449 (N_13449,N_13097,N_13113);
xor U13450 (N_13450,N_13065,N_13051);
nor U13451 (N_13451,N_13140,N_13128);
and U13452 (N_13452,N_13143,N_13159);
or U13453 (N_13453,N_13066,N_13152);
or U13454 (N_13454,N_13158,N_13244);
and U13455 (N_13455,N_13073,N_13082);
nand U13456 (N_13456,N_13065,N_13140);
or U13457 (N_13457,N_13095,N_13092);
and U13458 (N_13458,N_13219,N_13239);
or U13459 (N_13459,N_13057,N_13168);
nor U13460 (N_13460,N_13109,N_13005);
xnor U13461 (N_13461,N_13204,N_13231);
or U13462 (N_13462,N_13020,N_13132);
and U13463 (N_13463,N_13163,N_13017);
nor U13464 (N_13464,N_13073,N_13183);
xnor U13465 (N_13465,N_13115,N_13206);
xnor U13466 (N_13466,N_13055,N_13200);
nand U13467 (N_13467,N_13199,N_13109);
xnor U13468 (N_13468,N_13241,N_13029);
nand U13469 (N_13469,N_13235,N_13019);
or U13470 (N_13470,N_13150,N_13194);
and U13471 (N_13471,N_13025,N_13245);
or U13472 (N_13472,N_13240,N_13007);
nor U13473 (N_13473,N_13117,N_13238);
xnor U13474 (N_13474,N_13202,N_13248);
and U13475 (N_13475,N_13119,N_13080);
and U13476 (N_13476,N_13169,N_13124);
and U13477 (N_13477,N_13131,N_13063);
nor U13478 (N_13478,N_13007,N_13067);
nand U13479 (N_13479,N_13057,N_13133);
nand U13480 (N_13480,N_13221,N_13039);
or U13481 (N_13481,N_13159,N_13050);
nor U13482 (N_13482,N_13191,N_13100);
or U13483 (N_13483,N_13180,N_13134);
or U13484 (N_13484,N_13075,N_13045);
or U13485 (N_13485,N_13170,N_13113);
or U13486 (N_13486,N_13203,N_13051);
or U13487 (N_13487,N_13194,N_13126);
and U13488 (N_13488,N_13158,N_13216);
and U13489 (N_13489,N_13116,N_13024);
xnor U13490 (N_13490,N_13006,N_13023);
nand U13491 (N_13491,N_13101,N_13002);
nor U13492 (N_13492,N_13212,N_13039);
and U13493 (N_13493,N_13020,N_13220);
nand U13494 (N_13494,N_13139,N_13102);
xor U13495 (N_13495,N_13131,N_13001);
nor U13496 (N_13496,N_13236,N_13163);
or U13497 (N_13497,N_13086,N_13147);
nand U13498 (N_13498,N_13210,N_13230);
nor U13499 (N_13499,N_13010,N_13105);
nand U13500 (N_13500,N_13479,N_13330);
nand U13501 (N_13501,N_13304,N_13260);
or U13502 (N_13502,N_13427,N_13378);
nor U13503 (N_13503,N_13449,N_13490);
or U13504 (N_13504,N_13464,N_13388);
and U13505 (N_13505,N_13382,N_13476);
nor U13506 (N_13506,N_13424,N_13355);
xnor U13507 (N_13507,N_13328,N_13486);
or U13508 (N_13508,N_13422,N_13492);
nand U13509 (N_13509,N_13395,N_13253);
nand U13510 (N_13510,N_13359,N_13409);
nand U13511 (N_13511,N_13339,N_13438);
or U13512 (N_13512,N_13303,N_13307);
and U13513 (N_13513,N_13343,N_13284);
nand U13514 (N_13514,N_13285,N_13437);
xor U13515 (N_13515,N_13370,N_13419);
or U13516 (N_13516,N_13450,N_13394);
xor U13517 (N_13517,N_13410,N_13430);
nor U13518 (N_13518,N_13334,N_13400);
or U13519 (N_13519,N_13389,N_13418);
or U13520 (N_13520,N_13302,N_13365);
and U13521 (N_13521,N_13398,N_13273);
nor U13522 (N_13522,N_13270,N_13447);
xnor U13523 (N_13523,N_13368,N_13296);
xor U13524 (N_13524,N_13455,N_13458);
nand U13525 (N_13525,N_13351,N_13290);
nor U13526 (N_13526,N_13325,N_13357);
and U13527 (N_13527,N_13301,N_13429);
nor U13528 (N_13528,N_13411,N_13471);
nor U13529 (N_13529,N_13469,N_13448);
and U13530 (N_13530,N_13446,N_13277);
and U13531 (N_13531,N_13348,N_13250);
or U13532 (N_13532,N_13268,N_13261);
nor U13533 (N_13533,N_13435,N_13423);
and U13534 (N_13534,N_13344,N_13297);
xnor U13535 (N_13535,N_13392,N_13456);
xnor U13536 (N_13536,N_13279,N_13407);
nand U13537 (N_13537,N_13282,N_13298);
or U13538 (N_13538,N_13363,N_13477);
nor U13539 (N_13539,N_13482,N_13267);
or U13540 (N_13540,N_13300,N_13364);
or U13541 (N_13541,N_13292,N_13488);
or U13542 (N_13542,N_13366,N_13369);
nand U13543 (N_13543,N_13480,N_13416);
xnor U13544 (N_13544,N_13346,N_13428);
or U13545 (N_13545,N_13311,N_13467);
nor U13546 (N_13546,N_13322,N_13291);
xor U13547 (N_13547,N_13402,N_13465);
xor U13548 (N_13548,N_13276,N_13406);
or U13549 (N_13549,N_13256,N_13375);
nor U13550 (N_13550,N_13345,N_13452);
or U13551 (N_13551,N_13308,N_13367);
xor U13552 (N_13552,N_13404,N_13305);
or U13553 (N_13553,N_13352,N_13266);
nor U13554 (N_13554,N_13281,N_13376);
and U13555 (N_13555,N_13320,N_13444);
xnor U13556 (N_13556,N_13264,N_13373);
and U13557 (N_13557,N_13288,N_13272);
nor U13558 (N_13558,N_13439,N_13342);
nor U13559 (N_13559,N_13341,N_13251);
and U13560 (N_13560,N_13495,N_13472);
xnor U13561 (N_13561,N_13387,N_13318);
and U13562 (N_13562,N_13440,N_13417);
xor U13563 (N_13563,N_13385,N_13286);
xnor U13564 (N_13564,N_13313,N_13324);
and U13565 (N_13565,N_13489,N_13257);
or U13566 (N_13566,N_13425,N_13485);
and U13567 (N_13567,N_13280,N_13295);
or U13568 (N_13568,N_13453,N_13254);
xnor U13569 (N_13569,N_13274,N_13299);
nor U13570 (N_13570,N_13293,N_13316);
or U13571 (N_13571,N_13354,N_13294);
nand U13572 (N_13572,N_13319,N_13405);
xor U13573 (N_13573,N_13498,N_13326);
xnor U13574 (N_13574,N_13278,N_13321);
nor U13575 (N_13575,N_13413,N_13451);
nor U13576 (N_13576,N_13377,N_13432);
or U13577 (N_13577,N_13358,N_13384);
nor U13578 (N_13578,N_13493,N_13306);
xor U13579 (N_13579,N_13445,N_13317);
and U13580 (N_13580,N_13420,N_13252);
or U13581 (N_13581,N_13259,N_13323);
xor U13582 (N_13582,N_13460,N_13255);
xnor U13583 (N_13583,N_13466,N_13353);
nand U13584 (N_13584,N_13401,N_13399);
or U13585 (N_13585,N_13390,N_13258);
nand U13586 (N_13586,N_13478,N_13287);
and U13587 (N_13587,N_13309,N_13397);
or U13588 (N_13588,N_13473,N_13463);
and U13589 (N_13589,N_13391,N_13396);
and U13590 (N_13590,N_13421,N_13361);
or U13591 (N_13591,N_13338,N_13497);
nand U13592 (N_13592,N_13462,N_13356);
nor U13593 (N_13593,N_13380,N_13263);
xnor U13594 (N_13594,N_13374,N_13412);
nor U13595 (N_13595,N_13327,N_13362);
nor U13596 (N_13596,N_13426,N_13289);
nor U13597 (N_13597,N_13408,N_13350);
or U13598 (N_13598,N_13491,N_13265);
nand U13599 (N_13599,N_13349,N_13483);
or U13600 (N_13600,N_13271,N_13262);
or U13601 (N_13601,N_13494,N_13312);
or U13602 (N_13602,N_13433,N_13275);
nand U13603 (N_13603,N_13329,N_13347);
and U13604 (N_13604,N_13487,N_13371);
or U13605 (N_13605,N_13360,N_13496);
and U13606 (N_13606,N_13431,N_13442);
xor U13607 (N_13607,N_13372,N_13340);
and U13608 (N_13608,N_13403,N_13468);
nor U13609 (N_13609,N_13331,N_13335);
or U13610 (N_13610,N_13434,N_13475);
xor U13611 (N_13611,N_13283,N_13436);
nand U13612 (N_13612,N_13386,N_13470);
xor U13613 (N_13613,N_13337,N_13443);
or U13614 (N_13614,N_13454,N_13484);
nand U13615 (N_13615,N_13474,N_13499);
xnor U13616 (N_13616,N_13336,N_13459);
or U13617 (N_13617,N_13481,N_13333);
xor U13618 (N_13618,N_13310,N_13461);
or U13619 (N_13619,N_13269,N_13393);
nand U13620 (N_13620,N_13379,N_13332);
xnor U13621 (N_13621,N_13414,N_13315);
nand U13622 (N_13622,N_13381,N_13383);
nor U13623 (N_13623,N_13314,N_13457);
or U13624 (N_13624,N_13415,N_13441);
and U13625 (N_13625,N_13448,N_13374);
nand U13626 (N_13626,N_13424,N_13255);
or U13627 (N_13627,N_13295,N_13491);
or U13628 (N_13628,N_13330,N_13385);
and U13629 (N_13629,N_13490,N_13474);
and U13630 (N_13630,N_13296,N_13256);
nand U13631 (N_13631,N_13450,N_13376);
or U13632 (N_13632,N_13324,N_13494);
and U13633 (N_13633,N_13321,N_13399);
and U13634 (N_13634,N_13363,N_13324);
xnor U13635 (N_13635,N_13326,N_13383);
nand U13636 (N_13636,N_13426,N_13428);
nor U13637 (N_13637,N_13473,N_13332);
and U13638 (N_13638,N_13428,N_13482);
and U13639 (N_13639,N_13275,N_13355);
nor U13640 (N_13640,N_13307,N_13333);
nor U13641 (N_13641,N_13398,N_13454);
xor U13642 (N_13642,N_13481,N_13430);
or U13643 (N_13643,N_13421,N_13494);
or U13644 (N_13644,N_13255,N_13314);
and U13645 (N_13645,N_13280,N_13307);
nor U13646 (N_13646,N_13386,N_13422);
xnor U13647 (N_13647,N_13327,N_13349);
or U13648 (N_13648,N_13333,N_13495);
xor U13649 (N_13649,N_13371,N_13399);
nand U13650 (N_13650,N_13346,N_13426);
nor U13651 (N_13651,N_13408,N_13327);
and U13652 (N_13652,N_13415,N_13265);
nor U13653 (N_13653,N_13498,N_13304);
nand U13654 (N_13654,N_13482,N_13286);
and U13655 (N_13655,N_13472,N_13421);
or U13656 (N_13656,N_13466,N_13333);
nor U13657 (N_13657,N_13360,N_13330);
or U13658 (N_13658,N_13347,N_13388);
or U13659 (N_13659,N_13473,N_13355);
or U13660 (N_13660,N_13427,N_13282);
or U13661 (N_13661,N_13466,N_13352);
nor U13662 (N_13662,N_13393,N_13427);
and U13663 (N_13663,N_13424,N_13442);
xnor U13664 (N_13664,N_13490,N_13469);
nor U13665 (N_13665,N_13427,N_13355);
xor U13666 (N_13666,N_13486,N_13422);
nor U13667 (N_13667,N_13456,N_13335);
nor U13668 (N_13668,N_13252,N_13438);
xnor U13669 (N_13669,N_13451,N_13434);
or U13670 (N_13670,N_13458,N_13379);
and U13671 (N_13671,N_13465,N_13372);
nor U13672 (N_13672,N_13322,N_13361);
nand U13673 (N_13673,N_13277,N_13376);
nor U13674 (N_13674,N_13273,N_13368);
and U13675 (N_13675,N_13456,N_13372);
nor U13676 (N_13676,N_13251,N_13312);
or U13677 (N_13677,N_13473,N_13464);
xnor U13678 (N_13678,N_13473,N_13431);
nand U13679 (N_13679,N_13487,N_13268);
or U13680 (N_13680,N_13461,N_13429);
or U13681 (N_13681,N_13466,N_13497);
or U13682 (N_13682,N_13444,N_13262);
nor U13683 (N_13683,N_13332,N_13400);
and U13684 (N_13684,N_13453,N_13372);
nor U13685 (N_13685,N_13337,N_13338);
xor U13686 (N_13686,N_13303,N_13427);
and U13687 (N_13687,N_13398,N_13486);
xor U13688 (N_13688,N_13476,N_13415);
or U13689 (N_13689,N_13347,N_13353);
xor U13690 (N_13690,N_13431,N_13267);
or U13691 (N_13691,N_13333,N_13278);
nand U13692 (N_13692,N_13434,N_13459);
nor U13693 (N_13693,N_13459,N_13489);
and U13694 (N_13694,N_13298,N_13451);
nand U13695 (N_13695,N_13384,N_13285);
nor U13696 (N_13696,N_13403,N_13281);
xor U13697 (N_13697,N_13401,N_13426);
or U13698 (N_13698,N_13477,N_13301);
and U13699 (N_13699,N_13286,N_13389);
xor U13700 (N_13700,N_13343,N_13434);
nand U13701 (N_13701,N_13291,N_13250);
or U13702 (N_13702,N_13454,N_13466);
xnor U13703 (N_13703,N_13327,N_13366);
or U13704 (N_13704,N_13478,N_13446);
xor U13705 (N_13705,N_13411,N_13416);
and U13706 (N_13706,N_13381,N_13274);
or U13707 (N_13707,N_13484,N_13447);
nand U13708 (N_13708,N_13288,N_13373);
nor U13709 (N_13709,N_13286,N_13485);
or U13710 (N_13710,N_13307,N_13358);
xnor U13711 (N_13711,N_13361,N_13324);
or U13712 (N_13712,N_13441,N_13435);
and U13713 (N_13713,N_13395,N_13375);
or U13714 (N_13714,N_13331,N_13495);
and U13715 (N_13715,N_13321,N_13467);
and U13716 (N_13716,N_13381,N_13402);
and U13717 (N_13717,N_13489,N_13480);
nor U13718 (N_13718,N_13266,N_13297);
nand U13719 (N_13719,N_13312,N_13351);
or U13720 (N_13720,N_13492,N_13461);
nand U13721 (N_13721,N_13386,N_13356);
xnor U13722 (N_13722,N_13392,N_13273);
xnor U13723 (N_13723,N_13339,N_13437);
and U13724 (N_13724,N_13304,N_13394);
nor U13725 (N_13725,N_13335,N_13356);
or U13726 (N_13726,N_13440,N_13365);
or U13727 (N_13727,N_13391,N_13361);
or U13728 (N_13728,N_13268,N_13416);
and U13729 (N_13729,N_13288,N_13322);
or U13730 (N_13730,N_13281,N_13346);
and U13731 (N_13731,N_13447,N_13280);
xor U13732 (N_13732,N_13483,N_13448);
and U13733 (N_13733,N_13287,N_13322);
and U13734 (N_13734,N_13495,N_13490);
nor U13735 (N_13735,N_13379,N_13411);
xor U13736 (N_13736,N_13432,N_13415);
nand U13737 (N_13737,N_13309,N_13371);
nor U13738 (N_13738,N_13377,N_13304);
and U13739 (N_13739,N_13272,N_13251);
nor U13740 (N_13740,N_13351,N_13294);
or U13741 (N_13741,N_13446,N_13430);
nand U13742 (N_13742,N_13427,N_13394);
xnor U13743 (N_13743,N_13414,N_13314);
nand U13744 (N_13744,N_13490,N_13342);
and U13745 (N_13745,N_13304,N_13280);
and U13746 (N_13746,N_13466,N_13422);
and U13747 (N_13747,N_13286,N_13362);
and U13748 (N_13748,N_13304,N_13494);
and U13749 (N_13749,N_13256,N_13400);
or U13750 (N_13750,N_13571,N_13526);
nand U13751 (N_13751,N_13570,N_13589);
and U13752 (N_13752,N_13688,N_13670);
nor U13753 (N_13753,N_13523,N_13608);
and U13754 (N_13754,N_13647,N_13644);
xnor U13755 (N_13755,N_13576,N_13705);
or U13756 (N_13756,N_13702,N_13742);
xnor U13757 (N_13757,N_13538,N_13559);
or U13758 (N_13758,N_13569,N_13675);
and U13759 (N_13759,N_13633,N_13597);
and U13760 (N_13760,N_13619,N_13563);
xnor U13761 (N_13761,N_13717,N_13503);
or U13762 (N_13762,N_13522,N_13684);
xnor U13763 (N_13763,N_13550,N_13532);
or U13764 (N_13764,N_13720,N_13680);
and U13765 (N_13765,N_13690,N_13612);
and U13766 (N_13766,N_13507,N_13598);
and U13767 (N_13767,N_13554,N_13515);
nand U13768 (N_13768,N_13505,N_13689);
and U13769 (N_13769,N_13749,N_13723);
and U13770 (N_13770,N_13734,N_13708);
nor U13771 (N_13771,N_13737,N_13590);
or U13772 (N_13772,N_13635,N_13686);
nor U13773 (N_13773,N_13678,N_13582);
nand U13774 (N_13774,N_13724,N_13745);
and U13775 (N_13775,N_13714,N_13518);
or U13776 (N_13776,N_13676,N_13618);
nor U13777 (N_13777,N_13603,N_13606);
nand U13778 (N_13778,N_13551,N_13511);
or U13779 (N_13779,N_13533,N_13623);
or U13780 (N_13780,N_13525,N_13736);
and U13781 (N_13781,N_13561,N_13615);
nor U13782 (N_13782,N_13620,N_13501);
nand U13783 (N_13783,N_13659,N_13641);
xnor U13784 (N_13784,N_13663,N_13711);
or U13785 (N_13785,N_13510,N_13591);
xor U13786 (N_13786,N_13575,N_13669);
nor U13787 (N_13787,N_13642,N_13564);
or U13788 (N_13788,N_13624,N_13539);
and U13789 (N_13789,N_13548,N_13573);
and U13790 (N_13790,N_13691,N_13695);
nand U13791 (N_13791,N_13586,N_13668);
nor U13792 (N_13792,N_13656,N_13535);
xor U13793 (N_13793,N_13524,N_13580);
xor U13794 (N_13794,N_13739,N_13628);
or U13795 (N_13795,N_13517,N_13687);
nand U13796 (N_13796,N_13541,N_13562);
and U13797 (N_13797,N_13540,N_13648);
xnor U13798 (N_13798,N_13602,N_13611);
nand U13799 (N_13799,N_13701,N_13746);
xor U13800 (N_13800,N_13693,N_13643);
and U13801 (N_13801,N_13508,N_13662);
nor U13802 (N_13802,N_13747,N_13725);
and U13803 (N_13803,N_13528,N_13557);
nand U13804 (N_13804,N_13639,N_13629);
nand U13805 (N_13805,N_13574,N_13681);
and U13806 (N_13806,N_13732,N_13610);
and U13807 (N_13807,N_13596,N_13519);
xnor U13808 (N_13808,N_13592,N_13645);
nand U13809 (N_13809,N_13558,N_13545);
or U13810 (N_13810,N_13672,N_13500);
nor U13811 (N_13811,N_13738,N_13630);
nand U13812 (N_13812,N_13584,N_13527);
xnor U13813 (N_13813,N_13706,N_13555);
xor U13814 (N_13814,N_13609,N_13567);
nand U13815 (N_13815,N_13731,N_13604);
xor U13816 (N_13816,N_13617,N_13651);
nor U13817 (N_13817,N_13722,N_13613);
xor U13818 (N_13818,N_13700,N_13650);
or U13819 (N_13819,N_13568,N_13729);
nand U13820 (N_13820,N_13553,N_13677);
xnor U13821 (N_13821,N_13679,N_13735);
nand U13822 (N_13822,N_13572,N_13683);
nor U13823 (N_13823,N_13682,N_13657);
nor U13824 (N_13824,N_13716,N_13653);
nor U13825 (N_13825,N_13621,N_13649);
nand U13826 (N_13826,N_13529,N_13709);
and U13827 (N_13827,N_13730,N_13614);
nand U13828 (N_13828,N_13660,N_13585);
or U13829 (N_13829,N_13704,N_13546);
or U13830 (N_13830,N_13599,N_13566);
xor U13831 (N_13831,N_13626,N_13685);
nor U13832 (N_13832,N_13697,N_13552);
nor U13833 (N_13833,N_13696,N_13646);
nor U13834 (N_13834,N_13531,N_13547);
or U13835 (N_13835,N_13616,N_13521);
xnor U13836 (N_13836,N_13640,N_13520);
nor U13837 (N_13837,N_13587,N_13631);
nor U13838 (N_13838,N_13632,N_13713);
or U13839 (N_13839,N_13560,N_13694);
xor U13840 (N_13840,N_13605,N_13530);
and U13841 (N_13841,N_13671,N_13652);
nand U13842 (N_13842,N_13719,N_13542);
and U13843 (N_13843,N_13654,N_13544);
or U13844 (N_13844,N_13655,N_13740);
nand U13845 (N_13845,N_13673,N_13504);
nor U13846 (N_13846,N_13502,N_13658);
and U13847 (N_13847,N_13726,N_13579);
xnor U13848 (N_13848,N_13664,N_13625);
nor U13849 (N_13849,N_13595,N_13534);
xnor U13850 (N_13850,N_13607,N_13667);
and U13851 (N_13851,N_13594,N_13715);
or U13852 (N_13852,N_13537,N_13748);
xnor U13853 (N_13853,N_13512,N_13588);
or U13854 (N_13854,N_13578,N_13637);
or U13855 (N_13855,N_13593,N_13622);
or U13856 (N_13856,N_13733,N_13638);
xor U13857 (N_13857,N_13703,N_13727);
nor U13858 (N_13858,N_13661,N_13674);
nand U13859 (N_13859,N_13513,N_13516);
and U13860 (N_13860,N_13665,N_13581);
nor U13861 (N_13861,N_13556,N_13634);
nand U13862 (N_13862,N_13543,N_13601);
and U13863 (N_13863,N_13721,N_13536);
or U13864 (N_13864,N_13707,N_13509);
and U13865 (N_13865,N_13666,N_13514);
and U13866 (N_13866,N_13583,N_13577);
xnor U13867 (N_13867,N_13627,N_13710);
xor U13868 (N_13868,N_13712,N_13718);
or U13869 (N_13869,N_13565,N_13741);
nand U13870 (N_13870,N_13692,N_13636);
or U13871 (N_13871,N_13549,N_13699);
and U13872 (N_13872,N_13600,N_13728);
nor U13873 (N_13873,N_13506,N_13744);
and U13874 (N_13874,N_13743,N_13698);
or U13875 (N_13875,N_13528,N_13656);
nand U13876 (N_13876,N_13557,N_13738);
xnor U13877 (N_13877,N_13524,N_13629);
or U13878 (N_13878,N_13504,N_13611);
or U13879 (N_13879,N_13613,N_13522);
nor U13880 (N_13880,N_13635,N_13513);
or U13881 (N_13881,N_13717,N_13685);
nor U13882 (N_13882,N_13714,N_13680);
or U13883 (N_13883,N_13564,N_13568);
nor U13884 (N_13884,N_13733,N_13644);
and U13885 (N_13885,N_13636,N_13606);
and U13886 (N_13886,N_13547,N_13741);
nand U13887 (N_13887,N_13504,N_13704);
nor U13888 (N_13888,N_13623,N_13550);
xnor U13889 (N_13889,N_13572,N_13614);
and U13890 (N_13890,N_13568,N_13508);
xor U13891 (N_13891,N_13608,N_13634);
nand U13892 (N_13892,N_13575,N_13582);
nand U13893 (N_13893,N_13685,N_13536);
nand U13894 (N_13894,N_13564,N_13511);
or U13895 (N_13895,N_13587,N_13642);
and U13896 (N_13896,N_13568,N_13704);
nor U13897 (N_13897,N_13647,N_13631);
or U13898 (N_13898,N_13549,N_13520);
or U13899 (N_13899,N_13586,N_13729);
or U13900 (N_13900,N_13565,N_13685);
or U13901 (N_13901,N_13672,N_13576);
nor U13902 (N_13902,N_13589,N_13675);
xnor U13903 (N_13903,N_13545,N_13597);
nand U13904 (N_13904,N_13520,N_13560);
nor U13905 (N_13905,N_13646,N_13734);
or U13906 (N_13906,N_13511,N_13640);
and U13907 (N_13907,N_13580,N_13629);
nand U13908 (N_13908,N_13527,N_13616);
nand U13909 (N_13909,N_13637,N_13616);
and U13910 (N_13910,N_13689,N_13712);
and U13911 (N_13911,N_13635,N_13502);
and U13912 (N_13912,N_13724,N_13669);
nand U13913 (N_13913,N_13501,N_13685);
or U13914 (N_13914,N_13540,N_13670);
and U13915 (N_13915,N_13528,N_13507);
or U13916 (N_13916,N_13541,N_13710);
xor U13917 (N_13917,N_13692,N_13627);
xor U13918 (N_13918,N_13500,N_13539);
and U13919 (N_13919,N_13632,N_13529);
nand U13920 (N_13920,N_13684,N_13713);
nor U13921 (N_13921,N_13549,N_13727);
nand U13922 (N_13922,N_13507,N_13748);
and U13923 (N_13923,N_13689,N_13541);
nor U13924 (N_13924,N_13688,N_13587);
and U13925 (N_13925,N_13539,N_13555);
xor U13926 (N_13926,N_13614,N_13745);
xnor U13927 (N_13927,N_13619,N_13546);
nand U13928 (N_13928,N_13701,N_13622);
nand U13929 (N_13929,N_13712,N_13558);
nor U13930 (N_13930,N_13709,N_13565);
nor U13931 (N_13931,N_13575,N_13611);
nor U13932 (N_13932,N_13506,N_13712);
or U13933 (N_13933,N_13524,N_13743);
or U13934 (N_13934,N_13500,N_13741);
and U13935 (N_13935,N_13661,N_13742);
nor U13936 (N_13936,N_13575,N_13672);
nor U13937 (N_13937,N_13506,N_13588);
nand U13938 (N_13938,N_13633,N_13603);
xor U13939 (N_13939,N_13582,N_13518);
nor U13940 (N_13940,N_13721,N_13516);
nor U13941 (N_13941,N_13503,N_13579);
and U13942 (N_13942,N_13648,N_13610);
or U13943 (N_13943,N_13620,N_13622);
or U13944 (N_13944,N_13548,N_13555);
nor U13945 (N_13945,N_13512,N_13558);
nand U13946 (N_13946,N_13668,N_13706);
xnor U13947 (N_13947,N_13552,N_13680);
and U13948 (N_13948,N_13633,N_13573);
nand U13949 (N_13949,N_13746,N_13523);
nand U13950 (N_13950,N_13687,N_13545);
or U13951 (N_13951,N_13500,N_13615);
xor U13952 (N_13952,N_13733,N_13728);
or U13953 (N_13953,N_13626,N_13551);
xor U13954 (N_13954,N_13726,N_13685);
and U13955 (N_13955,N_13742,N_13561);
or U13956 (N_13956,N_13655,N_13656);
nor U13957 (N_13957,N_13679,N_13534);
or U13958 (N_13958,N_13649,N_13673);
or U13959 (N_13959,N_13638,N_13501);
xnor U13960 (N_13960,N_13604,N_13602);
or U13961 (N_13961,N_13595,N_13654);
or U13962 (N_13962,N_13516,N_13565);
nor U13963 (N_13963,N_13561,N_13587);
xor U13964 (N_13964,N_13525,N_13684);
or U13965 (N_13965,N_13627,N_13643);
nor U13966 (N_13966,N_13585,N_13732);
nand U13967 (N_13967,N_13639,N_13593);
and U13968 (N_13968,N_13609,N_13501);
nor U13969 (N_13969,N_13592,N_13738);
and U13970 (N_13970,N_13505,N_13643);
nor U13971 (N_13971,N_13612,N_13596);
xnor U13972 (N_13972,N_13596,N_13706);
and U13973 (N_13973,N_13516,N_13690);
and U13974 (N_13974,N_13667,N_13745);
xor U13975 (N_13975,N_13506,N_13675);
or U13976 (N_13976,N_13626,N_13566);
or U13977 (N_13977,N_13508,N_13567);
nor U13978 (N_13978,N_13668,N_13572);
and U13979 (N_13979,N_13659,N_13587);
and U13980 (N_13980,N_13577,N_13575);
xnor U13981 (N_13981,N_13567,N_13672);
xnor U13982 (N_13982,N_13569,N_13546);
nor U13983 (N_13983,N_13561,N_13553);
nand U13984 (N_13984,N_13711,N_13734);
nor U13985 (N_13985,N_13532,N_13739);
nand U13986 (N_13986,N_13618,N_13729);
or U13987 (N_13987,N_13711,N_13657);
and U13988 (N_13988,N_13566,N_13586);
or U13989 (N_13989,N_13579,N_13661);
nor U13990 (N_13990,N_13646,N_13578);
nand U13991 (N_13991,N_13536,N_13731);
nor U13992 (N_13992,N_13672,N_13735);
nand U13993 (N_13993,N_13622,N_13557);
nand U13994 (N_13994,N_13521,N_13654);
nand U13995 (N_13995,N_13710,N_13575);
nor U13996 (N_13996,N_13592,N_13648);
and U13997 (N_13997,N_13559,N_13604);
nor U13998 (N_13998,N_13730,N_13718);
or U13999 (N_13999,N_13569,N_13596);
xnor U14000 (N_14000,N_13982,N_13968);
and U14001 (N_14001,N_13759,N_13866);
nand U14002 (N_14002,N_13953,N_13904);
nand U14003 (N_14003,N_13776,N_13889);
xnor U14004 (N_14004,N_13951,N_13954);
nor U14005 (N_14005,N_13811,N_13870);
and U14006 (N_14006,N_13808,N_13823);
xnor U14007 (N_14007,N_13906,N_13958);
or U14008 (N_14008,N_13883,N_13816);
or U14009 (N_14009,N_13960,N_13765);
and U14010 (N_14010,N_13832,N_13859);
nor U14011 (N_14011,N_13821,N_13941);
xnor U14012 (N_14012,N_13983,N_13852);
and U14013 (N_14013,N_13931,N_13989);
and U14014 (N_14014,N_13986,N_13772);
and U14015 (N_14015,N_13908,N_13767);
or U14016 (N_14016,N_13981,N_13944);
nor U14017 (N_14017,N_13936,N_13812);
or U14018 (N_14018,N_13771,N_13871);
nand U14019 (N_14019,N_13798,N_13780);
and U14020 (N_14020,N_13804,N_13949);
nand U14021 (N_14021,N_13775,N_13948);
xor U14022 (N_14022,N_13881,N_13894);
xnor U14023 (N_14023,N_13916,N_13827);
xnor U14024 (N_14024,N_13991,N_13988);
or U14025 (N_14025,N_13930,N_13836);
and U14026 (N_14026,N_13878,N_13886);
nor U14027 (N_14027,N_13888,N_13807);
nor U14028 (N_14028,N_13751,N_13994);
nand U14029 (N_14029,N_13873,N_13795);
nor U14030 (N_14030,N_13861,N_13839);
nand U14031 (N_14031,N_13955,N_13834);
nand U14032 (N_14032,N_13814,N_13865);
and U14033 (N_14033,N_13992,N_13845);
or U14034 (N_14034,N_13914,N_13770);
nor U14035 (N_14035,N_13758,N_13867);
or U14036 (N_14036,N_13862,N_13921);
and U14037 (N_14037,N_13756,N_13782);
or U14038 (N_14038,N_13830,N_13912);
or U14039 (N_14039,N_13973,N_13840);
and U14040 (N_14040,N_13915,N_13764);
nand U14041 (N_14041,N_13882,N_13841);
nand U14042 (N_14042,N_13942,N_13920);
nor U14043 (N_14043,N_13879,N_13843);
nand U14044 (N_14044,N_13938,N_13909);
nor U14045 (N_14045,N_13802,N_13791);
nor U14046 (N_14046,N_13806,N_13831);
nand U14047 (N_14047,N_13974,N_13987);
nor U14048 (N_14048,N_13817,N_13937);
xnor U14049 (N_14049,N_13926,N_13887);
nor U14050 (N_14050,N_13940,N_13774);
nor U14051 (N_14051,N_13947,N_13863);
nor U14052 (N_14052,N_13826,N_13796);
or U14053 (N_14053,N_13825,N_13950);
xnor U14054 (N_14054,N_13956,N_13829);
nor U14055 (N_14055,N_13857,N_13877);
or U14056 (N_14056,N_13868,N_13922);
xnor U14057 (N_14057,N_13820,N_13833);
nor U14058 (N_14058,N_13925,N_13900);
or U14059 (N_14059,N_13896,N_13966);
xor U14060 (N_14060,N_13792,N_13847);
nand U14061 (N_14061,N_13917,N_13971);
nand U14062 (N_14062,N_13943,N_13952);
or U14063 (N_14063,N_13869,N_13837);
xor U14064 (N_14064,N_13998,N_13903);
nor U14065 (N_14065,N_13809,N_13924);
or U14066 (N_14066,N_13768,N_13898);
and U14067 (N_14067,N_13783,N_13850);
nand U14068 (N_14068,N_13893,N_13805);
nand U14069 (N_14069,N_13990,N_13786);
nor U14070 (N_14070,N_13853,N_13860);
and U14071 (N_14071,N_13975,N_13838);
or U14072 (N_14072,N_13962,N_13901);
and U14073 (N_14073,N_13763,N_13874);
and U14074 (N_14074,N_13781,N_13890);
xor U14075 (N_14075,N_13970,N_13815);
or U14076 (N_14076,N_13977,N_13935);
and U14077 (N_14077,N_13891,N_13846);
xor U14078 (N_14078,N_13761,N_13785);
xnor U14079 (N_14079,N_13919,N_13779);
nor U14080 (N_14080,N_13872,N_13910);
or U14081 (N_14081,N_13828,N_13911);
nand U14082 (N_14082,N_13803,N_13799);
nand U14083 (N_14083,N_13801,N_13884);
nand U14084 (N_14084,N_13961,N_13895);
nor U14085 (N_14085,N_13876,N_13789);
nor U14086 (N_14086,N_13972,N_13939);
nor U14087 (N_14087,N_13965,N_13993);
or U14088 (N_14088,N_13760,N_13923);
xor U14089 (N_14089,N_13848,N_13849);
xnor U14090 (N_14090,N_13907,N_13750);
and U14091 (N_14091,N_13856,N_13819);
or U14092 (N_14092,N_13754,N_13788);
xnor U14093 (N_14093,N_13946,N_13755);
nor U14094 (N_14094,N_13818,N_13855);
nor U14095 (N_14095,N_13793,N_13842);
and U14096 (N_14096,N_13757,N_13899);
nand U14097 (N_14097,N_13995,N_13753);
nor U14098 (N_14098,N_13854,N_13999);
nand U14099 (N_14099,N_13957,N_13766);
xnor U14100 (N_14100,N_13813,N_13835);
xnor U14101 (N_14101,N_13797,N_13969);
and U14102 (N_14102,N_13997,N_13976);
and U14103 (N_14103,N_13929,N_13794);
nand U14104 (N_14104,N_13985,N_13963);
nand U14105 (N_14105,N_13918,N_13800);
xnor U14106 (N_14106,N_13934,N_13787);
nand U14107 (N_14107,N_13880,N_13932);
and U14108 (N_14108,N_13790,N_13913);
nor U14109 (N_14109,N_13824,N_13967);
xor U14110 (N_14110,N_13844,N_13752);
or U14111 (N_14111,N_13773,N_13858);
nand U14112 (N_14112,N_13945,N_13875);
nor U14113 (N_14113,N_13933,N_13777);
or U14114 (N_14114,N_13964,N_13851);
or U14115 (N_14115,N_13959,N_13928);
nor U14116 (N_14116,N_13892,N_13978);
xor U14117 (N_14117,N_13784,N_13927);
or U14118 (N_14118,N_13885,N_13810);
xor U14119 (N_14119,N_13902,N_13905);
and U14120 (N_14120,N_13984,N_13769);
and U14121 (N_14121,N_13979,N_13897);
or U14122 (N_14122,N_13762,N_13778);
nor U14123 (N_14123,N_13996,N_13864);
or U14124 (N_14124,N_13822,N_13980);
or U14125 (N_14125,N_13916,N_13813);
xnor U14126 (N_14126,N_13836,N_13775);
nor U14127 (N_14127,N_13933,N_13925);
nor U14128 (N_14128,N_13799,N_13863);
nor U14129 (N_14129,N_13829,N_13933);
xnor U14130 (N_14130,N_13898,N_13971);
xnor U14131 (N_14131,N_13880,N_13876);
and U14132 (N_14132,N_13821,N_13750);
nand U14133 (N_14133,N_13912,N_13757);
xnor U14134 (N_14134,N_13944,N_13821);
xor U14135 (N_14135,N_13825,N_13770);
and U14136 (N_14136,N_13801,N_13798);
nand U14137 (N_14137,N_13881,N_13876);
nand U14138 (N_14138,N_13797,N_13917);
and U14139 (N_14139,N_13923,N_13870);
nor U14140 (N_14140,N_13958,N_13909);
nor U14141 (N_14141,N_13920,N_13778);
xor U14142 (N_14142,N_13889,N_13769);
xor U14143 (N_14143,N_13831,N_13868);
nand U14144 (N_14144,N_13953,N_13960);
nor U14145 (N_14145,N_13992,N_13925);
and U14146 (N_14146,N_13990,N_13780);
nor U14147 (N_14147,N_13760,N_13861);
or U14148 (N_14148,N_13761,N_13929);
nor U14149 (N_14149,N_13812,N_13998);
or U14150 (N_14150,N_13756,N_13811);
nand U14151 (N_14151,N_13939,N_13850);
nor U14152 (N_14152,N_13998,N_13981);
nor U14153 (N_14153,N_13839,N_13790);
nand U14154 (N_14154,N_13903,N_13965);
nand U14155 (N_14155,N_13765,N_13927);
or U14156 (N_14156,N_13902,N_13878);
nor U14157 (N_14157,N_13848,N_13924);
or U14158 (N_14158,N_13814,N_13893);
or U14159 (N_14159,N_13909,N_13850);
and U14160 (N_14160,N_13793,N_13766);
or U14161 (N_14161,N_13844,N_13762);
nand U14162 (N_14162,N_13991,N_13822);
xor U14163 (N_14163,N_13785,N_13981);
nor U14164 (N_14164,N_13937,N_13954);
nand U14165 (N_14165,N_13825,N_13865);
or U14166 (N_14166,N_13945,N_13853);
and U14167 (N_14167,N_13857,N_13828);
nand U14168 (N_14168,N_13798,N_13811);
and U14169 (N_14169,N_13836,N_13851);
nand U14170 (N_14170,N_13959,N_13782);
nand U14171 (N_14171,N_13853,N_13896);
or U14172 (N_14172,N_13875,N_13817);
and U14173 (N_14173,N_13961,N_13868);
nand U14174 (N_14174,N_13864,N_13990);
xor U14175 (N_14175,N_13766,N_13758);
and U14176 (N_14176,N_13759,N_13814);
nor U14177 (N_14177,N_13925,N_13881);
or U14178 (N_14178,N_13906,N_13767);
and U14179 (N_14179,N_13986,N_13894);
nand U14180 (N_14180,N_13852,N_13878);
or U14181 (N_14181,N_13827,N_13813);
or U14182 (N_14182,N_13953,N_13921);
nand U14183 (N_14183,N_13781,N_13897);
xor U14184 (N_14184,N_13945,N_13795);
nor U14185 (N_14185,N_13768,N_13852);
and U14186 (N_14186,N_13885,N_13952);
nand U14187 (N_14187,N_13930,N_13863);
nor U14188 (N_14188,N_13777,N_13952);
or U14189 (N_14189,N_13910,N_13835);
and U14190 (N_14190,N_13990,N_13836);
and U14191 (N_14191,N_13750,N_13849);
or U14192 (N_14192,N_13917,N_13958);
nor U14193 (N_14193,N_13957,N_13792);
nand U14194 (N_14194,N_13842,N_13780);
nor U14195 (N_14195,N_13955,N_13976);
nor U14196 (N_14196,N_13946,N_13778);
xnor U14197 (N_14197,N_13850,N_13864);
and U14198 (N_14198,N_13814,N_13855);
nor U14199 (N_14199,N_13822,N_13886);
xor U14200 (N_14200,N_13894,N_13891);
nor U14201 (N_14201,N_13758,N_13831);
nand U14202 (N_14202,N_13903,N_13762);
xor U14203 (N_14203,N_13949,N_13899);
nor U14204 (N_14204,N_13988,N_13857);
and U14205 (N_14205,N_13855,N_13951);
nand U14206 (N_14206,N_13982,N_13880);
and U14207 (N_14207,N_13851,N_13951);
and U14208 (N_14208,N_13968,N_13907);
or U14209 (N_14209,N_13880,N_13959);
nand U14210 (N_14210,N_13919,N_13904);
or U14211 (N_14211,N_13856,N_13842);
and U14212 (N_14212,N_13865,N_13853);
and U14213 (N_14213,N_13949,N_13806);
and U14214 (N_14214,N_13951,N_13828);
nor U14215 (N_14215,N_13787,N_13935);
xnor U14216 (N_14216,N_13819,N_13990);
nor U14217 (N_14217,N_13842,N_13992);
xor U14218 (N_14218,N_13906,N_13820);
xor U14219 (N_14219,N_13821,N_13950);
and U14220 (N_14220,N_13752,N_13758);
or U14221 (N_14221,N_13887,N_13784);
and U14222 (N_14222,N_13893,N_13979);
or U14223 (N_14223,N_13851,N_13823);
nor U14224 (N_14224,N_13839,N_13876);
nand U14225 (N_14225,N_13904,N_13782);
xnor U14226 (N_14226,N_13961,N_13970);
xor U14227 (N_14227,N_13755,N_13922);
nand U14228 (N_14228,N_13751,N_13910);
or U14229 (N_14229,N_13775,N_13893);
or U14230 (N_14230,N_13781,N_13917);
and U14231 (N_14231,N_13787,N_13866);
xnor U14232 (N_14232,N_13751,N_13963);
xor U14233 (N_14233,N_13946,N_13980);
nor U14234 (N_14234,N_13871,N_13792);
or U14235 (N_14235,N_13760,N_13860);
and U14236 (N_14236,N_13771,N_13973);
nor U14237 (N_14237,N_13925,N_13822);
nand U14238 (N_14238,N_13879,N_13789);
and U14239 (N_14239,N_13906,N_13932);
xnor U14240 (N_14240,N_13908,N_13850);
nand U14241 (N_14241,N_13826,N_13827);
xnor U14242 (N_14242,N_13942,N_13872);
or U14243 (N_14243,N_13906,N_13967);
nand U14244 (N_14244,N_13950,N_13752);
nand U14245 (N_14245,N_13965,N_13990);
and U14246 (N_14246,N_13956,N_13831);
nand U14247 (N_14247,N_13993,N_13914);
nor U14248 (N_14248,N_13924,N_13882);
or U14249 (N_14249,N_13895,N_13920);
or U14250 (N_14250,N_14009,N_14220);
or U14251 (N_14251,N_14125,N_14053);
and U14252 (N_14252,N_14033,N_14095);
or U14253 (N_14253,N_14234,N_14204);
nor U14254 (N_14254,N_14217,N_14044);
and U14255 (N_14255,N_14114,N_14133);
nor U14256 (N_14256,N_14112,N_14213);
or U14257 (N_14257,N_14101,N_14134);
and U14258 (N_14258,N_14149,N_14207);
nand U14259 (N_14259,N_14158,N_14135);
or U14260 (N_14260,N_14100,N_14071);
xor U14261 (N_14261,N_14006,N_14208);
nand U14262 (N_14262,N_14064,N_14067);
and U14263 (N_14263,N_14073,N_14247);
or U14264 (N_14264,N_14153,N_14235);
nor U14265 (N_14265,N_14242,N_14025);
xnor U14266 (N_14266,N_14188,N_14192);
nor U14267 (N_14267,N_14178,N_14078);
nor U14268 (N_14268,N_14055,N_14086);
and U14269 (N_14269,N_14040,N_14048);
xnor U14270 (N_14270,N_14168,N_14090);
and U14271 (N_14271,N_14120,N_14194);
or U14272 (N_14272,N_14110,N_14173);
and U14273 (N_14273,N_14218,N_14015);
nor U14274 (N_14274,N_14179,N_14076);
nor U14275 (N_14275,N_14057,N_14170);
and U14276 (N_14276,N_14130,N_14074);
nor U14277 (N_14277,N_14108,N_14243);
or U14278 (N_14278,N_14079,N_14199);
and U14279 (N_14279,N_14165,N_14138);
or U14280 (N_14280,N_14052,N_14177);
or U14281 (N_14281,N_14042,N_14087);
or U14282 (N_14282,N_14065,N_14206);
xor U14283 (N_14283,N_14231,N_14066);
xor U14284 (N_14284,N_14222,N_14148);
xor U14285 (N_14285,N_14146,N_14157);
nand U14286 (N_14286,N_14131,N_14142);
xnor U14287 (N_14287,N_14171,N_14163);
and U14288 (N_14288,N_14010,N_14062);
or U14289 (N_14289,N_14027,N_14096);
or U14290 (N_14290,N_14151,N_14164);
nand U14291 (N_14291,N_14059,N_14167);
nor U14292 (N_14292,N_14002,N_14223);
nor U14293 (N_14293,N_14014,N_14003);
nor U14294 (N_14294,N_14129,N_14012);
xnor U14295 (N_14295,N_14038,N_14032);
nor U14296 (N_14296,N_14099,N_14020);
or U14297 (N_14297,N_14245,N_14195);
nand U14298 (N_14298,N_14037,N_14080);
xnor U14299 (N_14299,N_14184,N_14019);
nor U14300 (N_14300,N_14126,N_14160);
xnor U14301 (N_14301,N_14034,N_14183);
or U14302 (N_14302,N_14116,N_14068);
xor U14303 (N_14303,N_14205,N_14132);
and U14304 (N_14304,N_14072,N_14169);
and U14305 (N_14305,N_14091,N_14202);
and U14306 (N_14306,N_14050,N_14175);
nand U14307 (N_14307,N_14196,N_14000);
or U14308 (N_14308,N_14239,N_14182);
xnor U14309 (N_14309,N_14144,N_14008);
and U14310 (N_14310,N_14180,N_14140);
and U14311 (N_14311,N_14161,N_14081);
or U14312 (N_14312,N_14249,N_14215);
or U14313 (N_14313,N_14021,N_14122);
and U14314 (N_14314,N_14233,N_14045);
nand U14315 (N_14315,N_14113,N_14229);
nand U14316 (N_14316,N_14221,N_14145);
nand U14317 (N_14317,N_14123,N_14022);
and U14318 (N_14318,N_14190,N_14241);
nand U14319 (N_14319,N_14075,N_14107);
or U14320 (N_14320,N_14041,N_14185);
xor U14321 (N_14321,N_14069,N_14085);
nor U14322 (N_14322,N_14056,N_14186);
or U14323 (N_14323,N_14106,N_14198);
nor U14324 (N_14324,N_14124,N_14121);
xnor U14325 (N_14325,N_14216,N_14211);
nor U14326 (N_14326,N_14007,N_14093);
xor U14327 (N_14327,N_14102,N_14028);
nand U14328 (N_14328,N_14083,N_14077);
nor U14329 (N_14329,N_14097,N_14230);
nand U14330 (N_14330,N_14043,N_14237);
or U14331 (N_14331,N_14029,N_14004);
and U14332 (N_14332,N_14094,N_14147);
nor U14333 (N_14333,N_14226,N_14200);
or U14334 (N_14334,N_14212,N_14162);
and U14335 (N_14335,N_14089,N_14219);
and U14336 (N_14336,N_14156,N_14154);
nand U14337 (N_14337,N_14039,N_14141);
nand U14338 (N_14338,N_14011,N_14103);
nand U14339 (N_14339,N_14115,N_14201);
and U14340 (N_14340,N_14139,N_14070);
or U14341 (N_14341,N_14127,N_14238);
or U14342 (N_14342,N_14018,N_14118);
nand U14343 (N_14343,N_14236,N_14001);
xnor U14344 (N_14344,N_14244,N_14152);
and U14345 (N_14345,N_14036,N_14054);
and U14346 (N_14346,N_14017,N_14031);
and U14347 (N_14347,N_14143,N_14246);
nand U14348 (N_14348,N_14203,N_14117);
xor U14349 (N_14349,N_14026,N_14193);
or U14350 (N_14350,N_14084,N_14248);
and U14351 (N_14351,N_14105,N_14024);
nand U14352 (N_14352,N_14061,N_14240);
nand U14353 (N_14353,N_14209,N_14047);
nand U14354 (N_14354,N_14109,N_14104);
nand U14355 (N_14355,N_14174,N_14232);
or U14356 (N_14356,N_14189,N_14176);
nor U14357 (N_14357,N_14128,N_14187);
xnor U14358 (N_14358,N_14111,N_14005);
xnor U14359 (N_14359,N_14092,N_14225);
nand U14360 (N_14360,N_14098,N_14228);
nand U14361 (N_14361,N_14046,N_14136);
xnor U14362 (N_14362,N_14224,N_14181);
and U14363 (N_14363,N_14058,N_14210);
xor U14364 (N_14364,N_14137,N_14159);
or U14365 (N_14365,N_14063,N_14013);
and U14366 (N_14366,N_14119,N_14172);
nor U14367 (N_14367,N_14214,N_14035);
nand U14368 (N_14368,N_14227,N_14030);
nand U14369 (N_14369,N_14088,N_14082);
xnor U14370 (N_14370,N_14049,N_14150);
or U14371 (N_14371,N_14060,N_14197);
or U14372 (N_14372,N_14191,N_14023);
nand U14373 (N_14373,N_14051,N_14166);
xnor U14374 (N_14374,N_14155,N_14016);
and U14375 (N_14375,N_14113,N_14030);
xnor U14376 (N_14376,N_14048,N_14015);
or U14377 (N_14377,N_14115,N_14240);
nand U14378 (N_14378,N_14202,N_14147);
nand U14379 (N_14379,N_14111,N_14025);
and U14380 (N_14380,N_14019,N_14208);
nor U14381 (N_14381,N_14087,N_14150);
xnor U14382 (N_14382,N_14214,N_14065);
and U14383 (N_14383,N_14145,N_14035);
nand U14384 (N_14384,N_14028,N_14196);
or U14385 (N_14385,N_14224,N_14147);
xor U14386 (N_14386,N_14212,N_14193);
nor U14387 (N_14387,N_14042,N_14173);
and U14388 (N_14388,N_14118,N_14180);
or U14389 (N_14389,N_14104,N_14229);
and U14390 (N_14390,N_14035,N_14231);
nor U14391 (N_14391,N_14030,N_14059);
xnor U14392 (N_14392,N_14014,N_14043);
or U14393 (N_14393,N_14056,N_14218);
or U14394 (N_14394,N_14175,N_14168);
and U14395 (N_14395,N_14195,N_14057);
nand U14396 (N_14396,N_14061,N_14150);
nand U14397 (N_14397,N_14076,N_14141);
or U14398 (N_14398,N_14211,N_14078);
and U14399 (N_14399,N_14124,N_14133);
xor U14400 (N_14400,N_14054,N_14046);
nand U14401 (N_14401,N_14228,N_14173);
xnor U14402 (N_14402,N_14168,N_14173);
and U14403 (N_14403,N_14102,N_14214);
and U14404 (N_14404,N_14186,N_14039);
nor U14405 (N_14405,N_14154,N_14078);
nand U14406 (N_14406,N_14122,N_14047);
xor U14407 (N_14407,N_14194,N_14142);
and U14408 (N_14408,N_14170,N_14189);
nand U14409 (N_14409,N_14205,N_14194);
nor U14410 (N_14410,N_14111,N_14067);
nor U14411 (N_14411,N_14100,N_14197);
nor U14412 (N_14412,N_14246,N_14000);
nand U14413 (N_14413,N_14131,N_14239);
and U14414 (N_14414,N_14009,N_14034);
nand U14415 (N_14415,N_14160,N_14061);
nand U14416 (N_14416,N_14022,N_14118);
and U14417 (N_14417,N_14233,N_14055);
xnor U14418 (N_14418,N_14163,N_14094);
or U14419 (N_14419,N_14234,N_14029);
or U14420 (N_14420,N_14116,N_14167);
xnor U14421 (N_14421,N_14013,N_14238);
and U14422 (N_14422,N_14103,N_14141);
and U14423 (N_14423,N_14171,N_14025);
or U14424 (N_14424,N_14018,N_14023);
nand U14425 (N_14425,N_14238,N_14026);
and U14426 (N_14426,N_14011,N_14188);
xnor U14427 (N_14427,N_14220,N_14231);
nor U14428 (N_14428,N_14140,N_14220);
nand U14429 (N_14429,N_14112,N_14049);
xnor U14430 (N_14430,N_14025,N_14055);
and U14431 (N_14431,N_14166,N_14174);
nor U14432 (N_14432,N_14023,N_14048);
nor U14433 (N_14433,N_14082,N_14236);
nor U14434 (N_14434,N_14100,N_14051);
nand U14435 (N_14435,N_14229,N_14135);
nand U14436 (N_14436,N_14187,N_14088);
nor U14437 (N_14437,N_14086,N_14108);
nand U14438 (N_14438,N_14000,N_14051);
and U14439 (N_14439,N_14228,N_14064);
or U14440 (N_14440,N_14157,N_14229);
xnor U14441 (N_14441,N_14147,N_14021);
and U14442 (N_14442,N_14127,N_14229);
nor U14443 (N_14443,N_14151,N_14176);
xor U14444 (N_14444,N_14227,N_14052);
nor U14445 (N_14445,N_14045,N_14221);
or U14446 (N_14446,N_14196,N_14227);
and U14447 (N_14447,N_14152,N_14249);
nor U14448 (N_14448,N_14243,N_14131);
nor U14449 (N_14449,N_14017,N_14233);
or U14450 (N_14450,N_14088,N_14165);
nand U14451 (N_14451,N_14126,N_14084);
nand U14452 (N_14452,N_14059,N_14247);
nand U14453 (N_14453,N_14187,N_14226);
or U14454 (N_14454,N_14137,N_14026);
or U14455 (N_14455,N_14146,N_14249);
and U14456 (N_14456,N_14078,N_14011);
nand U14457 (N_14457,N_14042,N_14129);
xnor U14458 (N_14458,N_14031,N_14129);
and U14459 (N_14459,N_14193,N_14135);
or U14460 (N_14460,N_14238,N_14157);
and U14461 (N_14461,N_14249,N_14049);
nand U14462 (N_14462,N_14110,N_14058);
nand U14463 (N_14463,N_14218,N_14189);
xnor U14464 (N_14464,N_14054,N_14146);
or U14465 (N_14465,N_14088,N_14116);
xor U14466 (N_14466,N_14061,N_14133);
nand U14467 (N_14467,N_14192,N_14137);
and U14468 (N_14468,N_14002,N_14016);
nor U14469 (N_14469,N_14058,N_14109);
nand U14470 (N_14470,N_14016,N_14130);
and U14471 (N_14471,N_14104,N_14237);
or U14472 (N_14472,N_14224,N_14038);
nand U14473 (N_14473,N_14070,N_14094);
and U14474 (N_14474,N_14182,N_14113);
nor U14475 (N_14475,N_14182,N_14228);
nor U14476 (N_14476,N_14016,N_14148);
nor U14477 (N_14477,N_14027,N_14233);
or U14478 (N_14478,N_14191,N_14213);
nand U14479 (N_14479,N_14121,N_14003);
nand U14480 (N_14480,N_14131,N_14208);
nor U14481 (N_14481,N_14212,N_14033);
nor U14482 (N_14482,N_14023,N_14203);
nand U14483 (N_14483,N_14040,N_14167);
and U14484 (N_14484,N_14169,N_14214);
and U14485 (N_14485,N_14013,N_14076);
xnor U14486 (N_14486,N_14109,N_14014);
nand U14487 (N_14487,N_14052,N_14050);
nor U14488 (N_14488,N_14024,N_14121);
nand U14489 (N_14489,N_14074,N_14118);
nand U14490 (N_14490,N_14172,N_14045);
and U14491 (N_14491,N_14038,N_14095);
xnor U14492 (N_14492,N_14218,N_14200);
nor U14493 (N_14493,N_14137,N_14115);
nand U14494 (N_14494,N_14161,N_14092);
nor U14495 (N_14495,N_14010,N_14036);
xor U14496 (N_14496,N_14000,N_14209);
nand U14497 (N_14497,N_14121,N_14082);
or U14498 (N_14498,N_14023,N_14053);
nor U14499 (N_14499,N_14032,N_14146);
nand U14500 (N_14500,N_14468,N_14298);
xnor U14501 (N_14501,N_14276,N_14417);
nor U14502 (N_14502,N_14410,N_14332);
nand U14503 (N_14503,N_14403,N_14493);
xnor U14504 (N_14504,N_14436,N_14443);
xor U14505 (N_14505,N_14408,N_14322);
nor U14506 (N_14506,N_14371,N_14350);
nand U14507 (N_14507,N_14455,N_14373);
and U14508 (N_14508,N_14255,N_14479);
and U14509 (N_14509,N_14307,N_14301);
nand U14510 (N_14510,N_14385,N_14454);
and U14511 (N_14511,N_14294,N_14377);
nor U14512 (N_14512,N_14426,N_14413);
and U14513 (N_14513,N_14415,N_14305);
xnor U14514 (N_14514,N_14324,N_14334);
nand U14515 (N_14515,N_14351,N_14388);
xor U14516 (N_14516,N_14459,N_14288);
xor U14517 (N_14517,N_14411,N_14353);
nand U14518 (N_14518,N_14318,N_14378);
nor U14519 (N_14519,N_14489,N_14375);
or U14520 (N_14520,N_14266,N_14354);
nand U14521 (N_14521,N_14262,N_14372);
and U14522 (N_14522,N_14390,N_14268);
nor U14523 (N_14523,N_14293,N_14337);
or U14524 (N_14524,N_14445,N_14333);
nor U14525 (N_14525,N_14289,N_14303);
xor U14526 (N_14526,N_14446,N_14453);
nor U14527 (N_14527,N_14323,N_14279);
nor U14528 (N_14528,N_14269,N_14496);
nor U14529 (N_14529,N_14250,N_14327);
nor U14530 (N_14530,N_14418,N_14290);
nor U14531 (N_14531,N_14484,N_14286);
nor U14532 (N_14532,N_14486,N_14430);
or U14533 (N_14533,N_14363,N_14437);
nor U14534 (N_14534,N_14365,N_14469);
nor U14535 (N_14535,N_14397,N_14358);
and U14536 (N_14536,N_14355,N_14304);
nand U14537 (N_14537,N_14259,N_14348);
nor U14538 (N_14538,N_14389,N_14423);
xnor U14539 (N_14539,N_14253,N_14257);
and U14540 (N_14540,N_14464,N_14435);
and U14541 (N_14541,N_14449,N_14414);
nand U14542 (N_14542,N_14312,N_14483);
nand U14543 (N_14543,N_14267,N_14499);
nand U14544 (N_14544,N_14431,N_14328);
xor U14545 (N_14545,N_14292,N_14405);
nand U14546 (N_14546,N_14462,N_14317);
and U14547 (N_14547,N_14452,N_14357);
nor U14548 (N_14548,N_14321,N_14297);
nor U14549 (N_14549,N_14367,N_14319);
and U14550 (N_14550,N_14391,N_14396);
nor U14551 (N_14551,N_14394,N_14458);
or U14552 (N_14552,N_14275,N_14370);
and U14553 (N_14553,N_14441,N_14299);
or U14554 (N_14554,N_14335,N_14368);
nand U14555 (N_14555,N_14252,N_14477);
and U14556 (N_14556,N_14326,N_14399);
nand U14557 (N_14557,N_14448,N_14444);
or U14558 (N_14558,N_14361,N_14395);
or U14559 (N_14559,N_14495,N_14482);
nand U14560 (N_14560,N_14256,N_14420);
xnor U14561 (N_14561,N_14472,N_14313);
nand U14562 (N_14562,N_14473,N_14341);
nor U14563 (N_14563,N_14382,N_14310);
and U14564 (N_14564,N_14331,N_14471);
nand U14565 (N_14565,N_14295,N_14284);
and U14566 (N_14566,N_14384,N_14460);
xor U14567 (N_14567,N_14416,N_14419);
xnor U14568 (N_14568,N_14342,N_14283);
nand U14569 (N_14569,N_14258,N_14308);
xnor U14570 (N_14570,N_14381,N_14466);
nor U14571 (N_14571,N_14362,N_14380);
nand U14572 (N_14572,N_14271,N_14254);
nor U14573 (N_14573,N_14470,N_14467);
and U14574 (N_14574,N_14442,N_14425);
or U14575 (N_14575,N_14315,N_14270);
nand U14576 (N_14576,N_14360,N_14424);
xor U14577 (N_14577,N_14386,N_14406);
or U14578 (N_14578,N_14329,N_14383);
xor U14579 (N_14579,N_14475,N_14277);
nand U14580 (N_14580,N_14407,N_14440);
xnor U14581 (N_14581,N_14490,N_14339);
and U14582 (N_14582,N_14369,N_14494);
xor U14583 (N_14583,N_14278,N_14392);
and U14584 (N_14584,N_14401,N_14359);
nand U14585 (N_14585,N_14487,N_14345);
xor U14586 (N_14586,N_14264,N_14480);
xnor U14587 (N_14587,N_14497,N_14447);
nand U14588 (N_14588,N_14439,N_14352);
or U14589 (N_14589,N_14461,N_14433);
xnor U14590 (N_14590,N_14478,N_14398);
or U14591 (N_14591,N_14402,N_14343);
xor U14592 (N_14592,N_14302,N_14488);
and U14593 (N_14593,N_14338,N_14265);
nor U14594 (N_14594,N_14393,N_14422);
and U14595 (N_14595,N_14314,N_14296);
nand U14596 (N_14596,N_14465,N_14316);
and U14597 (N_14597,N_14457,N_14412);
nand U14598 (N_14598,N_14320,N_14485);
xor U14599 (N_14599,N_14456,N_14349);
nand U14600 (N_14600,N_14273,N_14387);
xnor U14601 (N_14601,N_14404,N_14260);
nor U14602 (N_14602,N_14374,N_14463);
or U14603 (N_14603,N_14325,N_14340);
or U14604 (N_14604,N_14330,N_14481);
nand U14605 (N_14605,N_14280,N_14366);
and U14606 (N_14606,N_14491,N_14427);
and U14607 (N_14607,N_14300,N_14498);
nor U14608 (N_14608,N_14346,N_14311);
or U14609 (N_14609,N_14356,N_14336);
nand U14610 (N_14610,N_14281,N_14306);
nor U14611 (N_14611,N_14438,N_14451);
xnor U14612 (N_14612,N_14287,N_14400);
nor U14613 (N_14613,N_14421,N_14432);
xor U14614 (N_14614,N_14309,N_14450);
or U14615 (N_14615,N_14364,N_14282);
nor U14616 (N_14616,N_14428,N_14376);
nand U14617 (N_14617,N_14474,N_14492);
nor U14618 (N_14618,N_14344,N_14291);
and U14619 (N_14619,N_14347,N_14251);
nand U14620 (N_14620,N_14274,N_14272);
nor U14621 (N_14621,N_14285,N_14409);
nand U14622 (N_14622,N_14263,N_14379);
and U14623 (N_14623,N_14434,N_14476);
and U14624 (N_14624,N_14429,N_14261);
nand U14625 (N_14625,N_14328,N_14453);
or U14626 (N_14626,N_14431,N_14317);
nor U14627 (N_14627,N_14270,N_14339);
and U14628 (N_14628,N_14291,N_14465);
or U14629 (N_14629,N_14362,N_14484);
and U14630 (N_14630,N_14354,N_14314);
nor U14631 (N_14631,N_14250,N_14283);
xor U14632 (N_14632,N_14402,N_14279);
xnor U14633 (N_14633,N_14475,N_14302);
nand U14634 (N_14634,N_14453,N_14389);
xor U14635 (N_14635,N_14310,N_14494);
or U14636 (N_14636,N_14402,N_14328);
or U14637 (N_14637,N_14358,N_14398);
xnor U14638 (N_14638,N_14331,N_14275);
nand U14639 (N_14639,N_14384,N_14269);
xnor U14640 (N_14640,N_14250,N_14377);
nor U14641 (N_14641,N_14440,N_14485);
xor U14642 (N_14642,N_14402,N_14266);
or U14643 (N_14643,N_14465,N_14306);
or U14644 (N_14644,N_14412,N_14426);
nor U14645 (N_14645,N_14369,N_14426);
and U14646 (N_14646,N_14305,N_14495);
or U14647 (N_14647,N_14262,N_14473);
nand U14648 (N_14648,N_14353,N_14303);
nand U14649 (N_14649,N_14301,N_14393);
nor U14650 (N_14650,N_14273,N_14357);
or U14651 (N_14651,N_14408,N_14394);
and U14652 (N_14652,N_14494,N_14481);
nor U14653 (N_14653,N_14481,N_14478);
nor U14654 (N_14654,N_14277,N_14462);
nor U14655 (N_14655,N_14271,N_14275);
nor U14656 (N_14656,N_14434,N_14371);
nor U14657 (N_14657,N_14357,N_14429);
nor U14658 (N_14658,N_14392,N_14456);
xnor U14659 (N_14659,N_14321,N_14388);
and U14660 (N_14660,N_14495,N_14450);
or U14661 (N_14661,N_14268,N_14484);
or U14662 (N_14662,N_14290,N_14350);
nor U14663 (N_14663,N_14445,N_14302);
or U14664 (N_14664,N_14288,N_14440);
and U14665 (N_14665,N_14345,N_14433);
xor U14666 (N_14666,N_14494,N_14478);
or U14667 (N_14667,N_14343,N_14279);
nand U14668 (N_14668,N_14304,N_14453);
and U14669 (N_14669,N_14429,N_14445);
nor U14670 (N_14670,N_14314,N_14378);
or U14671 (N_14671,N_14365,N_14344);
nand U14672 (N_14672,N_14260,N_14302);
or U14673 (N_14673,N_14388,N_14412);
nor U14674 (N_14674,N_14311,N_14298);
xnor U14675 (N_14675,N_14315,N_14305);
or U14676 (N_14676,N_14494,N_14470);
nand U14677 (N_14677,N_14451,N_14491);
xor U14678 (N_14678,N_14373,N_14448);
xor U14679 (N_14679,N_14463,N_14484);
or U14680 (N_14680,N_14271,N_14341);
xor U14681 (N_14681,N_14410,N_14393);
and U14682 (N_14682,N_14416,N_14263);
or U14683 (N_14683,N_14308,N_14493);
xor U14684 (N_14684,N_14348,N_14301);
nor U14685 (N_14685,N_14289,N_14405);
xor U14686 (N_14686,N_14494,N_14292);
and U14687 (N_14687,N_14422,N_14341);
or U14688 (N_14688,N_14378,N_14292);
and U14689 (N_14689,N_14353,N_14349);
xor U14690 (N_14690,N_14291,N_14420);
nor U14691 (N_14691,N_14469,N_14494);
and U14692 (N_14692,N_14481,N_14447);
and U14693 (N_14693,N_14371,N_14335);
nor U14694 (N_14694,N_14462,N_14263);
nand U14695 (N_14695,N_14458,N_14372);
nor U14696 (N_14696,N_14483,N_14314);
or U14697 (N_14697,N_14265,N_14362);
or U14698 (N_14698,N_14313,N_14422);
or U14699 (N_14699,N_14308,N_14253);
nor U14700 (N_14700,N_14371,N_14494);
nand U14701 (N_14701,N_14298,N_14320);
nor U14702 (N_14702,N_14461,N_14342);
nand U14703 (N_14703,N_14459,N_14294);
nor U14704 (N_14704,N_14490,N_14294);
nor U14705 (N_14705,N_14395,N_14376);
and U14706 (N_14706,N_14432,N_14440);
and U14707 (N_14707,N_14322,N_14356);
nand U14708 (N_14708,N_14437,N_14371);
nand U14709 (N_14709,N_14371,N_14479);
xnor U14710 (N_14710,N_14380,N_14327);
and U14711 (N_14711,N_14461,N_14450);
and U14712 (N_14712,N_14361,N_14296);
nand U14713 (N_14713,N_14342,N_14355);
nor U14714 (N_14714,N_14423,N_14422);
nand U14715 (N_14715,N_14301,N_14369);
xnor U14716 (N_14716,N_14272,N_14357);
or U14717 (N_14717,N_14372,N_14408);
xnor U14718 (N_14718,N_14382,N_14276);
and U14719 (N_14719,N_14368,N_14455);
nor U14720 (N_14720,N_14250,N_14301);
and U14721 (N_14721,N_14336,N_14464);
nor U14722 (N_14722,N_14482,N_14444);
xnor U14723 (N_14723,N_14327,N_14480);
nand U14724 (N_14724,N_14358,N_14410);
nor U14725 (N_14725,N_14282,N_14474);
nor U14726 (N_14726,N_14482,N_14390);
nor U14727 (N_14727,N_14411,N_14295);
nor U14728 (N_14728,N_14412,N_14442);
nand U14729 (N_14729,N_14420,N_14377);
and U14730 (N_14730,N_14430,N_14446);
nor U14731 (N_14731,N_14468,N_14378);
nand U14732 (N_14732,N_14443,N_14441);
nand U14733 (N_14733,N_14395,N_14308);
and U14734 (N_14734,N_14441,N_14357);
or U14735 (N_14735,N_14358,N_14328);
or U14736 (N_14736,N_14312,N_14361);
nor U14737 (N_14737,N_14314,N_14373);
nor U14738 (N_14738,N_14330,N_14379);
nand U14739 (N_14739,N_14357,N_14266);
and U14740 (N_14740,N_14390,N_14267);
and U14741 (N_14741,N_14257,N_14272);
xnor U14742 (N_14742,N_14269,N_14368);
and U14743 (N_14743,N_14387,N_14382);
nor U14744 (N_14744,N_14367,N_14400);
nor U14745 (N_14745,N_14388,N_14384);
and U14746 (N_14746,N_14435,N_14490);
nor U14747 (N_14747,N_14435,N_14280);
xor U14748 (N_14748,N_14326,N_14286);
nor U14749 (N_14749,N_14291,N_14422);
or U14750 (N_14750,N_14620,N_14612);
or U14751 (N_14751,N_14574,N_14687);
nand U14752 (N_14752,N_14602,N_14582);
nor U14753 (N_14753,N_14586,N_14694);
nor U14754 (N_14754,N_14712,N_14597);
xnor U14755 (N_14755,N_14604,N_14724);
and U14756 (N_14756,N_14549,N_14576);
and U14757 (N_14757,N_14505,N_14606);
xnor U14758 (N_14758,N_14652,N_14584);
and U14759 (N_14759,N_14611,N_14721);
nor U14760 (N_14760,N_14568,N_14720);
nor U14761 (N_14761,N_14745,N_14595);
xor U14762 (N_14762,N_14587,N_14651);
nand U14763 (N_14763,N_14551,N_14544);
or U14764 (N_14764,N_14641,N_14748);
nor U14765 (N_14765,N_14592,N_14547);
xnor U14766 (N_14766,N_14525,N_14569);
and U14767 (N_14767,N_14617,N_14603);
and U14768 (N_14768,N_14645,N_14643);
nand U14769 (N_14769,N_14605,N_14662);
and U14770 (N_14770,N_14685,N_14545);
and U14771 (N_14771,N_14534,N_14577);
or U14772 (N_14772,N_14701,N_14580);
xnor U14773 (N_14773,N_14596,N_14664);
and U14774 (N_14774,N_14585,N_14559);
xor U14775 (N_14775,N_14507,N_14583);
nand U14776 (N_14776,N_14504,N_14625);
xor U14777 (N_14777,N_14570,N_14558);
and U14778 (N_14778,N_14706,N_14675);
nor U14779 (N_14779,N_14591,N_14621);
or U14780 (N_14780,N_14716,N_14635);
or U14781 (N_14781,N_14710,N_14711);
xnor U14782 (N_14782,N_14671,N_14502);
and U14783 (N_14783,N_14698,N_14571);
xor U14784 (N_14784,N_14689,N_14508);
or U14785 (N_14785,N_14561,N_14518);
or U14786 (N_14786,N_14658,N_14676);
or U14787 (N_14787,N_14679,N_14669);
xor U14788 (N_14788,N_14686,N_14734);
nand U14789 (N_14789,N_14510,N_14540);
xnor U14790 (N_14790,N_14736,N_14688);
xor U14791 (N_14791,N_14524,N_14536);
or U14792 (N_14792,N_14632,N_14601);
nand U14793 (N_14793,N_14554,N_14661);
xor U14794 (N_14794,N_14666,N_14619);
and U14795 (N_14795,N_14501,N_14727);
nand U14796 (N_14796,N_14573,N_14581);
nand U14797 (N_14797,N_14503,N_14695);
or U14798 (N_14798,N_14579,N_14644);
nor U14799 (N_14799,N_14743,N_14634);
nand U14800 (N_14800,N_14532,N_14512);
nand U14801 (N_14801,N_14722,N_14697);
xor U14802 (N_14802,N_14715,N_14672);
or U14803 (N_14803,N_14730,N_14589);
nand U14804 (N_14804,N_14673,N_14638);
xor U14805 (N_14805,N_14537,N_14511);
nand U14806 (N_14806,N_14640,N_14588);
or U14807 (N_14807,N_14514,N_14627);
xnor U14808 (N_14808,N_14656,N_14714);
xor U14809 (N_14809,N_14523,N_14509);
nand U14810 (N_14810,N_14531,N_14650);
xnor U14811 (N_14811,N_14705,N_14546);
and U14812 (N_14812,N_14723,N_14533);
or U14813 (N_14813,N_14553,N_14552);
nand U14814 (N_14814,N_14733,N_14657);
nand U14815 (N_14815,N_14667,N_14719);
xnor U14816 (N_14816,N_14648,N_14566);
xnor U14817 (N_14817,N_14642,N_14522);
nor U14818 (N_14818,N_14744,N_14654);
nor U14819 (N_14819,N_14636,N_14702);
or U14820 (N_14820,N_14646,N_14746);
nor U14821 (N_14821,N_14628,N_14622);
xnor U14822 (N_14822,N_14742,N_14665);
nor U14823 (N_14823,N_14680,N_14623);
xnor U14824 (N_14824,N_14629,N_14678);
or U14825 (N_14825,N_14739,N_14737);
nor U14826 (N_14826,N_14521,N_14562);
and U14827 (N_14827,N_14567,N_14613);
or U14828 (N_14828,N_14506,N_14709);
and U14829 (N_14829,N_14563,N_14653);
nor U14830 (N_14830,N_14526,N_14607);
nand U14831 (N_14831,N_14560,N_14631);
or U14832 (N_14832,N_14550,N_14557);
xor U14833 (N_14833,N_14616,N_14543);
or U14834 (N_14834,N_14647,N_14626);
or U14835 (N_14835,N_14699,N_14615);
and U14836 (N_14836,N_14528,N_14707);
nor U14837 (N_14837,N_14614,N_14572);
and U14838 (N_14838,N_14541,N_14538);
xnor U14839 (N_14839,N_14609,N_14683);
or U14840 (N_14840,N_14649,N_14691);
nor U14841 (N_14841,N_14513,N_14741);
or U14842 (N_14842,N_14708,N_14630);
or U14843 (N_14843,N_14735,N_14668);
and U14844 (N_14844,N_14693,N_14729);
and U14845 (N_14845,N_14618,N_14738);
nor U14846 (N_14846,N_14608,N_14725);
and U14847 (N_14847,N_14578,N_14598);
nand U14848 (N_14848,N_14565,N_14703);
nor U14849 (N_14849,N_14556,N_14515);
xor U14850 (N_14850,N_14520,N_14718);
and U14851 (N_14851,N_14594,N_14726);
nand U14852 (N_14852,N_14704,N_14713);
nand U14853 (N_14853,N_14749,N_14663);
xnor U14854 (N_14854,N_14624,N_14555);
and U14855 (N_14855,N_14747,N_14519);
nand U14856 (N_14856,N_14682,N_14681);
and U14857 (N_14857,N_14530,N_14670);
and U14858 (N_14858,N_14575,N_14690);
nand U14859 (N_14859,N_14610,N_14599);
xnor U14860 (N_14860,N_14548,N_14564);
nor U14861 (N_14861,N_14731,N_14535);
and U14862 (N_14862,N_14674,N_14717);
nand U14863 (N_14863,N_14539,N_14516);
and U14864 (N_14864,N_14517,N_14639);
nand U14865 (N_14865,N_14692,N_14659);
or U14866 (N_14866,N_14527,N_14684);
and U14867 (N_14867,N_14677,N_14637);
or U14868 (N_14868,N_14633,N_14732);
or U14869 (N_14869,N_14500,N_14655);
nor U14870 (N_14870,N_14740,N_14529);
or U14871 (N_14871,N_14593,N_14696);
or U14872 (N_14872,N_14728,N_14600);
or U14873 (N_14873,N_14590,N_14542);
xor U14874 (N_14874,N_14660,N_14700);
or U14875 (N_14875,N_14703,N_14741);
xnor U14876 (N_14876,N_14506,N_14594);
nand U14877 (N_14877,N_14552,N_14666);
xor U14878 (N_14878,N_14597,N_14514);
or U14879 (N_14879,N_14606,N_14563);
nor U14880 (N_14880,N_14529,N_14715);
or U14881 (N_14881,N_14729,N_14650);
nor U14882 (N_14882,N_14693,N_14680);
and U14883 (N_14883,N_14656,N_14735);
and U14884 (N_14884,N_14501,N_14605);
xor U14885 (N_14885,N_14709,N_14693);
and U14886 (N_14886,N_14695,N_14694);
and U14887 (N_14887,N_14589,N_14701);
xnor U14888 (N_14888,N_14659,N_14504);
or U14889 (N_14889,N_14542,N_14676);
nand U14890 (N_14890,N_14568,N_14583);
and U14891 (N_14891,N_14556,N_14526);
nor U14892 (N_14892,N_14714,N_14707);
nor U14893 (N_14893,N_14616,N_14724);
xor U14894 (N_14894,N_14701,N_14647);
or U14895 (N_14895,N_14514,N_14652);
and U14896 (N_14896,N_14628,N_14574);
xor U14897 (N_14897,N_14659,N_14729);
nand U14898 (N_14898,N_14601,N_14556);
or U14899 (N_14899,N_14623,N_14721);
and U14900 (N_14900,N_14537,N_14520);
nor U14901 (N_14901,N_14585,N_14744);
or U14902 (N_14902,N_14584,N_14650);
or U14903 (N_14903,N_14508,N_14679);
and U14904 (N_14904,N_14660,N_14707);
nand U14905 (N_14905,N_14528,N_14697);
xnor U14906 (N_14906,N_14701,N_14557);
nand U14907 (N_14907,N_14726,N_14640);
xor U14908 (N_14908,N_14685,N_14507);
and U14909 (N_14909,N_14739,N_14667);
nand U14910 (N_14910,N_14647,N_14680);
and U14911 (N_14911,N_14547,N_14733);
xor U14912 (N_14912,N_14545,N_14706);
nor U14913 (N_14913,N_14671,N_14635);
xnor U14914 (N_14914,N_14587,N_14726);
or U14915 (N_14915,N_14643,N_14647);
nor U14916 (N_14916,N_14637,N_14625);
or U14917 (N_14917,N_14628,N_14687);
nor U14918 (N_14918,N_14616,N_14515);
and U14919 (N_14919,N_14648,N_14641);
nor U14920 (N_14920,N_14602,N_14570);
and U14921 (N_14921,N_14602,N_14696);
nor U14922 (N_14922,N_14541,N_14630);
xor U14923 (N_14923,N_14673,N_14552);
or U14924 (N_14924,N_14632,N_14695);
nor U14925 (N_14925,N_14698,N_14566);
xor U14926 (N_14926,N_14536,N_14560);
nor U14927 (N_14927,N_14695,N_14669);
nand U14928 (N_14928,N_14653,N_14532);
or U14929 (N_14929,N_14733,N_14662);
nor U14930 (N_14930,N_14748,N_14683);
nor U14931 (N_14931,N_14711,N_14644);
xnor U14932 (N_14932,N_14737,N_14643);
xnor U14933 (N_14933,N_14745,N_14564);
xnor U14934 (N_14934,N_14618,N_14730);
nor U14935 (N_14935,N_14636,N_14625);
and U14936 (N_14936,N_14616,N_14628);
xnor U14937 (N_14937,N_14676,N_14580);
or U14938 (N_14938,N_14675,N_14569);
nor U14939 (N_14939,N_14748,N_14552);
nand U14940 (N_14940,N_14666,N_14719);
or U14941 (N_14941,N_14535,N_14555);
or U14942 (N_14942,N_14670,N_14697);
nor U14943 (N_14943,N_14728,N_14695);
nor U14944 (N_14944,N_14614,N_14556);
or U14945 (N_14945,N_14667,N_14727);
nand U14946 (N_14946,N_14640,N_14672);
nand U14947 (N_14947,N_14690,N_14528);
xor U14948 (N_14948,N_14638,N_14659);
nand U14949 (N_14949,N_14542,N_14702);
xor U14950 (N_14950,N_14609,N_14593);
xor U14951 (N_14951,N_14678,N_14649);
nor U14952 (N_14952,N_14704,N_14697);
and U14953 (N_14953,N_14600,N_14660);
or U14954 (N_14954,N_14662,N_14617);
or U14955 (N_14955,N_14535,N_14725);
xor U14956 (N_14956,N_14527,N_14625);
or U14957 (N_14957,N_14596,N_14733);
nand U14958 (N_14958,N_14585,N_14633);
nor U14959 (N_14959,N_14544,N_14611);
or U14960 (N_14960,N_14566,N_14662);
xnor U14961 (N_14961,N_14558,N_14578);
and U14962 (N_14962,N_14728,N_14541);
nand U14963 (N_14963,N_14563,N_14625);
nor U14964 (N_14964,N_14529,N_14697);
nand U14965 (N_14965,N_14707,N_14667);
or U14966 (N_14966,N_14726,N_14671);
and U14967 (N_14967,N_14581,N_14665);
and U14968 (N_14968,N_14551,N_14660);
xor U14969 (N_14969,N_14581,N_14656);
and U14970 (N_14970,N_14529,N_14517);
nor U14971 (N_14971,N_14642,N_14535);
nor U14972 (N_14972,N_14645,N_14664);
and U14973 (N_14973,N_14656,N_14546);
nand U14974 (N_14974,N_14729,N_14667);
nor U14975 (N_14975,N_14640,N_14641);
nor U14976 (N_14976,N_14526,N_14558);
nor U14977 (N_14977,N_14690,N_14599);
xnor U14978 (N_14978,N_14653,N_14657);
xor U14979 (N_14979,N_14583,N_14565);
xnor U14980 (N_14980,N_14627,N_14684);
nand U14981 (N_14981,N_14620,N_14587);
xnor U14982 (N_14982,N_14590,N_14575);
xnor U14983 (N_14983,N_14566,N_14705);
and U14984 (N_14984,N_14585,N_14561);
xor U14985 (N_14985,N_14574,N_14550);
xor U14986 (N_14986,N_14549,N_14584);
or U14987 (N_14987,N_14570,N_14590);
and U14988 (N_14988,N_14604,N_14729);
or U14989 (N_14989,N_14723,N_14677);
or U14990 (N_14990,N_14739,N_14697);
xor U14991 (N_14991,N_14605,N_14547);
or U14992 (N_14992,N_14696,N_14697);
and U14993 (N_14993,N_14655,N_14749);
nor U14994 (N_14994,N_14569,N_14560);
and U14995 (N_14995,N_14715,N_14661);
nor U14996 (N_14996,N_14649,N_14558);
or U14997 (N_14997,N_14552,N_14580);
nand U14998 (N_14998,N_14516,N_14517);
nor U14999 (N_14999,N_14575,N_14678);
xor U15000 (N_15000,N_14994,N_14916);
nor U15001 (N_15001,N_14964,N_14969);
nand U15002 (N_15002,N_14837,N_14775);
nand U15003 (N_15003,N_14892,N_14888);
and U15004 (N_15004,N_14933,N_14787);
nor U15005 (N_15005,N_14829,N_14909);
nand U15006 (N_15006,N_14901,N_14806);
nand U15007 (N_15007,N_14895,N_14820);
and U15008 (N_15008,N_14801,N_14936);
nor U15009 (N_15009,N_14790,N_14776);
nor U15010 (N_15010,N_14755,N_14822);
or U15011 (N_15011,N_14870,N_14867);
nor U15012 (N_15012,N_14952,N_14868);
nor U15013 (N_15013,N_14852,N_14921);
or U15014 (N_15014,N_14900,N_14973);
nand U15015 (N_15015,N_14762,N_14917);
nor U15016 (N_15016,N_14771,N_14983);
and U15017 (N_15017,N_14816,N_14944);
and U15018 (N_15018,N_14962,N_14919);
or U15019 (N_15019,N_14785,N_14751);
or U15020 (N_15020,N_14881,N_14815);
or U15021 (N_15021,N_14766,N_14835);
or U15022 (N_15022,N_14929,N_14890);
nand U15023 (N_15023,N_14946,N_14905);
or U15024 (N_15024,N_14911,N_14935);
and U15025 (N_15025,N_14864,N_14937);
or U15026 (N_15026,N_14851,N_14825);
nor U15027 (N_15027,N_14880,N_14834);
nand U15028 (N_15028,N_14780,N_14840);
nor U15029 (N_15029,N_14750,N_14841);
nand U15030 (N_15030,N_14800,N_14794);
and U15031 (N_15031,N_14889,N_14843);
nand U15032 (N_15032,N_14847,N_14989);
nor U15033 (N_15033,N_14949,N_14761);
nor U15034 (N_15034,N_14985,N_14891);
nor U15035 (N_15035,N_14797,N_14981);
or U15036 (N_15036,N_14902,N_14913);
and U15037 (N_15037,N_14967,N_14810);
nor U15038 (N_15038,N_14830,N_14886);
nand U15039 (N_15039,N_14966,N_14939);
and U15040 (N_15040,N_14930,N_14808);
nand U15041 (N_15041,N_14908,N_14999);
nor U15042 (N_15042,N_14791,N_14860);
and U15043 (N_15043,N_14986,N_14907);
nor U15044 (N_15044,N_14831,N_14804);
or U15045 (N_15045,N_14789,N_14849);
and U15046 (N_15046,N_14982,N_14887);
and U15047 (N_15047,N_14977,N_14769);
or U15048 (N_15048,N_14752,N_14846);
or U15049 (N_15049,N_14953,N_14920);
xnor U15050 (N_15050,N_14923,N_14811);
nand U15051 (N_15051,N_14996,N_14833);
nor U15052 (N_15052,N_14903,N_14926);
nor U15053 (N_15053,N_14987,N_14842);
or U15054 (N_15054,N_14948,N_14968);
nand U15055 (N_15055,N_14814,N_14875);
and U15056 (N_15056,N_14839,N_14878);
xnor U15057 (N_15057,N_14971,N_14813);
xor U15058 (N_15058,N_14898,N_14853);
nand U15059 (N_15059,N_14912,N_14854);
nor U15060 (N_15060,N_14786,N_14970);
nor U15061 (N_15061,N_14845,N_14947);
nand U15062 (N_15062,N_14956,N_14772);
nor U15063 (N_15063,N_14894,N_14865);
or U15064 (N_15064,N_14826,N_14945);
nand U15065 (N_15065,N_14979,N_14941);
and U15066 (N_15066,N_14836,N_14893);
or U15067 (N_15067,N_14988,N_14856);
nand U15068 (N_15068,N_14799,N_14992);
nand U15069 (N_15069,N_14897,N_14899);
or U15070 (N_15070,N_14803,N_14809);
nor U15071 (N_15071,N_14960,N_14765);
nand U15072 (N_15072,N_14998,N_14906);
or U15073 (N_15073,N_14774,N_14796);
nand U15074 (N_15074,N_14873,N_14757);
or U15075 (N_15075,N_14858,N_14884);
and U15076 (N_15076,N_14940,N_14980);
xor U15077 (N_15077,N_14753,N_14793);
xnor U15078 (N_15078,N_14764,N_14934);
and U15079 (N_15079,N_14759,N_14778);
or U15080 (N_15080,N_14975,N_14754);
xnor U15081 (N_15081,N_14871,N_14783);
or U15082 (N_15082,N_14914,N_14758);
or U15083 (N_15083,N_14844,N_14848);
nor U15084 (N_15084,N_14788,N_14876);
or U15085 (N_15085,N_14984,N_14925);
nand U15086 (N_15086,N_14861,N_14927);
nand U15087 (N_15087,N_14823,N_14874);
xor U15088 (N_15088,N_14859,N_14931);
nor U15089 (N_15089,N_14974,N_14792);
nor U15090 (N_15090,N_14805,N_14918);
nand U15091 (N_15091,N_14862,N_14756);
nor U15092 (N_15092,N_14812,N_14857);
nor U15093 (N_15093,N_14773,N_14869);
xor U15094 (N_15094,N_14954,N_14990);
xnor U15095 (N_15095,N_14777,N_14997);
nand U15096 (N_15096,N_14991,N_14827);
xor U15097 (N_15097,N_14817,N_14958);
nand U15098 (N_15098,N_14763,N_14957);
or U15099 (N_15099,N_14838,N_14781);
nand U15100 (N_15100,N_14782,N_14784);
or U15101 (N_15101,N_14938,N_14795);
xnor U15102 (N_15102,N_14882,N_14928);
nand U15103 (N_15103,N_14866,N_14767);
or U15104 (N_15104,N_14972,N_14879);
or U15105 (N_15105,N_14961,N_14819);
nor U15106 (N_15106,N_14850,N_14828);
or U15107 (N_15107,N_14832,N_14872);
xor U15108 (N_15108,N_14922,N_14779);
nor U15109 (N_15109,N_14965,N_14885);
or U15110 (N_15110,N_14924,N_14976);
xnor U15111 (N_15111,N_14915,N_14942);
or U15112 (N_15112,N_14877,N_14978);
and U15113 (N_15113,N_14950,N_14821);
xor U15114 (N_15114,N_14932,N_14768);
or U15115 (N_15115,N_14995,N_14959);
and U15116 (N_15116,N_14943,N_14963);
and U15117 (N_15117,N_14798,N_14863);
nor U15118 (N_15118,N_14910,N_14802);
xnor U15119 (N_15119,N_14824,N_14904);
nand U15120 (N_15120,N_14818,N_14760);
nor U15121 (N_15121,N_14955,N_14883);
or U15122 (N_15122,N_14993,N_14951);
or U15123 (N_15123,N_14896,N_14770);
and U15124 (N_15124,N_14855,N_14807);
xor U15125 (N_15125,N_14881,N_14993);
nand U15126 (N_15126,N_14797,N_14750);
and U15127 (N_15127,N_14912,N_14893);
nand U15128 (N_15128,N_14952,N_14904);
nor U15129 (N_15129,N_14835,N_14846);
nor U15130 (N_15130,N_14951,N_14826);
and U15131 (N_15131,N_14982,N_14896);
and U15132 (N_15132,N_14866,N_14937);
nor U15133 (N_15133,N_14833,N_14835);
nor U15134 (N_15134,N_14889,N_14803);
nor U15135 (N_15135,N_14838,N_14792);
and U15136 (N_15136,N_14862,N_14773);
xor U15137 (N_15137,N_14885,N_14937);
or U15138 (N_15138,N_14762,N_14951);
nand U15139 (N_15139,N_14903,N_14782);
nand U15140 (N_15140,N_14845,N_14898);
or U15141 (N_15141,N_14998,N_14865);
xnor U15142 (N_15142,N_14929,N_14817);
and U15143 (N_15143,N_14828,N_14774);
xor U15144 (N_15144,N_14825,N_14781);
nor U15145 (N_15145,N_14966,N_14929);
nor U15146 (N_15146,N_14974,N_14962);
and U15147 (N_15147,N_14778,N_14840);
and U15148 (N_15148,N_14966,N_14841);
or U15149 (N_15149,N_14953,N_14840);
or U15150 (N_15150,N_14904,N_14913);
xnor U15151 (N_15151,N_14856,N_14980);
and U15152 (N_15152,N_14773,N_14946);
or U15153 (N_15153,N_14760,N_14946);
xnor U15154 (N_15154,N_14868,N_14969);
nor U15155 (N_15155,N_14841,N_14765);
nand U15156 (N_15156,N_14753,N_14924);
and U15157 (N_15157,N_14881,N_14790);
nor U15158 (N_15158,N_14976,N_14951);
nor U15159 (N_15159,N_14754,N_14791);
nand U15160 (N_15160,N_14767,N_14854);
nand U15161 (N_15161,N_14971,N_14970);
nor U15162 (N_15162,N_14863,N_14960);
nand U15163 (N_15163,N_14876,N_14995);
and U15164 (N_15164,N_14925,N_14885);
nor U15165 (N_15165,N_14839,N_14968);
and U15166 (N_15166,N_14756,N_14963);
nor U15167 (N_15167,N_14756,N_14990);
xor U15168 (N_15168,N_14774,N_14753);
and U15169 (N_15169,N_14776,N_14972);
nor U15170 (N_15170,N_14793,N_14851);
nand U15171 (N_15171,N_14907,N_14899);
nand U15172 (N_15172,N_14980,N_14812);
nor U15173 (N_15173,N_14950,N_14884);
nand U15174 (N_15174,N_14959,N_14984);
nor U15175 (N_15175,N_14755,N_14950);
nor U15176 (N_15176,N_14790,N_14786);
nor U15177 (N_15177,N_14785,N_14912);
nand U15178 (N_15178,N_14873,N_14905);
xor U15179 (N_15179,N_14840,N_14917);
xor U15180 (N_15180,N_14753,N_14940);
nor U15181 (N_15181,N_14801,N_14979);
or U15182 (N_15182,N_14787,N_14807);
nor U15183 (N_15183,N_14860,N_14907);
and U15184 (N_15184,N_14909,N_14814);
nand U15185 (N_15185,N_14961,N_14949);
xor U15186 (N_15186,N_14954,N_14946);
nand U15187 (N_15187,N_14964,N_14837);
xnor U15188 (N_15188,N_14856,N_14906);
nor U15189 (N_15189,N_14786,N_14989);
or U15190 (N_15190,N_14944,N_14802);
or U15191 (N_15191,N_14995,N_14852);
or U15192 (N_15192,N_14855,N_14884);
nand U15193 (N_15193,N_14991,N_14868);
nand U15194 (N_15194,N_14877,N_14885);
xor U15195 (N_15195,N_14765,N_14838);
xor U15196 (N_15196,N_14855,N_14975);
nand U15197 (N_15197,N_14966,N_14792);
xnor U15198 (N_15198,N_14970,N_14943);
or U15199 (N_15199,N_14823,N_14783);
or U15200 (N_15200,N_14911,N_14773);
nor U15201 (N_15201,N_14807,N_14937);
and U15202 (N_15202,N_14922,N_14882);
nand U15203 (N_15203,N_14963,N_14818);
xor U15204 (N_15204,N_14761,N_14873);
nand U15205 (N_15205,N_14868,N_14886);
and U15206 (N_15206,N_14829,N_14805);
and U15207 (N_15207,N_14962,N_14996);
and U15208 (N_15208,N_14763,N_14869);
nor U15209 (N_15209,N_14870,N_14916);
xnor U15210 (N_15210,N_14766,N_14909);
and U15211 (N_15211,N_14988,N_14874);
xnor U15212 (N_15212,N_14957,N_14810);
nor U15213 (N_15213,N_14820,N_14930);
and U15214 (N_15214,N_14791,N_14811);
or U15215 (N_15215,N_14930,N_14827);
and U15216 (N_15216,N_14897,N_14823);
xnor U15217 (N_15217,N_14968,N_14854);
and U15218 (N_15218,N_14780,N_14980);
xnor U15219 (N_15219,N_14788,N_14958);
nand U15220 (N_15220,N_14752,N_14997);
or U15221 (N_15221,N_14873,N_14893);
xnor U15222 (N_15222,N_14980,N_14880);
nand U15223 (N_15223,N_14757,N_14795);
and U15224 (N_15224,N_14996,N_14943);
and U15225 (N_15225,N_14901,N_14940);
and U15226 (N_15226,N_14762,N_14882);
or U15227 (N_15227,N_14845,N_14920);
xor U15228 (N_15228,N_14874,N_14834);
or U15229 (N_15229,N_14931,N_14892);
and U15230 (N_15230,N_14783,N_14865);
nand U15231 (N_15231,N_14913,N_14910);
nor U15232 (N_15232,N_14955,N_14982);
and U15233 (N_15233,N_14858,N_14772);
or U15234 (N_15234,N_14768,N_14753);
nand U15235 (N_15235,N_14885,N_14984);
or U15236 (N_15236,N_14929,N_14872);
nor U15237 (N_15237,N_14867,N_14893);
nor U15238 (N_15238,N_14787,N_14844);
or U15239 (N_15239,N_14921,N_14904);
xor U15240 (N_15240,N_14842,N_14938);
nand U15241 (N_15241,N_14801,N_14875);
and U15242 (N_15242,N_14840,N_14908);
xnor U15243 (N_15243,N_14830,N_14973);
xnor U15244 (N_15244,N_14855,N_14777);
nor U15245 (N_15245,N_14936,N_14922);
xnor U15246 (N_15246,N_14917,N_14934);
xnor U15247 (N_15247,N_14948,N_14958);
or U15248 (N_15248,N_14868,N_14764);
nor U15249 (N_15249,N_14878,N_14814);
nand U15250 (N_15250,N_15237,N_15137);
or U15251 (N_15251,N_15185,N_15199);
and U15252 (N_15252,N_15187,N_15089);
nor U15253 (N_15253,N_15078,N_15160);
nand U15254 (N_15254,N_15061,N_15088);
nand U15255 (N_15255,N_15245,N_15030);
and U15256 (N_15256,N_15010,N_15121);
nor U15257 (N_15257,N_15198,N_15249);
xnor U15258 (N_15258,N_15114,N_15039);
nand U15259 (N_15259,N_15101,N_15075);
and U15260 (N_15260,N_15054,N_15164);
xnor U15261 (N_15261,N_15124,N_15184);
and U15262 (N_15262,N_15055,N_15023);
nor U15263 (N_15263,N_15177,N_15133);
nand U15264 (N_15264,N_15085,N_15144);
nand U15265 (N_15265,N_15041,N_15072);
xnor U15266 (N_15266,N_15169,N_15224);
and U15267 (N_15267,N_15231,N_15146);
xor U15268 (N_15268,N_15035,N_15062);
xor U15269 (N_15269,N_15194,N_15046);
nand U15270 (N_15270,N_15248,N_15097);
nor U15271 (N_15271,N_15213,N_15093);
nor U15272 (N_15272,N_15174,N_15135);
or U15273 (N_15273,N_15025,N_15090);
or U15274 (N_15274,N_15215,N_15212);
nand U15275 (N_15275,N_15189,N_15209);
or U15276 (N_15276,N_15107,N_15067);
and U15277 (N_15277,N_15206,N_15105);
nand U15278 (N_15278,N_15193,N_15110);
xnor U15279 (N_15279,N_15118,N_15115);
and U15280 (N_15280,N_15226,N_15175);
nor U15281 (N_15281,N_15017,N_15197);
nand U15282 (N_15282,N_15051,N_15071);
nor U15283 (N_15283,N_15087,N_15019);
xor U15284 (N_15284,N_15211,N_15241);
xor U15285 (N_15285,N_15070,N_15148);
and U15286 (N_15286,N_15021,N_15242);
and U15287 (N_15287,N_15000,N_15130);
nand U15288 (N_15288,N_15106,N_15120);
xnor U15289 (N_15289,N_15139,N_15034);
or U15290 (N_15290,N_15003,N_15228);
xnor U15291 (N_15291,N_15165,N_15040);
nand U15292 (N_15292,N_15079,N_15073);
nand U15293 (N_15293,N_15117,N_15082);
and U15294 (N_15294,N_15240,N_15014);
and U15295 (N_15295,N_15173,N_15108);
nand U15296 (N_15296,N_15168,N_15134);
or U15297 (N_15297,N_15200,N_15007);
and U15298 (N_15298,N_15140,N_15050);
and U15299 (N_15299,N_15220,N_15098);
nor U15300 (N_15300,N_15042,N_15151);
nor U15301 (N_15301,N_15233,N_15029);
xnor U15302 (N_15302,N_15103,N_15022);
nand U15303 (N_15303,N_15196,N_15147);
and U15304 (N_15304,N_15102,N_15027);
nand U15305 (N_15305,N_15008,N_15161);
and U15306 (N_15306,N_15011,N_15016);
nand U15307 (N_15307,N_15057,N_15203);
and U15308 (N_15308,N_15052,N_15020);
nor U15309 (N_15309,N_15013,N_15119);
xor U15310 (N_15310,N_15205,N_15192);
nand U15311 (N_15311,N_15063,N_15142);
xnor U15312 (N_15312,N_15032,N_15158);
xnor U15313 (N_15313,N_15081,N_15092);
nor U15314 (N_15314,N_15091,N_15186);
and U15315 (N_15315,N_15127,N_15038);
nand U15316 (N_15316,N_15179,N_15043);
xor U15317 (N_15317,N_15044,N_15112);
nor U15318 (N_15318,N_15170,N_15246);
or U15319 (N_15319,N_15128,N_15176);
xor U15320 (N_15320,N_15214,N_15218);
nor U15321 (N_15321,N_15084,N_15191);
xnor U15322 (N_15322,N_15180,N_15015);
and U15323 (N_15323,N_15138,N_15060);
and U15324 (N_15324,N_15152,N_15005);
xor U15325 (N_15325,N_15210,N_15068);
nor U15326 (N_15326,N_15064,N_15069);
and U15327 (N_15327,N_15178,N_15077);
nor U15328 (N_15328,N_15109,N_15111);
nand U15329 (N_15329,N_15153,N_15033);
nor U15330 (N_15330,N_15065,N_15154);
nand U15331 (N_15331,N_15244,N_15195);
and U15332 (N_15332,N_15056,N_15229);
nand U15333 (N_15333,N_15149,N_15236);
nand U15334 (N_15334,N_15126,N_15181);
or U15335 (N_15335,N_15002,N_15009);
nor U15336 (N_15336,N_15113,N_15141);
xor U15337 (N_15337,N_15156,N_15223);
nand U15338 (N_15338,N_15076,N_15096);
or U15339 (N_15339,N_15216,N_15125);
or U15340 (N_15340,N_15145,N_15190);
nor U15341 (N_15341,N_15235,N_15049);
nor U15342 (N_15342,N_15157,N_15183);
xnor U15343 (N_15343,N_15001,N_15188);
nand U15344 (N_15344,N_15047,N_15058);
or U15345 (N_15345,N_15162,N_15208);
nand U15346 (N_15346,N_15045,N_15159);
xor U15347 (N_15347,N_15132,N_15232);
and U15348 (N_15348,N_15024,N_15086);
xnor U15349 (N_15349,N_15182,N_15201);
or U15350 (N_15350,N_15122,N_15028);
nand U15351 (N_15351,N_15227,N_15116);
nor U15352 (N_15352,N_15074,N_15171);
nor U15353 (N_15353,N_15225,N_15166);
and U15354 (N_15354,N_15053,N_15204);
and U15355 (N_15355,N_15031,N_15004);
and U15356 (N_15356,N_15202,N_15239);
xnor U15357 (N_15357,N_15143,N_15129);
nor U15358 (N_15358,N_15163,N_15095);
and U15359 (N_15359,N_15247,N_15066);
nand U15360 (N_15360,N_15104,N_15217);
nor U15361 (N_15361,N_15238,N_15099);
nand U15362 (N_15362,N_15018,N_15123);
or U15363 (N_15363,N_15167,N_15207);
xnor U15364 (N_15364,N_15048,N_15012);
nor U15365 (N_15365,N_15219,N_15083);
and U15366 (N_15366,N_15136,N_15150);
nor U15367 (N_15367,N_15243,N_15037);
xor U15368 (N_15368,N_15094,N_15059);
nand U15369 (N_15369,N_15222,N_15221);
nor U15370 (N_15370,N_15006,N_15080);
or U15371 (N_15371,N_15100,N_15131);
or U15372 (N_15372,N_15036,N_15155);
xor U15373 (N_15373,N_15230,N_15172);
nand U15374 (N_15374,N_15026,N_15234);
nor U15375 (N_15375,N_15064,N_15100);
or U15376 (N_15376,N_15216,N_15217);
xor U15377 (N_15377,N_15068,N_15145);
nor U15378 (N_15378,N_15058,N_15089);
nand U15379 (N_15379,N_15177,N_15226);
nor U15380 (N_15380,N_15158,N_15205);
or U15381 (N_15381,N_15055,N_15202);
nand U15382 (N_15382,N_15017,N_15041);
xnor U15383 (N_15383,N_15047,N_15010);
nand U15384 (N_15384,N_15202,N_15194);
nor U15385 (N_15385,N_15159,N_15162);
nand U15386 (N_15386,N_15032,N_15054);
or U15387 (N_15387,N_15097,N_15054);
and U15388 (N_15388,N_15125,N_15046);
nand U15389 (N_15389,N_15205,N_15130);
nor U15390 (N_15390,N_15203,N_15194);
nor U15391 (N_15391,N_15167,N_15076);
xnor U15392 (N_15392,N_15100,N_15204);
xor U15393 (N_15393,N_15134,N_15084);
nand U15394 (N_15394,N_15212,N_15054);
and U15395 (N_15395,N_15049,N_15113);
or U15396 (N_15396,N_15011,N_15221);
nor U15397 (N_15397,N_15066,N_15011);
xnor U15398 (N_15398,N_15173,N_15123);
or U15399 (N_15399,N_15230,N_15223);
and U15400 (N_15400,N_15016,N_15064);
xnor U15401 (N_15401,N_15004,N_15086);
nand U15402 (N_15402,N_15246,N_15222);
nor U15403 (N_15403,N_15158,N_15221);
or U15404 (N_15404,N_15148,N_15159);
nor U15405 (N_15405,N_15173,N_15034);
nand U15406 (N_15406,N_15035,N_15190);
and U15407 (N_15407,N_15118,N_15110);
nand U15408 (N_15408,N_15152,N_15140);
nor U15409 (N_15409,N_15083,N_15029);
and U15410 (N_15410,N_15211,N_15025);
xor U15411 (N_15411,N_15156,N_15041);
and U15412 (N_15412,N_15240,N_15038);
nor U15413 (N_15413,N_15108,N_15198);
or U15414 (N_15414,N_15130,N_15094);
or U15415 (N_15415,N_15176,N_15038);
or U15416 (N_15416,N_15233,N_15239);
xor U15417 (N_15417,N_15214,N_15160);
xnor U15418 (N_15418,N_15240,N_15034);
and U15419 (N_15419,N_15007,N_15175);
and U15420 (N_15420,N_15101,N_15001);
xor U15421 (N_15421,N_15059,N_15116);
xnor U15422 (N_15422,N_15219,N_15100);
and U15423 (N_15423,N_15198,N_15233);
nor U15424 (N_15424,N_15127,N_15196);
and U15425 (N_15425,N_15124,N_15188);
and U15426 (N_15426,N_15217,N_15215);
and U15427 (N_15427,N_15162,N_15096);
nand U15428 (N_15428,N_15004,N_15151);
nand U15429 (N_15429,N_15111,N_15234);
nand U15430 (N_15430,N_15121,N_15179);
or U15431 (N_15431,N_15133,N_15030);
xor U15432 (N_15432,N_15170,N_15161);
nand U15433 (N_15433,N_15018,N_15094);
nor U15434 (N_15434,N_15204,N_15046);
xnor U15435 (N_15435,N_15100,N_15142);
nor U15436 (N_15436,N_15239,N_15073);
nand U15437 (N_15437,N_15031,N_15132);
nand U15438 (N_15438,N_15142,N_15184);
and U15439 (N_15439,N_15021,N_15244);
and U15440 (N_15440,N_15016,N_15192);
nor U15441 (N_15441,N_15127,N_15164);
or U15442 (N_15442,N_15103,N_15010);
nand U15443 (N_15443,N_15146,N_15227);
nor U15444 (N_15444,N_15181,N_15235);
xor U15445 (N_15445,N_15228,N_15197);
nor U15446 (N_15446,N_15028,N_15109);
or U15447 (N_15447,N_15070,N_15243);
and U15448 (N_15448,N_15032,N_15248);
nand U15449 (N_15449,N_15064,N_15004);
and U15450 (N_15450,N_15165,N_15020);
nand U15451 (N_15451,N_15233,N_15143);
or U15452 (N_15452,N_15078,N_15081);
and U15453 (N_15453,N_15017,N_15142);
and U15454 (N_15454,N_15201,N_15017);
nand U15455 (N_15455,N_15017,N_15108);
and U15456 (N_15456,N_15036,N_15064);
xor U15457 (N_15457,N_15238,N_15055);
or U15458 (N_15458,N_15003,N_15078);
nand U15459 (N_15459,N_15142,N_15104);
nor U15460 (N_15460,N_15154,N_15186);
xor U15461 (N_15461,N_15121,N_15193);
xnor U15462 (N_15462,N_15019,N_15080);
nor U15463 (N_15463,N_15000,N_15221);
or U15464 (N_15464,N_15028,N_15178);
xnor U15465 (N_15465,N_15235,N_15180);
and U15466 (N_15466,N_15116,N_15068);
nor U15467 (N_15467,N_15066,N_15234);
nand U15468 (N_15468,N_15019,N_15161);
and U15469 (N_15469,N_15199,N_15085);
nand U15470 (N_15470,N_15185,N_15118);
or U15471 (N_15471,N_15231,N_15170);
or U15472 (N_15472,N_15007,N_15181);
or U15473 (N_15473,N_15201,N_15240);
or U15474 (N_15474,N_15201,N_15155);
nor U15475 (N_15475,N_15218,N_15161);
or U15476 (N_15476,N_15228,N_15100);
nor U15477 (N_15477,N_15189,N_15095);
nor U15478 (N_15478,N_15136,N_15010);
nand U15479 (N_15479,N_15088,N_15052);
nor U15480 (N_15480,N_15163,N_15069);
nand U15481 (N_15481,N_15038,N_15189);
nor U15482 (N_15482,N_15030,N_15134);
or U15483 (N_15483,N_15185,N_15204);
nand U15484 (N_15484,N_15136,N_15121);
nor U15485 (N_15485,N_15049,N_15031);
or U15486 (N_15486,N_15048,N_15179);
nand U15487 (N_15487,N_15066,N_15015);
xnor U15488 (N_15488,N_15069,N_15140);
and U15489 (N_15489,N_15042,N_15184);
nor U15490 (N_15490,N_15176,N_15116);
nand U15491 (N_15491,N_15107,N_15207);
xor U15492 (N_15492,N_15240,N_15092);
nor U15493 (N_15493,N_15053,N_15185);
nand U15494 (N_15494,N_15000,N_15184);
or U15495 (N_15495,N_15005,N_15218);
and U15496 (N_15496,N_15167,N_15104);
or U15497 (N_15497,N_15077,N_15185);
or U15498 (N_15498,N_15085,N_15033);
nand U15499 (N_15499,N_15114,N_15185);
xnor U15500 (N_15500,N_15453,N_15358);
xnor U15501 (N_15501,N_15450,N_15250);
nand U15502 (N_15502,N_15407,N_15370);
or U15503 (N_15503,N_15394,N_15472);
or U15504 (N_15504,N_15259,N_15371);
nor U15505 (N_15505,N_15348,N_15436);
nand U15506 (N_15506,N_15486,N_15307);
or U15507 (N_15507,N_15417,N_15405);
or U15508 (N_15508,N_15253,N_15263);
nand U15509 (N_15509,N_15467,N_15313);
nor U15510 (N_15510,N_15306,N_15400);
nor U15511 (N_15511,N_15408,N_15320);
and U15512 (N_15512,N_15283,N_15430);
nand U15513 (N_15513,N_15470,N_15481);
or U15514 (N_15514,N_15369,N_15461);
and U15515 (N_15515,N_15254,N_15305);
or U15516 (N_15516,N_15491,N_15386);
or U15517 (N_15517,N_15361,N_15399);
nor U15518 (N_15518,N_15323,N_15438);
nand U15519 (N_15519,N_15398,N_15496);
and U15520 (N_15520,N_15387,N_15411);
or U15521 (N_15521,N_15356,N_15420);
nor U15522 (N_15522,N_15474,N_15458);
or U15523 (N_15523,N_15298,N_15376);
or U15524 (N_15524,N_15463,N_15375);
nand U15525 (N_15525,N_15485,N_15344);
and U15526 (N_15526,N_15360,N_15302);
or U15527 (N_15527,N_15428,N_15282);
xor U15528 (N_15528,N_15346,N_15395);
xor U15529 (N_15529,N_15340,N_15258);
nand U15530 (N_15530,N_15316,N_15431);
xor U15531 (N_15531,N_15286,N_15264);
nor U15532 (N_15532,N_15442,N_15418);
nand U15533 (N_15533,N_15489,N_15372);
nor U15534 (N_15534,N_15362,N_15350);
nand U15535 (N_15535,N_15357,N_15300);
xnor U15536 (N_15536,N_15331,N_15437);
nand U15537 (N_15537,N_15423,N_15368);
nor U15538 (N_15538,N_15349,N_15390);
and U15539 (N_15539,N_15385,N_15284);
nand U15540 (N_15540,N_15443,N_15303);
and U15541 (N_15541,N_15404,N_15318);
nand U15542 (N_15542,N_15290,N_15392);
and U15543 (N_15543,N_15364,N_15459);
nor U15544 (N_15544,N_15280,N_15338);
xor U15545 (N_15545,N_15476,N_15382);
or U15546 (N_15546,N_15359,N_15268);
nor U15547 (N_15547,N_15292,N_15273);
nand U15548 (N_15548,N_15339,N_15281);
and U15549 (N_15549,N_15389,N_15447);
nor U15550 (N_15550,N_15416,N_15285);
and U15551 (N_15551,N_15352,N_15373);
nor U15552 (N_15552,N_15388,N_15262);
nand U15553 (N_15553,N_15310,N_15278);
xor U15554 (N_15554,N_15335,N_15427);
nor U15555 (N_15555,N_15412,N_15363);
or U15556 (N_15556,N_15478,N_15435);
and U15557 (N_15557,N_15276,N_15299);
xor U15558 (N_15558,N_15308,N_15272);
or U15559 (N_15559,N_15311,N_15391);
xnor U15560 (N_15560,N_15469,N_15291);
nor U15561 (N_15561,N_15457,N_15462);
nor U15562 (N_15562,N_15499,N_15354);
xor U15563 (N_15563,N_15379,N_15434);
nand U15564 (N_15564,N_15410,N_15295);
nor U15565 (N_15565,N_15322,N_15465);
or U15566 (N_15566,N_15269,N_15256);
or U15567 (N_15567,N_15402,N_15275);
and U15568 (N_15568,N_15294,N_15460);
nor U15569 (N_15569,N_15381,N_15468);
xor U15570 (N_15570,N_15317,N_15332);
nor U15571 (N_15571,N_15304,N_15419);
or U15572 (N_15572,N_15498,N_15315);
or U15573 (N_15573,N_15367,N_15255);
and U15574 (N_15574,N_15270,N_15384);
nand U15575 (N_15575,N_15251,N_15330);
or U15576 (N_15576,N_15445,N_15342);
or U15577 (N_15577,N_15271,N_15347);
and U15578 (N_15578,N_15495,N_15464);
or U15579 (N_15579,N_15403,N_15477);
and U15580 (N_15580,N_15426,N_15260);
nor U15581 (N_15581,N_15380,N_15257);
or U15582 (N_15582,N_15482,N_15494);
xor U15583 (N_15583,N_15265,N_15433);
xor U15584 (N_15584,N_15440,N_15483);
nand U15585 (N_15585,N_15454,N_15393);
or U15586 (N_15586,N_15479,N_15296);
or U15587 (N_15587,N_15309,N_15456);
nand U15588 (N_15588,N_15415,N_15425);
nand U15589 (N_15589,N_15424,N_15378);
and U15590 (N_15590,N_15466,N_15343);
xor U15591 (N_15591,N_15473,N_15328);
xor U15592 (N_15592,N_15288,N_15488);
and U15593 (N_15593,N_15374,N_15324);
xor U15594 (N_15594,N_15429,N_15365);
or U15595 (N_15595,N_15321,N_15441);
nand U15596 (N_15596,N_15471,N_15439);
nand U15597 (N_15597,N_15396,N_15266);
nand U15598 (N_15598,N_15345,N_15487);
nor U15599 (N_15599,N_15314,N_15261);
nand U15600 (N_15600,N_15490,N_15401);
and U15601 (N_15601,N_15334,N_15326);
xor U15602 (N_15602,N_15252,N_15449);
xnor U15603 (N_15603,N_15422,N_15337);
xor U15604 (N_15604,N_15366,N_15414);
nor U15605 (N_15605,N_15409,N_15432);
or U15606 (N_15606,N_15383,N_15444);
nor U15607 (N_15607,N_15319,N_15274);
or U15608 (N_15608,N_15492,N_15325);
nor U15609 (N_15609,N_15297,N_15353);
or U15610 (N_15610,N_15448,N_15267);
nand U15611 (N_15611,N_15279,N_15277);
or U15612 (N_15612,N_15293,N_15287);
xnor U15613 (N_15613,N_15493,N_15312);
or U15614 (N_15614,N_15406,N_15327);
xnor U15615 (N_15615,N_15452,N_15336);
nand U15616 (N_15616,N_15475,N_15455);
nor U15617 (N_15617,N_15451,N_15480);
or U15618 (N_15618,N_15497,N_15446);
nor U15619 (N_15619,N_15484,N_15301);
and U15620 (N_15620,N_15397,N_15355);
nand U15621 (N_15621,N_15329,N_15351);
xnor U15622 (N_15622,N_15333,N_15341);
or U15623 (N_15623,N_15289,N_15421);
and U15624 (N_15624,N_15377,N_15413);
nor U15625 (N_15625,N_15323,N_15473);
xnor U15626 (N_15626,N_15390,N_15483);
nand U15627 (N_15627,N_15266,N_15470);
nor U15628 (N_15628,N_15279,N_15309);
and U15629 (N_15629,N_15259,N_15441);
or U15630 (N_15630,N_15288,N_15478);
nand U15631 (N_15631,N_15407,N_15463);
and U15632 (N_15632,N_15351,N_15314);
or U15633 (N_15633,N_15420,N_15451);
xnor U15634 (N_15634,N_15446,N_15391);
xor U15635 (N_15635,N_15260,N_15404);
xnor U15636 (N_15636,N_15414,N_15495);
nor U15637 (N_15637,N_15426,N_15418);
and U15638 (N_15638,N_15441,N_15442);
xnor U15639 (N_15639,N_15457,N_15497);
or U15640 (N_15640,N_15399,N_15301);
and U15641 (N_15641,N_15487,N_15362);
xor U15642 (N_15642,N_15303,N_15434);
nand U15643 (N_15643,N_15253,N_15259);
xnor U15644 (N_15644,N_15279,N_15401);
or U15645 (N_15645,N_15417,N_15283);
nand U15646 (N_15646,N_15449,N_15415);
nand U15647 (N_15647,N_15410,N_15402);
nor U15648 (N_15648,N_15418,N_15340);
and U15649 (N_15649,N_15475,N_15255);
and U15650 (N_15650,N_15423,N_15379);
xor U15651 (N_15651,N_15396,N_15317);
nor U15652 (N_15652,N_15451,N_15346);
nor U15653 (N_15653,N_15486,N_15499);
nor U15654 (N_15654,N_15385,N_15417);
xnor U15655 (N_15655,N_15274,N_15384);
and U15656 (N_15656,N_15270,N_15343);
nand U15657 (N_15657,N_15390,N_15307);
or U15658 (N_15658,N_15300,N_15432);
or U15659 (N_15659,N_15368,N_15487);
and U15660 (N_15660,N_15298,N_15450);
xnor U15661 (N_15661,N_15461,N_15252);
and U15662 (N_15662,N_15347,N_15453);
xor U15663 (N_15663,N_15376,N_15280);
xor U15664 (N_15664,N_15390,N_15393);
and U15665 (N_15665,N_15480,N_15310);
nand U15666 (N_15666,N_15268,N_15478);
nand U15667 (N_15667,N_15272,N_15277);
or U15668 (N_15668,N_15270,N_15361);
xnor U15669 (N_15669,N_15363,N_15432);
xnor U15670 (N_15670,N_15364,N_15318);
nor U15671 (N_15671,N_15296,N_15286);
or U15672 (N_15672,N_15462,N_15471);
nor U15673 (N_15673,N_15262,N_15495);
xnor U15674 (N_15674,N_15384,N_15408);
and U15675 (N_15675,N_15391,N_15275);
or U15676 (N_15676,N_15464,N_15497);
and U15677 (N_15677,N_15438,N_15258);
nand U15678 (N_15678,N_15428,N_15337);
nand U15679 (N_15679,N_15348,N_15282);
xor U15680 (N_15680,N_15374,N_15381);
xor U15681 (N_15681,N_15329,N_15364);
or U15682 (N_15682,N_15257,N_15477);
and U15683 (N_15683,N_15292,N_15380);
and U15684 (N_15684,N_15295,N_15467);
and U15685 (N_15685,N_15274,N_15290);
and U15686 (N_15686,N_15444,N_15471);
xnor U15687 (N_15687,N_15383,N_15494);
or U15688 (N_15688,N_15290,N_15393);
nand U15689 (N_15689,N_15485,N_15417);
and U15690 (N_15690,N_15317,N_15455);
and U15691 (N_15691,N_15420,N_15390);
xor U15692 (N_15692,N_15494,N_15347);
and U15693 (N_15693,N_15434,N_15286);
and U15694 (N_15694,N_15361,N_15455);
nand U15695 (N_15695,N_15474,N_15442);
nor U15696 (N_15696,N_15418,N_15328);
and U15697 (N_15697,N_15291,N_15437);
nand U15698 (N_15698,N_15476,N_15284);
nor U15699 (N_15699,N_15419,N_15458);
nor U15700 (N_15700,N_15307,N_15291);
and U15701 (N_15701,N_15352,N_15261);
nand U15702 (N_15702,N_15401,N_15352);
xnor U15703 (N_15703,N_15250,N_15440);
or U15704 (N_15704,N_15374,N_15267);
or U15705 (N_15705,N_15435,N_15291);
nand U15706 (N_15706,N_15446,N_15404);
xnor U15707 (N_15707,N_15486,N_15445);
xnor U15708 (N_15708,N_15446,N_15409);
or U15709 (N_15709,N_15473,N_15437);
and U15710 (N_15710,N_15408,N_15426);
nand U15711 (N_15711,N_15434,N_15344);
or U15712 (N_15712,N_15460,N_15321);
xor U15713 (N_15713,N_15282,N_15449);
xnor U15714 (N_15714,N_15365,N_15455);
nand U15715 (N_15715,N_15253,N_15368);
xor U15716 (N_15716,N_15301,N_15276);
nand U15717 (N_15717,N_15299,N_15361);
or U15718 (N_15718,N_15283,N_15404);
and U15719 (N_15719,N_15462,N_15491);
and U15720 (N_15720,N_15372,N_15482);
and U15721 (N_15721,N_15423,N_15266);
nand U15722 (N_15722,N_15292,N_15265);
xnor U15723 (N_15723,N_15384,N_15458);
xor U15724 (N_15724,N_15448,N_15405);
xor U15725 (N_15725,N_15294,N_15261);
xor U15726 (N_15726,N_15410,N_15355);
or U15727 (N_15727,N_15294,N_15327);
xor U15728 (N_15728,N_15387,N_15329);
nand U15729 (N_15729,N_15467,N_15326);
nor U15730 (N_15730,N_15294,N_15442);
xnor U15731 (N_15731,N_15432,N_15417);
and U15732 (N_15732,N_15373,N_15378);
nand U15733 (N_15733,N_15250,N_15431);
nor U15734 (N_15734,N_15405,N_15326);
or U15735 (N_15735,N_15368,N_15383);
or U15736 (N_15736,N_15360,N_15300);
or U15737 (N_15737,N_15492,N_15474);
and U15738 (N_15738,N_15284,N_15426);
nand U15739 (N_15739,N_15429,N_15425);
nand U15740 (N_15740,N_15468,N_15348);
nor U15741 (N_15741,N_15270,N_15324);
xor U15742 (N_15742,N_15286,N_15303);
nand U15743 (N_15743,N_15384,N_15388);
nand U15744 (N_15744,N_15405,N_15465);
nor U15745 (N_15745,N_15422,N_15254);
nor U15746 (N_15746,N_15396,N_15485);
xor U15747 (N_15747,N_15340,N_15462);
and U15748 (N_15748,N_15275,N_15321);
and U15749 (N_15749,N_15336,N_15387);
nand U15750 (N_15750,N_15686,N_15644);
xor U15751 (N_15751,N_15585,N_15716);
nor U15752 (N_15752,N_15720,N_15747);
or U15753 (N_15753,N_15661,N_15534);
nand U15754 (N_15754,N_15627,N_15626);
nor U15755 (N_15755,N_15609,N_15641);
xor U15756 (N_15756,N_15633,N_15666);
and U15757 (N_15757,N_15714,N_15547);
nor U15758 (N_15758,N_15517,N_15696);
or U15759 (N_15759,N_15637,N_15630);
xnor U15760 (N_15760,N_15733,N_15638);
or U15761 (N_15761,N_15566,N_15536);
or U15762 (N_15762,N_15724,N_15570);
nand U15763 (N_15763,N_15674,N_15516);
or U15764 (N_15764,N_15510,N_15657);
xnor U15765 (N_15765,N_15634,N_15734);
and U15766 (N_15766,N_15703,N_15655);
or U15767 (N_15767,N_15524,N_15581);
xor U15768 (N_15768,N_15613,N_15550);
and U15769 (N_15769,N_15717,N_15699);
xnor U15770 (N_15770,N_15684,N_15682);
nor U15771 (N_15771,N_15520,N_15571);
xor U15772 (N_15772,N_15515,N_15678);
or U15773 (N_15773,N_15688,N_15642);
nand U15774 (N_15774,N_15615,N_15672);
xor U15775 (N_15775,N_15692,N_15726);
nand U15776 (N_15776,N_15723,N_15731);
or U15777 (N_15777,N_15658,N_15691);
and U15778 (N_15778,N_15737,N_15681);
and U15779 (N_15779,N_15617,N_15710);
xor U15780 (N_15780,N_15586,N_15632);
xor U15781 (N_15781,N_15610,N_15549);
or U15782 (N_15782,N_15677,N_15667);
xor U15783 (N_15783,N_15687,N_15653);
and U15784 (N_15784,N_15537,N_15631);
and U15785 (N_15785,N_15577,N_15611);
and U15786 (N_15786,N_15584,N_15712);
or U15787 (N_15787,N_15521,N_15544);
xor U15788 (N_15788,N_15546,N_15560);
and U15789 (N_15789,N_15588,N_15522);
or U15790 (N_15790,N_15679,N_15513);
xnor U15791 (N_15791,N_15587,N_15551);
and U15792 (N_15792,N_15573,N_15680);
or U15793 (N_15793,N_15623,N_15695);
and U15794 (N_15794,N_15742,N_15545);
xnor U15795 (N_15795,N_15508,N_15523);
xnor U15796 (N_15796,N_15603,N_15740);
xor U15797 (N_15797,N_15507,N_15718);
or U15798 (N_15798,N_15505,N_15738);
xor U15799 (N_15799,N_15527,N_15745);
nand U15800 (N_15800,N_15599,N_15624);
or U15801 (N_15801,N_15572,N_15568);
nor U15802 (N_15802,N_15558,N_15539);
or U15803 (N_15803,N_15705,N_15622);
nor U15804 (N_15804,N_15713,N_15519);
nor U15805 (N_15805,N_15608,N_15746);
nor U15806 (N_15806,N_15582,N_15596);
or U15807 (N_15807,N_15620,N_15744);
nor U15808 (N_15808,N_15612,N_15739);
or U15809 (N_15809,N_15535,N_15518);
and U15810 (N_15810,N_15694,N_15664);
nand U15811 (N_15811,N_15643,N_15646);
nor U15812 (N_15812,N_15589,N_15619);
and U15813 (N_15813,N_15583,N_15567);
or U15814 (N_15814,N_15591,N_15690);
and U15815 (N_15815,N_15715,N_15662);
and U15816 (N_15816,N_15542,N_15594);
nor U15817 (N_15817,N_15698,N_15528);
and U15818 (N_15818,N_15654,N_15530);
nand U15819 (N_15819,N_15579,N_15529);
nor U15820 (N_15820,N_15649,N_15605);
and U15821 (N_15821,N_15748,N_15659);
nor U15822 (N_15822,N_15645,N_15629);
or U15823 (N_15823,N_15693,N_15636);
nor U15824 (N_15824,N_15741,N_15601);
and U15825 (N_15825,N_15554,N_15708);
xnor U15826 (N_15826,N_15541,N_15671);
or U15827 (N_15827,N_15514,N_15711);
and U15828 (N_15828,N_15697,N_15675);
nor U15829 (N_15829,N_15656,N_15721);
nand U15830 (N_15830,N_15700,N_15618);
nor U15831 (N_15831,N_15652,N_15743);
and U15832 (N_15832,N_15562,N_15525);
and U15833 (N_15833,N_15640,N_15729);
nor U15834 (N_15834,N_15668,N_15553);
or U15835 (N_15835,N_15595,N_15673);
or U15836 (N_15836,N_15732,N_15592);
nor U15837 (N_15837,N_15556,N_15735);
xnor U15838 (N_15838,N_15575,N_15559);
nor U15839 (N_15839,N_15580,N_15730);
xor U15840 (N_15840,N_15670,N_15548);
xnor U15841 (N_15841,N_15543,N_15651);
nand U15842 (N_15842,N_15701,N_15621);
and U15843 (N_15843,N_15563,N_15639);
and U15844 (N_15844,N_15531,N_15504);
nand U15845 (N_15845,N_15511,N_15574);
and U15846 (N_15846,N_15614,N_15578);
nand U15847 (N_15847,N_15555,N_15557);
xor U15848 (N_15848,N_15538,N_15606);
xnor U15849 (N_15849,N_15663,N_15593);
nand U15850 (N_15850,N_15533,N_15604);
or U15851 (N_15851,N_15512,N_15625);
nor U15852 (N_15852,N_15707,N_15683);
and U15853 (N_15853,N_15561,N_15564);
and U15854 (N_15854,N_15506,N_15736);
or U15855 (N_15855,N_15749,N_15502);
or U15856 (N_15856,N_15647,N_15576);
xor U15857 (N_15857,N_15725,N_15665);
or U15858 (N_15858,N_15532,N_15685);
xnor U15859 (N_15859,N_15590,N_15628);
xor U15860 (N_15860,N_15602,N_15719);
nand U15861 (N_15861,N_15540,N_15722);
nor U15862 (N_15862,N_15648,N_15616);
xor U15863 (N_15863,N_15706,N_15635);
nor U15864 (N_15864,N_15676,N_15660);
xnor U15865 (N_15865,N_15689,N_15500);
xnor U15866 (N_15866,N_15503,N_15501);
xnor U15867 (N_15867,N_15600,N_15597);
nor U15868 (N_15868,N_15565,N_15702);
and U15869 (N_15869,N_15607,N_15704);
nor U15870 (N_15870,N_15552,N_15509);
and U15871 (N_15871,N_15526,N_15709);
nand U15872 (N_15872,N_15728,N_15669);
nor U15873 (N_15873,N_15598,N_15727);
nor U15874 (N_15874,N_15650,N_15569);
nand U15875 (N_15875,N_15701,N_15721);
or U15876 (N_15876,N_15694,N_15558);
or U15877 (N_15877,N_15656,N_15724);
nand U15878 (N_15878,N_15562,N_15679);
nand U15879 (N_15879,N_15501,N_15505);
and U15880 (N_15880,N_15643,N_15555);
nor U15881 (N_15881,N_15621,N_15581);
nand U15882 (N_15882,N_15742,N_15612);
or U15883 (N_15883,N_15602,N_15630);
nor U15884 (N_15884,N_15732,N_15643);
nor U15885 (N_15885,N_15597,N_15554);
xor U15886 (N_15886,N_15728,N_15696);
and U15887 (N_15887,N_15703,N_15625);
nor U15888 (N_15888,N_15608,N_15612);
or U15889 (N_15889,N_15675,N_15662);
or U15890 (N_15890,N_15741,N_15645);
xnor U15891 (N_15891,N_15549,N_15515);
and U15892 (N_15892,N_15736,N_15699);
nand U15893 (N_15893,N_15543,N_15727);
nand U15894 (N_15894,N_15586,N_15649);
xor U15895 (N_15895,N_15616,N_15559);
xor U15896 (N_15896,N_15723,N_15644);
and U15897 (N_15897,N_15632,N_15688);
or U15898 (N_15898,N_15728,N_15532);
and U15899 (N_15899,N_15685,N_15547);
xor U15900 (N_15900,N_15571,N_15725);
or U15901 (N_15901,N_15508,N_15555);
or U15902 (N_15902,N_15722,N_15606);
or U15903 (N_15903,N_15679,N_15695);
xor U15904 (N_15904,N_15515,N_15654);
or U15905 (N_15905,N_15591,N_15597);
nand U15906 (N_15906,N_15606,N_15739);
or U15907 (N_15907,N_15619,N_15608);
and U15908 (N_15908,N_15672,N_15685);
nor U15909 (N_15909,N_15613,N_15620);
nand U15910 (N_15910,N_15674,N_15583);
nor U15911 (N_15911,N_15518,N_15741);
xnor U15912 (N_15912,N_15576,N_15549);
or U15913 (N_15913,N_15606,N_15567);
or U15914 (N_15914,N_15657,N_15641);
nand U15915 (N_15915,N_15599,N_15734);
nor U15916 (N_15916,N_15621,N_15663);
nand U15917 (N_15917,N_15654,N_15686);
or U15918 (N_15918,N_15680,N_15742);
xor U15919 (N_15919,N_15673,N_15723);
or U15920 (N_15920,N_15613,N_15689);
and U15921 (N_15921,N_15635,N_15606);
nand U15922 (N_15922,N_15581,N_15538);
or U15923 (N_15923,N_15582,N_15610);
nand U15924 (N_15924,N_15500,N_15611);
or U15925 (N_15925,N_15639,N_15636);
nor U15926 (N_15926,N_15689,N_15528);
and U15927 (N_15927,N_15686,N_15543);
xor U15928 (N_15928,N_15652,N_15663);
xnor U15929 (N_15929,N_15692,N_15686);
xor U15930 (N_15930,N_15579,N_15740);
nor U15931 (N_15931,N_15742,N_15542);
nor U15932 (N_15932,N_15506,N_15634);
nor U15933 (N_15933,N_15681,N_15571);
and U15934 (N_15934,N_15555,N_15674);
and U15935 (N_15935,N_15587,N_15673);
nor U15936 (N_15936,N_15734,N_15628);
xnor U15937 (N_15937,N_15712,N_15513);
or U15938 (N_15938,N_15670,N_15713);
nor U15939 (N_15939,N_15536,N_15647);
or U15940 (N_15940,N_15550,N_15596);
and U15941 (N_15941,N_15659,N_15736);
nor U15942 (N_15942,N_15736,N_15557);
and U15943 (N_15943,N_15551,N_15544);
or U15944 (N_15944,N_15646,N_15576);
xnor U15945 (N_15945,N_15745,N_15663);
and U15946 (N_15946,N_15698,N_15564);
nor U15947 (N_15947,N_15683,N_15611);
or U15948 (N_15948,N_15701,N_15559);
or U15949 (N_15949,N_15609,N_15582);
nand U15950 (N_15950,N_15650,N_15667);
nor U15951 (N_15951,N_15659,N_15609);
and U15952 (N_15952,N_15580,N_15733);
nand U15953 (N_15953,N_15520,N_15650);
or U15954 (N_15954,N_15677,N_15597);
nand U15955 (N_15955,N_15562,N_15690);
xnor U15956 (N_15956,N_15593,N_15586);
nor U15957 (N_15957,N_15736,N_15664);
and U15958 (N_15958,N_15578,N_15551);
or U15959 (N_15959,N_15737,N_15721);
nand U15960 (N_15960,N_15585,N_15612);
xor U15961 (N_15961,N_15525,N_15694);
and U15962 (N_15962,N_15742,N_15720);
and U15963 (N_15963,N_15630,N_15634);
nor U15964 (N_15964,N_15618,N_15525);
or U15965 (N_15965,N_15615,N_15543);
nor U15966 (N_15966,N_15690,N_15671);
xor U15967 (N_15967,N_15572,N_15559);
xor U15968 (N_15968,N_15708,N_15599);
nand U15969 (N_15969,N_15669,N_15544);
and U15970 (N_15970,N_15656,N_15541);
and U15971 (N_15971,N_15576,N_15734);
or U15972 (N_15972,N_15549,N_15709);
or U15973 (N_15973,N_15590,N_15711);
xnor U15974 (N_15974,N_15620,N_15681);
xor U15975 (N_15975,N_15529,N_15650);
or U15976 (N_15976,N_15541,N_15612);
and U15977 (N_15977,N_15681,N_15667);
or U15978 (N_15978,N_15709,N_15510);
nor U15979 (N_15979,N_15516,N_15518);
or U15980 (N_15980,N_15610,N_15546);
nand U15981 (N_15981,N_15500,N_15746);
or U15982 (N_15982,N_15571,N_15550);
nand U15983 (N_15983,N_15527,N_15558);
nand U15984 (N_15984,N_15682,N_15552);
or U15985 (N_15985,N_15688,N_15712);
nand U15986 (N_15986,N_15725,N_15519);
and U15987 (N_15987,N_15620,N_15721);
nor U15988 (N_15988,N_15563,N_15572);
nand U15989 (N_15989,N_15670,N_15664);
nand U15990 (N_15990,N_15650,N_15540);
xor U15991 (N_15991,N_15632,N_15560);
or U15992 (N_15992,N_15665,N_15546);
or U15993 (N_15993,N_15650,N_15563);
nand U15994 (N_15994,N_15513,N_15539);
or U15995 (N_15995,N_15732,N_15672);
or U15996 (N_15996,N_15677,N_15524);
xnor U15997 (N_15997,N_15554,N_15749);
and U15998 (N_15998,N_15592,N_15741);
or U15999 (N_15999,N_15510,N_15554);
nor U16000 (N_16000,N_15783,N_15932);
and U16001 (N_16001,N_15992,N_15801);
or U16002 (N_16002,N_15979,N_15848);
nor U16003 (N_16003,N_15876,N_15875);
and U16004 (N_16004,N_15974,N_15991);
or U16005 (N_16005,N_15755,N_15762);
nand U16006 (N_16006,N_15911,N_15832);
xor U16007 (N_16007,N_15931,N_15963);
or U16008 (N_16008,N_15920,N_15822);
nor U16009 (N_16009,N_15926,N_15786);
or U16010 (N_16010,N_15998,N_15781);
nand U16011 (N_16011,N_15784,N_15797);
xnor U16012 (N_16012,N_15942,N_15836);
nand U16013 (N_16013,N_15983,N_15857);
nor U16014 (N_16014,N_15937,N_15810);
and U16015 (N_16015,N_15774,N_15757);
and U16016 (N_16016,N_15856,N_15905);
nand U16017 (N_16017,N_15880,N_15816);
nand U16018 (N_16018,N_15791,N_15788);
and U16019 (N_16019,N_15819,N_15802);
nand U16020 (N_16020,N_15826,N_15956);
and U16021 (N_16021,N_15869,N_15862);
xnor U16022 (N_16022,N_15835,N_15897);
nand U16023 (N_16023,N_15989,N_15976);
and U16024 (N_16024,N_15975,N_15888);
xor U16025 (N_16025,N_15889,N_15868);
and U16026 (N_16026,N_15855,N_15866);
xnor U16027 (N_16027,N_15763,N_15940);
or U16028 (N_16028,N_15957,N_15910);
or U16029 (N_16029,N_15765,N_15767);
nand U16030 (N_16030,N_15815,N_15789);
nor U16031 (N_16031,N_15771,N_15874);
nor U16032 (N_16032,N_15837,N_15756);
nand U16033 (N_16033,N_15898,N_15846);
xor U16034 (N_16034,N_15800,N_15843);
nor U16035 (N_16035,N_15943,N_15923);
nor U16036 (N_16036,N_15944,N_15849);
nand U16037 (N_16037,N_15813,N_15904);
xor U16038 (N_16038,N_15808,N_15844);
nor U16039 (N_16039,N_15759,N_15833);
nor U16040 (N_16040,N_15871,N_15930);
and U16041 (N_16041,N_15891,N_15987);
nor U16042 (N_16042,N_15851,N_15914);
or U16043 (N_16043,N_15896,N_15929);
nand U16044 (N_16044,N_15997,N_15790);
or U16045 (N_16045,N_15761,N_15883);
xor U16046 (N_16046,N_15900,N_15913);
xor U16047 (N_16047,N_15919,N_15793);
and U16048 (N_16048,N_15973,N_15951);
xnor U16049 (N_16049,N_15994,N_15988);
or U16050 (N_16050,N_15894,N_15879);
nand U16051 (N_16051,N_15903,N_15782);
or U16052 (N_16052,N_15799,N_15938);
nor U16053 (N_16053,N_15870,N_15830);
xor U16054 (N_16054,N_15917,N_15778);
and U16055 (N_16055,N_15915,N_15850);
nor U16056 (N_16056,N_15758,N_15780);
and U16057 (N_16057,N_15787,N_15794);
or U16058 (N_16058,N_15985,N_15892);
xnor U16059 (N_16059,N_15847,N_15777);
nand U16060 (N_16060,N_15865,N_15751);
or U16061 (N_16061,N_15907,N_15820);
or U16062 (N_16062,N_15909,N_15864);
nand U16063 (N_16063,N_15982,N_15853);
and U16064 (N_16064,N_15860,N_15804);
or U16065 (N_16065,N_15953,N_15845);
or U16066 (N_16066,N_15936,N_15946);
and U16067 (N_16067,N_15773,N_15809);
nand U16068 (N_16068,N_15779,N_15811);
xnor U16069 (N_16069,N_15928,N_15927);
nand U16070 (N_16070,N_15854,N_15887);
or U16071 (N_16071,N_15966,N_15918);
or U16072 (N_16072,N_15775,N_15805);
nand U16073 (N_16073,N_15965,N_15803);
nor U16074 (N_16074,N_15993,N_15878);
and U16075 (N_16075,N_15945,N_15796);
nor U16076 (N_16076,N_15812,N_15838);
nor U16077 (N_16077,N_15828,N_15823);
or U16078 (N_16078,N_15881,N_15754);
nand U16079 (N_16079,N_15962,N_15960);
xor U16080 (N_16080,N_15901,N_15840);
or U16081 (N_16081,N_15884,N_15922);
or U16082 (N_16082,N_15980,N_15996);
or U16083 (N_16083,N_15934,N_15935);
xnor U16084 (N_16084,N_15798,N_15877);
and U16085 (N_16085,N_15999,N_15814);
xnor U16086 (N_16086,N_15916,N_15959);
or U16087 (N_16087,N_15949,N_15827);
nand U16088 (N_16088,N_15834,N_15842);
xor U16089 (N_16089,N_15852,N_15952);
nand U16090 (N_16090,N_15872,N_15825);
nor U16091 (N_16091,N_15968,N_15908);
nor U16092 (N_16092,N_15867,N_15776);
or U16093 (N_16093,N_15895,N_15939);
nand U16094 (N_16094,N_15839,N_15770);
xor U16095 (N_16095,N_15950,N_15752);
nand U16096 (N_16096,N_15955,N_15893);
nand U16097 (N_16097,N_15831,N_15970);
or U16098 (N_16098,N_15882,N_15990);
nor U16099 (N_16099,N_15902,N_15785);
or U16100 (N_16100,N_15795,N_15964);
nor U16101 (N_16101,N_15806,N_15863);
nor U16102 (N_16102,N_15792,N_15824);
nand U16103 (N_16103,N_15885,N_15764);
nand U16104 (N_16104,N_15941,N_15921);
nand U16105 (N_16105,N_15818,N_15972);
nor U16106 (N_16106,N_15924,N_15912);
nand U16107 (N_16107,N_15829,N_15995);
and U16108 (N_16108,N_15978,N_15954);
nand U16109 (N_16109,N_15768,N_15760);
nor U16110 (N_16110,N_15906,N_15961);
nand U16111 (N_16111,N_15861,N_15933);
nor U16112 (N_16112,N_15859,N_15899);
nor U16113 (N_16113,N_15750,N_15766);
or U16114 (N_16114,N_15948,N_15821);
nor U16115 (N_16115,N_15890,N_15886);
xor U16116 (N_16116,N_15841,N_15969);
xor U16117 (N_16117,N_15807,N_15858);
nor U16118 (N_16118,N_15967,N_15769);
xnor U16119 (N_16119,N_15817,N_15971);
nand U16120 (N_16120,N_15753,N_15873);
and U16121 (N_16121,N_15958,N_15981);
xnor U16122 (N_16122,N_15977,N_15986);
or U16123 (N_16123,N_15925,N_15772);
or U16124 (N_16124,N_15984,N_15947);
nand U16125 (N_16125,N_15899,N_15823);
or U16126 (N_16126,N_15988,N_15874);
and U16127 (N_16127,N_15794,N_15826);
nor U16128 (N_16128,N_15934,N_15890);
nand U16129 (N_16129,N_15953,N_15904);
nor U16130 (N_16130,N_15795,N_15876);
or U16131 (N_16131,N_15939,N_15817);
nand U16132 (N_16132,N_15975,N_15851);
xnor U16133 (N_16133,N_15947,N_15915);
or U16134 (N_16134,N_15790,N_15949);
or U16135 (N_16135,N_15903,N_15819);
and U16136 (N_16136,N_15874,N_15888);
and U16137 (N_16137,N_15829,N_15968);
nand U16138 (N_16138,N_15959,N_15973);
and U16139 (N_16139,N_15890,N_15833);
and U16140 (N_16140,N_15882,N_15790);
or U16141 (N_16141,N_15798,N_15925);
and U16142 (N_16142,N_15983,N_15843);
and U16143 (N_16143,N_15778,N_15876);
or U16144 (N_16144,N_15927,N_15966);
xor U16145 (N_16145,N_15880,N_15972);
nor U16146 (N_16146,N_15890,N_15922);
and U16147 (N_16147,N_15872,N_15778);
and U16148 (N_16148,N_15898,N_15951);
xor U16149 (N_16149,N_15988,N_15986);
and U16150 (N_16150,N_15891,N_15770);
or U16151 (N_16151,N_15752,N_15918);
xnor U16152 (N_16152,N_15921,N_15797);
nor U16153 (N_16153,N_15914,N_15894);
xnor U16154 (N_16154,N_15976,N_15755);
and U16155 (N_16155,N_15846,N_15809);
and U16156 (N_16156,N_15994,N_15978);
xnor U16157 (N_16157,N_15768,N_15853);
nor U16158 (N_16158,N_15856,N_15893);
or U16159 (N_16159,N_15768,N_15991);
and U16160 (N_16160,N_15981,N_15815);
or U16161 (N_16161,N_15913,N_15847);
nand U16162 (N_16162,N_15854,N_15830);
xor U16163 (N_16163,N_15781,N_15976);
xor U16164 (N_16164,N_15992,N_15855);
nor U16165 (N_16165,N_15953,N_15951);
nor U16166 (N_16166,N_15859,N_15920);
xnor U16167 (N_16167,N_15959,N_15996);
nor U16168 (N_16168,N_15828,N_15933);
nor U16169 (N_16169,N_15868,N_15977);
and U16170 (N_16170,N_15809,N_15896);
nand U16171 (N_16171,N_15905,N_15942);
and U16172 (N_16172,N_15985,N_15836);
nor U16173 (N_16173,N_15808,N_15989);
or U16174 (N_16174,N_15886,N_15779);
xnor U16175 (N_16175,N_15789,N_15757);
or U16176 (N_16176,N_15876,N_15802);
or U16177 (N_16177,N_15763,N_15778);
nand U16178 (N_16178,N_15898,N_15780);
and U16179 (N_16179,N_15914,N_15854);
nor U16180 (N_16180,N_15913,N_15998);
xor U16181 (N_16181,N_15898,N_15811);
nor U16182 (N_16182,N_15976,N_15961);
and U16183 (N_16183,N_15864,N_15868);
xnor U16184 (N_16184,N_15786,N_15785);
nor U16185 (N_16185,N_15875,N_15808);
nand U16186 (N_16186,N_15968,N_15909);
xor U16187 (N_16187,N_15863,N_15779);
and U16188 (N_16188,N_15810,N_15990);
nor U16189 (N_16189,N_15789,N_15863);
xor U16190 (N_16190,N_15993,N_15776);
xor U16191 (N_16191,N_15956,N_15846);
and U16192 (N_16192,N_15814,N_15761);
nor U16193 (N_16193,N_15912,N_15903);
nor U16194 (N_16194,N_15875,N_15869);
nand U16195 (N_16195,N_15767,N_15913);
nor U16196 (N_16196,N_15805,N_15819);
nor U16197 (N_16197,N_15979,N_15967);
nor U16198 (N_16198,N_15895,N_15926);
or U16199 (N_16199,N_15857,N_15848);
nor U16200 (N_16200,N_15995,N_15790);
xnor U16201 (N_16201,N_15883,N_15971);
or U16202 (N_16202,N_15930,N_15893);
and U16203 (N_16203,N_15900,N_15950);
nor U16204 (N_16204,N_15810,N_15837);
or U16205 (N_16205,N_15844,N_15793);
nor U16206 (N_16206,N_15922,N_15991);
nand U16207 (N_16207,N_15870,N_15838);
nand U16208 (N_16208,N_15864,N_15847);
nor U16209 (N_16209,N_15927,N_15839);
xnor U16210 (N_16210,N_15983,N_15930);
xor U16211 (N_16211,N_15999,N_15968);
or U16212 (N_16212,N_15803,N_15818);
or U16213 (N_16213,N_15954,N_15880);
nor U16214 (N_16214,N_15807,N_15835);
and U16215 (N_16215,N_15975,N_15906);
nor U16216 (N_16216,N_15957,N_15806);
and U16217 (N_16217,N_15895,N_15810);
nor U16218 (N_16218,N_15781,N_15826);
nand U16219 (N_16219,N_15780,N_15794);
or U16220 (N_16220,N_15916,N_15787);
xnor U16221 (N_16221,N_15791,N_15988);
nand U16222 (N_16222,N_15816,N_15855);
nand U16223 (N_16223,N_15896,N_15976);
nand U16224 (N_16224,N_15773,N_15796);
nand U16225 (N_16225,N_15990,N_15797);
xnor U16226 (N_16226,N_15968,N_15821);
nor U16227 (N_16227,N_15969,N_15948);
nand U16228 (N_16228,N_15903,N_15881);
nand U16229 (N_16229,N_15887,N_15781);
nor U16230 (N_16230,N_15779,N_15790);
nor U16231 (N_16231,N_15903,N_15930);
and U16232 (N_16232,N_15827,N_15777);
nor U16233 (N_16233,N_15775,N_15978);
nand U16234 (N_16234,N_15769,N_15953);
nor U16235 (N_16235,N_15981,N_15973);
nor U16236 (N_16236,N_15921,N_15967);
or U16237 (N_16237,N_15918,N_15781);
nor U16238 (N_16238,N_15755,N_15892);
or U16239 (N_16239,N_15770,N_15830);
nor U16240 (N_16240,N_15982,N_15886);
nor U16241 (N_16241,N_15951,N_15963);
nand U16242 (N_16242,N_15911,N_15961);
or U16243 (N_16243,N_15752,N_15870);
nand U16244 (N_16244,N_15914,N_15752);
or U16245 (N_16245,N_15942,N_15882);
nand U16246 (N_16246,N_15810,N_15906);
nor U16247 (N_16247,N_15792,N_15762);
nand U16248 (N_16248,N_15995,N_15893);
xnor U16249 (N_16249,N_15841,N_15893);
nand U16250 (N_16250,N_16180,N_16075);
or U16251 (N_16251,N_16245,N_16007);
nor U16252 (N_16252,N_16134,N_16239);
or U16253 (N_16253,N_16067,N_16157);
and U16254 (N_16254,N_16168,N_16128);
nand U16255 (N_16255,N_16154,N_16074);
or U16256 (N_16256,N_16191,N_16177);
nor U16257 (N_16257,N_16053,N_16217);
nand U16258 (N_16258,N_16035,N_16151);
or U16259 (N_16259,N_16167,N_16052);
nor U16260 (N_16260,N_16204,N_16008);
xnor U16261 (N_16261,N_16039,N_16083);
and U16262 (N_16262,N_16063,N_16159);
nand U16263 (N_16263,N_16044,N_16205);
or U16264 (N_16264,N_16169,N_16235);
nand U16265 (N_16265,N_16135,N_16155);
nor U16266 (N_16266,N_16006,N_16170);
xnor U16267 (N_16267,N_16133,N_16064);
or U16268 (N_16268,N_16149,N_16025);
xor U16269 (N_16269,N_16079,N_16101);
xnor U16270 (N_16270,N_16203,N_16209);
or U16271 (N_16271,N_16041,N_16090);
nor U16272 (N_16272,N_16118,N_16073);
nand U16273 (N_16273,N_16012,N_16196);
xnor U16274 (N_16274,N_16223,N_16152);
and U16275 (N_16275,N_16005,N_16032);
or U16276 (N_16276,N_16127,N_16001);
nand U16277 (N_16277,N_16094,N_16043);
xor U16278 (N_16278,N_16129,N_16026);
xor U16279 (N_16279,N_16247,N_16199);
or U16280 (N_16280,N_16059,N_16047);
nor U16281 (N_16281,N_16238,N_16153);
nor U16282 (N_16282,N_16027,N_16119);
nand U16283 (N_16283,N_16104,N_16172);
and U16284 (N_16284,N_16046,N_16194);
nor U16285 (N_16285,N_16219,N_16181);
or U16286 (N_16286,N_16056,N_16077);
nand U16287 (N_16287,N_16086,N_16085);
or U16288 (N_16288,N_16050,N_16174);
nor U16289 (N_16289,N_16145,N_16193);
or U16290 (N_16290,N_16054,N_16106);
and U16291 (N_16291,N_16200,N_16233);
or U16292 (N_16292,N_16211,N_16066);
nand U16293 (N_16293,N_16158,N_16126);
nand U16294 (N_16294,N_16092,N_16031);
and U16295 (N_16295,N_16117,N_16049);
xor U16296 (N_16296,N_16100,N_16230);
xnor U16297 (N_16297,N_16163,N_16232);
nor U16298 (N_16298,N_16014,N_16003);
xor U16299 (N_16299,N_16183,N_16173);
or U16300 (N_16300,N_16021,N_16146);
xor U16301 (N_16301,N_16091,N_16150);
xnor U16302 (N_16302,N_16078,N_16201);
xnor U16303 (N_16303,N_16057,N_16162);
xor U16304 (N_16304,N_16103,N_16136);
xor U16305 (N_16305,N_16130,N_16186);
nand U16306 (N_16306,N_16055,N_16185);
and U16307 (N_16307,N_16215,N_16143);
nor U16308 (N_16308,N_16022,N_16024);
nor U16309 (N_16309,N_16188,N_16226);
nand U16310 (N_16310,N_16089,N_16213);
nand U16311 (N_16311,N_16147,N_16198);
nand U16312 (N_16312,N_16176,N_16069);
xor U16313 (N_16313,N_16248,N_16095);
or U16314 (N_16314,N_16192,N_16034);
nor U16315 (N_16315,N_16225,N_16029);
nor U16316 (N_16316,N_16112,N_16244);
nand U16317 (N_16317,N_16033,N_16190);
and U16318 (N_16318,N_16220,N_16023);
nand U16319 (N_16319,N_16137,N_16108);
nor U16320 (N_16320,N_16000,N_16017);
or U16321 (N_16321,N_16207,N_16102);
xnor U16322 (N_16322,N_16110,N_16165);
or U16323 (N_16323,N_16124,N_16087);
nand U16324 (N_16324,N_16002,N_16060);
nor U16325 (N_16325,N_16015,N_16098);
xor U16326 (N_16326,N_16148,N_16122);
nand U16327 (N_16327,N_16229,N_16184);
nand U16328 (N_16328,N_16004,N_16156);
xnor U16329 (N_16329,N_16140,N_16061);
nand U16330 (N_16330,N_16097,N_16038);
xnor U16331 (N_16331,N_16120,N_16195);
nand U16332 (N_16332,N_16231,N_16093);
xor U16333 (N_16333,N_16020,N_16121);
nor U16334 (N_16334,N_16171,N_16018);
xnor U16335 (N_16335,N_16111,N_16212);
nand U16336 (N_16336,N_16142,N_16218);
or U16337 (N_16337,N_16189,N_16082);
xnor U16338 (N_16338,N_16125,N_16010);
and U16339 (N_16339,N_16115,N_16206);
xor U16340 (N_16340,N_16243,N_16227);
or U16341 (N_16341,N_16197,N_16081);
and U16342 (N_16342,N_16070,N_16048);
nand U16343 (N_16343,N_16065,N_16076);
or U16344 (N_16344,N_16062,N_16222);
nor U16345 (N_16345,N_16210,N_16242);
nand U16346 (N_16346,N_16249,N_16028);
and U16347 (N_16347,N_16088,N_16036);
xnor U16348 (N_16348,N_16161,N_16221);
xor U16349 (N_16349,N_16164,N_16160);
nand U16350 (N_16350,N_16224,N_16013);
or U16351 (N_16351,N_16109,N_16116);
and U16352 (N_16352,N_16175,N_16037);
or U16353 (N_16353,N_16009,N_16234);
and U16354 (N_16354,N_16246,N_16179);
nor U16355 (N_16355,N_16045,N_16241);
and U16356 (N_16356,N_16071,N_16019);
or U16357 (N_16357,N_16113,N_16011);
and U16358 (N_16358,N_16138,N_16107);
and U16359 (N_16359,N_16240,N_16096);
and U16360 (N_16360,N_16123,N_16068);
nand U16361 (N_16361,N_16141,N_16216);
nor U16362 (N_16362,N_16237,N_16099);
nor U16363 (N_16363,N_16139,N_16058);
or U16364 (N_16364,N_16166,N_16072);
nand U16365 (N_16365,N_16178,N_16187);
nor U16366 (N_16366,N_16114,N_16042);
or U16367 (N_16367,N_16144,N_16030);
xnor U16368 (N_16368,N_16202,N_16040);
xor U16369 (N_16369,N_16236,N_16105);
nand U16370 (N_16370,N_16080,N_16084);
nand U16371 (N_16371,N_16051,N_16208);
xor U16372 (N_16372,N_16131,N_16228);
and U16373 (N_16373,N_16214,N_16132);
and U16374 (N_16374,N_16182,N_16016);
and U16375 (N_16375,N_16190,N_16148);
nand U16376 (N_16376,N_16035,N_16198);
nand U16377 (N_16377,N_16096,N_16095);
nor U16378 (N_16378,N_16097,N_16123);
nand U16379 (N_16379,N_16157,N_16158);
or U16380 (N_16380,N_16245,N_16004);
xnor U16381 (N_16381,N_16146,N_16205);
xnor U16382 (N_16382,N_16244,N_16154);
or U16383 (N_16383,N_16051,N_16137);
and U16384 (N_16384,N_16053,N_16185);
xor U16385 (N_16385,N_16172,N_16015);
nor U16386 (N_16386,N_16096,N_16046);
nand U16387 (N_16387,N_16144,N_16050);
xnor U16388 (N_16388,N_16192,N_16035);
nand U16389 (N_16389,N_16092,N_16152);
or U16390 (N_16390,N_16009,N_16157);
or U16391 (N_16391,N_16247,N_16210);
xor U16392 (N_16392,N_16117,N_16156);
nor U16393 (N_16393,N_16134,N_16103);
and U16394 (N_16394,N_16162,N_16198);
nor U16395 (N_16395,N_16092,N_16190);
and U16396 (N_16396,N_16193,N_16089);
and U16397 (N_16397,N_16140,N_16226);
or U16398 (N_16398,N_16194,N_16202);
xor U16399 (N_16399,N_16031,N_16244);
and U16400 (N_16400,N_16011,N_16208);
nand U16401 (N_16401,N_16139,N_16186);
and U16402 (N_16402,N_16199,N_16032);
xor U16403 (N_16403,N_16100,N_16048);
nor U16404 (N_16404,N_16234,N_16237);
or U16405 (N_16405,N_16098,N_16151);
and U16406 (N_16406,N_16208,N_16120);
nor U16407 (N_16407,N_16024,N_16149);
or U16408 (N_16408,N_16043,N_16064);
nor U16409 (N_16409,N_16207,N_16114);
nand U16410 (N_16410,N_16209,N_16012);
or U16411 (N_16411,N_16027,N_16183);
and U16412 (N_16412,N_16064,N_16231);
or U16413 (N_16413,N_16081,N_16199);
xor U16414 (N_16414,N_16000,N_16103);
and U16415 (N_16415,N_16072,N_16187);
xor U16416 (N_16416,N_16010,N_16088);
and U16417 (N_16417,N_16086,N_16161);
nand U16418 (N_16418,N_16101,N_16009);
nor U16419 (N_16419,N_16185,N_16156);
or U16420 (N_16420,N_16003,N_16212);
xnor U16421 (N_16421,N_16039,N_16239);
xor U16422 (N_16422,N_16036,N_16097);
or U16423 (N_16423,N_16072,N_16191);
nand U16424 (N_16424,N_16086,N_16000);
and U16425 (N_16425,N_16078,N_16089);
xnor U16426 (N_16426,N_16208,N_16127);
and U16427 (N_16427,N_16076,N_16213);
or U16428 (N_16428,N_16129,N_16095);
and U16429 (N_16429,N_16126,N_16042);
or U16430 (N_16430,N_16063,N_16216);
and U16431 (N_16431,N_16241,N_16076);
nor U16432 (N_16432,N_16110,N_16198);
nor U16433 (N_16433,N_16177,N_16101);
and U16434 (N_16434,N_16103,N_16119);
nand U16435 (N_16435,N_16096,N_16154);
nand U16436 (N_16436,N_16072,N_16111);
nor U16437 (N_16437,N_16092,N_16213);
xor U16438 (N_16438,N_16055,N_16024);
and U16439 (N_16439,N_16158,N_16085);
nand U16440 (N_16440,N_16117,N_16016);
xnor U16441 (N_16441,N_16092,N_16047);
xor U16442 (N_16442,N_16194,N_16198);
nor U16443 (N_16443,N_16048,N_16208);
nand U16444 (N_16444,N_16035,N_16211);
and U16445 (N_16445,N_16191,N_16194);
and U16446 (N_16446,N_16245,N_16195);
or U16447 (N_16447,N_16197,N_16209);
nand U16448 (N_16448,N_16224,N_16229);
nand U16449 (N_16449,N_16009,N_16058);
or U16450 (N_16450,N_16242,N_16167);
and U16451 (N_16451,N_16114,N_16132);
nor U16452 (N_16452,N_16147,N_16195);
and U16453 (N_16453,N_16219,N_16195);
and U16454 (N_16454,N_16083,N_16182);
and U16455 (N_16455,N_16208,N_16010);
nor U16456 (N_16456,N_16192,N_16204);
or U16457 (N_16457,N_16037,N_16001);
xnor U16458 (N_16458,N_16189,N_16106);
or U16459 (N_16459,N_16144,N_16227);
and U16460 (N_16460,N_16227,N_16103);
nand U16461 (N_16461,N_16154,N_16050);
nor U16462 (N_16462,N_16065,N_16043);
nor U16463 (N_16463,N_16217,N_16044);
nand U16464 (N_16464,N_16126,N_16108);
nand U16465 (N_16465,N_16222,N_16003);
or U16466 (N_16466,N_16129,N_16066);
or U16467 (N_16467,N_16212,N_16175);
or U16468 (N_16468,N_16153,N_16052);
and U16469 (N_16469,N_16198,N_16091);
and U16470 (N_16470,N_16135,N_16184);
or U16471 (N_16471,N_16248,N_16242);
or U16472 (N_16472,N_16126,N_16111);
and U16473 (N_16473,N_16147,N_16174);
nand U16474 (N_16474,N_16056,N_16060);
nand U16475 (N_16475,N_16109,N_16044);
and U16476 (N_16476,N_16165,N_16034);
xnor U16477 (N_16477,N_16088,N_16039);
or U16478 (N_16478,N_16068,N_16141);
nor U16479 (N_16479,N_16138,N_16208);
and U16480 (N_16480,N_16131,N_16042);
nor U16481 (N_16481,N_16145,N_16245);
or U16482 (N_16482,N_16027,N_16058);
xnor U16483 (N_16483,N_16205,N_16077);
xnor U16484 (N_16484,N_16229,N_16043);
xnor U16485 (N_16485,N_16026,N_16099);
xor U16486 (N_16486,N_16057,N_16061);
nand U16487 (N_16487,N_16028,N_16072);
and U16488 (N_16488,N_16003,N_16112);
nand U16489 (N_16489,N_16158,N_16180);
nor U16490 (N_16490,N_16082,N_16170);
nor U16491 (N_16491,N_16226,N_16183);
or U16492 (N_16492,N_16085,N_16056);
or U16493 (N_16493,N_16014,N_16110);
nand U16494 (N_16494,N_16059,N_16188);
xor U16495 (N_16495,N_16120,N_16231);
and U16496 (N_16496,N_16208,N_16211);
xor U16497 (N_16497,N_16207,N_16178);
and U16498 (N_16498,N_16038,N_16238);
xnor U16499 (N_16499,N_16056,N_16097);
nand U16500 (N_16500,N_16299,N_16296);
nor U16501 (N_16501,N_16267,N_16498);
nand U16502 (N_16502,N_16282,N_16405);
xnor U16503 (N_16503,N_16321,N_16389);
nor U16504 (N_16504,N_16420,N_16312);
and U16505 (N_16505,N_16487,N_16399);
nor U16506 (N_16506,N_16464,N_16271);
nand U16507 (N_16507,N_16477,N_16258);
nand U16508 (N_16508,N_16264,N_16485);
xor U16509 (N_16509,N_16377,N_16311);
nor U16510 (N_16510,N_16346,N_16251);
nor U16511 (N_16511,N_16426,N_16491);
and U16512 (N_16512,N_16370,N_16497);
nor U16513 (N_16513,N_16330,N_16445);
xor U16514 (N_16514,N_16383,N_16489);
or U16515 (N_16515,N_16417,N_16373);
or U16516 (N_16516,N_16462,N_16252);
or U16517 (N_16517,N_16371,N_16364);
or U16518 (N_16518,N_16331,N_16307);
nor U16519 (N_16519,N_16463,N_16414);
or U16520 (N_16520,N_16315,N_16273);
nor U16521 (N_16521,N_16297,N_16400);
or U16522 (N_16522,N_16265,N_16272);
and U16523 (N_16523,N_16332,N_16355);
xor U16524 (N_16524,N_16286,N_16460);
nand U16525 (N_16525,N_16365,N_16304);
and U16526 (N_16526,N_16479,N_16260);
xor U16527 (N_16527,N_16368,N_16404);
or U16528 (N_16528,N_16429,N_16397);
and U16529 (N_16529,N_16480,N_16356);
and U16530 (N_16530,N_16478,N_16372);
or U16531 (N_16531,N_16309,N_16366);
xnor U16532 (N_16532,N_16352,N_16442);
nor U16533 (N_16533,N_16452,N_16351);
nand U16534 (N_16534,N_16493,N_16348);
nand U16535 (N_16535,N_16430,N_16283);
and U16536 (N_16536,N_16499,N_16415);
nand U16537 (N_16537,N_16341,N_16257);
nand U16538 (N_16538,N_16256,N_16329);
and U16539 (N_16539,N_16450,N_16278);
or U16540 (N_16540,N_16424,N_16314);
and U16541 (N_16541,N_16443,N_16350);
or U16542 (N_16542,N_16380,N_16461);
nor U16543 (N_16543,N_16320,N_16421);
and U16544 (N_16544,N_16358,N_16482);
xnor U16545 (N_16545,N_16467,N_16333);
nand U16546 (N_16546,N_16472,N_16281);
nor U16547 (N_16547,N_16268,N_16255);
nor U16548 (N_16548,N_16416,N_16409);
and U16549 (N_16549,N_16492,N_16446);
and U16550 (N_16550,N_16342,N_16301);
or U16551 (N_16551,N_16406,N_16340);
or U16552 (N_16552,N_16395,N_16471);
nand U16553 (N_16553,N_16481,N_16306);
nor U16554 (N_16554,N_16363,N_16486);
or U16555 (N_16555,N_16328,N_16376);
or U16556 (N_16556,N_16305,N_16466);
nor U16557 (N_16557,N_16313,N_16387);
xnor U16558 (N_16558,N_16474,N_16495);
nand U16559 (N_16559,N_16441,N_16419);
nor U16560 (N_16560,N_16459,N_16308);
xor U16561 (N_16561,N_16411,N_16469);
nor U16562 (N_16562,N_16334,N_16490);
and U16563 (N_16563,N_16434,N_16488);
nor U16564 (N_16564,N_16293,N_16440);
nand U16565 (N_16565,N_16401,N_16322);
and U16566 (N_16566,N_16349,N_16367);
nand U16567 (N_16567,N_16285,N_16473);
and U16568 (N_16568,N_16270,N_16403);
xnor U16569 (N_16569,N_16448,N_16253);
nor U16570 (N_16570,N_16337,N_16276);
xor U16571 (N_16571,N_16274,N_16475);
xor U16572 (N_16572,N_16410,N_16344);
or U16573 (N_16573,N_16303,N_16468);
and U16574 (N_16574,N_16439,N_16433);
nand U16575 (N_16575,N_16375,N_16269);
xnor U16576 (N_16576,N_16392,N_16318);
nand U16577 (N_16577,N_16388,N_16338);
and U16578 (N_16578,N_16279,N_16284);
xor U16579 (N_16579,N_16263,N_16451);
and U16580 (N_16580,N_16390,N_16412);
nor U16581 (N_16581,N_16425,N_16295);
and U16582 (N_16582,N_16394,N_16413);
and U16583 (N_16583,N_16277,N_16353);
and U16584 (N_16584,N_16302,N_16465);
and U16585 (N_16585,N_16250,N_16418);
nor U16586 (N_16586,N_16391,N_16432);
or U16587 (N_16587,N_16339,N_16453);
or U16588 (N_16588,N_16261,N_16357);
nor U16589 (N_16589,N_16436,N_16325);
nor U16590 (N_16590,N_16379,N_16292);
nand U16591 (N_16591,N_16431,N_16288);
xnor U16592 (N_16592,N_16361,N_16290);
nand U16593 (N_16593,N_16326,N_16362);
or U16594 (N_16594,N_16347,N_16407);
nor U16595 (N_16595,N_16384,N_16262);
or U16596 (N_16596,N_16275,N_16359);
nand U16597 (N_16597,N_16393,N_16343);
nand U16598 (N_16598,N_16335,N_16327);
nor U16599 (N_16599,N_16457,N_16437);
or U16600 (N_16600,N_16438,N_16402);
and U16601 (N_16601,N_16259,N_16444);
xnor U16602 (N_16602,N_16494,N_16317);
and U16603 (N_16603,N_16374,N_16449);
and U16604 (N_16604,N_16408,N_16447);
or U16605 (N_16605,N_16280,N_16354);
nor U16606 (N_16606,N_16254,N_16336);
nand U16607 (N_16607,N_16323,N_16287);
or U16608 (N_16608,N_16324,N_16427);
nor U16609 (N_16609,N_16294,N_16300);
nor U16610 (N_16610,N_16423,N_16470);
or U16611 (N_16611,N_16496,N_16454);
nor U16612 (N_16612,N_16382,N_16291);
nand U16613 (N_16613,N_16458,N_16381);
nor U16614 (N_16614,N_16316,N_16396);
nor U16615 (N_16615,N_16484,N_16476);
xor U16616 (N_16616,N_16298,N_16422);
and U16617 (N_16617,N_16385,N_16378);
and U16618 (N_16618,N_16266,N_16398);
nor U16619 (N_16619,N_16289,N_16360);
or U16620 (N_16620,N_16386,N_16435);
or U16621 (N_16621,N_16455,N_16310);
xnor U16622 (N_16622,N_16369,N_16483);
and U16623 (N_16623,N_16456,N_16345);
and U16624 (N_16624,N_16428,N_16319);
and U16625 (N_16625,N_16267,N_16375);
and U16626 (N_16626,N_16313,N_16331);
nand U16627 (N_16627,N_16288,N_16470);
and U16628 (N_16628,N_16407,N_16377);
and U16629 (N_16629,N_16445,N_16297);
or U16630 (N_16630,N_16440,N_16478);
xnor U16631 (N_16631,N_16336,N_16261);
nand U16632 (N_16632,N_16386,N_16252);
and U16633 (N_16633,N_16279,N_16322);
and U16634 (N_16634,N_16480,N_16359);
nand U16635 (N_16635,N_16297,N_16484);
xor U16636 (N_16636,N_16438,N_16433);
xor U16637 (N_16637,N_16269,N_16336);
or U16638 (N_16638,N_16306,N_16276);
nand U16639 (N_16639,N_16480,N_16284);
and U16640 (N_16640,N_16414,N_16496);
or U16641 (N_16641,N_16419,N_16432);
and U16642 (N_16642,N_16426,N_16264);
nand U16643 (N_16643,N_16331,N_16301);
nor U16644 (N_16644,N_16396,N_16394);
nor U16645 (N_16645,N_16396,N_16385);
nand U16646 (N_16646,N_16425,N_16251);
nand U16647 (N_16647,N_16314,N_16255);
and U16648 (N_16648,N_16467,N_16444);
nor U16649 (N_16649,N_16443,N_16373);
or U16650 (N_16650,N_16439,N_16470);
nor U16651 (N_16651,N_16384,N_16254);
xnor U16652 (N_16652,N_16376,N_16264);
nor U16653 (N_16653,N_16313,N_16356);
nand U16654 (N_16654,N_16336,N_16485);
and U16655 (N_16655,N_16253,N_16347);
xor U16656 (N_16656,N_16442,N_16356);
and U16657 (N_16657,N_16331,N_16327);
or U16658 (N_16658,N_16404,N_16284);
and U16659 (N_16659,N_16413,N_16440);
xnor U16660 (N_16660,N_16338,N_16251);
and U16661 (N_16661,N_16476,N_16378);
and U16662 (N_16662,N_16439,N_16446);
nor U16663 (N_16663,N_16286,N_16429);
and U16664 (N_16664,N_16419,N_16277);
nor U16665 (N_16665,N_16419,N_16331);
xor U16666 (N_16666,N_16466,N_16256);
and U16667 (N_16667,N_16324,N_16371);
xnor U16668 (N_16668,N_16298,N_16467);
or U16669 (N_16669,N_16451,N_16409);
xor U16670 (N_16670,N_16389,N_16455);
xnor U16671 (N_16671,N_16296,N_16390);
nor U16672 (N_16672,N_16377,N_16344);
xor U16673 (N_16673,N_16480,N_16408);
nand U16674 (N_16674,N_16453,N_16410);
nand U16675 (N_16675,N_16464,N_16493);
and U16676 (N_16676,N_16260,N_16265);
nor U16677 (N_16677,N_16475,N_16398);
and U16678 (N_16678,N_16436,N_16271);
and U16679 (N_16679,N_16402,N_16487);
or U16680 (N_16680,N_16495,N_16266);
and U16681 (N_16681,N_16425,N_16335);
and U16682 (N_16682,N_16308,N_16316);
nor U16683 (N_16683,N_16372,N_16288);
nand U16684 (N_16684,N_16408,N_16383);
nor U16685 (N_16685,N_16362,N_16409);
nand U16686 (N_16686,N_16278,N_16302);
nand U16687 (N_16687,N_16445,N_16423);
nor U16688 (N_16688,N_16267,N_16265);
or U16689 (N_16689,N_16373,N_16352);
nand U16690 (N_16690,N_16292,N_16348);
xor U16691 (N_16691,N_16296,N_16256);
xnor U16692 (N_16692,N_16267,N_16272);
and U16693 (N_16693,N_16471,N_16301);
xor U16694 (N_16694,N_16467,N_16440);
nor U16695 (N_16695,N_16355,N_16399);
nor U16696 (N_16696,N_16423,N_16382);
and U16697 (N_16697,N_16280,N_16375);
nand U16698 (N_16698,N_16310,N_16302);
nand U16699 (N_16699,N_16353,N_16342);
and U16700 (N_16700,N_16418,N_16284);
nand U16701 (N_16701,N_16381,N_16418);
or U16702 (N_16702,N_16398,N_16466);
nand U16703 (N_16703,N_16389,N_16275);
and U16704 (N_16704,N_16418,N_16290);
nand U16705 (N_16705,N_16374,N_16394);
xor U16706 (N_16706,N_16435,N_16394);
nand U16707 (N_16707,N_16278,N_16482);
and U16708 (N_16708,N_16349,N_16476);
xnor U16709 (N_16709,N_16444,N_16429);
and U16710 (N_16710,N_16356,N_16254);
nor U16711 (N_16711,N_16493,N_16346);
nor U16712 (N_16712,N_16410,N_16279);
nor U16713 (N_16713,N_16446,N_16389);
xor U16714 (N_16714,N_16419,N_16309);
nand U16715 (N_16715,N_16426,N_16342);
and U16716 (N_16716,N_16276,N_16457);
xor U16717 (N_16717,N_16362,N_16327);
or U16718 (N_16718,N_16459,N_16406);
nor U16719 (N_16719,N_16378,N_16414);
nand U16720 (N_16720,N_16401,N_16472);
and U16721 (N_16721,N_16440,N_16302);
and U16722 (N_16722,N_16429,N_16298);
and U16723 (N_16723,N_16267,N_16280);
or U16724 (N_16724,N_16294,N_16270);
nand U16725 (N_16725,N_16388,N_16418);
or U16726 (N_16726,N_16330,N_16328);
or U16727 (N_16727,N_16276,N_16415);
nand U16728 (N_16728,N_16260,N_16306);
and U16729 (N_16729,N_16468,N_16251);
xnor U16730 (N_16730,N_16485,N_16377);
xor U16731 (N_16731,N_16478,N_16477);
nand U16732 (N_16732,N_16472,N_16360);
nand U16733 (N_16733,N_16345,N_16359);
xnor U16734 (N_16734,N_16310,N_16458);
and U16735 (N_16735,N_16258,N_16275);
xnor U16736 (N_16736,N_16436,N_16279);
xor U16737 (N_16737,N_16321,N_16359);
or U16738 (N_16738,N_16304,N_16293);
nor U16739 (N_16739,N_16345,N_16305);
or U16740 (N_16740,N_16305,N_16357);
nor U16741 (N_16741,N_16468,N_16329);
nor U16742 (N_16742,N_16410,N_16415);
xor U16743 (N_16743,N_16469,N_16471);
nand U16744 (N_16744,N_16460,N_16459);
nand U16745 (N_16745,N_16413,N_16268);
and U16746 (N_16746,N_16361,N_16471);
xor U16747 (N_16747,N_16278,N_16416);
xnor U16748 (N_16748,N_16428,N_16483);
or U16749 (N_16749,N_16294,N_16381);
and U16750 (N_16750,N_16656,N_16512);
and U16751 (N_16751,N_16736,N_16623);
xor U16752 (N_16752,N_16675,N_16583);
nor U16753 (N_16753,N_16710,N_16741);
and U16754 (N_16754,N_16637,N_16638);
xnor U16755 (N_16755,N_16517,N_16700);
nand U16756 (N_16756,N_16545,N_16649);
and U16757 (N_16757,N_16734,N_16686);
xnor U16758 (N_16758,N_16664,N_16746);
xor U16759 (N_16759,N_16670,N_16588);
or U16760 (N_16760,N_16546,N_16612);
nand U16761 (N_16761,N_16504,N_16552);
and U16762 (N_16762,N_16555,N_16599);
or U16763 (N_16763,N_16674,N_16594);
nor U16764 (N_16764,N_16541,N_16662);
nor U16765 (N_16765,N_16596,N_16543);
or U16766 (N_16766,N_16742,N_16591);
or U16767 (N_16767,N_16696,N_16506);
nor U16768 (N_16768,N_16635,N_16622);
and U16769 (N_16769,N_16733,N_16522);
or U16770 (N_16770,N_16628,N_16540);
nor U16771 (N_16771,N_16502,N_16681);
or U16772 (N_16772,N_16557,N_16705);
nor U16773 (N_16773,N_16711,N_16568);
xor U16774 (N_16774,N_16747,N_16523);
nor U16775 (N_16775,N_16740,N_16593);
nor U16776 (N_16776,N_16515,N_16665);
nand U16777 (N_16777,N_16693,N_16634);
and U16778 (N_16778,N_16717,N_16718);
xnor U16779 (N_16779,N_16640,N_16566);
or U16780 (N_16780,N_16531,N_16564);
and U16781 (N_16781,N_16587,N_16537);
and U16782 (N_16782,N_16703,N_16626);
and U16783 (N_16783,N_16613,N_16639);
nor U16784 (N_16784,N_16614,N_16646);
or U16785 (N_16785,N_16644,N_16726);
or U16786 (N_16786,N_16544,N_16676);
and U16787 (N_16787,N_16709,N_16679);
and U16788 (N_16788,N_16601,N_16688);
and U16789 (N_16789,N_16536,N_16682);
xor U16790 (N_16790,N_16684,N_16694);
or U16791 (N_16791,N_16739,N_16632);
and U16792 (N_16792,N_16652,N_16542);
or U16793 (N_16793,N_16500,N_16749);
nand U16794 (N_16794,N_16650,N_16658);
nand U16795 (N_16795,N_16589,N_16559);
and U16796 (N_16796,N_16534,N_16680);
nand U16797 (N_16797,N_16714,N_16524);
xnor U16798 (N_16798,N_16701,N_16704);
xnor U16799 (N_16799,N_16551,N_16556);
nor U16800 (N_16800,N_16657,N_16526);
xnor U16801 (N_16801,N_16720,N_16732);
nor U16802 (N_16802,N_16737,N_16745);
nor U16803 (N_16803,N_16519,N_16610);
or U16804 (N_16804,N_16511,N_16507);
nor U16805 (N_16805,N_16663,N_16629);
nand U16806 (N_16806,N_16707,N_16532);
or U16807 (N_16807,N_16672,N_16579);
or U16808 (N_16808,N_16516,N_16563);
and U16809 (N_16809,N_16595,N_16721);
nand U16810 (N_16810,N_16631,N_16648);
xnor U16811 (N_16811,N_16748,N_16645);
and U16812 (N_16812,N_16607,N_16633);
or U16813 (N_16813,N_16730,N_16597);
or U16814 (N_16814,N_16509,N_16520);
nand U16815 (N_16815,N_16636,N_16529);
xnor U16816 (N_16816,N_16689,N_16659);
and U16817 (N_16817,N_16510,N_16653);
xor U16818 (N_16818,N_16615,N_16548);
and U16819 (N_16819,N_16617,N_16698);
xor U16820 (N_16820,N_16738,N_16687);
and U16821 (N_16821,N_16678,N_16619);
and U16822 (N_16822,N_16525,N_16729);
and U16823 (N_16823,N_16569,N_16582);
nand U16824 (N_16824,N_16744,N_16618);
xnor U16825 (N_16825,N_16671,N_16581);
nor U16826 (N_16826,N_16604,N_16553);
or U16827 (N_16827,N_16501,N_16685);
nor U16828 (N_16828,N_16735,N_16575);
nand U16829 (N_16829,N_16630,N_16702);
nor U16830 (N_16830,N_16655,N_16592);
nand U16831 (N_16831,N_16605,N_16625);
or U16832 (N_16832,N_16586,N_16715);
xnor U16833 (N_16833,N_16570,N_16716);
nor U16834 (N_16834,N_16609,N_16533);
nand U16835 (N_16835,N_16620,N_16725);
xor U16836 (N_16836,N_16578,N_16571);
nor U16837 (N_16837,N_16673,N_16724);
and U16838 (N_16838,N_16691,N_16572);
or U16839 (N_16839,N_16505,N_16728);
nor U16840 (N_16840,N_16527,N_16647);
nor U16841 (N_16841,N_16641,N_16577);
or U16842 (N_16842,N_16549,N_16667);
xor U16843 (N_16843,N_16683,N_16666);
or U16844 (N_16844,N_16567,N_16690);
xnor U16845 (N_16845,N_16606,N_16616);
or U16846 (N_16846,N_16603,N_16651);
xor U16847 (N_16847,N_16550,N_16621);
nand U16848 (N_16848,N_16598,N_16743);
or U16849 (N_16849,N_16660,N_16514);
nand U16850 (N_16850,N_16697,N_16654);
xnor U16851 (N_16851,N_16576,N_16668);
nor U16852 (N_16852,N_16590,N_16706);
xor U16853 (N_16853,N_16602,N_16627);
and U16854 (N_16854,N_16530,N_16503);
xnor U16855 (N_16855,N_16513,N_16538);
xnor U16856 (N_16856,N_16580,N_16677);
nand U16857 (N_16857,N_16560,N_16562);
xnor U16858 (N_16858,N_16508,N_16669);
nand U16859 (N_16859,N_16584,N_16528);
or U16860 (N_16860,N_16731,N_16692);
nand U16861 (N_16861,N_16722,N_16642);
and U16862 (N_16862,N_16727,N_16535);
or U16863 (N_16863,N_16719,N_16518);
xnor U16864 (N_16864,N_16723,N_16708);
xor U16865 (N_16865,N_16611,N_16521);
or U16866 (N_16866,N_16643,N_16608);
nand U16867 (N_16867,N_16712,N_16561);
or U16868 (N_16868,N_16624,N_16558);
xnor U16869 (N_16869,N_16600,N_16695);
xor U16870 (N_16870,N_16554,N_16547);
and U16871 (N_16871,N_16585,N_16713);
xnor U16872 (N_16872,N_16661,N_16565);
and U16873 (N_16873,N_16574,N_16573);
and U16874 (N_16874,N_16539,N_16699);
nand U16875 (N_16875,N_16641,N_16722);
and U16876 (N_16876,N_16556,N_16588);
and U16877 (N_16877,N_16570,N_16680);
nand U16878 (N_16878,N_16669,N_16671);
nor U16879 (N_16879,N_16550,N_16666);
and U16880 (N_16880,N_16677,N_16527);
nor U16881 (N_16881,N_16691,N_16650);
xor U16882 (N_16882,N_16672,N_16742);
or U16883 (N_16883,N_16611,N_16511);
xnor U16884 (N_16884,N_16714,N_16745);
nor U16885 (N_16885,N_16701,N_16626);
nand U16886 (N_16886,N_16697,N_16624);
nand U16887 (N_16887,N_16692,N_16661);
xnor U16888 (N_16888,N_16735,N_16705);
xnor U16889 (N_16889,N_16502,N_16503);
and U16890 (N_16890,N_16727,N_16519);
nor U16891 (N_16891,N_16663,N_16678);
and U16892 (N_16892,N_16539,N_16540);
and U16893 (N_16893,N_16526,N_16729);
nand U16894 (N_16894,N_16547,N_16679);
or U16895 (N_16895,N_16560,N_16637);
or U16896 (N_16896,N_16522,N_16528);
or U16897 (N_16897,N_16534,N_16707);
nor U16898 (N_16898,N_16509,N_16567);
and U16899 (N_16899,N_16538,N_16739);
and U16900 (N_16900,N_16692,N_16606);
and U16901 (N_16901,N_16648,N_16614);
and U16902 (N_16902,N_16648,N_16626);
and U16903 (N_16903,N_16572,N_16513);
or U16904 (N_16904,N_16518,N_16545);
nand U16905 (N_16905,N_16635,N_16667);
xor U16906 (N_16906,N_16597,N_16679);
xnor U16907 (N_16907,N_16653,N_16589);
xnor U16908 (N_16908,N_16536,N_16718);
nand U16909 (N_16909,N_16700,N_16530);
nor U16910 (N_16910,N_16505,N_16577);
and U16911 (N_16911,N_16674,N_16511);
nand U16912 (N_16912,N_16549,N_16581);
and U16913 (N_16913,N_16576,N_16611);
and U16914 (N_16914,N_16533,N_16584);
nand U16915 (N_16915,N_16554,N_16530);
or U16916 (N_16916,N_16591,N_16608);
nor U16917 (N_16917,N_16555,N_16529);
or U16918 (N_16918,N_16599,N_16629);
or U16919 (N_16919,N_16711,N_16650);
nor U16920 (N_16920,N_16564,N_16517);
nand U16921 (N_16921,N_16648,N_16586);
and U16922 (N_16922,N_16649,N_16604);
and U16923 (N_16923,N_16547,N_16677);
nor U16924 (N_16924,N_16708,N_16728);
or U16925 (N_16925,N_16601,N_16538);
nor U16926 (N_16926,N_16658,N_16522);
or U16927 (N_16927,N_16575,N_16520);
nand U16928 (N_16928,N_16583,N_16551);
nand U16929 (N_16929,N_16640,N_16715);
xnor U16930 (N_16930,N_16557,N_16742);
nand U16931 (N_16931,N_16649,N_16500);
nand U16932 (N_16932,N_16698,N_16620);
xor U16933 (N_16933,N_16740,N_16728);
xor U16934 (N_16934,N_16733,N_16623);
nor U16935 (N_16935,N_16717,N_16517);
and U16936 (N_16936,N_16572,N_16721);
nor U16937 (N_16937,N_16639,N_16533);
nor U16938 (N_16938,N_16614,N_16697);
nand U16939 (N_16939,N_16567,N_16626);
nor U16940 (N_16940,N_16581,N_16521);
nand U16941 (N_16941,N_16691,N_16705);
and U16942 (N_16942,N_16642,N_16525);
nor U16943 (N_16943,N_16511,N_16612);
and U16944 (N_16944,N_16744,N_16514);
nand U16945 (N_16945,N_16539,N_16563);
and U16946 (N_16946,N_16611,N_16585);
xor U16947 (N_16947,N_16694,N_16685);
xnor U16948 (N_16948,N_16548,N_16643);
and U16949 (N_16949,N_16530,N_16734);
nor U16950 (N_16950,N_16528,N_16730);
nor U16951 (N_16951,N_16724,N_16567);
and U16952 (N_16952,N_16642,N_16698);
xnor U16953 (N_16953,N_16721,N_16674);
xnor U16954 (N_16954,N_16628,N_16527);
nor U16955 (N_16955,N_16720,N_16581);
xor U16956 (N_16956,N_16532,N_16653);
nand U16957 (N_16957,N_16530,N_16505);
or U16958 (N_16958,N_16614,N_16514);
and U16959 (N_16959,N_16719,N_16520);
or U16960 (N_16960,N_16539,N_16709);
xor U16961 (N_16961,N_16694,N_16547);
nor U16962 (N_16962,N_16686,N_16641);
nand U16963 (N_16963,N_16547,N_16523);
nand U16964 (N_16964,N_16733,N_16655);
or U16965 (N_16965,N_16592,N_16748);
xnor U16966 (N_16966,N_16628,N_16533);
and U16967 (N_16967,N_16636,N_16542);
and U16968 (N_16968,N_16711,N_16635);
and U16969 (N_16969,N_16681,N_16699);
xor U16970 (N_16970,N_16620,N_16570);
nor U16971 (N_16971,N_16520,N_16678);
xor U16972 (N_16972,N_16541,N_16575);
and U16973 (N_16973,N_16691,N_16660);
xor U16974 (N_16974,N_16714,N_16605);
nor U16975 (N_16975,N_16644,N_16524);
or U16976 (N_16976,N_16636,N_16708);
xnor U16977 (N_16977,N_16585,N_16576);
and U16978 (N_16978,N_16664,N_16677);
nand U16979 (N_16979,N_16542,N_16519);
nand U16980 (N_16980,N_16676,N_16721);
nand U16981 (N_16981,N_16556,N_16531);
or U16982 (N_16982,N_16539,N_16696);
nand U16983 (N_16983,N_16740,N_16541);
or U16984 (N_16984,N_16593,N_16601);
and U16985 (N_16985,N_16622,N_16636);
or U16986 (N_16986,N_16580,N_16652);
xnor U16987 (N_16987,N_16528,N_16680);
and U16988 (N_16988,N_16692,N_16565);
or U16989 (N_16989,N_16633,N_16572);
or U16990 (N_16990,N_16625,N_16651);
nand U16991 (N_16991,N_16712,N_16553);
or U16992 (N_16992,N_16562,N_16614);
and U16993 (N_16993,N_16563,N_16700);
xor U16994 (N_16994,N_16519,N_16646);
nand U16995 (N_16995,N_16695,N_16690);
or U16996 (N_16996,N_16653,N_16608);
or U16997 (N_16997,N_16695,N_16585);
nand U16998 (N_16998,N_16576,N_16509);
xor U16999 (N_16999,N_16687,N_16600);
nor U17000 (N_17000,N_16912,N_16991);
or U17001 (N_17001,N_16803,N_16981);
nor U17002 (N_17002,N_16999,N_16920);
xor U17003 (N_17003,N_16961,N_16784);
nand U17004 (N_17004,N_16909,N_16882);
nor U17005 (N_17005,N_16960,N_16923);
nor U17006 (N_17006,N_16992,N_16852);
or U17007 (N_17007,N_16964,N_16770);
and U17008 (N_17008,N_16934,N_16775);
xnor U17009 (N_17009,N_16815,N_16821);
and U17010 (N_17010,N_16820,N_16758);
nand U17011 (N_17011,N_16845,N_16858);
xnor U17012 (N_17012,N_16759,N_16935);
nand U17013 (N_17013,N_16799,N_16841);
nand U17014 (N_17014,N_16965,N_16808);
nor U17015 (N_17015,N_16833,N_16809);
nor U17016 (N_17016,N_16949,N_16864);
and U17017 (N_17017,N_16823,N_16898);
xor U17018 (N_17018,N_16943,N_16811);
and U17019 (N_17019,N_16879,N_16971);
nor U17020 (N_17020,N_16886,N_16804);
and U17021 (N_17021,N_16884,N_16831);
xnor U17022 (N_17022,N_16945,N_16780);
nand U17023 (N_17023,N_16910,N_16914);
nor U17024 (N_17024,N_16752,N_16894);
nor U17025 (N_17025,N_16984,N_16973);
nand U17026 (N_17026,N_16851,N_16849);
or U17027 (N_17027,N_16847,N_16860);
nand U17028 (N_17028,N_16816,N_16777);
or U17029 (N_17029,N_16985,N_16765);
or U17030 (N_17030,N_16903,N_16883);
nor U17031 (N_17031,N_16940,N_16848);
nor U17032 (N_17032,N_16931,N_16774);
or U17033 (N_17033,N_16790,N_16873);
or U17034 (N_17034,N_16783,N_16834);
nand U17035 (N_17035,N_16768,N_16987);
and U17036 (N_17036,N_16776,N_16767);
nand U17037 (N_17037,N_16766,N_16927);
nor U17038 (N_17038,N_16812,N_16838);
nor U17039 (N_17039,N_16966,N_16798);
nand U17040 (N_17040,N_16807,N_16936);
nand U17041 (N_17041,N_16843,N_16980);
or U17042 (N_17042,N_16896,N_16832);
nor U17043 (N_17043,N_16990,N_16900);
nand U17044 (N_17044,N_16806,N_16950);
or U17045 (N_17045,N_16958,N_16818);
xnor U17046 (N_17046,N_16953,N_16760);
or U17047 (N_17047,N_16885,N_16926);
or U17048 (N_17048,N_16773,N_16750);
and U17049 (N_17049,N_16836,N_16897);
nand U17050 (N_17050,N_16788,N_16772);
nor U17051 (N_17051,N_16871,N_16976);
nor U17052 (N_17052,N_16874,N_16891);
xor U17053 (N_17053,N_16859,N_16918);
nor U17054 (N_17054,N_16881,N_16754);
nor U17055 (N_17055,N_16865,N_16974);
nor U17056 (N_17056,N_16877,N_16876);
xnor U17057 (N_17057,N_16822,N_16786);
nor U17058 (N_17058,N_16878,N_16906);
nand U17059 (N_17059,N_16866,N_16956);
nand U17060 (N_17060,N_16872,N_16781);
xnor U17061 (N_17061,N_16939,N_16805);
or U17062 (N_17062,N_16967,N_16929);
nor U17063 (N_17063,N_16793,N_16925);
xor U17064 (N_17064,N_16797,N_16997);
nand U17065 (N_17065,N_16800,N_16930);
and U17066 (N_17066,N_16917,N_16826);
or U17067 (N_17067,N_16868,N_16948);
and U17068 (N_17068,N_16972,N_16944);
or U17069 (N_17069,N_16893,N_16957);
nor U17070 (N_17070,N_16996,N_16861);
or U17071 (N_17071,N_16814,N_16937);
nor U17072 (N_17072,N_16938,N_16890);
xor U17073 (N_17073,N_16796,N_16817);
nor U17074 (N_17074,N_16795,N_16875);
xnor U17075 (N_17075,N_16867,N_16870);
or U17076 (N_17076,N_16954,N_16762);
or U17077 (N_17077,N_16978,N_16869);
nor U17078 (N_17078,N_16915,N_16846);
or U17079 (N_17079,N_16941,N_16769);
xor U17080 (N_17080,N_16888,N_16892);
xor U17081 (N_17081,N_16899,N_16993);
or U17082 (N_17082,N_16970,N_16764);
or U17083 (N_17083,N_16771,N_16975);
and U17084 (N_17084,N_16850,N_16791);
or U17085 (N_17085,N_16810,N_16844);
xor U17086 (N_17086,N_16801,N_16928);
and U17087 (N_17087,N_16907,N_16998);
or U17088 (N_17088,N_16813,N_16802);
nand U17089 (N_17089,N_16761,N_16751);
xnor U17090 (N_17090,N_16830,N_16842);
or U17091 (N_17091,N_16895,N_16983);
nand U17092 (N_17092,N_16778,N_16779);
or U17093 (N_17093,N_16753,N_16977);
xnor U17094 (N_17094,N_16787,N_16854);
nand U17095 (N_17095,N_16825,N_16756);
and U17096 (N_17096,N_16785,N_16947);
and U17097 (N_17097,N_16819,N_16889);
or U17098 (N_17098,N_16946,N_16913);
or U17099 (N_17099,N_16855,N_16880);
xnor U17100 (N_17100,N_16994,N_16919);
xnor U17101 (N_17101,N_16828,N_16789);
xnor U17102 (N_17102,N_16840,N_16863);
nand U17103 (N_17103,N_16839,N_16905);
and U17104 (N_17104,N_16827,N_16989);
or U17105 (N_17105,N_16922,N_16853);
nand U17106 (N_17106,N_16755,N_16951);
nor U17107 (N_17107,N_16952,N_16911);
nand U17108 (N_17108,N_16932,N_16942);
or U17109 (N_17109,N_16969,N_16782);
nand U17110 (N_17110,N_16988,N_16986);
and U17111 (N_17111,N_16968,N_16837);
or U17112 (N_17112,N_16757,N_16963);
nor U17113 (N_17113,N_16862,N_16829);
and U17114 (N_17114,N_16835,N_16904);
nand U17115 (N_17115,N_16921,N_16924);
xnor U17116 (N_17116,N_16959,N_16962);
and U17117 (N_17117,N_16763,N_16856);
and U17118 (N_17118,N_16857,N_16916);
nor U17119 (N_17119,N_16792,N_16979);
xor U17120 (N_17120,N_16955,N_16982);
and U17121 (N_17121,N_16902,N_16794);
and U17122 (N_17122,N_16824,N_16995);
or U17123 (N_17123,N_16901,N_16933);
and U17124 (N_17124,N_16908,N_16887);
nor U17125 (N_17125,N_16892,N_16955);
nor U17126 (N_17126,N_16964,N_16780);
or U17127 (N_17127,N_16925,N_16824);
nand U17128 (N_17128,N_16800,N_16776);
xor U17129 (N_17129,N_16985,N_16883);
nand U17130 (N_17130,N_16866,N_16815);
or U17131 (N_17131,N_16846,N_16907);
xnor U17132 (N_17132,N_16881,N_16905);
xor U17133 (N_17133,N_16966,N_16851);
xnor U17134 (N_17134,N_16818,N_16944);
nand U17135 (N_17135,N_16937,N_16891);
xnor U17136 (N_17136,N_16819,N_16826);
nor U17137 (N_17137,N_16877,N_16896);
nand U17138 (N_17138,N_16835,N_16864);
nand U17139 (N_17139,N_16871,N_16817);
xnor U17140 (N_17140,N_16860,N_16890);
xnor U17141 (N_17141,N_16757,N_16919);
nor U17142 (N_17142,N_16883,N_16930);
nand U17143 (N_17143,N_16791,N_16986);
or U17144 (N_17144,N_16770,N_16805);
nand U17145 (N_17145,N_16894,N_16870);
or U17146 (N_17146,N_16796,N_16798);
nand U17147 (N_17147,N_16881,N_16909);
nand U17148 (N_17148,N_16791,N_16981);
nor U17149 (N_17149,N_16756,N_16827);
xor U17150 (N_17150,N_16898,N_16791);
nor U17151 (N_17151,N_16807,N_16761);
nand U17152 (N_17152,N_16912,N_16989);
or U17153 (N_17153,N_16802,N_16818);
nor U17154 (N_17154,N_16800,N_16984);
xnor U17155 (N_17155,N_16971,N_16909);
and U17156 (N_17156,N_16978,N_16875);
nand U17157 (N_17157,N_16987,N_16757);
nor U17158 (N_17158,N_16848,N_16908);
nor U17159 (N_17159,N_16828,N_16984);
or U17160 (N_17160,N_16778,N_16856);
nand U17161 (N_17161,N_16852,N_16757);
xnor U17162 (N_17162,N_16868,N_16801);
and U17163 (N_17163,N_16825,N_16755);
and U17164 (N_17164,N_16974,N_16775);
nor U17165 (N_17165,N_16899,N_16975);
and U17166 (N_17166,N_16867,N_16998);
or U17167 (N_17167,N_16961,N_16822);
or U17168 (N_17168,N_16860,N_16762);
nor U17169 (N_17169,N_16904,N_16966);
xnor U17170 (N_17170,N_16930,N_16971);
and U17171 (N_17171,N_16988,N_16939);
xnor U17172 (N_17172,N_16852,N_16862);
nor U17173 (N_17173,N_16989,N_16762);
or U17174 (N_17174,N_16812,N_16814);
or U17175 (N_17175,N_16780,N_16912);
and U17176 (N_17176,N_16795,N_16947);
xnor U17177 (N_17177,N_16970,N_16815);
nand U17178 (N_17178,N_16951,N_16865);
or U17179 (N_17179,N_16891,N_16763);
nand U17180 (N_17180,N_16947,N_16917);
nor U17181 (N_17181,N_16997,N_16755);
nor U17182 (N_17182,N_16856,N_16982);
or U17183 (N_17183,N_16974,N_16811);
nand U17184 (N_17184,N_16990,N_16946);
xor U17185 (N_17185,N_16764,N_16913);
or U17186 (N_17186,N_16968,N_16947);
nand U17187 (N_17187,N_16916,N_16959);
and U17188 (N_17188,N_16847,N_16810);
nand U17189 (N_17189,N_16791,N_16768);
nand U17190 (N_17190,N_16795,N_16974);
and U17191 (N_17191,N_16826,N_16937);
or U17192 (N_17192,N_16876,N_16884);
or U17193 (N_17193,N_16900,N_16822);
xor U17194 (N_17194,N_16891,N_16888);
nor U17195 (N_17195,N_16864,N_16885);
nand U17196 (N_17196,N_16954,N_16958);
nand U17197 (N_17197,N_16947,N_16906);
nand U17198 (N_17198,N_16792,N_16818);
nand U17199 (N_17199,N_16798,N_16795);
and U17200 (N_17200,N_16799,N_16867);
and U17201 (N_17201,N_16989,N_16908);
nand U17202 (N_17202,N_16930,N_16937);
or U17203 (N_17203,N_16793,N_16869);
and U17204 (N_17204,N_16756,N_16952);
nor U17205 (N_17205,N_16755,N_16877);
xor U17206 (N_17206,N_16926,N_16960);
nand U17207 (N_17207,N_16923,N_16893);
nor U17208 (N_17208,N_16914,N_16873);
nor U17209 (N_17209,N_16760,N_16976);
nor U17210 (N_17210,N_16790,N_16914);
and U17211 (N_17211,N_16859,N_16777);
xor U17212 (N_17212,N_16824,N_16926);
and U17213 (N_17213,N_16818,N_16942);
and U17214 (N_17214,N_16848,N_16914);
nand U17215 (N_17215,N_16898,N_16847);
or U17216 (N_17216,N_16843,N_16998);
nand U17217 (N_17217,N_16869,N_16900);
or U17218 (N_17218,N_16812,N_16775);
nand U17219 (N_17219,N_16999,N_16886);
xnor U17220 (N_17220,N_16993,N_16887);
and U17221 (N_17221,N_16821,N_16862);
or U17222 (N_17222,N_16818,N_16917);
nand U17223 (N_17223,N_16948,N_16815);
nand U17224 (N_17224,N_16945,N_16840);
and U17225 (N_17225,N_16904,N_16878);
nand U17226 (N_17226,N_16864,N_16970);
and U17227 (N_17227,N_16825,N_16773);
nor U17228 (N_17228,N_16954,N_16845);
xnor U17229 (N_17229,N_16754,N_16753);
and U17230 (N_17230,N_16845,N_16948);
nand U17231 (N_17231,N_16812,N_16789);
or U17232 (N_17232,N_16846,N_16906);
xnor U17233 (N_17233,N_16893,N_16850);
nand U17234 (N_17234,N_16854,N_16859);
nand U17235 (N_17235,N_16818,N_16889);
nand U17236 (N_17236,N_16873,N_16991);
xor U17237 (N_17237,N_16970,N_16811);
and U17238 (N_17238,N_16863,N_16782);
nand U17239 (N_17239,N_16758,N_16828);
nor U17240 (N_17240,N_16817,N_16827);
nand U17241 (N_17241,N_16977,N_16990);
nor U17242 (N_17242,N_16753,N_16986);
xor U17243 (N_17243,N_16980,N_16788);
xnor U17244 (N_17244,N_16752,N_16889);
and U17245 (N_17245,N_16924,N_16992);
or U17246 (N_17246,N_16772,N_16887);
xnor U17247 (N_17247,N_16942,N_16821);
xor U17248 (N_17248,N_16752,N_16982);
xor U17249 (N_17249,N_16953,N_16998);
and U17250 (N_17250,N_17099,N_17085);
or U17251 (N_17251,N_17245,N_17210);
and U17252 (N_17252,N_17057,N_17223);
and U17253 (N_17253,N_17022,N_17158);
and U17254 (N_17254,N_17198,N_17144);
and U17255 (N_17255,N_17184,N_17215);
nand U17256 (N_17256,N_17146,N_17028);
nand U17257 (N_17257,N_17081,N_17208);
and U17258 (N_17258,N_17050,N_17202);
xor U17259 (N_17259,N_17197,N_17153);
xnor U17260 (N_17260,N_17093,N_17042);
nand U17261 (N_17261,N_17172,N_17008);
nor U17262 (N_17262,N_17178,N_17249);
xor U17263 (N_17263,N_17154,N_17044);
and U17264 (N_17264,N_17060,N_17024);
xnor U17265 (N_17265,N_17241,N_17043);
nor U17266 (N_17266,N_17181,N_17211);
and U17267 (N_17267,N_17062,N_17032);
nand U17268 (N_17268,N_17013,N_17142);
or U17269 (N_17269,N_17035,N_17069);
nand U17270 (N_17270,N_17082,N_17168);
xnor U17271 (N_17271,N_17243,N_17037);
nor U17272 (N_17272,N_17025,N_17229);
and U17273 (N_17273,N_17121,N_17130);
nand U17274 (N_17274,N_17117,N_17126);
nand U17275 (N_17275,N_17119,N_17075);
xnor U17276 (N_17276,N_17113,N_17125);
and U17277 (N_17277,N_17204,N_17040);
nand U17278 (N_17278,N_17000,N_17091);
xor U17279 (N_17279,N_17180,N_17054);
or U17280 (N_17280,N_17226,N_17072);
or U17281 (N_17281,N_17034,N_17015);
xor U17282 (N_17282,N_17122,N_17009);
nor U17283 (N_17283,N_17170,N_17156);
xor U17284 (N_17284,N_17128,N_17166);
xnor U17285 (N_17285,N_17095,N_17221);
and U17286 (N_17286,N_17020,N_17007);
and U17287 (N_17287,N_17182,N_17171);
or U17288 (N_17288,N_17058,N_17003);
xor U17289 (N_17289,N_17176,N_17030);
or U17290 (N_17290,N_17134,N_17029);
or U17291 (N_17291,N_17157,N_17212);
xor U17292 (N_17292,N_17098,N_17195);
and U17293 (N_17293,N_17149,N_17010);
or U17294 (N_17294,N_17228,N_17232);
or U17295 (N_17295,N_17186,N_17143);
nand U17296 (N_17296,N_17151,N_17021);
and U17297 (N_17297,N_17155,N_17086);
or U17298 (N_17298,N_17139,N_17097);
or U17299 (N_17299,N_17011,N_17111);
nand U17300 (N_17300,N_17071,N_17014);
xor U17301 (N_17301,N_17135,N_17234);
and U17302 (N_17302,N_17231,N_17136);
and U17303 (N_17303,N_17235,N_17053);
or U17304 (N_17304,N_17065,N_17005);
nor U17305 (N_17305,N_17206,N_17070);
xnor U17306 (N_17306,N_17141,N_17110);
nand U17307 (N_17307,N_17036,N_17045);
and U17308 (N_17308,N_17055,N_17052);
or U17309 (N_17309,N_17209,N_17114);
and U17310 (N_17310,N_17224,N_17179);
xor U17311 (N_17311,N_17064,N_17160);
nor U17312 (N_17312,N_17188,N_17150);
nor U17313 (N_17313,N_17063,N_17246);
nor U17314 (N_17314,N_17049,N_17088);
nand U17315 (N_17315,N_17078,N_17059);
and U17316 (N_17316,N_17192,N_17177);
nand U17317 (N_17317,N_17175,N_17006);
and U17318 (N_17318,N_17191,N_17076);
nor U17319 (N_17319,N_17163,N_17079);
nor U17320 (N_17320,N_17219,N_17001);
xnor U17321 (N_17321,N_17220,N_17193);
or U17322 (N_17322,N_17068,N_17239);
nor U17323 (N_17323,N_17048,N_17129);
nor U17324 (N_17324,N_17084,N_17124);
or U17325 (N_17325,N_17100,N_17018);
xnor U17326 (N_17326,N_17019,N_17087);
or U17327 (N_17327,N_17066,N_17218);
nor U17328 (N_17328,N_17033,N_17041);
nor U17329 (N_17329,N_17214,N_17047);
nor U17330 (N_17330,N_17199,N_17222);
and U17331 (N_17331,N_17238,N_17090);
nand U17332 (N_17332,N_17216,N_17138);
xor U17333 (N_17333,N_17038,N_17004);
nor U17334 (N_17334,N_17169,N_17161);
or U17335 (N_17335,N_17173,N_17116);
or U17336 (N_17336,N_17002,N_17167);
or U17337 (N_17337,N_17240,N_17190);
nor U17338 (N_17338,N_17164,N_17165);
nand U17339 (N_17339,N_17080,N_17200);
nor U17340 (N_17340,N_17105,N_17089);
and U17341 (N_17341,N_17207,N_17183);
xnor U17342 (N_17342,N_17104,N_17152);
xor U17343 (N_17343,N_17194,N_17148);
and U17344 (N_17344,N_17187,N_17233);
and U17345 (N_17345,N_17247,N_17108);
and U17346 (N_17346,N_17140,N_17230);
nor U17347 (N_17347,N_17123,N_17203);
xor U17348 (N_17348,N_17225,N_17106);
and U17349 (N_17349,N_17073,N_17092);
nand U17350 (N_17350,N_17103,N_17027);
or U17351 (N_17351,N_17056,N_17074);
or U17352 (N_17352,N_17147,N_17120);
or U17353 (N_17353,N_17236,N_17189);
nand U17354 (N_17354,N_17039,N_17159);
and U17355 (N_17355,N_17096,N_17109);
nor U17356 (N_17356,N_17026,N_17067);
and U17357 (N_17357,N_17196,N_17145);
or U17358 (N_17358,N_17061,N_17046);
or U17359 (N_17359,N_17174,N_17101);
nor U17360 (N_17360,N_17227,N_17244);
and U17361 (N_17361,N_17205,N_17115);
xnor U17362 (N_17362,N_17023,N_17102);
and U17363 (N_17363,N_17077,N_17248);
and U17364 (N_17364,N_17017,N_17201);
nor U17365 (N_17365,N_17083,N_17131);
nand U17366 (N_17366,N_17107,N_17213);
and U17367 (N_17367,N_17031,N_17127);
xnor U17368 (N_17368,N_17112,N_17132);
or U17369 (N_17369,N_17051,N_17237);
xnor U17370 (N_17370,N_17217,N_17012);
or U17371 (N_17371,N_17133,N_17094);
nor U17372 (N_17372,N_17185,N_17016);
and U17373 (N_17373,N_17162,N_17137);
and U17374 (N_17374,N_17118,N_17242);
nor U17375 (N_17375,N_17180,N_17055);
xor U17376 (N_17376,N_17030,N_17042);
nand U17377 (N_17377,N_17094,N_17185);
nand U17378 (N_17378,N_17065,N_17022);
or U17379 (N_17379,N_17151,N_17032);
or U17380 (N_17380,N_17134,N_17018);
xor U17381 (N_17381,N_17074,N_17082);
and U17382 (N_17382,N_17093,N_17049);
xnor U17383 (N_17383,N_17173,N_17197);
nor U17384 (N_17384,N_17173,N_17058);
nor U17385 (N_17385,N_17037,N_17171);
and U17386 (N_17386,N_17152,N_17189);
nor U17387 (N_17387,N_17081,N_17116);
nand U17388 (N_17388,N_17222,N_17226);
and U17389 (N_17389,N_17163,N_17228);
or U17390 (N_17390,N_17140,N_17246);
or U17391 (N_17391,N_17146,N_17128);
nor U17392 (N_17392,N_17085,N_17046);
xor U17393 (N_17393,N_17190,N_17130);
and U17394 (N_17394,N_17001,N_17207);
nand U17395 (N_17395,N_17132,N_17114);
nand U17396 (N_17396,N_17052,N_17070);
or U17397 (N_17397,N_17175,N_17061);
nor U17398 (N_17398,N_17038,N_17113);
xnor U17399 (N_17399,N_17103,N_17026);
and U17400 (N_17400,N_17190,N_17007);
or U17401 (N_17401,N_17087,N_17134);
or U17402 (N_17402,N_17066,N_17089);
xor U17403 (N_17403,N_17222,N_17248);
xor U17404 (N_17404,N_17096,N_17152);
nor U17405 (N_17405,N_17174,N_17059);
and U17406 (N_17406,N_17005,N_17123);
or U17407 (N_17407,N_17165,N_17031);
nand U17408 (N_17408,N_17030,N_17186);
xor U17409 (N_17409,N_17024,N_17019);
and U17410 (N_17410,N_17037,N_17162);
nor U17411 (N_17411,N_17207,N_17179);
or U17412 (N_17412,N_17072,N_17023);
and U17413 (N_17413,N_17094,N_17143);
xnor U17414 (N_17414,N_17002,N_17079);
nor U17415 (N_17415,N_17151,N_17055);
or U17416 (N_17416,N_17228,N_17178);
nand U17417 (N_17417,N_17019,N_17227);
nand U17418 (N_17418,N_17218,N_17178);
nand U17419 (N_17419,N_17133,N_17091);
nand U17420 (N_17420,N_17123,N_17201);
nand U17421 (N_17421,N_17080,N_17188);
nand U17422 (N_17422,N_17014,N_17096);
or U17423 (N_17423,N_17080,N_17132);
nor U17424 (N_17424,N_17174,N_17050);
and U17425 (N_17425,N_17064,N_17143);
and U17426 (N_17426,N_17086,N_17159);
xor U17427 (N_17427,N_17164,N_17067);
xor U17428 (N_17428,N_17020,N_17193);
nor U17429 (N_17429,N_17240,N_17137);
and U17430 (N_17430,N_17128,N_17021);
or U17431 (N_17431,N_17036,N_17040);
xor U17432 (N_17432,N_17170,N_17137);
nand U17433 (N_17433,N_17125,N_17025);
xor U17434 (N_17434,N_17025,N_17142);
xnor U17435 (N_17435,N_17008,N_17128);
and U17436 (N_17436,N_17187,N_17047);
nor U17437 (N_17437,N_17004,N_17024);
xnor U17438 (N_17438,N_17191,N_17147);
or U17439 (N_17439,N_17058,N_17075);
or U17440 (N_17440,N_17226,N_17201);
nor U17441 (N_17441,N_17099,N_17081);
nand U17442 (N_17442,N_17175,N_17118);
xnor U17443 (N_17443,N_17197,N_17045);
and U17444 (N_17444,N_17054,N_17208);
and U17445 (N_17445,N_17033,N_17161);
or U17446 (N_17446,N_17207,N_17005);
nor U17447 (N_17447,N_17121,N_17115);
or U17448 (N_17448,N_17069,N_17153);
nor U17449 (N_17449,N_17170,N_17214);
nor U17450 (N_17450,N_17098,N_17173);
xor U17451 (N_17451,N_17239,N_17111);
or U17452 (N_17452,N_17202,N_17159);
nand U17453 (N_17453,N_17060,N_17150);
nor U17454 (N_17454,N_17118,N_17148);
and U17455 (N_17455,N_17141,N_17176);
nor U17456 (N_17456,N_17219,N_17208);
xnor U17457 (N_17457,N_17133,N_17109);
and U17458 (N_17458,N_17018,N_17021);
nor U17459 (N_17459,N_17173,N_17206);
and U17460 (N_17460,N_17115,N_17105);
nand U17461 (N_17461,N_17034,N_17170);
nand U17462 (N_17462,N_17046,N_17094);
nand U17463 (N_17463,N_17182,N_17076);
nand U17464 (N_17464,N_17067,N_17041);
nor U17465 (N_17465,N_17187,N_17075);
xor U17466 (N_17466,N_17119,N_17159);
and U17467 (N_17467,N_17223,N_17201);
xnor U17468 (N_17468,N_17093,N_17142);
nor U17469 (N_17469,N_17174,N_17223);
or U17470 (N_17470,N_17201,N_17082);
nand U17471 (N_17471,N_17183,N_17198);
and U17472 (N_17472,N_17174,N_17235);
nand U17473 (N_17473,N_17241,N_17171);
and U17474 (N_17474,N_17229,N_17198);
xor U17475 (N_17475,N_17113,N_17044);
or U17476 (N_17476,N_17127,N_17054);
nor U17477 (N_17477,N_17167,N_17108);
and U17478 (N_17478,N_17056,N_17092);
or U17479 (N_17479,N_17244,N_17048);
nand U17480 (N_17480,N_17186,N_17079);
and U17481 (N_17481,N_17236,N_17053);
xor U17482 (N_17482,N_17102,N_17191);
nand U17483 (N_17483,N_17015,N_17122);
nor U17484 (N_17484,N_17058,N_17171);
and U17485 (N_17485,N_17079,N_17130);
nor U17486 (N_17486,N_17187,N_17012);
or U17487 (N_17487,N_17166,N_17083);
or U17488 (N_17488,N_17027,N_17161);
nand U17489 (N_17489,N_17130,N_17009);
nor U17490 (N_17490,N_17083,N_17171);
and U17491 (N_17491,N_17003,N_17022);
or U17492 (N_17492,N_17244,N_17101);
or U17493 (N_17493,N_17121,N_17089);
nand U17494 (N_17494,N_17115,N_17194);
xor U17495 (N_17495,N_17234,N_17039);
xor U17496 (N_17496,N_17227,N_17201);
xnor U17497 (N_17497,N_17096,N_17161);
nand U17498 (N_17498,N_17064,N_17183);
nand U17499 (N_17499,N_17090,N_17014);
or U17500 (N_17500,N_17354,N_17485);
nand U17501 (N_17501,N_17250,N_17325);
and U17502 (N_17502,N_17462,N_17257);
and U17503 (N_17503,N_17466,N_17261);
xnor U17504 (N_17504,N_17368,N_17469);
and U17505 (N_17505,N_17262,N_17381);
and U17506 (N_17506,N_17339,N_17323);
or U17507 (N_17507,N_17476,N_17451);
and U17508 (N_17508,N_17345,N_17346);
or U17509 (N_17509,N_17319,N_17364);
xnor U17510 (N_17510,N_17407,N_17461);
and U17511 (N_17511,N_17292,N_17498);
xnor U17512 (N_17512,N_17371,N_17444);
nor U17513 (N_17513,N_17265,N_17280);
nor U17514 (N_17514,N_17317,N_17380);
xnor U17515 (N_17515,N_17449,N_17360);
xnor U17516 (N_17516,N_17460,N_17430);
xnor U17517 (N_17517,N_17379,N_17489);
and U17518 (N_17518,N_17281,N_17409);
or U17519 (N_17519,N_17258,N_17412);
xor U17520 (N_17520,N_17434,N_17361);
and U17521 (N_17521,N_17482,N_17357);
xor U17522 (N_17522,N_17279,N_17473);
and U17523 (N_17523,N_17484,N_17336);
or U17524 (N_17524,N_17411,N_17415);
or U17525 (N_17525,N_17266,N_17429);
nand U17526 (N_17526,N_17278,N_17295);
nor U17527 (N_17527,N_17367,N_17495);
and U17528 (N_17528,N_17401,N_17387);
or U17529 (N_17529,N_17303,N_17352);
or U17530 (N_17530,N_17403,N_17329);
nand U17531 (N_17531,N_17400,N_17386);
nor U17532 (N_17532,N_17391,N_17457);
nor U17533 (N_17533,N_17486,N_17418);
or U17534 (N_17534,N_17388,N_17314);
nand U17535 (N_17535,N_17343,N_17491);
nand U17536 (N_17536,N_17350,N_17297);
or U17537 (N_17537,N_17471,N_17341);
and U17538 (N_17538,N_17494,N_17274);
nor U17539 (N_17539,N_17456,N_17299);
and U17540 (N_17540,N_17393,N_17335);
nor U17541 (N_17541,N_17284,N_17478);
nand U17542 (N_17542,N_17394,N_17253);
and U17543 (N_17543,N_17497,N_17291);
nor U17544 (N_17544,N_17472,N_17337);
xor U17545 (N_17545,N_17488,N_17334);
xor U17546 (N_17546,N_17384,N_17363);
nand U17547 (N_17547,N_17263,N_17269);
nand U17548 (N_17548,N_17358,N_17463);
or U17549 (N_17549,N_17277,N_17406);
nor U17550 (N_17550,N_17296,N_17397);
nand U17551 (N_17551,N_17419,N_17405);
nand U17552 (N_17552,N_17426,N_17382);
nand U17553 (N_17553,N_17356,N_17428);
or U17554 (N_17554,N_17294,N_17424);
nand U17555 (N_17555,N_17441,N_17435);
xnor U17556 (N_17556,N_17313,N_17378);
nand U17557 (N_17557,N_17342,N_17398);
nor U17558 (N_17558,N_17465,N_17458);
nor U17559 (N_17559,N_17286,N_17353);
xnor U17560 (N_17560,N_17302,N_17309);
and U17561 (N_17561,N_17300,N_17445);
xor U17562 (N_17562,N_17433,N_17321);
or U17563 (N_17563,N_17422,N_17453);
or U17564 (N_17564,N_17355,N_17328);
or U17565 (N_17565,N_17308,N_17413);
and U17566 (N_17566,N_17362,N_17268);
or U17567 (N_17567,N_17493,N_17331);
nor U17568 (N_17568,N_17327,N_17390);
xnor U17569 (N_17569,N_17320,N_17365);
nand U17570 (N_17570,N_17431,N_17298);
nor U17571 (N_17571,N_17282,N_17454);
or U17572 (N_17572,N_17402,N_17369);
or U17573 (N_17573,N_17370,N_17414);
nand U17574 (N_17574,N_17270,N_17450);
and U17575 (N_17575,N_17396,N_17487);
and U17576 (N_17576,N_17479,N_17492);
xnor U17577 (N_17577,N_17395,N_17264);
or U17578 (N_17578,N_17349,N_17490);
xor U17579 (N_17579,N_17307,N_17375);
or U17580 (N_17580,N_17276,N_17304);
or U17581 (N_17581,N_17417,N_17446);
and U17582 (N_17582,N_17275,N_17410);
xor U17583 (N_17583,N_17420,N_17448);
and U17584 (N_17584,N_17436,N_17322);
nor U17585 (N_17585,N_17464,N_17289);
or U17586 (N_17586,N_17427,N_17372);
or U17587 (N_17587,N_17338,N_17423);
nor U17588 (N_17588,N_17438,N_17283);
and U17589 (N_17589,N_17373,N_17481);
xor U17590 (N_17590,N_17315,N_17425);
xnor U17591 (N_17591,N_17359,N_17273);
xnor U17592 (N_17592,N_17340,N_17452);
xor U17593 (N_17593,N_17293,N_17290);
nand U17594 (N_17594,N_17383,N_17260);
and U17595 (N_17595,N_17399,N_17312);
nand U17596 (N_17596,N_17316,N_17252);
or U17597 (N_17597,N_17468,N_17271);
and U17598 (N_17598,N_17389,N_17377);
or U17599 (N_17599,N_17404,N_17374);
nand U17600 (N_17600,N_17459,N_17496);
or U17601 (N_17601,N_17256,N_17251);
nor U17602 (N_17602,N_17267,N_17474);
xor U17603 (N_17603,N_17310,N_17285);
or U17604 (N_17604,N_17288,N_17326);
xnor U17605 (N_17605,N_17287,N_17366);
xor U17606 (N_17606,N_17305,N_17467);
xor U17607 (N_17607,N_17477,N_17439);
or U17608 (N_17608,N_17330,N_17416);
and U17609 (N_17609,N_17311,N_17442);
and U17610 (N_17610,N_17347,N_17499);
nand U17611 (N_17611,N_17455,N_17324);
xnor U17612 (N_17612,N_17432,N_17254);
and U17613 (N_17613,N_17480,N_17351);
and U17614 (N_17614,N_17255,N_17344);
xor U17615 (N_17615,N_17318,N_17392);
and U17616 (N_17616,N_17376,N_17333);
or U17617 (N_17617,N_17272,N_17385);
or U17618 (N_17618,N_17443,N_17348);
or U17619 (N_17619,N_17408,N_17259);
nand U17620 (N_17620,N_17475,N_17437);
and U17621 (N_17621,N_17301,N_17306);
and U17622 (N_17622,N_17447,N_17483);
xor U17623 (N_17623,N_17421,N_17440);
and U17624 (N_17624,N_17470,N_17332);
nand U17625 (N_17625,N_17475,N_17317);
nand U17626 (N_17626,N_17421,N_17459);
nor U17627 (N_17627,N_17307,N_17339);
and U17628 (N_17628,N_17359,N_17262);
and U17629 (N_17629,N_17409,N_17491);
and U17630 (N_17630,N_17326,N_17458);
nor U17631 (N_17631,N_17344,N_17343);
xor U17632 (N_17632,N_17440,N_17409);
xnor U17633 (N_17633,N_17251,N_17379);
nand U17634 (N_17634,N_17452,N_17253);
or U17635 (N_17635,N_17436,N_17497);
nand U17636 (N_17636,N_17440,N_17403);
nor U17637 (N_17637,N_17494,N_17453);
xnor U17638 (N_17638,N_17371,N_17451);
nor U17639 (N_17639,N_17252,N_17321);
and U17640 (N_17640,N_17377,N_17495);
and U17641 (N_17641,N_17269,N_17266);
nand U17642 (N_17642,N_17439,N_17331);
or U17643 (N_17643,N_17401,N_17414);
and U17644 (N_17644,N_17484,N_17283);
and U17645 (N_17645,N_17451,N_17487);
or U17646 (N_17646,N_17464,N_17413);
xor U17647 (N_17647,N_17314,N_17279);
xnor U17648 (N_17648,N_17344,N_17356);
nor U17649 (N_17649,N_17281,N_17346);
nor U17650 (N_17650,N_17259,N_17492);
nand U17651 (N_17651,N_17341,N_17460);
nor U17652 (N_17652,N_17340,N_17493);
xor U17653 (N_17653,N_17385,N_17265);
nor U17654 (N_17654,N_17432,N_17454);
xor U17655 (N_17655,N_17474,N_17285);
or U17656 (N_17656,N_17274,N_17329);
or U17657 (N_17657,N_17406,N_17329);
nand U17658 (N_17658,N_17309,N_17498);
nor U17659 (N_17659,N_17448,N_17476);
xor U17660 (N_17660,N_17325,N_17259);
nor U17661 (N_17661,N_17266,N_17333);
and U17662 (N_17662,N_17448,N_17481);
and U17663 (N_17663,N_17324,N_17484);
nor U17664 (N_17664,N_17371,N_17422);
xor U17665 (N_17665,N_17371,N_17260);
nand U17666 (N_17666,N_17484,N_17314);
and U17667 (N_17667,N_17313,N_17344);
or U17668 (N_17668,N_17258,N_17323);
or U17669 (N_17669,N_17347,N_17262);
and U17670 (N_17670,N_17376,N_17476);
or U17671 (N_17671,N_17421,N_17446);
or U17672 (N_17672,N_17478,N_17404);
nand U17673 (N_17673,N_17419,N_17344);
and U17674 (N_17674,N_17315,N_17265);
and U17675 (N_17675,N_17288,N_17385);
nor U17676 (N_17676,N_17274,N_17431);
nor U17677 (N_17677,N_17482,N_17393);
nor U17678 (N_17678,N_17297,N_17325);
xor U17679 (N_17679,N_17267,N_17443);
nor U17680 (N_17680,N_17499,N_17256);
nand U17681 (N_17681,N_17332,N_17495);
or U17682 (N_17682,N_17331,N_17324);
nor U17683 (N_17683,N_17352,N_17276);
and U17684 (N_17684,N_17362,N_17256);
nor U17685 (N_17685,N_17419,N_17390);
nand U17686 (N_17686,N_17348,N_17388);
and U17687 (N_17687,N_17342,N_17360);
nor U17688 (N_17688,N_17371,N_17251);
xor U17689 (N_17689,N_17260,N_17342);
and U17690 (N_17690,N_17496,N_17373);
or U17691 (N_17691,N_17417,N_17254);
nand U17692 (N_17692,N_17444,N_17479);
nor U17693 (N_17693,N_17305,N_17262);
and U17694 (N_17694,N_17342,N_17409);
or U17695 (N_17695,N_17486,N_17455);
or U17696 (N_17696,N_17339,N_17487);
and U17697 (N_17697,N_17426,N_17326);
and U17698 (N_17698,N_17357,N_17307);
nand U17699 (N_17699,N_17485,N_17360);
or U17700 (N_17700,N_17476,N_17260);
nand U17701 (N_17701,N_17365,N_17380);
nor U17702 (N_17702,N_17258,N_17394);
nor U17703 (N_17703,N_17444,N_17311);
or U17704 (N_17704,N_17470,N_17312);
or U17705 (N_17705,N_17338,N_17493);
nor U17706 (N_17706,N_17487,N_17349);
nand U17707 (N_17707,N_17408,N_17389);
xnor U17708 (N_17708,N_17312,N_17488);
nor U17709 (N_17709,N_17405,N_17399);
xor U17710 (N_17710,N_17304,N_17386);
and U17711 (N_17711,N_17366,N_17347);
xnor U17712 (N_17712,N_17336,N_17255);
or U17713 (N_17713,N_17405,N_17356);
xnor U17714 (N_17714,N_17442,N_17392);
or U17715 (N_17715,N_17446,N_17365);
or U17716 (N_17716,N_17327,N_17388);
or U17717 (N_17717,N_17497,N_17277);
and U17718 (N_17718,N_17411,N_17423);
and U17719 (N_17719,N_17271,N_17369);
nand U17720 (N_17720,N_17452,N_17482);
or U17721 (N_17721,N_17417,N_17430);
nand U17722 (N_17722,N_17434,N_17419);
and U17723 (N_17723,N_17410,N_17309);
xor U17724 (N_17724,N_17448,N_17332);
nor U17725 (N_17725,N_17383,N_17251);
or U17726 (N_17726,N_17309,N_17473);
and U17727 (N_17727,N_17255,N_17444);
nor U17728 (N_17728,N_17327,N_17350);
or U17729 (N_17729,N_17270,N_17347);
or U17730 (N_17730,N_17255,N_17342);
or U17731 (N_17731,N_17356,N_17374);
and U17732 (N_17732,N_17389,N_17414);
or U17733 (N_17733,N_17253,N_17378);
nand U17734 (N_17734,N_17431,N_17484);
xor U17735 (N_17735,N_17463,N_17299);
nor U17736 (N_17736,N_17334,N_17380);
or U17737 (N_17737,N_17272,N_17321);
nor U17738 (N_17738,N_17429,N_17286);
and U17739 (N_17739,N_17432,N_17476);
nand U17740 (N_17740,N_17289,N_17319);
nand U17741 (N_17741,N_17396,N_17280);
and U17742 (N_17742,N_17370,N_17419);
nor U17743 (N_17743,N_17476,N_17378);
and U17744 (N_17744,N_17298,N_17254);
or U17745 (N_17745,N_17338,N_17276);
and U17746 (N_17746,N_17463,N_17359);
or U17747 (N_17747,N_17356,N_17287);
or U17748 (N_17748,N_17372,N_17265);
and U17749 (N_17749,N_17471,N_17447);
nor U17750 (N_17750,N_17724,N_17504);
and U17751 (N_17751,N_17643,N_17613);
xnor U17752 (N_17752,N_17733,N_17746);
or U17753 (N_17753,N_17521,N_17537);
and U17754 (N_17754,N_17742,N_17666);
and U17755 (N_17755,N_17561,N_17703);
nand U17756 (N_17756,N_17715,N_17551);
nor U17757 (N_17757,N_17570,N_17594);
or U17758 (N_17758,N_17667,N_17658);
nand U17759 (N_17759,N_17595,N_17529);
nand U17760 (N_17760,N_17527,N_17701);
and U17761 (N_17761,N_17720,N_17590);
nor U17762 (N_17762,N_17679,N_17502);
nand U17763 (N_17763,N_17705,N_17671);
nand U17764 (N_17764,N_17602,N_17525);
nand U17765 (N_17765,N_17545,N_17744);
and U17766 (N_17766,N_17543,N_17706);
and U17767 (N_17767,N_17695,N_17621);
and U17768 (N_17768,N_17597,N_17592);
and U17769 (N_17769,N_17653,N_17648);
nand U17770 (N_17770,N_17688,N_17712);
or U17771 (N_17771,N_17611,N_17513);
nand U17772 (N_17772,N_17532,N_17646);
nand U17773 (N_17773,N_17596,N_17748);
nor U17774 (N_17774,N_17636,N_17586);
nand U17775 (N_17775,N_17538,N_17540);
xor U17776 (N_17776,N_17503,N_17536);
or U17777 (N_17777,N_17605,N_17631);
xnor U17778 (N_17778,N_17740,N_17506);
or U17779 (N_17779,N_17673,N_17610);
nor U17780 (N_17780,N_17694,N_17584);
or U17781 (N_17781,N_17734,N_17573);
xnor U17782 (N_17782,N_17591,N_17635);
or U17783 (N_17783,N_17515,N_17736);
nand U17784 (N_17784,N_17574,N_17580);
xor U17785 (N_17785,N_17560,N_17689);
xnor U17786 (N_17786,N_17716,N_17566);
xnor U17787 (N_17787,N_17721,N_17517);
xor U17788 (N_17788,N_17735,N_17674);
nand U17789 (N_17789,N_17539,N_17691);
and U17790 (N_17790,N_17672,N_17678);
or U17791 (N_17791,N_17697,N_17656);
nand U17792 (N_17792,N_17509,N_17546);
xnor U17793 (N_17793,N_17550,N_17626);
and U17794 (N_17794,N_17585,N_17544);
or U17795 (N_17795,N_17582,N_17690);
or U17796 (N_17796,N_17711,N_17696);
nand U17797 (N_17797,N_17680,N_17661);
nor U17798 (N_17798,N_17670,N_17535);
nor U17799 (N_17799,N_17552,N_17718);
or U17800 (N_17800,N_17575,N_17554);
nand U17801 (N_17801,N_17511,N_17647);
xor U17802 (N_17802,N_17632,N_17624);
and U17803 (N_17803,N_17668,N_17524);
and U17804 (N_17804,N_17729,N_17641);
nor U17805 (N_17805,N_17514,N_17567);
or U17806 (N_17806,N_17604,N_17687);
and U17807 (N_17807,N_17642,N_17704);
nor U17808 (N_17808,N_17659,N_17702);
and U17809 (N_17809,N_17665,N_17533);
xnor U17810 (N_17810,N_17558,N_17583);
and U17811 (N_17811,N_17714,N_17739);
or U17812 (N_17812,N_17634,N_17660);
nor U17813 (N_17813,N_17588,N_17581);
or U17814 (N_17814,N_17662,N_17542);
nand U17815 (N_17815,N_17548,N_17587);
and U17816 (N_17816,N_17644,N_17708);
or U17817 (N_17817,N_17501,N_17505);
or U17818 (N_17818,N_17657,N_17518);
xnor U17819 (N_17819,N_17526,N_17738);
and U17820 (N_17820,N_17675,N_17625);
xor U17821 (N_17821,N_17622,N_17549);
or U17822 (N_17822,N_17599,N_17652);
or U17823 (N_17823,N_17512,N_17664);
and U17824 (N_17824,N_17645,N_17699);
or U17825 (N_17825,N_17609,N_17726);
and U17826 (N_17826,N_17614,N_17562);
xor U17827 (N_17827,N_17601,N_17743);
nand U17828 (N_17828,N_17685,N_17598);
and U17829 (N_17829,N_17654,N_17722);
xor U17830 (N_17830,N_17737,N_17516);
xor U17831 (N_17831,N_17682,N_17713);
nand U17832 (N_17832,N_17693,N_17572);
nor U17833 (N_17833,N_17676,N_17723);
nand U17834 (N_17834,N_17568,N_17618);
nand U17835 (N_17835,N_17619,N_17728);
nor U17836 (N_17836,N_17589,N_17633);
nor U17837 (N_17837,N_17727,N_17725);
and U17838 (N_17838,N_17640,N_17523);
and U17839 (N_17839,N_17651,N_17557);
nor U17840 (N_17840,N_17747,N_17510);
xor U17841 (N_17841,N_17745,N_17577);
nand U17842 (N_17842,N_17681,N_17522);
nor U17843 (N_17843,N_17617,N_17534);
and U17844 (N_17844,N_17629,N_17683);
or U17845 (N_17845,N_17707,N_17528);
nand U17846 (N_17846,N_17593,N_17547);
xnor U17847 (N_17847,N_17564,N_17563);
xnor U17848 (N_17848,N_17508,N_17556);
xnor U17849 (N_17849,N_17531,N_17741);
nor U17850 (N_17850,N_17616,N_17710);
nand U17851 (N_17851,N_17606,N_17639);
and U17852 (N_17852,N_17569,N_17520);
nand U17853 (N_17853,N_17541,N_17638);
nor U17854 (N_17854,N_17628,N_17698);
nor U17855 (N_17855,N_17717,N_17612);
or U17856 (N_17856,N_17709,N_17686);
and U17857 (N_17857,N_17507,N_17669);
xnor U17858 (N_17858,N_17637,N_17579);
or U17859 (N_17859,N_17555,N_17607);
and U17860 (N_17860,N_17630,N_17649);
xor U17861 (N_17861,N_17650,N_17730);
xor U17862 (N_17862,N_17603,N_17620);
nand U17863 (N_17863,N_17608,N_17615);
nor U17864 (N_17864,N_17565,N_17623);
and U17865 (N_17865,N_17731,N_17732);
or U17866 (N_17866,N_17530,N_17749);
nor U17867 (N_17867,N_17553,N_17677);
and U17868 (N_17868,N_17600,N_17692);
or U17869 (N_17869,N_17700,N_17571);
and U17870 (N_17870,N_17578,N_17684);
nor U17871 (N_17871,N_17719,N_17559);
and U17872 (N_17872,N_17627,N_17519);
nand U17873 (N_17873,N_17576,N_17655);
nor U17874 (N_17874,N_17663,N_17500);
nor U17875 (N_17875,N_17716,N_17588);
nor U17876 (N_17876,N_17553,N_17555);
and U17877 (N_17877,N_17539,N_17684);
xor U17878 (N_17878,N_17668,N_17664);
and U17879 (N_17879,N_17524,N_17745);
nand U17880 (N_17880,N_17662,N_17746);
xor U17881 (N_17881,N_17615,N_17521);
and U17882 (N_17882,N_17626,N_17696);
nor U17883 (N_17883,N_17702,N_17538);
nand U17884 (N_17884,N_17588,N_17602);
and U17885 (N_17885,N_17590,N_17628);
or U17886 (N_17886,N_17506,N_17661);
and U17887 (N_17887,N_17670,N_17503);
xnor U17888 (N_17888,N_17507,N_17544);
nand U17889 (N_17889,N_17680,N_17715);
nor U17890 (N_17890,N_17727,N_17572);
nand U17891 (N_17891,N_17619,N_17594);
or U17892 (N_17892,N_17609,N_17724);
and U17893 (N_17893,N_17705,N_17686);
nor U17894 (N_17894,N_17556,N_17703);
and U17895 (N_17895,N_17695,N_17564);
nor U17896 (N_17896,N_17625,N_17618);
and U17897 (N_17897,N_17747,N_17675);
nand U17898 (N_17898,N_17503,N_17682);
nand U17899 (N_17899,N_17649,N_17704);
nor U17900 (N_17900,N_17564,N_17644);
nand U17901 (N_17901,N_17614,N_17700);
nand U17902 (N_17902,N_17519,N_17738);
xor U17903 (N_17903,N_17547,N_17657);
nand U17904 (N_17904,N_17632,N_17500);
nor U17905 (N_17905,N_17518,N_17628);
nand U17906 (N_17906,N_17660,N_17744);
and U17907 (N_17907,N_17676,N_17508);
xor U17908 (N_17908,N_17692,N_17541);
nand U17909 (N_17909,N_17748,N_17718);
or U17910 (N_17910,N_17518,N_17693);
or U17911 (N_17911,N_17646,N_17652);
nor U17912 (N_17912,N_17581,N_17538);
nor U17913 (N_17913,N_17685,N_17580);
nor U17914 (N_17914,N_17586,N_17573);
and U17915 (N_17915,N_17579,N_17656);
nor U17916 (N_17916,N_17706,N_17724);
nand U17917 (N_17917,N_17570,N_17736);
nand U17918 (N_17918,N_17532,N_17685);
nor U17919 (N_17919,N_17538,N_17510);
or U17920 (N_17920,N_17560,N_17564);
and U17921 (N_17921,N_17543,N_17608);
xor U17922 (N_17922,N_17632,N_17569);
nor U17923 (N_17923,N_17743,N_17550);
and U17924 (N_17924,N_17707,N_17582);
xor U17925 (N_17925,N_17534,N_17601);
xor U17926 (N_17926,N_17666,N_17588);
and U17927 (N_17927,N_17668,N_17616);
or U17928 (N_17928,N_17635,N_17508);
and U17929 (N_17929,N_17534,N_17694);
xor U17930 (N_17930,N_17588,N_17545);
nor U17931 (N_17931,N_17604,N_17577);
xor U17932 (N_17932,N_17543,N_17578);
nand U17933 (N_17933,N_17530,N_17654);
nand U17934 (N_17934,N_17687,N_17549);
and U17935 (N_17935,N_17744,N_17560);
xor U17936 (N_17936,N_17681,N_17747);
nor U17937 (N_17937,N_17540,N_17519);
xor U17938 (N_17938,N_17669,N_17590);
xor U17939 (N_17939,N_17561,N_17530);
and U17940 (N_17940,N_17730,N_17557);
nor U17941 (N_17941,N_17742,N_17648);
xnor U17942 (N_17942,N_17703,N_17708);
xnor U17943 (N_17943,N_17741,N_17648);
or U17944 (N_17944,N_17746,N_17702);
nor U17945 (N_17945,N_17599,N_17739);
or U17946 (N_17946,N_17510,N_17662);
xnor U17947 (N_17947,N_17541,N_17558);
nor U17948 (N_17948,N_17591,N_17600);
or U17949 (N_17949,N_17523,N_17520);
xnor U17950 (N_17950,N_17627,N_17645);
and U17951 (N_17951,N_17621,N_17691);
xnor U17952 (N_17952,N_17625,N_17547);
and U17953 (N_17953,N_17589,N_17690);
nand U17954 (N_17954,N_17628,N_17714);
and U17955 (N_17955,N_17726,N_17695);
or U17956 (N_17956,N_17592,N_17693);
and U17957 (N_17957,N_17660,N_17523);
xor U17958 (N_17958,N_17622,N_17533);
nand U17959 (N_17959,N_17565,N_17704);
xnor U17960 (N_17960,N_17588,N_17573);
or U17961 (N_17961,N_17558,N_17682);
nor U17962 (N_17962,N_17687,N_17632);
or U17963 (N_17963,N_17681,N_17521);
and U17964 (N_17964,N_17713,N_17554);
nor U17965 (N_17965,N_17641,N_17733);
or U17966 (N_17966,N_17661,N_17635);
nand U17967 (N_17967,N_17550,N_17708);
nand U17968 (N_17968,N_17671,N_17680);
or U17969 (N_17969,N_17663,N_17725);
xnor U17970 (N_17970,N_17637,N_17739);
xnor U17971 (N_17971,N_17523,N_17643);
nand U17972 (N_17972,N_17595,N_17721);
nor U17973 (N_17973,N_17655,N_17641);
nand U17974 (N_17974,N_17574,N_17720);
xor U17975 (N_17975,N_17608,N_17530);
and U17976 (N_17976,N_17581,N_17612);
nand U17977 (N_17977,N_17527,N_17722);
nor U17978 (N_17978,N_17505,N_17667);
xnor U17979 (N_17979,N_17591,N_17573);
xor U17980 (N_17980,N_17534,N_17741);
xnor U17981 (N_17981,N_17668,N_17533);
xor U17982 (N_17982,N_17594,N_17507);
nor U17983 (N_17983,N_17673,N_17600);
and U17984 (N_17984,N_17521,N_17662);
xnor U17985 (N_17985,N_17629,N_17587);
or U17986 (N_17986,N_17586,N_17543);
or U17987 (N_17987,N_17530,N_17643);
nor U17988 (N_17988,N_17709,N_17704);
nand U17989 (N_17989,N_17629,N_17603);
xnor U17990 (N_17990,N_17692,N_17682);
and U17991 (N_17991,N_17517,N_17660);
or U17992 (N_17992,N_17671,N_17539);
nor U17993 (N_17993,N_17701,N_17518);
nand U17994 (N_17994,N_17678,N_17529);
nand U17995 (N_17995,N_17526,N_17539);
or U17996 (N_17996,N_17594,N_17711);
and U17997 (N_17997,N_17737,N_17637);
and U17998 (N_17998,N_17714,N_17525);
xor U17999 (N_17999,N_17618,N_17550);
and U18000 (N_18000,N_17808,N_17866);
nand U18001 (N_18001,N_17881,N_17963);
nor U18002 (N_18002,N_17806,N_17867);
and U18003 (N_18003,N_17843,N_17933);
nand U18004 (N_18004,N_17814,N_17753);
xor U18005 (N_18005,N_17918,N_17955);
nor U18006 (N_18006,N_17812,N_17770);
nand U18007 (N_18007,N_17829,N_17862);
xnor U18008 (N_18008,N_17844,N_17977);
and U18009 (N_18009,N_17868,N_17997);
nor U18010 (N_18010,N_17818,N_17995);
or U18011 (N_18011,N_17876,N_17830);
nor U18012 (N_18012,N_17809,N_17904);
or U18013 (N_18013,N_17785,N_17750);
xor U18014 (N_18014,N_17931,N_17973);
nand U18015 (N_18015,N_17765,N_17824);
xnor U18016 (N_18016,N_17822,N_17888);
xnor U18017 (N_18017,N_17902,N_17864);
nand U18018 (N_18018,N_17797,N_17762);
nor U18019 (N_18019,N_17869,N_17865);
and U18020 (N_18020,N_17805,N_17776);
nand U18021 (N_18021,N_17878,N_17924);
nand U18022 (N_18022,N_17959,N_17898);
xnor U18023 (N_18023,N_17919,N_17943);
and U18024 (N_18024,N_17858,N_17999);
nor U18025 (N_18025,N_17796,N_17758);
nand U18026 (N_18026,N_17828,N_17942);
nor U18027 (N_18027,N_17965,N_17978);
or U18028 (N_18028,N_17795,N_17875);
and U18029 (N_18029,N_17907,N_17948);
and U18030 (N_18030,N_17927,N_17981);
xor U18031 (N_18031,N_17764,N_17870);
xnor U18032 (N_18032,N_17816,N_17923);
nor U18033 (N_18033,N_17893,N_17825);
nor U18034 (N_18034,N_17968,N_17820);
or U18035 (N_18035,N_17873,N_17766);
or U18036 (N_18036,N_17921,N_17819);
nand U18037 (N_18037,N_17961,N_17944);
nand U18038 (N_18038,N_17979,N_17863);
or U18039 (N_18039,N_17794,N_17984);
nor U18040 (N_18040,N_17789,N_17859);
nor U18041 (N_18041,N_17953,N_17839);
or U18042 (N_18042,N_17767,N_17782);
or U18043 (N_18043,N_17817,N_17905);
nand U18044 (N_18044,N_17990,N_17799);
and U18045 (N_18045,N_17886,N_17772);
or U18046 (N_18046,N_17987,N_17771);
nand U18047 (N_18047,N_17930,N_17912);
or U18048 (N_18048,N_17952,N_17761);
and U18049 (N_18049,N_17976,N_17803);
xnor U18050 (N_18050,N_17848,N_17956);
xnor U18051 (N_18051,N_17926,N_17768);
or U18052 (N_18052,N_17983,N_17841);
or U18053 (N_18053,N_17985,N_17802);
xor U18054 (N_18054,N_17938,N_17853);
or U18055 (N_18055,N_17975,N_17890);
nor U18056 (N_18056,N_17856,N_17879);
nand U18057 (N_18057,N_17813,N_17897);
or U18058 (N_18058,N_17838,N_17754);
nand U18059 (N_18059,N_17996,N_17769);
nor U18060 (N_18060,N_17980,N_17954);
and U18061 (N_18061,N_17871,N_17986);
nor U18062 (N_18062,N_17752,N_17815);
and U18063 (N_18063,N_17757,N_17847);
xnor U18064 (N_18064,N_17945,N_17929);
or U18065 (N_18065,N_17874,N_17833);
xor U18066 (N_18066,N_17964,N_17860);
nor U18067 (N_18067,N_17906,N_17951);
xnor U18068 (N_18068,N_17779,N_17908);
xor U18069 (N_18069,N_17969,N_17861);
and U18070 (N_18070,N_17998,N_17884);
xor U18071 (N_18071,N_17936,N_17780);
nor U18072 (N_18072,N_17823,N_17751);
nor U18073 (N_18073,N_17826,N_17835);
and U18074 (N_18074,N_17774,N_17958);
xor U18075 (N_18075,N_17787,N_17894);
and U18076 (N_18076,N_17941,N_17900);
nand U18077 (N_18077,N_17916,N_17800);
nor U18078 (N_18078,N_17914,N_17821);
and U18079 (N_18079,N_17880,N_17777);
nor U18080 (N_18080,N_17892,N_17972);
and U18081 (N_18081,N_17887,N_17756);
nor U18082 (N_18082,N_17935,N_17837);
nor U18083 (N_18083,N_17934,N_17903);
nor U18084 (N_18084,N_17895,N_17940);
and U18085 (N_18085,N_17781,N_17889);
nor U18086 (N_18086,N_17970,N_17901);
and U18087 (N_18087,N_17915,N_17882);
xor U18088 (N_18088,N_17834,N_17836);
nand U18089 (N_18089,N_17920,N_17992);
and U18090 (N_18090,N_17791,N_17775);
xor U18091 (N_18091,N_17962,N_17760);
and U18092 (N_18092,N_17988,N_17946);
nand U18093 (N_18093,N_17845,N_17971);
nand U18094 (N_18094,N_17788,N_17872);
or U18095 (N_18095,N_17849,N_17891);
xor U18096 (N_18096,N_17851,N_17842);
or U18097 (N_18097,N_17798,N_17810);
nor U18098 (N_18098,N_17910,N_17932);
and U18099 (N_18099,N_17807,N_17804);
xnor U18100 (N_18100,N_17925,N_17854);
and U18101 (N_18101,N_17928,N_17885);
xnor U18102 (N_18102,N_17801,N_17755);
xor U18103 (N_18103,N_17939,N_17949);
xnor U18104 (N_18104,N_17982,N_17832);
nand U18105 (N_18105,N_17773,N_17883);
nor U18106 (N_18106,N_17967,N_17857);
nand U18107 (N_18107,N_17993,N_17974);
and U18108 (N_18108,N_17877,N_17917);
or U18109 (N_18109,N_17966,N_17778);
and U18110 (N_18110,N_17947,N_17759);
nand U18111 (N_18111,N_17790,N_17786);
nor U18112 (N_18112,N_17827,N_17784);
xor U18113 (N_18113,N_17846,N_17994);
nor U18114 (N_18114,N_17957,N_17909);
or U18115 (N_18115,N_17850,N_17793);
and U18116 (N_18116,N_17811,N_17989);
and U18117 (N_18117,N_17855,N_17913);
nand U18118 (N_18118,N_17911,N_17792);
and U18119 (N_18119,N_17840,N_17899);
and U18120 (N_18120,N_17783,N_17896);
nor U18121 (N_18121,N_17950,N_17991);
and U18122 (N_18122,N_17922,N_17852);
nor U18123 (N_18123,N_17937,N_17763);
nor U18124 (N_18124,N_17960,N_17831);
xor U18125 (N_18125,N_17844,N_17999);
and U18126 (N_18126,N_17936,N_17915);
nand U18127 (N_18127,N_17988,N_17842);
nand U18128 (N_18128,N_17987,N_17943);
or U18129 (N_18129,N_17815,N_17755);
and U18130 (N_18130,N_17821,N_17942);
and U18131 (N_18131,N_17795,N_17861);
nand U18132 (N_18132,N_17790,N_17966);
xor U18133 (N_18133,N_17919,N_17856);
nand U18134 (N_18134,N_17909,N_17828);
nor U18135 (N_18135,N_17825,N_17791);
and U18136 (N_18136,N_17785,N_17921);
nor U18137 (N_18137,N_17793,N_17989);
xor U18138 (N_18138,N_17964,N_17951);
and U18139 (N_18139,N_17897,N_17923);
and U18140 (N_18140,N_17758,N_17885);
nor U18141 (N_18141,N_17767,N_17841);
and U18142 (N_18142,N_17857,N_17801);
or U18143 (N_18143,N_17903,N_17925);
nand U18144 (N_18144,N_17928,N_17786);
nand U18145 (N_18145,N_17874,N_17940);
and U18146 (N_18146,N_17850,N_17846);
and U18147 (N_18147,N_17934,N_17909);
nand U18148 (N_18148,N_17931,N_17798);
and U18149 (N_18149,N_17878,N_17794);
xor U18150 (N_18150,N_17946,N_17791);
nor U18151 (N_18151,N_17895,N_17951);
or U18152 (N_18152,N_17908,N_17764);
nand U18153 (N_18153,N_17766,N_17951);
nor U18154 (N_18154,N_17816,N_17906);
xnor U18155 (N_18155,N_17929,N_17843);
nand U18156 (N_18156,N_17965,N_17788);
xnor U18157 (N_18157,N_17901,N_17832);
and U18158 (N_18158,N_17872,N_17909);
nand U18159 (N_18159,N_17835,N_17765);
or U18160 (N_18160,N_17889,N_17934);
xnor U18161 (N_18161,N_17925,N_17849);
xor U18162 (N_18162,N_17815,N_17951);
xnor U18163 (N_18163,N_17881,N_17844);
xnor U18164 (N_18164,N_17909,N_17842);
and U18165 (N_18165,N_17965,N_17980);
nand U18166 (N_18166,N_17783,N_17754);
or U18167 (N_18167,N_17833,N_17751);
nand U18168 (N_18168,N_17920,N_17760);
nand U18169 (N_18169,N_17910,N_17963);
or U18170 (N_18170,N_17934,N_17812);
nor U18171 (N_18171,N_17853,N_17858);
xor U18172 (N_18172,N_17962,N_17953);
or U18173 (N_18173,N_17914,N_17860);
and U18174 (N_18174,N_17796,N_17847);
and U18175 (N_18175,N_17794,N_17886);
xor U18176 (N_18176,N_17998,N_17924);
and U18177 (N_18177,N_17819,N_17935);
or U18178 (N_18178,N_17911,N_17952);
xnor U18179 (N_18179,N_17861,N_17982);
or U18180 (N_18180,N_17972,N_17891);
nand U18181 (N_18181,N_17812,N_17887);
nor U18182 (N_18182,N_17963,N_17854);
xor U18183 (N_18183,N_17821,N_17874);
nor U18184 (N_18184,N_17785,N_17885);
nand U18185 (N_18185,N_17781,N_17843);
and U18186 (N_18186,N_17923,N_17859);
nor U18187 (N_18187,N_17957,N_17754);
or U18188 (N_18188,N_17909,N_17910);
and U18189 (N_18189,N_17756,N_17926);
nand U18190 (N_18190,N_17994,N_17993);
nand U18191 (N_18191,N_17988,N_17849);
and U18192 (N_18192,N_17822,N_17873);
or U18193 (N_18193,N_17776,N_17858);
or U18194 (N_18194,N_17782,N_17879);
nor U18195 (N_18195,N_17828,N_17910);
nor U18196 (N_18196,N_17780,N_17996);
or U18197 (N_18197,N_17849,N_17959);
or U18198 (N_18198,N_17783,N_17990);
nor U18199 (N_18199,N_17779,N_17942);
nand U18200 (N_18200,N_17978,N_17751);
nand U18201 (N_18201,N_17902,N_17805);
or U18202 (N_18202,N_17833,N_17828);
nand U18203 (N_18203,N_17937,N_17910);
xor U18204 (N_18204,N_17968,N_17839);
nand U18205 (N_18205,N_17791,N_17840);
xnor U18206 (N_18206,N_17948,N_17938);
and U18207 (N_18207,N_17818,N_17912);
and U18208 (N_18208,N_17943,N_17868);
xor U18209 (N_18209,N_17933,N_17887);
and U18210 (N_18210,N_17913,N_17951);
nor U18211 (N_18211,N_17984,N_17795);
or U18212 (N_18212,N_17875,N_17801);
nand U18213 (N_18213,N_17796,N_17771);
nor U18214 (N_18214,N_17923,N_17941);
or U18215 (N_18215,N_17861,N_17949);
nor U18216 (N_18216,N_17884,N_17811);
nor U18217 (N_18217,N_17850,N_17955);
xor U18218 (N_18218,N_17756,N_17905);
and U18219 (N_18219,N_17828,N_17776);
and U18220 (N_18220,N_17961,N_17958);
nor U18221 (N_18221,N_17981,N_17944);
nor U18222 (N_18222,N_17930,N_17859);
and U18223 (N_18223,N_17990,N_17805);
nor U18224 (N_18224,N_17880,N_17899);
nor U18225 (N_18225,N_17820,N_17979);
and U18226 (N_18226,N_17904,N_17880);
and U18227 (N_18227,N_17773,N_17866);
nor U18228 (N_18228,N_17815,N_17941);
or U18229 (N_18229,N_17882,N_17757);
nor U18230 (N_18230,N_17827,N_17865);
or U18231 (N_18231,N_17881,N_17930);
xnor U18232 (N_18232,N_17934,N_17777);
nor U18233 (N_18233,N_17807,N_17831);
nand U18234 (N_18234,N_17982,N_17768);
and U18235 (N_18235,N_17904,N_17813);
xor U18236 (N_18236,N_17914,N_17773);
or U18237 (N_18237,N_17800,N_17897);
nand U18238 (N_18238,N_17943,N_17778);
nand U18239 (N_18239,N_17876,N_17917);
nor U18240 (N_18240,N_17774,N_17771);
nor U18241 (N_18241,N_17960,N_17996);
nor U18242 (N_18242,N_17931,N_17855);
nor U18243 (N_18243,N_17835,N_17886);
nand U18244 (N_18244,N_17981,N_17789);
nand U18245 (N_18245,N_17951,N_17912);
nor U18246 (N_18246,N_17802,N_17946);
or U18247 (N_18247,N_17822,N_17939);
nand U18248 (N_18248,N_17907,N_17962);
xnor U18249 (N_18249,N_17779,N_17919);
xor U18250 (N_18250,N_18078,N_18032);
nor U18251 (N_18251,N_18178,N_18224);
nand U18252 (N_18252,N_18128,N_18160);
or U18253 (N_18253,N_18238,N_18096);
and U18254 (N_18254,N_18107,N_18126);
xor U18255 (N_18255,N_18081,N_18165);
and U18256 (N_18256,N_18120,N_18073);
xor U18257 (N_18257,N_18146,N_18004);
and U18258 (N_18258,N_18228,N_18136);
and U18259 (N_18259,N_18132,N_18024);
or U18260 (N_18260,N_18048,N_18155);
or U18261 (N_18261,N_18234,N_18069);
nand U18262 (N_18262,N_18091,N_18205);
nor U18263 (N_18263,N_18212,N_18051);
nor U18264 (N_18264,N_18058,N_18077);
or U18265 (N_18265,N_18116,N_18198);
xnor U18266 (N_18266,N_18030,N_18074);
nor U18267 (N_18267,N_18218,N_18233);
or U18268 (N_18268,N_18214,N_18072);
or U18269 (N_18269,N_18225,N_18002);
and U18270 (N_18270,N_18190,N_18129);
nand U18271 (N_18271,N_18040,N_18079);
and U18272 (N_18272,N_18035,N_18020);
or U18273 (N_18273,N_18008,N_18085);
xor U18274 (N_18274,N_18093,N_18098);
and U18275 (N_18275,N_18039,N_18204);
nor U18276 (N_18276,N_18210,N_18090);
or U18277 (N_18277,N_18123,N_18153);
nor U18278 (N_18278,N_18112,N_18017);
nor U18279 (N_18279,N_18015,N_18157);
nor U18280 (N_18280,N_18215,N_18118);
xor U18281 (N_18281,N_18247,N_18082);
nor U18282 (N_18282,N_18203,N_18038);
and U18283 (N_18283,N_18242,N_18168);
nor U18284 (N_18284,N_18025,N_18170);
nor U18285 (N_18285,N_18135,N_18150);
or U18286 (N_18286,N_18166,N_18036);
or U18287 (N_18287,N_18089,N_18070);
xnor U18288 (N_18288,N_18200,N_18092);
and U18289 (N_18289,N_18053,N_18076);
nor U18290 (N_18290,N_18059,N_18216);
xor U18291 (N_18291,N_18029,N_18137);
nor U18292 (N_18292,N_18026,N_18033);
xor U18293 (N_18293,N_18066,N_18018);
nor U18294 (N_18294,N_18134,N_18094);
nor U18295 (N_18295,N_18144,N_18006);
xor U18296 (N_18296,N_18188,N_18141);
xnor U18297 (N_18297,N_18248,N_18009);
xnor U18298 (N_18298,N_18211,N_18088);
xor U18299 (N_18299,N_18162,N_18050);
xor U18300 (N_18300,N_18163,N_18223);
nand U18301 (N_18301,N_18231,N_18156);
nand U18302 (N_18302,N_18192,N_18063);
nor U18303 (N_18303,N_18044,N_18100);
nor U18304 (N_18304,N_18229,N_18101);
nor U18305 (N_18305,N_18011,N_18060);
and U18306 (N_18306,N_18005,N_18171);
xnor U18307 (N_18307,N_18142,N_18226);
and U18308 (N_18308,N_18235,N_18182);
or U18309 (N_18309,N_18027,N_18122);
xor U18310 (N_18310,N_18167,N_18189);
nand U18311 (N_18311,N_18103,N_18186);
xor U18312 (N_18312,N_18151,N_18174);
xor U18313 (N_18313,N_18193,N_18217);
and U18314 (N_18314,N_18086,N_18158);
xnor U18315 (N_18315,N_18199,N_18043);
nand U18316 (N_18316,N_18220,N_18000);
xor U18317 (N_18317,N_18104,N_18102);
and U18318 (N_18318,N_18049,N_18194);
nand U18319 (N_18319,N_18133,N_18239);
nand U18320 (N_18320,N_18164,N_18196);
or U18321 (N_18321,N_18046,N_18111);
nor U18322 (N_18322,N_18007,N_18185);
and U18323 (N_18323,N_18014,N_18172);
and U18324 (N_18324,N_18175,N_18110);
xor U18325 (N_18325,N_18125,N_18045);
or U18326 (N_18326,N_18176,N_18019);
and U18327 (N_18327,N_18221,N_18031);
and U18328 (N_18328,N_18139,N_18083);
nor U18329 (N_18329,N_18159,N_18109);
xnor U18330 (N_18330,N_18201,N_18023);
xor U18331 (N_18331,N_18181,N_18084);
or U18332 (N_18332,N_18012,N_18010);
or U18333 (N_18333,N_18149,N_18061);
or U18334 (N_18334,N_18105,N_18071);
and U18335 (N_18335,N_18246,N_18057);
and U18336 (N_18336,N_18117,N_18237);
nor U18337 (N_18337,N_18209,N_18173);
and U18338 (N_18338,N_18245,N_18152);
or U18339 (N_18339,N_18068,N_18113);
and U18340 (N_18340,N_18042,N_18114);
xnor U18341 (N_18341,N_18003,N_18145);
nand U18342 (N_18342,N_18227,N_18064);
and U18343 (N_18343,N_18184,N_18016);
nor U18344 (N_18344,N_18127,N_18095);
or U18345 (N_18345,N_18041,N_18021);
and U18346 (N_18346,N_18197,N_18138);
or U18347 (N_18347,N_18001,N_18028);
nand U18348 (N_18348,N_18065,N_18206);
or U18349 (N_18349,N_18148,N_18037);
nand U18350 (N_18350,N_18187,N_18055);
or U18351 (N_18351,N_18236,N_18240);
or U18352 (N_18352,N_18080,N_18207);
or U18353 (N_18353,N_18232,N_18241);
or U18354 (N_18354,N_18244,N_18075);
nand U18355 (N_18355,N_18179,N_18230);
xor U18356 (N_18356,N_18121,N_18108);
or U18357 (N_18357,N_18034,N_18154);
nand U18358 (N_18358,N_18143,N_18131);
xnor U18359 (N_18359,N_18169,N_18243);
nor U18360 (N_18360,N_18161,N_18130);
nand U18361 (N_18361,N_18213,N_18124);
xnor U18362 (N_18362,N_18056,N_18219);
nor U18363 (N_18363,N_18222,N_18183);
or U18364 (N_18364,N_18249,N_18191);
xnor U18365 (N_18365,N_18087,N_18202);
and U18366 (N_18366,N_18115,N_18052);
nor U18367 (N_18367,N_18054,N_18147);
or U18368 (N_18368,N_18047,N_18067);
nand U18369 (N_18369,N_18062,N_18195);
or U18370 (N_18370,N_18180,N_18177);
xnor U18371 (N_18371,N_18119,N_18208);
nand U18372 (N_18372,N_18022,N_18140);
xnor U18373 (N_18373,N_18099,N_18106);
nor U18374 (N_18374,N_18097,N_18013);
and U18375 (N_18375,N_18105,N_18173);
nand U18376 (N_18376,N_18248,N_18034);
nand U18377 (N_18377,N_18006,N_18170);
nand U18378 (N_18378,N_18079,N_18085);
and U18379 (N_18379,N_18178,N_18155);
or U18380 (N_18380,N_18162,N_18097);
and U18381 (N_18381,N_18067,N_18184);
or U18382 (N_18382,N_18047,N_18240);
or U18383 (N_18383,N_18095,N_18212);
xor U18384 (N_18384,N_18218,N_18186);
and U18385 (N_18385,N_18218,N_18197);
xnor U18386 (N_18386,N_18001,N_18042);
and U18387 (N_18387,N_18152,N_18082);
nand U18388 (N_18388,N_18107,N_18071);
nor U18389 (N_18389,N_18100,N_18146);
or U18390 (N_18390,N_18169,N_18096);
nor U18391 (N_18391,N_18114,N_18162);
nor U18392 (N_18392,N_18168,N_18120);
xor U18393 (N_18393,N_18127,N_18225);
nand U18394 (N_18394,N_18084,N_18129);
nor U18395 (N_18395,N_18246,N_18169);
xnor U18396 (N_18396,N_18072,N_18076);
xor U18397 (N_18397,N_18099,N_18062);
or U18398 (N_18398,N_18188,N_18178);
nor U18399 (N_18399,N_18187,N_18172);
or U18400 (N_18400,N_18024,N_18146);
nor U18401 (N_18401,N_18020,N_18174);
nand U18402 (N_18402,N_18168,N_18140);
and U18403 (N_18403,N_18019,N_18025);
or U18404 (N_18404,N_18193,N_18107);
and U18405 (N_18405,N_18042,N_18168);
nand U18406 (N_18406,N_18067,N_18065);
nor U18407 (N_18407,N_18148,N_18216);
xnor U18408 (N_18408,N_18249,N_18100);
nor U18409 (N_18409,N_18158,N_18149);
nor U18410 (N_18410,N_18007,N_18118);
nor U18411 (N_18411,N_18248,N_18056);
xor U18412 (N_18412,N_18224,N_18021);
xnor U18413 (N_18413,N_18206,N_18036);
nand U18414 (N_18414,N_18005,N_18230);
or U18415 (N_18415,N_18075,N_18173);
or U18416 (N_18416,N_18089,N_18119);
xnor U18417 (N_18417,N_18116,N_18234);
nand U18418 (N_18418,N_18069,N_18018);
nand U18419 (N_18419,N_18056,N_18051);
or U18420 (N_18420,N_18060,N_18219);
nor U18421 (N_18421,N_18090,N_18156);
nor U18422 (N_18422,N_18002,N_18178);
or U18423 (N_18423,N_18072,N_18078);
nor U18424 (N_18424,N_18029,N_18002);
nand U18425 (N_18425,N_18005,N_18065);
and U18426 (N_18426,N_18221,N_18198);
nor U18427 (N_18427,N_18244,N_18127);
nor U18428 (N_18428,N_18099,N_18173);
or U18429 (N_18429,N_18024,N_18162);
nor U18430 (N_18430,N_18202,N_18051);
nor U18431 (N_18431,N_18072,N_18168);
and U18432 (N_18432,N_18221,N_18086);
xor U18433 (N_18433,N_18074,N_18021);
or U18434 (N_18434,N_18190,N_18097);
xor U18435 (N_18435,N_18189,N_18003);
xnor U18436 (N_18436,N_18064,N_18245);
and U18437 (N_18437,N_18046,N_18155);
nor U18438 (N_18438,N_18102,N_18223);
nand U18439 (N_18439,N_18147,N_18135);
nand U18440 (N_18440,N_18134,N_18239);
nor U18441 (N_18441,N_18042,N_18206);
xor U18442 (N_18442,N_18000,N_18041);
nor U18443 (N_18443,N_18230,N_18232);
nand U18444 (N_18444,N_18045,N_18248);
or U18445 (N_18445,N_18014,N_18104);
xor U18446 (N_18446,N_18121,N_18103);
nor U18447 (N_18447,N_18170,N_18237);
xor U18448 (N_18448,N_18076,N_18174);
nor U18449 (N_18449,N_18065,N_18242);
or U18450 (N_18450,N_18091,N_18126);
nor U18451 (N_18451,N_18151,N_18047);
nor U18452 (N_18452,N_18049,N_18096);
xnor U18453 (N_18453,N_18034,N_18227);
nor U18454 (N_18454,N_18157,N_18120);
nand U18455 (N_18455,N_18179,N_18224);
nor U18456 (N_18456,N_18146,N_18143);
xnor U18457 (N_18457,N_18125,N_18200);
and U18458 (N_18458,N_18125,N_18236);
and U18459 (N_18459,N_18128,N_18110);
xor U18460 (N_18460,N_18144,N_18058);
xnor U18461 (N_18461,N_18216,N_18093);
nor U18462 (N_18462,N_18068,N_18175);
or U18463 (N_18463,N_18223,N_18169);
nand U18464 (N_18464,N_18026,N_18204);
xnor U18465 (N_18465,N_18121,N_18030);
and U18466 (N_18466,N_18213,N_18047);
nand U18467 (N_18467,N_18028,N_18086);
nand U18468 (N_18468,N_18189,N_18078);
xnor U18469 (N_18469,N_18243,N_18172);
and U18470 (N_18470,N_18054,N_18191);
or U18471 (N_18471,N_18110,N_18103);
xor U18472 (N_18472,N_18166,N_18022);
xnor U18473 (N_18473,N_18199,N_18070);
xnor U18474 (N_18474,N_18111,N_18177);
xor U18475 (N_18475,N_18109,N_18157);
nand U18476 (N_18476,N_18108,N_18177);
xnor U18477 (N_18477,N_18243,N_18205);
or U18478 (N_18478,N_18053,N_18110);
and U18479 (N_18479,N_18234,N_18172);
and U18480 (N_18480,N_18223,N_18108);
and U18481 (N_18481,N_18207,N_18222);
or U18482 (N_18482,N_18238,N_18002);
xnor U18483 (N_18483,N_18062,N_18053);
nor U18484 (N_18484,N_18071,N_18119);
nor U18485 (N_18485,N_18217,N_18132);
or U18486 (N_18486,N_18115,N_18073);
nand U18487 (N_18487,N_18165,N_18062);
nor U18488 (N_18488,N_18129,N_18249);
nor U18489 (N_18489,N_18027,N_18133);
nor U18490 (N_18490,N_18045,N_18220);
xnor U18491 (N_18491,N_18223,N_18089);
nor U18492 (N_18492,N_18122,N_18059);
or U18493 (N_18493,N_18133,N_18215);
nor U18494 (N_18494,N_18084,N_18106);
and U18495 (N_18495,N_18053,N_18008);
xnor U18496 (N_18496,N_18123,N_18219);
and U18497 (N_18497,N_18179,N_18163);
or U18498 (N_18498,N_18044,N_18065);
or U18499 (N_18499,N_18212,N_18115);
and U18500 (N_18500,N_18391,N_18363);
xor U18501 (N_18501,N_18464,N_18279);
nand U18502 (N_18502,N_18463,N_18474);
or U18503 (N_18503,N_18488,N_18297);
or U18504 (N_18504,N_18291,N_18361);
nand U18505 (N_18505,N_18389,N_18341);
xnor U18506 (N_18506,N_18357,N_18415);
nor U18507 (N_18507,N_18368,N_18430);
nor U18508 (N_18508,N_18328,N_18253);
nor U18509 (N_18509,N_18344,N_18492);
xnor U18510 (N_18510,N_18425,N_18440);
nor U18511 (N_18511,N_18252,N_18472);
and U18512 (N_18512,N_18358,N_18412);
xnor U18513 (N_18513,N_18446,N_18434);
and U18514 (N_18514,N_18406,N_18285);
or U18515 (N_18515,N_18410,N_18311);
xor U18516 (N_18516,N_18480,N_18481);
or U18517 (N_18517,N_18272,N_18382);
xnor U18518 (N_18518,N_18306,N_18466);
nor U18519 (N_18519,N_18438,N_18427);
or U18520 (N_18520,N_18444,N_18264);
nor U18521 (N_18521,N_18373,N_18342);
nor U18522 (N_18522,N_18270,N_18288);
or U18523 (N_18523,N_18477,N_18448);
or U18524 (N_18524,N_18330,N_18309);
nand U18525 (N_18525,N_18354,N_18433);
nor U18526 (N_18526,N_18296,N_18281);
nand U18527 (N_18527,N_18257,N_18413);
and U18528 (N_18528,N_18365,N_18303);
xnor U18529 (N_18529,N_18317,N_18258);
nor U18530 (N_18530,N_18462,N_18323);
nand U18531 (N_18531,N_18471,N_18426);
nor U18532 (N_18532,N_18315,N_18407);
nand U18533 (N_18533,N_18287,N_18429);
nand U18534 (N_18534,N_18326,N_18443);
or U18535 (N_18535,N_18305,N_18316);
or U18536 (N_18536,N_18355,N_18333);
and U18537 (N_18537,N_18467,N_18352);
or U18538 (N_18538,N_18479,N_18439);
and U18539 (N_18539,N_18353,N_18489);
nand U18540 (N_18540,N_18400,N_18418);
xor U18541 (N_18541,N_18451,N_18402);
xnor U18542 (N_18542,N_18308,N_18304);
nor U18543 (N_18543,N_18293,N_18367);
and U18544 (N_18544,N_18284,N_18310);
or U18545 (N_18545,N_18454,N_18324);
and U18546 (N_18546,N_18384,N_18445);
xnor U18547 (N_18547,N_18322,N_18436);
and U18548 (N_18548,N_18453,N_18460);
nor U18549 (N_18549,N_18499,N_18290);
nand U18550 (N_18550,N_18286,N_18314);
nor U18551 (N_18551,N_18278,N_18419);
and U18552 (N_18552,N_18461,N_18449);
and U18553 (N_18553,N_18485,N_18263);
nand U18554 (N_18554,N_18274,N_18280);
xnor U18555 (N_18555,N_18267,N_18331);
nand U18556 (N_18556,N_18478,N_18476);
and U18557 (N_18557,N_18452,N_18457);
nand U18558 (N_18558,N_18404,N_18401);
and U18559 (N_18559,N_18473,N_18374);
nand U18560 (N_18560,N_18254,N_18386);
and U18561 (N_18561,N_18298,N_18256);
nand U18562 (N_18562,N_18428,N_18356);
nand U18563 (N_18563,N_18276,N_18339);
xor U18564 (N_18564,N_18340,N_18362);
or U18565 (N_18565,N_18343,N_18295);
and U18566 (N_18566,N_18292,N_18403);
nand U18567 (N_18567,N_18302,N_18447);
xor U18568 (N_18568,N_18470,N_18366);
nor U18569 (N_18569,N_18456,N_18486);
nand U18570 (N_18570,N_18307,N_18450);
or U18571 (N_18571,N_18487,N_18411);
and U18572 (N_18572,N_18251,N_18318);
and U18573 (N_18573,N_18385,N_18498);
nand U18574 (N_18574,N_18469,N_18369);
or U18575 (N_18575,N_18283,N_18377);
xor U18576 (N_18576,N_18493,N_18387);
nor U18577 (N_18577,N_18437,N_18268);
xor U18578 (N_18578,N_18259,N_18379);
nor U18579 (N_18579,N_18392,N_18458);
or U18580 (N_18580,N_18408,N_18334);
xor U18581 (N_18581,N_18266,N_18261);
and U18582 (N_18582,N_18465,N_18442);
nand U18583 (N_18583,N_18347,N_18380);
and U18584 (N_18584,N_18475,N_18299);
and U18585 (N_18585,N_18255,N_18350);
xor U18586 (N_18586,N_18398,N_18381);
nor U18587 (N_18587,N_18420,N_18395);
and U18588 (N_18588,N_18273,N_18338);
or U18589 (N_18589,N_18277,N_18482);
xnor U18590 (N_18590,N_18289,N_18441);
and U18591 (N_18591,N_18271,N_18275);
and U18592 (N_18592,N_18496,N_18431);
or U18593 (N_18593,N_18390,N_18250);
and U18594 (N_18594,N_18397,N_18300);
and U18595 (N_18595,N_18459,N_18378);
and U18596 (N_18596,N_18265,N_18327);
xor U18597 (N_18597,N_18360,N_18320);
xor U18598 (N_18598,N_18346,N_18269);
xnor U18599 (N_18599,N_18325,N_18332);
or U18600 (N_18600,N_18371,N_18494);
nand U18601 (N_18601,N_18484,N_18421);
and U18602 (N_18602,N_18497,N_18370);
xnor U18603 (N_18603,N_18455,N_18336);
nor U18604 (N_18604,N_18348,N_18491);
xor U18605 (N_18605,N_18383,N_18282);
xor U18606 (N_18606,N_18393,N_18416);
nor U18607 (N_18607,N_18337,N_18409);
nand U18608 (N_18608,N_18423,N_18399);
or U18609 (N_18609,N_18313,N_18376);
nor U18610 (N_18610,N_18319,N_18301);
xor U18611 (N_18611,N_18435,N_18483);
or U18612 (N_18612,N_18364,N_18345);
and U18613 (N_18613,N_18351,N_18495);
nor U18614 (N_18614,N_18424,N_18260);
or U18615 (N_18615,N_18359,N_18396);
nor U18616 (N_18616,N_18335,N_18375);
nor U18617 (N_18617,N_18394,N_18432);
or U18618 (N_18618,N_18312,N_18422);
and U18619 (N_18619,N_18405,N_18468);
and U18620 (N_18620,N_18329,N_18372);
or U18621 (N_18621,N_18417,N_18388);
xor U18622 (N_18622,N_18321,N_18262);
xnor U18623 (N_18623,N_18294,N_18490);
or U18624 (N_18624,N_18414,N_18349);
or U18625 (N_18625,N_18370,N_18426);
and U18626 (N_18626,N_18359,N_18356);
and U18627 (N_18627,N_18305,N_18477);
nand U18628 (N_18628,N_18275,N_18313);
xnor U18629 (N_18629,N_18472,N_18373);
nor U18630 (N_18630,N_18288,N_18475);
xnor U18631 (N_18631,N_18364,N_18449);
nand U18632 (N_18632,N_18417,N_18343);
nand U18633 (N_18633,N_18498,N_18432);
nand U18634 (N_18634,N_18278,N_18326);
and U18635 (N_18635,N_18289,N_18464);
or U18636 (N_18636,N_18294,N_18463);
nand U18637 (N_18637,N_18287,N_18326);
nor U18638 (N_18638,N_18323,N_18357);
and U18639 (N_18639,N_18334,N_18447);
nand U18640 (N_18640,N_18379,N_18450);
or U18641 (N_18641,N_18308,N_18314);
nand U18642 (N_18642,N_18263,N_18471);
and U18643 (N_18643,N_18377,N_18455);
or U18644 (N_18644,N_18349,N_18254);
nor U18645 (N_18645,N_18391,N_18454);
and U18646 (N_18646,N_18323,N_18451);
and U18647 (N_18647,N_18451,N_18399);
xnor U18648 (N_18648,N_18284,N_18360);
nor U18649 (N_18649,N_18434,N_18415);
xor U18650 (N_18650,N_18450,N_18429);
nand U18651 (N_18651,N_18470,N_18266);
or U18652 (N_18652,N_18435,N_18334);
nand U18653 (N_18653,N_18378,N_18256);
xor U18654 (N_18654,N_18397,N_18380);
and U18655 (N_18655,N_18374,N_18322);
and U18656 (N_18656,N_18447,N_18430);
and U18657 (N_18657,N_18398,N_18323);
nor U18658 (N_18658,N_18410,N_18360);
nand U18659 (N_18659,N_18299,N_18326);
nand U18660 (N_18660,N_18314,N_18427);
nand U18661 (N_18661,N_18413,N_18314);
xnor U18662 (N_18662,N_18431,N_18284);
xnor U18663 (N_18663,N_18452,N_18495);
and U18664 (N_18664,N_18359,N_18292);
and U18665 (N_18665,N_18443,N_18415);
and U18666 (N_18666,N_18370,N_18374);
and U18667 (N_18667,N_18490,N_18482);
and U18668 (N_18668,N_18316,N_18487);
nand U18669 (N_18669,N_18366,N_18393);
nor U18670 (N_18670,N_18452,N_18496);
nand U18671 (N_18671,N_18454,N_18434);
and U18672 (N_18672,N_18452,N_18433);
and U18673 (N_18673,N_18258,N_18455);
nor U18674 (N_18674,N_18295,N_18321);
or U18675 (N_18675,N_18312,N_18470);
nand U18676 (N_18676,N_18372,N_18361);
nor U18677 (N_18677,N_18433,N_18268);
nand U18678 (N_18678,N_18337,N_18305);
or U18679 (N_18679,N_18494,N_18324);
and U18680 (N_18680,N_18275,N_18496);
xnor U18681 (N_18681,N_18268,N_18272);
and U18682 (N_18682,N_18467,N_18466);
xnor U18683 (N_18683,N_18453,N_18347);
nor U18684 (N_18684,N_18281,N_18331);
or U18685 (N_18685,N_18355,N_18405);
xnor U18686 (N_18686,N_18366,N_18461);
nor U18687 (N_18687,N_18317,N_18409);
nor U18688 (N_18688,N_18421,N_18416);
nand U18689 (N_18689,N_18405,N_18492);
xnor U18690 (N_18690,N_18363,N_18336);
xnor U18691 (N_18691,N_18379,N_18448);
xor U18692 (N_18692,N_18460,N_18410);
and U18693 (N_18693,N_18366,N_18262);
or U18694 (N_18694,N_18265,N_18483);
nand U18695 (N_18695,N_18258,N_18413);
or U18696 (N_18696,N_18441,N_18280);
nor U18697 (N_18697,N_18329,N_18484);
nand U18698 (N_18698,N_18309,N_18279);
nand U18699 (N_18699,N_18334,N_18305);
xor U18700 (N_18700,N_18349,N_18289);
and U18701 (N_18701,N_18270,N_18418);
or U18702 (N_18702,N_18384,N_18480);
xnor U18703 (N_18703,N_18381,N_18349);
xnor U18704 (N_18704,N_18428,N_18368);
or U18705 (N_18705,N_18464,N_18488);
nor U18706 (N_18706,N_18423,N_18462);
and U18707 (N_18707,N_18296,N_18492);
or U18708 (N_18708,N_18312,N_18328);
or U18709 (N_18709,N_18356,N_18388);
and U18710 (N_18710,N_18493,N_18276);
nand U18711 (N_18711,N_18482,N_18291);
xnor U18712 (N_18712,N_18476,N_18351);
nand U18713 (N_18713,N_18444,N_18252);
and U18714 (N_18714,N_18295,N_18274);
and U18715 (N_18715,N_18415,N_18350);
and U18716 (N_18716,N_18267,N_18464);
or U18717 (N_18717,N_18261,N_18461);
and U18718 (N_18718,N_18444,N_18401);
xnor U18719 (N_18719,N_18463,N_18492);
and U18720 (N_18720,N_18349,N_18288);
nor U18721 (N_18721,N_18311,N_18297);
xor U18722 (N_18722,N_18357,N_18280);
xor U18723 (N_18723,N_18315,N_18259);
nand U18724 (N_18724,N_18460,N_18449);
nand U18725 (N_18725,N_18353,N_18430);
xnor U18726 (N_18726,N_18405,N_18497);
or U18727 (N_18727,N_18301,N_18382);
nor U18728 (N_18728,N_18427,N_18259);
xor U18729 (N_18729,N_18455,N_18263);
and U18730 (N_18730,N_18488,N_18469);
and U18731 (N_18731,N_18498,N_18451);
xor U18732 (N_18732,N_18403,N_18429);
nor U18733 (N_18733,N_18341,N_18462);
nand U18734 (N_18734,N_18304,N_18432);
nand U18735 (N_18735,N_18463,N_18348);
nand U18736 (N_18736,N_18451,N_18459);
nor U18737 (N_18737,N_18293,N_18306);
nand U18738 (N_18738,N_18283,N_18254);
nor U18739 (N_18739,N_18434,N_18394);
nand U18740 (N_18740,N_18442,N_18437);
nand U18741 (N_18741,N_18263,N_18397);
and U18742 (N_18742,N_18316,N_18455);
nor U18743 (N_18743,N_18492,N_18481);
nand U18744 (N_18744,N_18408,N_18423);
xnor U18745 (N_18745,N_18436,N_18351);
nor U18746 (N_18746,N_18278,N_18271);
and U18747 (N_18747,N_18264,N_18302);
or U18748 (N_18748,N_18321,N_18329);
xor U18749 (N_18749,N_18276,N_18285);
xor U18750 (N_18750,N_18687,N_18541);
nand U18751 (N_18751,N_18633,N_18699);
nor U18752 (N_18752,N_18675,N_18516);
nand U18753 (N_18753,N_18522,N_18593);
nand U18754 (N_18754,N_18502,N_18707);
xnor U18755 (N_18755,N_18603,N_18583);
nand U18756 (N_18756,N_18734,N_18706);
and U18757 (N_18757,N_18591,N_18665);
nor U18758 (N_18758,N_18692,N_18544);
or U18759 (N_18759,N_18517,N_18681);
and U18760 (N_18760,N_18504,N_18555);
nor U18761 (N_18761,N_18545,N_18535);
xnor U18762 (N_18762,N_18639,N_18536);
xnor U18763 (N_18763,N_18712,N_18612);
or U18764 (N_18764,N_18745,N_18710);
nand U18765 (N_18765,N_18589,N_18653);
and U18766 (N_18766,N_18610,N_18747);
nor U18767 (N_18767,N_18521,N_18598);
and U18768 (N_18768,N_18514,N_18608);
nand U18769 (N_18769,N_18520,N_18671);
xnor U18770 (N_18770,N_18667,N_18731);
nor U18771 (N_18771,N_18732,N_18556);
and U18772 (N_18772,N_18640,N_18718);
nand U18773 (N_18773,N_18508,N_18743);
and U18774 (N_18774,N_18525,N_18550);
nand U18775 (N_18775,N_18519,N_18558);
and U18776 (N_18776,N_18597,N_18664);
and U18777 (N_18777,N_18551,N_18630);
and U18778 (N_18778,N_18552,N_18509);
nand U18779 (N_18779,N_18636,N_18742);
or U18780 (N_18780,N_18601,N_18625);
nor U18781 (N_18781,N_18627,N_18678);
xnor U18782 (N_18782,N_18562,N_18580);
xnor U18783 (N_18783,N_18534,N_18657);
nand U18784 (N_18784,N_18703,N_18565);
nand U18785 (N_18785,N_18513,N_18631);
nand U18786 (N_18786,N_18568,N_18663);
nor U18787 (N_18787,N_18694,N_18669);
and U18788 (N_18788,N_18547,N_18649);
or U18789 (N_18789,N_18739,N_18507);
xor U18790 (N_18790,N_18614,N_18559);
and U18791 (N_18791,N_18590,N_18740);
xnor U18792 (N_18792,N_18658,N_18646);
nand U18793 (N_18793,N_18634,N_18730);
xnor U18794 (N_18794,N_18673,N_18652);
or U18795 (N_18795,N_18683,N_18680);
xor U18796 (N_18796,N_18584,N_18713);
nand U18797 (N_18797,N_18659,N_18503);
nor U18798 (N_18798,N_18617,N_18599);
and U18799 (N_18799,N_18549,N_18576);
nand U18800 (N_18800,N_18575,N_18626);
nor U18801 (N_18801,N_18729,N_18564);
xor U18802 (N_18802,N_18684,N_18577);
or U18803 (N_18803,N_18648,N_18749);
nor U18804 (N_18804,N_18645,N_18725);
nand U18805 (N_18805,N_18720,N_18723);
nand U18806 (N_18806,N_18661,N_18537);
nand U18807 (N_18807,N_18515,N_18524);
and U18808 (N_18808,N_18727,N_18668);
nor U18809 (N_18809,N_18709,N_18691);
nand U18810 (N_18810,N_18643,N_18543);
and U18811 (N_18811,N_18682,N_18721);
nand U18812 (N_18812,N_18676,N_18578);
or U18813 (N_18813,N_18567,N_18621);
xor U18814 (N_18814,N_18728,N_18670);
nor U18815 (N_18815,N_18573,N_18604);
nor U18816 (N_18816,N_18609,N_18736);
nand U18817 (N_18817,N_18744,N_18554);
nor U18818 (N_18818,N_18719,N_18587);
and U18819 (N_18819,N_18585,N_18606);
or U18820 (N_18820,N_18654,N_18700);
nor U18821 (N_18821,N_18532,N_18655);
or U18822 (N_18822,N_18748,N_18738);
nand U18823 (N_18823,N_18602,N_18644);
nor U18824 (N_18824,N_18571,N_18641);
nand U18825 (N_18825,N_18560,N_18624);
or U18826 (N_18826,N_18701,N_18530);
nor U18827 (N_18827,N_18638,N_18500);
xor U18828 (N_18828,N_18656,N_18588);
nor U18829 (N_18829,N_18501,N_18613);
nand U18830 (N_18830,N_18733,N_18528);
nor U18831 (N_18831,N_18662,N_18622);
xnor U18832 (N_18832,N_18629,N_18632);
or U18833 (N_18833,N_18569,N_18726);
nand U18834 (N_18834,N_18505,N_18529);
nor U18835 (N_18835,N_18595,N_18582);
xnor U18836 (N_18836,N_18563,N_18735);
nand U18837 (N_18837,N_18581,N_18695);
and U18838 (N_18838,N_18533,N_18600);
and U18839 (N_18839,N_18538,N_18523);
and U18840 (N_18840,N_18708,N_18566);
nor U18841 (N_18841,N_18542,N_18686);
nand U18842 (N_18842,N_18650,N_18510);
or U18843 (N_18843,N_18572,N_18539);
nand U18844 (N_18844,N_18637,N_18557);
xnor U18845 (N_18845,N_18527,N_18619);
nor U18846 (N_18846,N_18689,N_18690);
nand U18847 (N_18847,N_18574,N_18628);
xnor U18848 (N_18848,N_18561,N_18746);
and U18849 (N_18849,N_18697,N_18586);
and U18850 (N_18850,N_18616,N_18531);
and U18851 (N_18851,N_18620,N_18715);
nor U18852 (N_18852,N_18685,N_18579);
nand U18853 (N_18853,N_18666,N_18696);
nand U18854 (N_18854,N_18506,N_18651);
xnor U18855 (N_18855,N_18512,N_18672);
nand U18856 (N_18856,N_18594,N_18688);
nor U18857 (N_18857,N_18553,N_18693);
or U18858 (N_18858,N_18526,N_18518);
and U18859 (N_18859,N_18679,N_18618);
nand U18860 (N_18860,N_18540,N_18741);
nor U18861 (N_18861,N_18511,N_18605);
xor U18862 (N_18862,N_18737,N_18722);
nand U18863 (N_18863,N_18635,N_18716);
or U18864 (N_18864,N_18570,N_18677);
and U18865 (N_18865,N_18611,N_18704);
xnor U18866 (N_18866,N_18647,N_18711);
nor U18867 (N_18867,N_18705,N_18698);
and U18868 (N_18868,N_18714,N_18623);
or U18869 (N_18869,N_18596,N_18607);
nor U18870 (N_18870,N_18724,N_18702);
or U18871 (N_18871,N_18674,N_18660);
and U18872 (N_18872,N_18592,N_18548);
nand U18873 (N_18873,N_18546,N_18615);
and U18874 (N_18874,N_18717,N_18642);
xor U18875 (N_18875,N_18515,N_18570);
xnor U18876 (N_18876,N_18558,N_18660);
nand U18877 (N_18877,N_18748,N_18650);
xor U18878 (N_18878,N_18676,N_18555);
or U18879 (N_18879,N_18568,N_18514);
and U18880 (N_18880,N_18591,N_18506);
or U18881 (N_18881,N_18654,N_18723);
xnor U18882 (N_18882,N_18579,N_18514);
and U18883 (N_18883,N_18661,N_18621);
nand U18884 (N_18884,N_18656,N_18747);
nor U18885 (N_18885,N_18528,N_18697);
nand U18886 (N_18886,N_18553,N_18584);
and U18887 (N_18887,N_18590,N_18687);
xnor U18888 (N_18888,N_18534,N_18546);
and U18889 (N_18889,N_18548,N_18728);
nand U18890 (N_18890,N_18628,N_18719);
and U18891 (N_18891,N_18544,N_18550);
nor U18892 (N_18892,N_18582,N_18561);
nand U18893 (N_18893,N_18723,N_18656);
or U18894 (N_18894,N_18702,N_18501);
or U18895 (N_18895,N_18596,N_18610);
nand U18896 (N_18896,N_18608,N_18642);
or U18897 (N_18897,N_18623,N_18520);
xnor U18898 (N_18898,N_18684,N_18551);
nor U18899 (N_18899,N_18567,N_18706);
or U18900 (N_18900,N_18599,N_18639);
or U18901 (N_18901,N_18620,N_18678);
nand U18902 (N_18902,N_18650,N_18531);
nor U18903 (N_18903,N_18514,N_18720);
or U18904 (N_18904,N_18650,N_18553);
and U18905 (N_18905,N_18538,N_18625);
or U18906 (N_18906,N_18652,N_18545);
and U18907 (N_18907,N_18742,N_18547);
nand U18908 (N_18908,N_18680,N_18642);
xor U18909 (N_18909,N_18579,N_18580);
nand U18910 (N_18910,N_18633,N_18728);
nor U18911 (N_18911,N_18736,N_18634);
nand U18912 (N_18912,N_18740,N_18596);
nor U18913 (N_18913,N_18614,N_18543);
xor U18914 (N_18914,N_18628,N_18582);
nor U18915 (N_18915,N_18637,N_18591);
nand U18916 (N_18916,N_18697,N_18618);
nand U18917 (N_18917,N_18553,N_18637);
nor U18918 (N_18918,N_18553,N_18705);
nor U18919 (N_18919,N_18513,N_18671);
and U18920 (N_18920,N_18554,N_18579);
nor U18921 (N_18921,N_18631,N_18636);
nor U18922 (N_18922,N_18628,N_18696);
or U18923 (N_18923,N_18697,N_18659);
nand U18924 (N_18924,N_18640,N_18589);
or U18925 (N_18925,N_18676,N_18660);
nor U18926 (N_18926,N_18527,N_18502);
and U18927 (N_18927,N_18581,N_18506);
xor U18928 (N_18928,N_18538,N_18723);
xor U18929 (N_18929,N_18614,N_18671);
xor U18930 (N_18930,N_18727,N_18720);
or U18931 (N_18931,N_18542,N_18720);
nand U18932 (N_18932,N_18574,N_18708);
or U18933 (N_18933,N_18543,N_18541);
nand U18934 (N_18934,N_18725,N_18522);
nand U18935 (N_18935,N_18625,N_18633);
or U18936 (N_18936,N_18593,N_18667);
xor U18937 (N_18937,N_18557,N_18709);
nand U18938 (N_18938,N_18580,N_18631);
or U18939 (N_18939,N_18539,N_18557);
nor U18940 (N_18940,N_18602,N_18507);
nand U18941 (N_18941,N_18640,N_18633);
nand U18942 (N_18942,N_18692,N_18682);
or U18943 (N_18943,N_18659,N_18663);
nor U18944 (N_18944,N_18622,N_18668);
nand U18945 (N_18945,N_18696,N_18715);
or U18946 (N_18946,N_18553,N_18704);
nand U18947 (N_18947,N_18536,N_18573);
nand U18948 (N_18948,N_18569,N_18596);
nand U18949 (N_18949,N_18557,N_18661);
xor U18950 (N_18950,N_18645,N_18723);
xnor U18951 (N_18951,N_18714,N_18718);
xor U18952 (N_18952,N_18662,N_18744);
nor U18953 (N_18953,N_18657,N_18636);
nor U18954 (N_18954,N_18537,N_18612);
xnor U18955 (N_18955,N_18730,N_18676);
nor U18956 (N_18956,N_18674,N_18713);
or U18957 (N_18957,N_18691,N_18657);
nor U18958 (N_18958,N_18740,N_18619);
xnor U18959 (N_18959,N_18727,N_18552);
nor U18960 (N_18960,N_18622,N_18707);
or U18961 (N_18961,N_18701,N_18512);
or U18962 (N_18962,N_18569,N_18636);
and U18963 (N_18963,N_18594,N_18506);
or U18964 (N_18964,N_18545,N_18557);
or U18965 (N_18965,N_18701,N_18541);
or U18966 (N_18966,N_18625,N_18726);
nand U18967 (N_18967,N_18521,N_18740);
nand U18968 (N_18968,N_18743,N_18559);
nor U18969 (N_18969,N_18747,N_18664);
nor U18970 (N_18970,N_18637,N_18639);
nor U18971 (N_18971,N_18646,N_18704);
nor U18972 (N_18972,N_18602,N_18604);
or U18973 (N_18973,N_18660,N_18574);
or U18974 (N_18974,N_18660,N_18695);
nand U18975 (N_18975,N_18602,N_18509);
xnor U18976 (N_18976,N_18503,N_18741);
nor U18977 (N_18977,N_18704,N_18614);
or U18978 (N_18978,N_18654,N_18533);
nor U18979 (N_18979,N_18526,N_18502);
and U18980 (N_18980,N_18578,N_18605);
nand U18981 (N_18981,N_18720,N_18593);
and U18982 (N_18982,N_18548,N_18520);
nor U18983 (N_18983,N_18623,N_18668);
xnor U18984 (N_18984,N_18613,N_18668);
nand U18985 (N_18985,N_18673,N_18507);
nor U18986 (N_18986,N_18690,N_18745);
nand U18987 (N_18987,N_18718,N_18726);
nand U18988 (N_18988,N_18602,N_18603);
xnor U18989 (N_18989,N_18728,N_18704);
and U18990 (N_18990,N_18584,N_18528);
xnor U18991 (N_18991,N_18721,N_18669);
or U18992 (N_18992,N_18566,N_18633);
and U18993 (N_18993,N_18640,N_18684);
and U18994 (N_18994,N_18690,N_18705);
nand U18995 (N_18995,N_18564,N_18552);
xor U18996 (N_18996,N_18711,N_18673);
or U18997 (N_18997,N_18658,N_18557);
or U18998 (N_18998,N_18619,N_18575);
nand U18999 (N_18999,N_18726,N_18695);
and U19000 (N_19000,N_18880,N_18761);
nand U19001 (N_19001,N_18895,N_18923);
and U19002 (N_19002,N_18860,N_18821);
and U19003 (N_19003,N_18938,N_18990);
xor U19004 (N_19004,N_18908,N_18898);
nand U19005 (N_19005,N_18809,N_18874);
nand U19006 (N_19006,N_18885,N_18919);
xor U19007 (N_19007,N_18765,N_18762);
xor U19008 (N_19008,N_18995,N_18883);
nor U19009 (N_19009,N_18818,N_18858);
and U19010 (N_19010,N_18778,N_18933);
or U19011 (N_19011,N_18960,N_18848);
and U19012 (N_19012,N_18944,N_18943);
or U19013 (N_19013,N_18962,N_18920);
xor U19014 (N_19014,N_18914,N_18915);
xnor U19015 (N_19015,N_18779,N_18911);
or U19016 (N_19016,N_18966,N_18863);
and U19017 (N_19017,N_18783,N_18992);
nand U19018 (N_19018,N_18973,N_18887);
nand U19019 (N_19019,N_18849,N_18822);
nand U19020 (N_19020,N_18906,N_18934);
or U19021 (N_19021,N_18871,N_18951);
and U19022 (N_19022,N_18835,N_18803);
xnor U19023 (N_19023,N_18903,N_18800);
nand U19024 (N_19024,N_18791,N_18836);
xor U19025 (N_19025,N_18958,N_18928);
and U19026 (N_19026,N_18987,N_18983);
xnor U19027 (N_19027,N_18812,N_18805);
or U19028 (N_19028,N_18961,N_18917);
or U19029 (N_19029,N_18769,N_18853);
or U19030 (N_19030,N_18937,N_18784);
xor U19031 (N_19031,N_18774,N_18757);
xor U19032 (N_19032,N_18855,N_18793);
nand U19033 (N_19033,N_18820,N_18845);
nand U19034 (N_19034,N_18879,N_18940);
or U19035 (N_19035,N_18891,N_18806);
and U19036 (N_19036,N_18974,N_18894);
or U19037 (N_19037,N_18807,N_18816);
nor U19038 (N_19038,N_18884,N_18921);
or U19039 (N_19039,N_18873,N_18946);
xnor U19040 (N_19040,N_18996,N_18764);
or U19041 (N_19041,N_18905,N_18956);
xor U19042 (N_19042,N_18890,N_18859);
xor U19043 (N_19043,N_18876,N_18815);
nor U19044 (N_19044,N_18814,N_18963);
nor U19045 (N_19045,N_18752,N_18794);
xor U19046 (N_19046,N_18952,N_18795);
nor U19047 (N_19047,N_18939,N_18922);
xnor U19048 (N_19048,N_18862,N_18900);
or U19049 (N_19049,N_18804,N_18837);
xor U19050 (N_19050,N_18770,N_18839);
xor U19051 (N_19051,N_18771,N_18870);
xnor U19052 (N_19052,N_18964,N_18912);
xor U19053 (N_19053,N_18833,N_18844);
and U19054 (N_19054,N_18947,N_18979);
nor U19055 (N_19055,N_18788,N_18932);
or U19056 (N_19056,N_18829,N_18948);
nand U19057 (N_19057,N_18767,N_18792);
and U19058 (N_19058,N_18864,N_18750);
xor U19059 (N_19059,N_18889,N_18929);
nor U19060 (N_19060,N_18872,N_18897);
xor U19061 (N_19061,N_18954,N_18957);
nand U19062 (N_19062,N_18828,N_18852);
xnor U19063 (N_19063,N_18758,N_18776);
nor U19064 (N_19064,N_18959,N_18824);
xnor U19065 (N_19065,N_18850,N_18976);
and U19066 (N_19066,N_18931,N_18991);
xnor U19067 (N_19067,N_18875,N_18888);
or U19068 (N_19068,N_18968,N_18772);
or U19069 (N_19069,N_18925,N_18949);
nor U19070 (N_19070,N_18866,N_18777);
and U19071 (N_19071,N_18927,N_18755);
and U19072 (N_19072,N_18902,N_18942);
nand U19073 (N_19073,N_18832,N_18945);
xnor U19074 (N_19074,N_18901,N_18913);
or U19075 (N_19075,N_18786,N_18856);
nand U19076 (N_19076,N_18978,N_18819);
and U19077 (N_19077,N_18984,N_18846);
and U19078 (N_19078,N_18838,N_18982);
xnor U19079 (N_19079,N_18965,N_18941);
xnor U19080 (N_19080,N_18910,N_18854);
or U19081 (N_19081,N_18997,N_18918);
xnor U19082 (N_19082,N_18878,N_18924);
or U19083 (N_19083,N_18787,N_18841);
or U19084 (N_19084,N_18851,N_18802);
and U19085 (N_19085,N_18753,N_18930);
xor U19086 (N_19086,N_18950,N_18789);
or U19087 (N_19087,N_18955,N_18751);
nor U19088 (N_19088,N_18988,N_18810);
nand U19089 (N_19089,N_18882,N_18986);
or U19090 (N_19090,N_18843,N_18834);
or U19091 (N_19091,N_18831,N_18798);
xnor U19092 (N_19092,N_18826,N_18904);
nor U19093 (N_19093,N_18896,N_18754);
and U19094 (N_19094,N_18989,N_18857);
or U19095 (N_19095,N_18909,N_18967);
and U19096 (N_19096,N_18823,N_18935);
or U19097 (N_19097,N_18808,N_18993);
and U19098 (N_19098,N_18907,N_18811);
xor U19099 (N_19099,N_18916,N_18893);
or U19100 (N_19100,N_18801,N_18980);
nor U19101 (N_19101,N_18813,N_18780);
and U19102 (N_19102,N_18781,N_18953);
nor U19103 (N_19103,N_18881,N_18899);
nand U19104 (N_19104,N_18766,N_18867);
xor U19105 (N_19105,N_18999,N_18768);
nor U19106 (N_19106,N_18775,N_18886);
or U19107 (N_19107,N_18981,N_18782);
nor U19108 (N_19108,N_18868,N_18825);
or U19109 (N_19109,N_18971,N_18969);
and U19110 (N_19110,N_18759,N_18865);
xnor U19111 (N_19111,N_18869,N_18994);
or U19112 (N_19112,N_18796,N_18760);
nand U19113 (N_19113,N_18847,N_18830);
nor U19114 (N_19114,N_18926,N_18977);
and U19115 (N_19115,N_18756,N_18892);
nor U19116 (N_19116,N_18985,N_18861);
nor U19117 (N_19117,N_18817,N_18840);
nor U19118 (N_19118,N_18842,N_18827);
and U19119 (N_19119,N_18790,N_18970);
and U19120 (N_19120,N_18797,N_18972);
and U19121 (N_19121,N_18763,N_18998);
and U19122 (N_19122,N_18877,N_18975);
nor U19123 (N_19123,N_18785,N_18773);
nor U19124 (N_19124,N_18799,N_18936);
nand U19125 (N_19125,N_18946,N_18774);
xor U19126 (N_19126,N_18802,N_18940);
or U19127 (N_19127,N_18762,N_18859);
or U19128 (N_19128,N_18765,N_18997);
xor U19129 (N_19129,N_18930,N_18838);
or U19130 (N_19130,N_18858,N_18808);
xor U19131 (N_19131,N_18990,N_18773);
nand U19132 (N_19132,N_18805,N_18981);
or U19133 (N_19133,N_18750,N_18840);
nand U19134 (N_19134,N_18935,N_18776);
nor U19135 (N_19135,N_18864,N_18963);
or U19136 (N_19136,N_18962,N_18988);
and U19137 (N_19137,N_18888,N_18846);
or U19138 (N_19138,N_18816,N_18881);
or U19139 (N_19139,N_18785,N_18812);
nor U19140 (N_19140,N_18945,N_18771);
nand U19141 (N_19141,N_18927,N_18864);
xor U19142 (N_19142,N_18780,N_18991);
nor U19143 (N_19143,N_18785,N_18792);
nand U19144 (N_19144,N_18960,N_18959);
or U19145 (N_19145,N_18826,N_18976);
nor U19146 (N_19146,N_18962,N_18845);
and U19147 (N_19147,N_18801,N_18814);
nand U19148 (N_19148,N_18924,N_18933);
or U19149 (N_19149,N_18834,N_18858);
and U19150 (N_19150,N_18982,N_18827);
and U19151 (N_19151,N_18791,N_18984);
nand U19152 (N_19152,N_18921,N_18989);
nor U19153 (N_19153,N_18921,N_18837);
xor U19154 (N_19154,N_18926,N_18894);
nand U19155 (N_19155,N_18894,N_18887);
nand U19156 (N_19156,N_18869,N_18793);
or U19157 (N_19157,N_18948,N_18800);
xnor U19158 (N_19158,N_18846,N_18827);
xnor U19159 (N_19159,N_18828,N_18815);
nor U19160 (N_19160,N_18863,N_18955);
xnor U19161 (N_19161,N_18770,N_18942);
and U19162 (N_19162,N_18980,N_18845);
xor U19163 (N_19163,N_18890,N_18960);
xor U19164 (N_19164,N_18806,N_18939);
and U19165 (N_19165,N_18823,N_18958);
or U19166 (N_19166,N_18856,N_18805);
or U19167 (N_19167,N_18798,N_18811);
nand U19168 (N_19168,N_18997,N_18991);
nor U19169 (N_19169,N_18954,N_18808);
xor U19170 (N_19170,N_18910,N_18931);
nor U19171 (N_19171,N_18831,N_18806);
xor U19172 (N_19172,N_18957,N_18871);
xnor U19173 (N_19173,N_18846,N_18800);
and U19174 (N_19174,N_18907,N_18866);
or U19175 (N_19175,N_18998,N_18782);
nor U19176 (N_19176,N_18937,N_18775);
or U19177 (N_19177,N_18869,N_18795);
xnor U19178 (N_19178,N_18952,N_18770);
or U19179 (N_19179,N_18905,N_18978);
xor U19180 (N_19180,N_18924,N_18830);
nor U19181 (N_19181,N_18961,N_18848);
nor U19182 (N_19182,N_18980,N_18969);
and U19183 (N_19183,N_18801,N_18990);
xnor U19184 (N_19184,N_18797,N_18884);
xor U19185 (N_19185,N_18781,N_18955);
nand U19186 (N_19186,N_18817,N_18789);
and U19187 (N_19187,N_18863,N_18988);
xor U19188 (N_19188,N_18774,N_18844);
nand U19189 (N_19189,N_18972,N_18864);
or U19190 (N_19190,N_18858,N_18908);
and U19191 (N_19191,N_18912,N_18830);
nor U19192 (N_19192,N_18894,N_18822);
xor U19193 (N_19193,N_18852,N_18916);
and U19194 (N_19194,N_18835,N_18753);
nor U19195 (N_19195,N_18916,N_18903);
and U19196 (N_19196,N_18752,N_18937);
nand U19197 (N_19197,N_18898,N_18766);
nor U19198 (N_19198,N_18881,N_18860);
nand U19199 (N_19199,N_18800,N_18787);
nor U19200 (N_19200,N_18993,N_18821);
nand U19201 (N_19201,N_18978,N_18754);
xnor U19202 (N_19202,N_18898,N_18798);
nand U19203 (N_19203,N_18982,N_18905);
nor U19204 (N_19204,N_18805,N_18775);
nand U19205 (N_19205,N_18912,N_18829);
or U19206 (N_19206,N_18845,N_18869);
xnor U19207 (N_19207,N_18981,N_18814);
nand U19208 (N_19208,N_18783,N_18947);
nand U19209 (N_19209,N_18801,N_18813);
or U19210 (N_19210,N_18885,N_18881);
or U19211 (N_19211,N_18923,N_18843);
or U19212 (N_19212,N_18845,N_18828);
and U19213 (N_19213,N_18952,N_18951);
nand U19214 (N_19214,N_18922,N_18834);
xor U19215 (N_19215,N_18941,N_18796);
and U19216 (N_19216,N_18780,N_18926);
nor U19217 (N_19217,N_18916,N_18844);
and U19218 (N_19218,N_18898,N_18855);
xnor U19219 (N_19219,N_18818,N_18830);
nand U19220 (N_19220,N_18972,N_18780);
and U19221 (N_19221,N_18924,N_18835);
nand U19222 (N_19222,N_18963,N_18806);
and U19223 (N_19223,N_18810,N_18985);
nand U19224 (N_19224,N_18768,N_18851);
xor U19225 (N_19225,N_18882,N_18901);
and U19226 (N_19226,N_18867,N_18801);
nand U19227 (N_19227,N_18976,N_18874);
nand U19228 (N_19228,N_18911,N_18958);
or U19229 (N_19229,N_18979,N_18793);
and U19230 (N_19230,N_18833,N_18934);
or U19231 (N_19231,N_18895,N_18936);
and U19232 (N_19232,N_18938,N_18995);
xnor U19233 (N_19233,N_18786,N_18808);
or U19234 (N_19234,N_18827,N_18990);
or U19235 (N_19235,N_18928,N_18919);
and U19236 (N_19236,N_18994,N_18817);
nor U19237 (N_19237,N_18916,N_18788);
nor U19238 (N_19238,N_18957,N_18963);
nand U19239 (N_19239,N_18937,N_18959);
or U19240 (N_19240,N_18780,N_18979);
nor U19241 (N_19241,N_18838,N_18843);
nor U19242 (N_19242,N_18890,N_18954);
xnor U19243 (N_19243,N_18800,N_18954);
nor U19244 (N_19244,N_18828,N_18769);
xor U19245 (N_19245,N_18774,N_18986);
nand U19246 (N_19246,N_18878,N_18799);
and U19247 (N_19247,N_18911,N_18915);
or U19248 (N_19248,N_18796,N_18826);
xor U19249 (N_19249,N_18967,N_18840);
or U19250 (N_19250,N_19190,N_19141);
or U19251 (N_19251,N_19133,N_19070);
or U19252 (N_19252,N_19225,N_19105);
or U19253 (N_19253,N_19204,N_19093);
or U19254 (N_19254,N_19248,N_19118);
nor U19255 (N_19255,N_19087,N_19142);
and U19256 (N_19256,N_19085,N_19163);
nand U19257 (N_19257,N_19223,N_19067);
nand U19258 (N_19258,N_19246,N_19078);
and U19259 (N_19259,N_19162,N_19226);
and U19260 (N_19260,N_19171,N_19138);
and U19261 (N_19261,N_19159,N_19164);
nand U19262 (N_19262,N_19015,N_19187);
xnor U19263 (N_19263,N_19022,N_19121);
nand U19264 (N_19264,N_19028,N_19043);
nand U19265 (N_19265,N_19013,N_19144);
nand U19266 (N_19266,N_19244,N_19151);
xnor U19267 (N_19267,N_19177,N_19030);
nor U19268 (N_19268,N_19023,N_19103);
or U19269 (N_19269,N_19107,N_19056);
xnor U19270 (N_19270,N_19068,N_19046);
or U19271 (N_19271,N_19036,N_19011);
nor U19272 (N_19272,N_19047,N_19100);
and U19273 (N_19273,N_19062,N_19205);
or U19274 (N_19274,N_19066,N_19038);
xor U19275 (N_19275,N_19074,N_19051);
nor U19276 (N_19276,N_19154,N_19014);
nand U19277 (N_19277,N_19218,N_19053);
nand U19278 (N_19278,N_19097,N_19137);
and U19279 (N_19279,N_19122,N_19000);
nand U19280 (N_19280,N_19196,N_19052);
nand U19281 (N_19281,N_19130,N_19195);
xor U19282 (N_19282,N_19149,N_19099);
xor U19283 (N_19283,N_19131,N_19071);
or U19284 (N_19284,N_19126,N_19239);
and U19285 (N_19285,N_19245,N_19181);
nand U19286 (N_19286,N_19170,N_19045);
nand U19287 (N_19287,N_19109,N_19102);
or U19288 (N_19288,N_19150,N_19192);
nand U19289 (N_19289,N_19228,N_19167);
nand U19290 (N_19290,N_19220,N_19098);
nand U19291 (N_19291,N_19242,N_19124);
nand U19292 (N_19292,N_19227,N_19147);
nor U19293 (N_19293,N_19233,N_19208);
or U19294 (N_19294,N_19157,N_19082);
nor U19295 (N_19295,N_19235,N_19210);
nand U19296 (N_19296,N_19217,N_19044);
and U19297 (N_19297,N_19219,N_19004);
nand U19298 (N_19298,N_19128,N_19001);
nand U19299 (N_19299,N_19092,N_19182);
and U19300 (N_19300,N_19174,N_19139);
and U19301 (N_19301,N_19104,N_19148);
xor U19302 (N_19302,N_19160,N_19143);
nor U19303 (N_19303,N_19005,N_19112);
and U19304 (N_19304,N_19063,N_19010);
xor U19305 (N_19305,N_19029,N_19117);
and U19306 (N_19306,N_19050,N_19125);
nor U19307 (N_19307,N_19090,N_19179);
and U19308 (N_19308,N_19194,N_19165);
xnor U19309 (N_19309,N_19035,N_19249);
and U19310 (N_19310,N_19055,N_19199);
xor U19311 (N_19311,N_19060,N_19230);
and U19312 (N_19312,N_19009,N_19158);
nand U19313 (N_19313,N_19207,N_19229);
nand U19314 (N_19314,N_19119,N_19012);
and U19315 (N_19315,N_19113,N_19057);
nand U19316 (N_19316,N_19037,N_19108);
nor U19317 (N_19317,N_19198,N_19115);
nand U19318 (N_19318,N_19006,N_19088);
and U19319 (N_19319,N_19079,N_19173);
nor U19320 (N_19320,N_19027,N_19084);
and U19321 (N_19321,N_19191,N_19156);
nor U19322 (N_19322,N_19202,N_19212);
and U19323 (N_19323,N_19058,N_19188);
nand U19324 (N_19324,N_19189,N_19214);
and U19325 (N_19325,N_19241,N_19193);
nor U19326 (N_19326,N_19236,N_19059);
or U19327 (N_19327,N_19178,N_19176);
xnor U19328 (N_19328,N_19080,N_19211);
nor U19329 (N_19329,N_19221,N_19215);
nor U19330 (N_19330,N_19213,N_19240);
nor U19331 (N_19331,N_19224,N_19183);
or U19332 (N_19332,N_19021,N_19110);
nor U19333 (N_19333,N_19209,N_19120);
xor U19334 (N_19334,N_19168,N_19129);
xor U19335 (N_19335,N_19152,N_19185);
or U19336 (N_19336,N_19106,N_19134);
nand U19337 (N_19337,N_19132,N_19003);
nor U19338 (N_19338,N_19018,N_19065);
xor U19339 (N_19339,N_19032,N_19089);
nand U19340 (N_19340,N_19123,N_19206);
and U19341 (N_19341,N_19020,N_19081);
xor U19342 (N_19342,N_19146,N_19140);
nor U19343 (N_19343,N_19072,N_19232);
nor U19344 (N_19344,N_19247,N_19116);
nand U19345 (N_19345,N_19049,N_19002);
nor U19346 (N_19346,N_19016,N_19025);
nor U19347 (N_19347,N_19184,N_19073);
or U19348 (N_19348,N_19155,N_19197);
nor U19349 (N_19349,N_19026,N_19096);
or U19350 (N_19350,N_19031,N_19007);
nor U19351 (N_19351,N_19094,N_19175);
xnor U19352 (N_19352,N_19161,N_19064);
nand U19353 (N_19353,N_19201,N_19075);
nand U19354 (N_19354,N_19200,N_19077);
nand U19355 (N_19355,N_19101,N_19238);
xor U19356 (N_19356,N_19033,N_19019);
nor U19357 (N_19357,N_19039,N_19186);
nand U19358 (N_19358,N_19095,N_19091);
nor U19359 (N_19359,N_19243,N_19017);
or U19360 (N_19360,N_19203,N_19216);
nor U19361 (N_19361,N_19136,N_19024);
or U19362 (N_19362,N_19222,N_19041);
nor U19363 (N_19363,N_19034,N_19237);
xor U19364 (N_19364,N_19048,N_19054);
and U19365 (N_19365,N_19008,N_19086);
or U19366 (N_19366,N_19169,N_19069);
and U19367 (N_19367,N_19127,N_19172);
xor U19368 (N_19368,N_19114,N_19153);
or U19369 (N_19369,N_19040,N_19111);
xnor U19370 (N_19370,N_19083,N_19061);
nor U19371 (N_19371,N_19166,N_19234);
or U19372 (N_19372,N_19042,N_19145);
nor U19373 (N_19373,N_19135,N_19231);
nand U19374 (N_19374,N_19076,N_19180);
nor U19375 (N_19375,N_19113,N_19015);
or U19376 (N_19376,N_19025,N_19099);
nand U19377 (N_19377,N_19115,N_19001);
nor U19378 (N_19378,N_19182,N_19170);
or U19379 (N_19379,N_19102,N_19019);
and U19380 (N_19380,N_19075,N_19144);
nand U19381 (N_19381,N_19174,N_19123);
and U19382 (N_19382,N_19111,N_19199);
and U19383 (N_19383,N_19047,N_19179);
or U19384 (N_19384,N_19244,N_19098);
and U19385 (N_19385,N_19064,N_19034);
nor U19386 (N_19386,N_19045,N_19146);
xor U19387 (N_19387,N_19193,N_19064);
or U19388 (N_19388,N_19013,N_19054);
or U19389 (N_19389,N_19016,N_19237);
xnor U19390 (N_19390,N_19199,N_19180);
nand U19391 (N_19391,N_19210,N_19100);
nand U19392 (N_19392,N_19237,N_19214);
xor U19393 (N_19393,N_19117,N_19175);
or U19394 (N_19394,N_19234,N_19130);
or U19395 (N_19395,N_19220,N_19126);
or U19396 (N_19396,N_19145,N_19024);
nand U19397 (N_19397,N_19068,N_19111);
or U19398 (N_19398,N_19127,N_19072);
or U19399 (N_19399,N_19195,N_19004);
nand U19400 (N_19400,N_19180,N_19137);
or U19401 (N_19401,N_19006,N_19157);
xor U19402 (N_19402,N_19138,N_19056);
or U19403 (N_19403,N_19231,N_19024);
xnor U19404 (N_19404,N_19045,N_19111);
or U19405 (N_19405,N_19201,N_19051);
nand U19406 (N_19406,N_19101,N_19077);
nand U19407 (N_19407,N_19156,N_19220);
nor U19408 (N_19408,N_19079,N_19062);
and U19409 (N_19409,N_19131,N_19198);
or U19410 (N_19410,N_19186,N_19111);
nand U19411 (N_19411,N_19198,N_19190);
or U19412 (N_19412,N_19083,N_19200);
and U19413 (N_19413,N_19166,N_19124);
nor U19414 (N_19414,N_19165,N_19033);
nand U19415 (N_19415,N_19155,N_19161);
nand U19416 (N_19416,N_19184,N_19126);
nand U19417 (N_19417,N_19177,N_19127);
and U19418 (N_19418,N_19110,N_19011);
nor U19419 (N_19419,N_19211,N_19106);
nor U19420 (N_19420,N_19244,N_19048);
or U19421 (N_19421,N_19063,N_19024);
and U19422 (N_19422,N_19186,N_19055);
xor U19423 (N_19423,N_19167,N_19049);
nand U19424 (N_19424,N_19056,N_19050);
nor U19425 (N_19425,N_19009,N_19052);
xor U19426 (N_19426,N_19216,N_19237);
nor U19427 (N_19427,N_19083,N_19097);
nand U19428 (N_19428,N_19027,N_19141);
or U19429 (N_19429,N_19119,N_19068);
nand U19430 (N_19430,N_19184,N_19215);
or U19431 (N_19431,N_19062,N_19042);
xor U19432 (N_19432,N_19007,N_19045);
and U19433 (N_19433,N_19072,N_19119);
or U19434 (N_19434,N_19028,N_19012);
xor U19435 (N_19435,N_19031,N_19083);
and U19436 (N_19436,N_19059,N_19174);
xor U19437 (N_19437,N_19101,N_19179);
or U19438 (N_19438,N_19006,N_19219);
nand U19439 (N_19439,N_19129,N_19046);
nor U19440 (N_19440,N_19232,N_19033);
nor U19441 (N_19441,N_19217,N_19247);
nand U19442 (N_19442,N_19043,N_19098);
and U19443 (N_19443,N_19195,N_19168);
or U19444 (N_19444,N_19194,N_19216);
and U19445 (N_19445,N_19198,N_19239);
and U19446 (N_19446,N_19001,N_19050);
and U19447 (N_19447,N_19059,N_19223);
or U19448 (N_19448,N_19020,N_19091);
nand U19449 (N_19449,N_19022,N_19023);
and U19450 (N_19450,N_19110,N_19186);
nor U19451 (N_19451,N_19075,N_19182);
or U19452 (N_19452,N_19114,N_19166);
xnor U19453 (N_19453,N_19223,N_19142);
or U19454 (N_19454,N_19172,N_19106);
nand U19455 (N_19455,N_19204,N_19120);
and U19456 (N_19456,N_19140,N_19181);
xor U19457 (N_19457,N_19034,N_19246);
nor U19458 (N_19458,N_19015,N_19049);
or U19459 (N_19459,N_19081,N_19105);
or U19460 (N_19460,N_19022,N_19015);
nand U19461 (N_19461,N_19007,N_19219);
xor U19462 (N_19462,N_19186,N_19096);
and U19463 (N_19463,N_19208,N_19128);
and U19464 (N_19464,N_19173,N_19159);
xnor U19465 (N_19465,N_19097,N_19063);
or U19466 (N_19466,N_19002,N_19200);
xor U19467 (N_19467,N_19213,N_19120);
and U19468 (N_19468,N_19131,N_19006);
nor U19469 (N_19469,N_19219,N_19127);
xnor U19470 (N_19470,N_19175,N_19148);
or U19471 (N_19471,N_19049,N_19018);
or U19472 (N_19472,N_19221,N_19166);
and U19473 (N_19473,N_19162,N_19234);
nor U19474 (N_19474,N_19172,N_19149);
or U19475 (N_19475,N_19039,N_19202);
xnor U19476 (N_19476,N_19117,N_19220);
xnor U19477 (N_19477,N_19142,N_19064);
nand U19478 (N_19478,N_19043,N_19172);
or U19479 (N_19479,N_19021,N_19131);
and U19480 (N_19480,N_19160,N_19002);
xor U19481 (N_19481,N_19034,N_19174);
or U19482 (N_19482,N_19105,N_19203);
and U19483 (N_19483,N_19127,N_19134);
xor U19484 (N_19484,N_19025,N_19064);
xnor U19485 (N_19485,N_19090,N_19026);
or U19486 (N_19486,N_19134,N_19116);
and U19487 (N_19487,N_19049,N_19175);
nor U19488 (N_19488,N_19245,N_19113);
nor U19489 (N_19489,N_19143,N_19082);
or U19490 (N_19490,N_19208,N_19043);
and U19491 (N_19491,N_19030,N_19049);
nor U19492 (N_19492,N_19156,N_19166);
nor U19493 (N_19493,N_19009,N_19029);
or U19494 (N_19494,N_19148,N_19246);
or U19495 (N_19495,N_19105,N_19012);
and U19496 (N_19496,N_19042,N_19047);
nor U19497 (N_19497,N_19137,N_19204);
or U19498 (N_19498,N_19022,N_19024);
or U19499 (N_19499,N_19012,N_19120);
nand U19500 (N_19500,N_19263,N_19467);
nor U19501 (N_19501,N_19349,N_19482);
xnor U19502 (N_19502,N_19446,N_19287);
and U19503 (N_19503,N_19381,N_19396);
and U19504 (N_19504,N_19356,N_19327);
or U19505 (N_19505,N_19335,N_19478);
xor U19506 (N_19506,N_19322,N_19357);
nor U19507 (N_19507,N_19435,N_19484);
xnor U19508 (N_19508,N_19398,N_19388);
or U19509 (N_19509,N_19450,N_19382);
and U19510 (N_19510,N_19419,N_19378);
and U19511 (N_19511,N_19294,N_19472);
or U19512 (N_19512,N_19466,N_19493);
xnor U19513 (N_19513,N_19289,N_19348);
xor U19514 (N_19514,N_19267,N_19333);
xor U19515 (N_19515,N_19344,N_19371);
nand U19516 (N_19516,N_19369,N_19256);
nor U19517 (N_19517,N_19417,N_19496);
nor U19518 (N_19518,N_19433,N_19367);
xor U19519 (N_19519,N_19332,N_19401);
and U19520 (N_19520,N_19431,N_19281);
nor U19521 (N_19521,N_19340,N_19261);
nor U19522 (N_19522,N_19265,N_19479);
and U19523 (N_19523,N_19451,N_19293);
and U19524 (N_19524,N_19481,N_19443);
nand U19525 (N_19525,N_19483,N_19291);
xnor U19526 (N_19526,N_19485,N_19355);
or U19527 (N_19527,N_19390,N_19439);
nand U19528 (N_19528,N_19480,N_19361);
and U19529 (N_19529,N_19288,N_19468);
and U19530 (N_19530,N_19441,N_19442);
or U19531 (N_19531,N_19331,N_19424);
nor U19532 (N_19532,N_19299,N_19470);
nand U19533 (N_19533,N_19422,N_19298);
xnor U19534 (N_19534,N_19314,N_19409);
nor U19535 (N_19535,N_19319,N_19475);
nand U19536 (N_19536,N_19423,N_19427);
and U19537 (N_19537,N_19347,N_19455);
nand U19538 (N_19538,N_19339,N_19350);
or U19539 (N_19539,N_19326,N_19460);
nor U19540 (N_19540,N_19488,N_19497);
and U19541 (N_19541,N_19386,N_19402);
nor U19542 (N_19542,N_19385,N_19305);
xnor U19543 (N_19543,N_19477,N_19285);
nor U19544 (N_19544,N_19308,N_19368);
xnor U19545 (N_19545,N_19315,N_19370);
xor U19546 (N_19546,N_19316,N_19410);
and U19547 (N_19547,N_19270,N_19336);
and U19548 (N_19548,N_19328,N_19320);
nor U19549 (N_19549,N_19275,N_19408);
or U19550 (N_19550,N_19429,N_19301);
or U19551 (N_19551,N_19359,N_19421);
xnor U19552 (N_19552,N_19334,N_19325);
xor U19553 (N_19553,N_19387,N_19250);
and U19554 (N_19554,N_19338,N_19395);
nor U19555 (N_19555,N_19329,N_19413);
xor U19556 (N_19556,N_19474,N_19399);
xor U19557 (N_19557,N_19364,N_19376);
and U19558 (N_19558,N_19414,N_19458);
nand U19559 (N_19559,N_19411,N_19318);
or U19560 (N_19560,N_19469,N_19363);
and U19561 (N_19561,N_19342,N_19486);
nand U19562 (N_19562,N_19274,N_19461);
nor U19563 (N_19563,N_19307,N_19377);
nor U19564 (N_19564,N_19276,N_19384);
nand U19565 (N_19565,N_19252,N_19254);
and U19566 (N_19566,N_19449,N_19393);
nand U19567 (N_19567,N_19290,N_19268);
nand U19568 (N_19568,N_19375,N_19297);
and U19569 (N_19569,N_19292,N_19306);
nor U19570 (N_19570,N_19277,N_19330);
nor U19571 (N_19571,N_19358,N_19445);
nor U19572 (N_19572,N_19444,N_19426);
nor U19573 (N_19573,N_19494,N_19491);
xor U19574 (N_19574,N_19490,N_19323);
nor U19575 (N_19575,N_19471,N_19313);
nor U19576 (N_19576,N_19264,N_19400);
nand U19577 (N_19577,N_19416,N_19403);
nand U19578 (N_19578,N_19459,N_19260);
nand U19579 (N_19579,N_19372,N_19452);
nand U19580 (N_19580,N_19391,N_19269);
nand U19581 (N_19581,N_19346,N_19352);
nor U19582 (N_19582,N_19262,N_19279);
or U19583 (N_19583,N_19311,N_19440);
or U19584 (N_19584,N_19282,N_19425);
and U19585 (N_19585,N_19300,N_19257);
nand U19586 (N_19586,N_19258,N_19354);
xor U19587 (N_19587,N_19351,N_19343);
xnor U19588 (N_19588,N_19374,N_19283);
and U19589 (N_19589,N_19495,N_19310);
nand U19590 (N_19590,N_19407,N_19380);
or U19591 (N_19591,N_19432,N_19420);
or U19592 (N_19592,N_19394,N_19366);
xor U19593 (N_19593,N_19284,N_19457);
or U19594 (N_19594,N_19296,N_19447);
and U19595 (N_19595,N_19389,N_19360);
or U19596 (N_19596,N_19453,N_19255);
or U19597 (N_19597,N_19272,N_19345);
and U19598 (N_19598,N_19304,N_19365);
and U19599 (N_19599,N_19302,N_19397);
and U19600 (N_19600,N_19324,N_19251);
and U19601 (N_19601,N_19259,N_19448);
nand U19602 (N_19602,N_19341,N_19271);
or U19603 (N_19603,N_19489,N_19379);
xor U19604 (N_19604,N_19499,N_19383);
xnor U19605 (N_19605,N_19465,N_19434);
xor U19606 (N_19606,N_19418,N_19286);
or U19607 (N_19607,N_19405,N_19373);
nand U19608 (N_19608,N_19303,N_19309);
nor U19609 (N_19609,N_19278,N_19454);
nor U19610 (N_19610,N_19464,N_19437);
nand U19611 (N_19611,N_19412,N_19463);
or U19612 (N_19612,N_19273,N_19321);
xor U19613 (N_19613,N_19312,N_19337);
nor U19614 (N_19614,N_19280,N_19430);
and U19615 (N_19615,N_19415,N_19456);
and U19616 (N_19616,N_19487,N_19406);
and U19617 (N_19617,N_19492,N_19462);
nand U19618 (N_19618,N_19353,N_19295);
xor U19619 (N_19619,N_19392,N_19317);
nor U19620 (N_19620,N_19476,N_19428);
and U19621 (N_19621,N_19266,N_19473);
and U19622 (N_19622,N_19404,N_19498);
xor U19623 (N_19623,N_19362,N_19436);
or U19624 (N_19624,N_19438,N_19253);
nor U19625 (N_19625,N_19478,N_19472);
or U19626 (N_19626,N_19383,N_19453);
and U19627 (N_19627,N_19362,N_19391);
xnor U19628 (N_19628,N_19332,N_19498);
or U19629 (N_19629,N_19495,N_19411);
xor U19630 (N_19630,N_19435,N_19421);
and U19631 (N_19631,N_19460,N_19485);
xnor U19632 (N_19632,N_19458,N_19257);
nand U19633 (N_19633,N_19451,N_19442);
or U19634 (N_19634,N_19411,N_19352);
nand U19635 (N_19635,N_19258,N_19387);
nor U19636 (N_19636,N_19286,N_19272);
nand U19637 (N_19637,N_19446,N_19473);
nand U19638 (N_19638,N_19271,N_19309);
nor U19639 (N_19639,N_19288,N_19367);
and U19640 (N_19640,N_19304,N_19289);
xnor U19641 (N_19641,N_19456,N_19309);
nand U19642 (N_19642,N_19389,N_19258);
and U19643 (N_19643,N_19262,N_19386);
xor U19644 (N_19644,N_19292,N_19361);
nor U19645 (N_19645,N_19461,N_19419);
nor U19646 (N_19646,N_19336,N_19389);
nor U19647 (N_19647,N_19467,N_19266);
or U19648 (N_19648,N_19365,N_19432);
nor U19649 (N_19649,N_19459,N_19483);
or U19650 (N_19650,N_19317,N_19490);
nand U19651 (N_19651,N_19329,N_19454);
xnor U19652 (N_19652,N_19471,N_19344);
or U19653 (N_19653,N_19352,N_19479);
xnor U19654 (N_19654,N_19310,N_19319);
nand U19655 (N_19655,N_19363,N_19293);
and U19656 (N_19656,N_19418,N_19343);
or U19657 (N_19657,N_19256,N_19321);
or U19658 (N_19658,N_19387,N_19333);
or U19659 (N_19659,N_19444,N_19488);
nand U19660 (N_19660,N_19356,N_19386);
or U19661 (N_19661,N_19473,N_19342);
and U19662 (N_19662,N_19394,N_19437);
xnor U19663 (N_19663,N_19253,N_19284);
nor U19664 (N_19664,N_19363,N_19305);
nand U19665 (N_19665,N_19258,N_19477);
or U19666 (N_19666,N_19300,N_19264);
or U19667 (N_19667,N_19454,N_19390);
xnor U19668 (N_19668,N_19408,N_19424);
and U19669 (N_19669,N_19460,N_19392);
xnor U19670 (N_19670,N_19302,N_19487);
nand U19671 (N_19671,N_19295,N_19345);
nand U19672 (N_19672,N_19456,N_19342);
nor U19673 (N_19673,N_19469,N_19298);
nor U19674 (N_19674,N_19418,N_19291);
xnor U19675 (N_19675,N_19401,N_19367);
nand U19676 (N_19676,N_19325,N_19375);
nor U19677 (N_19677,N_19296,N_19260);
nor U19678 (N_19678,N_19460,N_19466);
and U19679 (N_19679,N_19482,N_19252);
nand U19680 (N_19680,N_19448,N_19407);
nand U19681 (N_19681,N_19469,N_19262);
and U19682 (N_19682,N_19287,N_19335);
nand U19683 (N_19683,N_19377,N_19411);
xnor U19684 (N_19684,N_19411,N_19425);
nand U19685 (N_19685,N_19465,N_19328);
nand U19686 (N_19686,N_19333,N_19493);
or U19687 (N_19687,N_19364,N_19353);
xor U19688 (N_19688,N_19451,N_19279);
nor U19689 (N_19689,N_19353,N_19469);
nor U19690 (N_19690,N_19360,N_19399);
nand U19691 (N_19691,N_19367,N_19389);
nor U19692 (N_19692,N_19441,N_19380);
and U19693 (N_19693,N_19399,N_19331);
or U19694 (N_19694,N_19478,N_19307);
and U19695 (N_19695,N_19290,N_19447);
nand U19696 (N_19696,N_19401,N_19312);
or U19697 (N_19697,N_19260,N_19325);
nand U19698 (N_19698,N_19436,N_19355);
nand U19699 (N_19699,N_19320,N_19414);
nand U19700 (N_19700,N_19435,N_19345);
and U19701 (N_19701,N_19483,N_19252);
xor U19702 (N_19702,N_19420,N_19448);
and U19703 (N_19703,N_19285,N_19403);
or U19704 (N_19704,N_19499,N_19334);
and U19705 (N_19705,N_19379,N_19343);
nor U19706 (N_19706,N_19499,N_19472);
and U19707 (N_19707,N_19275,N_19291);
nand U19708 (N_19708,N_19399,N_19347);
xor U19709 (N_19709,N_19443,N_19421);
or U19710 (N_19710,N_19454,N_19377);
nor U19711 (N_19711,N_19450,N_19283);
xnor U19712 (N_19712,N_19462,N_19309);
xnor U19713 (N_19713,N_19289,N_19269);
or U19714 (N_19714,N_19410,N_19404);
or U19715 (N_19715,N_19354,N_19347);
and U19716 (N_19716,N_19421,N_19330);
and U19717 (N_19717,N_19336,N_19319);
nand U19718 (N_19718,N_19369,N_19349);
xnor U19719 (N_19719,N_19366,N_19411);
or U19720 (N_19720,N_19440,N_19421);
nand U19721 (N_19721,N_19381,N_19412);
and U19722 (N_19722,N_19366,N_19401);
nand U19723 (N_19723,N_19365,N_19427);
nor U19724 (N_19724,N_19289,N_19294);
xnor U19725 (N_19725,N_19294,N_19343);
or U19726 (N_19726,N_19367,N_19440);
or U19727 (N_19727,N_19329,N_19263);
nand U19728 (N_19728,N_19300,N_19450);
xor U19729 (N_19729,N_19405,N_19283);
nand U19730 (N_19730,N_19294,N_19298);
nand U19731 (N_19731,N_19415,N_19390);
xor U19732 (N_19732,N_19421,N_19476);
and U19733 (N_19733,N_19429,N_19449);
nand U19734 (N_19734,N_19474,N_19343);
xor U19735 (N_19735,N_19256,N_19322);
or U19736 (N_19736,N_19416,N_19394);
or U19737 (N_19737,N_19448,N_19267);
nor U19738 (N_19738,N_19420,N_19435);
and U19739 (N_19739,N_19451,N_19277);
or U19740 (N_19740,N_19448,N_19421);
xor U19741 (N_19741,N_19303,N_19409);
xor U19742 (N_19742,N_19489,N_19271);
xor U19743 (N_19743,N_19312,N_19258);
nor U19744 (N_19744,N_19323,N_19364);
xnor U19745 (N_19745,N_19339,N_19428);
and U19746 (N_19746,N_19405,N_19301);
nand U19747 (N_19747,N_19465,N_19390);
xor U19748 (N_19748,N_19494,N_19362);
nand U19749 (N_19749,N_19285,N_19265);
nand U19750 (N_19750,N_19714,N_19514);
xnor U19751 (N_19751,N_19698,N_19717);
nand U19752 (N_19752,N_19562,N_19630);
and U19753 (N_19753,N_19688,N_19639);
nand U19754 (N_19754,N_19604,N_19621);
and U19755 (N_19755,N_19590,N_19538);
xnor U19756 (N_19756,N_19536,N_19738);
and U19757 (N_19757,N_19610,N_19742);
xnor U19758 (N_19758,N_19715,N_19641);
nor U19759 (N_19759,N_19697,N_19693);
xnor U19760 (N_19760,N_19667,N_19707);
or U19761 (N_19761,N_19512,N_19623);
and U19762 (N_19762,N_19637,N_19664);
and U19763 (N_19763,N_19551,N_19612);
and U19764 (N_19764,N_19710,N_19704);
or U19765 (N_19765,N_19665,N_19656);
nor U19766 (N_19766,N_19689,N_19614);
nor U19767 (N_19767,N_19577,N_19617);
or U19768 (N_19768,N_19719,N_19530);
xnor U19769 (N_19769,N_19691,N_19725);
xnor U19770 (N_19770,N_19507,N_19699);
nor U19771 (N_19771,N_19560,N_19556);
xor U19772 (N_19772,N_19574,N_19650);
or U19773 (N_19773,N_19713,N_19554);
nand U19774 (N_19774,N_19526,N_19678);
and U19775 (N_19775,N_19631,N_19548);
and U19776 (N_19776,N_19607,N_19733);
and U19777 (N_19777,N_19745,N_19661);
or U19778 (N_19778,N_19675,N_19681);
nand U19779 (N_19779,N_19606,N_19726);
nand U19780 (N_19780,N_19647,N_19564);
nand U19781 (N_19781,N_19504,N_19660);
nor U19782 (N_19782,N_19748,N_19625);
and U19783 (N_19783,N_19674,N_19599);
xor U19784 (N_19784,N_19692,N_19558);
and U19785 (N_19785,N_19586,N_19722);
nor U19786 (N_19786,N_19735,N_19569);
nor U19787 (N_19787,N_19627,N_19505);
or U19788 (N_19788,N_19711,N_19701);
nand U19789 (N_19789,N_19723,N_19629);
nor U19790 (N_19790,N_19695,N_19508);
nor U19791 (N_19791,N_19712,N_19736);
nor U19792 (N_19792,N_19626,N_19608);
and U19793 (N_19793,N_19567,N_19533);
nor U19794 (N_19794,N_19522,N_19655);
xnor U19795 (N_19795,N_19615,N_19502);
nand U19796 (N_19796,N_19549,N_19624);
nor U19797 (N_19797,N_19720,N_19669);
and U19798 (N_19798,N_19525,N_19676);
nand U19799 (N_19799,N_19588,N_19593);
nand U19800 (N_19800,N_19500,N_19597);
and U19801 (N_19801,N_19649,N_19657);
nor U19802 (N_19802,N_19634,N_19563);
xnor U19803 (N_19803,N_19747,N_19523);
and U19804 (N_19804,N_19559,N_19513);
nand U19805 (N_19805,N_19611,N_19565);
xor U19806 (N_19806,N_19645,N_19552);
xor U19807 (N_19807,N_19557,N_19550);
and U19808 (N_19808,N_19658,N_19578);
or U19809 (N_19809,N_19737,N_19679);
nand U19810 (N_19810,N_19618,N_19584);
nand U19811 (N_19811,N_19594,N_19501);
nand U19812 (N_19812,N_19546,N_19687);
xor U19813 (N_19813,N_19587,N_19542);
and U19814 (N_19814,N_19603,N_19729);
or U19815 (N_19815,N_19696,N_19740);
or U19816 (N_19816,N_19709,N_19668);
and U19817 (N_19817,N_19648,N_19613);
and U19818 (N_19818,N_19638,N_19528);
or U19819 (N_19819,N_19732,N_19534);
nand U19820 (N_19820,N_19568,N_19702);
and U19821 (N_19821,N_19553,N_19561);
nand U19822 (N_19822,N_19666,N_19671);
nand U19823 (N_19823,N_19616,N_19589);
xnor U19824 (N_19824,N_19677,N_19690);
xor U19825 (N_19825,N_19598,N_19601);
xnor U19826 (N_19826,N_19581,N_19700);
and U19827 (N_19827,N_19663,N_19596);
nor U19828 (N_19828,N_19566,N_19516);
or U19829 (N_19829,N_19591,N_19555);
nand U19830 (N_19830,N_19686,N_19672);
nand U19831 (N_19831,N_19673,N_19519);
nand U19832 (N_19832,N_19600,N_19537);
xnor U19833 (N_19833,N_19576,N_19592);
or U19834 (N_19834,N_19570,N_19595);
nand U19835 (N_19835,N_19620,N_19541);
xnor U19836 (N_19836,N_19743,N_19705);
nor U19837 (N_19837,N_19544,N_19716);
and U19838 (N_19838,N_19746,N_19585);
nand U19839 (N_19839,N_19506,N_19741);
nand U19840 (N_19840,N_19540,N_19529);
and U19841 (N_19841,N_19524,N_19543);
and U19842 (N_19842,N_19662,N_19531);
nor U19843 (N_19843,N_19582,N_19646);
or U19844 (N_19844,N_19535,N_19683);
or U19845 (N_19845,N_19632,N_19628);
nand U19846 (N_19846,N_19680,N_19708);
or U19847 (N_19847,N_19527,N_19642);
xor U19848 (N_19848,N_19602,N_19659);
and U19849 (N_19849,N_19744,N_19734);
nor U19850 (N_19850,N_19517,N_19739);
or U19851 (N_19851,N_19730,N_19653);
nor U19852 (N_19852,N_19518,N_19703);
and U19853 (N_19853,N_19575,N_19572);
and U19854 (N_19854,N_19503,N_19635);
xnor U19855 (N_19855,N_19651,N_19640);
nand U19856 (N_19856,N_19605,N_19643);
nand U19857 (N_19857,N_19511,N_19521);
and U19858 (N_19858,N_19579,N_19670);
and U19859 (N_19859,N_19724,N_19636);
nor U19860 (N_19860,N_19622,N_19510);
nor U19861 (N_19861,N_19654,N_19706);
nor U19862 (N_19862,N_19539,N_19644);
nor U19863 (N_19863,N_19571,N_19619);
xor U19864 (N_19864,N_19573,N_19652);
and U19865 (N_19865,N_19633,N_19532);
xnor U19866 (N_19866,N_19684,N_19728);
nand U19867 (N_19867,N_19685,N_19694);
xor U19868 (N_19868,N_19545,N_19580);
or U19869 (N_19869,N_19682,N_19583);
or U19870 (N_19870,N_19727,N_19731);
xnor U19871 (N_19871,N_19609,N_19547);
nand U19872 (N_19872,N_19718,N_19721);
xor U19873 (N_19873,N_19509,N_19515);
or U19874 (N_19874,N_19749,N_19520);
and U19875 (N_19875,N_19692,N_19540);
nand U19876 (N_19876,N_19590,N_19737);
xnor U19877 (N_19877,N_19504,N_19617);
nor U19878 (N_19878,N_19549,N_19589);
and U19879 (N_19879,N_19565,N_19641);
and U19880 (N_19880,N_19508,N_19639);
xor U19881 (N_19881,N_19530,N_19666);
xor U19882 (N_19882,N_19577,N_19673);
xor U19883 (N_19883,N_19549,N_19508);
and U19884 (N_19884,N_19634,N_19518);
and U19885 (N_19885,N_19719,N_19698);
nor U19886 (N_19886,N_19727,N_19708);
and U19887 (N_19887,N_19630,N_19555);
nand U19888 (N_19888,N_19583,N_19553);
nor U19889 (N_19889,N_19665,N_19601);
and U19890 (N_19890,N_19646,N_19634);
xnor U19891 (N_19891,N_19740,N_19569);
or U19892 (N_19892,N_19626,N_19576);
and U19893 (N_19893,N_19697,N_19731);
nor U19894 (N_19894,N_19580,N_19644);
nand U19895 (N_19895,N_19668,N_19640);
xor U19896 (N_19896,N_19633,N_19552);
or U19897 (N_19897,N_19648,N_19654);
or U19898 (N_19898,N_19666,N_19573);
and U19899 (N_19899,N_19663,N_19699);
nor U19900 (N_19900,N_19505,N_19714);
or U19901 (N_19901,N_19539,N_19529);
or U19902 (N_19902,N_19540,N_19737);
and U19903 (N_19903,N_19510,N_19516);
or U19904 (N_19904,N_19717,N_19578);
xor U19905 (N_19905,N_19647,N_19524);
or U19906 (N_19906,N_19655,N_19579);
nor U19907 (N_19907,N_19685,N_19553);
and U19908 (N_19908,N_19559,N_19651);
nand U19909 (N_19909,N_19543,N_19643);
and U19910 (N_19910,N_19623,N_19712);
nor U19911 (N_19911,N_19576,N_19612);
or U19912 (N_19912,N_19670,N_19655);
nand U19913 (N_19913,N_19703,N_19670);
or U19914 (N_19914,N_19718,N_19523);
or U19915 (N_19915,N_19710,N_19621);
and U19916 (N_19916,N_19524,N_19696);
or U19917 (N_19917,N_19646,N_19527);
or U19918 (N_19918,N_19512,N_19646);
and U19919 (N_19919,N_19545,N_19532);
nor U19920 (N_19920,N_19718,N_19547);
or U19921 (N_19921,N_19563,N_19544);
nand U19922 (N_19922,N_19748,N_19687);
and U19923 (N_19923,N_19510,N_19709);
xor U19924 (N_19924,N_19625,N_19564);
nand U19925 (N_19925,N_19699,N_19682);
or U19926 (N_19926,N_19712,N_19544);
nand U19927 (N_19927,N_19745,N_19593);
nor U19928 (N_19928,N_19627,N_19534);
or U19929 (N_19929,N_19623,N_19709);
xor U19930 (N_19930,N_19514,N_19704);
xnor U19931 (N_19931,N_19505,N_19709);
xor U19932 (N_19932,N_19667,N_19746);
or U19933 (N_19933,N_19714,N_19694);
and U19934 (N_19934,N_19526,N_19570);
nand U19935 (N_19935,N_19698,N_19707);
or U19936 (N_19936,N_19537,N_19683);
nor U19937 (N_19937,N_19580,N_19615);
xor U19938 (N_19938,N_19542,N_19724);
nand U19939 (N_19939,N_19684,N_19673);
nor U19940 (N_19940,N_19620,N_19595);
nand U19941 (N_19941,N_19643,N_19732);
or U19942 (N_19942,N_19656,N_19730);
nand U19943 (N_19943,N_19733,N_19513);
and U19944 (N_19944,N_19596,N_19617);
and U19945 (N_19945,N_19556,N_19668);
nand U19946 (N_19946,N_19541,N_19601);
nand U19947 (N_19947,N_19710,N_19676);
xnor U19948 (N_19948,N_19719,N_19689);
xor U19949 (N_19949,N_19627,N_19609);
and U19950 (N_19950,N_19640,N_19539);
nor U19951 (N_19951,N_19710,N_19615);
nor U19952 (N_19952,N_19603,N_19732);
xor U19953 (N_19953,N_19744,N_19680);
and U19954 (N_19954,N_19572,N_19536);
nor U19955 (N_19955,N_19506,N_19701);
nor U19956 (N_19956,N_19601,N_19594);
or U19957 (N_19957,N_19531,N_19550);
or U19958 (N_19958,N_19643,N_19603);
nand U19959 (N_19959,N_19653,N_19613);
nor U19960 (N_19960,N_19743,N_19734);
nand U19961 (N_19961,N_19590,N_19690);
nand U19962 (N_19962,N_19599,N_19574);
xnor U19963 (N_19963,N_19527,N_19613);
xnor U19964 (N_19964,N_19695,N_19732);
or U19965 (N_19965,N_19743,N_19586);
nor U19966 (N_19966,N_19579,N_19562);
xor U19967 (N_19967,N_19591,N_19706);
nand U19968 (N_19968,N_19602,N_19501);
xor U19969 (N_19969,N_19525,N_19608);
nand U19970 (N_19970,N_19671,N_19640);
or U19971 (N_19971,N_19687,N_19592);
xor U19972 (N_19972,N_19577,N_19644);
or U19973 (N_19973,N_19671,N_19545);
nor U19974 (N_19974,N_19542,N_19546);
nor U19975 (N_19975,N_19746,N_19745);
and U19976 (N_19976,N_19653,N_19660);
and U19977 (N_19977,N_19638,N_19518);
nor U19978 (N_19978,N_19584,N_19688);
and U19979 (N_19979,N_19564,N_19598);
nor U19980 (N_19980,N_19727,N_19628);
nand U19981 (N_19981,N_19607,N_19646);
xor U19982 (N_19982,N_19746,N_19547);
nand U19983 (N_19983,N_19598,N_19637);
or U19984 (N_19984,N_19669,N_19536);
or U19985 (N_19985,N_19533,N_19511);
or U19986 (N_19986,N_19551,N_19689);
or U19987 (N_19987,N_19513,N_19540);
xor U19988 (N_19988,N_19605,N_19675);
or U19989 (N_19989,N_19502,N_19662);
nand U19990 (N_19990,N_19608,N_19619);
nand U19991 (N_19991,N_19615,N_19690);
and U19992 (N_19992,N_19744,N_19704);
and U19993 (N_19993,N_19555,N_19525);
xnor U19994 (N_19994,N_19706,N_19542);
nor U19995 (N_19995,N_19697,N_19727);
xor U19996 (N_19996,N_19614,N_19546);
xnor U19997 (N_19997,N_19633,N_19558);
or U19998 (N_19998,N_19700,N_19518);
nand U19999 (N_19999,N_19665,N_19644);
or U20000 (N_20000,N_19856,N_19827);
nor U20001 (N_20001,N_19810,N_19845);
nand U20002 (N_20002,N_19945,N_19991);
xnor U20003 (N_20003,N_19999,N_19787);
and U20004 (N_20004,N_19910,N_19886);
nor U20005 (N_20005,N_19826,N_19985);
xor U20006 (N_20006,N_19891,N_19915);
xor U20007 (N_20007,N_19987,N_19939);
nand U20008 (N_20008,N_19896,N_19873);
and U20009 (N_20009,N_19997,N_19981);
nor U20010 (N_20010,N_19913,N_19956);
xnor U20011 (N_20011,N_19778,N_19828);
nor U20012 (N_20012,N_19862,N_19859);
and U20013 (N_20013,N_19898,N_19989);
nor U20014 (N_20014,N_19951,N_19766);
and U20015 (N_20015,N_19751,N_19941);
xnor U20016 (N_20016,N_19835,N_19995);
nor U20017 (N_20017,N_19978,N_19962);
and U20018 (N_20018,N_19935,N_19803);
and U20019 (N_20019,N_19922,N_19868);
or U20020 (N_20020,N_19963,N_19954);
or U20021 (N_20021,N_19850,N_19974);
xor U20022 (N_20022,N_19966,N_19755);
and U20023 (N_20023,N_19964,N_19914);
or U20024 (N_20024,N_19878,N_19967);
nor U20025 (N_20025,N_19846,N_19952);
nand U20026 (N_20026,N_19816,N_19905);
nand U20027 (N_20027,N_19793,N_19775);
xnor U20028 (N_20028,N_19938,N_19806);
nand U20029 (N_20029,N_19866,N_19921);
xnor U20030 (N_20030,N_19830,N_19979);
nor U20031 (N_20031,N_19882,N_19943);
nand U20032 (N_20032,N_19777,N_19942);
nand U20033 (N_20033,N_19757,N_19770);
nand U20034 (N_20034,N_19871,N_19976);
nand U20035 (N_20035,N_19900,N_19799);
xnor U20036 (N_20036,N_19853,N_19811);
xor U20037 (N_20037,N_19959,N_19791);
xor U20038 (N_20038,N_19877,N_19761);
nand U20039 (N_20039,N_19968,N_19788);
nand U20040 (N_20040,N_19818,N_19771);
xnor U20041 (N_20041,N_19798,N_19795);
nor U20042 (N_20042,N_19919,N_19925);
xnor U20043 (N_20043,N_19909,N_19836);
or U20044 (N_20044,N_19769,N_19960);
nor U20045 (N_20045,N_19837,N_19800);
xnor U20046 (N_20046,N_19948,N_19955);
and U20047 (N_20047,N_19903,N_19809);
and U20048 (N_20048,N_19988,N_19773);
and U20049 (N_20049,N_19867,N_19932);
nor U20050 (N_20050,N_19977,N_19872);
nand U20051 (N_20051,N_19764,N_19881);
xor U20052 (N_20052,N_19883,N_19944);
xnor U20053 (N_20053,N_19840,N_19958);
and U20054 (N_20054,N_19933,N_19753);
and U20055 (N_20055,N_19897,N_19879);
or U20056 (N_20056,N_19975,N_19953);
or U20057 (N_20057,N_19807,N_19970);
or U20058 (N_20058,N_19920,N_19779);
and U20059 (N_20059,N_19923,N_19829);
xor U20060 (N_20060,N_19885,N_19961);
xor U20061 (N_20061,N_19785,N_19834);
nor U20062 (N_20062,N_19860,N_19847);
nand U20063 (N_20063,N_19855,N_19801);
xor U20064 (N_20064,N_19814,N_19813);
xor U20065 (N_20065,N_19880,N_19822);
nor U20066 (N_20066,N_19869,N_19858);
and U20067 (N_20067,N_19950,N_19783);
nand U20068 (N_20068,N_19864,N_19812);
nand U20069 (N_20069,N_19917,N_19780);
nand U20070 (N_20070,N_19865,N_19884);
and U20071 (N_20071,N_19888,N_19969);
xnor U20072 (N_20072,N_19931,N_19762);
nor U20073 (N_20073,N_19870,N_19758);
nand U20074 (N_20074,N_19823,N_19894);
xnor U20075 (N_20075,N_19875,N_19852);
xnor U20076 (N_20076,N_19851,N_19998);
nor U20077 (N_20077,N_19750,N_19763);
nor U20078 (N_20078,N_19902,N_19817);
or U20079 (N_20079,N_19876,N_19973);
nor U20080 (N_20080,N_19936,N_19874);
xor U20081 (N_20081,N_19887,N_19984);
nand U20082 (N_20082,N_19831,N_19992);
nor U20083 (N_20083,N_19849,N_19857);
nand U20084 (N_20084,N_19792,N_19971);
nand U20085 (N_20085,N_19794,N_19899);
or U20086 (N_20086,N_19754,N_19756);
or U20087 (N_20087,N_19996,N_19893);
and U20088 (N_20088,N_19927,N_19796);
nor U20089 (N_20089,N_19924,N_19765);
nand U20090 (N_20090,N_19843,N_19947);
and U20091 (N_20091,N_19832,N_19782);
or U20092 (N_20092,N_19772,N_19928);
nor U20093 (N_20093,N_19918,N_19912);
xor U20094 (N_20094,N_19982,N_19789);
and U20095 (N_20095,N_19752,N_19957);
nand U20096 (N_20096,N_19930,N_19842);
xor U20097 (N_20097,N_19781,N_19838);
nor U20098 (N_20098,N_19890,N_19805);
nor U20099 (N_20099,N_19784,N_19926);
or U20100 (N_20100,N_19895,N_19802);
and U20101 (N_20101,N_19937,N_19916);
nand U20102 (N_20102,N_19949,N_19861);
and U20103 (N_20103,N_19892,N_19993);
xnor U20104 (N_20104,N_19904,N_19833);
and U20105 (N_20105,N_19863,N_19854);
nor U20106 (N_20106,N_19819,N_19776);
nor U20107 (N_20107,N_19990,N_19821);
xnor U20108 (N_20108,N_19824,N_19848);
nand U20109 (N_20109,N_19972,N_19759);
nor U20110 (N_20110,N_19825,N_19929);
and U20111 (N_20111,N_19760,N_19911);
and U20112 (N_20112,N_19797,N_19786);
or U20113 (N_20113,N_19906,N_19889);
xor U20114 (N_20114,N_19841,N_19965);
nor U20115 (N_20115,N_19808,N_19980);
or U20116 (N_20116,N_19983,N_19839);
and U20117 (N_20117,N_19844,N_19986);
or U20118 (N_20118,N_19946,N_19768);
xnor U20119 (N_20119,N_19767,N_19940);
or U20120 (N_20120,N_19994,N_19804);
nand U20121 (N_20121,N_19901,N_19815);
and U20122 (N_20122,N_19774,N_19820);
nand U20123 (N_20123,N_19790,N_19934);
and U20124 (N_20124,N_19907,N_19908);
and U20125 (N_20125,N_19799,N_19890);
or U20126 (N_20126,N_19826,N_19760);
and U20127 (N_20127,N_19932,N_19925);
and U20128 (N_20128,N_19982,N_19792);
xor U20129 (N_20129,N_19973,N_19818);
or U20130 (N_20130,N_19984,N_19756);
nor U20131 (N_20131,N_19904,N_19785);
nand U20132 (N_20132,N_19957,N_19905);
nor U20133 (N_20133,N_19990,N_19953);
nor U20134 (N_20134,N_19915,N_19975);
xor U20135 (N_20135,N_19910,N_19856);
xor U20136 (N_20136,N_19778,N_19974);
nor U20137 (N_20137,N_19753,N_19840);
nand U20138 (N_20138,N_19859,N_19891);
nand U20139 (N_20139,N_19957,N_19917);
xnor U20140 (N_20140,N_19978,N_19954);
and U20141 (N_20141,N_19821,N_19904);
and U20142 (N_20142,N_19753,N_19901);
nand U20143 (N_20143,N_19887,N_19982);
nand U20144 (N_20144,N_19950,N_19921);
or U20145 (N_20145,N_19874,N_19912);
nand U20146 (N_20146,N_19780,N_19757);
xnor U20147 (N_20147,N_19763,N_19751);
xor U20148 (N_20148,N_19865,N_19863);
nor U20149 (N_20149,N_19957,N_19954);
or U20150 (N_20150,N_19912,N_19792);
nand U20151 (N_20151,N_19994,N_19962);
nand U20152 (N_20152,N_19764,N_19902);
xor U20153 (N_20153,N_19926,N_19783);
or U20154 (N_20154,N_19823,N_19956);
nor U20155 (N_20155,N_19880,N_19866);
xor U20156 (N_20156,N_19815,N_19802);
or U20157 (N_20157,N_19980,N_19767);
nor U20158 (N_20158,N_19949,N_19854);
xor U20159 (N_20159,N_19964,N_19913);
nand U20160 (N_20160,N_19753,N_19885);
nand U20161 (N_20161,N_19938,N_19898);
or U20162 (N_20162,N_19824,N_19997);
and U20163 (N_20163,N_19912,N_19953);
xnor U20164 (N_20164,N_19829,N_19877);
xor U20165 (N_20165,N_19914,N_19979);
xor U20166 (N_20166,N_19889,N_19920);
nand U20167 (N_20167,N_19846,N_19816);
and U20168 (N_20168,N_19782,N_19969);
or U20169 (N_20169,N_19829,N_19818);
xor U20170 (N_20170,N_19921,N_19805);
xnor U20171 (N_20171,N_19851,N_19996);
xnor U20172 (N_20172,N_19778,N_19960);
and U20173 (N_20173,N_19827,N_19820);
nor U20174 (N_20174,N_19874,N_19762);
nor U20175 (N_20175,N_19876,N_19981);
and U20176 (N_20176,N_19999,N_19995);
xor U20177 (N_20177,N_19869,N_19803);
or U20178 (N_20178,N_19766,N_19797);
nand U20179 (N_20179,N_19768,N_19962);
and U20180 (N_20180,N_19886,N_19765);
xnor U20181 (N_20181,N_19903,N_19780);
nand U20182 (N_20182,N_19994,N_19753);
or U20183 (N_20183,N_19772,N_19856);
and U20184 (N_20184,N_19943,N_19912);
nor U20185 (N_20185,N_19851,N_19788);
xor U20186 (N_20186,N_19880,N_19863);
and U20187 (N_20187,N_19773,N_19832);
and U20188 (N_20188,N_19974,N_19834);
and U20189 (N_20189,N_19978,N_19824);
nand U20190 (N_20190,N_19875,N_19978);
nor U20191 (N_20191,N_19978,N_19973);
nor U20192 (N_20192,N_19752,N_19764);
or U20193 (N_20193,N_19883,N_19979);
xnor U20194 (N_20194,N_19958,N_19929);
nor U20195 (N_20195,N_19970,N_19750);
and U20196 (N_20196,N_19943,N_19848);
xnor U20197 (N_20197,N_19879,N_19940);
nor U20198 (N_20198,N_19839,N_19999);
or U20199 (N_20199,N_19823,N_19884);
and U20200 (N_20200,N_19930,N_19835);
xor U20201 (N_20201,N_19824,N_19982);
xor U20202 (N_20202,N_19908,N_19847);
nand U20203 (N_20203,N_19778,N_19922);
or U20204 (N_20204,N_19877,N_19772);
nor U20205 (N_20205,N_19854,N_19769);
nand U20206 (N_20206,N_19873,N_19759);
or U20207 (N_20207,N_19863,N_19785);
and U20208 (N_20208,N_19950,N_19850);
nor U20209 (N_20209,N_19910,N_19835);
nor U20210 (N_20210,N_19823,N_19869);
and U20211 (N_20211,N_19802,N_19850);
xnor U20212 (N_20212,N_19869,N_19947);
xnor U20213 (N_20213,N_19794,N_19983);
nor U20214 (N_20214,N_19853,N_19926);
nor U20215 (N_20215,N_19950,N_19927);
xor U20216 (N_20216,N_19824,N_19767);
and U20217 (N_20217,N_19901,N_19915);
nor U20218 (N_20218,N_19844,N_19935);
nor U20219 (N_20219,N_19783,N_19819);
or U20220 (N_20220,N_19800,N_19955);
and U20221 (N_20221,N_19754,N_19805);
nor U20222 (N_20222,N_19926,N_19756);
and U20223 (N_20223,N_19753,N_19785);
xnor U20224 (N_20224,N_19899,N_19922);
nor U20225 (N_20225,N_19868,N_19926);
nor U20226 (N_20226,N_19784,N_19763);
and U20227 (N_20227,N_19980,N_19893);
and U20228 (N_20228,N_19874,N_19983);
and U20229 (N_20229,N_19925,N_19751);
or U20230 (N_20230,N_19930,N_19873);
nand U20231 (N_20231,N_19784,N_19802);
and U20232 (N_20232,N_19876,N_19755);
and U20233 (N_20233,N_19955,N_19961);
xnor U20234 (N_20234,N_19912,N_19774);
nor U20235 (N_20235,N_19801,N_19925);
or U20236 (N_20236,N_19797,N_19901);
nor U20237 (N_20237,N_19842,N_19759);
xor U20238 (N_20238,N_19806,N_19875);
xnor U20239 (N_20239,N_19959,N_19958);
xor U20240 (N_20240,N_19791,N_19887);
or U20241 (N_20241,N_19816,N_19792);
nand U20242 (N_20242,N_19798,N_19877);
or U20243 (N_20243,N_19792,N_19787);
and U20244 (N_20244,N_19855,N_19838);
or U20245 (N_20245,N_19839,N_19870);
xnor U20246 (N_20246,N_19835,N_19975);
and U20247 (N_20247,N_19759,N_19950);
and U20248 (N_20248,N_19918,N_19792);
nor U20249 (N_20249,N_19757,N_19826);
or U20250 (N_20250,N_20104,N_20184);
nor U20251 (N_20251,N_20171,N_20097);
or U20252 (N_20252,N_20223,N_20238);
nand U20253 (N_20253,N_20198,N_20149);
xnor U20254 (N_20254,N_20248,N_20233);
and U20255 (N_20255,N_20086,N_20058);
or U20256 (N_20256,N_20022,N_20009);
nand U20257 (N_20257,N_20066,N_20245);
or U20258 (N_20258,N_20016,N_20225);
nor U20259 (N_20259,N_20150,N_20134);
and U20260 (N_20260,N_20031,N_20051);
nand U20261 (N_20261,N_20242,N_20197);
xnor U20262 (N_20262,N_20012,N_20181);
xnor U20263 (N_20263,N_20115,N_20231);
nand U20264 (N_20264,N_20002,N_20214);
or U20265 (N_20265,N_20189,N_20083);
xor U20266 (N_20266,N_20064,N_20000);
nor U20267 (N_20267,N_20162,N_20121);
and U20268 (N_20268,N_20030,N_20174);
and U20269 (N_20269,N_20019,N_20176);
nand U20270 (N_20270,N_20026,N_20232);
xnor U20271 (N_20271,N_20216,N_20228);
nand U20272 (N_20272,N_20136,N_20156);
or U20273 (N_20273,N_20206,N_20201);
or U20274 (N_20274,N_20117,N_20032);
nand U20275 (N_20275,N_20109,N_20106);
nand U20276 (N_20276,N_20133,N_20240);
nand U20277 (N_20277,N_20132,N_20166);
nor U20278 (N_20278,N_20151,N_20160);
or U20279 (N_20279,N_20220,N_20173);
or U20280 (N_20280,N_20118,N_20027);
xor U20281 (N_20281,N_20013,N_20023);
xnor U20282 (N_20282,N_20138,N_20243);
nand U20283 (N_20283,N_20141,N_20237);
xnor U20284 (N_20284,N_20059,N_20247);
nand U20285 (N_20285,N_20089,N_20142);
or U20286 (N_20286,N_20050,N_20111);
and U20287 (N_20287,N_20192,N_20061);
or U20288 (N_20288,N_20124,N_20249);
nor U20289 (N_20289,N_20230,N_20036);
xor U20290 (N_20290,N_20195,N_20035);
nor U20291 (N_20291,N_20046,N_20208);
and U20292 (N_20292,N_20041,N_20018);
or U20293 (N_20293,N_20167,N_20082);
nand U20294 (N_20294,N_20053,N_20090);
nand U20295 (N_20295,N_20094,N_20112);
xor U20296 (N_20296,N_20123,N_20105);
or U20297 (N_20297,N_20054,N_20037);
and U20298 (N_20298,N_20034,N_20212);
and U20299 (N_20299,N_20049,N_20187);
or U20300 (N_20300,N_20017,N_20159);
nand U20301 (N_20301,N_20099,N_20244);
nor U20302 (N_20302,N_20199,N_20024);
and U20303 (N_20303,N_20003,N_20163);
and U20304 (N_20304,N_20188,N_20021);
or U20305 (N_20305,N_20144,N_20045);
nand U20306 (N_20306,N_20113,N_20088);
nand U20307 (N_20307,N_20186,N_20185);
or U20308 (N_20308,N_20219,N_20165);
or U20309 (N_20309,N_20081,N_20010);
xnor U20310 (N_20310,N_20127,N_20205);
xnor U20311 (N_20311,N_20043,N_20079);
nor U20312 (N_20312,N_20137,N_20029);
nor U20313 (N_20313,N_20011,N_20014);
nand U20314 (N_20314,N_20005,N_20147);
nor U20315 (N_20315,N_20221,N_20170);
and U20316 (N_20316,N_20075,N_20073);
nor U20317 (N_20317,N_20120,N_20067);
xnor U20318 (N_20318,N_20196,N_20047);
or U20319 (N_20319,N_20179,N_20152);
nand U20320 (N_20320,N_20103,N_20068);
and U20321 (N_20321,N_20204,N_20085);
and U20322 (N_20322,N_20241,N_20096);
or U20323 (N_20323,N_20114,N_20234);
xnor U20324 (N_20324,N_20055,N_20062);
nand U20325 (N_20325,N_20153,N_20190);
and U20326 (N_20326,N_20063,N_20169);
xor U20327 (N_20327,N_20191,N_20217);
nor U20328 (N_20328,N_20060,N_20007);
nand U20329 (N_20329,N_20227,N_20044);
xnor U20330 (N_20330,N_20071,N_20119);
xnor U20331 (N_20331,N_20056,N_20178);
nor U20332 (N_20332,N_20102,N_20177);
or U20333 (N_20333,N_20182,N_20135);
and U20334 (N_20334,N_20222,N_20125);
nor U20335 (N_20335,N_20207,N_20098);
or U20336 (N_20336,N_20004,N_20146);
or U20337 (N_20337,N_20130,N_20143);
xor U20338 (N_20338,N_20076,N_20048);
nand U20339 (N_20339,N_20140,N_20101);
and U20340 (N_20340,N_20084,N_20224);
and U20341 (N_20341,N_20052,N_20042);
nand U20342 (N_20342,N_20025,N_20200);
nor U20343 (N_20343,N_20038,N_20108);
or U20344 (N_20344,N_20065,N_20229);
or U20345 (N_20345,N_20092,N_20175);
nor U20346 (N_20346,N_20006,N_20057);
xor U20347 (N_20347,N_20039,N_20020);
and U20348 (N_20348,N_20116,N_20209);
nor U20349 (N_20349,N_20074,N_20239);
nor U20350 (N_20350,N_20033,N_20145);
and U20351 (N_20351,N_20131,N_20128);
nand U20352 (N_20352,N_20122,N_20211);
nand U20353 (N_20353,N_20235,N_20040);
and U20354 (N_20354,N_20087,N_20246);
and U20355 (N_20355,N_20100,N_20180);
xnor U20356 (N_20356,N_20139,N_20078);
nand U20357 (N_20357,N_20183,N_20213);
nor U20358 (N_20358,N_20226,N_20148);
xor U20359 (N_20359,N_20015,N_20210);
or U20360 (N_20360,N_20008,N_20129);
or U20361 (N_20361,N_20203,N_20093);
nand U20362 (N_20362,N_20028,N_20091);
nor U20363 (N_20363,N_20194,N_20215);
xnor U20364 (N_20364,N_20110,N_20168);
nor U20365 (N_20365,N_20157,N_20236);
xor U20366 (N_20366,N_20158,N_20070);
xor U20367 (N_20367,N_20172,N_20218);
or U20368 (N_20368,N_20155,N_20095);
xor U20369 (N_20369,N_20154,N_20069);
and U20370 (N_20370,N_20164,N_20080);
or U20371 (N_20371,N_20193,N_20001);
xor U20372 (N_20372,N_20072,N_20202);
nor U20373 (N_20373,N_20107,N_20126);
or U20374 (N_20374,N_20077,N_20161);
xnor U20375 (N_20375,N_20115,N_20056);
xnor U20376 (N_20376,N_20103,N_20056);
nand U20377 (N_20377,N_20146,N_20202);
nand U20378 (N_20378,N_20095,N_20176);
nor U20379 (N_20379,N_20071,N_20189);
xnor U20380 (N_20380,N_20014,N_20020);
or U20381 (N_20381,N_20013,N_20099);
nand U20382 (N_20382,N_20242,N_20065);
xnor U20383 (N_20383,N_20225,N_20058);
nor U20384 (N_20384,N_20011,N_20067);
or U20385 (N_20385,N_20154,N_20186);
nand U20386 (N_20386,N_20088,N_20132);
xor U20387 (N_20387,N_20187,N_20078);
and U20388 (N_20388,N_20173,N_20125);
nand U20389 (N_20389,N_20118,N_20140);
or U20390 (N_20390,N_20107,N_20214);
xor U20391 (N_20391,N_20177,N_20083);
or U20392 (N_20392,N_20003,N_20198);
nor U20393 (N_20393,N_20012,N_20199);
and U20394 (N_20394,N_20098,N_20140);
nor U20395 (N_20395,N_20004,N_20086);
and U20396 (N_20396,N_20085,N_20135);
xnor U20397 (N_20397,N_20098,N_20068);
nand U20398 (N_20398,N_20247,N_20034);
nand U20399 (N_20399,N_20134,N_20098);
or U20400 (N_20400,N_20123,N_20119);
or U20401 (N_20401,N_20129,N_20082);
xnor U20402 (N_20402,N_20116,N_20185);
nand U20403 (N_20403,N_20054,N_20124);
and U20404 (N_20404,N_20079,N_20111);
and U20405 (N_20405,N_20212,N_20176);
nand U20406 (N_20406,N_20225,N_20111);
and U20407 (N_20407,N_20201,N_20087);
or U20408 (N_20408,N_20143,N_20171);
and U20409 (N_20409,N_20119,N_20018);
xnor U20410 (N_20410,N_20011,N_20041);
or U20411 (N_20411,N_20078,N_20046);
xnor U20412 (N_20412,N_20020,N_20170);
nor U20413 (N_20413,N_20100,N_20125);
and U20414 (N_20414,N_20083,N_20138);
or U20415 (N_20415,N_20083,N_20182);
nor U20416 (N_20416,N_20003,N_20030);
or U20417 (N_20417,N_20092,N_20023);
xnor U20418 (N_20418,N_20022,N_20158);
nor U20419 (N_20419,N_20130,N_20202);
or U20420 (N_20420,N_20093,N_20212);
or U20421 (N_20421,N_20239,N_20223);
nand U20422 (N_20422,N_20184,N_20203);
nor U20423 (N_20423,N_20041,N_20187);
and U20424 (N_20424,N_20025,N_20090);
xor U20425 (N_20425,N_20069,N_20062);
xor U20426 (N_20426,N_20028,N_20152);
nor U20427 (N_20427,N_20114,N_20044);
xnor U20428 (N_20428,N_20125,N_20249);
nor U20429 (N_20429,N_20091,N_20163);
xnor U20430 (N_20430,N_20003,N_20179);
nor U20431 (N_20431,N_20003,N_20133);
or U20432 (N_20432,N_20137,N_20161);
and U20433 (N_20433,N_20125,N_20198);
or U20434 (N_20434,N_20085,N_20148);
nand U20435 (N_20435,N_20170,N_20146);
or U20436 (N_20436,N_20215,N_20243);
and U20437 (N_20437,N_20158,N_20121);
xor U20438 (N_20438,N_20099,N_20175);
or U20439 (N_20439,N_20082,N_20022);
nand U20440 (N_20440,N_20012,N_20242);
or U20441 (N_20441,N_20143,N_20004);
or U20442 (N_20442,N_20186,N_20092);
nor U20443 (N_20443,N_20041,N_20245);
nand U20444 (N_20444,N_20195,N_20058);
xor U20445 (N_20445,N_20173,N_20141);
or U20446 (N_20446,N_20169,N_20121);
xnor U20447 (N_20447,N_20100,N_20241);
nand U20448 (N_20448,N_20166,N_20154);
or U20449 (N_20449,N_20219,N_20223);
nand U20450 (N_20450,N_20218,N_20081);
xnor U20451 (N_20451,N_20225,N_20079);
nor U20452 (N_20452,N_20141,N_20048);
and U20453 (N_20453,N_20135,N_20079);
or U20454 (N_20454,N_20192,N_20076);
nand U20455 (N_20455,N_20204,N_20125);
and U20456 (N_20456,N_20008,N_20074);
xnor U20457 (N_20457,N_20065,N_20217);
or U20458 (N_20458,N_20025,N_20091);
and U20459 (N_20459,N_20008,N_20057);
and U20460 (N_20460,N_20034,N_20160);
nor U20461 (N_20461,N_20142,N_20008);
xor U20462 (N_20462,N_20066,N_20041);
nor U20463 (N_20463,N_20056,N_20090);
and U20464 (N_20464,N_20206,N_20230);
xor U20465 (N_20465,N_20021,N_20228);
nand U20466 (N_20466,N_20081,N_20024);
nand U20467 (N_20467,N_20001,N_20168);
or U20468 (N_20468,N_20235,N_20065);
or U20469 (N_20469,N_20215,N_20150);
nor U20470 (N_20470,N_20087,N_20207);
or U20471 (N_20471,N_20176,N_20071);
xor U20472 (N_20472,N_20022,N_20241);
or U20473 (N_20473,N_20069,N_20247);
nor U20474 (N_20474,N_20000,N_20104);
and U20475 (N_20475,N_20036,N_20234);
nand U20476 (N_20476,N_20110,N_20206);
and U20477 (N_20477,N_20208,N_20163);
or U20478 (N_20478,N_20076,N_20089);
and U20479 (N_20479,N_20237,N_20171);
xor U20480 (N_20480,N_20208,N_20184);
and U20481 (N_20481,N_20213,N_20170);
or U20482 (N_20482,N_20248,N_20070);
nand U20483 (N_20483,N_20161,N_20247);
xnor U20484 (N_20484,N_20132,N_20209);
xnor U20485 (N_20485,N_20150,N_20009);
nand U20486 (N_20486,N_20163,N_20022);
nor U20487 (N_20487,N_20222,N_20208);
nor U20488 (N_20488,N_20008,N_20091);
or U20489 (N_20489,N_20194,N_20156);
nor U20490 (N_20490,N_20055,N_20104);
xnor U20491 (N_20491,N_20152,N_20043);
nor U20492 (N_20492,N_20096,N_20169);
xor U20493 (N_20493,N_20087,N_20053);
xor U20494 (N_20494,N_20194,N_20012);
nor U20495 (N_20495,N_20147,N_20211);
or U20496 (N_20496,N_20073,N_20063);
nor U20497 (N_20497,N_20131,N_20140);
nand U20498 (N_20498,N_20059,N_20128);
or U20499 (N_20499,N_20018,N_20113);
or U20500 (N_20500,N_20312,N_20499);
nor U20501 (N_20501,N_20498,N_20339);
xor U20502 (N_20502,N_20300,N_20348);
nand U20503 (N_20503,N_20252,N_20428);
nand U20504 (N_20504,N_20250,N_20293);
or U20505 (N_20505,N_20266,N_20386);
and U20506 (N_20506,N_20264,N_20280);
or U20507 (N_20507,N_20257,N_20490);
or U20508 (N_20508,N_20469,N_20452);
nand U20509 (N_20509,N_20302,N_20290);
nand U20510 (N_20510,N_20425,N_20279);
xnor U20511 (N_20511,N_20430,N_20324);
nor U20512 (N_20512,N_20352,N_20396);
and U20513 (N_20513,N_20391,N_20400);
nor U20514 (N_20514,N_20294,N_20460);
and U20515 (N_20515,N_20454,N_20307);
or U20516 (N_20516,N_20416,N_20328);
or U20517 (N_20517,N_20314,N_20346);
nand U20518 (N_20518,N_20447,N_20433);
nor U20519 (N_20519,N_20390,N_20273);
and U20520 (N_20520,N_20381,N_20358);
or U20521 (N_20521,N_20253,N_20353);
and U20522 (N_20522,N_20341,N_20363);
and U20523 (N_20523,N_20393,N_20372);
xor U20524 (N_20524,N_20354,N_20464);
nor U20525 (N_20525,N_20449,N_20423);
xor U20526 (N_20526,N_20258,N_20301);
and U20527 (N_20527,N_20477,N_20255);
and U20528 (N_20528,N_20355,N_20376);
nor U20529 (N_20529,N_20407,N_20441);
or U20530 (N_20530,N_20344,N_20493);
or U20531 (N_20531,N_20395,N_20463);
nor U20532 (N_20532,N_20335,N_20359);
or U20533 (N_20533,N_20424,N_20459);
and U20534 (N_20534,N_20487,N_20458);
and U20535 (N_20535,N_20491,N_20329);
nand U20536 (N_20536,N_20436,N_20319);
and U20537 (N_20537,N_20313,N_20256);
xor U20538 (N_20538,N_20488,N_20369);
and U20539 (N_20539,N_20262,N_20326);
or U20540 (N_20540,N_20251,N_20412);
or U20541 (N_20541,N_20349,N_20289);
nand U20542 (N_20542,N_20343,N_20371);
nor U20543 (N_20543,N_20479,N_20385);
and U20544 (N_20544,N_20277,N_20299);
nand U20545 (N_20545,N_20271,N_20304);
and U20546 (N_20546,N_20404,N_20426);
or U20547 (N_20547,N_20429,N_20383);
nand U20548 (N_20548,N_20411,N_20380);
or U20549 (N_20549,N_20345,N_20443);
nor U20550 (N_20550,N_20492,N_20421);
xor U20551 (N_20551,N_20378,N_20461);
and U20552 (N_20552,N_20403,N_20422);
nand U20553 (N_20553,N_20288,N_20342);
and U20554 (N_20554,N_20496,N_20254);
nand U20555 (N_20555,N_20474,N_20432);
xor U20556 (N_20556,N_20274,N_20322);
xnor U20557 (N_20557,N_20309,N_20455);
nor U20558 (N_20558,N_20406,N_20413);
and U20559 (N_20559,N_20476,N_20286);
nor U20560 (N_20560,N_20350,N_20334);
nor U20561 (N_20561,N_20295,N_20483);
nor U20562 (N_20562,N_20442,N_20331);
or U20563 (N_20563,N_20445,N_20332);
or U20564 (N_20564,N_20473,N_20357);
or U20565 (N_20565,N_20269,N_20272);
and U20566 (N_20566,N_20471,N_20296);
xnor U20567 (N_20567,N_20306,N_20282);
or U20568 (N_20568,N_20472,N_20270);
xnor U20569 (N_20569,N_20318,N_20316);
nand U20570 (N_20570,N_20401,N_20291);
or U20571 (N_20571,N_20267,N_20420);
nand U20572 (N_20572,N_20340,N_20410);
and U20573 (N_20573,N_20261,N_20361);
or U20574 (N_20574,N_20408,N_20435);
nand U20575 (N_20575,N_20311,N_20275);
nor U20576 (N_20576,N_20480,N_20268);
xor U20577 (N_20577,N_20325,N_20482);
nor U20578 (N_20578,N_20418,N_20285);
xor U20579 (N_20579,N_20467,N_20281);
nand U20580 (N_20580,N_20494,N_20298);
xor U20581 (N_20581,N_20437,N_20481);
xor U20582 (N_20582,N_20405,N_20263);
nand U20583 (N_20583,N_20427,N_20305);
nand U20584 (N_20584,N_20387,N_20439);
nand U20585 (N_20585,N_20370,N_20453);
nor U20586 (N_20586,N_20475,N_20457);
and U20587 (N_20587,N_20392,N_20336);
or U20588 (N_20588,N_20497,N_20470);
or U20589 (N_20589,N_20402,N_20415);
nand U20590 (N_20590,N_20398,N_20362);
or U20591 (N_20591,N_20397,N_20260);
nor U20592 (N_20592,N_20434,N_20366);
or U20593 (N_20593,N_20446,N_20283);
and U20594 (N_20594,N_20409,N_20303);
and U20595 (N_20595,N_20373,N_20323);
and U20596 (N_20596,N_20259,N_20438);
and U20597 (N_20597,N_20310,N_20364);
nand U20598 (N_20598,N_20287,N_20478);
xnor U20599 (N_20599,N_20374,N_20388);
xnor U20600 (N_20600,N_20444,N_20347);
and U20601 (N_20601,N_20495,N_20360);
xnor U20602 (N_20602,N_20466,N_20375);
nor U20603 (N_20603,N_20484,N_20321);
or U20604 (N_20604,N_20394,N_20333);
xnor U20605 (N_20605,N_20382,N_20384);
nand U20606 (N_20606,N_20448,N_20489);
or U20607 (N_20607,N_20297,N_20417);
xor U20608 (N_20608,N_20337,N_20465);
nor U20609 (N_20609,N_20265,N_20414);
or U20610 (N_20610,N_20486,N_20338);
nand U20611 (N_20611,N_20351,N_20292);
and U20612 (N_20612,N_20419,N_20367);
and U20613 (N_20613,N_20451,N_20278);
xnor U20614 (N_20614,N_20327,N_20315);
and U20615 (N_20615,N_20276,N_20308);
xnor U20616 (N_20616,N_20330,N_20320);
and U20617 (N_20617,N_20317,N_20284);
and U20618 (N_20618,N_20456,N_20377);
nand U20619 (N_20619,N_20450,N_20368);
xnor U20620 (N_20620,N_20468,N_20365);
and U20621 (N_20621,N_20389,N_20399);
nand U20622 (N_20622,N_20379,N_20356);
and U20623 (N_20623,N_20485,N_20440);
nor U20624 (N_20624,N_20431,N_20462);
nor U20625 (N_20625,N_20479,N_20419);
and U20626 (N_20626,N_20348,N_20447);
and U20627 (N_20627,N_20498,N_20397);
xnor U20628 (N_20628,N_20342,N_20442);
nand U20629 (N_20629,N_20369,N_20387);
nand U20630 (N_20630,N_20468,N_20358);
nor U20631 (N_20631,N_20319,N_20332);
and U20632 (N_20632,N_20419,N_20348);
nor U20633 (N_20633,N_20274,N_20440);
or U20634 (N_20634,N_20263,N_20276);
and U20635 (N_20635,N_20344,N_20290);
or U20636 (N_20636,N_20287,N_20277);
and U20637 (N_20637,N_20320,N_20480);
and U20638 (N_20638,N_20409,N_20485);
xnor U20639 (N_20639,N_20377,N_20453);
xor U20640 (N_20640,N_20472,N_20386);
xor U20641 (N_20641,N_20344,N_20422);
and U20642 (N_20642,N_20329,N_20406);
xor U20643 (N_20643,N_20301,N_20382);
xnor U20644 (N_20644,N_20413,N_20488);
nor U20645 (N_20645,N_20270,N_20437);
xnor U20646 (N_20646,N_20396,N_20425);
nor U20647 (N_20647,N_20489,N_20493);
or U20648 (N_20648,N_20260,N_20371);
nor U20649 (N_20649,N_20422,N_20416);
or U20650 (N_20650,N_20421,N_20279);
or U20651 (N_20651,N_20320,N_20491);
and U20652 (N_20652,N_20371,N_20389);
xnor U20653 (N_20653,N_20438,N_20378);
nand U20654 (N_20654,N_20474,N_20270);
and U20655 (N_20655,N_20350,N_20421);
and U20656 (N_20656,N_20417,N_20273);
nand U20657 (N_20657,N_20387,N_20266);
xor U20658 (N_20658,N_20296,N_20350);
nor U20659 (N_20659,N_20494,N_20330);
nand U20660 (N_20660,N_20443,N_20414);
xnor U20661 (N_20661,N_20291,N_20460);
xnor U20662 (N_20662,N_20375,N_20326);
nor U20663 (N_20663,N_20259,N_20307);
nor U20664 (N_20664,N_20442,N_20251);
or U20665 (N_20665,N_20488,N_20426);
nand U20666 (N_20666,N_20374,N_20462);
or U20667 (N_20667,N_20389,N_20483);
nand U20668 (N_20668,N_20477,N_20374);
or U20669 (N_20669,N_20477,N_20313);
and U20670 (N_20670,N_20498,N_20279);
nand U20671 (N_20671,N_20393,N_20407);
and U20672 (N_20672,N_20260,N_20268);
or U20673 (N_20673,N_20367,N_20352);
or U20674 (N_20674,N_20489,N_20488);
and U20675 (N_20675,N_20469,N_20473);
nand U20676 (N_20676,N_20448,N_20479);
nand U20677 (N_20677,N_20461,N_20455);
nor U20678 (N_20678,N_20378,N_20264);
and U20679 (N_20679,N_20499,N_20303);
nor U20680 (N_20680,N_20318,N_20427);
and U20681 (N_20681,N_20383,N_20495);
and U20682 (N_20682,N_20261,N_20412);
nor U20683 (N_20683,N_20276,N_20372);
and U20684 (N_20684,N_20497,N_20339);
nand U20685 (N_20685,N_20415,N_20269);
xor U20686 (N_20686,N_20452,N_20450);
and U20687 (N_20687,N_20349,N_20278);
nand U20688 (N_20688,N_20307,N_20283);
and U20689 (N_20689,N_20255,N_20473);
xor U20690 (N_20690,N_20328,N_20320);
nand U20691 (N_20691,N_20406,N_20484);
or U20692 (N_20692,N_20480,N_20385);
xnor U20693 (N_20693,N_20410,N_20423);
or U20694 (N_20694,N_20362,N_20431);
or U20695 (N_20695,N_20372,N_20334);
or U20696 (N_20696,N_20493,N_20477);
or U20697 (N_20697,N_20372,N_20309);
and U20698 (N_20698,N_20355,N_20268);
nor U20699 (N_20699,N_20494,N_20417);
nand U20700 (N_20700,N_20470,N_20319);
or U20701 (N_20701,N_20425,N_20272);
xor U20702 (N_20702,N_20364,N_20262);
and U20703 (N_20703,N_20344,N_20308);
xnor U20704 (N_20704,N_20315,N_20441);
nor U20705 (N_20705,N_20363,N_20399);
or U20706 (N_20706,N_20477,N_20487);
and U20707 (N_20707,N_20310,N_20257);
xor U20708 (N_20708,N_20269,N_20497);
nand U20709 (N_20709,N_20444,N_20253);
and U20710 (N_20710,N_20370,N_20388);
nand U20711 (N_20711,N_20387,N_20416);
nand U20712 (N_20712,N_20382,N_20339);
or U20713 (N_20713,N_20300,N_20389);
or U20714 (N_20714,N_20324,N_20480);
and U20715 (N_20715,N_20459,N_20354);
xnor U20716 (N_20716,N_20462,N_20339);
nor U20717 (N_20717,N_20402,N_20489);
and U20718 (N_20718,N_20284,N_20390);
or U20719 (N_20719,N_20391,N_20338);
or U20720 (N_20720,N_20372,N_20287);
xnor U20721 (N_20721,N_20437,N_20434);
and U20722 (N_20722,N_20272,N_20477);
or U20723 (N_20723,N_20262,N_20324);
xnor U20724 (N_20724,N_20365,N_20298);
nand U20725 (N_20725,N_20288,N_20251);
xor U20726 (N_20726,N_20321,N_20461);
or U20727 (N_20727,N_20462,N_20470);
xor U20728 (N_20728,N_20320,N_20282);
nor U20729 (N_20729,N_20478,N_20490);
and U20730 (N_20730,N_20323,N_20328);
nor U20731 (N_20731,N_20375,N_20476);
or U20732 (N_20732,N_20357,N_20394);
xnor U20733 (N_20733,N_20394,N_20292);
and U20734 (N_20734,N_20268,N_20273);
nor U20735 (N_20735,N_20486,N_20287);
xnor U20736 (N_20736,N_20345,N_20376);
nor U20737 (N_20737,N_20283,N_20302);
nor U20738 (N_20738,N_20435,N_20267);
and U20739 (N_20739,N_20433,N_20317);
and U20740 (N_20740,N_20460,N_20412);
and U20741 (N_20741,N_20457,N_20468);
and U20742 (N_20742,N_20494,N_20485);
xor U20743 (N_20743,N_20495,N_20462);
xor U20744 (N_20744,N_20365,N_20296);
nor U20745 (N_20745,N_20315,N_20499);
and U20746 (N_20746,N_20356,N_20302);
and U20747 (N_20747,N_20492,N_20473);
nand U20748 (N_20748,N_20438,N_20328);
nor U20749 (N_20749,N_20460,N_20302);
or U20750 (N_20750,N_20501,N_20600);
nand U20751 (N_20751,N_20680,N_20529);
xor U20752 (N_20752,N_20579,N_20537);
nor U20753 (N_20753,N_20731,N_20748);
nand U20754 (N_20754,N_20690,N_20666);
or U20755 (N_20755,N_20715,N_20504);
and U20756 (N_20756,N_20611,N_20624);
nor U20757 (N_20757,N_20658,N_20694);
nor U20758 (N_20758,N_20638,N_20719);
xnor U20759 (N_20759,N_20635,N_20587);
or U20760 (N_20760,N_20558,N_20548);
and U20761 (N_20761,N_20502,N_20565);
nand U20762 (N_20762,N_20569,N_20514);
and U20763 (N_20763,N_20656,N_20683);
nor U20764 (N_20764,N_20653,N_20534);
xor U20765 (N_20765,N_20512,N_20516);
xor U20766 (N_20766,N_20636,N_20571);
xnor U20767 (N_20767,N_20519,N_20556);
nand U20768 (N_20768,N_20667,N_20745);
nor U20769 (N_20769,N_20539,N_20732);
xor U20770 (N_20770,N_20729,N_20520);
xor U20771 (N_20771,N_20621,N_20639);
or U20772 (N_20772,N_20524,N_20688);
or U20773 (N_20773,N_20597,N_20659);
nand U20774 (N_20774,N_20628,N_20612);
xnor U20775 (N_20775,N_20660,N_20640);
nand U20776 (N_20776,N_20541,N_20708);
and U20777 (N_20777,N_20623,N_20697);
nor U20778 (N_20778,N_20675,N_20677);
or U20779 (N_20779,N_20725,N_20546);
xnor U20780 (N_20780,N_20665,N_20506);
or U20781 (N_20781,N_20630,N_20509);
nand U20782 (N_20782,N_20596,N_20500);
nand U20783 (N_20783,N_20563,N_20610);
and U20784 (N_20784,N_20648,N_20695);
and U20785 (N_20785,N_20508,N_20625);
nand U20786 (N_20786,N_20654,N_20644);
nor U20787 (N_20787,N_20568,N_20613);
and U20788 (N_20788,N_20586,N_20560);
or U20789 (N_20789,N_20589,N_20723);
nand U20790 (N_20790,N_20521,N_20574);
nand U20791 (N_20791,N_20713,N_20605);
or U20792 (N_20792,N_20561,N_20669);
nand U20793 (N_20793,N_20535,N_20704);
and U20794 (N_20794,N_20622,N_20620);
or U20795 (N_20795,N_20661,N_20533);
and U20796 (N_20796,N_20646,N_20642);
or U20797 (N_20797,N_20671,N_20673);
nand U20798 (N_20798,N_20663,N_20550);
nand U20799 (N_20799,N_20637,N_20617);
nor U20800 (N_20800,N_20738,N_20627);
and U20801 (N_20801,N_20554,N_20701);
or U20802 (N_20802,N_20632,N_20581);
nor U20803 (N_20803,N_20517,N_20580);
xor U20804 (N_20804,N_20721,N_20538);
nand U20805 (N_20805,N_20532,N_20528);
nand U20806 (N_20806,N_20530,N_20536);
xnor U20807 (N_20807,N_20549,N_20607);
nor U20808 (N_20808,N_20650,N_20740);
or U20809 (N_20809,N_20712,N_20689);
and U20810 (N_20810,N_20647,N_20576);
nand U20811 (N_20811,N_20583,N_20547);
xor U20812 (N_20812,N_20746,N_20686);
or U20813 (N_20813,N_20573,N_20591);
nand U20814 (N_20814,N_20742,N_20649);
xnor U20815 (N_20815,N_20633,N_20720);
nand U20816 (N_20816,N_20747,N_20567);
xor U20817 (N_20817,N_20555,N_20737);
nand U20818 (N_20818,N_20590,N_20582);
or U20819 (N_20819,N_20734,N_20629);
nand U20820 (N_20820,N_20735,N_20657);
or U20821 (N_20821,N_20552,N_20749);
xor U20822 (N_20822,N_20526,N_20566);
nand U20823 (N_20823,N_20578,N_20736);
xnor U20824 (N_20824,N_20544,N_20743);
and U20825 (N_20825,N_20614,N_20684);
and U20826 (N_20826,N_20577,N_20739);
and U20827 (N_20827,N_20706,N_20730);
or U20828 (N_20828,N_20615,N_20601);
nor U20829 (N_20829,N_20559,N_20603);
xor U20830 (N_20830,N_20678,N_20726);
and U20831 (N_20831,N_20662,N_20540);
nand U20832 (N_20832,N_20513,N_20553);
nor U20833 (N_20833,N_20598,N_20592);
and U20834 (N_20834,N_20702,N_20733);
xnor U20835 (N_20835,N_20626,N_20588);
or U20836 (N_20836,N_20652,N_20542);
or U20837 (N_20837,N_20631,N_20602);
or U20838 (N_20838,N_20645,N_20584);
or U20839 (N_20839,N_20741,N_20608);
and U20840 (N_20840,N_20515,N_20672);
nand U20841 (N_20841,N_20545,N_20682);
and U20842 (N_20842,N_20510,N_20594);
and U20843 (N_20843,N_20685,N_20717);
or U20844 (N_20844,N_20655,N_20531);
xnor U20845 (N_20845,N_20505,N_20543);
or U20846 (N_20846,N_20709,N_20522);
and U20847 (N_20847,N_20705,N_20693);
and U20848 (N_20848,N_20507,N_20714);
or U20849 (N_20849,N_20595,N_20503);
nor U20850 (N_20850,N_20609,N_20616);
nand U20851 (N_20851,N_20681,N_20618);
or U20852 (N_20852,N_20728,N_20679);
or U20853 (N_20853,N_20716,N_20527);
nor U20854 (N_20854,N_20711,N_20619);
or U20855 (N_20855,N_20641,N_20700);
nor U20856 (N_20856,N_20724,N_20674);
nor U20857 (N_20857,N_20557,N_20643);
and U20858 (N_20858,N_20698,N_20718);
and U20859 (N_20859,N_20703,N_20692);
or U20860 (N_20860,N_20668,N_20518);
nor U20861 (N_20861,N_20523,N_20599);
nand U20862 (N_20862,N_20634,N_20593);
or U20863 (N_20863,N_20511,N_20562);
nand U20864 (N_20864,N_20676,N_20670);
and U20865 (N_20865,N_20604,N_20707);
xnor U20866 (N_20866,N_20722,N_20651);
or U20867 (N_20867,N_20710,N_20687);
or U20868 (N_20868,N_20664,N_20691);
and U20869 (N_20869,N_20572,N_20575);
xnor U20870 (N_20870,N_20551,N_20606);
nor U20871 (N_20871,N_20696,N_20727);
and U20872 (N_20872,N_20585,N_20525);
xnor U20873 (N_20873,N_20564,N_20699);
and U20874 (N_20874,N_20570,N_20744);
or U20875 (N_20875,N_20705,N_20614);
xnor U20876 (N_20876,N_20528,N_20698);
or U20877 (N_20877,N_20590,N_20524);
xnor U20878 (N_20878,N_20622,N_20698);
or U20879 (N_20879,N_20527,N_20614);
xor U20880 (N_20880,N_20710,N_20696);
or U20881 (N_20881,N_20663,N_20554);
nand U20882 (N_20882,N_20745,N_20645);
xor U20883 (N_20883,N_20564,N_20714);
xor U20884 (N_20884,N_20558,N_20637);
and U20885 (N_20885,N_20565,N_20680);
or U20886 (N_20886,N_20639,N_20562);
xnor U20887 (N_20887,N_20642,N_20719);
or U20888 (N_20888,N_20530,N_20528);
nand U20889 (N_20889,N_20652,N_20654);
or U20890 (N_20890,N_20570,N_20689);
nor U20891 (N_20891,N_20583,N_20627);
and U20892 (N_20892,N_20641,N_20621);
nor U20893 (N_20893,N_20530,N_20697);
nor U20894 (N_20894,N_20549,N_20537);
nor U20895 (N_20895,N_20631,N_20606);
or U20896 (N_20896,N_20701,N_20685);
xnor U20897 (N_20897,N_20716,N_20561);
and U20898 (N_20898,N_20716,N_20692);
nand U20899 (N_20899,N_20532,N_20510);
or U20900 (N_20900,N_20529,N_20606);
nor U20901 (N_20901,N_20524,N_20527);
nor U20902 (N_20902,N_20560,N_20716);
or U20903 (N_20903,N_20669,N_20547);
and U20904 (N_20904,N_20586,N_20641);
nand U20905 (N_20905,N_20742,N_20566);
and U20906 (N_20906,N_20745,N_20616);
and U20907 (N_20907,N_20548,N_20703);
nand U20908 (N_20908,N_20639,N_20528);
or U20909 (N_20909,N_20570,N_20715);
nor U20910 (N_20910,N_20519,N_20564);
xnor U20911 (N_20911,N_20598,N_20509);
nor U20912 (N_20912,N_20633,N_20511);
nand U20913 (N_20913,N_20638,N_20606);
xnor U20914 (N_20914,N_20704,N_20728);
and U20915 (N_20915,N_20637,N_20690);
xnor U20916 (N_20916,N_20674,N_20567);
nor U20917 (N_20917,N_20596,N_20714);
nor U20918 (N_20918,N_20608,N_20621);
and U20919 (N_20919,N_20689,N_20643);
xor U20920 (N_20920,N_20663,N_20649);
nand U20921 (N_20921,N_20514,N_20693);
or U20922 (N_20922,N_20608,N_20570);
nand U20923 (N_20923,N_20505,N_20617);
or U20924 (N_20924,N_20534,N_20564);
xnor U20925 (N_20925,N_20749,N_20520);
nor U20926 (N_20926,N_20702,N_20709);
nand U20927 (N_20927,N_20559,N_20598);
nand U20928 (N_20928,N_20529,N_20548);
and U20929 (N_20929,N_20575,N_20624);
nand U20930 (N_20930,N_20644,N_20631);
or U20931 (N_20931,N_20729,N_20564);
or U20932 (N_20932,N_20514,N_20511);
nor U20933 (N_20933,N_20506,N_20732);
nor U20934 (N_20934,N_20688,N_20711);
nor U20935 (N_20935,N_20749,N_20576);
xor U20936 (N_20936,N_20559,N_20680);
nor U20937 (N_20937,N_20583,N_20717);
nand U20938 (N_20938,N_20735,N_20596);
nor U20939 (N_20939,N_20743,N_20597);
or U20940 (N_20940,N_20728,N_20639);
nand U20941 (N_20941,N_20696,N_20639);
nand U20942 (N_20942,N_20748,N_20683);
and U20943 (N_20943,N_20629,N_20556);
and U20944 (N_20944,N_20535,N_20665);
nand U20945 (N_20945,N_20566,N_20715);
or U20946 (N_20946,N_20621,N_20704);
or U20947 (N_20947,N_20638,N_20501);
and U20948 (N_20948,N_20588,N_20717);
and U20949 (N_20949,N_20747,N_20576);
xor U20950 (N_20950,N_20638,N_20704);
xnor U20951 (N_20951,N_20623,N_20576);
nand U20952 (N_20952,N_20577,N_20559);
nor U20953 (N_20953,N_20557,N_20559);
nor U20954 (N_20954,N_20668,N_20587);
or U20955 (N_20955,N_20536,N_20687);
or U20956 (N_20956,N_20566,N_20677);
nor U20957 (N_20957,N_20747,N_20521);
xor U20958 (N_20958,N_20535,N_20614);
or U20959 (N_20959,N_20660,N_20606);
xnor U20960 (N_20960,N_20581,N_20523);
or U20961 (N_20961,N_20678,N_20590);
nand U20962 (N_20962,N_20645,N_20629);
nor U20963 (N_20963,N_20558,N_20723);
or U20964 (N_20964,N_20641,N_20557);
or U20965 (N_20965,N_20721,N_20675);
xnor U20966 (N_20966,N_20661,N_20681);
or U20967 (N_20967,N_20666,N_20511);
xor U20968 (N_20968,N_20628,N_20517);
and U20969 (N_20969,N_20749,N_20554);
nand U20970 (N_20970,N_20658,N_20514);
xor U20971 (N_20971,N_20542,N_20651);
and U20972 (N_20972,N_20654,N_20723);
or U20973 (N_20973,N_20579,N_20539);
xor U20974 (N_20974,N_20746,N_20658);
or U20975 (N_20975,N_20637,N_20664);
and U20976 (N_20976,N_20642,N_20639);
nor U20977 (N_20977,N_20597,N_20641);
and U20978 (N_20978,N_20532,N_20613);
or U20979 (N_20979,N_20712,N_20576);
and U20980 (N_20980,N_20546,N_20706);
or U20981 (N_20981,N_20560,N_20645);
nor U20982 (N_20982,N_20679,N_20508);
and U20983 (N_20983,N_20725,N_20612);
nand U20984 (N_20984,N_20565,N_20726);
nand U20985 (N_20985,N_20650,N_20687);
or U20986 (N_20986,N_20732,N_20727);
nor U20987 (N_20987,N_20567,N_20518);
and U20988 (N_20988,N_20652,N_20681);
and U20989 (N_20989,N_20543,N_20719);
and U20990 (N_20990,N_20687,N_20574);
xnor U20991 (N_20991,N_20522,N_20639);
nor U20992 (N_20992,N_20710,N_20745);
and U20993 (N_20993,N_20694,N_20591);
or U20994 (N_20994,N_20686,N_20606);
xor U20995 (N_20995,N_20689,N_20682);
nand U20996 (N_20996,N_20577,N_20699);
nor U20997 (N_20997,N_20745,N_20598);
nand U20998 (N_20998,N_20600,N_20634);
nor U20999 (N_20999,N_20725,N_20714);
nor U21000 (N_21000,N_20806,N_20962);
nor U21001 (N_21001,N_20927,N_20984);
and U21002 (N_21002,N_20968,N_20940);
nand U21003 (N_21003,N_20914,N_20773);
nand U21004 (N_21004,N_20793,N_20903);
nand U21005 (N_21005,N_20847,N_20807);
or U21006 (N_21006,N_20846,N_20926);
nand U21007 (N_21007,N_20804,N_20783);
or U21008 (N_21008,N_20976,N_20959);
nand U21009 (N_21009,N_20821,N_20960);
or U21010 (N_21010,N_20757,N_20994);
or U21011 (N_21011,N_20938,N_20974);
xor U21012 (N_21012,N_20859,N_20857);
nand U21013 (N_21013,N_20870,N_20890);
nand U21014 (N_21014,N_20751,N_20882);
or U21015 (N_21015,N_20839,N_20834);
nor U21016 (N_21016,N_20887,N_20812);
nand U21017 (N_21017,N_20969,N_20842);
nor U21018 (N_21018,N_20893,N_20860);
or U21019 (N_21019,N_20805,N_20851);
nand U21020 (N_21020,N_20843,N_20918);
or U21021 (N_21021,N_20845,N_20904);
and U21022 (N_21022,N_20767,N_20891);
and U21023 (N_21023,N_20786,N_20935);
nand U21024 (N_21024,N_20817,N_20791);
nor U21025 (N_21025,N_20928,N_20937);
nor U21026 (N_21026,N_20874,N_20779);
and U21027 (N_21027,N_20795,N_20753);
nor U21028 (N_21028,N_20957,N_20840);
or U21029 (N_21029,N_20983,N_20943);
or U21030 (N_21030,N_20979,N_20966);
or U21031 (N_21031,N_20799,N_20873);
or U21032 (N_21032,N_20796,N_20770);
xnor U21033 (N_21033,N_20958,N_20950);
nor U21034 (N_21034,N_20837,N_20929);
and U21035 (N_21035,N_20965,N_20765);
nor U21036 (N_21036,N_20856,N_20872);
and U21037 (N_21037,N_20869,N_20910);
nand U21038 (N_21038,N_20798,N_20861);
or U21039 (N_21039,N_20772,N_20794);
or U21040 (N_21040,N_20788,N_20768);
nor U21041 (N_21041,N_20780,N_20932);
and U21042 (N_21042,N_20972,N_20758);
nor U21043 (N_21043,N_20916,N_20769);
or U21044 (N_21044,N_20899,N_20792);
and U21045 (N_21045,N_20832,N_20921);
nor U21046 (N_21046,N_20999,N_20875);
or U21047 (N_21047,N_20951,N_20803);
or U21048 (N_21048,N_20800,N_20953);
and U21049 (N_21049,N_20895,N_20900);
or U21050 (N_21050,N_20920,N_20771);
xnor U21051 (N_21051,N_20970,N_20981);
nand U21052 (N_21052,N_20995,N_20930);
and U21053 (N_21053,N_20978,N_20977);
nor U21054 (N_21054,N_20942,N_20755);
nand U21055 (N_21055,N_20776,N_20853);
nor U21056 (N_21056,N_20975,N_20781);
and U21057 (N_21057,N_20876,N_20829);
nor U21058 (N_21058,N_20766,N_20801);
xnor U21059 (N_21059,N_20988,N_20892);
and U21060 (N_21060,N_20946,N_20863);
xor U21061 (N_21061,N_20990,N_20790);
nor U21062 (N_21062,N_20756,N_20764);
nand U21063 (N_21063,N_20858,N_20996);
nor U21064 (N_21064,N_20980,N_20924);
or U21065 (N_21065,N_20825,N_20964);
xnor U21066 (N_21066,N_20867,N_20778);
xnor U21067 (N_21067,N_20784,N_20868);
or U21068 (N_21068,N_20855,N_20952);
and U21069 (N_21069,N_20922,N_20949);
xor U21070 (N_21070,N_20917,N_20802);
nand U21071 (N_21071,N_20810,N_20787);
nand U21072 (N_21072,N_20998,N_20844);
nor U21073 (N_21073,N_20907,N_20831);
nor U21074 (N_21074,N_20886,N_20823);
nand U21075 (N_21075,N_20785,N_20775);
nand U21076 (N_21076,N_20815,N_20809);
and U21077 (N_21077,N_20912,N_20945);
nand U21078 (N_21078,N_20889,N_20885);
nand U21079 (N_21079,N_20936,N_20763);
nor U21080 (N_21080,N_20754,N_20985);
or U21081 (N_21081,N_20838,N_20987);
or U21082 (N_21082,N_20841,N_20854);
and U21083 (N_21083,N_20948,N_20866);
and U21084 (N_21084,N_20963,N_20818);
or U21085 (N_21085,N_20750,N_20849);
or U21086 (N_21086,N_20761,N_20789);
or U21087 (N_21087,N_20902,N_20947);
xnor U21088 (N_21088,N_20894,N_20967);
xor U21089 (N_21089,N_20816,N_20760);
xnor U21090 (N_21090,N_20880,N_20906);
nor U21091 (N_21091,N_20934,N_20782);
or U21092 (N_21092,N_20897,N_20797);
xor U21093 (N_21093,N_20811,N_20759);
nand U21094 (N_21094,N_20905,N_20898);
nand U21095 (N_21095,N_20955,N_20852);
or U21096 (N_21096,N_20956,N_20919);
nor U21097 (N_21097,N_20865,N_20909);
nand U21098 (N_21098,N_20774,N_20813);
or U21099 (N_21099,N_20835,N_20989);
and U21100 (N_21100,N_20993,N_20944);
and U21101 (N_21101,N_20991,N_20871);
nor U21102 (N_21102,N_20941,N_20884);
nand U21103 (N_21103,N_20819,N_20864);
and U21104 (N_21104,N_20814,N_20881);
nand U21105 (N_21105,N_20808,N_20822);
nor U21106 (N_21106,N_20836,N_20826);
nand U21107 (N_21107,N_20992,N_20828);
or U21108 (N_21108,N_20908,N_20762);
xnor U21109 (N_21109,N_20877,N_20827);
nand U21110 (N_21110,N_20830,N_20878);
and U21111 (N_21111,N_20777,N_20833);
or U21112 (N_21112,N_20901,N_20888);
and U21113 (N_21113,N_20883,N_20923);
or U21114 (N_21114,N_20925,N_20961);
xnor U21115 (N_21115,N_20896,N_20850);
and U21116 (N_21116,N_20982,N_20911);
or U21117 (N_21117,N_20931,N_20862);
nand U21118 (N_21118,N_20913,N_20939);
nand U21119 (N_21119,N_20997,N_20820);
nor U21120 (N_21120,N_20752,N_20879);
nand U21121 (N_21121,N_20986,N_20971);
nor U21122 (N_21122,N_20933,N_20973);
nand U21123 (N_21123,N_20915,N_20824);
nor U21124 (N_21124,N_20848,N_20954);
xnor U21125 (N_21125,N_20806,N_20755);
or U21126 (N_21126,N_20837,N_20860);
or U21127 (N_21127,N_20989,N_20854);
or U21128 (N_21128,N_20982,N_20975);
or U21129 (N_21129,N_20915,N_20944);
nand U21130 (N_21130,N_20942,N_20874);
or U21131 (N_21131,N_20900,N_20844);
nand U21132 (N_21132,N_20907,N_20864);
nor U21133 (N_21133,N_20915,N_20803);
xor U21134 (N_21134,N_20943,N_20782);
or U21135 (N_21135,N_20911,N_20788);
nor U21136 (N_21136,N_20853,N_20759);
nor U21137 (N_21137,N_20830,N_20936);
nand U21138 (N_21138,N_20863,N_20804);
and U21139 (N_21139,N_20875,N_20750);
nor U21140 (N_21140,N_20862,N_20892);
nor U21141 (N_21141,N_20838,N_20954);
nand U21142 (N_21142,N_20829,N_20788);
and U21143 (N_21143,N_20753,N_20761);
or U21144 (N_21144,N_20950,N_20858);
nand U21145 (N_21145,N_20977,N_20761);
nand U21146 (N_21146,N_20937,N_20959);
nor U21147 (N_21147,N_20849,N_20763);
nor U21148 (N_21148,N_20833,N_20864);
nor U21149 (N_21149,N_20971,N_20984);
or U21150 (N_21150,N_20795,N_20816);
xnor U21151 (N_21151,N_20874,N_20973);
xnor U21152 (N_21152,N_20968,N_20950);
nor U21153 (N_21153,N_20880,N_20966);
or U21154 (N_21154,N_20991,N_20920);
nand U21155 (N_21155,N_20933,N_20962);
nor U21156 (N_21156,N_20838,N_20898);
nand U21157 (N_21157,N_20784,N_20963);
nor U21158 (N_21158,N_20763,N_20793);
or U21159 (N_21159,N_20824,N_20903);
xnor U21160 (N_21160,N_20954,N_20921);
nor U21161 (N_21161,N_20819,N_20800);
or U21162 (N_21162,N_20777,N_20764);
nand U21163 (N_21163,N_20905,N_20936);
nor U21164 (N_21164,N_20939,N_20882);
or U21165 (N_21165,N_20814,N_20764);
nor U21166 (N_21166,N_20962,N_20971);
nor U21167 (N_21167,N_20870,N_20970);
xor U21168 (N_21168,N_20885,N_20960);
xor U21169 (N_21169,N_20809,N_20851);
xor U21170 (N_21170,N_20924,N_20753);
nor U21171 (N_21171,N_20887,N_20775);
and U21172 (N_21172,N_20888,N_20907);
nand U21173 (N_21173,N_20879,N_20871);
nor U21174 (N_21174,N_20881,N_20920);
xnor U21175 (N_21175,N_20940,N_20797);
and U21176 (N_21176,N_20959,N_20828);
nand U21177 (N_21177,N_20983,N_20802);
and U21178 (N_21178,N_20898,N_20815);
and U21179 (N_21179,N_20957,N_20834);
nand U21180 (N_21180,N_20919,N_20830);
and U21181 (N_21181,N_20985,N_20838);
and U21182 (N_21182,N_20805,N_20795);
nor U21183 (N_21183,N_20939,N_20813);
nor U21184 (N_21184,N_20995,N_20795);
nor U21185 (N_21185,N_20884,N_20945);
and U21186 (N_21186,N_20895,N_20771);
and U21187 (N_21187,N_20817,N_20770);
and U21188 (N_21188,N_20925,N_20885);
xnor U21189 (N_21189,N_20949,N_20840);
or U21190 (N_21190,N_20967,N_20972);
and U21191 (N_21191,N_20792,N_20776);
xor U21192 (N_21192,N_20792,N_20845);
or U21193 (N_21193,N_20955,N_20837);
nand U21194 (N_21194,N_20939,N_20988);
nand U21195 (N_21195,N_20875,N_20932);
and U21196 (N_21196,N_20939,N_20868);
nand U21197 (N_21197,N_20843,N_20943);
and U21198 (N_21198,N_20811,N_20843);
nand U21199 (N_21199,N_20899,N_20912);
or U21200 (N_21200,N_20788,N_20876);
or U21201 (N_21201,N_20982,N_20851);
xnor U21202 (N_21202,N_20938,N_20849);
xnor U21203 (N_21203,N_20763,N_20751);
and U21204 (N_21204,N_20926,N_20911);
nor U21205 (N_21205,N_20872,N_20971);
nor U21206 (N_21206,N_20783,N_20989);
nor U21207 (N_21207,N_20798,N_20819);
or U21208 (N_21208,N_20795,N_20803);
and U21209 (N_21209,N_20829,N_20976);
xnor U21210 (N_21210,N_20850,N_20946);
and U21211 (N_21211,N_20925,N_20774);
or U21212 (N_21212,N_20906,N_20964);
and U21213 (N_21213,N_20812,N_20978);
nand U21214 (N_21214,N_20959,N_20866);
xor U21215 (N_21215,N_20856,N_20877);
and U21216 (N_21216,N_20975,N_20836);
nand U21217 (N_21217,N_20964,N_20888);
or U21218 (N_21218,N_20858,N_20794);
nand U21219 (N_21219,N_20905,N_20821);
or U21220 (N_21220,N_20796,N_20987);
and U21221 (N_21221,N_20843,N_20870);
nand U21222 (N_21222,N_20800,N_20841);
or U21223 (N_21223,N_20873,N_20874);
and U21224 (N_21224,N_20891,N_20955);
or U21225 (N_21225,N_20990,N_20754);
nand U21226 (N_21226,N_20831,N_20979);
nand U21227 (N_21227,N_20823,N_20872);
and U21228 (N_21228,N_20967,N_20961);
nand U21229 (N_21229,N_20814,N_20924);
nor U21230 (N_21230,N_20791,N_20871);
nor U21231 (N_21231,N_20817,N_20940);
xnor U21232 (N_21232,N_20875,N_20788);
nor U21233 (N_21233,N_20956,N_20885);
nor U21234 (N_21234,N_20752,N_20777);
and U21235 (N_21235,N_20853,N_20820);
nor U21236 (N_21236,N_20769,N_20974);
nor U21237 (N_21237,N_20990,N_20891);
and U21238 (N_21238,N_20907,N_20792);
and U21239 (N_21239,N_20997,N_20795);
or U21240 (N_21240,N_20987,N_20821);
or U21241 (N_21241,N_20807,N_20876);
xnor U21242 (N_21242,N_20926,N_20932);
xnor U21243 (N_21243,N_20777,N_20942);
nand U21244 (N_21244,N_20816,N_20825);
nand U21245 (N_21245,N_20753,N_20991);
nor U21246 (N_21246,N_20894,N_20835);
xor U21247 (N_21247,N_20848,N_20930);
nor U21248 (N_21248,N_20962,N_20856);
nand U21249 (N_21249,N_20929,N_20882);
or U21250 (N_21250,N_21114,N_21053);
or U21251 (N_21251,N_21202,N_21017);
nor U21252 (N_21252,N_21227,N_21090);
nand U21253 (N_21253,N_21076,N_21146);
or U21254 (N_21254,N_21224,N_21191);
nor U21255 (N_21255,N_21074,N_21150);
xor U21256 (N_21256,N_21171,N_21080);
nand U21257 (N_21257,N_21218,N_21194);
nand U21258 (N_21258,N_21063,N_21046);
nand U21259 (N_21259,N_21144,N_21073);
xnor U21260 (N_21260,N_21098,N_21054);
xor U21261 (N_21261,N_21170,N_21044);
and U21262 (N_21262,N_21151,N_21147);
and U21263 (N_21263,N_21056,N_21031);
and U21264 (N_21264,N_21215,N_21152);
and U21265 (N_21265,N_21043,N_21200);
and U21266 (N_21266,N_21166,N_21084);
or U21267 (N_21267,N_21005,N_21030);
xor U21268 (N_21268,N_21069,N_21059);
nor U21269 (N_21269,N_21220,N_21101);
or U21270 (N_21270,N_21001,N_21235);
nand U21271 (N_21271,N_21123,N_21142);
nor U21272 (N_21272,N_21126,N_21103);
nand U21273 (N_21273,N_21110,N_21164);
nor U21274 (N_21274,N_21032,N_21217);
or U21275 (N_21275,N_21072,N_21230);
xnor U21276 (N_21276,N_21109,N_21118);
nor U21277 (N_21277,N_21130,N_21096);
nand U21278 (N_21278,N_21242,N_21003);
xnor U21279 (N_21279,N_21033,N_21189);
xnor U21280 (N_21280,N_21047,N_21165);
and U21281 (N_21281,N_21140,N_21183);
nor U21282 (N_21282,N_21248,N_21206);
nand U21283 (N_21283,N_21006,N_21068);
and U21284 (N_21284,N_21184,N_21111);
or U21285 (N_21285,N_21079,N_21014);
nand U21286 (N_21286,N_21214,N_21018);
and U21287 (N_21287,N_21040,N_21204);
xnor U21288 (N_21288,N_21015,N_21112);
nor U21289 (N_21289,N_21237,N_21244);
xor U21290 (N_21290,N_21163,N_21167);
and U21291 (N_21291,N_21102,N_21182);
xnor U21292 (N_21292,N_21061,N_21125);
or U21293 (N_21293,N_21203,N_21067);
nand U21294 (N_21294,N_21233,N_21105);
nor U21295 (N_21295,N_21197,N_21190);
or U21296 (N_21296,N_21236,N_21077);
or U21297 (N_21297,N_21120,N_21087);
or U21298 (N_21298,N_21023,N_21139);
nand U21299 (N_21299,N_21060,N_21249);
nor U21300 (N_21300,N_21134,N_21199);
nor U21301 (N_21301,N_21222,N_21036);
xnor U21302 (N_21302,N_21124,N_21231);
nor U21303 (N_21303,N_21177,N_21207);
nand U21304 (N_21304,N_21025,N_21135);
nor U21305 (N_21305,N_21116,N_21221);
nor U21306 (N_21306,N_21175,N_21119);
or U21307 (N_21307,N_21219,N_21121);
and U21308 (N_21308,N_21049,N_21095);
nand U21309 (N_21309,N_21172,N_21245);
or U21310 (N_21310,N_21195,N_21065);
or U21311 (N_21311,N_21037,N_21012);
nor U21312 (N_21312,N_21078,N_21137);
and U21313 (N_21313,N_21019,N_21066);
and U21314 (N_21314,N_21070,N_21192);
or U21315 (N_21315,N_21020,N_21161);
xor U21316 (N_21316,N_21106,N_21154);
nand U21317 (N_21317,N_21000,N_21026);
xnor U21318 (N_21318,N_21100,N_21108);
or U21319 (N_21319,N_21062,N_21243);
or U21320 (N_21320,N_21010,N_21246);
nand U21321 (N_21321,N_21193,N_21013);
and U21322 (N_21322,N_21022,N_21082);
nor U21323 (N_21323,N_21145,N_21158);
nand U21324 (N_21324,N_21050,N_21099);
or U21325 (N_21325,N_21104,N_21240);
nor U21326 (N_21326,N_21028,N_21041);
nor U21327 (N_21327,N_21174,N_21122);
and U21328 (N_21328,N_21086,N_21058);
and U21329 (N_21329,N_21178,N_21093);
and U21330 (N_21330,N_21129,N_21107);
nand U21331 (N_21331,N_21034,N_21075);
and U21332 (N_21332,N_21148,N_21016);
or U21333 (N_21333,N_21160,N_21132);
nor U21334 (N_21334,N_21157,N_21051);
or U21335 (N_21335,N_21039,N_21057);
and U21336 (N_21336,N_21186,N_21127);
or U21337 (N_21337,N_21173,N_21210);
and U21338 (N_21338,N_21064,N_21185);
nor U21339 (N_21339,N_21029,N_21089);
nor U21340 (N_21340,N_21117,N_21238);
nand U21341 (N_21341,N_21212,N_21187);
or U21342 (N_21342,N_21228,N_21027);
nand U21343 (N_21343,N_21223,N_21247);
nand U21344 (N_21344,N_21181,N_21113);
nor U21345 (N_21345,N_21226,N_21138);
and U21346 (N_21346,N_21209,N_21133);
nand U21347 (N_21347,N_21168,N_21198);
xnor U21348 (N_21348,N_21241,N_21035);
xnor U21349 (N_21349,N_21004,N_21211);
and U21350 (N_21350,N_21169,N_21196);
or U21351 (N_21351,N_21131,N_21055);
nand U21352 (N_21352,N_21052,N_21143);
nand U21353 (N_21353,N_21225,N_21085);
nor U21354 (N_21354,N_21071,N_21011);
nor U21355 (N_21355,N_21081,N_21149);
nand U21356 (N_21356,N_21156,N_21179);
or U21357 (N_21357,N_21216,N_21136);
nand U21358 (N_21358,N_21083,N_21205);
nor U21359 (N_21359,N_21176,N_21159);
xor U21360 (N_21360,N_21092,N_21024);
or U21361 (N_21361,N_21021,N_21097);
and U21362 (N_21362,N_21091,N_21048);
or U21363 (N_21363,N_21232,N_21008);
and U21364 (N_21364,N_21229,N_21201);
and U21365 (N_21365,N_21239,N_21155);
or U21366 (N_21366,N_21213,N_21038);
nand U21367 (N_21367,N_21088,N_21234);
or U21368 (N_21368,N_21162,N_21208);
xnor U21369 (N_21369,N_21042,N_21188);
and U21370 (N_21370,N_21094,N_21115);
nor U21371 (N_21371,N_21153,N_21128);
xor U21372 (N_21372,N_21180,N_21007);
nor U21373 (N_21373,N_21009,N_21141);
xor U21374 (N_21374,N_21002,N_21045);
xnor U21375 (N_21375,N_21162,N_21177);
nor U21376 (N_21376,N_21093,N_21051);
or U21377 (N_21377,N_21238,N_21083);
xnor U21378 (N_21378,N_21056,N_21142);
xnor U21379 (N_21379,N_21130,N_21153);
nand U21380 (N_21380,N_21213,N_21097);
or U21381 (N_21381,N_21188,N_21144);
or U21382 (N_21382,N_21103,N_21129);
and U21383 (N_21383,N_21097,N_21198);
or U21384 (N_21384,N_21180,N_21207);
nor U21385 (N_21385,N_21223,N_21070);
xnor U21386 (N_21386,N_21194,N_21161);
xor U21387 (N_21387,N_21223,N_21068);
and U21388 (N_21388,N_21030,N_21019);
and U21389 (N_21389,N_21168,N_21186);
xor U21390 (N_21390,N_21192,N_21008);
xnor U21391 (N_21391,N_21225,N_21119);
and U21392 (N_21392,N_21123,N_21213);
nand U21393 (N_21393,N_21228,N_21031);
xor U21394 (N_21394,N_21229,N_21133);
or U21395 (N_21395,N_21137,N_21231);
nand U21396 (N_21396,N_21014,N_21065);
nor U21397 (N_21397,N_21041,N_21246);
or U21398 (N_21398,N_21065,N_21133);
nor U21399 (N_21399,N_21040,N_21033);
nor U21400 (N_21400,N_21173,N_21106);
nand U21401 (N_21401,N_21117,N_21004);
nand U21402 (N_21402,N_21199,N_21030);
or U21403 (N_21403,N_21108,N_21116);
or U21404 (N_21404,N_21126,N_21117);
or U21405 (N_21405,N_21125,N_21075);
or U21406 (N_21406,N_21089,N_21125);
nand U21407 (N_21407,N_21165,N_21200);
and U21408 (N_21408,N_21048,N_21114);
nor U21409 (N_21409,N_21218,N_21135);
xnor U21410 (N_21410,N_21173,N_21227);
xnor U21411 (N_21411,N_21071,N_21193);
nand U21412 (N_21412,N_21086,N_21063);
xor U21413 (N_21413,N_21198,N_21165);
nand U21414 (N_21414,N_21121,N_21227);
xnor U21415 (N_21415,N_21176,N_21226);
xnor U21416 (N_21416,N_21053,N_21039);
and U21417 (N_21417,N_21239,N_21029);
nand U21418 (N_21418,N_21237,N_21168);
and U21419 (N_21419,N_21170,N_21237);
xor U21420 (N_21420,N_21216,N_21011);
nand U21421 (N_21421,N_21243,N_21106);
xnor U21422 (N_21422,N_21138,N_21195);
or U21423 (N_21423,N_21148,N_21215);
and U21424 (N_21424,N_21223,N_21225);
xor U21425 (N_21425,N_21041,N_21157);
or U21426 (N_21426,N_21108,N_21120);
or U21427 (N_21427,N_21163,N_21138);
nor U21428 (N_21428,N_21036,N_21160);
or U21429 (N_21429,N_21066,N_21162);
xnor U21430 (N_21430,N_21041,N_21059);
nand U21431 (N_21431,N_21151,N_21120);
nand U21432 (N_21432,N_21129,N_21196);
nor U21433 (N_21433,N_21213,N_21192);
and U21434 (N_21434,N_21242,N_21109);
nor U21435 (N_21435,N_21160,N_21112);
nand U21436 (N_21436,N_21093,N_21120);
or U21437 (N_21437,N_21110,N_21081);
nand U21438 (N_21438,N_21223,N_21147);
nor U21439 (N_21439,N_21000,N_21043);
or U21440 (N_21440,N_21209,N_21174);
nor U21441 (N_21441,N_21056,N_21070);
and U21442 (N_21442,N_21002,N_21155);
or U21443 (N_21443,N_21042,N_21045);
nor U21444 (N_21444,N_21021,N_21020);
nand U21445 (N_21445,N_21212,N_21176);
xor U21446 (N_21446,N_21015,N_21111);
xor U21447 (N_21447,N_21129,N_21046);
nand U21448 (N_21448,N_21156,N_21067);
and U21449 (N_21449,N_21109,N_21092);
or U21450 (N_21450,N_21094,N_21004);
nand U21451 (N_21451,N_21239,N_21172);
xnor U21452 (N_21452,N_21098,N_21053);
and U21453 (N_21453,N_21218,N_21078);
or U21454 (N_21454,N_21126,N_21083);
nand U21455 (N_21455,N_21001,N_21116);
xor U21456 (N_21456,N_21049,N_21127);
nor U21457 (N_21457,N_21141,N_21069);
and U21458 (N_21458,N_21174,N_21038);
nand U21459 (N_21459,N_21135,N_21114);
and U21460 (N_21460,N_21109,N_21200);
and U21461 (N_21461,N_21229,N_21058);
xnor U21462 (N_21462,N_21197,N_21186);
and U21463 (N_21463,N_21117,N_21122);
and U21464 (N_21464,N_21169,N_21116);
or U21465 (N_21465,N_21244,N_21227);
or U21466 (N_21466,N_21227,N_21011);
nand U21467 (N_21467,N_21109,N_21102);
or U21468 (N_21468,N_21160,N_21212);
xnor U21469 (N_21469,N_21171,N_21168);
xnor U21470 (N_21470,N_21164,N_21101);
nor U21471 (N_21471,N_21141,N_21066);
or U21472 (N_21472,N_21112,N_21006);
nor U21473 (N_21473,N_21101,N_21188);
nand U21474 (N_21474,N_21186,N_21228);
xor U21475 (N_21475,N_21122,N_21107);
and U21476 (N_21476,N_21097,N_21118);
xnor U21477 (N_21477,N_21215,N_21218);
or U21478 (N_21478,N_21197,N_21130);
nor U21479 (N_21479,N_21166,N_21225);
and U21480 (N_21480,N_21207,N_21066);
and U21481 (N_21481,N_21106,N_21130);
nor U21482 (N_21482,N_21229,N_21161);
and U21483 (N_21483,N_21200,N_21015);
and U21484 (N_21484,N_21110,N_21097);
nor U21485 (N_21485,N_21139,N_21082);
nand U21486 (N_21486,N_21147,N_21225);
xor U21487 (N_21487,N_21102,N_21237);
and U21488 (N_21488,N_21232,N_21011);
xnor U21489 (N_21489,N_21106,N_21131);
and U21490 (N_21490,N_21181,N_21178);
xor U21491 (N_21491,N_21145,N_21058);
nor U21492 (N_21492,N_21100,N_21171);
nand U21493 (N_21493,N_21207,N_21225);
and U21494 (N_21494,N_21161,N_21181);
or U21495 (N_21495,N_21097,N_21081);
and U21496 (N_21496,N_21231,N_21032);
or U21497 (N_21497,N_21086,N_21049);
xnor U21498 (N_21498,N_21165,N_21009);
xnor U21499 (N_21499,N_21226,N_21143);
xor U21500 (N_21500,N_21419,N_21444);
or U21501 (N_21501,N_21317,N_21445);
nor U21502 (N_21502,N_21499,N_21463);
nor U21503 (N_21503,N_21433,N_21399);
xor U21504 (N_21504,N_21353,N_21251);
nor U21505 (N_21505,N_21367,N_21314);
or U21506 (N_21506,N_21359,N_21405);
and U21507 (N_21507,N_21311,N_21328);
nand U21508 (N_21508,N_21360,N_21490);
xnor U21509 (N_21509,N_21392,N_21466);
nand U21510 (N_21510,N_21361,N_21436);
xor U21511 (N_21511,N_21291,N_21438);
xor U21512 (N_21512,N_21269,N_21415);
nand U21513 (N_21513,N_21297,N_21351);
nand U21514 (N_21514,N_21458,N_21322);
nor U21515 (N_21515,N_21364,N_21397);
or U21516 (N_21516,N_21471,N_21497);
and U21517 (N_21517,N_21274,N_21289);
and U21518 (N_21518,N_21264,N_21315);
or U21519 (N_21519,N_21409,N_21293);
nor U21520 (N_21520,N_21334,N_21395);
and U21521 (N_21521,N_21457,N_21262);
nor U21522 (N_21522,N_21331,N_21414);
xnor U21523 (N_21523,N_21485,N_21418);
nor U21524 (N_21524,N_21330,N_21365);
and U21525 (N_21525,N_21337,N_21381);
or U21526 (N_21526,N_21408,N_21451);
and U21527 (N_21527,N_21257,N_21336);
nand U21528 (N_21528,N_21493,N_21424);
or U21529 (N_21529,N_21373,N_21390);
nand U21530 (N_21530,N_21253,N_21344);
or U21531 (N_21531,N_21265,N_21413);
nor U21532 (N_21532,N_21431,N_21343);
nand U21533 (N_21533,N_21294,N_21271);
nand U21534 (N_21534,N_21400,N_21372);
nand U21535 (N_21535,N_21292,N_21290);
and U21536 (N_21536,N_21422,N_21449);
and U21537 (N_21537,N_21350,N_21358);
nand U21538 (N_21538,N_21492,N_21455);
or U21539 (N_21539,N_21299,N_21446);
and U21540 (N_21540,N_21308,N_21417);
or U21541 (N_21541,N_21430,N_21281);
xor U21542 (N_21542,N_21491,N_21377);
nor U21543 (N_21543,N_21420,N_21263);
and U21544 (N_21544,N_21355,N_21439);
or U21545 (N_21545,N_21326,N_21329);
nor U21546 (N_21546,N_21483,N_21488);
and U21547 (N_21547,N_21324,N_21283);
or U21548 (N_21548,N_21478,N_21305);
xor U21549 (N_21549,N_21423,N_21440);
nor U21550 (N_21550,N_21312,N_21345);
xnor U21551 (N_21551,N_21270,N_21354);
nand U21552 (N_21552,N_21432,N_21303);
or U21553 (N_21553,N_21278,N_21277);
xor U21554 (N_21554,N_21272,N_21412);
xor U21555 (N_21555,N_21429,N_21275);
xnor U21556 (N_21556,N_21452,N_21487);
or U21557 (N_21557,N_21321,N_21309);
nor U21558 (N_21558,N_21260,N_21407);
xnor U21559 (N_21559,N_21347,N_21482);
xor U21560 (N_21560,N_21472,N_21267);
nand U21561 (N_21561,N_21443,N_21301);
nand U21562 (N_21562,N_21268,N_21435);
and U21563 (N_21563,N_21398,N_21302);
and U21564 (N_21564,N_21475,N_21374);
or U21565 (N_21565,N_21284,N_21421);
nor U21566 (N_21566,N_21286,N_21468);
nand U21567 (N_21567,N_21348,N_21287);
nor U21568 (N_21568,N_21363,N_21403);
nand U21569 (N_21569,N_21448,N_21496);
nand U21570 (N_21570,N_21410,N_21335);
nand U21571 (N_21571,N_21319,N_21416);
or U21572 (N_21572,N_21386,N_21349);
nor U21573 (N_21573,N_21387,N_21474);
nand U21574 (N_21574,N_21383,N_21484);
xnor U21575 (N_21575,N_21323,N_21279);
xor U21576 (N_21576,N_21385,N_21467);
and U21577 (N_21577,N_21261,N_21368);
and U21578 (N_21578,N_21434,N_21252);
nor U21579 (N_21579,N_21453,N_21380);
or U21580 (N_21580,N_21425,N_21307);
xor U21581 (N_21581,N_21370,N_21406);
nor U21582 (N_21582,N_21295,N_21288);
xnor U21583 (N_21583,N_21428,N_21391);
and U21584 (N_21584,N_21459,N_21357);
and U21585 (N_21585,N_21376,N_21481);
nand U21586 (N_21586,N_21285,N_21341);
or U21587 (N_21587,N_21402,N_21476);
and U21588 (N_21588,N_21450,N_21469);
or U21589 (N_21589,N_21282,N_21366);
nand U21590 (N_21590,N_21300,N_21494);
nand U21591 (N_21591,N_21339,N_21441);
xnor U21592 (N_21592,N_21427,N_21479);
or U21593 (N_21593,N_21460,N_21384);
xor U21594 (N_21594,N_21379,N_21498);
and U21595 (N_21595,N_21382,N_21352);
nand U21596 (N_21596,N_21325,N_21371);
xnor U21597 (N_21597,N_21259,N_21495);
or U21598 (N_21598,N_21276,N_21346);
nor U21599 (N_21599,N_21470,N_21394);
nand U21600 (N_21600,N_21333,N_21316);
or U21601 (N_21601,N_21369,N_21393);
or U21602 (N_21602,N_21356,N_21456);
or U21603 (N_21603,N_21465,N_21426);
xnor U21604 (N_21604,N_21462,N_21486);
and U21605 (N_21605,N_21362,N_21280);
or U21606 (N_21606,N_21310,N_21298);
nor U21607 (N_21607,N_21461,N_21375);
nor U21608 (N_21608,N_21258,N_21388);
or U21609 (N_21609,N_21332,N_21254);
nand U21610 (N_21610,N_21342,N_21273);
or U21611 (N_21611,N_21296,N_21454);
and U21612 (N_21612,N_21340,N_21306);
and U21613 (N_21613,N_21396,N_21338);
and U21614 (N_21614,N_21473,N_21477);
nor U21615 (N_21615,N_21304,N_21442);
and U21616 (N_21616,N_21489,N_21437);
xor U21617 (N_21617,N_21464,N_21389);
or U21618 (N_21618,N_21401,N_21313);
nor U21619 (N_21619,N_21378,N_21320);
nand U21620 (N_21620,N_21266,N_21250);
or U21621 (N_21621,N_21411,N_21318);
and U21622 (N_21622,N_21447,N_21404);
and U21623 (N_21623,N_21256,N_21255);
and U21624 (N_21624,N_21327,N_21480);
nor U21625 (N_21625,N_21419,N_21434);
or U21626 (N_21626,N_21397,N_21253);
nor U21627 (N_21627,N_21339,N_21276);
and U21628 (N_21628,N_21324,N_21442);
xor U21629 (N_21629,N_21407,N_21351);
nand U21630 (N_21630,N_21256,N_21320);
or U21631 (N_21631,N_21383,N_21448);
and U21632 (N_21632,N_21435,N_21358);
xnor U21633 (N_21633,N_21305,N_21463);
or U21634 (N_21634,N_21438,N_21406);
and U21635 (N_21635,N_21251,N_21252);
or U21636 (N_21636,N_21330,N_21441);
nor U21637 (N_21637,N_21325,N_21465);
nand U21638 (N_21638,N_21409,N_21253);
and U21639 (N_21639,N_21352,N_21359);
and U21640 (N_21640,N_21480,N_21358);
xnor U21641 (N_21641,N_21403,N_21308);
xor U21642 (N_21642,N_21406,N_21361);
nand U21643 (N_21643,N_21344,N_21446);
xor U21644 (N_21644,N_21336,N_21356);
nor U21645 (N_21645,N_21420,N_21481);
and U21646 (N_21646,N_21426,N_21307);
nor U21647 (N_21647,N_21460,N_21269);
and U21648 (N_21648,N_21426,N_21342);
and U21649 (N_21649,N_21485,N_21360);
nand U21650 (N_21650,N_21276,N_21277);
nor U21651 (N_21651,N_21499,N_21373);
and U21652 (N_21652,N_21310,N_21449);
nand U21653 (N_21653,N_21250,N_21492);
nor U21654 (N_21654,N_21336,N_21404);
nand U21655 (N_21655,N_21476,N_21491);
nand U21656 (N_21656,N_21417,N_21441);
xor U21657 (N_21657,N_21287,N_21264);
and U21658 (N_21658,N_21271,N_21360);
nor U21659 (N_21659,N_21341,N_21335);
xor U21660 (N_21660,N_21268,N_21471);
xor U21661 (N_21661,N_21397,N_21441);
xor U21662 (N_21662,N_21287,N_21278);
xor U21663 (N_21663,N_21459,N_21294);
and U21664 (N_21664,N_21499,N_21300);
or U21665 (N_21665,N_21365,N_21358);
and U21666 (N_21666,N_21455,N_21473);
or U21667 (N_21667,N_21311,N_21386);
xnor U21668 (N_21668,N_21350,N_21291);
xnor U21669 (N_21669,N_21463,N_21346);
nand U21670 (N_21670,N_21476,N_21251);
or U21671 (N_21671,N_21447,N_21476);
xnor U21672 (N_21672,N_21423,N_21340);
nand U21673 (N_21673,N_21363,N_21491);
and U21674 (N_21674,N_21275,N_21417);
and U21675 (N_21675,N_21376,N_21350);
nor U21676 (N_21676,N_21490,N_21339);
and U21677 (N_21677,N_21345,N_21307);
nor U21678 (N_21678,N_21404,N_21327);
nand U21679 (N_21679,N_21386,N_21416);
and U21680 (N_21680,N_21323,N_21459);
nand U21681 (N_21681,N_21305,N_21484);
xnor U21682 (N_21682,N_21366,N_21328);
and U21683 (N_21683,N_21431,N_21479);
nand U21684 (N_21684,N_21349,N_21341);
or U21685 (N_21685,N_21289,N_21414);
nand U21686 (N_21686,N_21395,N_21326);
nand U21687 (N_21687,N_21477,N_21376);
nand U21688 (N_21688,N_21293,N_21337);
or U21689 (N_21689,N_21291,N_21491);
nor U21690 (N_21690,N_21373,N_21404);
xor U21691 (N_21691,N_21309,N_21307);
nor U21692 (N_21692,N_21352,N_21367);
or U21693 (N_21693,N_21252,N_21443);
nor U21694 (N_21694,N_21495,N_21329);
nand U21695 (N_21695,N_21493,N_21477);
nand U21696 (N_21696,N_21261,N_21434);
or U21697 (N_21697,N_21303,N_21433);
and U21698 (N_21698,N_21490,N_21472);
or U21699 (N_21699,N_21321,N_21346);
or U21700 (N_21700,N_21464,N_21494);
or U21701 (N_21701,N_21498,N_21340);
nor U21702 (N_21702,N_21336,N_21286);
nand U21703 (N_21703,N_21496,N_21475);
and U21704 (N_21704,N_21275,N_21390);
nand U21705 (N_21705,N_21467,N_21280);
nor U21706 (N_21706,N_21495,N_21473);
nand U21707 (N_21707,N_21349,N_21434);
and U21708 (N_21708,N_21412,N_21299);
or U21709 (N_21709,N_21331,N_21468);
nand U21710 (N_21710,N_21327,N_21309);
and U21711 (N_21711,N_21477,N_21362);
and U21712 (N_21712,N_21327,N_21269);
and U21713 (N_21713,N_21328,N_21327);
xor U21714 (N_21714,N_21338,N_21316);
or U21715 (N_21715,N_21275,N_21320);
and U21716 (N_21716,N_21327,N_21413);
xnor U21717 (N_21717,N_21453,N_21288);
nor U21718 (N_21718,N_21338,N_21292);
nor U21719 (N_21719,N_21466,N_21419);
nor U21720 (N_21720,N_21286,N_21290);
and U21721 (N_21721,N_21441,N_21292);
nand U21722 (N_21722,N_21485,N_21428);
nor U21723 (N_21723,N_21473,N_21287);
or U21724 (N_21724,N_21496,N_21446);
nand U21725 (N_21725,N_21434,N_21495);
or U21726 (N_21726,N_21339,N_21491);
or U21727 (N_21727,N_21414,N_21423);
nor U21728 (N_21728,N_21486,N_21403);
nor U21729 (N_21729,N_21272,N_21331);
xor U21730 (N_21730,N_21260,N_21434);
xor U21731 (N_21731,N_21337,N_21452);
or U21732 (N_21732,N_21273,N_21461);
and U21733 (N_21733,N_21429,N_21365);
nand U21734 (N_21734,N_21492,N_21269);
nand U21735 (N_21735,N_21294,N_21326);
nor U21736 (N_21736,N_21388,N_21255);
xnor U21737 (N_21737,N_21296,N_21344);
nor U21738 (N_21738,N_21432,N_21310);
or U21739 (N_21739,N_21362,N_21490);
nor U21740 (N_21740,N_21321,N_21271);
xnor U21741 (N_21741,N_21284,N_21258);
or U21742 (N_21742,N_21441,N_21306);
nand U21743 (N_21743,N_21495,N_21263);
nand U21744 (N_21744,N_21436,N_21417);
and U21745 (N_21745,N_21473,N_21317);
nor U21746 (N_21746,N_21453,N_21438);
xnor U21747 (N_21747,N_21465,N_21340);
and U21748 (N_21748,N_21466,N_21351);
nor U21749 (N_21749,N_21330,N_21282);
xor U21750 (N_21750,N_21502,N_21616);
and U21751 (N_21751,N_21727,N_21570);
and U21752 (N_21752,N_21552,N_21587);
xor U21753 (N_21753,N_21688,N_21659);
and U21754 (N_21754,N_21746,N_21588);
or U21755 (N_21755,N_21531,N_21579);
nor U21756 (N_21756,N_21709,N_21742);
xnor U21757 (N_21757,N_21529,N_21654);
nor U21758 (N_21758,N_21622,N_21655);
xnor U21759 (N_21759,N_21607,N_21568);
and U21760 (N_21760,N_21586,N_21601);
and U21761 (N_21761,N_21603,N_21639);
and U21762 (N_21762,N_21533,N_21676);
nor U21763 (N_21763,N_21744,N_21610);
nand U21764 (N_21764,N_21681,N_21702);
xor U21765 (N_21765,N_21695,N_21594);
or U21766 (N_21766,N_21566,N_21582);
nand U21767 (N_21767,N_21577,N_21630);
xnor U21768 (N_21768,N_21706,N_21649);
nor U21769 (N_21769,N_21697,N_21698);
or U21770 (N_21770,N_21503,N_21521);
and U21771 (N_21771,N_21538,N_21737);
xnor U21772 (N_21772,N_21735,N_21627);
nor U21773 (N_21773,N_21572,N_21584);
nor U21774 (N_21774,N_21560,N_21625);
xor U21775 (N_21775,N_21725,N_21501);
nor U21776 (N_21776,N_21683,N_21699);
or U21777 (N_21777,N_21621,N_21575);
or U21778 (N_21778,N_21648,N_21554);
and U21779 (N_21779,N_21544,N_21642);
xnor U21780 (N_21780,N_21679,N_21666);
nor U21781 (N_21781,N_21524,N_21717);
and U21782 (N_21782,N_21653,N_21705);
or U21783 (N_21783,N_21637,N_21580);
xor U21784 (N_21784,N_21530,N_21656);
or U21785 (N_21785,N_21674,N_21661);
or U21786 (N_21786,N_21585,N_21628);
or U21787 (N_21787,N_21743,N_21693);
nor U21788 (N_21788,N_21636,N_21712);
nor U21789 (N_21789,N_21686,N_21605);
or U21790 (N_21790,N_21513,N_21730);
xor U21791 (N_21791,N_21663,N_21564);
and U21792 (N_21792,N_21711,N_21741);
and U21793 (N_21793,N_21546,N_21547);
or U21794 (N_21794,N_21640,N_21714);
nor U21795 (N_21795,N_21549,N_21728);
nor U21796 (N_21796,N_21684,N_21551);
or U21797 (N_21797,N_21632,N_21687);
or U21798 (N_21798,N_21731,N_21729);
and U21799 (N_21799,N_21583,N_21668);
and U21800 (N_21800,N_21534,N_21617);
or U21801 (N_21801,N_21520,N_21680);
nand U21802 (N_21802,N_21608,N_21677);
xor U21803 (N_21803,N_21660,N_21581);
and U21804 (N_21804,N_21669,N_21671);
xnor U21805 (N_21805,N_21623,N_21536);
nand U21806 (N_21806,N_21545,N_21635);
nor U21807 (N_21807,N_21541,N_21614);
or U21808 (N_21808,N_21690,N_21626);
and U21809 (N_21809,N_21716,N_21510);
or U21810 (N_21810,N_21553,N_21733);
xnor U21811 (N_21811,N_21696,N_21539);
and U21812 (N_21812,N_21540,N_21723);
nor U21813 (N_21813,N_21567,N_21664);
nor U21814 (N_21814,N_21682,N_21562);
nor U21815 (N_21815,N_21708,N_21747);
and U21816 (N_21816,N_21740,N_21634);
xor U21817 (N_21817,N_21619,N_21555);
xnor U21818 (N_21818,N_21609,N_21631);
and U21819 (N_21819,N_21550,N_21611);
nor U21820 (N_21820,N_21645,N_21672);
or U21821 (N_21821,N_21739,N_21597);
and U21822 (N_21822,N_21595,N_21719);
and U21823 (N_21823,N_21596,N_21678);
and U21824 (N_21824,N_21647,N_21745);
or U21825 (N_21825,N_21514,N_21720);
and U21826 (N_21826,N_21537,N_21576);
and U21827 (N_21827,N_21673,N_21593);
nor U21828 (N_21828,N_21641,N_21500);
and U21829 (N_21829,N_21559,N_21694);
xor U21830 (N_21830,N_21732,N_21578);
and U21831 (N_21831,N_21624,N_21509);
nand U21832 (N_21832,N_21561,N_21526);
xor U21833 (N_21833,N_21713,N_21511);
xor U21834 (N_21834,N_21504,N_21573);
nand U21835 (N_21835,N_21589,N_21600);
nand U21836 (N_21836,N_21701,N_21689);
and U21837 (N_21837,N_21508,N_21704);
nor U21838 (N_21838,N_21633,N_21722);
nor U21839 (N_21839,N_21571,N_21703);
xor U21840 (N_21840,N_21604,N_21665);
and U21841 (N_21841,N_21506,N_21726);
xnor U21842 (N_21842,N_21592,N_21662);
xnor U21843 (N_21843,N_21721,N_21646);
nor U21844 (N_21844,N_21618,N_21543);
xor U21845 (N_21845,N_21527,N_21724);
nand U21846 (N_21846,N_21715,N_21700);
xor U21847 (N_21847,N_21738,N_21651);
nand U21848 (N_21848,N_21535,N_21749);
xnor U21849 (N_21849,N_21670,N_21563);
xnor U21850 (N_21850,N_21691,N_21602);
or U21851 (N_21851,N_21505,N_21734);
and U21852 (N_21852,N_21548,N_21612);
xor U21853 (N_21853,N_21590,N_21606);
and U21854 (N_21854,N_21569,N_21599);
nand U21855 (N_21855,N_21620,N_21629);
or U21856 (N_21856,N_21644,N_21518);
nand U21857 (N_21857,N_21748,N_21558);
nand U21858 (N_21858,N_21613,N_21525);
nor U21859 (N_21859,N_21615,N_21652);
nand U21860 (N_21860,N_21591,N_21515);
and U21861 (N_21861,N_21685,N_21519);
and U21862 (N_21862,N_21542,N_21523);
nor U21863 (N_21863,N_21692,N_21556);
and U21864 (N_21864,N_21736,N_21517);
nand U21865 (N_21865,N_21718,N_21650);
or U21866 (N_21866,N_21707,N_21528);
nand U21867 (N_21867,N_21532,N_21710);
xnor U21868 (N_21868,N_21565,N_21557);
or U21869 (N_21869,N_21507,N_21638);
and U21870 (N_21870,N_21516,N_21598);
nor U21871 (N_21871,N_21657,N_21574);
or U21872 (N_21872,N_21522,N_21667);
nand U21873 (N_21873,N_21643,N_21675);
and U21874 (N_21874,N_21658,N_21512);
or U21875 (N_21875,N_21574,N_21557);
nand U21876 (N_21876,N_21619,N_21690);
or U21877 (N_21877,N_21723,N_21551);
nand U21878 (N_21878,N_21677,N_21678);
xor U21879 (N_21879,N_21725,N_21535);
nor U21880 (N_21880,N_21522,N_21546);
or U21881 (N_21881,N_21649,N_21574);
or U21882 (N_21882,N_21572,N_21686);
nor U21883 (N_21883,N_21512,N_21598);
nand U21884 (N_21884,N_21578,N_21733);
or U21885 (N_21885,N_21580,N_21525);
and U21886 (N_21886,N_21661,N_21626);
nand U21887 (N_21887,N_21705,N_21566);
xnor U21888 (N_21888,N_21608,N_21538);
nand U21889 (N_21889,N_21509,N_21697);
nor U21890 (N_21890,N_21719,N_21647);
nor U21891 (N_21891,N_21722,N_21502);
nand U21892 (N_21892,N_21717,N_21537);
or U21893 (N_21893,N_21732,N_21665);
and U21894 (N_21894,N_21692,N_21705);
xor U21895 (N_21895,N_21645,N_21514);
nand U21896 (N_21896,N_21683,N_21706);
and U21897 (N_21897,N_21503,N_21746);
and U21898 (N_21898,N_21664,N_21659);
nand U21899 (N_21899,N_21643,N_21647);
or U21900 (N_21900,N_21572,N_21545);
and U21901 (N_21901,N_21559,N_21636);
or U21902 (N_21902,N_21741,N_21621);
or U21903 (N_21903,N_21735,N_21720);
xor U21904 (N_21904,N_21533,N_21553);
and U21905 (N_21905,N_21626,N_21562);
or U21906 (N_21906,N_21736,N_21524);
xnor U21907 (N_21907,N_21714,N_21521);
nor U21908 (N_21908,N_21672,N_21510);
and U21909 (N_21909,N_21546,N_21564);
or U21910 (N_21910,N_21582,N_21664);
or U21911 (N_21911,N_21573,N_21629);
and U21912 (N_21912,N_21679,N_21526);
xnor U21913 (N_21913,N_21567,N_21701);
or U21914 (N_21914,N_21707,N_21578);
nand U21915 (N_21915,N_21616,N_21514);
nand U21916 (N_21916,N_21610,N_21644);
nor U21917 (N_21917,N_21611,N_21609);
or U21918 (N_21918,N_21511,N_21562);
xnor U21919 (N_21919,N_21595,N_21710);
and U21920 (N_21920,N_21744,N_21506);
nor U21921 (N_21921,N_21538,N_21536);
nor U21922 (N_21922,N_21615,N_21630);
xor U21923 (N_21923,N_21551,N_21711);
nand U21924 (N_21924,N_21514,N_21508);
or U21925 (N_21925,N_21719,N_21729);
or U21926 (N_21926,N_21715,N_21530);
nor U21927 (N_21927,N_21614,N_21742);
or U21928 (N_21928,N_21516,N_21543);
or U21929 (N_21929,N_21689,N_21584);
xnor U21930 (N_21930,N_21607,N_21749);
nand U21931 (N_21931,N_21542,N_21681);
or U21932 (N_21932,N_21640,N_21503);
xnor U21933 (N_21933,N_21598,N_21545);
xor U21934 (N_21934,N_21640,N_21616);
nand U21935 (N_21935,N_21529,N_21580);
or U21936 (N_21936,N_21522,N_21543);
nor U21937 (N_21937,N_21638,N_21532);
or U21938 (N_21938,N_21567,N_21570);
nor U21939 (N_21939,N_21641,N_21508);
nand U21940 (N_21940,N_21702,N_21732);
nand U21941 (N_21941,N_21555,N_21510);
xor U21942 (N_21942,N_21725,N_21588);
xor U21943 (N_21943,N_21664,N_21541);
nand U21944 (N_21944,N_21603,N_21727);
nand U21945 (N_21945,N_21502,N_21644);
xnor U21946 (N_21946,N_21708,N_21595);
or U21947 (N_21947,N_21500,N_21510);
nor U21948 (N_21948,N_21599,N_21639);
or U21949 (N_21949,N_21517,N_21580);
xnor U21950 (N_21950,N_21629,N_21540);
and U21951 (N_21951,N_21534,N_21542);
or U21952 (N_21952,N_21660,N_21714);
nand U21953 (N_21953,N_21631,N_21575);
and U21954 (N_21954,N_21668,N_21651);
nor U21955 (N_21955,N_21747,N_21693);
and U21956 (N_21956,N_21589,N_21554);
xor U21957 (N_21957,N_21649,N_21717);
nor U21958 (N_21958,N_21553,N_21528);
nor U21959 (N_21959,N_21732,N_21662);
nor U21960 (N_21960,N_21576,N_21692);
and U21961 (N_21961,N_21680,N_21503);
and U21962 (N_21962,N_21522,N_21624);
and U21963 (N_21963,N_21572,N_21588);
or U21964 (N_21964,N_21709,N_21713);
nor U21965 (N_21965,N_21698,N_21504);
xor U21966 (N_21966,N_21513,N_21636);
and U21967 (N_21967,N_21589,N_21517);
or U21968 (N_21968,N_21654,N_21602);
or U21969 (N_21969,N_21597,N_21689);
and U21970 (N_21970,N_21636,N_21686);
nand U21971 (N_21971,N_21686,N_21642);
and U21972 (N_21972,N_21683,N_21617);
or U21973 (N_21973,N_21690,N_21652);
xor U21974 (N_21974,N_21545,N_21663);
nor U21975 (N_21975,N_21683,N_21506);
and U21976 (N_21976,N_21739,N_21515);
or U21977 (N_21977,N_21675,N_21661);
nor U21978 (N_21978,N_21713,N_21625);
xor U21979 (N_21979,N_21588,N_21616);
nand U21980 (N_21980,N_21582,N_21731);
or U21981 (N_21981,N_21546,N_21599);
nand U21982 (N_21982,N_21684,N_21602);
and U21983 (N_21983,N_21505,N_21743);
nand U21984 (N_21984,N_21680,N_21718);
nor U21985 (N_21985,N_21742,N_21640);
and U21986 (N_21986,N_21637,N_21629);
xor U21987 (N_21987,N_21644,N_21685);
nand U21988 (N_21988,N_21703,N_21560);
or U21989 (N_21989,N_21534,N_21567);
nor U21990 (N_21990,N_21567,N_21738);
nor U21991 (N_21991,N_21661,N_21632);
nand U21992 (N_21992,N_21653,N_21697);
xor U21993 (N_21993,N_21550,N_21653);
nand U21994 (N_21994,N_21749,N_21662);
or U21995 (N_21995,N_21600,N_21531);
and U21996 (N_21996,N_21631,N_21678);
nand U21997 (N_21997,N_21597,N_21729);
xnor U21998 (N_21998,N_21659,N_21626);
nand U21999 (N_21999,N_21723,N_21693);
nand U22000 (N_22000,N_21964,N_21779);
xnor U22001 (N_22001,N_21761,N_21960);
or U22002 (N_22002,N_21888,N_21774);
nand U22003 (N_22003,N_21777,N_21974);
nor U22004 (N_22004,N_21771,N_21948);
nand U22005 (N_22005,N_21917,N_21752);
nand U22006 (N_22006,N_21928,N_21953);
or U22007 (N_22007,N_21983,N_21858);
or U22008 (N_22008,N_21995,N_21821);
nor U22009 (N_22009,N_21932,N_21780);
nor U22010 (N_22010,N_21866,N_21889);
nand U22011 (N_22011,N_21907,N_21944);
nor U22012 (N_22012,N_21908,N_21835);
or U22013 (N_22013,N_21768,N_21934);
and U22014 (N_22014,N_21999,N_21895);
nand U22015 (N_22015,N_21776,N_21825);
nor U22016 (N_22016,N_21970,N_21819);
nand U22017 (N_22017,N_21894,N_21962);
nor U22018 (N_22018,N_21941,N_21765);
xnor U22019 (N_22019,N_21860,N_21820);
nor U22020 (N_22020,N_21946,N_21919);
nand U22021 (N_22021,N_21816,N_21753);
and U22022 (N_22022,N_21906,N_21814);
and U22023 (N_22023,N_21916,N_21885);
xor U22024 (N_22024,N_21950,N_21817);
nor U22025 (N_22025,N_21940,N_21833);
xnor U22026 (N_22026,N_21802,N_21959);
nand U22027 (N_22027,N_21979,N_21797);
and U22028 (N_22028,N_21849,N_21818);
xor U22029 (N_22029,N_21790,N_21968);
nor U22030 (N_22030,N_21961,N_21963);
xor U22031 (N_22031,N_21881,N_21982);
nand U22032 (N_22032,N_21939,N_21873);
nor U22033 (N_22033,N_21750,N_21846);
and U22034 (N_22034,N_21856,N_21764);
and U22035 (N_22035,N_21839,N_21875);
or U22036 (N_22036,N_21954,N_21792);
xor U22037 (N_22037,N_21929,N_21770);
nand U22038 (N_22038,N_21911,N_21924);
and U22039 (N_22039,N_21871,N_21972);
or U22040 (N_22040,N_21813,N_21997);
xor U22041 (N_22041,N_21931,N_21864);
xnor U22042 (N_22042,N_21957,N_21829);
or U22043 (N_22043,N_21943,N_21925);
nor U22044 (N_22044,N_21773,N_21836);
nor U22045 (N_22045,N_21902,N_21874);
nand U22046 (N_22046,N_21901,N_21955);
xnor U22047 (N_22047,N_21843,N_21884);
and U22048 (N_22048,N_21949,N_21868);
nor U22049 (N_22049,N_21857,N_21980);
nand U22050 (N_22050,N_21930,N_21945);
nor U22051 (N_22051,N_21956,N_21832);
xor U22052 (N_22052,N_21996,N_21879);
and U22053 (N_22053,N_21851,N_21897);
and U22054 (N_22054,N_21891,N_21926);
nor U22055 (N_22055,N_21883,N_21806);
xor U22056 (N_22056,N_21967,N_21772);
xnor U22057 (N_22057,N_21903,N_21751);
and U22058 (N_22058,N_21815,N_21905);
and U22059 (N_22059,N_21998,N_21759);
and U22060 (N_22060,N_21852,N_21775);
xnor U22061 (N_22061,N_21870,N_21847);
xor U22062 (N_22062,N_21799,N_21992);
and U22063 (N_22063,N_21990,N_21840);
nand U22064 (N_22064,N_21981,N_21803);
xnor U22065 (N_22065,N_21826,N_21882);
and U22066 (N_22066,N_21854,N_21984);
nor U22067 (N_22067,N_21876,N_21760);
nand U22068 (N_22068,N_21952,N_21975);
and U22069 (N_22069,N_21850,N_21947);
or U22070 (N_22070,N_21805,N_21862);
nor U22071 (N_22071,N_21795,N_21786);
xor U22072 (N_22072,N_21969,N_21844);
and U22073 (N_22073,N_21782,N_21793);
or U22074 (N_22074,N_21785,N_21918);
nand U22075 (N_22075,N_21767,N_21878);
nor U22076 (N_22076,N_21827,N_21892);
nor U22077 (N_22077,N_21778,N_21783);
nand U22078 (N_22078,N_21796,N_21763);
xor U22079 (N_22079,N_21937,N_21807);
nor U22080 (N_22080,N_21828,N_21987);
and U22081 (N_22081,N_21958,N_21804);
nor U22082 (N_22082,N_21993,N_21973);
nand U22083 (N_22083,N_21798,N_21808);
and U22084 (N_22084,N_21867,N_21985);
nand U22085 (N_22085,N_21838,N_21914);
xor U22086 (N_22086,N_21912,N_21830);
nand U22087 (N_22087,N_21855,N_21800);
or U22088 (N_22088,N_21971,N_21794);
and U22089 (N_22089,N_21923,N_21935);
nor U22090 (N_22090,N_21757,N_21801);
or U22091 (N_22091,N_21756,N_21877);
and U22092 (N_22092,N_21824,N_21848);
or U22093 (N_22093,N_21841,N_21754);
and U22094 (N_22094,N_21787,N_21904);
xor U22095 (N_22095,N_21938,N_21890);
or U22096 (N_22096,N_21927,N_21872);
nor U22097 (N_22097,N_21965,N_21976);
nor U22098 (N_22098,N_21766,N_21896);
xnor U22099 (N_22099,N_21812,N_21988);
and U22100 (N_22100,N_21789,N_21791);
xor U22101 (N_22101,N_21863,N_21809);
or U22102 (N_22102,N_21845,N_21922);
and U22103 (N_22103,N_21966,N_21853);
or U22104 (N_22104,N_21788,N_21936);
and U22105 (N_22105,N_21822,N_21977);
nor U22106 (N_22106,N_21758,N_21865);
nor U22107 (N_22107,N_21811,N_21755);
or U22108 (N_22108,N_21869,N_21886);
and U22109 (N_22109,N_21986,N_21769);
nand U22110 (N_22110,N_21910,N_21762);
or U22111 (N_22111,N_21989,N_21810);
nand U22112 (N_22112,N_21861,N_21837);
and U22113 (N_22113,N_21951,N_21915);
and U22114 (N_22114,N_21994,N_21893);
and U22115 (N_22115,N_21898,N_21784);
nor U22116 (N_22116,N_21842,N_21921);
and U22117 (N_22117,N_21978,N_21834);
nand U22118 (N_22118,N_21942,N_21899);
nor U22119 (N_22119,N_21900,N_21991);
and U22120 (N_22120,N_21909,N_21913);
or U22121 (N_22121,N_21920,N_21887);
or U22122 (N_22122,N_21880,N_21823);
or U22123 (N_22123,N_21831,N_21933);
xor U22124 (N_22124,N_21859,N_21781);
and U22125 (N_22125,N_21869,N_21819);
or U22126 (N_22126,N_21874,N_21821);
xnor U22127 (N_22127,N_21815,N_21959);
and U22128 (N_22128,N_21838,N_21878);
or U22129 (N_22129,N_21804,N_21955);
xor U22130 (N_22130,N_21893,N_21937);
nor U22131 (N_22131,N_21848,N_21833);
xnor U22132 (N_22132,N_21916,N_21752);
nand U22133 (N_22133,N_21936,N_21856);
or U22134 (N_22134,N_21886,N_21768);
nor U22135 (N_22135,N_21999,N_21966);
nor U22136 (N_22136,N_21781,N_21782);
nand U22137 (N_22137,N_21921,N_21839);
nand U22138 (N_22138,N_21945,N_21779);
or U22139 (N_22139,N_21919,N_21911);
or U22140 (N_22140,N_21883,N_21820);
nor U22141 (N_22141,N_21916,N_21819);
xor U22142 (N_22142,N_21893,N_21850);
nand U22143 (N_22143,N_21920,N_21966);
and U22144 (N_22144,N_21900,N_21910);
and U22145 (N_22145,N_21836,N_21852);
nand U22146 (N_22146,N_21753,N_21994);
xor U22147 (N_22147,N_21939,N_21842);
nor U22148 (N_22148,N_21915,N_21770);
nor U22149 (N_22149,N_21832,N_21910);
xor U22150 (N_22150,N_21826,N_21803);
nand U22151 (N_22151,N_21964,N_21934);
nand U22152 (N_22152,N_21944,N_21751);
or U22153 (N_22153,N_21994,N_21873);
nand U22154 (N_22154,N_21884,N_21780);
and U22155 (N_22155,N_21807,N_21967);
or U22156 (N_22156,N_21880,N_21756);
or U22157 (N_22157,N_21957,N_21964);
xnor U22158 (N_22158,N_21919,N_21908);
xor U22159 (N_22159,N_21790,N_21781);
nand U22160 (N_22160,N_21964,N_21909);
xor U22161 (N_22161,N_21988,N_21902);
xor U22162 (N_22162,N_21922,N_21901);
or U22163 (N_22163,N_21808,N_21883);
or U22164 (N_22164,N_21950,N_21753);
nand U22165 (N_22165,N_21763,N_21787);
or U22166 (N_22166,N_21756,N_21941);
nor U22167 (N_22167,N_21837,N_21941);
nand U22168 (N_22168,N_21857,N_21793);
nor U22169 (N_22169,N_21818,N_21809);
or U22170 (N_22170,N_21843,N_21833);
xnor U22171 (N_22171,N_21918,N_21889);
nor U22172 (N_22172,N_21979,N_21866);
nor U22173 (N_22173,N_21762,N_21907);
and U22174 (N_22174,N_21931,N_21940);
nor U22175 (N_22175,N_21937,N_21802);
nor U22176 (N_22176,N_21871,N_21944);
or U22177 (N_22177,N_21962,N_21938);
and U22178 (N_22178,N_21848,N_21873);
or U22179 (N_22179,N_21898,N_21884);
or U22180 (N_22180,N_21776,N_21912);
or U22181 (N_22181,N_21941,N_21972);
nor U22182 (N_22182,N_21849,N_21773);
or U22183 (N_22183,N_21831,N_21805);
nand U22184 (N_22184,N_21899,N_21920);
and U22185 (N_22185,N_21815,N_21856);
and U22186 (N_22186,N_21846,N_21979);
or U22187 (N_22187,N_21765,N_21771);
nor U22188 (N_22188,N_21957,N_21904);
nand U22189 (N_22189,N_21874,N_21791);
nand U22190 (N_22190,N_21765,N_21768);
nor U22191 (N_22191,N_21923,N_21857);
xor U22192 (N_22192,N_21930,N_21807);
or U22193 (N_22193,N_21806,N_21753);
and U22194 (N_22194,N_21783,N_21830);
nor U22195 (N_22195,N_21785,N_21750);
nor U22196 (N_22196,N_21885,N_21960);
nor U22197 (N_22197,N_21765,N_21836);
and U22198 (N_22198,N_21823,N_21879);
nand U22199 (N_22199,N_21848,N_21957);
and U22200 (N_22200,N_21914,N_21988);
or U22201 (N_22201,N_21883,N_21865);
or U22202 (N_22202,N_21811,N_21871);
nor U22203 (N_22203,N_21898,N_21984);
nand U22204 (N_22204,N_21984,N_21915);
nor U22205 (N_22205,N_21770,N_21917);
nand U22206 (N_22206,N_21845,N_21882);
nor U22207 (N_22207,N_21818,N_21988);
or U22208 (N_22208,N_21953,N_21897);
nor U22209 (N_22209,N_21841,N_21776);
and U22210 (N_22210,N_21991,N_21770);
or U22211 (N_22211,N_21948,N_21781);
and U22212 (N_22212,N_21791,N_21898);
xnor U22213 (N_22213,N_21958,N_21862);
nand U22214 (N_22214,N_21989,N_21942);
and U22215 (N_22215,N_21877,N_21875);
or U22216 (N_22216,N_21863,N_21993);
or U22217 (N_22217,N_21850,N_21897);
or U22218 (N_22218,N_21881,N_21900);
nor U22219 (N_22219,N_21760,N_21909);
nand U22220 (N_22220,N_21780,N_21907);
xnor U22221 (N_22221,N_21988,N_21800);
nor U22222 (N_22222,N_21875,N_21901);
nand U22223 (N_22223,N_21790,N_21892);
or U22224 (N_22224,N_21842,N_21982);
nor U22225 (N_22225,N_21962,N_21880);
xnor U22226 (N_22226,N_21769,N_21833);
and U22227 (N_22227,N_21867,N_21758);
nand U22228 (N_22228,N_21889,N_21854);
or U22229 (N_22229,N_21793,N_21859);
xor U22230 (N_22230,N_21806,N_21950);
xor U22231 (N_22231,N_21939,N_21972);
xnor U22232 (N_22232,N_21943,N_21777);
and U22233 (N_22233,N_21793,N_21906);
or U22234 (N_22234,N_21853,N_21828);
nor U22235 (N_22235,N_21929,N_21950);
or U22236 (N_22236,N_21979,N_21930);
nor U22237 (N_22237,N_21977,N_21760);
nand U22238 (N_22238,N_21790,N_21872);
nor U22239 (N_22239,N_21762,N_21771);
xnor U22240 (N_22240,N_21761,N_21949);
and U22241 (N_22241,N_21838,N_21756);
or U22242 (N_22242,N_21953,N_21963);
nand U22243 (N_22243,N_21861,N_21996);
nand U22244 (N_22244,N_21899,N_21806);
nor U22245 (N_22245,N_21980,N_21840);
nor U22246 (N_22246,N_21768,N_21792);
nand U22247 (N_22247,N_21773,N_21805);
xor U22248 (N_22248,N_21757,N_21750);
nand U22249 (N_22249,N_21951,N_21868);
nand U22250 (N_22250,N_22043,N_22137);
or U22251 (N_22251,N_22049,N_22177);
xor U22252 (N_22252,N_22216,N_22112);
and U22253 (N_22253,N_22138,N_22057);
nor U22254 (N_22254,N_22183,N_22228);
or U22255 (N_22255,N_22077,N_22052);
or U22256 (N_22256,N_22106,N_22086);
nor U22257 (N_22257,N_22211,N_22224);
and U22258 (N_22258,N_22185,N_22209);
nor U22259 (N_22259,N_22023,N_22125);
nor U22260 (N_22260,N_22160,N_22175);
nor U22261 (N_22261,N_22114,N_22219);
or U22262 (N_22262,N_22107,N_22127);
and U22263 (N_22263,N_22198,N_22234);
nand U22264 (N_22264,N_22191,N_22117);
and U22265 (N_22265,N_22136,N_22172);
nand U22266 (N_22266,N_22018,N_22141);
or U22267 (N_22267,N_22024,N_22012);
or U22268 (N_22268,N_22105,N_22072);
and U22269 (N_22269,N_22226,N_22020);
nand U22270 (N_22270,N_22184,N_22215);
or U22271 (N_22271,N_22048,N_22133);
or U22272 (N_22272,N_22092,N_22235);
and U22273 (N_22273,N_22101,N_22067);
nand U22274 (N_22274,N_22233,N_22025);
xor U22275 (N_22275,N_22139,N_22030);
or U22276 (N_22276,N_22080,N_22021);
nor U22277 (N_22277,N_22028,N_22222);
and U22278 (N_22278,N_22016,N_22123);
or U22279 (N_22279,N_22203,N_22208);
and U22280 (N_22280,N_22008,N_22121);
nor U22281 (N_22281,N_22095,N_22238);
xnor U22282 (N_22282,N_22161,N_22195);
xor U22283 (N_22283,N_22026,N_22201);
or U22284 (N_22284,N_22082,N_22156);
xor U22285 (N_22285,N_22249,N_22190);
or U22286 (N_22286,N_22015,N_22071);
or U22287 (N_22287,N_22243,N_22115);
nor U22288 (N_22288,N_22056,N_22070);
nor U22289 (N_22289,N_22035,N_22239);
and U22290 (N_22290,N_22229,N_22162);
or U22291 (N_22291,N_22083,N_22240);
xnor U22292 (N_22292,N_22084,N_22174);
or U22293 (N_22293,N_22181,N_22019);
nand U22294 (N_22294,N_22093,N_22073);
nor U22295 (N_22295,N_22068,N_22186);
nor U22296 (N_22296,N_22000,N_22140);
xnor U22297 (N_22297,N_22173,N_22055);
nor U22298 (N_22298,N_22041,N_22230);
nand U22299 (N_22299,N_22031,N_22011);
nand U22300 (N_22300,N_22091,N_22065);
nand U22301 (N_22301,N_22124,N_22061);
and U22302 (N_22302,N_22007,N_22126);
nor U22303 (N_22303,N_22128,N_22003);
nor U22304 (N_22304,N_22247,N_22168);
and U22305 (N_22305,N_22188,N_22204);
and U22306 (N_22306,N_22079,N_22058);
nand U22307 (N_22307,N_22152,N_22163);
nor U22308 (N_22308,N_22166,N_22097);
and U22309 (N_22309,N_22075,N_22225);
nor U22310 (N_22310,N_22116,N_22081);
and U22311 (N_22311,N_22148,N_22036);
or U22312 (N_22312,N_22147,N_22194);
or U22313 (N_22313,N_22214,N_22223);
xor U22314 (N_22314,N_22033,N_22189);
nor U22315 (N_22315,N_22078,N_22113);
xor U22316 (N_22316,N_22199,N_22119);
nor U22317 (N_22317,N_22221,N_22046);
nor U22318 (N_22318,N_22010,N_22034);
nand U22319 (N_22319,N_22220,N_22038);
xnor U22320 (N_22320,N_22153,N_22197);
and U22321 (N_22321,N_22088,N_22232);
and U22322 (N_22322,N_22131,N_22245);
nor U22323 (N_22323,N_22060,N_22098);
xnor U22324 (N_22324,N_22085,N_22096);
and U22325 (N_22325,N_22159,N_22146);
nor U22326 (N_22326,N_22029,N_22142);
xnor U22327 (N_22327,N_22066,N_22017);
xor U22328 (N_22328,N_22179,N_22210);
xnor U22329 (N_22329,N_22165,N_22054);
nand U22330 (N_22330,N_22178,N_22242);
nand U22331 (N_22331,N_22145,N_22196);
or U22332 (N_22332,N_22205,N_22231);
nand U22333 (N_22333,N_22089,N_22039);
or U22334 (N_22334,N_22149,N_22212);
and U22335 (N_22335,N_22180,N_22244);
or U22336 (N_22336,N_22013,N_22192);
nor U22337 (N_22337,N_22135,N_22170);
nand U22338 (N_22338,N_22014,N_22155);
and U22339 (N_22339,N_22206,N_22169);
nand U22340 (N_22340,N_22108,N_22171);
nand U22341 (N_22341,N_22246,N_22059);
or U22342 (N_22342,N_22087,N_22120);
and U22343 (N_22343,N_22104,N_22045);
and U22344 (N_22344,N_22090,N_22006);
nor U22345 (N_22345,N_22050,N_22109);
or U22346 (N_22346,N_22009,N_22001);
xor U22347 (N_22347,N_22042,N_22094);
and U22348 (N_22348,N_22047,N_22236);
and U22349 (N_22349,N_22110,N_22074);
nand U22350 (N_22350,N_22241,N_22051);
xor U22351 (N_22351,N_22182,N_22218);
nor U22352 (N_22352,N_22134,N_22217);
nor U22353 (N_22353,N_22111,N_22164);
nand U22354 (N_22354,N_22237,N_22044);
or U22355 (N_22355,N_22002,N_22143);
nand U22356 (N_22356,N_22130,N_22103);
and U22357 (N_22357,N_22032,N_22154);
nor U22358 (N_22358,N_22213,N_22040);
or U22359 (N_22359,N_22202,N_22022);
or U22360 (N_22360,N_22150,N_22167);
xnor U22361 (N_22361,N_22158,N_22100);
and U22362 (N_22362,N_22064,N_22063);
or U22363 (N_22363,N_22248,N_22053);
and U22364 (N_22364,N_22037,N_22193);
xor U22365 (N_22365,N_22187,N_22129);
xnor U22366 (N_22366,N_22062,N_22144);
nor U22367 (N_22367,N_22157,N_22118);
and U22368 (N_22368,N_22122,N_22069);
or U22369 (N_22369,N_22227,N_22176);
or U22370 (N_22370,N_22132,N_22151);
nand U22371 (N_22371,N_22076,N_22005);
or U22372 (N_22372,N_22102,N_22200);
and U22373 (N_22373,N_22004,N_22099);
nand U22374 (N_22374,N_22027,N_22207);
and U22375 (N_22375,N_22062,N_22205);
or U22376 (N_22376,N_22180,N_22229);
or U22377 (N_22377,N_22041,N_22246);
nor U22378 (N_22378,N_22023,N_22152);
xor U22379 (N_22379,N_22074,N_22098);
nand U22380 (N_22380,N_22055,N_22233);
xnor U22381 (N_22381,N_22147,N_22197);
or U22382 (N_22382,N_22046,N_22014);
xor U22383 (N_22383,N_22191,N_22097);
and U22384 (N_22384,N_22141,N_22034);
nand U22385 (N_22385,N_22104,N_22119);
nor U22386 (N_22386,N_22108,N_22198);
nor U22387 (N_22387,N_22212,N_22060);
and U22388 (N_22388,N_22233,N_22209);
xnor U22389 (N_22389,N_22036,N_22177);
or U22390 (N_22390,N_22012,N_22248);
or U22391 (N_22391,N_22211,N_22212);
xnor U22392 (N_22392,N_22162,N_22089);
or U22393 (N_22393,N_22172,N_22022);
xor U22394 (N_22394,N_22233,N_22105);
or U22395 (N_22395,N_22180,N_22045);
and U22396 (N_22396,N_22126,N_22051);
nand U22397 (N_22397,N_22135,N_22044);
or U22398 (N_22398,N_22197,N_22143);
nand U22399 (N_22399,N_22070,N_22132);
xnor U22400 (N_22400,N_22069,N_22116);
or U22401 (N_22401,N_22029,N_22043);
and U22402 (N_22402,N_22234,N_22107);
and U22403 (N_22403,N_22174,N_22243);
nor U22404 (N_22404,N_22066,N_22184);
nand U22405 (N_22405,N_22014,N_22099);
and U22406 (N_22406,N_22104,N_22207);
and U22407 (N_22407,N_22143,N_22125);
nand U22408 (N_22408,N_22161,N_22017);
nand U22409 (N_22409,N_22001,N_22170);
nand U22410 (N_22410,N_22207,N_22218);
nor U22411 (N_22411,N_22009,N_22170);
or U22412 (N_22412,N_22189,N_22072);
xor U22413 (N_22413,N_22006,N_22139);
and U22414 (N_22414,N_22240,N_22219);
and U22415 (N_22415,N_22247,N_22074);
nand U22416 (N_22416,N_22015,N_22216);
and U22417 (N_22417,N_22113,N_22195);
nand U22418 (N_22418,N_22103,N_22092);
xor U22419 (N_22419,N_22081,N_22240);
nand U22420 (N_22420,N_22020,N_22179);
and U22421 (N_22421,N_22207,N_22145);
and U22422 (N_22422,N_22190,N_22038);
xor U22423 (N_22423,N_22101,N_22152);
nor U22424 (N_22424,N_22223,N_22091);
xor U22425 (N_22425,N_22054,N_22022);
nand U22426 (N_22426,N_22057,N_22246);
xnor U22427 (N_22427,N_22005,N_22190);
nand U22428 (N_22428,N_22059,N_22148);
nor U22429 (N_22429,N_22175,N_22068);
nand U22430 (N_22430,N_22223,N_22067);
or U22431 (N_22431,N_22159,N_22076);
and U22432 (N_22432,N_22195,N_22235);
xnor U22433 (N_22433,N_22110,N_22169);
nand U22434 (N_22434,N_22133,N_22116);
xnor U22435 (N_22435,N_22133,N_22054);
or U22436 (N_22436,N_22199,N_22197);
nor U22437 (N_22437,N_22160,N_22041);
or U22438 (N_22438,N_22030,N_22067);
and U22439 (N_22439,N_22127,N_22068);
and U22440 (N_22440,N_22110,N_22234);
and U22441 (N_22441,N_22220,N_22019);
and U22442 (N_22442,N_22224,N_22235);
xnor U22443 (N_22443,N_22060,N_22153);
nor U22444 (N_22444,N_22014,N_22181);
nor U22445 (N_22445,N_22055,N_22077);
xnor U22446 (N_22446,N_22179,N_22123);
or U22447 (N_22447,N_22062,N_22204);
nand U22448 (N_22448,N_22145,N_22052);
nand U22449 (N_22449,N_22044,N_22178);
nor U22450 (N_22450,N_22133,N_22199);
or U22451 (N_22451,N_22205,N_22109);
xor U22452 (N_22452,N_22136,N_22190);
nand U22453 (N_22453,N_22013,N_22057);
xor U22454 (N_22454,N_22205,N_22203);
xnor U22455 (N_22455,N_22169,N_22247);
and U22456 (N_22456,N_22153,N_22140);
and U22457 (N_22457,N_22098,N_22247);
nor U22458 (N_22458,N_22209,N_22205);
nor U22459 (N_22459,N_22022,N_22223);
nor U22460 (N_22460,N_22174,N_22176);
nor U22461 (N_22461,N_22017,N_22192);
xnor U22462 (N_22462,N_22181,N_22165);
xor U22463 (N_22463,N_22091,N_22176);
nor U22464 (N_22464,N_22178,N_22241);
or U22465 (N_22465,N_22139,N_22004);
and U22466 (N_22466,N_22105,N_22060);
nand U22467 (N_22467,N_22008,N_22130);
and U22468 (N_22468,N_22049,N_22043);
xor U22469 (N_22469,N_22175,N_22199);
nor U22470 (N_22470,N_22169,N_22012);
nand U22471 (N_22471,N_22213,N_22017);
or U22472 (N_22472,N_22148,N_22241);
xnor U22473 (N_22473,N_22041,N_22240);
and U22474 (N_22474,N_22191,N_22177);
nand U22475 (N_22475,N_22015,N_22021);
nand U22476 (N_22476,N_22102,N_22105);
and U22477 (N_22477,N_22172,N_22101);
and U22478 (N_22478,N_22109,N_22206);
xor U22479 (N_22479,N_22123,N_22189);
and U22480 (N_22480,N_22139,N_22196);
and U22481 (N_22481,N_22070,N_22025);
nor U22482 (N_22482,N_22029,N_22210);
xnor U22483 (N_22483,N_22066,N_22210);
or U22484 (N_22484,N_22039,N_22225);
xnor U22485 (N_22485,N_22168,N_22055);
or U22486 (N_22486,N_22170,N_22033);
xor U22487 (N_22487,N_22195,N_22224);
and U22488 (N_22488,N_22059,N_22222);
and U22489 (N_22489,N_22082,N_22153);
nand U22490 (N_22490,N_22022,N_22038);
and U22491 (N_22491,N_22037,N_22013);
or U22492 (N_22492,N_22181,N_22053);
xor U22493 (N_22493,N_22152,N_22133);
xor U22494 (N_22494,N_22060,N_22185);
xor U22495 (N_22495,N_22108,N_22189);
and U22496 (N_22496,N_22181,N_22186);
and U22497 (N_22497,N_22079,N_22119);
nand U22498 (N_22498,N_22085,N_22242);
nand U22499 (N_22499,N_22192,N_22113);
and U22500 (N_22500,N_22269,N_22305);
nor U22501 (N_22501,N_22471,N_22302);
xor U22502 (N_22502,N_22392,N_22328);
nor U22503 (N_22503,N_22426,N_22339);
and U22504 (N_22504,N_22356,N_22289);
nor U22505 (N_22505,N_22263,N_22495);
nand U22506 (N_22506,N_22274,N_22474);
nand U22507 (N_22507,N_22341,N_22286);
nand U22508 (N_22508,N_22414,N_22368);
nor U22509 (N_22509,N_22303,N_22325);
or U22510 (N_22510,N_22281,N_22454);
nand U22511 (N_22511,N_22373,N_22321);
nand U22512 (N_22512,N_22367,N_22313);
nand U22513 (N_22513,N_22369,N_22372);
nand U22514 (N_22514,N_22479,N_22461);
xnor U22515 (N_22515,N_22482,N_22485);
xor U22516 (N_22516,N_22265,N_22428);
nand U22517 (N_22517,N_22353,N_22312);
nor U22518 (N_22518,N_22273,N_22472);
xor U22519 (N_22519,N_22278,N_22293);
and U22520 (N_22520,N_22361,N_22359);
nor U22521 (N_22521,N_22282,N_22387);
nor U22522 (N_22522,N_22491,N_22345);
nor U22523 (N_22523,N_22316,N_22434);
nand U22524 (N_22524,N_22447,N_22453);
and U22525 (N_22525,N_22407,N_22425);
or U22526 (N_22526,N_22393,N_22486);
xnor U22527 (N_22527,N_22354,N_22351);
nor U22528 (N_22528,N_22431,N_22450);
xor U22529 (N_22529,N_22259,N_22371);
nor U22530 (N_22530,N_22498,N_22430);
nor U22531 (N_22531,N_22399,N_22390);
nor U22532 (N_22532,N_22350,N_22412);
and U22533 (N_22533,N_22264,N_22365);
nor U22534 (N_22534,N_22421,N_22406);
and U22535 (N_22535,N_22441,N_22487);
nand U22536 (N_22536,N_22277,N_22255);
xor U22537 (N_22537,N_22420,N_22287);
nand U22538 (N_22538,N_22308,N_22307);
nor U22539 (N_22539,N_22352,N_22291);
or U22540 (N_22540,N_22301,N_22309);
nand U22541 (N_22541,N_22357,N_22314);
or U22542 (N_22542,N_22283,N_22256);
or U22543 (N_22543,N_22298,N_22419);
and U22544 (N_22544,N_22438,N_22452);
nand U22545 (N_22545,N_22375,N_22388);
or U22546 (N_22546,N_22409,N_22318);
nor U22547 (N_22547,N_22451,N_22266);
nor U22548 (N_22548,N_22327,N_22370);
nand U22549 (N_22549,N_22460,N_22284);
and U22550 (N_22550,N_22443,N_22310);
and U22551 (N_22551,N_22459,N_22422);
nor U22552 (N_22552,N_22366,N_22427);
or U22553 (N_22553,N_22257,N_22488);
nand U22554 (N_22554,N_22376,N_22338);
nand U22555 (N_22555,N_22383,N_22483);
nor U22556 (N_22556,N_22386,N_22444);
or U22557 (N_22557,N_22466,N_22411);
or U22558 (N_22558,N_22496,N_22396);
nor U22559 (N_22559,N_22465,N_22299);
xor U22560 (N_22560,N_22268,N_22464);
nor U22561 (N_22561,N_22455,N_22404);
and U22562 (N_22562,N_22276,N_22279);
xor U22563 (N_22563,N_22480,N_22457);
xor U22564 (N_22564,N_22362,N_22349);
or U22565 (N_22565,N_22262,N_22330);
nor U22566 (N_22566,N_22253,N_22448);
or U22567 (N_22567,N_22382,N_22467);
or U22568 (N_22568,N_22272,N_22499);
and U22569 (N_22569,N_22463,N_22381);
and U22570 (N_22570,N_22324,N_22334);
xnor U22571 (N_22571,N_22343,N_22418);
nand U22572 (N_22572,N_22384,N_22473);
nor U22573 (N_22573,N_22340,N_22477);
nor U22574 (N_22574,N_22481,N_22379);
xor U22575 (N_22575,N_22360,N_22333);
or U22576 (N_22576,N_22319,N_22267);
or U22577 (N_22577,N_22413,N_22304);
nand U22578 (N_22578,N_22374,N_22335);
xor U22579 (N_22579,N_22292,N_22449);
xnor U22580 (N_22580,N_22497,N_22423);
nand U22581 (N_22581,N_22462,N_22342);
and U22582 (N_22582,N_22363,N_22400);
or U22583 (N_22583,N_22469,N_22440);
xor U22584 (N_22584,N_22252,N_22271);
xnor U22585 (N_22585,N_22493,N_22322);
nand U22586 (N_22586,N_22300,N_22401);
and U22587 (N_22587,N_22378,N_22346);
or U22588 (N_22588,N_22397,N_22410);
nor U22589 (N_22589,N_22288,N_22320);
or U22590 (N_22590,N_22389,N_22439);
or U22591 (N_22591,N_22332,N_22317);
nor U22592 (N_22592,N_22385,N_22476);
xnor U22593 (N_22593,N_22394,N_22331);
xor U22594 (N_22594,N_22403,N_22395);
nand U22595 (N_22595,N_22250,N_22280);
xor U22596 (N_22596,N_22417,N_22458);
or U22597 (N_22597,N_22416,N_22408);
nand U22598 (N_22598,N_22391,N_22475);
xnor U22599 (N_22599,N_22377,N_22294);
xnor U22600 (N_22600,N_22275,N_22297);
nor U22601 (N_22601,N_22442,N_22261);
and U22602 (N_22602,N_22270,N_22435);
nand U22603 (N_22603,N_22344,N_22337);
nand U22604 (N_22604,N_22402,N_22437);
xnor U22605 (N_22605,N_22424,N_22311);
nor U22606 (N_22606,N_22484,N_22296);
or U22607 (N_22607,N_22348,N_22290);
or U22608 (N_22608,N_22478,N_22260);
xor U22609 (N_22609,N_22433,N_22315);
nor U22610 (N_22610,N_22405,N_22445);
nor U22611 (N_22611,N_22285,N_22494);
xnor U22612 (N_22612,N_22326,N_22306);
and U22613 (N_22613,N_22489,N_22398);
and U22614 (N_22614,N_22347,N_22446);
and U22615 (N_22615,N_22468,N_22355);
xnor U22616 (N_22616,N_22251,N_22295);
xnor U22617 (N_22617,N_22323,N_22436);
xnor U22618 (N_22618,N_22329,N_22364);
nand U22619 (N_22619,N_22490,N_22358);
xnor U22620 (N_22620,N_22258,N_22415);
nor U22621 (N_22621,N_22336,N_22470);
and U22622 (N_22622,N_22380,N_22254);
xnor U22623 (N_22623,N_22429,N_22432);
or U22624 (N_22624,N_22456,N_22492);
and U22625 (N_22625,N_22480,N_22359);
xor U22626 (N_22626,N_22371,N_22435);
or U22627 (N_22627,N_22265,N_22404);
nor U22628 (N_22628,N_22495,N_22253);
nor U22629 (N_22629,N_22383,N_22272);
nor U22630 (N_22630,N_22292,N_22404);
and U22631 (N_22631,N_22449,N_22331);
and U22632 (N_22632,N_22453,N_22496);
or U22633 (N_22633,N_22402,N_22318);
and U22634 (N_22634,N_22450,N_22270);
and U22635 (N_22635,N_22476,N_22463);
nand U22636 (N_22636,N_22351,N_22444);
nand U22637 (N_22637,N_22302,N_22300);
and U22638 (N_22638,N_22366,N_22287);
xnor U22639 (N_22639,N_22359,N_22454);
nor U22640 (N_22640,N_22446,N_22318);
nor U22641 (N_22641,N_22378,N_22416);
or U22642 (N_22642,N_22413,N_22403);
xnor U22643 (N_22643,N_22440,N_22274);
or U22644 (N_22644,N_22358,N_22478);
nand U22645 (N_22645,N_22390,N_22466);
nand U22646 (N_22646,N_22493,N_22343);
or U22647 (N_22647,N_22448,N_22484);
nand U22648 (N_22648,N_22254,N_22420);
nand U22649 (N_22649,N_22316,N_22326);
xnor U22650 (N_22650,N_22256,N_22378);
nor U22651 (N_22651,N_22317,N_22365);
and U22652 (N_22652,N_22410,N_22275);
nand U22653 (N_22653,N_22396,N_22408);
nand U22654 (N_22654,N_22434,N_22477);
and U22655 (N_22655,N_22306,N_22443);
or U22656 (N_22656,N_22496,N_22428);
nor U22657 (N_22657,N_22262,N_22353);
xor U22658 (N_22658,N_22330,N_22465);
xor U22659 (N_22659,N_22451,N_22311);
or U22660 (N_22660,N_22336,N_22258);
nand U22661 (N_22661,N_22488,N_22479);
and U22662 (N_22662,N_22360,N_22378);
nor U22663 (N_22663,N_22350,N_22470);
xnor U22664 (N_22664,N_22281,N_22282);
or U22665 (N_22665,N_22307,N_22489);
nor U22666 (N_22666,N_22393,N_22446);
xnor U22667 (N_22667,N_22473,N_22478);
nand U22668 (N_22668,N_22349,N_22458);
or U22669 (N_22669,N_22307,N_22374);
nand U22670 (N_22670,N_22401,N_22477);
and U22671 (N_22671,N_22287,N_22372);
or U22672 (N_22672,N_22398,N_22459);
and U22673 (N_22673,N_22292,N_22267);
xor U22674 (N_22674,N_22263,N_22283);
xor U22675 (N_22675,N_22275,N_22298);
xnor U22676 (N_22676,N_22296,N_22482);
xor U22677 (N_22677,N_22380,N_22483);
xor U22678 (N_22678,N_22252,N_22430);
or U22679 (N_22679,N_22386,N_22333);
nand U22680 (N_22680,N_22344,N_22487);
xnor U22681 (N_22681,N_22468,N_22426);
xnor U22682 (N_22682,N_22369,N_22360);
nand U22683 (N_22683,N_22376,N_22343);
and U22684 (N_22684,N_22443,N_22455);
nor U22685 (N_22685,N_22320,N_22279);
or U22686 (N_22686,N_22453,N_22332);
xor U22687 (N_22687,N_22452,N_22349);
and U22688 (N_22688,N_22311,N_22325);
nor U22689 (N_22689,N_22257,N_22424);
nor U22690 (N_22690,N_22481,N_22392);
xnor U22691 (N_22691,N_22424,N_22326);
or U22692 (N_22692,N_22371,N_22457);
or U22693 (N_22693,N_22361,N_22254);
xnor U22694 (N_22694,N_22319,N_22276);
nand U22695 (N_22695,N_22327,N_22448);
nand U22696 (N_22696,N_22444,N_22317);
nor U22697 (N_22697,N_22415,N_22400);
or U22698 (N_22698,N_22414,N_22376);
nor U22699 (N_22699,N_22316,N_22308);
or U22700 (N_22700,N_22471,N_22309);
or U22701 (N_22701,N_22403,N_22409);
nand U22702 (N_22702,N_22462,N_22335);
nor U22703 (N_22703,N_22419,N_22378);
or U22704 (N_22704,N_22346,N_22342);
nand U22705 (N_22705,N_22381,N_22333);
xor U22706 (N_22706,N_22271,N_22317);
xnor U22707 (N_22707,N_22312,N_22288);
nor U22708 (N_22708,N_22414,N_22327);
nand U22709 (N_22709,N_22497,N_22293);
and U22710 (N_22710,N_22361,N_22471);
and U22711 (N_22711,N_22450,N_22487);
xor U22712 (N_22712,N_22345,N_22260);
nand U22713 (N_22713,N_22253,N_22376);
or U22714 (N_22714,N_22407,N_22270);
nand U22715 (N_22715,N_22489,N_22362);
and U22716 (N_22716,N_22385,N_22353);
or U22717 (N_22717,N_22492,N_22281);
and U22718 (N_22718,N_22325,N_22430);
and U22719 (N_22719,N_22342,N_22357);
and U22720 (N_22720,N_22285,N_22490);
and U22721 (N_22721,N_22295,N_22481);
and U22722 (N_22722,N_22396,N_22403);
and U22723 (N_22723,N_22473,N_22466);
nor U22724 (N_22724,N_22438,N_22281);
nand U22725 (N_22725,N_22319,N_22415);
or U22726 (N_22726,N_22358,N_22305);
nor U22727 (N_22727,N_22328,N_22298);
or U22728 (N_22728,N_22479,N_22295);
xnor U22729 (N_22729,N_22342,N_22395);
xnor U22730 (N_22730,N_22277,N_22413);
or U22731 (N_22731,N_22444,N_22435);
or U22732 (N_22732,N_22391,N_22471);
and U22733 (N_22733,N_22456,N_22403);
and U22734 (N_22734,N_22399,N_22491);
xor U22735 (N_22735,N_22328,N_22252);
and U22736 (N_22736,N_22257,N_22382);
or U22737 (N_22737,N_22493,N_22258);
and U22738 (N_22738,N_22477,N_22369);
nor U22739 (N_22739,N_22445,N_22434);
nand U22740 (N_22740,N_22371,N_22362);
nand U22741 (N_22741,N_22486,N_22473);
nor U22742 (N_22742,N_22395,N_22289);
xor U22743 (N_22743,N_22300,N_22256);
nor U22744 (N_22744,N_22330,N_22449);
and U22745 (N_22745,N_22273,N_22492);
or U22746 (N_22746,N_22310,N_22326);
nor U22747 (N_22747,N_22255,N_22363);
nor U22748 (N_22748,N_22416,N_22288);
and U22749 (N_22749,N_22453,N_22484);
and U22750 (N_22750,N_22718,N_22599);
nand U22751 (N_22751,N_22564,N_22666);
and U22752 (N_22752,N_22701,N_22542);
nor U22753 (N_22753,N_22672,N_22622);
xnor U22754 (N_22754,N_22545,N_22706);
or U22755 (N_22755,N_22661,N_22653);
nor U22756 (N_22756,N_22699,N_22620);
xor U22757 (N_22757,N_22698,N_22595);
nor U22758 (N_22758,N_22736,N_22514);
and U22759 (N_22759,N_22727,N_22517);
and U22760 (N_22760,N_22726,N_22566);
nor U22761 (N_22761,N_22535,N_22586);
and U22762 (N_22762,N_22747,N_22612);
or U22763 (N_22763,N_22683,N_22597);
or U22764 (N_22764,N_22518,N_22516);
and U22765 (N_22765,N_22697,N_22615);
xor U22766 (N_22766,N_22580,N_22745);
and U22767 (N_22767,N_22630,N_22607);
nor U22768 (N_22768,N_22515,N_22700);
nor U22769 (N_22769,N_22705,N_22558);
and U22770 (N_22770,N_22505,N_22647);
xnor U22771 (N_22771,N_22560,N_22714);
and U22772 (N_22772,N_22569,N_22660);
nand U22773 (N_22773,N_22601,N_22685);
and U22774 (N_22774,N_22712,N_22682);
or U22775 (N_22775,N_22675,N_22592);
nor U22776 (N_22776,N_22567,N_22507);
or U22777 (N_22777,N_22674,N_22688);
nor U22778 (N_22778,N_22539,N_22663);
and U22779 (N_22779,N_22528,N_22687);
xnor U22780 (N_22780,N_22561,N_22578);
xor U22781 (N_22781,N_22526,N_22725);
or U22782 (N_22782,N_22636,N_22704);
or U22783 (N_22783,N_22676,N_22737);
nor U22784 (N_22784,N_22593,N_22533);
xnor U22785 (N_22785,N_22664,N_22695);
nand U22786 (N_22786,N_22531,N_22551);
nor U22787 (N_22787,N_22740,N_22713);
and U22788 (N_22788,N_22632,N_22555);
xnor U22789 (N_22789,N_22694,N_22568);
and U22790 (N_22790,N_22502,N_22691);
and U22791 (N_22791,N_22588,N_22540);
and U22792 (N_22792,N_22696,N_22521);
and U22793 (N_22793,N_22719,N_22731);
or U22794 (N_22794,N_22667,N_22641);
nor U22795 (N_22795,N_22741,N_22656);
xor U22796 (N_22796,N_22638,N_22673);
nand U22797 (N_22797,N_22626,N_22614);
nor U22798 (N_22798,N_22609,N_22639);
nor U22799 (N_22799,N_22742,N_22534);
xnor U22800 (N_22800,N_22541,N_22654);
xnor U22801 (N_22801,N_22648,N_22583);
or U22802 (N_22802,N_22585,N_22681);
nand U22803 (N_22803,N_22732,N_22651);
or U22804 (N_22804,N_22523,N_22710);
xor U22805 (N_22805,N_22657,N_22512);
and U22806 (N_22806,N_22670,N_22572);
or U22807 (N_22807,N_22532,N_22543);
nand U22808 (N_22808,N_22680,N_22716);
and U22809 (N_22809,N_22658,N_22734);
xnor U22810 (N_22810,N_22621,N_22721);
nand U22811 (N_22811,N_22552,N_22684);
xnor U22812 (N_22812,N_22735,N_22616);
nand U22813 (N_22813,N_22686,N_22678);
xnor U22814 (N_22814,N_22503,N_22631);
xor U22815 (N_22815,N_22645,N_22584);
and U22816 (N_22816,N_22562,N_22605);
xor U22817 (N_22817,N_22511,N_22510);
nand U22818 (N_22818,N_22744,N_22557);
xnor U22819 (N_22819,N_22722,N_22627);
or U22820 (N_22820,N_22619,N_22633);
or U22821 (N_22821,N_22548,N_22635);
xor U22822 (N_22822,N_22743,N_22573);
nand U22823 (N_22823,N_22519,N_22628);
nor U22824 (N_22824,N_22554,N_22500);
or U22825 (N_22825,N_22708,N_22668);
and U22826 (N_22826,N_22662,N_22623);
nor U22827 (N_22827,N_22563,N_22629);
or U22828 (N_22828,N_22677,N_22506);
xor U22829 (N_22829,N_22618,N_22637);
nand U22830 (N_22830,N_22652,N_22729);
and U22831 (N_22831,N_22610,N_22574);
nor U22832 (N_22832,N_22600,N_22581);
nor U22833 (N_22833,N_22707,N_22702);
or U22834 (N_22834,N_22692,N_22749);
xor U22835 (N_22835,N_22748,N_22738);
or U22836 (N_22836,N_22739,N_22709);
xor U22837 (N_22837,N_22570,N_22634);
and U22838 (N_22838,N_22642,N_22650);
and U22839 (N_22839,N_22659,N_22591);
xnor U22840 (N_22840,N_22550,N_22596);
nand U22841 (N_22841,N_22504,N_22723);
nand U22842 (N_22842,N_22524,N_22576);
xor U22843 (N_22843,N_22693,N_22538);
or U22844 (N_22844,N_22703,N_22669);
nor U22845 (N_22845,N_22640,N_22547);
or U22846 (N_22846,N_22603,N_22655);
and U22847 (N_22847,N_22544,N_22529);
nor U22848 (N_22848,N_22644,N_22689);
and U22849 (N_22849,N_22608,N_22587);
or U22850 (N_22850,N_22513,N_22690);
xnor U22851 (N_22851,N_22598,N_22646);
nand U22852 (N_22852,N_22537,N_22522);
and U22853 (N_22853,N_22575,N_22679);
and U22854 (N_22854,N_22509,N_22602);
and U22855 (N_22855,N_22613,N_22746);
nor U22856 (N_22856,N_22671,N_22546);
and U22857 (N_22857,N_22617,N_22525);
nand U22858 (N_22858,N_22549,N_22643);
and U22859 (N_22859,N_22530,N_22611);
nand U22860 (N_22860,N_22606,N_22536);
nor U22861 (N_22861,N_22604,N_22565);
or U22862 (N_22862,N_22582,N_22571);
or U22863 (N_22863,N_22556,N_22553);
or U22864 (N_22864,N_22579,N_22577);
nand U22865 (N_22865,N_22589,N_22733);
xor U22866 (N_22866,N_22625,N_22559);
or U22867 (N_22867,N_22715,N_22665);
or U22868 (N_22868,N_22730,N_22728);
nor U22869 (N_22869,N_22590,N_22649);
nand U22870 (N_22870,N_22508,N_22527);
and U22871 (N_22871,N_22720,N_22520);
and U22872 (N_22872,N_22624,N_22501);
nand U22873 (N_22873,N_22717,N_22724);
or U22874 (N_22874,N_22711,N_22594);
or U22875 (N_22875,N_22652,N_22564);
and U22876 (N_22876,N_22682,N_22710);
and U22877 (N_22877,N_22604,N_22648);
or U22878 (N_22878,N_22640,N_22674);
nor U22879 (N_22879,N_22574,N_22587);
nand U22880 (N_22880,N_22656,N_22677);
nand U22881 (N_22881,N_22564,N_22571);
nand U22882 (N_22882,N_22689,N_22548);
xor U22883 (N_22883,N_22723,N_22663);
and U22884 (N_22884,N_22582,N_22512);
or U22885 (N_22885,N_22562,N_22569);
nor U22886 (N_22886,N_22722,N_22660);
xnor U22887 (N_22887,N_22744,N_22578);
nand U22888 (N_22888,N_22626,N_22526);
nor U22889 (N_22889,N_22662,N_22710);
nor U22890 (N_22890,N_22538,N_22739);
and U22891 (N_22891,N_22534,N_22628);
nand U22892 (N_22892,N_22615,N_22539);
or U22893 (N_22893,N_22576,N_22697);
or U22894 (N_22894,N_22609,N_22592);
xor U22895 (N_22895,N_22715,N_22660);
or U22896 (N_22896,N_22706,N_22654);
and U22897 (N_22897,N_22619,N_22535);
nand U22898 (N_22898,N_22690,N_22571);
nor U22899 (N_22899,N_22746,N_22740);
xnor U22900 (N_22900,N_22580,N_22571);
nand U22901 (N_22901,N_22745,N_22626);
and U22902 (N_22902,N_22542,N_22632);
or U22903 (N_22903,N_22703,N_22586);
or U22904 (N_22904,N_22609,N_22684);
or U22905 (N_22905,N_22547,N_22615);
nor U22906 (N_22906,N_22685,N_22669);
nand U22907 (N_22907,N_22715,N_22698);
and U22908 (N_22908,N_22503,N_22668);
and U22909 (N_22909,N_22624,N_22634);
nand U22910 (N_22910,N_22600,N_22708);
and U22911 (N_22911,N_22507,N_22506);
and U22912 (N_22912,N_22507,N_22731);
nor U22913 (N_22913,N_22697,N_22695);
and U22914 (N_22914,N_22628,N_22539);
and U22915 (N_22915,N_22586,N_22711);
nor U22916 (N_22916,N_22666,N_22743);
nor U22917 (N_22917,N_22663,N_22688);
and U22918 (N_22918,N_22531,N_22687);
nor U22919 (N_22919,N_22747,N_22631);
nand U22920 (N_22920,N_22619,N_22567);
nand U22921 (N_22921,N_22541,N_22731);
and U22922 (N_22922,N_22507,N_22685);
nor U22923 (N_22923,N_22694,N_22527);
xnor U22924 (N_22924,N_22724,N_22559);
or U22925 (N_22925,N_22706,N_22619);
or U22926 (N_22926,N_22582,N_22577);
xor U22927 (N_22927,N_22527,N_22725);
or U22928 (N_22928,N_22748,N_22661);
and U22929 (N_22929,N_22674,N_22661);
and U22930 (N_22930,N_22624,N_22716);
or U22931 (N_22931,N_22631,N_22748);
nand U22932 (N_22932,N_22556,N_22520);
nor U22933 (N_22933,N_22692,N_22570);
and U22934 (N_22934,N_22607,N_22565);
and U22935 (N_22935,N_22574,N_22509);
or U22936 (N_22936,N_22667,N_22546);
xnor U22937 (N_22937,N_22738,N_22679);
nand U22938 (N_22938,N_22734,N_22547);
xnor U22939 (N_22939,N_22729,N_22711);
nand U22940 (N_22940,N_22724,N_22694);
or U22941 (N_22941,N_22522,N_22730);
and U22942 (N_22942,N_22703,N_22568);
nor U22943 (N_22943,N_22532,N_22743);
xnor U22944 (N_22944,N_22654,N_22513);
nand U22945 (N_22945,N_22621,N_22554);
and U22946 (N_22946,N_22524,N_22639);
nand U22947 (N_22947,N_22558,N_22550);
nand U22948 (N_22948,N_22669,N_22661);
nand U22949 (N_22949,N_22715,N_22580);
and U22950 (N_22950,N_22680,N_22551);
or U22951 (N_22951,N_22741,N_22541);
and U22952 (N_22952,N_22517,N_22742);
nor U22953 (N_22953,N_22619,N_22638);
nand U22954 (N_22954,N_22730,N_22532);
xor U22955 (N_22955,N_22581,N_22503);
or U22956 (N_22956,N_22664,N_22744);
and U22957 (N_22957,N_22671,N_22702);
nor U22958 (N_22958,N_22557,N_22715);
and U22959 (N_22959,N_22620,N_22569);
nor U22960 (N_22960,N_22719,N_22517);
xnor U22961 (N_22961,N_22625,N_22572);
xnor U22962 (N_22962,N_22658,N_22633);
nand U22963 (N_22963,N_22586,N_22579);
or U22964 (N_22964,N_22515,N_22546);
xor U22965 (N_22965,N_22558,N_22627);
or U22966 (N_22966,N_22714,N_22723);
and U22967 (N_22967,N_22624,N_22519);
nand U22968 (N_22968,N_22661,N_22613);
nor U22969 (N_22969,N_22682,N_22749);
xor U22970 (N_22970,N_22746,N_22602);
nand U22971 (N_22971,N_22539,N_22664);
or U22972 (N_22972,N_22598,N_22706);
nor U22973 (N_22973,N_22638,N_22692);
xor U22974 (N_22974,N_22593,N_22554);
xor U22975 (N_22975,N_22645,N_22712);
nand U22976 (N_22976,N_22592,N_22670);
nand U22977 (N_22977,N_22509,N_22713);
nand U22978 (N_22978,N_22734,N_22674);
or U22979 (N_22979,N_22508,N_22576);
and U22980 (N_22980,N_22660,N_22662);
xor U22981 (N_22981,N_22672,N_22649);
and U22982 (N_22982,N_22678,N_22698);
and U22983 (N_22983,N_22564,N_22552);
and U22984 (N_22984,N_22520,N_22739);
or U22985 (N_22985,N_22686,N_22553);
nand U22986 (N_22986,N_22511,N_22591);
xnor U22987 (N_22987,N_22693,N_22601);
or U22988 (N_22988,N_22635,N_22714);
nand U22989 (N_22989,N_22712,N_22626);
xnor U22990 (N_22990,N_22719,N_22590);
xnor U22991 (N_22991,N_22736,N_22619);
nor U22992 (N_22992,N_22534,N_22510);
nand U22993 (N_22993,N_22693,N_22612);
nor U22994 (N_22994,N_22634,N_22639);
and U22995 (N_22995,N_22506,N_22619);
nand U22996 (N_22996,N_22524,N_22635);
nand U22997 (N_22997,N_22594,N_22593);
or U22998 (N_22998,N_22599,N_22636);
or U22999 (N_22999,N_22574,N_22531);
nor U23000 (N_23000,N_22864,N_22922);
xnor U23001 (N_23001,N_22945,N_22860);
xor U23002 (N_23002,N_22784,N_22828);
nor U23003 (N_23003,N_22752,N_22939);
nand U23004 (N_23004,N_22954,N_22770);
and U23005 (N_23005,N_22978,N_22889);
nor U23006 (N_23006,N_22785,N_22903);
and U23007 (N_23007,N_22776,N_22862);
and U23008 (N_23008,N_22799,N_22859);
or U23009 (N_23009,N_22975,N_22805);
xor U23010 (N_23010,N_22790,N_22817);
xor U23011 (N_23011,N_22820,N_22809);
nand U23012 (N_23012,N_22991,N_22901);
and U23013 (N_23013,N_22824,N_22750);
xor U23014 (N_23014,N_22965,N_22890);
and U23015 (N_23015,N_22916,N_22923);
nand U23016 (N_23016,N_22947,N_22793);
nand U23017 (N_23017,N_22842,N_22830);
nand U23018 (N_23018,N_22777,N_22974);
and U23019 (N_23019,N_22818,N_22867);
nand U23020 (N_23020,N_22825,N_22982);
or U23021 (N_23021,N_22840,N_22891);
nand U23022 (N_23022,N_22815,N_22869);
and U23023 (N_23023,N_22783,N_22804);
nor U23024 (N_23024,N_22969,N_22936);
or U23025 (N_23025,N_22894,N_22893);
nand U23026 (N_23026,N_22873,N_22792);
or U23027 (N_23027,N_22786,N_22768);
nor U23028 (N_23028,N_22794,N_22765);
nor U23029 (N_23029,N_22838,N_22959);
and U23030 (N_23030,N_22915,N_22773);
and U23031 (N_23031,N_22902,N_22900);
and U23032 (N_23032,N_22920,N_22841);
or U23033 (N_23033,N_22823,N_22906);
nand U23034 (N_23034,N_22928,N_22912);
and U23035 (N_23035,N_22941,N_22992);
and U23036 (N_23036,N_22801,N_22904);
nand U23037 (N_23037,N_22997,N_22846);
xnor U23038 (N_23038,N_22896,N_22753);
nand U23039 (N_23039,N_22810,N_22751);
xnor U23040 (N_23040,N_22913,N_22881);
nand U23041 (N_23041,N_22987,N_22821);
nor U23042 (N_23042,N_22865,N_22995);
xor U23043 (N_23043,N_22882,N_22921);
and U23044 (N_23044,N_22791,N_22892);
xor U23045 (N_23045,N_22899,N_22955);
or U23046 (N_23046,N_22871,N_22835);
and U23047 (N_23047,N_22850,N_22837);
nor U23048 (N_23048,N_22877,N_22872);
or U23049 (N_23049,N_22852,N_22973);
or U23050 (N_23050,N_22989,N_22875);
nand U23051 (N_23051,N_22976,N_22851);
nand U23052 (N_23052,N_22878,N_22764);
nor U23053 (N_23053,N_22962,N_22970);
xor U23054 (N_23054,N_22834,N_22988);
nand U23055 (N_23055,N_22827,N_22762);
xor U23056 (N_23056,N_22931,N_22935);
or U23057 (N_23057,N_22953,N_22910);
nand U23058 (N_23058,N_22845,N_22814);
and U23059 (N_23059,N_22863,N_22769);
xor U23060 (N_23060,N_22957,N_22886);
xnor U23061 (N_23061,N_22986,N_22868);
and U23062 (N_23062,N_22934,N_22958);
nand U23063 (N_23063,N_22797,N_22933);
or U23064 (N_23064,N_22788,N_22844);
nand U23065 (N_23065,N_22984,N_22937);
nor U23066 (N_23066,N_22908,N_22993);
or U23067 (N_23067,N_22806,N_22968);
or U23068 (N_23068,N_22907,N_22780);
nor U23069 (N_23069,N_22996,N_22966);
nor U23070 (N_23070,N_22858,N_22767);
nand U23071 (N_23071,N_22870,N_22798);
nand U23072 (N_23072,N_22924,N_22983);
and U23073 (N_23073,N_22898,N_22774);
nor U23074 (N_23074,N_22778,N_22926);
nand U23075 (N_23075,N_22949,N_22905);
nand U23076 (N_23076,N_22763,N_22880);
xnor U23077 (N_23077,N_22857,N_22883);
and U23078 (N_23078,N_22961,N_22861);
nand U23079 (N_23079,N_22772,N_22839);
or U23080 (N_23080,N_22849,N_22779);
nor U23081 (N_23081,N_22816,N_22950);
nor U23082 (N_23082,N_22888,N_22795);
nor U23083 (N_23083,N_22807,N_22925);
xor U23084 (N_23084,N_22874,N_22999);
and U23085 (N_23085,N_22853,N_22836);
nor U23086 (N_23086,N_22981,N_22759);
nand U23087 (N_23087,N_22775,N_22812);
and U23088 (N_23088,N_22832,N_22932);
nand U23089 (N_23089,N_22876,N_22787);
or U23090 (N_23090,N_22866,N_22960);
or U23091 (N_23091,N_22942,N_22944);
nand U23092 (N_23092,N_22964,N_22972);
nor U23093 (N_23093,N_22796,N_22847);
nand U23094 (N_23094,N_22994,N_22887);
nor U23095 (N_23095,N_22940,N_22761);
or U23096 (N_23096,N_22758,N_22967);
and U23097 (N_23097,N_22819,N_22843);
nor U23098 (N_23098,N_22971,N_22990);
nor U23099 (N_23099,N_22948,N_22956);
nand U23100 (N_23100,N_22808,N_22854);
xnor U23101 (N_23101,N_22855,N_22757);
or U23102 (N_23102,N_22909,N_22914);
xnor U23103 (N_23103,N_22979,N_22771);
and U23104 (N_23104,N_22980,N_22811);
xnor U23105 (N_23105,N_22756,N_22833);
or U23106 (N_23106,N_22813,N_22831);
or U23107 (N_23107,N_22803,N_22781);
or U23108 (N_23108,N_22822,N_22951);
nor U23109 (N_23109,N_22927,N_22755);
or U23110 (N_23110,N_22884,N_22917);
nor U23111 (N_23111,N_22998,N_22938);
xor U23112 (N_23112,N_22911,N_22897);
nor U23113 (N_23113,N_22802,N_22895);
nor U23114 (N_23114,N_22929,N_22946);
nor U23115 (N_23115,N_22826,N_22963);
or U23116 (N_23116,N_22760,N_22885);
and U23117 (N_23117,N_22952,N_22977);
and U23118 (N_23118,N_22985,N_22919);
or U23119 (N_23119,N_22879,N_22789);
or U23120 (N_23120,N_22754,N_22782);
nor U23121 (N_23121,N_22766,N_22848);
or U23122 (N_23122,N_22930,N_22943);
xnor U23123 (N_23123,N_22800,N_22829);
nand U23124 (N_23124,N_22856,N_22918);
nor U23125 (N_23125,N_22854,N_22893);
nor U23126 (N_23126,N_22997,N_22992);
nand U23127 (N_23127,N_22947,N_22903);
or U23128 (N_23128,N_22888,N_22997);
nand U23129 (N_23129,N_22878,N_22941);
or U23130 (N_23130,N_22880,N_22975);
nor U23131 (N_23131,N_22890,N_22911);
and U23132 (N_23132,N_22820,N_22828);
nand U23133 (N_23133,N_22865,N_22948);
nand U23134 (N_23134,N_22842,N_22943);
nor U23135 (N_23135,N_22869,N_22852);
xor U23136 (N_23136,N_22992,N_22801);
or U23137 (N_23137,N_22761,N_22987);
xnor U23138 (N_23138,N_22941,N_22776);
and U23139 (N_23139,N_22847,N_22999);
and U23140 (N_23140,N_22931,N_22978);
and U23141 (N_23141,N_22831,N_22982);
and U23142 (N_23142,N_22935,N_22843);
nor U23143 (N_23143,N_22783,N_22843);
nand U23144 (N_23144,N_22856,N_22891);
nor U23145 (N_23145,N_22904,N_22848);
or U23146 (N_23146,N_22981,N_22851);
and U23147 (N_23147,N_22803,N_22945);
nor U23148 (N_23148,N_22933,N_22943);
nand U23149 (N_23149,N_22973,N_22950);
and U23150 (N_23150,N_22884,N_22772);
nand U23151 (N_23151,N_22815,N_22882);
nor U23152 (N_23152,N_22826,N_22821);
nand U23153 (N_23153,N_22770,N_22955);
nand U23154 (N_23154,N_22756,N_22951);
nor U23155 (N_23155,N_22957,N_22902);
nand U23156 (N_23156,N_22777,N_22859);
or U23157 (N_23157,N_22936,N_22764);
or U23158 (N_23158,N_22964,N_22963);
and U23159 (N_23159,N_22938,N_22939);
or U23160 (N_23160,N_22892,N_22920);
and U23161 (N_23161,N_22796,N_22913);
and U23162 (N_23162,N_22755,N_22916);
and U23163 (N_23163,N_22895,N_22790);
xor U23164 (N_23164,N_22912,N_22837);
xnor U23165 (N_23165,N_22983,N_22895);
xor U23166 (N_23166,N_22761,N_22833);
nand U23167 (N_23167,N_22764,N_22810);
and U23168 (N_23168,N_22812,N_22831);
nand U23169 (N_23169,N_22860,N_22972);
xnor U23170 (N_23170,N_22866,N_22986);
and U23171 (N_23171,N_22925,N_22946);
nand U23172 (N_23172,N_22945,N_22768);
nand U23173 (N_23173,N_22919,N_22843);
nor U23174 (N_23174,N_22945,N_22841);
or U23175 (N_23175,N_22758,N_22881);
nand U23176 (N_23176,N_22805,N_22790);
nor U23177 (N_23177,N_22858,N_22924);
nor U23178 (N_23178,N_22770,N_22914);
nand U23179 (N_23179,N_22957,N_22787);
or U23180 (N_23180,N_22860,N_22873);
nand U23181 (N_23181,N_22800,N_22792);
xor U23182 (N_23182,N_22797,N_22764);
xor U23183 (N_23183,N_22927,N_22898);
and U23184 (N_23184,N_22971,N_22948);
or U23185 (N_23185,N_22962,N_22980);
or U23186 (N_23186,N_22888,N_22788);
nand U23187 (N_23187,N_22771,N_22991);
or U23188 (N_23188,N_22926,N_22971);
and U23189 (N_23189,N_22756,N_22853);
xnor U23190 (N_23190,N_22856,N_22940);
nor U23191 (N_23191,N_22792,N_22876);
and U23192 (N_23192,N_22776,N_22990);
xor U23193 (N_23193,N_22947,N_22791);
nand U23194 (N_23194,N_22906,N_22996);
nand U23195 (N_23195,N_22830,N_22992);
nand U23196 (N_23196,N_22912,N_22827);
or U23197 (N_23197,N_22880,N_22971);
nand U23198 (N_23198,N_22834,N_22951);
nor U23199 (N_23199,N_22858,N_22770);
xor U23200 (N_23200,N_22880,N_22832);
nor U23201 (N_23201,N_22921,N_22765);
nor U23202 (N_23202,N_22989,N_22884);
nand U23203 (N_23203,N_22881,N_22900);
and U23204 (N_23204,N_22902,N_22916);
and U23205 (N_23205,N_22879,N_22754);
and U23206 (N_23206,N_22790,N_22765);
nor U23207 (N_23207,N_22799,N_22971);
xor U23208 (N_23208,N_22819,N_22760);
or U23209 (N_23209,N_22850,N_22821);
or U23210 (N_23210,N_22849,N_22755);
nand U23211 (N_23211,N_22859,N_22774);
or U23212 (N_23212,N_22820,N_22998);
nor U23213 (N_23213,N_22812,N_22807);
xnor U23214 (N_23214,N_22930,N_22868);
nor U23215 (N_23215,N_22774,N_22998);
or U23216 (N_23216,N_22816,N_22917);
nand U23217 (N_23217,N_22848,N_22989);
xor U23218 (N_23218,N_22935,N_22813);
xor U23219 (N_23219,N_22915,N_22993);
nor U23220 (N_23220,N_22765,N_22941);
nand U23221 (N_23221,N_22853,N_22868);
or U23222 (N_23222,N_22837,N_22861);
nand U23223 (N_23223,N_22828,N_22846);
xor U23224 (N_23224,N_22996,N_22922);
and U23225 (N_23225,N_22818,N_22920);
xor U23226 (N_23226,N_22785,N_22796);
xor U23227 (N_23227,N_22820,N_22786);
and U23228 (N_23228,N_22833,N_22805);
or U23229 (N_23229,N_22961,N_22995);
nand U23230 (N_23230,N_22790,N_22993);
nor U23231 (N_23231,N_22845,N_22915);
nor U23232 (N_23232,N_22941,N_22846);
nand U23233 (N_23233,N_22848,N_22877);
xnor U23234 (N_23234,N_22756,N_22868);
nor U23235 (N_23235,N_22975,N_22917);
nand U23236 (N_23236,N_22950,N_22997);
and U23237 (N_23237,N_22838,N_22875);
nand U23238 (N_23238,N_22772,N_22847);
nor U23239 (N_23239,N_22929,N_22801);
nor U23240 (N_23240,N_22977,N_22871);
nor U23241 (N_23241,N_22884,N_22760);
xnor U23242 (N_23242,N_22760,N_22893);
nand U23243 (N_23243,N_22846,N_22854);
or U23244 (N_23244,N_22853,N_22978);
and U23245 (N_23245,N_22839,N_22783);
or U23246 (N_23246,N_22975,N_22865);
xor U23247 (N_23247,N_22963,N_22992);
and U23248 (N_23248,N_22759,N_22877);
xor U23249 (N_23249,N_22926,N_22789);
nand U23250 (N_23250,N_23169,N_23208);
nand U23251 (N_23251,N_23108,N_23072);
nand U23252 (N_23252,N_23155,N_23148);
nor U23253 (N_23253,N_23179,N_23074);
or U23254 (N_23254,N_23113,N_23156);
nor U23255 (N_23255,N_23233,N_23094);
or U23256 (N_23256,N_23191,N_23050);
nor U23257 (N_23257,N_23023,N_23246);
xor U23258 (N_23258,N_23249,N_23006);
or U23259 (N_23259,N_23151,N_23175);
and U23260 (N_23260,N_23088,N_23157);
and U23261 (N_23261,N_23171,N_23062);
nor U23262 (N_23262,N_23209,N_23036);
nand U23263 (N_23263,N_23007,N_23055);
xnor U23264 (N_23264,N_23207,N_23183);
and U23265 (N_23265,N_23044,N_23166);
or U23266 (N_23266,N_23231,N_23133);
xor U23267 (N_23267,N_23187,N_23118);
or U23268 (N_23268,N_23182,N_23032);
nand U23269 (N_23269,N_23004,N_23145);
nand U23270 (N_23270,N_23200,N_23135);
nor U23271 (N_23271,N_23170,N_23185);
nor U23272 (N_23272,N_23221,N_23218);
and U23273 (N_23273,N_23026,N_23122);
xnor U23274 (N_23274,N_23079,N_23142);
nand U23275 (N_23275,N_23011,N_23053);
nor U23276 (N_23276,N_23212,N_23103);
xor U23277 (N_23277,N_23150,N_23238);
xor U23278 (N_23278,N_23025,N_23049);
or U23279 (N_23279,N_23019,N_23205);
nand U23280 (N_23280,N_23139,N_23125);
xnor U23281 (N_23281,N_23093,N_23137);
or U23282 (N_23282,N_23092,N_23048);
or U23283 (N_23283,N_23102,N_23115);
nand U23284 (N_23284,N_23227,N_23104);
nand U23285 (N_23285,N_23162,N_23146);
nor U23286 (N_23286,N_23159,N_23203);
xor U23287 (N_23287,N_23215,N_23127);
nand U23288 (N_23288,N_23041,N_23248);
xor U23289 (N_23289,N_23097,N_23144);
nand U23290 (N_23290,N_23022,N_23232);
nor U23291 (N_23291,N_23163,N_23095);
nor U23292 (N_23292,N_23016,N_23174);
and U23293 (N_23293,N_23134,N_23210);
xor U23294 (N_23294,N_23172,N_23199);
xnor U23295 (N_23295,N_23120,N_23213);
and U23296 (N_23296,N_23061,N_23229);
nor U23297 (N_23297,N_23021,N_23136);
xor U23298 (N_23298,N_23167,N_23168);
and U23299 (N_23299,N_23027,N_23116);
or U23300 (N_23300,N_23081,N_23119);
and U23301 (N_23301,N_23214,N_23003);
nor U23302 (N_23302,N_23077,N_23222);
and U23303 (N_23303,N_23070,N_23180);
or U23304 (N_23304,N_23206,N_23177);
and U23305 (N_23305,N_23043,N_23076);
nor U23306 (N_23306,N_23176,N_23018);
nor U23307 (N_23307,N_23065,N_23158);
or U23308 (N_23308,N_23105,N_23005);
xnor U23309 (N_23309,N_23189,N_23178);
and U23310 (N_23310,N_23236,N_23066);
or U23311 (N_23311,N_23243,N_23059);
or U23312 (N_23312,N_23201,N_23010);
and U23313 (N_23313,N_23031,N_23117);
or U23314 (N_23314,N_23051,N_23078);
nor U23315 (N_23315,N_23217,N_23219);
xnor U23316 (N_23316,N_23245,N_23064);
xor U23317 (N_23317,N_23247,N_23198);
and U23318 (N_23318,N_23153,N_23143);
and U23319 (N_23319,N_23235,N_23126);
xnor U23320 (N_23320,N_23190,N_23035);
nor U23321 (N_23321,N_23039,N_23195);
and U23322 (N_23322,N_23000,N_23196);
and U23323 (N_23323,N_23058,N_23147);
and U23324 (N_23324,N_23047,N_23193);
xnor U23325 (N_23325,N_23071,N_23098);
xor U23326 (N_23326,N_23224,N_23056);
nor U23327 (N_23327,N_23067,N_23054);
or U23328 (N_23328,N_23015,N_23140);
and U23329 (N_23329,N_23164,N_23086);
and U23330 (N_23330,N_23211,N_23090);
and U23331 (N_23331,N_23240,N_23197);
xor U23332 (N_23332,N_23068,N_23040);
and U23333 (N_23333,N_23083,N_23087);
xor U23334 (N_23334,N_23112,N_23091);
or U23335 (N_23335,N_23152,N_23225);
nor U23336 (N_23336,N_23063,N_23013);
or U23337 (N_23337,N_23202,N_23111);
or U23338 (N_23338,N_23029,N_23165);
and U23339 (N_23339,N_23106,N_23138);
nor U23340 (N_23340,N_23234,N_23080);
and U23341 (N_23341,N_23042,N_23130);
nor U23342 (N_23342,N_23160,N_23024);
and U23343 (N_23343,N_23107,N_23033);
or U23344 (N_23344,N_23096,N_23109);
or U23345 (N_23345,N_23001,N_23131);
nor U23346 (N_23346,N_23161,N_23194);
nand U23347 (N_23347,N_23237,N_23014);
nand U23348 (N_23348,N_23192,N_23220);
and U23349 (N_23349,N_23181,N_23052);
xor U23350 (N_23350,N_23244,N_23008);
nand U23351 (N_23351,N_23114,N_23204);
nor U23352 (N_23352,N_23017,N_23045);
and U23353 (N_23353,N_23141,N_23020);
or U23354 (N_23354,N_23060,N_23123);
nand U23355 (N_23355,N_23030,N_23149);
xor U23356 (N_23356,N_23002,N_23057);
and U23357 (N_23357,N_23230,N_23012);
nand U23358 (N_23358,N_23188,N_23099);
xor U23359 (N_23359,N_23154,N_23028);
xnor U23360 (N_23360,N_23228,N_23242);
nand U23361 (N_23361,N_23101,N_23223);
or U23362 (N_23362,N_23034,N_23084);
nand U23363 (N_23363,N_23173,N_23226);
nand U23364 (N_23364,N_23216,N_23089);
and U23365 (N_23365,N_23186,N_23038);
or U23366 (N_23366,N_23037,N_23129);
and U23367 (N_23367,N_23121,N_23110);
or U23368 (N_23368,N_23132,N_23124);
nor U23369 (N_23369,N_23069,N_23128);
nand U23370 (N_23370,N_23085,N_23239);
nand U23371 (N_23371,N_23082,N_23241);
and U23372 (N_23372,N_23073,N_23009);
or U23373 (N_23373,N_23075,N_23184);
or U23374 (N_23374,N_23100,N_23046);
or U23375 (N_23375,N_23076,N_23145);
nor U23376 (N_23376,N_23124,N_23204);
and U23377 (N_23377,N_23208,N_23143);
xor U23378 (N_23378,N_23055,N_23056);
and U23379 (N_23379,N_23057,N_23137);
nor U23380 (N_23380,N_23239,N_23153);
xor U23381 (N_23381,N_23131,N_23196);
nand U23382 (N_23382,N_23225,N_23132);
nor U23383 (N_23383,N_23120,N_23183);
nor U23384 (N_23384,N_23249,N_23051);
and U23385 (N_23385,N_23022,N_23100);
nand U23386 (N_23386,N_23181,N_23051);
or U23387 (N_23387,N_23086,N_23215);
or U23388 (N_23388,N_23102,N_23065);
or U23389 (N_23389,N_23150,N_23236);
nor U23390 (N_23390,N_23116,N_23173);
xnor U23391 (N_23391,N_23229,N_23056);
or U23392 (N_23392,N_23166,N_23247);
xnor U23393 (N_23393,N_23160,N_23018);
nand U23394 (N_23394,N_23246,N_23194);
nor U23395 (N_23395,N_23156,N_23029);
xor U23396 (N_23396,N_23010,N_23032);
and U23397 (N_23397,N_23107,N_23108);
and U23398 (N_23398,N_23153,N_23161);
xnor U23399 (N_23399,N_23009,N_23199);
xor U23400 (N_23400,N_23183,N_23031);
nand U23401 (N_23401,N_23019,N_23058);
and U23402 (N_23402,N_23105,N_23221);
and U23403 (N_23403,N_23095,N_23108);
nand U23404 (N_23404,N_23047,N_23230);
or U23405 (N_23405,N_23091,N_23074);
nor U23406 (N_23406,N_23034,N_23029);
nand U23407 (N_23407,N_23067,N_23138);
nor U23408 (N_23408,N_23143,N_23220);
xor U23409 (N_23409,N_23181,N_23215);
and U23410 (N_23410,N_23218,N_23028);
or U23411 (N_23411,N_23050,N_23087);
xnor U23412 (N_23412,N_23172,N_23248);
nor U23413 (N_23413,N_23005,N_23074);
or U23414 (N_23414,N_23000,N_23092);
nand U23415 (N_23415,N_23179,N_23240);
or U23416 (N_23416,N_23058,N_23092);
nand U23417 (N_23417,N_23019,N_23104);
and U23418 (N_23418,N_23031,N_23232);
xor U23419 (N_23419,N_23246,N_23231);
and U23420 (N_23420,N_23124,N_23058);
nand U23421 (N_23421,N_23158,N_23097);
or U23422 (N_23422,N_23057,N_23223);
xor U23423 (N_23423,N_23156,N_23166);
nor U23424 (N_23424,N_23043,N_23074);
xor U23425 (N_23425,N_23179,N_23143);
xor U23426 (N_23426,N_23044,N_23051);
nor U23427 (N_23427,N_23061,N_23209);
xor U23428 (N_23428,N_23242,N_23249);
and U23429 (N_23429,N_23121,N_23047);
and U23430 (N_23430,N_23001,N_23049);
and U23431 (N_23431,N_23004,N_23205);
or U23432 (N_23432,N_23180,N_23030);
nor U23433 (N_23433,N_23113,N_23168);
nor U23434 (N_23434,N_23094,N_23245);
nand U23435 (N_23435,N_23060,N_23042);
nor U23436 (N_23436,N_23183,N_23140);
and U23437 (N_23437,N_23193,N_23228);
and U23438 (N_23438,N_23010,N_23014);
nor U23439 (N_23439,N_23001,N_23096);
and U23440 (N_23440,N_23137,N_23008);
xor U23441 (N_23441,N_23147,N_23127);
or U23442 (N_23442,N_23112,N_23072);
nor U23443 (N_23443,N_23106,N_23226);
nand U23444 (N_23444,N_23137,N_23040);
xnor U23445 (N_23445,N_23171,N_23232);
xnor U23446 (N_23446,N_23107,N_23188);
nor U23447 (N_23447,N_23149,N_23176);
and U23448 (N_23448,N_23132,N_23100);
nand U23449 (N_23449,N_23022,N_23175);
and U23450 (N_23450,N_23030,N_23101);
nor U23451 (N_23451,N_23207,N_23138);
and U23452 (N_23452,N_23083,N_23230);
nor U23453 (N_23453,N_23030,N_23099);
or U23454 (N_23454,N_23089,N_23001);
xnor U23455 (N_23455,N_23093,N_23118);
or U23456 (N_23456,N_23227,N_23236);
nand U23457 (N_23457,N_23041,N_23174);
nand U23458 (N_23458,N_23216,N_23177);
and U23459 (N_23459,N_23224,N_23120);
nand U23460 (N_23460,N_23159,N_23130);
or U23461 (N_23461,N_23190,N_23178);
xnor U23462 (N_23462,N_23044,N_23146);
nand U23463 (N_23463,N_23125,N_23144);
or U23464 (N_23464,N_23002,N_23102);
xnor U23465 (N_23465,N_23101,N_23116);
nor U23466 (N_23466,N_23053,N_23080);
nand U23467 (N_23467,N_23196,N_23189);
and U23468 (N_23468,N_23221,N_23223);
or U23469 (N_23469,N_23200,N_23220);
nand U23470 (N_23470,N_23080,N_23099);
nand U23471 (N_23471,N_23231,N_23215);
nor U23472 (N_23472,N_23000,N_23115);
nand U23473 (N_23473,N_23184,N_23137);
nor U23474 (N_23474,N_23101,N_23004);
nor U23475 (N_23475,N_23145,N_23138);
xor U23476 (N_23476,N_23037,N_23071);
nor U23477 (N_23477,N_23151,N_23022);
or U23478 (N_23478,N_23247,N_23117);
nand U23479 (N_23479,N_23033,N_23043);
and U23480 (N_23480,N_23177,N_23049);
nor U23481 (N_23481,N_23124,N_23074);
xor U23482 (N_23482,N_23229,N_23068);
and U23483 (N_23483,N_23085,N_23140);
nor U23484 (N_23484,N_23198,N_23096);
nor U23485 (N_23485,N_23184,N_23172);
nand U23486 (N_23486,N_23086,N_23162);
nor U23487 (N_23487,N_23227,N_23062);
xor U23488 (N_23488,N_23051,N_23062);
xor U23489 (N_23489,N_23175,N_23248);
nand U23490 (N_23490,N_23139,N_23126);
and U23491 (N_23491,N_23096,N_23008);
or U23492 (N_23492,N_23137,N_23156);
or U23493 (N_23493,N_23110,N_23118);
nand U23494 (N_23494,N_23083,N_23014);
nand U23495 (N_23495,N_23154,N_23064);
and U23496 (N_23496,N_23204,N_23009);
or U23497 (N_23497,N_23076,N_23137);
or U23498 (N_23498,N_23118,N_23128);
nand U23499 (N_23499,N_23183,N_23105);
or U23500 (N_23500,N_23461,N_23447);
nor U23501 (N_23501,N_23473,N_23275);
nand U23502 (N_23502,N_23493,N_23403);
nand U23503 (N_23503,N_23302,N_23332);
nor U23504 (N_23504,N_23353,N_23365);
xnor U23505 (N_23505,N_23456,N_23494);
xor U23506 (N_23506,N_23422,N_23391);
or U23507 (N_23507,N_23417,N_23415);
or U23508 (N_23508,N_23257,N_23326);
nand U23509 (N_23509,N_23289,N_23449);
and U23510 (N_23510,N_23484,N_23342);
nor U23511 (N_23511,N_23262,N_23250);
or U23512 (N_23512,N_23467,N_23421);
nand U23513 (N_23513,N_23260,N_23310);
nand U23514 (N_23514,N_23475,N_23393);
xnor U23515 (N_23515,N_23282,N_23253);
and U23516 (N_23516,N_23448,N_23256);
nor U23517 (N_23517,N_23407,N_23396);
xor U23518 (N_23518,N_23291,N_23371);
and U23519 (N_23519,N_23290,N_23278);
and U23520 (N_23520,N_23347,N_23344);
or U23521 (N_23521,N_23444,N_23468);
and U23522 (N_23522,N_23434,N_23496);
xor U23523 (N_23523,N_23269,N_23384);
nand U23524 (N_23524,N_23352,N_23273);
and U23525 (N_23525,N_23258,N_23462);
nand U23526 (N_23526,N_23427,N_23404);
xor U23527 (N_23527,N_23374,N_23433);
nor U23528 (N_23528,N_23418,N_23478);
nand U23529 (N_23529,N_23349,N_23408);
and U23530 (N_23530,N_23387,N_23416);
or U23531 (N_23531,N_23409,N_23259);
nor U23532 (N_23532,N_23399,N_23499);
nand U23533 (N_23533,N_23370,N_23450);
nor U23534 (N_23534,N_23363,N_23361);
and U23535 (N_23535,N_23451,N_23491);
and U23536 (N_23536,N_23277,N_23312);
or U23537 (N_23537,N_23263,N_23339);
nor U23538 (N_23538,N_23308,N_23364);
xnor U23539 (N_23539,N_23319,N_23329);
or U23540 (N_23540,N_23476,N_23483);
nand U23541 (N_23541,N_23330,N_23428);
nand U23542 (N_23542,N_23360,N_23410);
nor U23543 (N_23543,N_23272,N_23276);
nor U23544 (N_23544,N_23401,N_23279);
xnor U23545 (N_23545,N_23252,N_23293);
xor U23546 (N_23546,N_23327,N_23285);
nand U23547 (N_23547,N_23299,N_23367);
or U23548 (N_23548,N_23379,N_23498);
nor U23549 (N_23549,N_23255,N_23333);
and U23550 (N_23550,N_23322,N_23446);
and U23551 (N_23551,N_23264,N_23430);
or U23552 (N_23552,N_23495,N_23459);
nand U23553 (N_23553,N_23348,N_23389);
or U23554 (N_23554,N_23429,N_23472);
nand U23555 (N_23555,N_23423,N_23378);
or U23556 (N_23556,N_23270,N_23454);
or U23557 (N_23557,N_23377,N_23355);
nand U23558 (N_23558,N_23400,N_23437);
xor U23559 (N_23559,N_23373,N_23338);
xor U23560 (N_23560,N_23296,N_23479);
and U23561 (N_23561,N_23311,N_23354);
or U23562 (N_23562,N_23366,N_23283);
nand U23563 (N_23563,N_23426,N_23394);
nor U23564 (N_23564,N_23414,N_23323);
nor U23565 (N_23565,N_23280,N_23411);
and U23566 (N_23566,N_23424,N_23318);
nor U23567 (N_23567,N_23439,N_23435);
or U23568 (N_23568,N_23304,N_23492);
xnor U23569 (N_23569,N_23261,N_23469);
and U23570 (N_23570,N_23324,N_23369);
xnor U23571 (N_23571,N_23301,N_23268);
nand U23572 (N_23572,N_23436,N_23341);
xor U23573 (N_23573,N_23345,N_23376);
or U23574 (N_23574,N_23266,N_23406);
nand U23575 (N_23575,N_23337,N_23490);
nor U23576 (N_23576,N_23271,N_23357);
nand U23577 (N_23577,N_23316,N_23488);
or U23578 (N_23578,N_23481,N_23317);
xor U23579 (N_23579,N_23300,N_23368);
xor U23580 (N_23580,N_23489,N_23265);
xor U23581 (N_23581,N_23432,N_23390);
xor U23582 (N_23582,N_23482,N_23474);
or U23583 (N_23583,N_23381,N_23325);
nor U23584 (N_23584,N_23440,N_23477);
xor U23585 (N_23585,N_23425,N_23438);
nand U23586 (N_23586,N_23284,N_23497);
and U23587 (N_23587,N_23457,N_23287);
nand U23588 (N_23588,N_23386,N_23463);
nor U23589 (N_23589,N_23356,N_23362);
and U23590 (N_23590,N_23458,N_23346);
nor U23591 (N_23591,N_23288,N_23350);
and U23592 (N_23592,N_23420,N_23292);
nor U23593 (N_23593,N_23382,N_23385);
nor U23594 (N_23594,N_23334,N_23331);
nor U23595 (N_23595,N_23460,N_23254);
and U23596 (N_23596,N_23295,N_23313);
nor U23597 (N_23597,N_23297,N_23452);
xor U23598 (N_23598,N_23306,N_23395);
xor U23599 (N_23599,N_23397,N_23485);
and U23600 (N_23600,N_23464,N_23281);
nor U23601 (N_23601,N_23286,N_23413);
and U23602 (N_23602,N_23487,N_23466);
and U23603 (N_23603,N_23303,N_23358);
and U23604 (N_23604,N_23314,N_23298);
nor U23605 (N_23605,N_23336,N_23392);
and U23606 (N_23606,N_23470,N_23471);
nand U23607 (N_23607,N_23274,N_23402);
nand U23608 (N_23608,N_23480,N_23294);
xor U23609 (N_23609,N_23453,N_23320);
xnor U23610 (N_23610,N_23441,N_23465);
and U23611 (N_23611,N_23335,N_23380);
xor U23612 (N_23612,N_23305,N_23405);
nor U23613 (N_23613,N_23351,N_23251);
and U23614 (N_23614,N_23328,N_23309);
nor U23615 (N_23615,N_23431,N_23359);
and U23616 (N_23616,N_23315,N_23455);
nor U23617 (N_23617,N_23442,N_23443);
and U23618 (N_23618,N_23383,N_23419);
xor U23619 (N_23619,N_23388,N_23486);
nand U23620 (N_23620,N_23343,N_23340);
nor U23621 (N_23621,N_23375,N_23267);
nor U23622 (N_23622,N_23307,N_23372);
and U23623 (N_23623,N_23398,N_23321);
or U23624 (N_23624,N_23445,N_23412);
nand U23625 (N_23625,N_23409,N_23483);
nor U23626 (N_23626,N_23332,N_23319);
xor U23627 (N_23627,N_23358,N_23285);
and U23628 (N_23628,N_23461,N_23432);
and U23629 (N_23629,N_23439,N_23349);
xnor U23630 (N_23630,N_23331,N_23406);
xnor U23631 (N_23631,N_23316,N_23402);
xor U23632 (N_23632,N_23263,N_23377);
nand U23633 (N_23633,N_23465,N_23397);
nor U23634 (N_23634,N_23462,N_23441);
nand U23635 (N_23635,N_23273,N_23396);
nor U23636 (N_23636,N_23408,N_23463);
xnor U23637 (N_23637,N_23498,N_23393);
nand U23638 (N_23638,N_23321,N_23292);
and U23639 (N_23639,N_23429,N_23302);
xnor U23640 (N_23640,N_23466,N_23362);
xor U23641 (N_23641,N_23345,N_23279);
and U23642 (N_23642,N_23381,N_23291);
nor U23643 (N_23643,N_23469,N_23259);
nor U23644 (N_23644,N_23395,N_23415);
or U23645 (N_23645,N_23287,N_23325);
xor U23646 (N_23646,N_23295,N_23469);
and U23647 (N_23647,N_23463,N_23375);
nor U23648 (N_23648,N_23470,N_23368);
and U23649 (N_23649,N_23262,N_23441);
nand U23650 (N_23650,N_23466,N_23429);
and U23651 (N_23651,N_23344,N_23473);
nand U23652 (N_23652,N_23319,N_23349);
and U23653 (N_23653,N_23282,N_23267);
and U23654 (N_23654,N_23420,N_23439);
nor U23655 (N_23655,N_23379,N_23484);
nand U23656 (N_23656,N_23413,N_23407);
nand U23657 (N_23657,N_23407,N_23439);
or U23658 (N_23658,N_23274,N_23487);
nor U23659 (N_23659,N_23267,N_23483);
nand U23660 (N_23660,N_23312,N_23492);
or U23661 (N_23661,N_23361,N_23399);
or U23662 (N_23662,N_23353,N_23401);
and U23663 (N_23663,N_23321,N_23393);
and U23664 (N_23664,N_23378,N_23464);
nand U23665 (N_23665,N_23458,N_23392);
or U23666 (N_23666,N_23324,N_23279);
xnor U23667 (N_23667,N_23446,N_23486);
nand U23668 (N_23668,N_23261,N_23446);
or U23669 (N_23669,N_23321,N_23332);
or U23670 (N_23670,N_23427,N_23479);
xor U23671 (N_23671,N_23358,N_23289);
nor U23672 (N_23672,N_23437,N_23293);
nand U23673 (N_23673,N_23374,N_23349);
and U23674 (N_23674,N_23346,N_23495);
xnor U23675 (N_23675,N_23280,N_23432);
and U23676 (N_23676,N_23467,N_23322);
nor U23677 (N_23677,N_23466,N_23268);
xor U23678 (N_23678,N_23322,N_23303);
xnor U23679 (N_23679,N_23460,N_23349);
and U23680 (N_23680,N_23402,N_23496);
nor U23681 (N_23681,N_23343,N_23414);
nand U23682 (N_23682,N_23402,N_23429);
or U23683 (N_23683,N_23317,N_23297);
nand U23684 (N_23684,N_23497,N_23425);
xnor U23685 (N_23685,N_23383,N_23343);
or U23686 (N_23686,N_23336,N_23351);
nand U23687 (N_23687,N_23433,N_23469);
and U23688 (N_23688,N_23376,N_23326);
nand U23689 (N_23689,N_23346,N_23347);
nor U23690 (N_23690,N_23283,N_23423);
or U23691 (N_23691,N_23252,N_23422);
nor U23692 (N_23692,N_23393,N_23373);
xor U23693 (N_23693,N_23472,N_23377);
or U23694 (N_23694,N_23398,N_23291);
and U23695 (N_23695,N_23362,N_23495);
nand U23696 (N_23696,N_23438,N_23313);
or U23697 (N_23697,N_23308,N_23285);
and U23698 (N_23698,N_23366,N_23411);
nand U23699 (N_23699,N_23489,N_23451);
nand U23700 (N_23700,N_23478,N_23407);
nand U23701 (N_23701,N_23401,N_23449);
nor U23702 (N_23702,N_23279,N_23314);
nor U23703 (N_23703,N_23392,N_23253);
xor U23704 (N_23704,N_23277,N_23313);
or U23705 (N_23705,N_23494,N_23488);
nand U23706 (N_23706,N_23276,N_23292);
or U23707 (N_23707,N_23492,N_23329);
nor U23708 (N_23708,N_23357,N_23307);
nand U23709 (N_23709,N_23422,N_23430);
nor U23710 (N_23710,N_23324,N_23257);
and U23711 (N_23711,N_23292,N_23274);
nand U23712 (N_23712,N_23426,N_23263);
nor U23713 (N_23713,N_23478,N_23383);
and U23714 (N_23714,N_23252,N_23329);
or U23715 (N_23715,N_23298,N_23422);
and U23716 (N_23716,N_23260,N_23460);
nor U23717 (N_23717,N_23331,N_23354);
and U23718 (N_23718,N_23448,N_23304);
and U23719 (N_23719,N_23359,N_23497);
nand U23720 (N_23720,N_23445,N_23265);
nor U23721 (N_23721,N_23298,N_23418);
xnor U23722 (N_23722,N_23447,N_23469);
nand U23723 (N_23723,N_23267,N_23390);
or U23724 (N_23724,N_23412,N_23496);
nand U23725 (N_23725,N_23338,N_23263);
or U23726 (N_23726,N_23341,N_23321);
xor U23727 (N_23727,N_23462,N_23329);
or U23728 (N_23728,N_23257,N_23310);
xnor U23729 (N_23729,N_23276,N_23470);
and U23730 (N_23730,N_23354,N_23396);
and U23731 (N_23731,N_23440,N_23257);
and U23732 (N_23732,N_23482,N_23443);
xor U23733 (N_23733,N_23438,N_23427);
nor U23734 (N_23734,N_23388,N_23454);
and U23735 (N_23735,N_23321,N_23314);
nand U23736 (N_23736,N_23357,N_23367);
and U23737 (N_23737,N_23464,N_23447);
nand U23738 (N_23738,N_23458,N_23474);
nor U23739 (N_23739,N_23491,N_23494);
or U23740 (N_23740,N_23402,N_23455);
or U23741 (N_23741,N_23352,N_23386);
nor U23742 (N_23742,N_23316,N_23412);
nand U23743 (N_23743,N_23409,N_23340);
xor U23744 (N_23744,N_23343,N_23305);
nand U23745 (N_23745,N_23407,N_23418);
xnor U23746 (N_23746,N_23259,N_23283);
nor U23747 (N_23747,N_23461,N_23336);
xnor U23748 (N_23748,N_23259,N_23351);
nand U23749 (N_23749,N_23359,N_23415);
nand U23750 (N_23750,N_23604,N_23690);
and U23751 (N_23751,N_23528,N_23667);
nand U23752 (N_23752,N_23566,N_23668);
and U23753 (N_23753,N_23509,N_23717);
nand U23754 (N_23754,N_23647,N_23674);
or U23755 (N_23755,N_23658,N_23738);
or U23756 (N_23756,N_23543,N_23636);
nand U23757 (N_23757,N_23575,N_23714);
or U23758 (N_23758,N_23531,N_23665);
nand U23759 (N_23759,N_23663,N_23680);
and U23760 (N_23760,N_23578,N_23689);
and U23761 (N_23761,N_23541,N_23726);
nor U23762 (N_23762,N_23641,N_23632);
or U23763 (N_23763,N_23615,N_23530);
or U23764 (N_23764,N_23623,N_23540);
and U23765 (N_23765,N_23748,N_23722);
or U23766 (N_23766,N_23691,N_23570);
nand U23767 (N_23767,N_23662,N_23605);
xor U23768 (N_23768,N_23695,N_23661);
xnor U23769 (N_23769,N_23573,N_23542);
nand U23770 (N_23770,N_23525,N_23624);
xor U23771 (N_23771,N_23548,N_23526);
nor U23772 (N_23772,N_23514,N_23574);
and U23773 (N_23773,N_23683,N_23622);
xnor U23774 (N_23774,N_23720,N_23634);
or U23775 (N_23775,N_23594,N_23589);
nand U23776 (N_23776,N_23715,N_23627);
nand U23777 (N_23777,N_23535,N_23611);
nand U23778 (N_23778,N_23602,N_23723);
xnor U23779 (N_23779,N_23648,N_23697);
or U23780 (N_23780,N_23709,N_23679);
xor U23781 (N_23781,N_23568,N_23638);
xor U23782 (N_23782,N_23686,N_23549);
nand U23783 (N_23783,N_23698,N_23546);
or U23784 (N_23784,N_23544,N_23737);
and U23785 (N_23785,N_23584,N_23564);
xnor U23786 (N_23786,N_23593,N_23713);
or U23787 (N_23787,N_23506,N_23613);
xor U23788 (N_23788,N_23612,N_23742);
xor U23789 (N_23789,N_23736,N_23744);
nand U23790 (N_23790,N_23687,N_23743);
and U23791 (N_23791,N_23576,N_23505);
nor U23792 (N_23792,N_23553,N_23614);
and U23793 (N_23793,N_23577,N_23693);
nand U23794 (N_23794,N_23741,N_23705);
or U23795 (N_23795,N_23617,N_23512);
or U23796 (N_23796,N_23702,N_23579);
or U23797 (N_23797,N_23708,N_23650);
nor U23798 (N_23798,N_23590,N_23716);
nand U23799 (N_23799,N_23607,N_23625);
nor U23800 (N_23800,N_23610,N_23601);
nand U23801 (N_23801,N_23652,N_23700);
nand U23802 (N_23802,N_23732,N_23740);
and U23803 (N_23803,N_23630,N_23729);
and U23804 (N_23804,N_23633,N_23563);
xnor U23805 (N_23805,N_23596,N_23735);
xnor U23806 (N_23806,N_23699,N_23646);
or U23807 (N_23807,N_23677,N_23519);
or U23808 (N_23808,N_23500,N_23582);
and U23809 (N_23809,N_23508,N_23725);
xor U23810 (N_23810,N_23556,N_23524);
nor U23811 (N_23811,N_23644,N_23696);
nor U23812 (N_23812,N_23501,N_23597);
or U23813 (N_23813,N_23598,N_23682);
and U23814 (N_23814,N_23704,N_23694);
xor U23815 (N_23815,N_23621,N_23599);
or U23816 (N_23816,N_23551,N_23557);
or U23817 (N_23817,N_23739,N_23560);
nand U23818 (N_23818,N_23547,N_23583);
or U23819 (N_23819,N_23731,N_23626);
nor U23820 (N_23820,N_23718,N_23609);
xnor U23821 (N_23821,N_23504,N_23676);
xnor U23822 (N_23822,N_23628,N_23639);
and U23823 (N_23823,N_23672,N_23527);
nand U23824 (N_23824,N_23719,N_23538);
and U23825 (N_23825,N_23710,N_23520);
or U23826 (N_23826,N_23730,N_23503);
nor U23827 (N_23827,N_23635,N_23747);
and U23828 (N_23828,N_23685,N_23684);
xnor U23829 (N_23829,N_23706,N_23569);
and U23830 (N_23830,N_23532,N_23688);
and U23831 (N_23831,N_23517,N_23643);
or U23832 (N_23832,N_23550,N_23513);
or U23833 (N_23833,N_23681,N_23561);
xor U23834 (N_23834,N_23734,N_23659);
xnor U23835 (N_23835,N_23586,N_23522);
xnor U23836 (N_23836,N_23746,N_23510);
nand U23837 (N_23837,N_23537,N_23728);
or U23838 (N_23838,N_23619,N_23585);
xnor U23839 (N_23839,N_23515,N_23631);
nand U23840 (N_23840,N_23595,N_23592);
xnor U23841 (N_23841,N_23657,N_23701);
nand U23842 (N_23842,N_23580,N_23536);
or U23843 (N_23843,N_23533,N_23507);
xor U23844 (N_23844,N_23523,N_23711);
and U23845 (N_23845,N_23678,N_23673);
xnor U23846 (N_23846,N_23660,N_23671);
or U23847 (N_23847,N_23581,N_23502);
and U23848 (N_23848,N_23649,N_23637);
nor U23849 (N_23849,N_23608,N_23554);
and U23850 (N_23850,N_23651,N_23518);
and U23851 (N_23851,N_23534,N_23600);
and U23852 (N_23852,N_23616,N_23521);
nor U23853 (N_23853,N_23749,N_23555);
nor U23854 (N_23854,N_23645,N_23511);
and U23855 (N_23855,N_23545,N_23552);
and U23856 (N_23856,N_23539,N_23603);
nand U23857 (N_23857,N_23675,N_23588);
nor U23858 (N_23858,N_23559,N_23733);
and U23859 (N_23859,N_23707,N_23618);
or U23860 (N_23860,N_23692,N_23558);
and U23861 (N_23861,N_23572,N_23656);
nor U23862 (N_23862,N_23606,N_23629);
nand U23863 (N_23863,N_23669,N_23745);
xnor U23864 (N_23864,N_23565,N_23703);
nor U23865 (N_23865,N_23640,N_23567);
or U23866 (N_23866,N_23724,N_23529);
xor U23867 (N_23867,N_23620,N_23670);
nand U23868 (N_23868,N_23516,N_23712);
nor U23869 (N_23869,N_23727,N_23571);
nor U23870 (N_23870,N_23653,N_23587);
nor U23871 (N_23871,N_23642,N_23655);
or U23872 (N_23872,N_23664,N_23562);
and U23873 (N_23873,N_23654,N_23591);
xor U23874 (N_23874,N_23666,N_23721);
or U23875 (N_23875,N_23650,N_23567);
nand U23876 (N_23876,N_23618,N_23738);
xor U23877 (N_23877,N_23559,N_23515);
xor U23878 (N_23878,N_23689,N_23631);
nand U23879 (N_23879,N_23641,N_23715);
and U23880 (N_23880,N_23701,N_23576);
nor U23881 (N_23881,N_23537,N_23609);
or U23882 (N_23882,N_23614,N_23558);
nand U23883 (N_23883,N_23514,N_23645);
nor U23884 (N_23884,N_23565,N_23500);
or U23885 (N_23885,N_23516,N_23618);
nand U23886 (N_23886,N_23521,N_23636);
nand U23887 (N_23887,N_23620,N_23501);
nand U23888 (N_23888,N_23548,N_23535);
xor U23889 (N_23889,N_23625,N_23630);
and U23890 (N_23890,N_23628,N_23632);
nand U23891 (N_23891,N_23744,N_23611);
and U23892 (N_23892,N_23638,N_23523);
xnor U23893 (N_23893,N_23520,N_23709);
nor U23894 (N_23894,N_23568,N_23506);
or U23895 (N_23895,N_23630,N_23662);
nand U23896 (N_23896,N_23726,N_23590);
or U23897 (N_23897,N_23520,N_23634);
xnor U23898 (N_23898,N_23567,N_23604);
xor U23899 (N_23899,N_23551,N_23609);
nand U23900 (N_23900,N_23710,N_23624);
xor U23901 (N_23901,N_23553,N_23665);
xor U23902 (N_23902,N_23586,N_23566);
xor U23903 (N_23903,N_23748,N_23627);
or U23904 (N_23904,N_23641,N_23673);
or U23905 (N_23905,N_23748,N_23672);
or U23906 (N_23906,N_23572,N_23652);
and U23907 (N_23907,N_23577,N_23642);
nor U23908 (N_23908,N_23539,N_23650);
nand U23909 (N_23909,N_23744,N_23746);
or U23910 (N_23910,N_23703,N_23610);
xor U23911 (N_23911,N_23683,N_23584);
nand U23912 (N_23912,N_23638,N_23697);
nand U23913 (N_23913,N_23682,N_23575);
and U23914 (N_23914,N_23662,N_23573);
nand U23915 (N_23915,N_23568,N_23671);
nand U23916 (N_23916,N_23735,N_23538);
nand U23917 (N_23917,N_23624,N_23502);
xor U23918 (N_23918,N_23533,N_23541);
nor U23919 (N_23919,N_23510,N_23668);
or U23920 (N_23920,N_23705,N_23719);
xor U23921 (N_23921,N_23607,N_23696);
xor U23922 (N_23922,N_23589,N_23724);
xor U23923 (N_23923,N_23519,N_23646);
nand U23924 (N_23924,N_23592,N_23708);
nor U23925 (N_23925,N_23672,N_23699);
nand U23926 (N_23926,N_23618,N_23531);
or U23927 (N_23927,N_23721,N_23635);
nand U23928 (N_23928,N_23734,N_23500);
and U23929 (N_23929,N_23529,N_23633);
or U23930 (N_23930,N_23559,N_23547);
or U23931 (N_23931,N_23515,N_23508);
xnor U23932 (N_23932,N_23689,N_23691);
nand U23933 (N_23933,N_23677,N_23675);
nor U23934 (N_23934,N_23566,N_23729);
nor U23935 (N_23935,N_23514,N_23724);
and U23936 (N_23936,N_23742,N_23729);
or U23937 (N_23937,N_23647,N_23587);
nand U23938 (N_23938,N_23725,N_23556);
or U23939 (N_23939,N_23500,N_23611);
or U23940 (N_23940,N_23657,N_23554);
nor U23941 (N_23941,N_23527,N_23595);
nor U23942 (N_23942,N_23591,N_23609);
nand U23943 (N_23943,N_23612,N_23614);
nand U23944 (N_23944,N_23749,N_23739);
nor U23945 (N_23945,N_23682,N_23749);
and U23946 (N_23946,N_23623,N_23599);
nor U23947 (N_23947,N_23694,N_23591);
xnor U23948 (N_23948,N_23657,N_23607);
or U23949 (N_23949,N_23636,N_23643);
or U23950 (N_23950,N_23638,N_23574);
xor U23951 (N_23951,N_23573,N_23528);
or U23952 (N_23952,N_23670,N_23527);
nand U23953 (N_23953,N_23538,N_23548);
xor U23954 (N_23954,N_23579,N_23661);
nor U23955 (N_23955,N_23620,N_23645);
nor U23956 (N_23956,N_23648,N_23669);
xnor U23957 (N_23957,N_23624,N_23615);
and U23958 (N_23958,N_23683,N_23718);
or U23959 (N_23959,N_23522,N_23600);
nor U23960 (N_23960,N_23746,N_23636);
nor U23961 (N_23961,N_23707,N_23682);
nand U23962 (N_23962,N_23625,N_23599);
nor U23963 (N_23963,N_23653,N_23685);
nor U23964 (N_23964,N_23685,N_23632);
or U23965 (N_23965,N_23644,N_23692);
or U23966 (N_23966,N_23521,N_23653);
xnor U23967 (N_23967,N_23694,N_23650);
or U23968 (N_23968,N_23557,N_23692);
and U23969 (N_23969,N_23746,N_23640);
nand U23970 (N_23970,N_23685,N_23665);
nor U23971 (N_23971,N_23657,N_23518);
nor U23972 (N_23972,N_23512,N_23527);
xnor U23973 (N_23973,N_23572,N_23680);
or U23974 (N_23974,N_23710,N_23631);
xor U23975 (N_23975,N_23644,N_23619);
nand U23976 (N_23976,N_23738,N_23518);
nand U23977 (N_23977,N_23538,N_23500);
nor U23978 (N_23978,N_23719,N_23731);
nand U23979 (N_23979,N_23584,N_23700);
xor U23980 (N_23980,N_23737,N_23699);
and U23981 (N_23981,N_23620,N_23564);
and U23982 (N_23982,N_23735,N_23649);
xor U23983 (N_23983,N_23580,N_23745);
nor U23984 (N_23984,N_23699,N_23609);
nand U23985 (N_23985,N_23722,N_23737);
nand U23986 (N_23986,N_23749,N_23609);
and U23987 (N_23987,N_23581,N_23684);
and U23988 (N_23988,N_23521,N_23681);
or U23989 (N_23989,N_23616,N_23675);
and U23990 (N_23990,N_23730,N_23654);
nor U23991 (N_23991,N_23724,N_23698);
and U23992 (N_23992,N_23594,N_23580);
and U23993 (N_23993,N_23740,N_23560);
nor U23994 (N_23994,N_23599,N_23704);
and U23995 (N_23995,N_23505,N_23634);
nand U23996 (N_23996,N_23536,N_23641);
nor U23997 (N_23997,N_23548,N_23543);
and U23998 (N_23998,N_23720,N_23521);
nor U23999 (N_23999,N_23649,N_23644);
and U24000 (N_24000,N_23917,N_23775);
nand U24001 (N_24001,N_23810,N_23918);
xor U24002 (N_24002,N_23855,N_23912);
nor U24003 (N_24003,N_23943,N_23893);
nor U24004 (N_24004,N_23859,N_23803);
xnor U24005 (N_24005,N_23846,N_23920);
nor U24006 (N_24006,N_23947,N_23833);
nor U24007 (N_24007,N_23925,N_23852);
or U24008 (N_24008,N_23974,N_23930);
nor U24009 (N_24009,N_23984,N_23802);
nor U24010 (N_24010,N_23907,N_23760);
nand U24011 (N_24011,N_23877,N_23841);
and U24012 (N_24012,N_23789,N_23892);
nand U24013 (N_24013,N_23993,N_23823);
and U24014 (N_24014,N_23781,N_23985);
nand U24015 (N_24015,N_23771,N_23766);
nand U24016 (N_24016,N_23792,N_23902);
or U24017 (N_24017,N_23765,N_23929);
or U24018 (N_24018,N_23853,N_23777);
and U24019 (N_24019,N_23991,N_23934);
or U24020 (N_24020,N_23961,N_23960);
and U24021 (N_24021,N_23774,N_23849);
nor U24022 (N_24022,N_23845,N_23981);
xor U24023 (N_24023,N_23860,N_23957);
nand U24024 (N_24024,N_23913,N_23834);
xnor U24025 (N_24025,N_23868,N_23759);
or U24026 (N_24026,N_23851,N_23903);
nor U24027 (N_24027,N_23832,N_23779);
xor U24028 (N_24028,N_23905,N_23915);
nand U24029 (N_24029,N_23945,N_23768);
and U24030 (N_24030,N_23844,N_23795);
nand U24031 (N_24031,N_23786,N_23797);
xor U24032 (N_24032,N_23835,N_23872);
nor U24033 (N_24033,N_23848,N_23939);
xnor U24034 (N_24034,N_23978,N_23898);
xor U24035 (N_24035,N_23858,N_23911);
and U24036 (N_24036,N_23926,N_23773);
nor U24037 (N_24037,N_23990,N_23887);
and U24038 (N_24038,N_23935,N_23964);
or U24039 (N_24039,N_23975,N_23850);
xor U24040 (N_24040,N_23752,N_23890);
nand U24041 (N_24041,N_23980,N_23944);
xnor U24042 (N_24042,N_23989,N_23966);
or U24043 (N_24043,N_23962,N_23826);
nand U24044 (N_24044,N_23937,N_23970);
xnor U24045 (N_24045,N_23891,N_23783);
or U24046 (N_24046,N_23971,N_23817);
nand U24047 (N_24047,N_23922,N_23942);
nor U24048 (N_24048,N_23916,N_23825);
nor U24049 (N_24049,N_23987,N_23979);
or U24050 (N_24050,N_23798,N_23956);
and U24051 (N_24051,N_23908,N_23847);
nand U24052 (N_24052,N_23862,N_23914);
nor U24053 (N_24053,N_23867,N_23936);
and U24054 (N_24054,N_23818,N_23808);
nor U24055 (N_24055,N_23910,N_23959);
nor U24056 (N_24056,N_23923,N_23963);
xor U24057 (N_24057,N_23756,N_23787);
xnor U24058 (N_24058,N_23793,N_23873);
and U24059 (N_24059,N_23986,N_23900);
nand U24060 (N_24060,N_23932,N_23751);
nor U24061 (N_24061,N_23794,N_23958);
xnor U24062 (N_24062,N_23837,N_23824);
xnor U24063 (N_24063,N_23888,N_23965);
nand U24064 (N_24064,N_23763,N_23885);
nand U24065 (N_24065,N_23857,N_23805);
and U24066 (N_24066,N_23899,N_23784);
xor U24067 (N_24067,N_23820,N_23778);
nand U24068 (N_24068,N_23950,N_23982);
or U24069 (N_24069,N_23828,N_23843);
or U24070 (N_24070,N_23830,N_23968);
and U24071 (N_24071,N_23772,N_23806);
or U24072 (N_24072,N_23755,N_23791);
or U24073 (N_24073,N_23758,N_23870);
nand U24074 (N_24074,N_23938,N_23995);
nand U24075 (N_24075,N_23799,N_23941);
nor U24076 (N_24076,N_23776,N_23865);
or U24077 (N_24077,N_23953,N_23750);
and U24078 (N_24078,N_23796,N_23909);
nor U24079 (N_24079,N_23842,N_23761);
xor U24080 (N_24080,N_23901,N_23889);
xor U24081 (N_24081,N_23969,N_23822);
or U24082 (N_24082,N_23933,N_23897);
nor U24083 (N_24083,N_23764,N_23998);
xnor U24084 (N_24084,N_23973,N_23790);
xor U24085 (N_24085,N_23829,N_23866);
or U24086 (N_24086,N_23800,N_23996);
nor U24087 (N_24087,N_23886,N_23831);
or U24088 (N_24088,N_23811,N_23770);
nand U24089 (N_24089,N_23946,N_23875);
and U24090 (N_24090,N_23972,N_23785);
nand U24091 (N_24091,N_23882,N_23954);
nand U24092 (N_24092,N_23904,N_23992);
nor U24093 (N_24093,N_23921,N_23884);
nand U24094 (N_24094,N_23854,N_23864);
nand U24095 (N_24095,N_23879,N_23769);
and U24096 (N_24096,N_23827,N_23815);
xnor U24097 (N_24097,N_23839,N_23952);
nand U24098 (N_24098,N_23931,N_23955);
and U24099 (N_24099,N_23782,N_23780);
and U24100 (N_24100,N_23951,N_23988);
or U24101 (N_24101,N_23919,N_23876);
and U24102 (N_24102,N_23812,N_23753);
nor U24103 (N_24103,N_23883,N_23807);
or U24104 (N_24104,N_23874,N_23895);
nor U24105 (N_24105,N_23836,N_23809);
nand U24106 (N_24106,N_23821,N_23927);
nor U24107 (N_24107,N_23906,N_23896);
and U24108 (N_24108,N_23940,N_23928);
xnor U24109 (N_24109,N_23871,N_23948);
or U24110 (N_24110,N_23924,N_23819);
and U24111 (N_24111,N_23869,N_23983);
xnor U24112 (N_24112,N_23894,N_23994);
and U24113 (N_24113,N_23814,N_23856);
or U24114 (N_24114,N_23804,N_23967);
nor U24115 (N_24115,N_23813,N_23861);
nand U24116 (N_24116,N_23757,N_23881);
or U24117 (N_24117,N_23949,N_23762);
and U24118 (N_24118,N_23801,N_23976);
nor U24119 (N_24119,N_23880,N_23788);
nand U24120 (N_24120,N_23997,N_23999);
and U24121 (N_24121,N_23863,N_23767);
and U24122 (N_24122,N_23840,N_23816);
or U24123 (N_24123,N_23977,N_23878);
nand U24124 (N_24124,N_23838,N_23754);
or U24125 (N_24125,N_23847,N_23760);
nor U24126 (N_24126,N_23811,N_23921);
or U24127 (N_24127,N_23852,N_23781);
nand U24128 (N_24128,N_23797,N_23904);
and U24129 (N_24129,N_23889,N_23997);
nor U24130 (N_24130,N_23827,N_23912);
and U24131 (N_24131,N_23779,N_23763);
nor U24132 (N_24132,N_23817,N_23973);
nand U24133 (N_24133,N_23777,N_23964);
nor U24134 (N_24134,N_23867,N_23934);
nand U24135 (N_24135,N_23877,N_23772);
xnor U24136 (N_24136,N_23983,N_23803);
nand U24137 (N_24137,N_23991,N_23813);
nand U24138 (N_24138,N_23817,N_23952);
xnor U24139 (N_24139,N_23768,N_23993);
nor U24140 (N_24140,N_23968,N_23841);
and U24141 (N_24141,N_23877,N_23955);
nor U24142 (N_24142,N_23937,N_23948);
or U24143 (N_24143,N_23761,N_23923);
nor U24144 (N_24144,N_23924,N_23953);
nor U24145 (N_24145,N_23998,N_23914);
and U24146 (N_24146,N_23835,N_23830);
nor U24147 (N_24147,N_23921,N_23975);
nor U24148 (N_24148,N_23818,N_23983);
nand U24149 (N_24149,N_23940,N_23826);
nand U24150 (N_24150,N_23965,N_23916);
nor U24151 (N_24151,N_23760,N_23783);
nand U24152 (N_24152,N_23991,N_23772);
nor U24153 (N_24153,N_23970,N_23785);
xnor U24154 (N_24154,N_23898,N_23998);
nor U24155 (N_24155,N_23831,N_23800);
nand U24156 (N_24156,N_23982,N_23837);
or U24157 (N_24157,N_23790,N_23945);
xnor U24158 (N_24158,N_23942,N_23790);
nand U24159 (N_24159,N_23946,N_23822);
or U24160 (N_24160,N_23984,N_23797);
or U24161 (N_24161,N_23823,N_23932);
and U24162 (N_24162,N_23909,N_23989);
nand U24163 (N_24163,N_23889,N_23788);
and U24164 (N_24164,N_23925,N_23842);
xor U24165 (N_24165,N_23947,N_23910);
and U24166 (N_24166,N_23975,N_23808);
xnor U24167 (N_24167,N_23929,N_23901);
and U24168 (N_24168,N_23930,N_23808);
nand U24169 (N_24169,N_23979,N_23928);
and U24170 (N_24170,N_23829,N_23835);
or U24171 (N_24171,N_23961,N_23828);
or U24172 (N_24172,N_23942,N_23823);
nor U24173 (N_24173,N_23866,N_23991);
and U24174 (N_24174,N_23977,N_23967);
xor U24175 (N_24175,N_23893,N_23971);
nor U24176 (N_24176,N_23983,N_23856);
or U24177 (N_24177,N_23934,N_23756);
and U24178 (N_24178,N_23981,N_23799);
xor U24179 (N_24179,N_23959,N_23759);
nand U24180 (N_24180,N_23980,N_23891);
xor U24181 (N_24181,N_23910,N_23812);
or U24182 (N_24182,N_23837,N_23855);
xor U24183 (N_24183,N_23980,N_23788);
nor U24184 (N_24184,N_23912,N_23967);
or U24185 (N_24185,N_23750,N_23851);
nor U24186 (N_24186,N_23849,N_23899);
nor U24187 (N_24187,N_23872,N_23771);
xnor U24188 (N_24188,N_23825,N_23941);
or U24189 (N_24189,N_23819,N_23975);
and U24190 (N_24190,N_23831,N_23950);
and U24191 (N_24191,N_23772,N_23808);
nor U24192 (N_24192,N_23850,N_23892);
and U24193 (N_24193,N_23830,N_23753);
or U24194 (N_24194,N_23941,N_23947);
xor U24195 (N_24195,N_23967,N_23784);
and U24196 (N_24196,N_23860,N_23912);
or U24197 (N_24197,N_23784,N_23939);
nor U24198 (N_24198,N_23973,N_23977);
nor U24199 (N_24199,N_23761,N_23937);
or U24200 (N_24200,N_23823,N_23913);
nor U24201 (N_24201,N_23788,N_23886);
nor U24202 (N_24202,N_23989,N_23884);
and U24203 (N_24203,N_23755,N_23978);
and U24204 (N_24204,N_23951,N_23934);
xor U24205 (N_24205,N_23818,N_23751);
and U24206 (N_24206,N_23873,N_23782);
nand U24207 (N_24207,N_23866,N_23849);
and U24208 (N_24208,N_23978,N_23766);
and U24209 (N_24209,N_23771,N_23892);
xor U24210 (N_24210,N_23795,N_23962);
or U24211 (N_24211,N_23804,N_23875);
xor U24212 (N_24212,N_23955,N_23893);
xnor U24213 (N_24213,N_23883,N_23854);
nand U24214 (N_24214,N_23859,N_23934);
nand U24215 (N_24215,N_23866,N_23912);
nor U24216 (N_24216,N_23872,N_23751);
nand U24217 (N_24217,N_23899,N_23856);
and U24218 (N_24218,N_23856,N_23900);
nand U24219 (N_24219,N_23837,N_23817);
nor U24220 (N_24220,N_23801,N_23868);
nor U24221 (N_24221,N_23990,N_23995);
xnor U24222 (N_24222,N_23806,N_23819);
or U24223 (N_24223,N_23918,N_23758);
nor U24224 (N_24224,N_23806,N_23969);
or U24225 (N_24225,N_23927,N_23809);
or U24226 (N_24226,N_23958,N_23796);
nor U24227 (N_24227,N_23836,N_23949);
xnor U24228 (N_24228,N_23835,N_23799);
and U24229 (N_24229,N_23923,N_23949);
nor U24230 (N_24230,N_23756,N_23869);
nor U24231 (N_24231,N_23794,N_23929);
xnor U24232 (N_24232,N_23770,N_23828);
nor U24233 (N_24233,N_23794,N_23872);
xor U24234 (N_24234,N_23887,N_23756);
and U24235 (N_24235,N_23997,N_23905);
nand U24236 (N_24236,N_23984,N_23969);
nand U24237 (N_24237,N_23759,N_23985);
and U24238 (N_24238,N_23940,N_23980);
or U24239 (N_24239,N_23991,N_23905);
or U24240 (N_24240,N_23925,N_23826);
xor U24241 (N_24241,N_23773,N_23754);
xnor U24242 (N_24242,N_23777,N_23985);
nand U24243 (N_24243,N_23788,N_23976);
or U24244 (N_24244,N_23933,N_23962);
and U24245 (N_24245,N_23918,N_23966);
or U24246 (N_24246,N_23994,N_23900);
xnor U24247 (N_24247,N_23847,N_23829);
or U24248 (N_24248,N_23985,N_23888);
or U24249 (N_24249,N_23795,N_23790);
or U24250 (N_24250,N_24003,N_24218);
nand U24251 (N_24251,N_24000,N_24086);
nand U24252 (N_24252,N_24200,N_24100);
xnor U24253 (N_24253,N_24018,N_24175);
nor U24254 (N_24254,N_24079,N_24230);
nor U24255 (N_24255,N_24211,N_24249);
nand U24256 (N_24256,N_24215,N_24064);
nand U24257 (N_24257,N_24062,N_24063);
nand U24258 (N_24258,N_24007,N_24113);
and U24259 (N_24259,N_24101,N_24219);
and U24260 (N_24260,N_24024,N_24241);
nand U24261 (N_24261,N_24121,N_24157);
and U24262 (N_24262,N_24025,N_24061);
nor U24263 (N_24263,N_24149,N_24033);
xnor U24264 (N_24264,N_24123,N_24115);
nand U24265 (N_24265,N_24049,N_24232);
xnor U24266 (N_24266,N_24088,N_24132);
and U24267 (N_24267,N_24236,N_24122);
or U24268 (N_24268,N_24098,N_24070);
or U24269 (N_24269,N_24134,N_24119);
or U24270 (N_24270,N_24147,N_24233);
xor U24271 (N_24271,N_24205,N_24248);
and U24272 (N_24272,N_24028,N_24083);
and U24273 (N_24273,N_24231,N_24164);
nor U24274 (N_24274,N_24111,N_24243);
and U24275 (N_24275,N_24234,N_24103);
xnor U24276 (N_24276,N_24220,N_24131);
and U24277 (N_24277,N_24207,N_24170);
or U24278 (N_24278,N_24117,N_24019);
and U24279 (N_24279,N_24116,N_24084);
nor U24280 (N_24280,N_24209,N_24180);
xnor U24281 (N_24281,N_24161,N_24091);
nor U24282 (N_24282,N_24069,N_24060);
nor U24283 (N_24283,N_24129,N_24081);
nor U24284 (N_24284,N_24167,N_24176);
or U24285 (N_24285,N_24050,N_24102);
nand U24286 (N_24286,N_24125,N_24216);
or U24287 (N_24287,N_24139,N_24008);
nand U24288 (N_24288,N_24197,N_24108);
xor U24289 (N_24289,N_24204,N_24169);
nor U24290 (N_24290,N_24052,N_24127);
and U24291 (N_24291,N_24178,N_24151);
xor U24292 (N_24292,N_24144,N_24191);
and U24293 (N_24293,N_24206,N_24153);
and U24294 (N_24294,N_24208,N_24022);
and U24295 (N_24295,N_24030,N_24198);
nor U24296 (N_24296,N_24226,N_24174);
nand U24297 (N_24297,N_24203,N_24145);
xor U24298 (N_24298,N_24156,N_24228);
nand U24299 (N_24299,N_24173,N_24239);
nor U24300 (N_24300,N_24080,N_24212);
xnor U24301 (N_24301,N_24133,N_24192);
nand U24302 (N_24302,N_24048,N_24087);
xnor U24303 (N_24303,N_24237,N_24009);
and U24304 (N_24304,N_24155,N_24181);
or U24305 (N_24305,N_24242,N_24213);
and U24306 (N_24306,N_24128,N_24136);
nand U24307 (N_24307,N_24221,N_24214);
or U24308 (N_24308,N_24006,N_24012);
nand U24309 (N_24309,N_24097,N_24002);
xnor U24310 (N_24310,N_24029,N_24059);
and U24311 (N_24311,N_24229,N_24107);
and U24312 (N_24312,N_24001,N_24126);
and U24313 (N_24313,N_24158,N_24057);
xnor U24314 (N_24314,N_24020,N_24021);
nor U24315 (N_24315,N_24152,N_24055);
xor U24316 (N_24316,N_24053,N_24124);
nor U24317 (N_24317,N_24043,N_24046);
xor U24318 (N_24318,N_24160,N_24166);
xnor U24319 (N_24319,N_24013,N_24159);
or U24320 (N_24320,N_24227,N_24068);
or U24321 (N_24321,N_24168,N_24118);
nor U24322 (N_24322,N_24142,N_24224);
xor U24323 (N_24323,N_24032,N_24141);
nand U24324 (N_24324,N_24225,N_24105);
xor U24325 (N_24325,N_24195,N_24040);
nor U24326 (N_24326,N_24073,N_24165);
xor U24327 (N_24327,N_24172,N_24035);
nand U24328 (N_24328,N_24065,N_24184);
nand U24329 (N_24329,N_24005,N_24016);
or U24330 (N_24330,N_24189,N_24036);
nand U24331 (N_24331,N_24041,N_24201);
xnor U24332 (N_24332,N_24187,N_24182);
or U24333 (N_24333,N_24199,N_24137);
and U24334 (N_24334,N_24183,N_24077);
and U24335 (N_24335,N_24039,N_24120);
xnor U24336 (N_24336,N_24140,N_24202);
or U24337 (N_24337,N_24054,N_24114);
or U24338 (N_24338,N_24190,N_24096);
nor U24339 (N_24339,N_24162,N_24004);
or U24340 (N_24340,N_24092,N_24179);
xor U24341 (N_24341,N_24094,N_24067);
or U24342 (N_24342,N_24240,N_24130);
nor U24343 (N_24343,N_24217,N_24010);
or U24344 (N_24344,N_24047,N_24148);
nor U24345 (N_24345,N_24247,N_24223);
and U24346 (N_24346,N_24109,N_24194);
nor U24347 (N_24347,N_24196,N_24154);
nor U24348 (N_24348,N_24074,N_24076);
nor U24349 (N_24349,N_24163,N_24186);
xor U24350 (N_24350,N_24246,N_24056);
nor U24351 (N_24351,N_24095,N_24066);
xor U24352 (N_24352,N_24037,N_24222);
or U24353 (N_24353,N_24210,N_24089);
nor U24354 (N_24354,N_24017,N_24245);
or U24355 (N_24355,N_24171,N_24090);
nor U24356 (N_24356,N_24026,N_24072);
xnor U24357 (N_24357,N_24244,N_24031);
or U24358 (N_24358,N_24099,N_24150);
nand U24359 (N_24359,N_24071,N_24075);
and U24360 (N_24360,N_24038,N_24106);
nor U24361 (N_24361,N_24104,N_24177);
nand U24362 (N_24362,N_24044,N_24085);
or U24363 (N_24363,N_24093,N_24188);
nor U24364 (N_24364,N_24193,N_24135);
xor U24365 (N_24365,N_24143,N_24042);
xnor U24366 (N_24366,N_24011,N_24082);
and U24367 (N_24367,N_24238,N_24015);
xor U24368 (N_24368,N_24058,N_24027);
nand U24369 (N_24369,N_24014,N_24138);
nand U24370 (N_24370,N_24045,N_24235);
and U24371 (N_24371,N_24185,N_24034);
or U24372 (N_24372,N_24078,N_24146);
or U24373 (N_24373,N_24110,N_24112);
and U24374 (N_24374,N_24051,N_24023);
nor U24375 (N_24375,N_24213,N_24184);
nor U24376 (N_24376,N_24083,N_24248);
or U24377 (N_24377,N_24109,N_24026);
or U24378 (N_24378,N_24182,N_24035);
and U24379 (N_24379,N_24144,N_24230);
or U24380 (N_24380,N_24152,N_24036);
or U24381 (N_24381,N_24050,N_24164);
nand U24382 (N_24382,N_24200,N_24180);
and U24383 (N_24383,N_24231,N_24144);
nor U24384 (N_24384,N_24076,N_24155);
and U24385 (N_24385,N_24061,N_24089);
nor U24386 (N_24386,N_24077,N_24163);
nand U24387 (N_24387,N_24036,N_24000);
or U24388 (N_24388,N_24186,N_24234);
xor U24389 (N_24389,N_24149,N_24163);
or U24390 (N_24390,N_24155,N_24196);
xnor U24391 (N_24391,N_24055,N_24141);
and U24392 (N_24392,N_24061,N_24207);
nor U24393 (N_24393,N_24129,N_24037);
nor U24394 (N_24394,N_24132,N_24044);
nor U24395 (N_24395,N_24030,N_24077);
or U24396 (N_24396,N_24057,N_24039);
or U24397 (N_24397,N_24245,N_24217);
nor U24398 (N_24398,N_24039,N_24166);
and U24399 (N_24399,N_24181,N_24004);
or U24400 (N_24400,N_24182,N_24216);
and U24401 (N_24401,N_24193,N_24126);
and U24402 (N_24402,N_24094,N_24114);
or U24403 (N_24403,N_24237,N_24032);
nor U24404 (N_24404,N_24110,N_24186);
and U24405 (N_24405,N_24242,N_24151);
or U24406 (N_24406,N_24236,N_24148);
or U24407 (N_24407,N_24206,N_24055);
or U24408 (N_24408,N_24216,N_24091);
nand U24409 (N_24409,N_24197,N_24017);
or U24410 (N_24410,N_24068,N_24007);
and U24411 (N_24411,N_24139,N_24186);
xnor U24412 (N_24412,N_24011,N_24092);
or U24413 (N_24413,N_24215,N_24139);
xor U24414 (N_24414,N_24224,N_24050);
or U24415 (N_24415,N_24079,N_24012);
nor U24416 (N_24416,N_24030,N_24039);
nor U24417 (N_24417,N_24143,N_24156);
xor U24418 (N_24418,N_24057,N_24070);
xnor U24419 (N_24419,N_24045,N_24091);
nand U24420 (N_24420,N_24127,N_24020);
nand U24421 (N_24421,N_24244,N_24056);
and U24422 (N_24422,N_24166,N_24075);
and U24423 (N_24423,N_24014,N_24033);
and U24424 (N_24424,N_24114,N_24142);
xnor U24425 (N_24425,N_24007,N_24221);
xnor U24426 (N_24426,N_24001,N_24035);
xor U24427 (N_24427,N_24100,N_24056);
xnor U24428 (N_24428,N_24031,N_24065);
nand U24429 (N_24429,N_24183,N_24221);
and U24430 (N_24430,N_24175,N_24028);
nor U24431 (N_24431,N_24208,N_24153);
xnor U24432 (N_24432,N_24235,N_24108);
nand U24433 (N_24433,N_24232,N_24149);
xor U24434 (N_24434,N_24050,N_24129);
xnor U24435 (N_24435,N_24042,N_24167);
or U24436 (N_24436,N_24022,N_24075);
and U24437 (N_24437,N_24131,N_24177);
or U24438 (N_24438,N_24059,N_24205);
nor U24439 (N_24439,N_24071,N_24100);
nand U24440 (N_24440,N_24169,N_24085);
or U24441 (N_24441,N_24037,N_24068);
nand U24442 (N_24442,N_24138,N_24166);
nor U24443 (N_24443,N_24028,N_24089);
xnor U24444 (N_24444,N_24114,N_24246);
nor U24445 (N_24445,N_24076,N_24087);
xor U24446 (N_24446,N_24072,N_24148);
xor U24447 (N_24447,N_24208,N_24231);
and U24448 (N_24448,N_24040,N_24019);
or U24449 (N_24449,N_24060,N_24233);
and U24450 (N_24450,N_24214,N_24154);
nor U24451 (N_24451,N_24074,N_24036);
and U24452 (N_24452,N_24008,N_24169);
or U24453 (N_24453,N_24107,N_24223);
xor U24454 (N_24454,N_24040,N_24113);
and U24455 (N_24455,N_24201,N_24106);
nor U24456 (N_24456,N_24144,N_24093);
xor U24457 (N_24457,N_24048,N_24156);
nand U24458 (N_24458,N_24213,N_24010);
xnor U24459 (N_24459,N_24028,N_24112);
nand U24460 (N_24460,N_24200,N_24058);
and U24461 (N_24461,N_24163,N_24207);
or U24462 (N_24462,N_24192,N_24221);
or U24463 (N_24463,N_24238,N_24065);
and U24464 (N_24464,N_24240,N_24196);
xnor U24465 (N_24465,N_24093,N_24205);
xnor U24466 (N_24466,N_24152,N_24068);
and U24467 (N_24467,N_24091,N_24165);
xor U24468 (N_24468,N_24192,N_24082);
nand U24469 (N_24469,N_24085,N_24017);
nand U24470 (N_24470,N_24162,N_24200);
and U24471 (N_24471,N_24154,N_24090);
or U24472 (N_24472,N_24066,N_24004);
nor U24473 (N_24473,N_24229,N_24002);
xor U24474 (N_24474,N_24119,N_24237);
xnor U24475 (N_24475,N_24065,N_24193);
or U24476 (N_24476,N_24053,N_24138);
or U24477 (N_24477,N_24027,N_24135);
nor U24478 (N_24478,N_24243,N_24225);
xor U24479 (N_24479,N_24121,N_24088);
xor U24480 (N_24480,N_24113,N_24183);
xor U24481 (N_24481,N_24171,N_24188);
xor U24482 (N_24482,N_24179,N_24194);
xor U24483 (N_24483,N_24225,N_24127);
xor U24484 (N_24484,N_24228,N_24024);
nor U24485 (N_24485,N_24231,N_24131);
nand U24486 (N_24486,N_24080,N_24170);
nand U24487 (N_24487,N_24036,N_24196);
nand U24488 (N_24488,N_24130,N_24203);
nand U24489 (N_24489,N_24119,N_24100);
xor U24490 (N_24490,N_24000,N_24182);
or U24491 (N_24491,N_24149,N_24059);
xnor U24492 (N_24492,N_24178,N_24041);
or U24493 (N_24493,N_24066,N_24110);
and U24494 (N_24494,N_24237,N_24019);
nand U24495 (N_24495,N_24055,N_24065);
and U24496 (N_24496,N_24029,N_24145);
or U24497 (N_24497,N_24047,N_24193);
or U24498 (N_24498,N_24070,N_24181);
nand U24499 (N_24499,N_24059,N_24148);
nand U24500 (N_24500,N_24411,N_24414);
and U24501 (N_24501,N_24291,N_24379);
or U24502 (N_24502,N_24283,N_24285);
nor U24503 (N_24503,N_24482,N_24415);
or U24504 (N_24504,N_24355,N_24276);
xnor U24505 (N_24505,N_24401,N_24445);
and U24506 (N_24506,N_24461,N_24406);
xnor U24507 (N_24507,N_24363,N_24494);
nor U24508 (N_24508,N_24436,N_24441);
xor U24509 (N_24509,N_24358,N_24469);
or U24510 (N_24510,N_24396,N_24498);
nor U24511 (N_24511,N_24356,N_24299);
nand U24512 (N_24512,N_24274,N_24269);
xor U24513 (N_24513,N_24470,N_24349);
or U24514 (N_24514,N_24280,N_24279);
nand U24515 (N_24515,N_24474,N_24380);
nand U24516 (N_24516,N_24298,N_24359);
or U24517 (N_24517,N_24386,N_24362);
nand U24518 (N_24518,N_24389,N_24427);
nor U24519 (N_24519,N_24378,N_24265);
xnor U24520 (N_24520,N_24278,N_24457);
and U24521 (N_24521,N_24388,N_24263);
nand U24522 (N_24522,N_24485,N_24486);
and U24523 (N_24523,N_24403,N_24431);
or U24524 (N_24524,N_24323,N_24348);
nand U24525 (N_24525,N_24442,N_24476);
and U24526 (N_24526,N_24357,N_24400);
and U24527 (N_24527,N_24277,N_24337);
or U24528 (N_24528,N_24463,N_24250);
nor U24529 (N_24529,N_24271,N_24308);
nand U24530 (N_24530,N_24360,N_24381);
nor U24531 (N_24531,N_24484,N_24303);
nand U24532 (N_24532,N_24350,N_24292);
and U24533 (N_24533,N_24423,N_24275);
nand U24534 (N_24534,N_24254,N_24439);
xnor U24535 (N_24535,N_24446,N_24343);
nand U24536 (N_24536,N_24438,N_24493);
xor U24537 (N_24537,N_24429,N_24432);
nand U24538 (N_24538,N_24377,N_24306);
nor U24539 (N_24539,N_24252,N_24453);
and U24540 (N_24540,N_24335,N_24339);
nor U24541 (N_24541,N_24405,N_24284);
nor U24542 (N_24542,N_24328,N_24322);
nand U24543 (N_24543,N_24309,N_24253);
or U24544 (N_24544,N_24426,N_24404);
nor U24545 (N_24545,N_24365,N_24327);
or U24546 (N_24546,N_24496,N_24273);
nand U24547 (N_24547,N_24394,N_24490);
nand U24548 (N_24548,N_24384,N_24326);
and U24549 (N_24549,N_24440,N_24304);
nand U24550 (N_24550,N_24251,N_24383);
or U24551 (N_24551,N_24324,N_24458);
nor U24552 (N_24552,N_24397,N_24402);
nor U24553 (N_24553,N_24311,N_24325);
xor U24554 (N_24554,N_24419,N_24302);
nor U24555 (N_24555,N_24422,N_24434);
and U24556 (N_24556,N_24368,N_24312);
xnor U24557 (N_24557,N_24366,N_24424);
and U24558 (N_24558,N_24336,N_24407);
xnor U24559 (N_24559,N_24315,N_24433);
or U24560 (N_24560,N_24468,N_24459);
nor U24561 (N_24561,N_24499,N_24479);
and U24562 (N_24562,N_24385,N_24286);
and U24563 (N_24563,N_24370,N_24449);
nor U24564 (N_24564,N_24492,N_24314);
or U24565 (N_24565,N_24487,N_24342);
or U24566 (N_24566,N_24294,N_24451);
or U24567 (N_24567,N_24488,N_24387);
and U24568 (N_24568,N_24320,N_24465);
and U24569 (N_24569,N_24460,N_24382);
or U24570 (N_24570,N_24354,N_24412);
nor U24571 (N_24571,N_24256,N_24310);
xor U24572 (N_24572,N_24437,N_24443);
nand U24573 (N_24573,N_24420,N_24466);
nor U24574 (N_24574,N_24416,N_24464);
nor U24575 (N_24575,N_24307,N_24361);
and U24576 (N_24576,N_24425,N_24471);
nor U24577 (N_24577,N_24255,N_24421);
nor U24578 (N_24578,N_24301,N_24448);
nand U24579 (N_24579,N_24316,N_24317);
xor U24580 (N_24580,N_24266,N_24353);
nor U24581 (N_24581,N_24371,N_24462);
nor U24582 (N_24582,N_24417,N_24296);
and U24583 (N_24583,N_24364,N_24418);
nand U24584 (N_24584,N_24341,N_24305);
nand U24585 (N_24585,N_24376,N_24295);
or U24586 (N_24586,N_24321,N_24467);
xnor U24587 (N_24587,N_24264,N_24345);
nand U24588 (N_24588,N_24456,N_24331);
nand U24589 (N_24589,N_24447,N_24290);
nor U24590 (N_24590,N_24413,N_24289);
nor U24591 (N_24591,N_24347,N_24393);
nand U24592 (N_24592,N_24344,N_24287);
and U24593 (N_24593,N_24390,N_24282);
nor U24594 (N_24594,N_24473,N_24257);
and U24595 (N_24595,N_24259,N_24332);
xnor U24596 (N_24596,N_24351,N_24497);
xnor U24597 (N_24597,N_24340,N_24293);
or U24598 (N_24598,N_24338,N_24270);
xnor U24599 (N_24599,N_24261,N_24267);
or U24600 (N_24600,N_24435,N_24330);
or U24601 (N_24601,N_24333,N_24281);
and U24602 (N_24602,N_24409,N_24334);
or U24603 (N_24603,N_24408,N_24483);
or U24604 (N_24604,N_24319,N_24297);
nand U24605 (N_24605,N_24430,N_24472);
and U24606 (N_24606,N_24374,N_24367);
nand U24607 (N_24607,N_24489,N_24477);
nor U24608 (N_24608,N_24478,N_24313);
nand U24609 (N_24609,N_24392,N_24455);
nor U24610 (N_24610,N_24268,N_24262);
or U24611 (N_24611,N_24352,N_24318);
nand U24612 (N_24612,N_24375,N_24300);
nand U24613 (N_24613,N_24329,N_24475);
xnor U24614 (N_24614,N_24258,N_24452);
nand U24615 (N_24615,N_24480,N_24399);
xor U24616 (N_24616,N_24481,N_24395);
nor U24617 (N_24617,N_24288,N_24391);
nand U24618 (N_24618,N_24491,N_24369);
nor U24619 (N_24619,N_24410,N_24428);
nor U24620 (N_24620,N_24454,N_24346);
and U24621 (N_24621,N_24444,N_24398);
or U24622 (N_24622,N_24450,N_24495);
nand U24623 (N_24623,N_24373,N_24272);
or U24624 (N_24624,N_24260,N_24372);
or U24625 (N_24625,N_24407,N_24419);
nand U24626 (N_24626,N_24450,N_24496);
nor U24627 (N_24627,N_24314,N_24391);
and U24628 (N_24628,N_24437,N_24274);
nor U24629 (N_24629,N_24399,N_24295);
and U24630 (N_24630,N_24294,N_24470);
or U24631 (N_24631,N_24442,N_24369);
xnor U24632 (N_24632,N_24267,N_24462);
or U24633 (N_24633,N_24497,N_24454);
nor U24634 (N_24634,N_24398,N_24414);
or U24635 (N_24635,N_24380,N_24363);
and U24636 (N_24636,N_24377,N_24477);
nor U24637 (N_24637,N_24284,N_24368);
nand U24638 (N_24638,N_24437,N_24350);
xnor U24639 (N_24639,N_24326,N_24473);
nor U24640 (N_24640,N_24426,N_24391);
and U24641 (N_24641,N_24250,N_24441);
nor U24642 (N_24642,N_24354,N_24480);
nand U24643 (N_24643,N_24484,N_24458);
xor U24644 (N_24644,N_24303,N_24362);
nor U24645 (N_24645,N_24344,N_24376);
nand U24646 (N_24646,N_24315,N_24392);
and U24647 (N_24647,N_24339,N_24322);
or U24648 (N_24648,N_24393,N_24304);
nand U24649 (N_24649,N_24356,N_24488);
and U24650 (N_24650,N_24434,N_24274);
or U24651 (N_24651,N_24337,N_24418);
and U24652 (N_24652,N_24469,N_24404);
xor U24653 (N_24653,N_24469,N_24461);
nor U24654 (N_24654,N_24256,N_24332);
or U24655 (N_24655,N_24298,N_24312);
xor U24656 (N_24656,N_24393,N_24419);
or U24657 (N_24657,N_24492,N_24471);
nor U24658 (N_24658,N_24388,N_24280);
and U24659 (N_24659,N_24492,N_24265);
nand U24660 (N_24660,N_24393,N_24313);
nor U24661 (N_24661,N_24267,N_24419);
xor U24662 (N_24662,N_24418,N_24357);
nor U24663 (N_24663,N_24495,N_24443);
or U24664 (N_24664,N_24359,N_24339);
or U24665 (N_24665,N_24423,N_24340);
or U24666 (N_24666,N_24262,N_24395);
nand U24667 (N_24667,N_24322,N_24336);
nand U24668 (N_24668,N_24327,N_24443);
nand U24669 (N_24669,N_24262,N_24398);
xnor U24670 (N_24670,N_24350,N_24287);
or U24671 (N_24671,N_24397,N_24327);
or U24672 (N_24672,N_24337,N_24268);
or U24673 (N_24673,N_24258,N_24298);
and U24674 (N_24674,N_24475,N_24399);
xor U24675 (N_24675,N_24343,N_24325);
or U24676 (N_24676,N_24495,N_24380);
nand U24677 (N_24677,N_24313,N_24285);
and U24678 (N_24678,N_24432,N_24260);
nand U24679 (N_24679,N_24305,N_24421);
xor U24680 (N_24680,N_24322,N_24352);
or U24681 (N_24681,N_24317,N_24437);
nand U24682 (N_24682,N_24375,N_24341);
and U24683 (N_24683,N_24484,N_24302);
xnor U24684 (N_24684,N_24483,N_24347);
nor U24685 (N_24685,N_24378,N_24371);
or U24686 (N_24686,N_24355,N_24282);
nor U24687 (N_24687,N_24446,N_24270);
xor U24688 (N_24688,N_24352,N_24347);
or U24689 (N_24689,N_24384,N_24295);
xnor U24690 (N_24690,N_24455,N_24433);
or U24691 (N_24691,N_24455,N_24356);
and U24692 (N_24692,N_24264,N_24252);
or U24693 (N_24693,N_24405,N_24379);
and U24694 (N_24694,N_24322,N_24378);
and U24695 (N_24695,N_24471,N_24436);
and U24696 (N_24696,N_24371,N_24271);
nand U24697 (N_24697,N_24400,N_24331);
nor U24698 (N_24698,N_24445,N_24388);
and U24699 (N_24699,N_24291,N_24489);
and U24700 (N_24700,N_24401,N_24471);
xor U24701 (N_24701,N_24342,N_24385);
nand U24702 (N_24702,N_24378,N_24498);
xor U24703 (N_24703,N_24272,N_24469);
xnor U24704 (N_24704,N_24338,N_24425);
or U24705 (N_24705,N_24420,N_24287);
nand U24706 (N_24706,N_24487,N_24307);
xor U24707 (N_24707,N_24448,N_24495);
xor U24708 (N_24708,N_24333,N_24291);
or U24709 (N_24709,N_24251,N_24469);
nor U24710 (N_24710,N_24257,N_24259);
nor U24711 (N_24711,N_24448,N_24482);
xor U24712 (N_24712,N_24347,N_24388);
and U24713 (N_24713,N_24302,N_24442);
nor U24714 (N_24714,N_24333,N_24413);
and U24715 (N_24715,N_24390,N_24472);
xor U24716 (N_24716,N_24347,N_24422);
and U24717 (N_24717,N_24308,N_24330);
nor U24718 (N_24718,N_24327,N_24252);
nand U24719 (N_24719,N_24373,N_24477);
xnor U24720 (N_24720,N_24324,N_24432);
xnor U24721 (N_24721,N_24341,N_24329);
and U24722 (N_24722,N_24354,N_24469);
xnor U24723 (N_24723,N_24264,N_24316);
nor U24724 (N_24724,N_24329,N_24494);
nor U24725 (N_24725,N_24378,N_24454);
nor U24726 (N_24726,N_24375,N_24274);
or U24727 (N_24727,N_24473,N_24422);
nor U24728 (N_24728,N_24442,N_24398);
or U24729 (N_24729,N_24324,N_24272);
and U24730 (N_24730,N_24293,N_24405);
xnor U24731 (N_24731,N_24412,N_24355);
or U24732 (N_24732,N_24323,N_24497);
nand U24733 (N_24733,N_24495,N_24447);
or U24734 (N_24734,N_24457,N_24439);
or U24735 (N_24735,N_24323,N_24333);
nand U24736 (N_24736,N_24351,N_24329);
and U24737 (N_24737,N_24340,N_24413);
nor U24738 (N_24738,N_24483,N_24495);
nand U24739 (N_24739,N_24396,N_24383);
xor U24740 (N_24740,N_24478,N_24446);
nor U24741 (N_24741,N_24478,N_24345);
xor U24742 (N_24742,N_24385,N_24489);
and U24743 (N_24743,N_24361,N_24407);
or U24744 (N_24744,N_24431,N_24469);
or U24745 (N_24745,N_24441,N_24292);
xor U24746 (N_24746,N_24259,N_24364);
xnor U24747 (N_24747,N_24444,N_24356);
xor U24748 (N_24748,N_24314,N_24446);
or U24749 (N_24749,N_24473,N_24301);
nand U24750 (N_24750,N_24544,N_24632);
nor U24751 (N_24751,N_24526,N_24642);
nand U24752 (N_24752,N_24576,N_24725);
nand U24753 (N_24753,N_24540,N_24686);
or U24754 (N_24754,N_24638,N_24527);
or U24755 (N_24755,N_24690,N_24665);
and U24756 (N_24756,N_24649,N_24625);
and U24757 (N_24757,N_24730,N_24747);
or U24758 (N_24758,N_24663,N_24709);
xor U24759 (N_24759,N_24640,N_24685);
xor U24760 (N_24760,N_24566,N_24716);
and U24761 (N_24761,N_24683,N_24697);
or U24762 (N_24762,N_24541,N_24729);
nor U24763 (N_24763,N_24557,N_24620);
or U24764 (N_24764,N_24538,N_24517);
and U24765 (N_24765,N_24512,N_24609);
nand U24766 (N_24766,N_24562,N_24667);
xor U24767 (N_24767,N_24728,N_24732);
xnor U24768 (N_24768,N_24570,N_24536);
and U24769 (N_24769,N_24706,N_24639);
xnor U24770 (N_24770,N_24584,N_24623);
nor U24771 (N_24771,N_24513,N_24585);
nor U24772 (N_24772,N_24553,N_24572);
nor U24773 (N_24773,N_24741,N_24646);
nand U24774 (N_24774,N_24662,N_24519);
nor U24775 (N_24775,N_24508,N_24565);
nand U24776 (N_24776,N_24731,N_24657);
xnor U24777 (N_24777,N_24594,N_24645);
xor U24778 (N_24778,N_24677,N_24534);
or U24779 (N_24779,N_24539,N_24637);
xor U24780 (N_24780,N_24511,N_24647);
nand U24781 (N_24781,N_24571,N_24717);
nor U24782 (N_24782,N_24669,N_24722);
and U24783 (N_24783,N_24636,N_24727);
or U24784 (N_24784,N_24676,N_24695);
and U24785 (N_24785,N_24664,N_24693);
and U24786 (N_24786,N_24615,N_24740);
or U24787 (N_24787,N_24605,N_24506);
nand U24788 (N_24788,N_24711,N_24533);
nand U24789 (N_24789,N_24656,N_24633);
or U24790 (N_24790,N_24688,N_24713);
xnor U24791 (N_24791,N_24653,N_24558);
nor U24792 (N_24792,N_24680,N_24612);
xor U24793 (N_24793,N_24682,N_24660);
or U24794 (N_24794,N_24520,N_24654);
or U24795 (N_24795,N_24661,N_24575);
or U24796 (N_24796,N_24611,N_24525);
and U24797 (N_24797,N_24503,N_24554);
xor U24798 (N_24798,N_24710,N_24581);
or U24799 (N_24799,N_24604,N_24691);
and U24800 (N_24800,N_24616,N_24749);
and U24801 (N_24801,N_24687,N_24715);
nor U24802 (N_24802,N_24546,N_24628);
or U24803 (N_24803,N_24744,N_24641);
nor U24804 (N_24804,N_24668,N_24543);
xnor U24805 (N_24805,N_24704,N_24535);
or U24806 (N_24806,N_24681,N_24733);
nand U24807 (N_24807,N_24745,N_24505);
and U24808 (N_24808,N_24521,N_24726);
nor U24809 (N_24809,N_24537,N_24679);
nand U24810 (N_24810,N_24718,N_24607);
nand U24811 (N_24811,N_24591,N_24569);
nand U24812 (N_24812,N_24593,N_24696);
or U24813 (N_24813,N_24651,N_24689);
or U24814 (N_24814,N_24705,N_24626);
or U24815 (N_24815,N_24671,N_24721);
and U24816 (N_24816,N_24698,N_24719);
or U24817 (N_24817,N_24714,N_24587);
and U24818 (N_24818,N_24550,N_24617);
xor U24819 (N_24819,N_24724,N_24723);
nor U24820 (N_24820,N_24630,N_24600);
or U24821 (N_24821,N_24518,N_24573);
nor U24822 (N_24822,N_24528,N_24545);
xor U24823 (N_24823,N_24603,N_24507);
and U24824 (N_24824,N_24748,N_24595);
nand U24825 (N_24825,N_24532,N_24580);
and U24826 (N_24826,N_24684,N_24670);
nand U24827 (N_24827,N_24501,N_24516);
nor U24828 (N_24828,N_24598,N_24524);
xnor U24829 (N_24829,N_24700,N_24602);
and U24830 (N_24830,N_24699,N_24586);
and U24831 (N_24831,N_24694,N_24629);
xnor U24832 (N_24832,N_24658,N_24561);
or U24833 (N_24833,N_24555,N_24502);
nor U24834 (N_24834,N_24627,N_24522);
and U24835 (N_24835,N_24552,N_24601);
nor U24836 (N_24836,N_24675,N_24592);
nand U24837 (N_24837,N_24589,N_24606);
or U24838 (N_24838,N_24578,N_24734);
and U24839 (N_24839,N_24579,N_24622);
xor U24840 (N_24840,N_24510,N_24701);
nor U24841 (N_24841,N_24652,N_24547);
nand U24842 (N_24842,N_24597,N_24530);
nor U24843 (N_24843,N_24631,N_24703);
or U24844 (N_24844,N_24738,N_24549);
or U24845 (N_24845,N_24500,N_24574);
and U24846 (N_24846,N_24596,N_24610);
or U24847 (N_24847,N_24659,N_24736);
nor U24848 (N_24848,N_24514,N_24735);
xor U24849 (N_24849,N_24583,N_24621);
or U24850 (N_24850,N_24608,N_24582);
xor U24851 (N_24851,N_24613,N_24542);
nor U24852 (N_24852,N_24563,N_24634);
xor U24853 (N_24853,N_24666,N_24531);
nor U24854 (N_24854,N_24515,N_24504);
or U24855 (N_24855,N_24712,N_24559);
and U24856 (N_24856,N_24567,N_24692);
nor U24857 (N_24857,N_24577,N_24548);
xor U24858 (N_24858,N_24564,N_24707);
xnor U24859 (N_24859,N_24648,N_24529);
xnor U24860 (N_24860,N_24590,N_24737);
or U24861 (N_24861,N_24708,N_24673);
and U24862 (N_24862,N_24509,N_24739);
and U24863 (N_24863,N_24618,N_24655);
nor U24864 (N_24864,N_24624,N_24614);
and U24865 (N_24865,N_24588,N_24560);
nor U24866 (N_24866,N_24644,N_24743);
and U24867 (N_24867,N_24619,N_24672);
or U24868 (N_24868,N_24674,N_24720);
xor U24869 (N_24869,N_24746,N_24643);
and U24870 (N_24870,N_24523,N_24678);
and U24871 (N_24871,N_24702,N_24742);
or U24872 (N_24872,N_24635,N_24551);
and U24873 (N_24873,N_24556,N_24568);
nand U24874 (N_24874,N_24650,N_24599);
or U24875 (N_24875,N_24599,N_24588);
nand U24876 (N_24876,N_24636,N_24681);
nor U24877 (N_24877,N_24717,N_24661);
or U24878 (N_24878,N_24731,N_24713);
or U24879 (N_24879,N_24716,N_24562);
xnor U24880 (N_24880,N_24519,N_24625);
xor U24881 (N_24881,N_24634,N_24684);
or U24882 (N_24882,N_24554,N_24749);
nor U24883 (N_24883,N_24692,N_24503);
nor U24884 (N_24884,N_24603,N_24644);
or U24885 (N_24885,N_24654,N_24559);
or U24886 (N_24886,N_24607,N_24561);
nand U24887 (N_24887,N_24659,N_24528);
nand U24888 (N_24888,N_24702,N_24578);
nand U24889 (N_24889,N_24525,N_24507);
nand U24890 (N_24890,N_24666,N_24709);
nor U24891 (N_24891,N_24739,N_24607);
xnor U24892 (N_24892,N_24519,N_24618);
xor U24893 (N_24893,N_24665,N_24575);
xor U24894 (N_24894,N_24588,N_24655);
nor U24895 (N_24895,N_24619,N_24657);
nand U24896 (N_24896,N_24745,N_24667);
xor U24897 (N_24897,N_24640,N_24696);
xnor U24898 (N_24898,N_24571,N_24560);
or U24899 (N_24899,N_24738,N_24574);
or U24900 (N_24900,N_24693,N_24623);
nor U24901 (N_24901,N_24672,N_24599);
xnor U24902 (N_24902,N_24570,N_24669);
or U24903 (N_24903,N_24537,N_24741);
xor U24904 (N_24904,N_24562,N_24647);
nand U24905 (N_24905,N_24662,N_24511);
and U24906 (N_24906,N_24669,N_24658);
and U24907 (N_24907,N_24648,N_24708);
nand U24908 (N_24908,N_24743,N_24708);
or U24909 (N_24909,N_24540,N_24735);
nand U24910 (N_24910,N_24614,N_24643);
nor U24911 (N_24911,N_24664,N_24571);
or U24912 (N_24912,N_24734,N_24709);
nand U24913 (N_24913,N_24557,N_24662);
and U24914 (N_24914,N_24613,N_24603);
or U24915 (N_24915,N_24515,N_24552);
nor U24916 (N_24916,N_24696,N_24660);
nor U24917 (N_24917,N_24720,N_24550);
or U24918 (N_24918,N_24749,N_24544);
xor U24919 (N_24919,N_24713,N_24700);
or U24920 (N_24920,N_24682,N_24573);
xnor U24921 (N_24921,N_24621,N_24522);
xnor U24922 (N_24922,N_24624,N_24740);
and U24923 (N_24923,N_24596,N_24535);
xor U24924 (N_24924,N_24594,N_24619);
and U24925 (N_24925,N_24708,N_24711);
nand U24926 (N_24926,N_24542,N_24749);
or U24927 (N_24927,N_24629,N_24701);
nor U24928 (N_24928,N_24558,N_24518);
nand U24929 (N_24929,N_24709,N_24501);
nor U24930 (N_24930,N_24690,N_24615);
and U24931 (N_24931,N_24611,N_24737);
nand U24932 (N_24932,N_24586,N_24682);
xor U24933 (N_24933,N_24559,N_24683);
nand U24934 (N_24934,N_24742,N_24708);
and U24935 (N_24935,N_24705,N_24509);
xnor U24936 (N_24936,N_24745,N_24734);
nand U24937 (N_24937,N_24651,N_24509);
nand U24938 (N_24938,N_24623,N_24512);
nand U24939 (N_24939,N_24565,N_24654);
nor U24940 (N_24940,N_24501,N_24605);
and U24941 (N_24941,N_24727,N_24719);
xnor U24942 (N_24942,N_24533,N_24568);
and U24943 (N_24943,N_24650,N_24707);
and U24944 (N_24944,N_24700,N_24723);
nand U24945 (N_24945,N_24749,N_24507);
nor U24946 (N_24946,N_24668,N_24695);
and U24947 (N_24947,N_24552,N_24537);
and U24948 (N_24948,N_24687,N_24671);
xnor U24949 (N_24949,N_24600,N_24606);
and U24950 (N_24950,N_24524,N_24618);
xor U24951 (N_24951,N_24707,N_24699);
xor U24952 (N_24952,N_24737,N_24582);
nor U24953 (N_24953,N_24569,N_24749);
xor U24954 (N_24954,N_24734,N_24637);
nand U24955 (N_24955,N_24651,N_24599);
nand U24956 (N_24956,N_24618,N_24573);
nand U24957 (N_24957,N_24551,N_24652);
or U24958 (N_24958,N_24676,N_24714);
nor U24959 (N_24959,N_24589,N_24576);
xnor U24960 (N_24960,N_24620,N_24748);
xnor U24961 (N_24961,N_24691,N_24606);
nand U24962 (N_24962,N_24510,N_24692);
nor U24963 (N_24963,N_24505,N_24726);
or U24964 (N_24964,N_24578,N_24673);
or U24965 (N_24965,N_24555,N_24582);
xor U24966 (N_24966,N_24734,N_24659);
or U24967 (N_24967,N_24546,N_24648);
nor U24968 (N_24968,N_24648,N_24558);
or U24969 (N_24969,N_24679,N_24510);
nor U24970 (N_24970,N_24738,N_24512);
nand U24971 (N_24971,N_24665,N_24536);
nor U24972 (N_24972,N_24505,N_24706);
xor U24973 (N_24973,N_24530,N_24587);
and U24974 (N_24974,N_24574,N_24513);
and U24975 (N_24975,N_24651,N_24536);
nand U24976 (N_24976,N_24558,N_24658);
and U24977 (N_24977,N_24740,N_24747);
or U24978 (N_24978,N_24638,N_24561);
nand U24979 (N_24979,N_24660,N_24661);
or U24980 (N_24980,N_24530,N_24675);
nor U24981 (N_24981,N_24613,N_24632);
and U24982 (N_24982,N_24577,N_24511);
nand U24983 (N_24983,N_24540,N_24601);
and U24984 (N_24984,N_24514,N_24578);
or U24985 (N_24985,N_24699,N_24522);
xor U24986 (N_24986,N_24686,N_24567);
nand U24987 (N_24987,N_24521,N_24532);
nand U24988 (N_24988,N_24702,N_24739);
and U24989 (N_24989,N_24518,N_24667);
nor U24990 (N_24990,N_24529,N_24742);
nor U24991 (N_24991,N_24550,N_24667);
nor U24992 (N_24992,N_24716,N_24711);
and U24993 (N_24993,N_24537,N_24690);
nand U24994 (N_24994,N_24587,N_24637);
and U24995 (N_24995,N_24585,N_24710);
and U24996 (N_24996,N_24530,N_24606);
or U24997 (N_24997,N_24502,N_24516);
xnor U24998 (N_24998,N_24532,N_24684);
and U24999 (N_24999,N_24555,N_24641);
nor U25000 (N_25000,N_24928,N_24926);
nand U25001 (N_25001,N_24758,N_24831);
nand U25002 (N_25002,N_24810,N_24863);
and U25003 (N_25003,N_24833,N_24891);
or U25004 (N_25004,N_24756,N_24793);
nor U25005 (N_25005,N_24823,N_24857);
nand U25006 (N_25006,N_24826,N_24875);
xnor U25007 (N_25007,N_24750,N_24865);
xor U25008 (N_25008,N_24901,N_24805);
and U25009 (N_25009,N_24807,N_24950);
nor U25010 (N_25010,N_24917,N_24965);
nand U25011 (N_25011,N_24874,N_24999);
and U25012 (N_25012,N_24754,N_24936);
and U25013 (N_25013,N_24890,N_24829);
or U25014 (N_25014,N_24952,N_24860);
and U25015 (N_25015,N_24771,N_24939);
nor U25016 (N_25016,N_24900,N_24905);
xor U25017 (N_25017,N_24790,N_24902);
or U25018 (N_25018,N_24904,N_24947);
or U25019 (N_25019,N_24920,N_24861);
xnor U25020 (N_25020,N_24931,N_24948);
nor U25021 (N_25021,N_24795,N_24883);
and U25022 (N_25022,N_24963,N_24791);
nor U25023 (N_25023,N_24832,N_24751);
or U25024 (N_25024,N_24766,N_24982);
nand U25025 (N_25025,N_24755,N_24856);
nor U25026 (N_25026,N_24765,N_24946);
nor U25027 (N_25027,N_24867,N_24851);
nor U25028 (N_25028,N_24984,N_24786);
and U25029 (N_25029,N_24797,N_24888);
or U25030 (N_25030,N_24842,N_24814);
or U25031 (N_25031,N_24945,N_24896);
nand U25032 (N_25032,N_24998,N_24876);
nand U25033 (N_25033,N_24953,N_24873);
nor U25034 (N_25034,N_24824,N_24837);
xor U25035 (N_25035,N_24942,N_24898);
nor U25036 (N_25036,N_24803,N_24869);
or U25037 (N_25037,N_24944,N_24987);
xnor U25038 (N_25038,N_24897,N_24835);
and U25039 (N_25039,N_24990,N_24783);
and U25040 (N_25040,N_24956,N_24862);
and U25041 (N_25041,N_24870,N_24752);
nor U25042 (N_25042,N_24997,N_24911);
xnor U25043 (N_25043,N_24762,N_24871);
xor U25044 (N_25044,N_24817,N_24794);
nor U25045 (N_25045,N_24916,N_24877);
nand U25046 (N_25046,N_24922,N_24992);
nor U25047 (N_25047,N_24886,N_24976);
and U25048 (N_25048,N_24859,N_24971);
xnor U25049 (N_25049,N_24907,N_24789);
or U25050 (N_25050,N_24830,N_24772);
nor U25051 (N_25051,N_24769,N_24968);
or U25052 (N_25052,N_24966,N_24813);
xor U25053 (N_25053,N_24887,N_24819);
xnor U25054 (N_25054,N_24845,N_24913);
xnor U25055 (N_25055,N_24885,N_24753);
nor U25056 (N_25056,N_24800,N_24878);
xnor U25057 (N_25057,N_24903,N_24855);
or U25058 (N_25058,N_24972,N_24767);
or U25059 (N_25059,N_24843,N_24937);
xnor U25060 (N_25060,N_24778,N_24957);
nor U25061 (N_25061,N_24760,N_24989);
xor U25062 (N_25062,N_24784,N_24864);
nand U25063 (N_25063,N_24825,N_24774);
nor U25064 (N_25064,N_24983,N_24995);
or U25065 (N_25065,N_24785,N_24974);
xnor U25066 (N_25066,N_24960,N_24884);
xor U25067 (N_25067,N_24941,N_24923);
xor U25068 (N_25068,N_24872,N_24930);
or U25069 (N_25069,N_24844,N_24943);
nand U25070 (N_25070,N_24763,N_24802);
and U25071 (N_25071,N_24777,N_24940);
xnor U25072 (N_25072,N_24882,N_24759);
nor U25073 (N_25073,N_24969,N_24918);
xor U25074 (N_25074,N_24840,N_24848);
nor U25075 (N_25075,N_24933,N_24836);
and U25076 (N_25076,N_24852,N_24838);
nor U25077 (N_25077,N_24906,N_24993);
and U25078 (N_25078,N_24799,N_24964);
and U25079 (N_25079,N_24975,N_24775);
nor U25080 (N_25080,N_24914,N_24949);
and U25081 (N_25081,N_24812,N_24955);
xor U25082 (N_25082,N_24776,N_24881);
nand U25083 (N_25083,N_24757,N_24994);
and U25084 (N_25084,N_24980,N_24816);
or U25085 (N_25085,N_24868,N_24927);
xor U25086 (N_25086,N_24996,N_24818);
nand U25087 (N_25087,N_24796,N_24787);
xnor U25088 (N_25088,N_24951,N_24827);
xor U25089 (N_25089,N_24921,N_24915);
nor U25090 (N_25090,N_24821,N_24978);
nor U25091 (N_25091,N_24973,N_24853);
xor U25092 (N_25092,N_24962,N_24909);
xor U25093 (N_25093,N_24822,N_24924);
nand U25094 (N_25094,N_24985,N_24792);
and U25095 (N_25095,N_24764,N_24908);
nand U25096 (N_25096,N_24910,N_24834);
nor U25097 (N_25097,N_24815,N_24761);
nor U25098 (N_25098,N_24954,N_24806);
and U25099 (N_25099,N_24991,N_24970);
or U25100 (N_25100,N_24979,N_24899);
or U25101 (N_25101,N_24811,N_24770);
nor U25102 (N_25102,N_24798,N_24849);
or U25103 (N_25103,N_24894,N_24892);
nor U25104 (N_25104,N_24929,N_24820);
xnor U25105 (N_25105,N_24773,N_24977);
or U25106 (N_25106,N_24801,N_24854);
and U25107 (N_25107,N_24934,N_24893);
xnor U25108 (N_25108,N_24958,N_24850);
nand U25109 (N_25109,N_24932,N_24839);
and U25110 (N_25110,N_24809,N_24959);
or U25111 (N_25111,N_24919,N_24866);
or U25112 (N_25112,N_24808,N_24858);
nand U25113 (N_25113,N_24779,N_24879);
or U25114 (N_25114,N_24782,N_24780);
or U25115 (N_25115,N_24925,N_24889);
xor U25116 (N_25116,N_24967,N_24912);
and U25117 (N_25117,N_24935,N_24895);
nand U25118 (N_25118,N_24828,N_24880);
and U25119 (N_25119,N_24988,N_24847);
and U25120 (N_25120,N_24781,N_24981);
or U25121 (N_25121,N_24938,N_24768);
xor U25122 (N_25122,N_24841,N_24804);
xnor U25123 (N_25123,N_24846,N_24986);
nor U25124 (N_25124,N_24788,N_24961);
nor U25125 (N_25125,N_24841,N_24837);
nand U25126 (N_25126,N_24773,N_24815);
xor U25127 (N_25127,N_24881,N_24949);
xnor U25128 (N_25128,N_24786,N_24809);
xnor U25129 (N_25129,N_24960,N_24932);
or U25130 (N_25130,N_24973,N_24929);
and U25131 (N_25131,N_24772,N_24847);
or U25132 (N_25132,N_24971,N_24839);
xnor U25133 (N_25133,N_24983,N_24774);
or U25134 (N_25134,N_24890,N_24757);
nand U25135 (N_25135,N_24819,N_24853);
nor U25136 (N_25136,N_24852,N_24877);
or U25137 (N_25137,N_24754,N_24821);
nand U25138 (N_25138,N_24962,N_24977);
nor U25139 (N_25139,N_24971,N_24887);
and U25140 (N_25140,N_24944,N_24827);
nor U25141 (N_25141,N_24843,N_24994);
nand U25142 (N_25142,N_24845,N_24830);
nor U25143 (N_25143,N_24869,N_24877);
and U25144 (N_25144,N_24894,N_24988);
and U25145 (N_25145,N_24886,N_24755);
nand U25146 (N_25146,N_24816,N_24822);
nor U25147 (N_25147,N_24817,N_24829);
nand U25148 (N_25148,N_24919,N_24802);
and U25149 (N_25149,N_24810,N_24768);
and U25150 (N_25150,N_24909,N_24894);
and U25151 (N_25151,N_24806,N_24933);
nor U25152 (N_25152,N_24940,N_24854);
and U25153 (N_25153,N_24837,N_24977);
or U25154 (N_25154,N_24876,N_24852);
or U25155 (N_25155,N_24902,N_24862);
xor U25156 (N_25156,N_24761,N_24819);
xor U25157 (N_25157,N_24849,N_24787);
xnor U25158 (N_25158,N_24825,N_24822);
and U25159 (N_25159,N_24824,N_24944);
nor U25160 (N_25160,N_24829,N_24865);
xor U25161 (N_25161,N_24998,N_24852);
nand U25162 (N_25162,N_24846,N_24913);
xor U25163 (N_25163,N_24810,N_24997);
nor U25164 (N_25164,N_24871,N_24798);
nor U25165 (N_25165,N_24965,N_24772);
and U25166 (N_25166,N_24980,N_24851);
and U25167 (N_25167,N_24914,N_24872);
and U25168 (N_25168,N_24986,N_24989);
and U25169 (N_25169,N_24909,N_24864);
and U25170 (N_25170,N_24854,N_24952);
or U25171 (N_25171,N_24967,N_24843);
or U25172 (N_25172,N_24754,N_24824);
nand U25173 (N_25173,N_24868,N_24770);
xnor U25174 (N_25174,N_24861,N_24883);
xnor U25175 (N_25175,N_24997,N_24955);
or U25176 (N_25176,N_24975,N_24839);
xnor U25177 (N_25177,N_24990,N_24947);
nor U25178 (N_25178,N_24891,N_24766);
nor U25179 (N_25179,N_24823,N_24791);
and U25180 (N_25180,N_24780,N_24762);
xor U25181 (N_25181,N_24914,N_24834);
and U25182 (N_25182,N_24997,N_24776);
nor U25183 (N_25183,N_24944,N_24837);
nand U25184 (N_25184,N_24831,N_24951);
nor U25185 (N_25185,N_24814,N_24760);
xnor U25186 (N_25186,N_24914,N_24916);
nor U25187 (N_25187,N_24979,N_24760);
or U25188 (N_25188,N_24791,N_24797);
xor U25189 (N_25189,N_24836,N_24818);
nor U25190 (N_25190,N_24924,N_24913);
or U25191 (N_25191,N_24770,N_24853);
or U25192 (N_25192,N_24971,N_24801);
nor U25193 (N_25193,N_24894,N_24817);
xor U25194 (N_25194,N_24931,N_24913);
nand U25195 (N_25195,N_24992,N_24758);
nor U25196 (N_25196,N_24962,N_24767);
nand U25197 (N_25197,N_24928,N_24823);
nand U25198 (N_25198,N_24835,N_24986);
xor U25199 (N_25199,N_24893,N_24850);
nand U25200 (N_25200,N_24931,N_24768);
or U25201 (N_25201,N_24943,N_24868);
nand U25202 (N_25202,N_24862,N_24886);
or U25203 (N_25203,N_24815,N_24758);
nor U25204 (N_25204,N_24984,N_24966);
nor U25205 (N_25205,N_24937,N_24962);
xor U25206 (N_25206,N_24958,N_24864);
nand U25207 (N_25207,N_24874,N_24887);
nand U25208 (N_25208,N_24932,N_24887);
and U25209 (N_25209,N_24953,N_24941);
or U25210 (N_25210,N_24875,N_24966);
or U25211 (N_25211,N_24894,N_24860);
xnor U25212 (N_25212,N_24823,N_24912);
and U25213 (N_25213,N_24768,N_24906);
nor U25214 (N_25214,N_24871,N_24808);
nor U25215 (N_25215,N_24823,N_24993);
xor U25216 (N_25216,N_24971,N_24879);
and U25217 (N_25217,N_24950,N_24870);
nand U25218 (N_25218,N_24992,N_24866);
nor U25219 (N_25219,N_24900,N_24985);
or U25220 (N_25220,N_24889,N_24954);
and U25221 (N_25221,N_24943,N_24806);
nand U25222 (N_25222,N_24818,N_24938);
nor U25223 (N_25223,N_24884,N_24944);
and U25224 (N_25224,N_24850,N_24962);
or U25225 (N_25225,N_24928,N_24935);
nand U25226 (N_25226,N_24773,N_24939);
xor U25227 (N_25227,N_24842,N_24811);
xor U25228 (N_25228,N_24787,N_24910);
nand U25229 (N_25229,N_24829,N_24775);
and U25230 (N_25230,N_24788,N_24857);
or U25231 (N_25231,N_24949,N_24956);
or U25232 (N_25232,N_24913,N_24860);
nor U25233 (N_25233,N_24768,N_24816);
xor U25234 (N_25234,N_24879,N_24878);
nor U25235 (N_25235,N_24896,N_24964);
and U25236 (N_25236,N_24951,N_24820);
nand U25237 (N_25237,N_24878,N_24758);
or U25238 (N_25238,N_24919,N_24891);
nand U25239 (N_25239,N_24951,N_24805);
or U25240 (N_25240,N_24992,N_24945);
nor U25241 (N_25241,N_24956,N_24934);
nand U25242 (N_25242,N_24796,N_24944);
nor U25243 (N_25243,N_24829,N_24783);
and U25244 (N_25244,N_24821,N_24971);
or U25245 (N_25245,N_24837,N_24852);
or U25246 (N_25246,N_24940,N_24990);
nor U25247 (N_25247,N_24768,N_24785);
nand U25248 (N_25248,N_24787,N_24808);
or U25249 (N_25249,N_24781,N_24994);
nor U25250 (N_25250,N_25014,N_25082);
nand U25251 (N_25251,N_25152,N_25195);
nand U25252 (N_25252,N_25235,N_25008);
or U25253 (N_25253,N_25029,N_25180);
nand U25254 (N_25254,N_25228,N_25208);
or U25255 (N_25255,N_25081,N_25074);
nor U25256 (N_25256,N_25194,N_25158);
xor U25257 (N_25257,N_25080,N_25185);
xor U25258 (N_25258,N_25100,N_25056);
or U25259 (N_25259,N_25226,N_25116);
nor U25260 (N_25260,N_25247,N_25097);
or U25261 (N_25261,N_25034,N_25010);
or U25262 (N_25262,N_25012,N_25045);
nor U25263 (N_25263,N_25069,N_25085);
and U25264 (N_25264,N_25087,N_25248);
or U25265 (N_25265,N_25172,N_25162);
nand U25266 (N_25266,N_25213,N_25057);
or U25267 (N_25267,N_25019,N_25217);
nor U25268 (N_25268,N_25063,N_25109);
xnor U25269 (N_25269,N_25126,N_25143);
and U25270 (N_25270,N_25234,N_25086);
xor U25271 (N_25271,N_25090,N_25117);
or U25272 (N_25272,N_25223,N_25161);
nor U25273 (N_25273,N_25121,N_25134);
nor U25274 (N_25274,N_25065,N_25214);
xnor U25275 (N_25275,N_25037,N_25233);
or U25276 (N_25276,N_25036,N_25089);
nor U25277 (N_25277,N_25154,N_25104);
or U25278 (N_25278,N_25098,N_25030);
xnor U25279 (N_25279,N_25165,N_25220);
xor U25280 (N_25280,N_25093,N_25201);
or U25281 (N_25281,N_25106,N_25011);
nand U25282 (N_25282,N_25148,N_25105);
nand U25283 (N_25283,N_25039,N_25151);
xnor U25284 (N_25284,N_25237,N_25156);
and U25285 (N_25285,N_25055,N_25038);
and U25286 (N_25286,N_25227,N_25033);
or U25287 (N_25287,N_25197,N_25127);
nand U25288 (N_25288,N_25130,N_25108);
or U25289 (N_25289,N_25068,N_25198);
nand U25290 (N_25290,N_25142,N_25187);
xnor U25291 (N_25291,N_25167,N_25112);
nand U25292 (N_25292,N_25219,N_25169);
or U25293 (N_25293,N_25231,N_25072);
nor U25294 (N_25294,N_25230,N_25009);
nand U25295 (N_25295,N_25168,N_25027);
and U25296 (N_25296,N_25079,N_25204);
and U25297 (N_25297,N_25184,N_25005);
nand U25298 (N_25298,N_25196,N_25071);
nor U25299 (N_25299,N_25173,N_25041);
nor U25300 (N_25300,N_25249,N_25075);
and U25301 (N_25301,N_25192,N_25017);
nand U25302 (N_25302,N_25094,N_25114);
nor U25303 (N_25303,N_25132,N_25001);
xnor U25304 (N_25304,N_25031,N_25244);
nor U25305 (N_25305,N_25129,N_25091);
or U25306 (N_25306,N_25178,N_25175);
nand U25307 (N_25307,N_25243,N_25177);
or U25308 (N_25308,N_25170,N_25006);
nor U25309 (N_25309,N_25061,N_25174);
and U25310 (N_25310,N_25042,N_25125);
or U25311 (N_25311,N_25115,N_25200);
nand U25312 (N_25312,N_25035,N_25157);
or U25313 (N_25313,N_25164,N_25051);
or U25314 (N_25314,N_25147,N_25003);
nand U25315 (N_25315,N_25242,N_25216);
or U25316 (N_25316,N_25120,N_25007);
nor U25317 (N_25317,N_25040,N_25203);
and U25318 (N_25318,N_25206,N_25189);
nand U25319 (N_25319,N_25163,N_25171);
nand U25320 (N_25320,N_25190,N_25224);
xnor U25321 (N_25321,N_25060,N_25021);
and U25322 (N_25322,N_25054,N_25043);
xor U25323 (N_25323,N_25016,N_25092);
nor U25324 (N_25324,N_25077,N_25133);
xor U25325 (N_25325,N_25084,N_25212);
nand U25326 (N_25326,N_25229,N_25053);
nor U25327 (N_25327,N_25241,N_25245);
and U25328 (N_25328,N_25066,N_25179);
xnor U25329 (N_25329,N_25232,N_25131);
and U25330 (N_25330,N_25225,N_25102);
xnor U25331 (N_25331,N_25062,N_25070);
and U25332 (N_25332,N_25078,N_25236);
nand U25333 (N_25333,N_25160,N_25015);
nand U25334 (N_25334,N_25150,N_25183);
and U25335 (N_25335,N_25095,N_25122);
nor U25336 (N_25336,N_25064,N_25155);
and U25337 (N_25337,N_25159,N_25026);
or U25338 (N_25338,N_25099,N_25018);
or U25339 (N_25339,N_25211,N_25210);
nor U25340 (N_25340,N_25144,N_25149);
and U25341 (N_25341,N_25145,N_25146);
or U25342 (N_25342,N_25119,N_25000);
nand U25343 (N_25343,N_25222,N_25181);
nand U25344 (N_25344,N_25140,N_25118);
nor U25345 (N_25345,N_25137,N_25193);
and U25346 (N_25346,N_25088,N_25028);
and U25347 (N_25347,N_25020,N_25207);
or U25348 (N_25348,N_25024,N_25059);
and U25349 (N_25349,N_25110,N_25246);
and U25350 (N_25350,N_25101,N_25141);
xor U25351 (N_25351,N_25046,N_25103);
xnor U25352 (N_25352,N_25073,N_25067);
nand U25353 (N_25353,N_25153,N_25218);
nand U25354 (N_25354,N_25023,N_25044);
nor U25355 (N_25355,N_25139,N_25215);
nor U25356 (N_25356,N_25025,N_25050);
and U25357 (N_25357,N_25138,N_25188);
or U25358 (N_25358,N_25111,N_25113);
nand U25359 (N_25359,N_25022,N_25047);
xnor U25360 (N_25360,N_25083,N_25209);
or U25361 (N_25361,N_25002,N_25032);
or U25362 (N_25362,N_25124,N_25096);
xor U25363 (N_25363,N_25221,N_25166);
xnor U25364 (N_25364,N_25004,N_25238);
xor U25365 (N_25365,N_25123,N_25202);
xor U25366 (N_25366,N_25239,N_25186);
xor U25367 (N_25367,N_25191,N_25048);
or U25368 (N_25368,N_25013,N_25136);
and U25369 (N_25369,N_25049,N_25182);
nand U25370 (N_25370,N_25058,N_25205);
xor U25371 (N_25371,N_25128,N_25240);
nor U25372 (N_25372,N_25076,N_25199);
xor U25373 (N_25373,N_25052,N_25135);
and U25374 (N_25374,N_25107,N_25176);
xnor U25375 (N_25375,N_25114,N_25055);
xor U25376 (N_25376,N_25136,N_25209);
nand U25377 (N_25377,N_25212,N_25226);
nor U25378 (N_25378,N_25104,N_25215);
nand U25379 (N_25379,N_25085,N_25108);
nand U25380 (N_25380,N_25082,N_25216);
xnor U25381 (N_25381,N_25063,N_25019);
nand U25382 (N_25382,N_25206,N_25070);
nor U25383 (N_25383,N_25035,N_25030);
nand U25384 (N_25384,N_25111,N_25033);
and U25385 (N_25385,N_25104,N_25087);
nand U25386 (N_25386,N_25015,N_25089);
and U25387 (N_25387,N_25233,N_25201);
and U25388 (N_25388,N_25061,N_25151);
and U25389 (N_25389,N_25145,N_25026);
or U25390 (N_25390,N_25081,N_25215);
or U25391 (N_25391,N_25230,N_25071);
xor U25392 (N_25392,N_25138,N_25217);
nand U25393 (N_25393,N_25012,N_25227);
or U25394 (N_25394,N_25091,N_25082);
xnor U25395 (N_25395,N_25002,N_25161);
nand U25396 (N_25396,N_25024,N_25249);
or U25397 (N_25397,N_25126,N_25048);
nand U25398 (N_25398,N_25043,N_25180);
nand U25399 (N_25399,N_25087,N_25210);
or U25400 (N_25400,N_25173,N_25011);
xor U25401 (N_25401,N_25104,N_25159);
nand U25402 (N_25402,N_25005,N_25126);
nor U25403 (N_25403,N_25031,N_25192);
nor U25404 (N_25404,N_25162,N_25130);
or U25405 (N_25405,N_25041,N_25016);
and U25406 (N_25406,N_25172,N_25119);
and U25407 (N_25407,N_25208,N_25011);
xor U25408 (N_25408,N_25041,N_25020);
nor U25409 (N_25409,N_25117,N_25180);
and U25410 (N_25410,N_25009,N_25222);
nor U25411 (N_25411,N_25059,N_25210);
and U25412 (N_25412,N_25083,N_25038);
xor U25413 (N_25413,N_25066,N_25068);
xor U25414 (N_25414,N_25135,N_25200);
nor U25415 (N_25415,N_25127,N_25099);
xor U25416 (N_25416,N_25012,N_25222);
and U25417 (N_25417,N_25030,N_25216);
or U25418 (N_25418,N_25042,N_25248);
nand U25419 (N_25419,N_25036,N_25083);
or U25420 (N_25420,N_25018,N_25203);
nor U25421 (N_25421,N_25097,N_25134);
and U25422 (N_25422,N_25032,N_25028);
xor U25423 (N_25423,N_25036,N_25175);
xor U25424 (N_25424,N_25234,N_25096);
xnor U25425 (N_25425,N_25169,N_25132);
nor U25426 (N_25426,N_25247,N_25086);
or U25427 (N_25427,N_25092,N_25137);
nor U25428 (N_25428,N_25098,N_25231);
xnor U25429 (N_25429,N_25086,N_25201);
nor U25430 (N_25430,N_25224,N_25150);
nor U25431 (N_25431,N_25145,N_25091);
and U25432 (N_25432,N_25216,N_25116);
or U25433 (N_25433,N_25063,N_25086);
nand U25434 (N_25434,N_25103,N_25174);
xnor U25435 (N_25435,N_25117,N_25164);
nand U25436 (N_25436,N_25096,N_25039);
or U25437 (N_25437,N_25074,N_25003);
and U25438 (N_25438,N_25141,N_25103);
nand U25439 (N_25439,N_25154,N_25246);
xor U25440 (N_25440,N_25152,N_25013);
nand U25441 (N_25441,N_25209,N_25170);
nor U25442 (N_25442,N_25173,N_25125);
nand U25443 (N_25443,N_25217,N_25125);
xnor U25444 (N_25444,N_25159,N_25177);
or U25445 (N_25445,N_25069,N_25014);
nand U25446 (N_25446,N_25058,N_25102);
xnor U25447 (N_25447,N_25155,N_25051);
nor U25448 (N_25448,N_25161,N_25107);
xor U25449 (N_25449,N_25158,N_25136);
xnor U25450 (N_25450,N_25187,N_25231);
nand U25451 (N_25451,N_25102,N_25139);
nor U25452 (N_25452,N_25190,N_25196);
or U25453 (N_25453,N_25172,N_25208);
or U25454 (N_25454,N_25187,N_25245);
xor U25455 (N_25455,N_25235,N_25037);
and U25456 (N_25456,N_25055,N_25043);
and U25457 (N_25457,N_25129,N_25137);
nor U25458 (N_25458,N_25068,N_25000);
and U25459 (N_25459,N_25246,N_25203);
or U25460 (N_25460,N_25010,N_25227);
or U25461 (N_25461,N_25074,N_25078);
xor U25462 (N_25462,N_25182,N_25096);
nor U25463 (N_25463,N_25090,N_25223);
and U25464 (N_25464,N_25233,N_25147);
xor U25465 (N_25465,N_25198,N_25060);
nor U25466 (N_25466,N_25201,N_25177);
nor U25467 (N_25467,N_25101,N_25021);
nand U25468 (N_25468,N_25138,N_25122);
xor U25469 (N_25469,N_25174,N_25122);
nor U25470 (N_25470,N_25023,N_25058);
or U25471 (N_25471,N_25153,N_25131);
xnor U25472 (N_25472,N_25240,N_25180);
nand U25473 (N_25473,N_25128,N_25188);
nor U25474 (N_25474,N_25191,N_25244);
and U25475 (N_25475,N_25160,N_25135);
nand U25476 (N_25476,N_25076,N_25036);
xnor U25477 (N_25477,N_25176,N_25083);
nor U25478 (N_25478,N_25027,N_25075);
nand U25479 (N_25479,N_25166,N_25201);
nor U25480 (N_25480,N_25186,N_25163);
xor U25481 (N_25481,N_25039,N_25009);
and U25482 (N_25482,N_25087,N_25121);
xor U25483 (N_25483,N_25048,N_25154);
nor U25484 (N_25484,N_25209,N_25172);
and U25485 (N_25485,N_25083,N_25220);
and U25486 (N_25486,N_25091,N_25121);
and U25487 (N_25487,N_25154,N_25114);
nand U25488 (N_25488,N_25094,N_25040);
nand U25489 (N_25489,N_25178,N_25214);
xor U25490 (N_25490,N_25036,N_25167);
or U25491 (N_25491,N_25162,N_25095);
nand U25492 (N_25492,N_25023,N_25234);
and U25493 (N_25493,N_25174,N_25150);
or U25494 (N_25494,N_25219,N_25150);
nand U25495 (N_25495,N_25225,N_25078);
xnor U25496 (N_25496,N_25009,N_25219);
nand U25497 (N_25497,N_25197,N_25056);
and U25498 (N_25498,N_25172,N_25127);
and U25499 (N_25499,N_25116,N_25147);
nand U25500 (N_25500,N_25458,N_25366);
or U25501 (N_25501,N_25394,N_25470);
or U25502 (N_25502,N_25473,N_25362);
nor U25503 (N_25503,N_25280,N_25281);
nand U25504 (N_25504,N_25369,N_25256);
and U25505 (N_25505,N_25445,N_25254);
or U25506 (N_25506,N_25498,N_25252);
or U25507 (N_25507,N_25389,N_25487);
and U25508 (N_25508,N_25271,N_25469);
nand U25509 (N_25509,N_25456,N_25272);
and U25510 (N_25510,N_25301,N_25294);
or U25511 (N_25511,N_25435,N_25467);
or U25512 (N_25512,N_25411,N_25448);
or U25513 (N_25513,N_25332,N_25292);
xor U25514 (N_25514,N_25431,N_25494);
and U25515 (N_25515,N_25270,N_25402);
nand U25516 (N_25516,N_25443,N_25282);
nor U25517 (N_25517,N_25263,N_25380);
or U25518 (N_25518,N_25387,N_25264);
xnor U25519 (N_25519,N_25315,N_25462);
nand U25520 (N_25520,N_25339,N_25317);
or U25521 (N_25521,N_25419,N_25365);
or U25522 (N_25522,N_25348,N_25491);
nor U25523 (N_25523,N_25440,N_25259);
and U25524 (N_25524,N_25401,N_25261);
or U25525 (N_25525,N_25396,N_25316);
nor U25526 (N_25526,N_25363,N_25475);
xnor U25527 (N_25527,N_25482,N_25437);
and U25528 (N_25528,N_25426,N_25346);
nor U25529 (N_25529,N_25367,N_25432);
xor U25530 (N_25530,N_25405,N_25488);
nand U25531 (N_25531,N_25409,N_25283);
and U25532 (N_25532,N_25327,N_25388);
and U25533 (N_25533,N_25260,N_25342);
nand U25534 (N_25534,N_25433,N_25353);
xnor U25535 (N_25535,N_25313,N_25345);
nand U25536 (N_25536,N_25321,N_25421);
or U25537 (N_25537,N_25459,N_25429);
nand U25538 (N_25538,N_25464,N_25335);
or U25539 (N_25539,N_25299,N_25490);
and U25540 (N_25540,N_25434,N_25293);
and U25541 (N_25541,N_25323,N_25436);
or U25542 (N_25542,N_25308,N_25287);
or U25543 (N_25543,N_25331,N_25472);
or U25544 (N_25544,N_25251,N_25476);
nor U25545 (N_25545,N_25408,N_25414);
xor U25546 (N_25546,N_25398,N_25305);
and U25547 (N_25547,N_25262,N_25463);
nor U25548 (N_25548,N_25274,N_25314);
nand U25549 (N_25549,N_25413,N_25350);
or U25550 (N_25550,N_25360,N_25297);
and U25551 (N_25551,N_25286,N_25338);
and U25552 (N_25552,N_25306,N_25382);
nand U25553 (N_25553,N_25478,N_25372);
nor U25554 (N_25554,N_25361,N_25311);
and U25555 (N_25555,N_25291,N_25474);
nor U25556 (N_25556,N_25495,N_25406);
nor U25557 (N_25557,N_25275,N_25298);
nor U25558 (N_25558,N_25452,N_25442);
nor U25559 (N_25559,N_25253,N_25358);
or U25560 (N_25560,N_25289,N_25438);
xor U25561 (N_25561,N_25352,N_25393);
and U25562 (N_25562,N_25391,N_25412);
nand U25563 (N_25563,N_25480,N_25325);
nand U25564 (N_25564,N_25334,N_25343);
nor U25565 (N_25565,N_25479,N_25385);
nor U25566 (N_25566,N_25492,N_25303);
xor U25567 (N_25567,N_25277,N_25466);
or U25568 (N_25568,N_25320,N_25288);
nand U25569 (N_25569,N_25446,N_25304);
xnor U25570 (N_25570,N_25395,N_25255);
and U25571 (N_25571,N_25290,N_25450);
nor U25572 (N_25572,N_25424,N_25376);
nor U25573 (N_25573,N_25453,N_25307);
nand U25574 (N_25574,N_25266,N_25422);
nor U25575 (N_25575,N_25379,N_25423);
nand U25576 (N_25576,N_25399,N_25383);
xor U25577 (N_25577,N_25444,N_25425);
xor U25578 (N_25578,N_25499,N_25344);
nand U25579 (N_25579,N_25460,N_25356);
and U25580 (N_25580,N_25430,N_25310);
nor U25581 (N_25581,N_25333,N_25373);
or U25582 (N_25582,N_25378,N_25324);
xnor U25583 (N_25583,N_25454,N_25349);
and U25584 (N_25584,N_25329,N_25357);
nor U25585 (N_25585,N_25328,N_25269);
xor U25586 (N_25586,N_25319,N_25265);
nand U25587 (N_25587,N_25347,N_25485);
or U25588 (N_25588,N_25447,N_25354);
xor U25589 (N_25589,N_25340,N_25497);
xnor U25590 (N_25590,N_25420,N_25471);
and U25591 (N_25591,N_25455,N_25489);
nand U25592 (N_25592,N_25410,N_25461);
or U25593 (N_25593,N_25381,N_25359);
nor U25594 (N_25594,N_25400,N_25322);
or U25595 (N_25595,N_25364,N_25428);
or U25596 (N_25596,N_25415,N_25465);
and U25597 (N_25597,N_25337,N_25375);
nand U25598 (N_25598,N_25493,N_25302);
or U25599 (N_25599,N_25392,N_25377);
and U25600 (N_25600,N_25427,N_25407);
nand U25601 (N_25601,N_25457,N_25257);
xor U25602 (N_25602,N_25451,N_25258);
and U25603 (N_25603,N_25355,N_25468);
and U25604 (N_25604,N_25449,N_25483);
xor U25605 (N_25605,N_25384,N_25390);
nor U25606 (N_25606,N_25300,N_25295);
nand U25607 (N_25607,N_25374,N_25278);
or U25608 (N_25608,N_25397,N_25296);
or U25609 (N_25609,N_25273,N_25351);
nor U25610 (N_25610,N_25368,N_25404);
xnor U25611 (N_25611,N_25268,N_25341);
nor U25612 (N_25612,N_25279,N_25439);
and U25613 (N_25613,N_25330,N_25416);
xnor U25614 (N_25614,N_25403,N_25417);
xnor U25615 (N_25615,N_25486,N_25267);
nand U25616 (N_25616,N_25496,N_25386);
nor U25617 (N_25617,N_25276,N_25312);
xnor U25618 (N_25618,N_25484,N_25336);
and U25619 (N_25619,N_25250,N_25285);
nand U25620 (N_25620,N_25441,N_25326);
nor U25621 (N_25621,N_25477,N_25284);
xnor U25622 (N_25622,N_25370,N_25371);
and U25623 (N_25623,N_25418,N_25481);
nand U25624 (N_25624,N_25309,N_25318);
and U25625 (N_25625,N_25328,N_25408);
and U25626 (N_25626,N_25296,N_25318);
nand U25627 (N_25627,N_25305,N_25386);
xor U25628 (N_25628,N_25382,N_25394);
nand U25629 (N_25629,N_25418,N_25268);
and U25630 (N_25630,N_25463,N_25390);
xor U25631 (N_25631,N_25445,N_25291);
nand U25632 (N_25632,N_25342,N_25410);
xnor U25633 (N_25633,N_25457,N_25499);
nand U25634 (N_25634,N_25278,N_25333);
or U25635 (N_25635,N_25265,N_25440);
nand U25636 (N_25636,N_25350,N_25329);
nand U25637 (N_25637,N_25293,N_25267);
xnor U25638 (N_25638,N_25416,N_25328);
nand U25639 (N_25639,N_25264,N_25456);
xnor U25640 (N_25640,N_25384,N_25405);
or U25641 (N_25641,N_25331,N_25268);
xor U25642 (N_25642,N_25359,N_25263);
and U25643 (N_25643,N_25305,N_25468);
and U25644 (N_25644,N_25332,N_25266);
and U25645 (N_25645,N_25405,N_25393);
nor U25646 (N_25646,N_25327,N_25334);
nand U25647 (N_25647,N_25394,N_25316);
nand U25648 (N_25648,N_25291,N_25440);
and U25649 (N_25649,N_25464,N_25410);
and U25650 (N_25650,N_25356,N_25317);
nand U25651 (N_25651,N_25456,N_25363);
and U25652 (N_25652,N_25367,N_25427);
or U25653 (N_25653,N_25469,N_25371);
nand U25654 (N_25654,N_25344,N_25480);
and U25655 (N_25655,N_25455,N_25397);
and U25656 (N_25656,N_25339,N_25391);
xnor U25657 (N_25657,N_25336,N_25257);
or U25658 (N_25658,N_25264,N_25401);
and U25659 (N_25659,N_25301,N_25465);
nand U25660 (N_25660,N_25367,N_25403);
or U25661 (N_25661,N_25281,N_25466);
nor U25662 (N_25662,N_25435,N_25319);
nor U25663 (N_25663,N_25336,N_25337);
and U25664 (N_25664,N_25347,N_25492);
nor U25665 (N_25665,N_25328,N_25334);
and U25666 (N_25666,N_25421,N_25473);
nand U25667 (N_25667,N_25461,N_25335);
nor U25668 (N_25668,N_25444,N_25251);
xnor U25669 (N_25669,N_25322,N_25430);
nor U25670 (N_25670,N_25302,N_25362);
or U25671 (N_25671,N_25440,N_25364);
nor U25672 (N_25672,N_25381,N_25288);
nor U25673 (N_25673,N_25491,N_25477);
and U25674 (N_25674,N_25354,N_25423);
nor U25675 (N_25675,N_25380,N_25362);
nand U25676 (N_25676,N_25487,N_25476);
nor U25677 (N_25677,N_25368,N_25405);
nor U25678 (N_25678,N_25271,N_25329);
nor U25679 (N_25679,N_25363,N_25425);
nand U25680 (N_25680,N_25415,N_25337);
nor U25681 (N_25681,N_25274,N_25412);
nand U25682 (N_25682,N_25376,N_25381);
or U25683 (N_25683,N_25300,N_25433);
nand U25684 (N_25684,N_25405,N_25490);
nor U25685 (N_25685,N_25464,N_25483);
nand U25686 (N_25686,N_25281,N_25316);
or U25687 (N_25687,N_25415,N_25470);
nor U25688 (N_25688,N_25372,N_25440);
and U25689 (N_25689,N_25354,N_25397);
or U25690 (N_25690,N_25494,N_25353);
xor U25691 (N_25691,N_25475,N_25291);
xor U25692 (N_25692,N_25387,N_25449);
xnor U25693 (N_25693,N_25286,N_25393);
xnor U25694 (N_25694,N_25498,N_25253);
nor U25695 (N_25695,N_25465,N_25429);
and U25696 (N_25696,N_25457,N_25461);
xor U25697 (N_25697,N_25359,N_25354);
nor U25698 (N_25698,N_25387,N_25345);
nor U25699 (N_25699,N_25303,N_25426);
or U25700 (N_25700,N_25294,N_25346);
or U25701 (N_25701,N_25313,N_25452);
xnor U25702 (N_25702,N_25251,N_25432);
nand U25703 (N_25703,N_25466,N_25388);
or U25704 (N_25704,N_25461,N_25416);
nand U25705 (N_25705,N_25348,N_25393);
xnor U25706 (N_25706,N_25275,N_25347);
nand U25707 (N_25707,N_25422,N_25361);
and U25708 (N_25708,N_25358,N_25351);
xnor U25709 (N_25709,N_25313,N_25421);
or U25710 (N_25710,N_25424,N_25333);
or U25711 (N_25711,N_25331,N_25259);
xor U25712 (N_25712,N_25467,N_25268);
xnor U25713 (N_25713,N_25418,N_25420);
and U25714 (N_25714,N_25415,N_25320);
xor U25715 (N_25715,N_25425,N_25346);
or U25716 (N_25716,N_25283,N_25400);
and U25717 (N_25717,N_25490,N_25464);
xor U25718 (N_25718,N_25306,N_25257);
nor U25719 (N_25719,N_25315,N_25267);
nand U25720 (N_25720,N_25378,N_25261);
xor U25721 (N_25721,N_25417,N_25268);
or U25722 (N_25722,N_25452,N_25373);
nand U25723 (N_25723,N_25276,N_25436);
or U25724 (N_25724,N_25479,N_25363);
or U25725 (N_25725,N_25365,N_25460);
and U25726 (N_25726,N_25480,N_25370);
nor U25727 (N_25727,N_25361,N_25409);
nand U25728 (N_25728,N_25280,N_25329);
nor U25729 (N_25729,N_25312,N_25452);
xnor U25730 (N_25730,N_25369,N_25315);
nor U25731 (N_25731,N_25468,N_25304);
and U25732 (N_25732,N_25455,N_25382);
nor U25733 (N_25733,N_25312,N_25424);
nand U25734 (N_25734,N_25451,N_25476);
xnor U25735 (N_25735,N_25284,N_25329);
and U25736 (N_25736,N_25444,N_25467);
nand U25737 (N_25737,N_25486,N_25320);
and U25738 (N_25738,N_25456,N_25423);
and U25739 (N_25739,N_25453,N_25418);
nand U25740 (N_25740,N_25468,N_25334);
and U25741 (N_25741,N_25295,N_25397);
nor U25742 (N_25742,N_25253,N_25357);
or U25743 (N_25743,N_25479,N_25446);
nor U25744 (N_25744,N_25388,N_25282);
nand U25745 (N_25745,N_25378,N_25262);
and U25746 (N_25746,N_25358,N_25285);
xor U25747 (N_25747,N_25343,N_25435);
or U25748 (N_25748,N_25414,N_25359);
xnor U25749 (N_25749,N_25439,N_25330);
nand U25750 (N_25750,N_25523,N_25603);
and U25751 (N_25751,N_25536,N_25596);
xnor U25752 (N_25752,N_25711,N_25532);
nor U25753 (N_25753,N_25599,N_25721);
or U25754 (N_25754,N_25724,N_25692);
xor U25755 (N_25755,N_25537,N_25632);
xnor U25756 (N_25756,N_25510,N_25633);
nand U25757 (N_25757,N_25549,N_25747);
nor U25758 (N_25758,N_25624,N_25635);
xor U25759 (N_25759,N_25584,N_25616);
xor U25760 (N_25760,N_25521,N_25547);
nor U25761 (N_25761,N_25503,N_25703);
nor U25762 (N_25762,N_25557,N_25745);
nand U25763 (N_25763,N_25589,N_25627);
or U25764 (N_25764,N_25680,N_25625);
nor U25765 (N_25765,N_25687,N_25585);
or U25766 (N_25766,N_25615,N_25689);
nand U25767 (N_25767,N_25611,N_25511);
nor U25768 (N_25768,N_25554,N_25727);
nor U25769 (N_25769,N_25746,N_25592);
or U25770 (N_25770,N_25588,N_25507);
and U25771 (N_25771,N_25606,N_25561);
and U25772 (N_25772,N_25518,N_25617);
and U25773 (N_25773,N_25720,N_25505);
nand U25774 (N_25774,N_25736,N_25709);
xor U25775 (N_25775,N_25701,N_25671);
or U25776 (N_25776,N_25545,N_25567);
xnor U25777 (N_25777,N_25504,N_25659);
or U25778 (N_25778,N_25691,N_25652);
and U25779 (N_25779,N_25639,N_25686);
and U25780 (N_25780,N_25621,N_25656);
and U25781 (N_25781,N_25675,N_25683);
nand U25782 (N_25782,N_25684,N_25710);
and U25783 (N_25783,N_25718,N_25682);
nand U25784 (N_25784,N_25548,N_25574);
xnor U25785 (N_25785,N_25622,N_25660);
xor U25786 (N_25786,N_25594,N_25642);
xor U25787 (N_25787,N_25716,N_25502);
or U25788 (N_25788,N_25693,N_25665);
nor U25789 (N_25789,N_25577,N_25733);
and U25790 (N_25790,N_25552,N_25732);
or U25791 (N_25791,N_25560,N_25590);
or U25792 (N_25792,N_25559,N_25737);
xor U25793 (N_25793,N_25661,N_25556);
nand U25794 (N_25794,N_25581,N_25512);
or U25795 (N_25795,N_25517,N_25648);
and U25796 (N_25796,N_25714,N_25658);
and U25797 (N_25797,N_25742,N_25728);
nand U25798 (N_25798,N_25748,N_25593);
or U25799 (N_25799,N_25651,N_25534);
nand U25800 (N_25800,N_25685,N_25717);
and U25801 (N_25801,N_25664,N_25631);
and U25802 (N_25802,N_25629,N_25605);
or U25803 (N_25803,N_25725,N_25630);
nor U25804 (N_25804,N_25530,N_25529);
xnor U25805 (N_25805,N_25587,N_25653);
or U25806 (N_25806,N_25515,N_25620);
nor U25807 (N_25807,N_25579,N_25739);
and U25808 (N_25808,N_25602,N_25525);
xnor U25809 (N_25809,N_25520,N_25688);
and U25810 (N_25810,N_25583,N_25668);
and U25811 (N_25811,N_25667,N_25508);
nand U25812 (N_25812,N_25726,N_25647);
nand U25813 (N_25813,N_25609,N_25705);
or U25814 (N_25814,N_25713,N_25626);
and U25815 (N_25815,N_25608,N_25575);
nor U25816 (N_25816,N_25550,N_25558);
nor U25817 (N_25817,N_25506,N_25731);
or U25818 (N_25818,N_25679,N_25519);
nor U25819 (N_25819,N_25514,N_25578);
or U25820 (N_25820,N_25663,N_25636);
xnor U25821 (N_25821,N_25734,N_25538);
nor U25822 (N_25822,N_25723,N_25531);
nor U25823 (N_25823,N_25528,N_25570);
and U25824 (N_25824,N_25553,N_25551);
xnor U25825 (N_25825,N_25522,N_25566);
nor U25826 (N_25826,N_25613,N_25641);
or U25827 (N_25827,N_25740,N_25696);
nor U25828 (N_25828,N_25712,N_25681);
nand U25829 (N_25829,N_25700,N_25612);
nand U25830 (N_25830,N_25535,N_25623);
or U25831 (N_25831,N_25513,N_25640);
nor U25832 (N_25832,N_25601,N_25618);
xnor U25833 (N_25833,N_25614,N_25673);
xnor U25834 (N_25834,N_25509,N_25657);
and U25835 (N_25835,N_25540,N_25695);
and U25836 (N_25836,N_25634,N_25743);
and U25837 (N_25837,N_25741,N_25676);
and U25838 (N_25838,N_25674,N_25730);
and U25839 (N_25839,N_25697,N_25638);
nor U25840 (N_25840,N_25654,N_25546);
xor U25841 (N_25841,N_25637,N_25662);
or U25842 (N_25842,N_25643,N_25543);
or U25843 (N_25843,N_25644,N_25500);
and U25844 (N_25844,N_25524,N_25738);
xor U25845 (N_25845,N_25544,N_25569);
xnor U25846 (N_25846,N_25600,N_25670);
or U25847 (N_25847,N_25672,N_25516);
nor U25848 (N_25848,N_25573,N_25649);
and U25849 (N_25849,N_25708,N_25580);
or U25850 (N_25850,N_25576,N_25735);
nor U25851 (N_25851,N_25722,N_25555);
or U25852 (N_25852,N_25607,N_25702);
or U25853 (N_25853,N_25565,N_25650);
or U25854 (N_25854,N_25646,N_25729);
nand U25855 (N_25855,N_25690,N_25645);
nor U25856 (N_25856,N_25563,N_25572);
and U25857 (N_25857,N_25704,N_25591);
and U25858 (N_25858,N_25597,N_25666);
nand U25859 (N_25859,N_25586,N_25598);
or U25860 (N_25860,N_25694,N_25604);
and U25861 (N_25861,N_25699,N_25719);
or U25862 (N_25862,N_25749,N_25564);
and U25863 (N_25863,N_25678,N_25571);
and U25864 (N_25864,N_25539,N_25533);
xnor U25865 (N_25865,N_25526,N_25568);
nand U25866 (N_25866,N_25619,N_25669);
xnor U25867 (N_25867,N_25655,N_25541);
and U25868 (N_25868,N_25715,N_25582);
and U25869 (N_25869,N_25542,N_25595);
or U25870 (N_25870,N_25706,N_25698);
nand U25871 (N_25871,N_25501,N_25628);
or U25872 (N_25872,N_25562,N_25527);
nand U25873 (N_25873,N_25744,N_25677);
and U25874 (N_25874,N_25610,N_25707);
nor U25875 (N_25875,N_25681,N_25651);
nor U25876 (N_25876,N_25713,N_25636);
nand U25877 (N_25877,N_25667,N_25532);
and U25878 (N_25878,N_25661,N_25590);
xor U25879 (N_25879,N_25692,N_25528);
and U25880 (N_25880,N_25652,N_25581);
and U25881 (N_25881,N_25616,N_25627);
and U25882 (N_25882,N_25573,N_25643);
or U25883 (N_25883,N_25700,N_25710);
or U25884 (N_25884,N_25606,N_25654);
and U25885 (N_25885,N_25541,N_25743);
or U25886 (N_25886,N_25588,N_25655);
nor U25887 (N_25887,N_25505,N_25603);
and U25888 (N_25888,N_25705,N_25695);
or U25889 (N_25889,N_25536,N_25503);
or U25890 (N_25890,N_25661,N_25619);
and U25891 (N_25891,N_25701,N_25738);
and U25892 (N_25892,N_25598,N_25511);
nand U25893 (N_25893,N_25627,N_25661);
and U25894 (N_25894,N_25608,N_25586);
or U25895 (N_25895,N_25630,N_25711);
xor U25896 (N_25896,N_25665,N_25662);
and U25897 (N_25897,N_25562,N_25631);
xnor U25898 (N_25898,N_25697,N_25513);
xor U25899 (N_25899,N_25552,N_25571);
nor U25900 (N_25900,N_25685,N_25544);
and U25901 (N_25901,N_25579,N_25602);
xor U25902 (N_25902,N_25684,N_25740);
nand U25903 (N_25903,N_25666,N_25640);
or U25904 (N_25904,N_25516,N_25690);
xor U25905 (N_25905,N_25732,N_25584);
xnor U25906 (N_25906,N_25573,N_25519);
and U25907 (N_25907,N_25607,N_25603);
xnor U25908 (N_25908,N_25726,N_25595);
xnor U25909 (N_25909,N_25595,N_25743);
and U25910 (N_25910,N_25663,N_25524);
nand U25911 (N_25911,N_25542,N_25543);
nor U25912 (N_25912,N_25533,N_25547);
and U25913 (N_25913,N_25680,N_25579);
nand U25914 (N_25914,N_25628,N_25573);
nor U25915 (N_25915,N_25700,N_25682);
nor U25916 (N_25916,N_25707,N_25622);
and U25917 (N_25917,N_25501,N_25705);
and U25918 (N_25918,N_25732,N_25583);
and U25919 (N_25919,N_25597,N_25694);
nor U25920 (N_25920,N_25562,N_25715);
or U25921 (N_25921,N_25723,N_25675);
xor U25922 (N_25922,N_25595,N_25530);
nor U25923 (N_25923,N_25704,N_25688);
and U25924 (N_25924,N_25724,N_25661);
xor U25925 (N_25925,N_25508,N_25723);
nor U25926 (N_25926,N_25522,N_25631);
nor U25927 (N_25927,N_25525,N_25515);
or U25928 (N_25928,N_25663,N_25747);
nor U25929 (N_25929,N_25655,N_25530);
nor U25930 (N_25930,N_25558,N_25570);
nor U25931 (N_25931,N_25633,N_25573);
xnor U25932 (N_25932,N_25591,N_25681);
xnor U25933 (N_25933,N_25725,N_25705);
xnor U25934 (N_25934,N_25694,N_25738);
or U25935 (N_25935,N_25554,N_25533);
xor U25936 (N_25936,N_25647,N_25662);
and U25937 (N_25937,N_25647,N_25747);
nor U25938 (N_25938,N_25556,N_25720);
nor U25939 (N_25939,N_25598,N_25550);
or U25940 (N_25940,N_25599,N_25686);
nand U25941 (N_25941,N_25642,N_25628);
or U25942 (N_25942,N_25608,N_25726);
nor U25943 (N_25943,N_25525,N_25678);
and U25944 (N_25944,N_25596,N_25600);
or U25945 (N_25945,N_25739,N_25526);
and U25946 (N_25946,N_25510,N_25515);
or U25947 (N_25947,N_25732,N_25699);
nand U25948 (N_25948,N_25508,N_25592);
nor U25949 (N_25949,N_25544,N_25627);
and U25950 (N_25950,N_25625,N_25538);
xnor U25951 (N_25951,N_25693,N_25690);
or U25952 (N_25952,N_25541,N_25567);
or U25953 (N_25953,N_25504,N_25506);
xnor U25954 (N_25954,N_25563,N_25560);
or U25955 (N_25955,N_25711,N_25703);
or U25956 (N_25956,N_25715,N_25741);
nand U25957 (N_25957,N_25612,N_25577);
nand U25958 (N_25958,N_25644,N_25662);
and U25959 (N_25959,N_25508,N_25583);
and U25960 (N_25960,N_25629,N_25616);
and U25961 (N_25961,N_25586,N_25589);
nand U25962 (N_25962,N_25580,N_25572);
nor U25963 (N_25963,N_25709,N_25595);
xnor U25964 (N_25964,N_25687,N_25524);
xor U25965 (N_25965,N_25642,N_25737);
and U25966 (N_25966,N_25627,N_25505);
nand U25967 (N_25967,N_25563,N_25629);
xor U25968 (N_25968,N_25622,N_25644);
nand U25969 (N_25969,N_25598,N_25514);
nand U25970 (N_25970,N_25533,N_25690);
or U25971 (N_25971,N_25570,N_25578);
and U25972 (N_25972,N_25731,N_25555);
xor U25973 (N_25973,N_25702,N_25543);
and U25974 (N_25974,N_25625,N_25748);
nor U25975 (N_25975,N_25699,N_25594);
and U25976 (N_25976,N_25743,N_25504);
or U25977 (N_25977,N_25727,N_25670);
or U25978 (N_25978,N_25638,N_25626);
nor U25979 (N_25979,N_25531,N_25719);
xor U25980 (N_25980,N_25643,N_25652);
or U25981 (N_25981,N_25742,N_25732);
and U25982 (N_25982,N_25500,N_25585);
nand U25983 (N_25983,N_25732,N_25643);
nand U25984 (N_25984,N_25520,N_25618);
or U25985 (N_25985,N_25693,N_25701);
nand U25986 (N_25986,N_25546,N_25605);
nand U25987 (N_25987,N_25612,N_25560);
xnor U25988 (N_25988,N_25537,N_25546);
xnor U25989 (N_25989,N_25557,N_25648);
nor U25990 (N_25990,N_25601,N_25734);
nor U25991 (N_25991,N_25735,N_25541);
and U25992 (N_25992,N_25703,N_25585);
xor U25993 (N_25993,N_25639,N_25685);
nand U25994 (N_25994,N_25575,N_25728);
nor U25995 (N_25995,N_25722,N_25659);
nand U25996 (N_25996,N_25679,N_25706);
nand U25997 (N_25997,N_25740,N_25561);
xor U25998 (N_25998,N_25608,N_25534);
nand U25999 (N_25999,N_25509,N_25548);
nand U26000 (N_26000,N_25891,N_25964);
or U26001 (N_26001,N_25876,N_25822);
xnor U26002 (N_26002,N_25843,N_25942);
nor U26003 (N_26003,N_25943,N_25773);
nand U26004 (N_26004,N_25811,N_25852);
xor U26005 (N_26005,N_25805,N_25982);
nor U26006 (N_26006,N_25798,N_25838);
nor U26007 (N_26007,N_25884,N_25904);
nor U26008 (N_26008,N_25810,N_25757);
and U26009 (N_26009,N_25901,N_25927);
nand U26010 (N_26010,N_25823,N_25941);
xnor U26011 (N_26011,N_25799,N_25778);
nand U26012 (N_26012,N_25958,N_25952);
nor U26013 (N_26013,N_25863,N_25989);
nand U26014 (N_26014,N_25839,N_25909);
nor U26015 (N_26015,N_25923,N_25753);
xor U26016 (N_26016,N_25750,N_25922);
nand U26017 (N_26017,N_25974,N_25968);
xnor U26018 (N_26018,N_25883,N_25987);
nand U26019 (N_26019,N_25981,N_25813);
and U26020 (N_26020,N_25944,N_25864);
nor U26021 (N_26021,N_25767,N_25930);
nand U26022 (N_26022,N_25874,N_25758);
nand U26023 (N_26023,N_25882,N_25996);
nor U26024 (N_26024,N_25752,N_25853);
nand U26025 (N_26025,N_25950,N_25755);
or U26026 (N_26026,N_25800,N_25803);
xnor U26027 (N_26027,N_25812,N_25972);
nand U26028 (N_26028,N_25781,N_25907);
and U26029 (N_26029,N_25910,N_25973);
nor U26030 (N_26030,N_25845,N_25848);
xnor U26031 (N_26031,N_25993,N_25826);
and U26032 (N_26032,N_25854,N_25946);
or U26033 (N_26033,N_25992,N_25963);
and U26034 (N_26034,N_25908,N_25881);
nand U26035 (N_26035,N_25977,N_25980);
nor U26036 (N_26036,N_25937,N_25868);
xnor U26037 (N_26037,N_25970,N_25962);
and U26038 (N_26038,N_25960,N_25903);
nand U26039 (N_26039,N_25762,N_25979);
and U26040 (N_26040,N_25784,N_25855);
nand U26041 (N_26041,N_25873,N_25985);
nor U26042 (N_26042,N_25774,N_25788);
xor U26043 (N_26043,N_25949,N_25911);
nor U26044 (N_26044,N_25835,N_25956);
nor U26045 (N_26045,N_25875,N_25790);
nand U26046 (N_26046,N_25915,N_25897);
or U26047 (N_26047,N_25841,N_25828);
xor U26048 (N_26048,N_25751,N_25804);
nand U26049 (N_26049,N_25861,N_25877);
or U26050 (N_26050,N_25765,N_25975);
xnor U26051 (N_26051,N_25865,N_25959);
or U26052 (N_26052,N_25791,N_25953);
nor U26053 (N_26053,N_25797,N_25764);
and U26054 (N_26054,N_25933,N_25991);
and U26055 (N_26055,N_25756,N_25986);
nand U26056 (N_26056,N_25997,N_25815);
nand U26057 (N_26057,N_25928,N_25916);
nor U26058 (N_26058,N_25990,N_25776);
nand U26059 (N_26059,N_25809,N_25779);
nor U26060 (N_26060,N_25772,N_25796);
and U26061 (N_26061,N_25777,N_25871);
or U26062 (N_26062,N_25880,N_25760);
or U26063 (N_26063,N_25917,N_25846);
nand U26064 (N_26064,N_25830,N_25939);
xor U26065 (N_26065,N_25870,N_25821);
nor U26066 (N_26066,N_25971,N_25999);
nor U26067 (N_26067,N_25894,N_25770);
or U26068 (N_26068,N_25820,N_25879);
and U26069 (N_26069,N_25878,N_25951);
nor U26070 (N_26070,N_25983,N_25890);
nand U26071 (N_26071,N_25806,N_25925);
nand U26072 (N_26072,N_25886,N_25988);
or U26073 (N_26073,N_25787,N_25827);
or U26074 (N_26074,N_25892,N_25836);
or U26075 (N_26075,N_25931,N_25783);
xor U26076 (N_26076,N_25965,N_25786);
xnor U26077 (N_26077,N_25947,N_25817);
nand U26078 (N_26078,N_25802,N_25775);
or U26079 (N_26079,N_25814,N_25899);
or U26080 (N_26080,N_25921,N_25795);
nor U26081 (N_26081,N_25829,N_25766);
xor U26082 (N_26082,N_25860,N_25789);
or U26083 (N_26083,N_25780,N_25831);
nor U26084 (N_26084,N_25867,N_25938);
or U26085 (N_26085,N_25936,N_25888);
xor U26086 (N_26086,N_25998,N_25819);
nand U26087 (N_26087,N_25954,N_25763);
nand U26088 (N_26088,N_25906,N_25898);
and U26089 (N_26089,N_25862,N_25818);
and U26090 (N_26090,N_25895,N_25832);
and U26091 (N_26091,N_25816,N_25842);
and U26092 (N_26092,N_25857,N_25978);
nand U26093 (N_26093,N_25896,N_25754);
xnor U26094 (N_26094,N_25900,N_25833);
or U26095 (N_26095,N_25966,N_25995);
or U26096 (N_26096,N_25926,N_25793);
nand U26097 (N_26097,N_25849,N_25924);
xnor U26098 (N_26098,N_25994,N_25825);
nand U26099 (N_26099,N_25856,N_25759);
nand U26100 (N_26100,N_25792,N_25955);
xnor U26101 (N_26101,N_25794,N_25887);
nor U26102 (N_26102,N_25914,N_25967);
or U26103 (N_26103,N_25957,N_25844);
and U26104 (N_26104,N_25769,N_25919);
xnor U26105 (N_26105,N_25934,N_25859);
and U26106 (N_26106,N_25824,N_25840);
nand U26107 (N_26107,N_25984,N_25976);
nor U26108 (N_26108,N_25929,N_25935);
or U26109 (N_26109,N_25869,N_25858);
or U26110 (N_26110,N_25885,N_25850);
xor U26111 (N_26111,N_25961,N_25851);
nor U26112 (N_26112,N_25834,N_25837);
xnor U26113 (N_26113,N_25771,N_25801);
or U26114 (N_26114,N_25889,N_25847);
xnor U26115 (N_26115,N_25902,N_25918);
and U26116 (N_26116,N_25913,N_25808);
or U26117 (N_26117,N_25807,N_25948);
nand U26118 (N_26118,N_25866,N_25782);
nand U26119 (N_26119,N_25768,N_25940);
nand U26120 (N_26120,N_25932,N_25905);
or U26121 (N_26121,N_25945,N_25920);
xor U26122 (N_26122,N_25872,N_25761);
nand U26123 (N_26123,N_25893,N_25969);
and U26124 (N_26124,N_25785,N_25912);
nand U26125 (N_26125,N_25809,N_25778);
or U26126 (N_26126,N_25758,N_25869);
xnor U26127 (N_26127,N_25994,N_25875);
xnor U26128 (N_26128,N_25905,N_25877);
nor U26129 (N_26129,N_25920,N_25830);
and U26130 (N_26130,N_25867,N_25917);
and U26131 (N_26131,N_25864,N_25888);
nand U26132 (N_26132,N_25809,N_25773);
nor U26133 (N_26133,N_25970,N_25785);
or U26134 (N_26134,N_25933,N_25819);
or U26135 (N_26135,N_25849,N_25853);
or U26136 (N_26136,N_25864,N_25936);
nand U26137 (N_26137,N_25889,N_25910);
nand U26138 (N_26138,N_25778,N_25768);
and U26139 (N_26139,N_25883,N_25875);
and U26140 (N_26140,N_25838,N_25941);
xnor U26141 (N_26141,N_25756,N_25766);
xnor U26142 (N_26142,N_25896,N_25977);
xor U26143 (N_26143,N_25839,N_25812);
xnor U26144 (N_26144,N_25898,N_25908);
nand U26145 (N_26145,N_25893,N_25936);
nand U26146 (N_26146,N_25989,N_25953);
xor U26147 (N_26147,N_25875,N_25849);
nand U26148 (N_26148,N_25858,N_25817);
nand U26149 (N_26149,N_25896,N_25809);
nand U26150 (N_26150,N_25794,N_25859);
or U26151 (N_26151,N_25885,N_25767);
nor U26152 (N_26152,N_25886,N_25861);
nand U26153 (N_26153,N_25791,N_25843);
and U26154 (N_26154,N_25778,N_25919);
xnor U26155 (N_26155,N_25936,N_25818);
nor U26156 (N_26156,N_25929,N_25856);
nand U26157 (N_26157,N_25782,N_25805);
xor U26158 (N_26158,N_25875,N_25835);
and U26159 (N_26159,N_25929,N_25926);
nor U26160 (N_26160,N_25812,N_25926);
and U26161 (N_26161,N_25949,N_25905);
and U26162 (N_26162,N_25900,N_25785);
and U26163 (N_26163,N_25782,N_25847);
and U26164 (N_26164,N_25913,N_25854);
and U26165 (N_26165,N_25751,N_25845);
xor U26166 (N_26166,N_25935,N_25913);
nand U26167 (N_26167,N_25753,N_25855);
and U26168 (N_26168,N_25759,N_25906);
xnor U26169 (N_26169,N_25768,N_25926);
and U26170 (N_26170,N_25857,N_25913);
nand U26171 (N_26171,N_25983,N_25892);
xor U26172 (N_26172,N_25954,N_25817);
nor U26173 (N_26173,N_25805,N_25789);
and U26174 (N_26174,N_25850,N_25956);
nor U26175 (N_26175,N_25905,N_25797);
or U26176 (N_26176,N_25998,N_25910);
or U26177 (N_26177,N_25798,N_25840);
or U26178 (N_26178,N_25767,N_25773);
nand U26179 (N_26179,N_25926,N_25813);
nand U26180 (N_26180,N_25901,N_25977);
and U26181 (N_26181,N_25899,N_25894);
nand U26182 (N_26182,N_25822,N_25921);
or U26183 (N_26183,N_25917,N_25771);
nand U26184 (N_26184,N_25860,N_25934);
or U26185 (N_26185,N_25794,N_25910);
and U26186 (N_26186,N_25759,N_25914);
nand U26187 (N_26187,N_25970,N_25927);
nor U26188 (N_26188,N_25937,N_25922);
nor U26189 (N_26189,N_25947,N_25914);
or U26190 (N_26190,N_25984,N_25988);
or U26191 (N_26191,N_25865,N_25974);
and U26192 (N_26192,N_25836,N_25853);
xnor U26193 (N_26193,N_25827,N_25792);
nor U26194 (N_26194,N_25964,N_25872);
xor U26195 (N_26195,N_25823,N_25851);
nand U26196 (N_26196,N_25864,N_25832);
nand U26197 (N_26197,N_25853,N_25851);
xor U26198 (N_26198,N_25808,N_25891);
xnor U26199 (N_26199,N_25923,N_25960);
and U26200 (N_26200,N_25826,N_25913);
nand U26201 (N_26201,N_25836,N_25816);
nand U26202 (N_26202,N_25830,N_25790);
xor U26203 (N_26203,N_25827,N_25824);
xor U26204 (N_26204,N_25843,N_25764);
or U26205 (N_26205,N_25904,N_25775);
nor U26206 (N_26206,N_25989,N_25792);
nor U26207 (N_26207,N_25793,N_25886);
nor U26208 (N_26208,N_25932,N_25953);
or U26209 (N_26209,N_25864,N_25752);
nor U26210 (N_26210,N_25880,N_25831);
or U26211 (N_26211,N_25935,N_25901);
and U26212 (N_26212,N_25989,N_25825);
xnor U26213 (N_26213,N_25956,N_25789);
nand U26214 (N_26214,N_25843,N_25754);
and U26215 (N_26215,N_25992,N_25866);
and U26216 (N_26216,N_25914,N_25957);
nor U26217 (N_26217,N_25977,N_25809);
or U26218 (N_26218,N_25867,N_25872);
xor U26219 (N_26219,N_25984,N_25967);
or U26220 (N_26220,N_25949,N_25980);
nand U26221 (N_26221,N_25823,N_25944);
or U26222 (N_26222,N_25850,N_25888);
or U26223 (N_26223,N_25870,N_25936);
and U26224 (N_26224,N_25925,N_25973);
or U26225 (N_26225,N_25772,N_25917);
xor U26226 (N_26226,N_25911,N_25876);
xnor U26227 (N_26227,N_25883,N_25996);
and U26228 (N_26228,N_25879,N_25974);
or U26229 (N_26229,N_25897,N_25783);
nor U26230 (N_26230,N_25762,N_25835);
nor U26231 (N_26231,N_25766,N_25771);
xnor U26232 (N_26232,N_25836,N_25939);
or U26233 (N_26233,N_25879,N_25842);
and U26234 (N_26234,N_25799,N_25851);
or U26235 (N_26235,N_25895,N_25864);
or U26236 (N_26236,N_25757,N_25798);
nor U26237 (N_26237,N_25955,N_25993);
and U26238 (N_26238,N_25856,N_25997);
nor U26239 (N_26239,N_25811,N_25839);
and U26240 (N_26240,N_25783,N_25837);
nor U26241 (N_26241,N_25976,N_25917);
or U26242 (N_26242,N_25995,N_25871);
xor U26243 (N_26243,N_25819,N_25856);
xnor U26244 (N_26244,N_25886,N_25786);
nand U26245 (N_26245,N_25805,N_25757);
or U26246 (N_26246,N_25956,N_25978);
nand U26247 (N_26247,N_25985,N_25840);
or U26248 (N_26248,N_25875,N_25782);
and U26249 (N_26249,N_25831,N_25972);
nor U26250 (N_26250,N_26190,N_26182);
and U26251 (N_26251,N_26152,N_26174);
nand U26252 (N_26252,N_26109,N_26185);
xor U26253 (N_26253,N_26036,N_26214);
xor U26254 (N_26254,N_26111,N_26249);
nor U26255 (N_26255,N_26072,N_26162);
or U26256 (N_26256,N_26010,N_26047);
nor U26257 (N_26257,N_26150,N_26153);
nand U26258 (N_26258,N_26195,N_26158);
nand U26259 (N_26259,N_26045,N_26227);
nor U26260 (N_26260,N_26240,N_26246);
nand U26261 (N_26261,N_26007,N_26101);
xnor U26262 (N_26262,N_26188,N_26141);
nor U26263 (N_26263,N_26247,N_26201);
or U26264 (N_26264,N_26066,N_26120);
or U26265 (N_26265,N_26049,N_26118);
xnor U26266 (N_26266,N_26226,N_26017);
and U26267 (N_26267,N_26027,N_26064);
or U26268 (N_26268,N_26128,N_26187);
and U26269 (N_26269,N_26197,N_26107);
nand U26270 (N_26270,N_26044,N_26229);
and U26271 (N_26271,N_26167,N_26024);
xor U26272 (N_26272,N_26077,N_26157);
and U26273 (N_26273,N_26029,N_26223);
nor U26274 (N_26274,N_26159,N_26209);
nand U26275 (N_26275,N_26138,N_26183);
or U26276 (N_26276,N_26095,N_26089);
nand U26277 (N_26277,N_26000,N_26173);
and U26278 (N_26278,N_26030,N_26222);
xor U26279 (N_26279,N_26093,N_26203);
nor U26280 (N_26280,N_26059,N_26042);
nor U26281 (N_26281,N_26147,N_26091);
nand U26282 (N_26282,N_26228,N_26211);
xnor U26283 (N_26283,N_26056,N_26114);
and U26284 (N_26284,N_26090,N_26244);
or U26285 (N_26285,N_26053,N_26076);
or U26286 (N_26286,N_26062,N_26115);
xor U26287 (N_26287,N_26117,N_26225);
xor U26288 (N_26288,N_26163,N_26026);
nand U26289 (N_26289,N_26212,N_26164);
nor U26290 (N_26290,N_26097,N_26236);
nor U26291 (N_26291,N_26065,N_26204);
and U26292 (N_26292,N_26224,N_26035);
nand U26293 (N_26293,N_26092,N_26189);
nor U26294 (N_26294,N_26184,N_26051);
or U26295 (N_26295,N_26177,N_26126);
and U26296 (N_26296,N_26046,N_26081);
nand U26297 (N_26297,N_26140,N_26181);
xor U26298 (N_26298,N_26116,N_26219);
xnor U26299 (N_26299,N_26106,N_26038);
xor U26300 (N_26300,N_26242,N_26198);
and U26301 (N_26301,N_26144,N_26063);
nand U26302 (N_26302,N_26043,N_26052);
nand U26303 (N_26303,N_26176,N_26192);
or U26304 (N_26304,N_26136,N_26206);
nor U26305 (N_26305,N_26196,N_26112);
xnor U26306 (N_26306,N_26025,N_26216);
nor U26307 (N_26307,N_26071,N_26175);
or U26308 (N_26308,N_26166,N_26032);
and U26309 (N_26309,N_26087,N_26001);
or U26310 (N_26310,N_26146,N_26127);
xnor U26311 (N_26311,N_26019,N_26202);
xnor U26312 (N_26312,N_26149,N_26179);
and U26313 (N_26313,N_26137,N_26217);
nor U26314 (N_26314,N_26180,N_26105);
nor U26315 (N_26315,N_26145,N_26134);
nand U26316 (N_26316,N_26034,N_26133);
and U26317 (N_26317,N_26067,N_26012);
xnor U26318 (N_26318,N_26013,N_26080);
and U26319 (N_26319,N_26155,N_26088);
or U26320 (N_26320,N_26135,N_26213);
and U26321 (N_26321,N_26110,N_26069);
nand U26322 (N_26322,N_26113,N_26186);
nand U26323 (N_26323,N_26078,N_26004);
xor U26324 (N_26324,N_26011,N_26099);
and U26325 (N_26325,N_26108,N_26058);
xor U26326 (N_26326,N_26083,N_26124);
and U26327 (N_26327,N_26129,N_26057);
nand U26328 (N_26328,N_26094,N_26243);
nor U26329 (N_26329,N_26003,N_26160);
or U26330 (N_26330,N_26104,N_26205);
and U26331 (N_26331,N_26241,N_26130);
and U26332 (N_26332,N_26230,N_26154);
xnor U26333 (N_26333,N_26054,N_26170);
nor U26334 (N_26334,N_26075,N_26018);
nor U26335 (N_26335,N_26239,N_26237);
xor U26336 (N_26336,N_26123,N_26208);
and U26337 (N_26337,N_26048,N_26148);
nor U26338 (N_26338,N_26121,N_26207);
nor U26339 (N_26339,N_26232,N_26015);
and U26340 (N_26340,N_26014,N_26008);
xnor U26341 (N_26341,N_26022,N_26070);
and U26342 (N_26342,N_26098,N_26096);
xor U26343 (N_26343,N_26200,N_26031);
nand U26344 (N_26344,N_26169,N_26142);
nor U26345 (N_26345,N_26002,N_26191);
and U26346 (N_26346,N_26139,N_26021);
nand U26347 (N_26347,N_26082,N_26132);
and U26348 (N_26348,N_26016,N_26068);
or U26349 (N_26349,N_26055,N_26235);
or U26350 (N_26350,N_26061,N_26005);
nand U26351 (N_26351,N_26073,N_26009);
xor U26352 (N_26352,N_26218,N_26100);
nand U26353 (N_26353,N_26033,N_26037);
or U26354 (N_26354,N_26221,N_26193);
nor U26355 (N_26355,N_26194,N_26171);
nor U26356 (N_26356,N_26039,N_26040);
nor U26357 (N_26357,N_26103,N_26238);
nor U26358 (N_26358,N_26143,N_26172);
and U26359 (N_26359,N_26178,N_26234);
nor U26360 (N_26360,N_26210,N_26245);
xor U26361 (N_26361,N_26084,N_26125);
nand U26362 (N_26362,N_26165,N_26215);
and U26363 (N_26363,N_26233,N_26050);
xnor U26364 (N_26364,N_26168,N_26060);
or U26365 (N_26365,N_26020,N_26151);
or U26366 (N_26366,N_26006,N_26086);
or U26367 (N_26367,N_26248,N_26041);
xnor U26368 (N_26368,N_26199,N_26074);
and U26369 (N_26369,N_26220,N_26131);
nor U26370 (N_26370,N_26085,N_26161);
and U26371 (N_26371,N_26102,N_26122);
nand U26372 (N_26372,N_26156,N_26119);
or U26373 (N_26373,N_26028,N_26231);
nor U26374 (N_26374,N_26023,N_26079);
nor U26375 (N_26375,N_26150,N_26147);
or U26376 (N_26376,N_26062,N_26184);
xor U26377 (N_26377,N_26203,N_26006);
or U26378 (N_26378,N_26150,N_26008);
nand U26379 (N_26379,N_26154,N_26011);
nand U26380 (N_26380,N_26040,N_26046);
and U26381 (N_26381,N_26090,N_26070);
or U26382 (N_26382,N_26017,N_26042);
or U26383 (N_26383,N_26074,N_26219);
and U26384 (N_26384,N_26070,N_26071);
or U26385 (N_26385,N_26055,N_26022);
and U26386 (N_26386,N_26098,N_26088);
or U26387 (N_26387,N_26248,N_26114);
and U26388 (N_26388,N_26198,N_26231);
and U26389 (N_26389,N_26097,N_26113);
nand U26390 (N_26390,N_26156,N_26035);
and U26391 (N_26391,N_26185,N_26069);
or U26392 (N_26392,N_26071,N_26147);
or U26393 (N_26393,N_26196,N_26119);
and U26394 (N_26394,N_26044,N_26031);
nand U26395 (N_26395,N_26163,N_26142);
or U26396 (N_26396,N_26076,N_26197);
nor U26397 (N_26397,N_26165,N_26205);
and U26398 (N_26398,N_26184,N_26128);
nor U26399 (N_26399,N_26130,N_26168);
and U26400 (N_26400,N_26157,N_26190);
nor U26401 (N_26401,N_26033,N_26002);
or U26402 (N_26402,N_26111,N_26086);
or U26403 (N_26403,N_26006,N_26039);
and U26404 (N_26404,N_26188,N_26097);
and U26405 (N_26405,N_26139,N_26053);
nand U26406 (N_26406,N_26041,N_26175);
nor U26407 (N_26407,N_26174,N_26154);
or U26408 (N_26408,N_26040,N_26164);
nor U26409 (N_26409,N_26138,N_26201);
xnor U26410 (N_26410,N_26202,N_26129);
and U26411 (N_26411,N_26180,N_26109);
nand U26412 (N_26412,N_26184,N_26109);
xnor U26413 (N_26413,N_26137,N_26140);
xnor U26414 (N_26414,N_26129,N_26021);
or U26415 (N_26415,N_26089,N_26065);
nor U26416 (N_26416,N_26181,N_26145);
or U26417 (N_26417,N_26022,N_26134);
or U26418 (N_26418,N_26024,N_26108);
xnor U26419 (N_26419,N_26196,N_26222);
and U26420 (N_26420,N_26229,N_26238);
and U26421 (N_26421,N_26245,N_26171);
nand U26422 (N_26422,N_26052,N_26204);
and U26423 (N_26423,N_26142,N_26134);
nand U26424 (N_26424,N_26017,N_26069);
nor U26425 (N_26425,N_26235,N_26101);
nor U26426 (N_26426,N_26229,N_26221);
xnor U26427 (N_26427,N_26108,N_26090);
nor U26428 (N_26428,N_26242,N_26209);
nor U26429 (N_26429,N_26013,N_26055);
and U26430 (N_26430,N_26103,N_26187);
nand U26431 (N_26431,N_26064,N_26044);
nor U26432 (N_26432,N_26140,N_26120);
and U26433 (N_26433,N_26190,N_26070);
and U26434 (N_26434,N_26093,N_26097);
or U26435 (N_26435,N_26001,N_26109);
xnor U26436 (N_26436,N_26220,N_26241);
or U26437 (N_26437,N_26142,N_26006);
and U26438 (N_26438,N_26079,N_26044);
xor U26439 (N_26439,N_26025,N_26195);
nor U26440 (N_26440,N_26177,N_26133);
nand U26441 (N_26441,N_26049,N_26050);
nor U26442 (N_26442,N_26053,N_26047);
and U26443 (N_26443,N_26216,N_26162);
and U26444 (N_26444,N_26247,N_26093);
nand U26445 (N_26445,N_26137,N_26034);
and U26446 (N_26446,N_26248,N_26002);
and U26447 (N_26447,N_26151,N_26141);
and U26448 (N_26448,N_26022,N_26216);
xnor U26449 (N_26449,N_26187,N_26223);
xor U26450 (N_26450,N_26033,N_26235);
xnor U26451 (N_26451,N_26237,N_26176);
nand U26452 (N_26452,N_26199,N_26164);
or U26453 (N_26453,N_26223,N_26073);
and U26454 (N_26454,N_26207,N_26116);
nand U26455 (N_26455,N_26084,N_26070);
xnor U26456 (N_26456,N_26097,N_26062);
or U26457 (N_26457,N_26135,N_26001);
and U26458 (N_26458,N_26120,N_26247);
and U26459 (N_26459,N_26008,N_26124);
xnor U26460 (N_26460,N_26211,N_26090);
and U26461 (N_26461,N_26080,N_26090);
nor U26462 (N_26462,N_26026,N_26006);
nor U26463 (N_26463,N_26009,N_26209);
or U26464 (N_26464,N_26221,N_26144);
and U26465 (N_26465,N_26008,N_26201);
xnor U26466 (N_26466,N_26090,N_26100);
nor U26467 (N_26467,N_26003,N_26246);
nand U26468 (N_26468,N_26016,N_26235);
and U26469 (N_26469,N_26182,N_26003);
and U26470 (N_26470,N_26057,N_26201);
or U26471 (N_26471,N_26208,N_26071);
xor U26472 (N_26472,N_26191,N_26222);
nand U26473 (N_26473,N_26085,N_26063);
and U26474 (N_26474,N_26110,N_26099);
and U26475 (N_26475,N_26245,N_26021);
nor U26476 (N_26476,N_26081,N_26118);
nor U26477 (N_26477,N_26182,N_26122);
xor U26478 (N_26478,N_26005,N_26103);
or U26479 (N_26479,N_26010,N_26126);
nor U26480 (N_26480,N_26051,N_26002);
and U26481 (N_26481,N_26021,N_26061);
or U26482 (N_26482,N_26234,N_26149);
or U26483 (N_26483,N_26083,N_26068);
nor U26484 (N_26484,N_26132,N_26232);
xnor U26485 (N_26485,N_26038,N_26046);
and U26486 (N_26486,N_26098,N_26005);
nand U26487 (N_26487,N_26150,N_26194);
xnor U26488 (N_26488,N_26071,N_26033);
and U26489 (N_26489,N_26039,N_26232);
or U26490 (N_26490,N_26248,N_26145);
and U26491 (N_26491,N_26090,N_26046);
nand U26492 (N_26492,N_26200,N_26245);
nor U26493 (N_26493,N_26185,N_26057);
nand U26494 (N_26494,N_26171,N_26035);
or U26495 (N_26495,N_26067,N_26021);
and U26496 (N_26496,N_26125,N_26099);
or U26497 (N_26497,N_26210,N_26018);
xnor U26498 (N_26498,N_26208,N_26028);
xor U26499 (N_26499,N_26226,N_26163);
nand U26500 (N_26500,N_26294,N_26333);
nor U26501 (N_26501,N_26388,N_26390);
nand U26502 (N_26502,N_26356,N_26282);
or U26503 (N_26503,N_26331,N_26469);
nor U26504 (N_26504,N_26339,N_26461);
nor U26505 (N_26505,N_26369,N_26314);
nor U26506 (N_26506,N_26342,N_26481);
and U26507 (N_26507,N_26363,N_26269);
xnor U26508 (N_26508,N_26274,N_26465);
xor U26509 (N_26509,N_26328,N_26422);
nand U26510 (N_26510,N_26479,N_26425);
nor U26511 (N_26511,N_26478,N_26371);
xor U26512 (N_26512,N_26340,N_26301);
nand U26513 (N_26513,N_26399,N_26495);
xnor U26514 (N_26514,N_26493,N_26497);
xor U26515 (N_26515,N_26321,N_26401);
xor U26516 (N_26516,N_26262,N_26375);
nand U26517 (N_26517,N_26365,N_26421);
nand U26518 (N_26518,N_26451,N_26286);
nand U26519 (N_26519,N_26499,N_26473);
nand U26520 (N_26520,N_26487,N_26416);
xnor U26521 (N_26521,N_26475,N_26347);
and U26522 (N_26522,N_26440,N_26482);
nand U26523 (N_26523,N_26311,N_26443);
and U26524 (N_26524,N_26281,N_26251);
and U26525 (N_26525,N_26306,N_26455);
and U26526 (N_26526,N_26277,N_26368);
nor U26527 (N_26527,N_26472,N_26442);
xnor U26528 (N_26528,N_26403,N_26329);
or U26529 (N_26529,N_26305,N_26374);
nand U26530 (N_26530,N_26485,N_26322);
and U26531 (N_26531,N_26386,N_26407);
or U26532 (N_26532,N_26253,N_26480);
xnor U26533 (N_26533,N_26323,N_26438);
nor U26534 (N_26534,N_26373,N_26498);
nand U26535 (N_26535,N_26441,N_26255);
or U26536 (N_26536,N_26405,N_26418);
xor U26537 (N_26537,N_26477,N_26355);
and U26538 (N_26538,N_26275,N_26335);
and U26539 (N_26539,N_26467,N_26254);
or U26540 (N_26540,N_26488,N_26258);
nand U26541 (N_26541,N_26494,N_26291);
xor U26542 (N_26542,N_26423,N_26300);
or U26543 (N_26543,N_26400,N_26460);
nor U26544 (N_26544,N_26264,N_26332);
xnor U26545 (N_26545,N_26256,N_26476);
nor U26546 (N_26546,N_26378,N_26382);
nor U26547 (N_26547,N_26450,N_26344);
nor U26548 (N_26548,N_26336,N_26353);
and U26549 (N_26549,N_26325,N_26289);
and U26550 (N_26550,N_26268,N_26419);
or U26551 (N_26551,N_26470,N_26427);
nor U26552 (N_26552,N_26361,N_26439);
or U26553 (N_26553,N_26394,N_26430);
or U26554 (N_26554,N_26413,N_26297);
or U26555 (N_26555,N_26393,N_26313);
or U26556 (N_26556,N_26298,N_26257);
nand U26557 (N_26557,N_26428,N_26341);
nand U26558 (N_26558,N_26383,N_26452);
or U26559 (N_26559,N_26354,N_26272);
or U26560 (N_26560,N_26360,N_26446);
nor U26561 (N_26561,N_26259,N_26310);
nor U26562 (N_26562,N_26349,N_26327);
nand U26563 (N_26563,N_26395,N_26273);
xnor U26564 (N_26564,N_26402,N_26364);
xor U26565 (N_26565,N_26411,N_26424);
and U26566 (N_26566,N_26320,N_26486);
and U26567 (N_26567,N_26457,N_26397);
or U26568 (N_26568,N_26433,N_26389);
or U26569 (N_26569,N_26284,N_26276);
and U26570 (N_26570,N_26362,N_26449);
nor U26571 (N_26571,N_26448,N_26324);
and U26572 (N_26572,N_26287,N_26279);
xnor U26573 (N_26573,N_26444,N_26285);
nor U26574 (N_26574,N_26464,N_26316);
and U26575 (N_26575,N_26270,N_26415);
and U26576 (N_26576,N_26417,N_26263);
nand U26577 (N_26577,N_26358,N_26466);
xor U26578 (N_26578,N_26343,N_26437);
nor U26579 (N_26579,N_26379,N_26346);
and U26580 (N_26580,N_26459,N_26490);
and U26581 (N_26581,N_26456,N_26345);
nor U26582 (N_26582,N_26414,N_26408);
or U26583 (N_26583,N_26391,N_26376);
xnor U26584 (N_26584,N_26271,N_26319);
nor U26585 (N_26585,N_26283,N_26260);
and U26586 (N_26586,N_26392,N_26303);
nand U26587 (N_26587,N_26435,N_26410);
nand U26588 (N_26588,N_26445,N_26454);
and U26589 (N_26589,N_26484,N_26409);
nor U26590 (N_26590,N_26315,N_26492);
and U26591 (N_26591,N_26468,N_26267);
nand U26592 (N_26592,N_26398,N_26462);
nand U26593 (N_26593,N_26252,N_26337);
or U26594 (N_26594,N_26309,N_26302);
or U26595 (N_26595,N_26483,N_26385);
or U26596 (N_26596,N_26491,N_26463);
and U26597 (N_26597,N_26288,N_26278);
or U26598 (N_26598,N_26261,N_26292);
and U26599 (N_26599,N_26326,N_26359);
and U26600 (N_26600,N_26447,N_26295);
xor U26601 (N_26601,N_26250,N_26351);
nor U26602 (N_26602,N_26429,N_26366);
and U26603 (N_26603,N_26304,N_26265);
or U26604 (N_26604,N_26307,N_26384);
xor U26605 (N_26605,N_26404,N_26471);
xor U26606 (N_26606,N_26299,N_26431);
nand U26607 (N_26607,N_26330,N_26338);
or U26608 (N_26608,N_26318,N_26312);
xor U26609 (N_26609,N_26308,N_26489);
and U26610 (N_26610,N_26317,N_26387);
and U26611 (N_26611,N_26396,N_26357);
and U26612 (N_26612,N_26334,N_26496);
xor U26613 (N_26613,N_26426,N_26474);
nor U26614 (N_26614,N_26290,N_26412);
xnor U26615 (N_26615,N_26380,N_26432);
xnor U26616 (N_26616,N_26352,N_26434);
and U26617 (N_26617,N_26348,N_26381);
and U26618 (N_26618,N_26296,N_26372);
nor U26619 (N_26619,N_26406,N_26293);
nand U26620 (N_26620,N_26458,N_26350);
or U26621 (N_26621,N_26266,N_26420);
and U26622 (N_26622,N_26370,N_26436);
xnor U26623 (N_26623,N_26367,N_26280);
nand U26624 (N_26624,N_26377,N_26453);
nand U26625 (N_26625,N_26404,N_26434);
nor U26626 (N_26626,N_26366,N_26445);
and U26627 (N_26627,N_26475,N_26384);
or U26628 (N_26628,N_26437,N_26368);
xor U26629 (N_26629,N_26334,N_26324);
and U26630 (N_26630,N_26456,N_26426);
xor U26631 (N_26631,N_26300,N_26277);
or U26632 (N_26632,N_26421,N_26265);
and U26633 (N_26633,N_26299,N_26484);
or U26634 (N_26634,N_26295,N_26279);
xor U26635 (N_26635,N_26491,N_26455);
and U26636 (N_26636,N_26415,N_26284);
xnor U26637 (N_26637,N_26322,N_26282);
nand U26638 (N_26638,N_26479,N_26291);
nor U26639 (N_26639,N_26272,N_26299);
nand U26640 (N_26640,N_26394,N_26315);
or U26641 (N_26641,N_26273,N_26492);
nand U26642 (N_26642,N_26482,N_26273);
and U26643 (N_26643,N_26330,N_26272);
nand U26644 (N_26644,N_26279,N_26293);
nor U26645 (N_26645,N_26441,N_26444);
and U26646 (N_26646,N_26396,N_26322);
nand U26647 (N_26647,N_26382,N_26494);
xnor U26648 (N_26648,N_26452,N_26448);
xnor U26649 (N_26649,N_26325,N_26373);
nor U26650 (N_26650,N_26354,N_26497);
or U26651 (N_26651,N_26387,N_26298);
nand U26652 (N_26652,N_26357,N_26329);
nor U26653 (N_26653,N_26467,N_26269);
or U26654 (N_26654,N_26495,N_26338);
and U26655 (N_26655,N_26393,N_26272);
and U26656 (N_26656,N_26263,N_26472);
and U26657 (N_26657,N_26359,N_26471);
nor U26658 (N_26658,N_26411,N_26354);
xnor U26659 (N_26659,N_26305,N_26345);
and U26660 (N_26660,N_26370,N_26441);
or U26661 (N_26661,N_26426,N_26463);
xnor U26662 (N_26662,N_26383,N_26308);
xor U26663 (N_26663,N_26473,N_26250);
or U26664 (N_26664,N_26454,N_26306);
and U26665 (N_26665,N_26498,N_26353);
xnor U26666 (N_26666,N_26330,N_26434);
nand U26667 (N_26667,N_26405,N_26345);
or U26668 (N_26668,N_26298,N_26340);
and U26669 (N_26669,N_26426,N_26344);
nor U26670 (N_26670,N_26346,N_26454);
and U26671 (N_26671,N_26467,N_26371);
nand U26672 (N_26672,N_26461,N_26459);
and U26673 (N_26673,N_26470,N_26283);
nand U26674 (N_26674,N_26473,N_26306);
xnor U26675 (N_26675,N_26457,N_26371);
and U26676 (N_26676,N_26373,N_26379);
xor U26677 (N_26677,N_26307,N_26419);
nand U26678 (N_26678,N_26275,N_26364);
xor U26679 (N_26679,N_26302,N_26496);
or U26680 (N_26680,N_26391,N_26270);
and U26681 (N_26681,N_26479,N_26268);
nor U26682 (N_26682,N_26430,N_26434);
and U26683 (N_26683,N_26481,N_26476);
xnor U26684 (N_26684,N_26389,N_26325);
xor U26685 (N_26685,N_26447,N_26481);
nand U26686 (N_26686,N_26399,N_26345);
or U26687 (N_26687,N_26476,N_26271);
xnor U26688 (N_26688,N_26378,N_26269);
xnor U26689 (N_26689,N_26425,N_26477);
or U26690 (N_26690,N_26275,N_26399);
xor U26691 (N_26691,N_26472,N_26302);
and U26692 (N_26692,N_26288,N_26390);
or U26693 (N_26693,N_26308,N_26296);
or U26694 (N_26694,N_26378,N_26270);
xnor U26695 (N_26695,N_26406,N_26331);
xor U26696 (N_26696,N_26464,N_26251);
nand U26697 (N_26697,N_26408,N_26283);
nand U26698 (N_26698,N_26423,N_26461);
xor U26699 (N_26699,N_26283,N_26447);
xor U26700 (N_26700,N_26430,N_26263);
and U26701 (N_26701,N_26496,N_26438);
and U26702 (N_26702,N_26272,N_26388);
or U26703 (N_26703,N_26458,N_26452);
and U26704 (N_26704,N_26385,N_26373);
and U26705 (N_26705,N_26265,N_26287);
nand U26706 (N_26706,N_26408,N_26456);
and U26707 (N_26707,N_26407,N_26290);
nand U26708 (N_26708,N_26389,N_26384);
or U26709 (N_26709,N_26482,N_26299);
nor U26710 (N_26710,N_26281,N_26252);
nor U26711 (N_26711,N_26479,N_26279);
xnor U26712 (N_26712,N_26314,N_26266);
xnor U26713 (N_26713,N_26401,N_26379);
xnor U26714 (N_26714,N_26330,N_26310);
or U26715 (N_26715,N_26346,N_26263);
and U26716 (N_26716,N_26293,N_26375);
nor U26717 (N_26717,N_26359,N_26438);
nor U26718 (N_26718,N_26441,N_26266);
nand U26719 (N_26719,N_26337,N_26265);
nand U26720 (N_26720,N_26322,N_26441);
nor U26721 (N_26721,N_26474,N_26425);
xnor U26722 (N_26722,N_26350,N_26262);
nor U26723 (N_26723,N_26316,N_26386);
xor U26724 (N_26724,N_26308,N_26445);
xnor U26725 (N_26725,N_26450,N_26491);
nand U26726 (N_26726,N_26357,N_26279);
nand U26727 (N_26727,N_26352,N_26487);
xor U26728 (N_26728,N_26279,N_26419);
and U26729 (N_26729,N_26450,N_26374);
and U26730 (N_26730,N_26262,N_26357);
or U26731 (N_26731,N_26339,N_26295);
xnor U26732 (N_26732,N_26362,N_26460);
xor U26733 (N_26733,N_26491,N_26355);
and U26734 (N_26734,N_26282,N_26402);
and U26735 (N_26735,N_26356,N_26348);
and U26736 (N_26736,N_26445,N_26411);
nand U26737 (N_26737,N_26395,N_26442);
xor U26738 (N_26738,N_26261,N_26368);
nor U26739 (N_26739,N_26304,N_26477);
xor U26740 (N_26740,N_26456,N_26370);
nor U26741 (N_26741,N_26498,N_26411);
or U26742 (N_26742,N_26263,N_26403);
xnor U26743 (N_26743,N_26378,N_26485);
xor U26744 (N_26744,N_26349,N_26398);
xnor U26745 (N_26745,N_26499,N_26350);
and U26746 (N_26746,N_26335,N_26311);
xor U26747 (N_26747,N_26268,N_26440);
or U26748 (N_26748,N_26302,N_26263);
xor U26749 (N_26749,N_26339,N_26485);
or U26750 (N_26750,N_26617,N_26525);
or U26751 (N_26751,N_26744,N_26508);
and U26752 (N_26752,N_26502,N_26602);
or U26753 (N_26753,N_26505,N_26665);
xnor U26754 (N_26754,N_26741,N_26703);
nand U26755 (N_26755,N_26664,N_26714);
and U26756 (N_26756,N_26728,N_26524);
nor U26757 (N_26757,N_26645,N_26609);
xnor U26758 (N_26758,N_26635,N_26732);
xor U26759 (N_26759,N_26712,N_26662);
xor U26760 (N_26760,N_26667,N_26646);
and U26761 (N_26761,N_26700,N_26581);
nand U26762 (N_26762,N_26641,N_26650);
and U26763 (N_26763,N_26659,N_26556);
and U26764 (N_26764,N_26591,N_26637);
and U26765 (N_26765,N_26518,N_26716);
and U26766 (N_26766,N_26632,N_26739);
xor U26767 (N_26767,N_26653,N_26689);
nor U26768 (N_26768,N_26674,N_26707);
xnor U26769 (N_26769,N_26742,N_26672);
nor U26770 (N_26770,N_26542,N_26569);
xnor U26771 (N_26771,N_26663,N_26532);
or U26772 (N_26772,N_26746,N_26634);
and U26773 (N_26773,N_26629,N_26511);
nor U26774 (N_26774,N_26683,N_26509);
xnor U26775 (N_26775,N_26638,N_26530);
xor U26776 (N_26776,N_26579,N_26610);
nor U26777 (N_26777,N_26685,N_26584);
and U26778 (N_26778,N_26574,N_26737);
nand U26779 (N_26779,N_26592,N_26690);
and U26780 (N_26780,N_26708,N_26553);
xnor U26781 (N_26781,N_26723,N_26506);
or U26782 (N_26782,N_26595,N_26545);
xnor U26783 (N_26783,N_26531,N_26538);
or U26784 (N_26784,N_26567,N_26673);
and U26785 (N_26785,N_26533,N_26586);
and U26786 (N_26786,N_26697,N_26701);
nor U26787 (N_26787,N_26516,N_26604);
xor U26788 (N_26788,N_26546,N_26601);
or U26789 (N_26789,N_26588,N_26564);
or U26790 (N_26790,N_26565,N_26523);
and U26791 (N_26791,N_26717,N_26513);
or U26792 (N_26792,N_26563,N_26749);
xnor U26793 (N_26793,N_26585,N_26668);
and U26794 (N_26794,N_26642,N_26711);
nor U26795 (N_26795,N_26576,N_26593);
xnor U26796 (N_26796,N_26608,N_26702);
or U26797 (N_26797,N_26643,N_26692);
and U26798 (N_26798,N_26639,N_26544);
xnor U26799 (N_26799,N_26649,N_26693);
and U26800 (N_26800,N_26729,N_26730);
or U26801 (N_26801,N_26535,N_26679);
nor U26802 (N_26802,N_26687,N_26706);
nor U26803 (N_26803,N_26521,N_26626);
xnor U26804 (N_26804,N_26627,N_26677);
xnor U26805 (N_26805,N_26636,N_26630);
xor U26806 (N_26806,N_26731,N_26724);
and U26807 (N_26807,N_26612,N_26589);
nor U26808 (N_26808,N_26587,N_26590);
or U26809 (N_26809,N_26503,N_26644);
nor U26810 (N_26810,N_26621,N_26721);
xnor U26811 (N_26811,N_26705,N_26522);
and U26812 (N_26812,N_26571,N_26615);
xnor U26813 (N_26813,N_26596,N_26657);
and U26814 (N_26814,N_26540,N_26572);
or U26815 (N_26815,N_26566,N_26560);
and U26816 (N_26816,N_26552,N_26620);
or U26817 (N_26817,N_26558,N_26583);
nor U26818 (N_26818,N_26678,N_26651);
and U26819 (N_26819,N_26570,N_26512);
or U26820 (N_26820,N_26733,N_26594);
or U26821 (N_26821,N_26537,N_26656);
nor U26822 (N_26822,N_26725,N_26534);
nand U26823 (N_26823,N_26727,N_26557);
or U26824 (N_26824,N_26600,N_26682);
nor U26825 (N_26825,N_26688,N_26676);
nor U26826 (N_26826,N_26666,N_26625);
nand U26827 (N_26827,N_26658,N_26536);
xnor U26828 (N_26828,N_26517,N_26623);
xnor U26829 (N_26829,N_26691,N_26541);
and U26830 (N_26830,N_26514,N_26501);
and U26831 (N_26831,N_26554,N_26680);
or U26832 (N_26832,N_26510,N_26709);
xor U26833 (N_26833,N_26527,N_26736);
or U26834 (N_26834,N_26622,N_26713);
nor U26835 (N_26835,N_26580,N_26726);
nand U26836 (N_26836,N_26597,N_26548);
xnor U26837 (N_26837,N_26743,N_26599);
nand U26838 (N_26838,N_26740,N_26628);
and U26839 (N_26839,N_26647,N_26515);
nor U26840 (N_26840,N_26507,N_26555);
nor U26841 (N_26841,N_26547,N_26652);
nand U26842 (N_26842,N_26520,N_26539);
nand U26843 (N_26843,N_26519,N_26578);
and U26844 (N_26844,N_26607,N_26562);
xnor U26845 (N_26845,N_26543,N_26661);
nor U26846 (N_26846,N_26734,N_26698);
nor U26847 (N_26847,N_26738,N_26718);
xnor U26848 (N_26848,N_26670,N_26695);
nor U26849 (N_26849,N_26660,N_26550);
or U26850 (N_26850,N_26616,N_26526);
nand U26851 (N_26851,N_26722,N_26719);
or U26852 (N_26852,N_26624,N_26748);
nand U26853 (N_26853,N_26747,N_26582);
or U26854 (N_26854,N_26575,N_26648);
or U26855 (N_26855,N_26603,N_26675);
xnor U26856 (N_26856,N_26669,N_26671);
nor U26857 (N_26857,N_26619,N_26500);
nor U26858 (N_26858,N_26745,N_26614);
and U26859 (N_26859,N_26529,N_26577);
nand U26860 (N_26860,N_26720,N_26598);
nor U26861 (N_26861,N_26654,N_26561);
nand U26862 (N_26862,N_26696,N_26694);
and U26863 (N_26863,N_26613,N_26605);
nand U26864 (N_26864,N_26633,N_26504);
nor U26865 (N_26865,N_26684,N_26611);
xor U26866 (N_26866,N_26528,N_26686);
and U26867 (N_26867,N_26681,N_26573);
xor U26868 (N_26868,N_26735,N_26715);
nand U26869 (N_26869,N_26618,N_26631);
and U26870 (N_26870,N_26551,N_26655);
nor U26871 (N_26871,N_26559,N_26704);
xnor U26872 (N_26872,N_26710,N_26549);
xnor U26873 (N_26873,N_26568,N_26699);
or U26874 (N_26874,N_26606,N_26640);
or U26875 (N_26875,N_26653,N_26733);
and U26876 (N_26876,N_26741,N_26748);
nand U26877 (N_26877,N_26566,N_26675);
nand U26878 (N_26878,N_26641,N_26575);
nand U26879 (N_26879,N_26732,N_26690);
and U26880 (N_26880,N_26571,N_26624);
nand U26881 (N_26881,N_26526,N_26675);
or U26882 (N_26882,N_26665,N_26637);
xor U26883 (N_26883,N_26566,N_26643);
nand U26884 (N_26884,N_26582,N_26657);
nor U26885 (N_26885,N_26582,N_26561);
xor U26886 (N_26886,N_26740,N_26721);
xor U26887 (N_26887,N_26638,N_26639);
nand U26888 (N_26888,N_26611,N_26592);
nor U26889 (N_26889,N_26558,N_26598);
xnor U26890 (N_26890,N_26649,N_26705);
nor U26891 (N_26891,N_26738,N_26586);
nor U26892 (N_26892,N_26725,N_26586);
nor U26893 (N_26893,N_26674,N_26578);
nor U26894 (N_26894,N_26561,N_26670);
nand U26895 (N_26895,N_26725,N_26532);
nand U26896 (N_26896,N_26568,N_26527);
xor U26897 (N_26897,N_26722,N_26554);
nor U26898 (N_26898,N_26554,N_26687);
or U26899 (N_26899,N_26638,N_26550);
or U26900 (N_26900,N_26560,N_26624);
nor U26901 (N_26901,N_26570,N_26711);
nand U26902 (N_26902,N_26615,N_26702);
nand U26903 (N_26903,N_26746,N_26607);
nand U26904 (N_26904,N_26524,N_26629);
xor U26905 (N_26905,N_26731,N_26734);
or U26906 (N_26906,N_26569,N_26568);
nand U26907 (N_26907,N_26683,N_26560);
nor U26908 (N_26908,N_26615,N_26714);
or U26909 (N_26909,N_26591,N_26729);
nand U26910 (N_26910,N_26642,N_26634);
or U26911 (N_26911,N_26506,N_26517);
nand U26912 (N_26912,N_26515,N_26520);
nand U26913 (N_26913,N_26586,N_26677);
xnor U26914 (N_26914,N_26581,N_26509);
and U26915 (N_26915,N_26697,N_26733);
nor U26916 (N_26916,N_26530,N_26720);
and U26917 (N_26917,N_26700,N_26618);
xor U26918 (N_26918,N_26671,N_26733);
xor U26919 (N_26919,N_26606,N_26594);
nor U26920 (N_26920,N_26526,N_26678);
xnor U26921 (N_26921,N_26732,N_26550);
or U26922 (N_26922,N_26510,N_26670);
nand U26923 (N_26923,N_26733,N_26672);
nor U26924 (N_26924,N_26559,N_26522);
xor U26925 (N_26925,N_26714,N_26745);
xor U26926 (N_26926,N_26725,N_26707);
and U26927 (N_26927,N_26738,N_26500);
xor U26928 (N_26928,N_26514,N_26673);
nor U26929 (N_26929,N_26635,N_26537);
nand U26930 (N_26930,N_26643,N_26572);
xnor U26931 (N_26931,N_26581,N_26726);
xor U26932 (N_26932,N_26658,N_26593);
and U26933 (N_26933,N_26744,N_26716);
nor U26934 (N_26934,N_26621,N_26545);
xor U26935 (N_26935,N_26691,N_26674);
or U26936 (N_26936,N_26742,N_26567);
xnor U26937 (N_26937,N_26564,N_26672);
xnor U26938 (N_26938,N_26515,N_26671);
and U26939 (N_26939,N_26658,N_26671);
nor U26940 (N_26940,N_26634,N_26695);
nor U26941 (N_26941,N_26548,N_26602);
nand U26942 (N_26942,N_26561,N_26645);
xor U26943 (N_26943,N_26588,N_26583);
nor U26944 (N_26944,N_26718,N_26712);
xor U26945 (N_26945,N_26676,N_26592);
or U26946 (N_26946,N_26680,N_26514);
nand U26947 (N_26947,N_26547,N_26556);
or U26948 (N_26948,N_26735,N_26555);
xnor U26949 (N_26949,N_26604,N_26698);
xor U26950 (N_26950,N_26698,N_26507);
or U26951 (N_26951,N_26665,N_26627);
nand U26952 (N_26952,N_26693,N_26643);
nor U26953 (N_26953,N_26611,N_26735);
or U26954 (N_26954,N_26519,N_26677);
xor U26955 (N_26955,N_26666,N_26513);
or U26956 (N_26956,N_26591,N_26576);
nand U26957 (N_26957,N_26507,N_26534);
and U26958 (N_26958,N_26654,N_26525);
nor U26959 (N_26959,N_26748,N_26644);
nand U26960 (N_26960,N_26500,N_26588);
and U26961 (N_26961,N_26595,N_26531);
nand U26962 (N_26962,N_26713,N_26740);
or U26963 (N_26963,N_26502,N_26609);
nor U26964 (N_26964,N_26525,N_26662);
xnor U26965 (N_26965,N_26666,N_26576);
xor U26966 (N_26966,N_26677,N_26550);
xor U26967 (N_26967,N_26669,N_26632);
nand U26968 (N_26968,N_26521,N_26730);
or U26969 (N_26969,N_26520,N_26714);
xnor U26970 (N_26970,N_26711,N_26691);
nand U26971 (N_26971,N_26708,N_26726);
and U26972 (N_26972,N_26720,N_26653);
and U26973 (N_26973,N_26637,N_26612);
nand U26974 (N_26974,N_26504,N_26718);
nor U26975 (N_26975,N_26612,N_26621);
or U26976 (N_26976,N_26562,N_26621);
and U26977 (N_26977,N_26721,N_26567);
or U26978 (N_26978,N_26572,N_26626);
and U26979 (N_26979,N_26601,N_26514);
and U26980 (N_26980,N_26560,N_26606);
nor U26981 (N_26981,N_26502,N_26717);
and U26982 (N_26982,N_26555,N_26619);
nor U26983 (N_26983,N_26678,N_26705);
xor U26984 (N_26984,N_26741,N_26516);
nor U26985 (N_26985,N_26728,N_26511);
or U26986 (N_26986,N_26640,N_26646);
or U26987 (N_26987,N_26601,N_26561);
nand U26988 (N_26988,N_26620,N_26574);
or U26989 (N_26989,N_26740,N_26532);
and U26990 (N_26990,N_26558,N_26690);
nand U26991 (N_26991,N_26737,N_26599);
nand U26992 (N_26992,N_26618,N_26702);
and U26993 (N_26993,N_26721,N_26611);
nor U26994 (N_26994,N_26523,N_26607);
xor U26995 (N_26995,N_26739,N_26592);
nand U26996 (N_26996,N_26609,N_26691);
nor U26997 (N_26997,N_26602,N_26729);
xnor U26998 (N_26998,N_26595,N_26652);
xnor U26999 (N_26999,N_26727,N_26721);
and U27000 (N_27000,N_26783,N_26826);
or U27001 (N_27001,N_26863,N_26838);
or U27002 (N_27002,N_26792,N_26823);
xnor U27003 (N_27003,N_26868,N_26989);
or U27004 (N_27004,N_26885,N_26836);
or U27005 (N_27005,N_26846,N_26842);
xnor U27006 (N_27006,N_26858,N_26897);
xnor U27007 (N_27007,N_26948,N_26793);
xor U27008 (N_27008,N_26772,N_26787);
xnor U27009 (N_27009,N_26961,N_26788);
xor U27010 (N_27010,N_26796,N_26778);
or U27011 (N_27011,N_26827,N_26881);
nand U27012 (N_27012,N_26790,N_26845);
nor U27013 (N_27013,N_26806,N_26862);
or U27014 (N_27014,N_26817,N_26883);
nand U27015 (N_27015,N_26913,N_26887);
nand U27016 (N_27016,N_26981,N_26857);
xnor U27017 (N_27017,N_26960,N_26946);
xor U27018 (N_27018,N_26853,N_26821);
and U27019 (N_27019,N_26894,N_26751);
nand U27020 (N_27020,N_26971,N_26917);
and U27021 (N_27021,N_26794,N_26910);
and U27022 (N_27022,N_26799,N_26819);
and U27023 (N_27023,N_26770,N_26983);
nor U27024 (N_27024,N_26984,N_26802);
xor U27025 (N_27025,N_26810,N_26861);
and U27026 (N_27026,N_26992,N_26972);
xnor U27027 (N_27027,N_26963,N_26764);
xnor U27028 (N_27028,N_26822,N_26976);
xnor U27029 (N_27029,N_26965,N_26878);
or U27030 (N_27030,N_26974,N_26997);
or U27031 (N_27031,N_26982,N_26918);
nor U27032 (N_27032,N_26791,N_26988);
nor U27033 (N_27033,N_26860,N_26904);
or U27034 (N_27034,N_26767,N_26801);
xnor U27035 (N_27035,N_26927,N_26760);
and U27036 (N_27036,N_26835,N_26933);
nor U27037 (N_27037,N_26815,N_26876);
nor U27038 (N_27038,N_26763,N_26759);
nand U27039 (N_27039,N_26813,N_26816);
nand U27040 (N_27040,N_26884,N_26985);
nor U27041 (N_27041,N_26930,N_26964);
or U27042 (N_27042,N_26777,N_26951);
nand U27043 (N_27043,N_26761,N_26755);
nor U27044 (N_27044,N_26756,N_26766);
nand U27045 (N_27045,N_26784,N_26758);
nor U27046 (N_27046,N_26824,N_26837);
nor U27047 (N_27047,N_26786,N_26956);
nand U27048 (N_27048,N_26891,N_26780);
nand U27049 (N_27049,N_26768,N_26914);
nor U27050 (N_27050,N_26993,N_26898);
and U27051 (N_27051,N_26803,N_26915);
nand U27052 (N_27052,N_26925,N_26829);
and U27053 (N_27053,N_26966,N_26931);
nand U27054 (N_27054,N_26909,N_26926);
and U27055 (N_27055,N_26944,N_26991);
xor U27056 (N_27056,N_26832,N_26916);
nand U27057 (N_27057,N_26875,N_26773);
xnor U27058 (N_27058,N_26919,N_26874);
or U27059 (N_27059,N_26980,N_26882);
nor U27060 (N_27060,N_26762,N_26908);
nand U27061 (N_27061,N_26830,N_26978);
nor U27062 (N_27062,N_26812,N_26831);
nand U27063 (N_27063,N_26934,N_26949);
and U27064 (N_27064,N_26940,N_26912);
xnor U27065 (N_27065,N_26929,N_26871);
or U27066 (N_27066,N_26795,N_26844);
and U27067 (N_27067,N_26945,N_26798);
xor U27068 (N_27068,N_26892,N_26809);
and U27069 (N_27069,N_26888,N_26754);
and U27070 (N_27070,N_26952,N_26872);
xnor U27071 (N_27071,N_26779,N_26865);
nand U27072 (N_27072,N_26957,N_26805);
or U27073 (N_27073,N_26828,N_26833);
nand U27074 (N_27074,N_26859,N_26849);
or U27075 (N_27075,N_26851,N_26870);
or U27076 (N_27076,N_26975,N_26750);
nor U27077 (N_27077,N_26848,N_26895);
or U27078 (N_27078,N_26811,N_26901);
nor U27079 (N_27079,N_26911,N_26947);
nand U27080 (N_27080,N_26995,N_26843);
and U27081 (N_27081,N_26970,N_26825);
or U27082 (N_27082,N_26757,N_26869);
nor U27083 (N_27083,N_26800,N_26864);
nor U27084 (N_27084,N_26998,N_26903);
and U27085 (N_27085,N_26937,N_26866);
and U27086 (N_27086,N_26797,N_26775);
and U27087 (N_27087,N_26873,N_26808);
nand U27088 (N_27088,N_26880,N_26990);
nand U27089 (N_27089,N_26774,N_26932);
and U27090 (N_27090,N_26820,N_26906);
and U27091 (N_27091,N_26924,N_26855);
nand U27092 (N_27092,N_26852,N_26785);
nor U27093 (N_27093,N_26789,N_26905);
or U27094 (N_27094,N_26781,N_26896);
and U27095 (N_27095,N_26955,N_26839);
and U27096 (N_27096,N_26804,N_26753);
or U27097 (N_27097,N_26907,N_26938);
or U27098 (N_27098,N_26877,N_26850);
nand U27099 (N_27099,N_26943,N_26935);
and U27100 (N_27100,N_26967,N_26886);
nand U27101 (N_27101,N_26818,N_26986);
xnor U27102 (N_27102,N_26902,N_26889);
nor U27103 (N_27103,N_26941,N_26893);
or U27104 (N_27104,N_26900,N_26994);
xnor U27105 (N_27105,N_26939,N_26953);
nor U27106 (N_27106,N_26807,N_26856);
nor U27107 (N_27107,N_26847,N_26841);
nand U27108 (N_27108,N_26840,N_26834);
and U27109 (N_27109,N_26867,N_26928);
and U27110 (N_27110,N_26969,N_26999);
or U27111 (N_27111,N_26950,N_26765);
xor U27112 (N_27112,N_26769,N_26922);
xor U27113 (N_27113,N_26954,N_26959);
nand U27114 (N_27114,N_26987,N_26920);
xnor U27115 (N_27115,N_26782,N_26776);
nand U27116 (N_27116,N_26771,N_26977);
or U27117 (N_27117,N_26979,N_26958);
nor U27118 (N_27118,N_26890,N_26814);
or U27119 (N_27119,N_26996,N_26879);
nor U27120 (N_27120,N_26854,N_26899);
xor U27121 (N_27121,N_26923,N_26942);
nor U27122 (N_27122,N_26973,N_26962);
and U27123 (N_27123,N_26752,N_26936);
and U27124 (N_27124,N_26968,N_26921);
nor U27125 (N_27125,N_26790,N_26863);
xor U27126 (N_27126,N_26932,N_26897);
nand U27127 (N_27127,N_26953,N_26980);
nor U27128 (N_27128,N_26796,N_26892);
or U27129 (N_27129,N_26941,N_26898);
and U27130 (N_27130,N_26862,N_26838);
nand U27131 (N_27131,N_26998,N_26755);
nand U27132 (N_27132,N_26959,N_26808);
and U27133 (N_27133,N_26875,N_26825);
nor U27134 (N_27134,N_26834,N_26782);
xnor U27135 (N_27135,N_26897,N_26871);
nor U27136 (N_27136,N_26792,N_26787);
or U27137 (N_27137,N_26837,N_26896);
nand U27138 (N_27138,N_26868,N_26819);
nor U27139 (N_27139,N_26813,N_26852);
nor U27140 (N_27140,N_26985,N_26766);
or U27141 (N_27141,N_26830,N_26894);
nand U27142 (N_27142,N_26987,N_26857);
or U27143 (N_27143,N_26838,N_26920);
nor U27144 (N_27144,N_26850,N_26849);
nor U27145 (N_27145,N_26773,N_26802);
nand U27146 (N_27146,N_26797,N_26951);
xnor U27147 (N_27147,N_26939,N_26929);
or U27148 (N_27148,N_26977,N_26941);
nor U27149 (N_27149,N_26877,N_26900);
and U27150 (N_27150,N_26906,N_26931);
xor U27151 (N_27151,N_26861,N_26763);
and U27152 (N_27152,N_26872,N_26914);
xor U27153 (N_27153,N_26913,N_26809);
or U27154 (N_27154,N_26769,N_26775);
xor U27155 (N_27155,N_26855,N_26993);
and U27156 (N_27156,N_26905,N_26837);
nand U27157 (N_27157,N_26768,N_26987);
and U27158 (N_27158,N_26972,N_26911);
or U27159 (N_27159,N_26959,N_26847);
xnor U27160 (N_27160,N_26937,N_26786);
or U27161 (N_27161,N_26916,N_26936);
xnor U27162 (N_27162,N_26874,N_26779);
nor U27163 (N_27163,N_26995,N_26943);
nor U27164 (N_27164,N_26790,N_26977);
xor U27165 (N_27165,N_26856,N_26834);
nand U27166 (N_27166,N_26903,N_26931);
or U27167 (N_27167,N_26857,N_26891);
nand U27168 (N_27168,N_26875,N_26902);
nand U27169 (N_27169,N_26783,N_26790);
and U27170 (N_27170,N_26801,N_26864);
or U27171 (N_27171,N_26972,N_26858);
nor U27172 (N_27172,N_26757,N_26837);
xor U27173 (N_27173,N_26973,N_26930);
and U27174 (N_27174,N_26967,N_26806);
nor U27175 (N_27175,N_26949,N_26890);
nand U27176 (N_27176,N_26896,N_26992);
nor U27177 (N_27177,N_26866,N_26918);
or U27178 (N_27178,N_26791,N_26867);
nor U27179 (N_27179,N_26825,N_26819);
xnor U27180 (N_27180,N_26794,N_26895);
or U27181 (N_27181,N_26984,N_26834);
nor U27182 (N_27182,N_26823,N_26967);
and U27183 (N_27183,N_26942,N_26899);
xnor U27184 (N_27184,N_26774,N_26938);
and U27185 (N_27185,N_26915,N_26758);
xnor U27186 (N_27186,N_26912,N_26973);
nor U27187 (N_27187,N_26958,N_26925);
xnor U27188 (N_27188,N_26884,N_26859);
nand U27189 (N_27189,N_26841,N_26833);
and U27190 (N_27190,N_26817,N_26938);
and U27191 (N_27191,N_26971,N_26849);
or U27192 (N_27192,N_26789,N_26916);
nand U27193 (N_27193,N_26946,N_26951);
or U27194 (N_27194,N_26915,N_26904);
nor U27195 (N_27195,N_26934,N_26877);
nand U27196 (N_27196,N_26750,N_26973);
or U27197 (N_27197,N_26968,N_26759);
or U27198 (N_27198,N_26803,N_26966);
and U27199 (N_27199,N_26756,N_26988);
and U27200 (N_27200,N_26966,N_26946);
nand U27201 (N_27201,N_26779,N_26760);
and U27202 (N_27202,N_26773,N_26956);
nor U27203 (N_27203,N_26963,N_26796);
nor U27204 (N_27204,N_26889,N_26993);
nand U27205 (N_27205,N_26915,N_26808);
and U27206 (N_27206,N_26921,N_26897);
or U27207 (N_27207,N_26886,N_26963);
or U27208 (N_27208,N_26954,N_26853);
nor U27209 (N_27209,N_26827,N_26839);
nand U27210 (N_27210,N_26891,N_26843);
xor U27211 (N_27211,N_26870,N_26858);
xor U27212 (N_27212,N_26999,N_26850);
nand U27213 (N_27213,N_26779,N_26895);
nor U27214 (N_27214,N_26797,N_26771);
or U27215 (N_27215,N_26900,N_26842);
or U27216 (N_27216,N_26750,N_26926);
nand U27217 (N_27217,N_26820,N_26780);
and U27218 (N_27218,N_26880,N_26765);
xnor U27219 (N_27219,N_26914,N_26951);
and U27220 (N_27220,N_26803,N_26784);
nand U27221 (N_27221,N_26852,N_26948);
or U27222 (N_27222,N_26984,N_26862);
nand U27223 (N_27223,N_26856,N_26813);
nand U27224 (N_27224,N_26961,N_26825);
nor U27225 (N_27225,N_26880,N_26903);
and U27226 (N_27226,N_26975,N_26988);
nor U27227 (N_27227,N_26824,N_26828);
and U27228 (N_27228,N_26849,N_26861);
nand U27229 (N_27229,N_26821,N_26840);
nand U27230 (N_27230,N_26835,N_26942);
or U27231 (N_27231,N_26817,N_26859);
nand U27232 (N_27232,N_26877,N_26868);
xnor U27233 (N_27233,N_26907,N_26902);
or U27234 (N_27234,N_26775,N_26854);
and U27235 (N_27235,N_26795,N_26981);
xnor U27236 (N_27236,N_26792,N_26881);
and U27237 (N_27237,N_26954,N_26988);
nand U27238 (N_27238,N_26993,N_26776);
or U27239 (N_27239,N_26875,N_26895);
or U27240 (N_27240,N_26915,N_26762);
or U27241 (N_27241,N_26753,N_26787);
nor U27242 (N_27242,N_26770,N_26910);
or U27243 (N_27243,N_26772,N_26861);
nor U27244 (N_27244,N_26786,N_26929);
nor U27245 (N_27245,N_26899,N_26901);
nand U27246 (N_27246,N_26942,N_26844);
or U27247 (N_27247,N_26999,N_26845);
xor U27248 (N_27248,N_26961,N_26991);
xnor U27249 (N_27249,N_26820,N_26874);
or U27250 (N_27250,N_27166,N_27120);
nor U27251 (N_27251,N_27031,N_27129);
or U27252 (N_27252,N_27030,N_27176);
and U27253 (N_27253,N_27091,N_27192);
or U27254 (N_27254,N_27237,N_27130);
xor U27255 (N_27255,N_27184,N_27000);
xnor U27256 (N_27256,N_27137,N_27038);
or U27257 (N_27257,N_27169,N_27108);
nand U27258 (N_27258,N_27160,N_27238);
xnor U27259 (N_27259,N_27004,N_27001);
or U27260 (N_27260,N_27113,N_27118);
or U27261 (N_27261,N_27049,N_27249);
and U27262 (N_27262,N_27224,N_27021);
or U27263 (N_27263,N_27047,N_27051);
nor U27264 (N_27264,N_27082,N_27058);
or U27265 (N_27265,N_27102,N_27125);
nor U27266 (N_27266,N_27141,N_27189);
nor U27267 (N_27267,N_27167,N_27024);
xor U27268 (N_27268,N_27029,N_27046);
nand U27269 (N_27269,N_27225,N_27239);
or U27270 (N_27270,N_27101,N_27069);
nand U27271 (N_27271,N_27041,N_27213);
nor U27272 (N_27272,N_27203,N_27015);
xor U27273 (N_27273,N_27144,N_27119);
nand U27274 (N_27274,N_27035,N_27218);
nand U27275 (N_27275,N_27084,N_27171);
nand U27276 (N_27276,N_27116,N_27009);
nand U27277 (N_27277,N_27240,N_27052);
or U27278 (N_27278,N_27121,N_27020);
and U27279 (N_27279,N_27190,N_27164);
nand U27280 (N_27280,N_27180,N_27065);
nand U27281 (N_27281,N_27114,N_27241);
or U27282 (N_27282,N_27078,N_27017);
xor U27283 (N_27283,N_27221,N_27191);
nand U27284 (N_27284,N_27086,N_27011);
and U27285 (N_27285,N_27196,N_27093);
nor U27286 (N_27286,N_27138,N_27215);
nand U27287 (N_27287,N_27162,N_27083);
xnor U27288 (N_27288,N_27127,N_27103);
and U27289 (N_27289,N_27008,N_27076);
nand U27290 (N_27290,N_27195,N_27136);
nor U27291 (N_27291,N_27060,N_27112);
and U27292 (N_27292,N_27111,N_27064);
nor U27293 (N_27293,N_27036,N_27117);
nor U27294 (N_27294,N_27159,N_27068);
or U27295 (N_27295,N_27085,N_27207);
or U27296 (N_27296,N_27100,N_27227);
xor U27297 (N_27297,N_27134,N_27057);
nand U27298 (N_27298,N_27002,N_27095);
or U27299 (N_27299,N_27182,N_27204);
or U27300 (N_27300,N_27247,N_27080);
or U27301 (N_27301,N_27026,N_27006);
nand U27302 (N_27302,N_27188,N_27105);
xor U27303 (N_27303,N_27056,N_27124);
and U27304 (N_27304,N_27061,N_27214);
nand U27305 (N_27305,N_27220,N_27199);
or U27306 (N_27306,N_27205,N_27208);
xor U27307 (N_27307,N_27153,N_27151);
xnor U27308 (N_27308,N_27054,N_27206);
and U27309 (N_27309,N_27135,N_27132);
and U27310 (N_27310,N_27107,N_27194);
xnor U27311 (N_27311,N_27244,N_27200);
nand U27312 (N_27312,N_27071,N_27109);
nand U27313 (N_27313,N_27033,N_27094);
and U27314 (N_27314,N_27219,N_27175);
xor U27315 (N_27315,N_27187,N_27045);
nand U27316 (N_27316,N_27181,N_27073);
nand U27317 (N_27317,N_27028,N_27016);
nor U27318 (N_27318,N_27027,N_27212);
xor U27319 (N_27319,N_27098,N_27186);
and U27320 (N_27320,N_27217,N_27092);
and U27321 (N_27321,N_27022,N_27178);
xnor U27322 (N_27322,N_27014,N_27236);
nand U27323 (N_27323,N_27123,N_27172);
nor U27324 (N_27324,N_27210,N_27165);
nand U27325 (N_27325,N_27089,N_27242);
nand U27326 (N_27326,N_27059,N_27122);
xnor U27327 (N_27327,N_27079,N_27232);
xor U27328 (N_27328,N_27097,N_27104);
or U27329 (N_27329,N_27106,N_27081);
or U27330 (N_27330,N_27158,N_27146);
or U27331 (N_27331,N_27099,N_27032);
and U27332 (N_27332,N_27235,N_27044);
nand U27333 (N_27333,N_27183,N_27063);
nand U27334 (N_27334,N_27040,N_27163);
xnor U27335 (N_27335,N_27179,N_27126);
nand U27336 (N_27336,N_27177,N_27007);
or U27337 (N_27337,N_27228,N_27019);
or U27338 (N_27338,N_27070,N_27211);
xnor U27339 (N_27339,N_27154,N_27230);
or U27340 (N_27340,N_27096,N_27013);
xnor U27341 (N_27341,N_27090,N_27088);
nand U27342 (N_27342,N_27050,N_27197);
and U27343 (N_27343,N_27245,N_27005);
nor U27344 (N_27344,N_27012,N_27209);
xnor U27345 (N_27345,N_27170,N_27145);
nand U27346 (N_27346,N_27131,N_27087);
nand U27347 (N_27347,N_27223,N_27226);
xor U27348 (N_27348,N_27143,N_27043);
or U27349 (N_27349,N_27025,N_27133);
nand U27350 (N_27350,N_27168,N_27075);
xor U27351 (N_27351,N_27039,N_27140);
xnor U27352 (N_27352,N_27161,N_27048);
and U27353 (N_27353,N_27034,N_27147);
and U27354 (N_27354,N_27067,N_27066);
xor U27355 (N_27355,N_27156,N_27243);
nand U27356 (N_27356,N_27198,N_27077);
xor U27357 (N_27357,N_27233,N_27037);
nand U27358 (N_27358,N_27231,N_27216);
or U27359 (N_27359,N_27010,N_27018);
nand U27360 (N_27360,N_27142,N_27248);
xor U27361 (N_27361,N_27193,N_27115);
nor U27362 (N_27362,N_27023,N_27173);
nand U27363 (N_27363,N_27155,N_27110);
and U27364 (N_27364,N_27202,N_27139);
nand U27365 (N_27365,N_27201,N_27074);
nor U27366 (N_27366,N_27055,N_27053);
and U27367 (N_27367,N_27234,N_27174);
xor U27368 (N_27368,N_27222,N_27042);
nor U27369 (N_27369,N_27128,N_27150);
nand U27370 (N_27370,N_27185,N_27246);
or U27371 (N_27371,N_27148,N_27062);
nand U27372 (N_27372,N_27229,N_27003);
and U27373 (N_27373,N_27157,N_27152);
nor U27374 (N_27374,N_27149,N_27072);
and U27375 (N_27375,N_27045,N_27004);
xor U27376 (N_27376,N_27228,N_27081);
nor U27377 (N_27377,N_27019,N_27242);
nor U27378 (N_27378,N_27234,N_27123);
and U27379 (N_27379,N_27066,N_27144);
xor U27380 (N_27380,N_27185,N_27033);
nand U27381 (N_27381,N_27216,N_27236);
nor U27382 (N_27382,N_27116,N_27200);
and U27383 (N_27383,N_27166,N_27186);
and U27384 (N_27384,N_27016,N_27162);
nand U27385 (N_27385,N_27110,N_27146);
and U27386 (N_27386,N_27249,N_27128);
nand U27387 (N_27387,N_27205,N_27018);
and U27388 (N_27388,N_27208,N_27192);
xor U27389 (N_27389,N_27003,N_27151);
and U27390 (N_27390,N_27181,N_27052);
xor U27391 (N_27391,N_27043,N_27175);
nand U27392 (N_27392,N_27066,N_27232);
or U27393 (N_27393,N_27224,N_27183);
nor U27394 (N_27394,N_27093,N_27100);
xnor U27395 (N_27395,N_27221,N_27177);
nor U27396 (N_27396,N_27233,N_27221);
nand U27397 (N_27397,N_27086,N_27232);
or U27398 (N_27398,N_27056,N_27246);
or U27399 (N_27399,N_27039,N_27167);
nor U27400 (N_27400,N_27045,N_27048);
or U27401 (N_27401,N_27137,N_27204);
and U27402 (N_27402,N_27127,N_27155);
or U27403 (N_27403,N_27192,N_27160);
nand U27404 (N_27404,N_27082,N_27211);
and U27405 (N_27405,N_27053,N_27132);
nor U27406 (N_27406,N_27153,N_27185);
xor U27407 (N_27407,N_27089,N_27002);
or U27408 (N_27408,N_27059,N_27070);
and U27409 (N_27409,N_27224,N_27054);
or U27410 (N_27410,N_27230,N_27085);
xnor U27411 (N_27411,N_27037,N_27144);
nor U27412 (N_27412,N_27146,N_27099);
nor U27413 (N_27413,N_27131,N_27026);
and U27414 (N_27414,N_27249,N_27218);
nand U27415 (N_27415,N_27231,N_27056);
or U27416 (N_27416,N_27005,N_27042);
and U27417 (N_27417,N_27184,N_27108);
and U27418 (N_27418,N_27114,N_27005);
nor U27419 (N_27419,N_27037,N_27126);
and U27420 (N_27420,N_27149,N_27169);
and U27421 (N_27421,N_27103,N_27129);
or U27422 (N_27422,N_27003,N_27005);
nand U27423 (N_27423,N_27019,N_27219);
and U27424 (N_27424,N_27028,N_27139);
xnor U27425 (N_27425,N_27053,N_27200);
and U27426 (N_27426,N_27192,N_27105);
nand U27427 (N_27427,N_27173,N_27090);
or U27428 (N_27428,N_27095,N_27152);
xor U27429 (N_27429,N_27089,N_27139);
nor U27430 (N_27430,N_27077,N_27025);
nand U27431 (N_27431,N_27236,N_27135);
xor U27432 (N_27432,N_27217,N_27218);
nor U27433 (N_27433,N_27220,N_27132);
and U27434 (N_27434,N_27217,N_27026);
xor U27435 (N_27435,N_27113,N_27197);
and U27436 (N_27436,N_27153,N_27165);
nand U27437 (N_27437,N_27076,N_27037);
nor U27438 (N_27438,N_27243,N_27083);
nand U27439 (N_27439,N_27043,N_27227);
and U27440 (N_27440,N_27230,N_27239);
nor U27441 (N_27441,N_27162,N_27238);
nand U27442 (N_27442,N_27065,N_27049);
xor U27443 (N_27443,N_27182,N_27062);
nor U27444 (N_27444,N_27195,N_27180);
or U27445 (N_27445,N_27226,N_27164);
nand U27446 (N_27446,N_27008,N_27018);
or U27447 (N_27447,N_27102,N_27078);
and U27448 (N_27448,N_27013,N_27097);
nor U27449 (N_27449,N_27223,N_27073);
or U27450 (N_27450,N_27224,N_27127);
nor U27451 (N_27451,N_27088,N_27102);
xnor U27452 (N_27452,N_27156,N_27085);
nand U27453 (N_27453,N_27125,N_27137);
and U27454 (N_27454,N_27078,N_27214);
and U27455 (N_27455,N_27128,N_27171);
or U27456 (N_27456,N_27111,N_27049);
xor U27457 (N_27457,N_27223,N_27248);
nor U27458 (N_27458,N_27115,N_27150);
and U27459 (N_27459,N_27215,N_27164);
xnor U27460 (N_27460,N_27171,N_27010);
xnor U27461 (N_27461,N_27109,N_27011);
nor U27462 (N_27462,N_27243,N_27195);
nand U27463 (N_27463,N_27159,N_27122);
nor U27464 (N_27464,N_27245,N_27118);
nand U27465 (N_27465,N_27131,N_27085);
nand U27466 (N_27466,N_27086,N_27111);
or U27467 (N_27467,N_27237,N_27144);
or U27468 (N_27468,N_27081,N_27249);
nor U27469 (N_27469,N_27187,N_27095);
nand U27470 (N_27470,N_27168,N_27166);
xor U27471 (N_27471,N_27198,N_27093);
nor U27472 (N_27472,N_27210,N_27053);
nor U27473 (N_27473,N_27239,N_27063);
nor U27474 (N_27474,N_27166,N_27005);
or U27475 (N_27475,N_27174,N_27109);
nand U27476 (N_27476,N_27166,N_27030);
and U27477 (N_27477,N_27168,N_27055);
xor U27478 (N_27478,N_27126,N_27198);
nand U27479 (N_27479,N_27170,N_27191);
xnor U27480 (N_27480,N_27080,N_27074);
nor U27481 (N_27481,N_27116,N_27086);
or U27482 (N_27482,N_27132,N_27008);
and U27483 (N_27483,N_27138,N_27014);
xnor U27484 (N_27484,N_27181,N_27064);
nor U27485 (N_27485,N_27160,N_27180);
nand U27486 (N_27486,N_27175,N_27039);
nor U27487 (N_27487,N_27229,N_27196);
nand U27488 (N_27488,N_27216,N_27058);
xnor U27489 (N_27489,N_27035,N_27028);
or U27490 (N_27490,N_27035,N_27072);
xor U27491 (N_27491,N_27202,N_27154);
xor U27492 (N_27492,N_27121,N_27030);
or U27493 (N_27493,N_27238,N_27087);
and U27494 (N_27494,N_27009,N_27199);
nand U27495 (N_27495,N_27061,N_27131);
nand U27496 (N_27496,N_27052,N_27203);
xnor U27497 (N_27497,N_27115,N_27187);
or U27498 (N_27498,N_27066,N_27150);
xor U27499 (N_27499,N_27195,N_27025);
xnor U27500 (N_27500,N_27263,N_27323);
or U27501 (N_27501,N_27450,N_27304);
nor U27502 (N_27502,N_27496,N_27362);
or U27503 (N_27503,N_27381,N_27281);
or U27504 (N_27504,N_27451,N_27486);
xnor U27505 (N_27505,N_27345,N_27459);
or U27506 (N_27506,N_27260,N_27359);
or U27507 (N_27507,N_27422,N_27366);
and U27508 (N_27508,N_27485,N_27467);
and U27509 (N_27509,N_27404,N_27465);
xor U27510 (N_27510,N_27406,N_27448);
and U27511 (N_27511,N_27273,N_27355);
or U27512 (N_27512,N_27363,N_27456);
nor U27513 (N_27513,N_27285,N_27369);
or U27514 (N_27514,N_27311,N_27343);
and U27515 (N_27515,N_27305,N_27474);
nor U27516 (N_27516,N_27418,N_27307);
and U27517 (N_27517,N_27278,N_27440);
or U27518 (N_27518,N_27457,N_27443);
and U27519 (N_27519,N_27360,N_27405);
xor U27520 (N_27520,N_27371,N_27267);
nor U27521 (N_27521,N_27268,N_27379);
nor U27522 (N_27522,N_27387,N_27331);
nor U27523 (N_27523,N_27365,N_27472);
and U27524 (N_27524,N_27478,N_27468);
and U27525 (N_27525,N_27453,N_27292);
or U27526 (N_27526,N_27430,N_27463);
or U27527 (N_27527,N_27253,N_27390);
and U27528 (N_27528,N_27491,N_27403);
nor U27529 (N_27529,N_27279,N_27287);
or U27530 (N_27530,N_27352,N_27255);
nand U27531 (N_27531,N_27481,N_27367);
nand U27532 (N_27532,N_27476,N_27291);
xnor U27533 (N_27533,N_27330,N_27421);
or U27534 (N_27534,N_27386,N_27332);
xnor U27535 (N_27535,N_27286,N_27393);
xnor U27536 (N_27536,N_27283,N_27340);
and U27537 (N_27537,N_27257,N_27460);
xnor U27538 (N_27538,N_27334,N_27270);
or U27539 (N_27539,N_27316,N_27497);
nor U27540 (N_27540,N_27389,N_27266);
and U27541 (N_27541,N_27301,N_27464);
or U27542 (N_27542,N_27347,N_27319);
or U27543 (N_27543,N_27261,N_27274);
and U27544 (N_27544,N_27484,N_27428);
and U27545 (N_27545,N_27425,N_27452);
nor U27546 (N_27546,N_27350,N_27402);
nand U27547 (N_27547,N_27300,N_27349);
or U27548 (N_27548,N_27419,N_27473);
nor U27549 (N_27549,N_27313,N_27407);
nand U27550 (N_27550,N_27437,N_27272);
xor U27551 (N_27551,N_27470,N_27434);
and U27552 (N_27552,N_27490,N_27326);
and U27553 (N_27553,N_27251,N_27455);
and U27554 (N_27554,N_27364,N_27454);
nand U27555 (N_27555,N_27436,N_27494);
xnor U27556 (N_27556,N_27401,N_27294);
nor U27557 (N_27557,N_27320,N_27357);
or U27558 (N_27558,N_27482,N_27314);
nor U27559 (N_27559,N_27312,N_27383);
nor U27560 (N_27560,N_27375,N_27321);
nand U27561 (N_27561,N_27318,N_27271);
nand U27562 (N_27562,N_27397,N_27299);
or U27563 (N_27563,N_27374,N_27414);
and U27564 (N_27564,N_27471,N_27342);
or U27565 (N_27565,N_27259,N_27475);
nand U27566 (N_27566,N_27391,N_27308);
nor U27567 (N_27567,N_27410,N_27256);
nor U27568 (N_27568,N_27358,N_27493);
nand U27569 (N_27569,N_27339,N_27395);
and U27570 (N_27570,N_27447,N_27409);
or U27571 (N_27571,N_27444,N_27322);
xnor U27572 (N_27572,N_27317,N_27495);
xor U27573 (N_27573,N_27341,N_27297);
nor U27574 (N_27574,N_27327,N_27400);
or U27575 (N_27575,N_27439,N_27426);
and U27576 (N_27576,N_27427,N_27431);
nand U27577 (N_27577,N_27250,N_27396);
nor U27578 (N_27578,N_27296,N_27373);
or U27579 (N_27579,N_27435,N_27380);
nand U27580 (N_27580,N_27315,N_27282);
nor U27581 (N_27581,N_27290,N_27462);
nand U27582 (N_27582,N_27392,N_27337);
nand U27583 (N_27583,N_27492,N_27498);
nand U27584 (N_27584,N_27277,N_27398);
or U27585 (N_27585,N_27412,N_27328);
or U27586 (N_27586,N_27310,N_27420);
nand U27587 (N_27587,N_27372,N_27370);
xnor U27588 (N_27588,N_27446,N_27442);
nand U27589 (N_27589,N_27254,N_27399);
nor U27590 (N_27590,N_27388,N_27354);
nor U27591 (N_27591,N_27346,N_27264);
or U27592 (N_27592,N_27353,N_27329);
or U27593 (N_27593,N_27262,N_27458);
or U27594 (N_27594,N_27411,N_27351);
xor U27595 (N_27595,N_27432,N_27269);
nand U27596 (N_27596,N_27356,N_27284);
nor U27597 (N_27597,N_27480,N_27258);
and U27598 (N_27598,N_27309,N_27348);
xnor U27599 (N_27599,N_27477,N_27376);
xnor U27600 (N_27600,N_27479,N_27413);
nor U27601 (N_27601,N_27441,N_27378);
nor U27602 (N_27602,N_27295,N_27489);
and U27603 (N_27603,N_27449,N_27461);
and U27604 (N_27604,N_27333,N_27384);
and U27605 (N_27605,N_27433,N_27288);
nand U27606 (N_27606,N_27293,N_27280);
nor U27607 (N_27607,N_27416,N_27275);
nand U27608 (N_27608,N_27424,N_27289);
nand U27609 (N_27609,N_27302,N_27487);
xnor U27610 (N_27610,N_27298,N_27483);
xnor U27611 (N_27611,N_27276,N_27265);
or U27612 (N_27612,N_27394,N_27303);
or U27613 (N_27613,N_27368,N_27445);
and U27614 (N_27614,N_27499,N_27335);
xnor U27615 (N_27615,N_27344,N_27423);
or U27616 (N_27616,N_27338,N_27252);
xnor U27617 (N_27617,N_27385,N_27336);
nand U27618 (N_27618,N_27306,N_27429);
or U27619 (N_27619,N_27377,N_27382);
and U27620 (N_27620,N_27438,N_27361);
or U27621 (N_27621,N_27324,N_27408);
or U27622 (N_27622,N_27466,N_27417);
nor U27623 (N_27623,N_27469,N_27488);
and U27624 (N_27624,N_27325,N_27415);
or U27625 (N_27625,N_27414,N_27291);
and U27626 (N_27626,N_27482,N_27293);
and U27627 (N_27627,N_27314,N_27402);
and U27628 (N_27628,N_27353,N_27370);
or U27629 (N_27629,N_27463,N_27438);
or U27630 (N_27630,N_27385,N_27267);
nor U27631 (N_27631,N_27366,N_27265);
xnor U27632 (N_27632,N_27354,N_27417);
or U27633 (N_27633,N_27280,N_27444);
nor U27634 (N_27634,N_27412,N_27429);
nand U27635 (N_27635,N_27299,N_27289);
or U27636 (N_27636,N_27343,N_27432);
nand U27637 (N_27637,N_27375,N_27497);
or U27638 (N_27638,N_27468,N_27394);
nand U27639 (N_27639,N_27488,N_27329);
nand U27640 (N_27640,N_27383,N_27286);
nor U27641 (N_27641,N_27322,N_27337);
or U27642 (N_27642,N_27432,N_27375);
nand U27643 (N_27643,N_27492,N_27340);
nor U27644 (N_27644,N_27399,N_27260);
xnor U27645 (N_27645,N_27487,N_27356);
or U27646 (N_27646,N_27373,N_27325);
nand U27647 (N_27647,N_27342,N_27302);
xor U27648 (N_27648,N_27370,N_27426);
xnor U27649 (N_27649,N_27469,N_27433);
nand U27650 (N_27650,N_27347,N_27294);
or U27651 (N_27651,N_27463,N_27344);
xor U27652 (N_27652,N_27304,N_27279);
nand U27653 (N_27653,N_27253,N_27313);
and U27654 (N_27654,N_27394,N_27487);
nand U27655 (N_27655,N_27341,N_27426);
xnor U27656 (N_27656,N_27437,N_27420);
and U27657 (N_27657,N_27267,N_27467);
nand U27658 (N_27658,N_27409,N_27499);
and U27659 (N_27659,N_27342,N_27345);
and U27660 (N_27660,N_27410,N_27291);
xor U27661 (N_27661,N_27427,N_27493);
nor U27662 (N_27662,N_27289,N_27316);
xnor U27663 (N_27663,N_27295,N_27477);
xor U27664 (N_27664,N_27398,N_27366);
nor U27665 (N_27665,N_27438,N_27296);
nand U27666 (N_27666,N_27268,N_27460);
or U27667 (N_27667,N_27404,N_27348);
nand U27668 (N_27668,N_27388,N_27261);
nand U27669 (N_27669,N_27392,N_27484);
nor U27670 (N_27670,N_27440,N_27488);
xor U27671 (N_27671,N_27259,N_27497);
nand U27672 (N_27672,N_27409,N_27406);
nand U27673 (N_27673,N_27290,N_27366);
xnor U27674 (N_27674,N_27293,N_27324);
xor U27675 (N_27675,N_27394,N_27414);
nor U27676 (N_27676,N_27358,N_27352);
or U27677 (N_27677,N_27493,N_27335);
nand U27678 (N_27678,N_27377,N_27423);
and U27679 (N_27679,N_27256,N_27472);
xor U27680 (N_27680,N_27309,N_27444);
and U27681 (N_27681,N_27262,N_27325);
xor U27682 (N_27682,N_27345,N_27291);
or U27683 (N_27683,N_27467,N_27498);
xnor U27684 (N_27684,N_27350,N_27286);
nor U27685 (N_27685,N_27490,N_27292);
nand U27686 (N_27686,N_27279,N_27466);
or U27687 (N_27687,N_27349,N_27493);
or U27688 (N_27688,N_27433,N_27293);
and U27689 (N_27689,N_27350,N_27309);
nor U27690 (N_27690,N_27253,N_27472);
nor U27691 (N_27691,N_27288,N_27392);
nand U27692 (N_27692,N_27250,N_27471);
and U27693 (N_27693,N_27386,N_27306);
nor U27694 (N_27694,N_27326,N_27315);
and U27695 (N_27695,N_27356,N_27426);
xor U27696 (N_27696,N_27281,N_27428);
or U27697 (N_27697,N_27396,N_27399);
nor U27698 (N_27698,N_27376,N_27293);
and U27699 (N_27699,N_27310,N_27479);
nor U27700 (N_27700,N_27316,N_27322);
nand U27701 (N_27701,N_27323,N_27352);
nand U27702 (N_27702,N_27311,N_27318);
nand U27703 (N_27703,N_27273,N_27466);
and U27704 (N_27704,N_27410,N_27422);
nor U27705 (N_27705,N_27354,N_27483);
or U27706 (N_27706,N_27347,N_27373);
and U27707 (N_27707,N_27426,N_27490);
nor U27708 (N_27708,N_27399,N_27492);
xor U27709 (N_27709,N_27434,N_27318);
or U27710 (N_27710,N_27488,N_27431);
and U27711 (N_27711,N_27448,N_27266);
or U27712 (N_27712,N_27484,N_27322);
nor U27713 (N_27713,N_27304,N_27493);
xnor U27714 (N_27714,N_27263,N_27295);
nor U27715 (N_27715,N_27474,N_27365);
or U27716 (N_27716,N_27393,N_27311);
and U27717 (N_27717,N_27367,N_27499);
and U27718 (N_27718,N_27343,N_27428);
xnor U27719 (N_27719,N_27424,N_27454);
xnor U27720 (N_27720,N_27336,N_27317);
nor U27721 (N_27721,N_27358,N_27463);
nand U27722 (N_27722,N_27416,N_27278);
and U27723 (N_27723,N_27319,N_27475);
nand U27724 (N_27724,N_27319,N_27258);
or U27725 (N_27725,N_27481,N_27467);
or U27726 (N_27726,N_27361,N_27293);
nor U27727 (N_27727,N_27280,N_27480);
nor U27728 (N_27728,N_27339,N_27497);
and U27729 (N_27729,N_27257,N_27453);
xor U27730 (N_27730,N_27403,N_27265);
nand U27731 (N_27731,N_27276,N_27391);
nand U27732 (N_27732,N_27485,N_27464);
nand U27733 (N_27733,N_27288,N_27306);
nand U27734 (N_27734,N_27352,N_27367);
nand U27735 (N_27735,N_27340,N_27339);
and U27736 (N_27736,N_27308,N_27495);
and U27737 (N_27737,N_27323,N_27455);
nand U27738 (N_27738,N_27342,N_27487);
nand U27739 (N_27739,N_27330,N_27286);
and U27740 (N_27740,N_27363,N_27266);
or U27741 (N_27741,N_27407,N_27263);
nand U27742 (N_27742,N_27317,N_27396);
and U27743 (N_27743,N_27270,N_27282);
nand U27744 (N_27744,N_27399,N_27270);
nand U27745 (N_27745,N_27316,N_27344);
and U27746 (N_27746,N_27362,N_27296);
xor U27747 (N_27747,N_27283,N_27454);
and U27748 (N_27748,N_27259,N_27341);
and U27749 (N_27749,N_27379,N_27264);
nor U27750 (N_27750,N_27740,N_27619);
and U27751 (N_27751,N_27700,N_27509);
or U27752 (N_27752,N_27669,N_27527);
nor U27753 (N_27753,N_27691,N_27713);
or U27754 (N_27754,N_27729,N_27589);
and U27755 (N_27755,N_27648,N_27654);
nand U27756 (N_27756,N_27635,N_27668);
nand U27757 (N_27757,N_27709,N_27597);
or U27758 (N_27758,N_27550,N_27566);
or U27759 (N_27759,N_27657,N_27575);
and U27760 (N_27760,N_27693,N_27698);
xnor U27761 (N_27761,N_27683,N_27677);
or U27762 (N_27762,N_27518,N_27651);
or U27763 (N_27763,N_27570,N_27632);
nor U27764 (N_27764,N_27702,N_27731);
and U27765 (N_27765,N_27689,N_27584);
and U27766 (N_27766,N_27736,N_27524);
nor U27767 (N_27767,N_27580,N_27665);
or U27768 (N_27768,N_27551,N_27673);
nand U27769 (N_27769,N_27701,N_27722);
nor U27770 (N_27770,N_27607,N_27561);
nor U27771 (N_27771,N_27644,N_27525);
nor U27772 (N_27772,N_27517,N_27549);
xnor U27773 (N_27773,N_27563,N_27643);
and U27774 (N_27774,N_27650,N_27539);
nand U27775 (N_27775,N_27558,N_27707);
nor U27776 (N_27776,N_27610,N_27557);
nand U27777 (N_27777,N_27600,N_27547);
xnor U27778 (N_27778,N_27695,N_27641);
xnor U27779 (N_27779,N_27679,N_27714);
and U27780 (N_27780,N_27726,N_27605);
xnor U27781 (N_27781,N_27741,N_27744);
nor U27782 (N_27782,N_27749,N_27661);
and U27783 (N_27783,N_27581,N_27667);
or U27784 (N_27784,N_27652,N_27615);
or U27785 (N_27785,N_27687,N_27569);
xor U27786 (N_27786,N_27670,N_27634);
nand U27787 (N_27787,N_27653,N_27717);
nor U27788 (N_27788,N_27672,N_27576);
nand U27789 (N_27789,N_27628,N_27636);
nor U27790 (N_27790,N_27624,N_27617);
xor U27791 (N_27791,N_27505,N_27737);
nor U27792 (N_27792,N_27572,N_27681);
xnor U27793 (N_27793,N_27533,N_27703);
xnor U27794 (N_27794,N_27523,N_27692);
xnor U27795 (N_27795,N_27627,N_27606);
nor U27796 (N_27796,N_27500,N_27649);
xnor U27797 (N_27797,N_27564,N_27603);
or U27798 (N_27798,N_27540,N_27526);
or U27799 (N_27799,N_27633,N_27507);
nor U27800 (N_27800,N_27658,N_27529);
and U27801 (N_27801,N_27697,N_27577);
nand U27802 (N_27802,N_27743,N_27711);
nor U27803 (N_27803,N_27536,N_27554);
nor U27804 (N_27804,N_27516,N_27594);
and U27805 (N_27805,N_27625,N_27515);
nand U27806 (N_27806,N_27716,N_27694);
nand U27807 (N_27807,N_27637,N_27696);
xnor U27808 (N_27808,N_27715,N_27640);
and U27809 (N_27809,N_27638,N_27586);
xor U27810 (N_27810,N_27590,N_27646);
or U27811 (N_27811,N_27676,N_27656);
and U27812 (N_27812,N_27647,N_27645);
nor U27813 (N_27813,N_27562,N_27735);
and U27814 (N_27814,N_27612,N_27506);
nor U27815 (N_27815,N_27655,N_27521);
or U27816 (N_27816,N_27623,N_27574);
nor U27817 (N_27817,N_27732,N_27601);
xnor U27818 (N_27818,N_27614,N_27739);
xnor U27819 (N_27819,N_27721,N_27690);
and U27820 (N_27820,N_27537,N_27556);
nand U27821 (N_27821,N_27510,N_27542);
or U27822 (N_27822,N_27583,N_27560);
nand U27823 (N_27823,N_27728,N_27546);
nor U27824 (N_27824,N_27503,N_27553);
nand U27825 (N_27825,N_27543,N_27592);
and U27826 (N_27826,N_27666,N_27530);
nor U27827 (N_27827,N_27680,N_27704);
xnor U27828 (N_27828,N_27686,N_27559);
nor U27829 (N_27829,N_27512,N_27659);
nor U27830 (N_27830,N_27678,N_27520);
nor U27831 (N_27831,N_27538,N_27664);
and U27832 (N_27832,N_27591,N_27568);
and U27833 (N_27833,N_27682,N_27579);
and U27834 (N_27834,N_27688,N_27708);
nand U27835 (N_27835,N_27508,N_27571);
and U27836 (N_27836,N_27596,N_27587);
xor U27837 (N_27837,N_27671,N_27642);
and U27838 (N_27838,N_27725,N_27541);
nor U27839 (N_27839,N_27502,N_27733);
xnor U27840 (N_27840,N_27660,N_27675);
xor U27841 (N_27841,N_27519,N_27511);
xnor U27842 (N_27842,N_27548,N_27723);
and U27843 (N_27843,N_27609,N_27684);
or U27844 (N_27844,N_27620,N_27626);
or U27845 (N_27845,N_27712,N_27674);
nand U27846 (N_27846,N_27618,N_27528);
xor U27847 (N_27847,N_27738,N_27629);
and U27848 (N_27848,N_27724,N_27706);
and U27849 (N_27849,N_27685,N_27598);
nor U27850 (N_27850,N_27555,N_27532);
nand U27851 (N_27851,N_27534,N_27746);
nand U27852 (N_27852,N_27501,N_27595);
nor U27853 (N_27853,N_27565,N_27720);
xor U27854 (N_27854,N_27593,N_27699);
xnor U27855 (N_27855,N_27705,N_27582);
nand U27856 (N_27856,N_27514,N_27727);
and U27857 (N_27857,N_27588,N_27639);
nor U27858 (N_27858,N_27745,N_27730);
xor U27859 (N_27859,N_27545,N_27622);
or U27860 (N_27860,N_27585,N_27567);
nand U27861 (N_27861,N_27631,N_27742);
xnor U27862 (N_27862,N_27578,N_27710);
or U27863 (N_27863,N_27608,N_27719);
or U27864 (N_27864,N_27616,N_27604);
nor U27865 (N_27865,N_27613,N_27531);
or U27866 (N_27866,N_27602,N_27544);
and U27867 (N_27867,N_27513,N_27663);
and U27868 (N_27868,N_27662,N_27734);
nand U27869 (N_27869,N_27522,N_27630);
xnor U27870 (N_27870,N_27621,N_27573);
or U27871 (N_27871,N_27748,N_27535);
or U27872 (N_27872,N_27552,N_27504);
xor U27873 (N_27873,N_27599,N_27611);
or U27874 (N_27874,N_27747,N_27718);
xnor U27875 (N_27875,N_27548,N_27705);
nand U27876 (N_27876,N_27730,N_27568);
xnor U27877 (N_27877,N_27591,N_27669);
nand U27878 (N_27878,N_27526,N_27567);
and U27879 (N_27879,N_27747,N_27560);
nand U27880 (N_27880,N_27721,N_27646);
or U27881 (N_27881,N_27734,N_27565);
xor U27882 (N_27882,N_27700,N_27745);
xor U27883 (N_27883,N_27741,N_27628);
and U27884 (N_27884,N_27748,N_27740);
or U27885 (N_27885,N_27692,N_27568);
or U27886 (N_27886,N_27612,N_27626);
nor U27887 (N_27887,N_27729,N_27747);
nor U27888 (N_27888,N_27525,N_27747);
and U27889 (N_27889,N_27718,N_27713);
nor U27890 (N_27890,N_27615,N_27508);
xnor U27891 (N_27891,N_27506,N_27584);
xor U27892 (N_27892,N_27735,N_27582);
nand U27893 (N_27893,N_27732,N_27683);
nor U27894 (N_27894,N_27513,N_27685);
nor U27895 (N_27895,N_27707,N_27697);
or U27896 (N_27896,N_27693,N_27586);
nand U27897 (N_27897,N_27610,N_27630);
xnor U27898 (N_27898,N_27704,N_27621);
xor U27899 (N_27899,N_27633,N_27700);
xnor U27900 (N_27900,N_27527,N_27511);
nor U27901 (N_27901,N_27523,N_27544);
xor U27902 (N_27902,N_27725,N_27592);
or U27903 (N_27903,N_27601,N_27730);
nand U27904 (N_27904,N_27589,N_27745);
and U27905 (N_27905,N_27657,N_27708);
xor U27906 (N_27906,N_27502,N_27659);
or U27907 (N_27907,N_27689,N_27616);
nand U27908 (N_27908,N_27619,N_27522);
or U27909 (N_27909,N_27608,N_27696);
or U27910 (N_27910,N_27725,N_27523);
or U27911 (N_27911,N_27610,N_27503);
xnor U27912 (N_27912,N_27626,N_27704);
xor U27913 (N_27913,N_27712,N_27510);
nor U27914 (N_27914,N_27618,N_27553);
xor U27915 (N_27915,N_27566,N_27684);
nor U27916 (N_27916,N_27668,N_27541);
and U27917 (N_27917,N_27524,N_27680);
or U27918 (N_27918,N_27693,N_27577);
xor U27919 (N_27919,N_27735,N_27517);
and U27920 (N_27920,N_27725,N_27517);
xnor U27921 (N_27921,N_27554,N_27691);
xnor U27922 (N_27922,N_27528,N_27649);
or U27923 (N_27923,N_27627,N_27573);
xor U27924 (N_27924,N_27744,N_27611);
xnor U27925 (N_27925,N_27512,N_27648);
nand U27926 (N_27926,N_27506,N_27690);
and U27927 (N_27927,N_27610,N_27663);
or U27928 (N_27928,N_27727,N_27661);
xnor U27929 (N_27929,N_27635,N_27544);
xnor U27930 (N_27930,N_27575,N_27687);
or U27931 (N_27931,N_27560,N_27618);
nand U27932 (N_27932,N_27672,N_27564);
xnor U27933 (N_27933,N_27594,N_27511);
nor U27934 (N_27934,N_27733,N_27605);
nand U27935 (N_27935,N_27694,N_27543);
xnor U27936 (N_27936,N_27693,N_27583);
nand U27937 (N_27937,N_27726,N_27603);
nand U27938 (N_27938,N_27532,N_27727);
and U27939 (N_27939,N_27627,N_27694);
or U27940 (N_27940,N_27533,N_27661);
nand U27941 (N_27941,N_27680,N_27611);
xor U27942 (N_27942,N_27700,N_27649);
nand U27943 (N_27943,N_27612,N_27668);
xnor U27944 (N_27944,N_27566,N_27544);
xor U27945 (N_27945,N_27686,N_27713);
xnor U27946 (N_27946,N_27650,N_27524);
xor U27947 (N_27947,N_27688,N_27529);
and U27948 (N_27948,N_27602,N_27684);
nor U27949 (N_27949,N_27580,N_27518);
and U27950 (N_27950,N_27665,N_27720);
nor U27951 (N_27951,N_27727,N_27662);
or U27952 (N_27952,N_27710,N_27734);
and U27953 (N_27953,N_27649,N_27713);
nor U27954 (N_27954,N_27613,N_27541);
and U27955 (N_27955,N_27723,N_27705);
xor U27956 (N_27956,N_27521,N_27732);
and U27957 (N_27957,N_27590,N_27625);
nand U27958 (N_27958,N_27531,N_27577);
and U27959 (N_27959,N_27660,N_27670);
or U27960 (N_27960,N_27616,N_27534);
xnor U27961 (N_27961,N_27693,N_27595);
xor U27962 (N_27962,N_27627,N_27593);
and U27963 (N_27963,N_27511,N_27545);
nand U27964 (N_27964,N_27714,N_27547);
nand U27965 (N_27965,N_27500,N_27566);
or U27966 (N_27966,N_27586,N_27685);
nor U27967 (N_27967,N_27717,N_27695);
xnor U27968 (N_27968,N_27682,N_27595);
nor U27969 (N_27969,N_27725,N_27526);
xnor U27970 (N_27970,N_27691,N_27536);
nor U27971 (N_27971,N_27635,N_27659);
xor U27972 (N_27972,N_27591,N_27645);
xnor U27973 (N_27973,N_27623,N_27555);
and U27974 (N_27974,N_27543,N_27611);
or U27975 (N_27975,N_27521,N_27525);
or U27976 (N_27976,N_27627,N_27605);
and U27977 (N_27977,N_27725,N_27602);
and U27978 (N_27978,N_27551,N_27730);
and U27979 (N_27979,N_27655,N_27686);
nor U27980 (N_27980,N_27703,N_27646);
nand U27981 (N_27981,N_27655,N_27506);
nor U27982 (N_27982,N_27626,N_27615);
xnor U27983 (N_27983,N_27591,N_27663);
nor U27984 (N_27984,N_27620,N_27710);
and U27985 (N_27985,N_27595,N_27592);
nand U27986 (N_27986,N_27662,N_27621);
and U27987 (N_27987,N_27565,N_27563);
xnor U27988 (N_27988,N_27570,N_27568);
and U27989 (N_27989,N_27630,N_27543);
or U27990 (N_27990,N_27621,N_27726);
nor U27991 (N_27991,N_27642,N_27719);
and U27992 (N_27992,N_27561,N_27553);
and U27993 (N_27993,N_27506,N_27665);
nor U27994 (N_27994,N_27664,N_27607);
and U27995 (N_27995,N_27670,N_27745);
nor U27996 (N_27996,N_27645,N_27518);
nand U27997 (N_27997,N_27652,N_27693);
and U27998 (N_27998,N_27656,N_27690);
nand U27999 (N_27999,N_27557,N_27697);
nand U28000 (N_28000,N_27797,N_27980);
nor U28001 (N_28001,N_27801,N_27815);
xor U28002 (N_28002,N_27832,N_27972);
nand U28003 (N_28003,N_27768,N_27885);
or U28004 (N_28004,N_27756,N_27944);
nor U28005 (N_28005,N_27953,N_27952);
xnor U28006 (N_28006,N_27989,N_27910);
and U28007 (N_28007,N_27785,N_27852);
xnor U28008 (N_28008,N_27977,N_27878);
and U28009 (N_28009,N_27882,N_27967);
xnor U28010 (N_28010,N_27820,N_27920);
and U28011 (N_28011,N_27915,N_27779);
nor U28012 (N_28012,N_27931,N_27862);
and U28013 (N_28013,N_27788,N_27771);
nand U28014 (N_28014,N_27908,N_27764);
and U28015 (N_28015,N_27906,N_27757);
nand U28016 (N_28016,N_27772,N_27750);
or U28017 (N_28017,N_27775,N_27760);
and U28018 (N_28018,N_27751,N_27899);
nor U28019 (N_28019,N_27867,N_27848);
xor U28020 (N_28020,N_27816,N_27805);
or U28021 (N_28021,N_27941,N_27802);
xnor U28022 (N_28022,N_27793,N_27965);
nor U28023 (N_28023,N_27819,N_27752);
nand U28024 (N_28024,N_27928,N_27790);
and U28025 (N_28025,N_27803,N_27861);
nand U28026 (N_28026,N_27940,N_27942);
nand U28027 (N_28027,N_27971,N_27887);
nand U28028 (N_28028,N_27782,N_27813);
or U28029 (N_28029,N_27930,N_27886);
or U28030 (N_28030,N_27880,N_27812);
and U28031 (N_28031,N_27976,N_27870);
nor U28032 (N_28032,N_27824,N_27973);
or U28033 (N_28033,N_27925,N_27759);
nand U28034 (N_28034,N_27798,N_27868);
and U28035 (N_28035,N_27776,N_27901);
nor U28036 (N_28036,N_27766,N_27800);
xnor U28037 (N_28037,N_27836,N_27844);
nor U28038 (N_28038,N_27834,N_27979);
nand U28039 (N_28039,N_27799,N_27831);
nor U28040 (N_28040,N_27854,N_27767);
xnor U28041 (N_28041,N_27804,N_27957);
or U28042 (N_28042,N_27839,N_27961);
xnor U28043 (N_28043,N_27784,N_27835);
nand U28044 (N_28044,N_27778,N_27795);
xor U28045 (N_28045,N_27917,N_27898);
nand U28046 (N_28046,N_27875,N_27966);
nor U28047 (N_28047,N_27933,N_27946);
xor U28048 (N_28048,N_27765,N_27845);
nand U28049 (N_28049,N_27863,N_27769);
and U28050 (N_28050,N_27825,N_27897);
and U28051 (N_28051,N_27807,N_27913);
or U28052 (N_28052,N_27932,N_27828);
and U28053 (N_28053,N_27787,N_27811);
or U28054 (N_28054,N_27838,N_27753);
and U28055 (N_28055,N_27903,N_27949);
or U28056 (N_28056,N_27890,N_27960);
nor U28057 (N_28057,N_27964,N_27853);
xor U28058 (N_28058,N_27794,N_27851);
nand U28059 (N_28059,N_27874,N_27859);
or U28060 (N_28060,N_27916,N_27873);
xnor U28061 (N_28061,N_27919,N_27809);
and U28062 (N_28062,N_27981,N_27783);
xnor U28063 (N_28063,N_27758,N_27796);
nor U28064 (N_28064,N_27770,N_27755);
and U28065 (N_28065,N_27914,N_27921);
nand U28066 (N_28066,N_27892,N_27888);
nand U28067 (N_28067,N_27881,N_27902);
nor U28068 (N_28068,N_27959,N_27904);
nor U28069 (N_28069,N_27761,N_27999);
nor U28070 (N_28070,N_27991,N_27936);
xnor U28071 (N_28071,N_27947,N_27840);
nand U28072 (N_28072,N_27958,N_27833);
or U28073 (N_28073,N_27970,N_27791);
nand U28074 (N_28074,N_27968,N_27763);
or U28075 (N_28075,N_27963,N_27808);
nor U28076 (N_28076,N_27889,N_27855);
and U28077 (N_28077,N_27884,N_27792);
or U28078 (N_28078,N_27948,N_27927);
and U28079 (N_28079,N_27907,N_27975);
or U28080 (N_28080,N_27985,N_27860);
nand U28081 (N_28081,N_27955,N_27909);
nand U28082 (N_28082,N_27945,N_27956);
or U28083 (N_28083,N_27923,N_27935);
or U28084 (N_28084,N_27969,N_27918);
or U28085 (N_28085,N_27894,N_27939);
and U28086 (N_28086,N_27857,N_27777);
nand U28087 (N_28087,N_27974,N_27864);
nand U28088 (N_28088,N_27986,N_27774);
nor U28089 (N_28089,N_27982,N_27994);
or U28090 (N_28090,N_27806,N_27841);
nand U28091 (N_28091,N_27950,N_27871);
or U28092 (N_28092,N_27905,N_27786);
nand U28093 (N_28093,N_27879,N_27983);
nand U28094 (N_28094,N_27843,N_27988);
or U28095 (N_28095,N_27865,N_27869);
nand U28096 (N_28096,N_27866,N_27876);
xor U28097 (N_28097,N_27842,N_27962);
nand U28098 (N_28098,N_27997,N_27996);
and U28099 (N_28099,N_27822,N_27847);
nor U28100 (N_28100,N_27827,N_27837);
nand U28101 (N_28101,N_27810,N_27850);
or U28102 (N_28102,N_27995,N_27922);
or U28103 (N_28103,N_27830,N_27829);
or U28104 (N_28104,N_27987,N_27912);
xnor U28105 (N_28105,N_27877,N_27990);
and U28106 (N_28106,N_27849,N_27891);
or U28107 (N_28107,N_27856,N_27938);
nor U28108 (N_28108,N_27911,N_27814);
xor U28109 (N_28109,N_27773,N_27883);
and U28110 (N_28110,N_27872,N_27993);
or U28111 (N_28111,N_27943,N_27951);
xnor U28112 (N_28112,N_27821,N_27893);
nand U28113 (N_28113,N_27817,N_27754);
and U28114 (N_28114,N_27818,N_27781);
and U28115 (N_28115,N_27900,N_27780);
xor U28116 (N_28116,N_27846,N_27826);
nor U28117 (N_28117,N_27789,N_27992);
or U28118 (N_28118,N_27998,N_27924);
nand U28119 (N_28119,N_27954,N_27926);
xor U28120 (N_28120,N_27929,N_27858);
and U28121 (N_28121,N_27937,N_27978);
or U28122 (N_28122,N_27984,N_27762);
xor U28123 (N_28123,N_27823,N_27896);
and U28124 (N_28124,N_27895,N_27934);
or U28125 (N_28125,N_27866,N_27861);
nor U28126 (N_28126,N_27938,N_27964);
nand U28127 (N_28127,N_27929,N_27942);
xor U28128 (N_28128,N_27874,N_27811);
xnor U28129 (N_28129,N_27977,N_27763);
xnor U28130 (N_28130,N_27806,N_27867);
xnor U28131 (N_28131,N_27855,N_27907);
or U28132 (N_28132,N_27873,N_27945);
nor U28133 (N_28133,N_27969,N_27834);
xnor U28134 (N_28134,N_27809,N_27987);
xor U28135 (N_28135,N_27876,N_27972);
or U28136 (N_28136,N_27918,N_27865);
nand U28137 (N_28137,N_27872,N_27970);
or U28138 (N_28138,N_27842,N_27880);
nand U28139 (N_28139,N_27952,N_27792);
and U28140 (N_28140,N_27975,N_27957);
and U28141 (N_28141,N_27772,N_27811);
nor U28142 (N_28142,N_27835,N_27960);
xnor U28143 (N_28143,N_27941,N_27840);
and U28144 (N_28144,N_27990,N_27907);
nand U28145 (N_28145,N_27811,N_27893);
and U28146 (N_28146,N_27768,N_27875);
nand U28147 (N_28147,N_27868,N_27875);
or U28148 (N_28148,N_27882,N_27907);
or U28149 (N_28149,N_27773,N_27804);
nand U28150 (N_28150,N_27864,N_27834);
nor U28151 (N_28151,N_27801,N_27791);
or U28152 (N_28152,N_27966,N_27932);
xor U28153 (N_28153,N_27853,N_27984);
or U28154 (N_28154,N_27923,N_27957);
nor U28155 (N_28155,N_27932,N_27976);
nor U28156 (N_28156,N_27958,N_27767);
nor U28157 (N_28157,N_27754,N_27921);
xor U28158 (N_28158,N_27771,N_27972);
nor U28159 (N_28159,N_27902,N_27820);
or U28160 (N_28160,N_27769,N_27854);
nor U28161 (N_28161,N_27935,N_27776);
nand U28162 (N_28162,N_27916,N_27850);
xnor U28163 (N_28163,N_27769,N_27834);
nand U28164 (N_28164,N_27898,N_27759);
or U28165 (N_28165,N_27752,N_27998);
nand U28166 (N_28166,N_27816,N_27942);
nor U28167 (N_28167,N_27882,N_27968);
and U28168 (N_28168,N_27854,N_27750);
or U28169 (N_28169,N_27959,N_27797);
nand U28170 (N_28170,N_27997,N_27796);
nand U28171 (N_28171,N_27753,N_27783);
or U28172 (N_28172,N_27933,N_27886);
nor U28173 (N_28173,N_27948,N_27962);
or U28174 (N_28174,N_27786,N_27954);
nor U28175 (N_28175,N_27789,N_27869);
and U28176 (N_28176,N_27759,N_27792);
nand U28177 (N_28177,N_27775,N_27962);
nand U28178 (N_28178,N_27865,N_27985);
nand U28179 (N_28179,N_27972,N_27890);
or U28180 (N_28180,N_27808,N_27980);
or U28181 (N_28181,N_27819,N_27938);
or U28182 (N_28182,N_27917,N_27871);
xor U28183 (N_28183,N_27825,N_27909);
xor U28184 (N_28184,N_27884,N_27995);
xor U28185 (N_28185,N_27914,N_27828);
or U28186 (N_28186,N_27885,N_27754);
nor U28187 (N_28187,N_27979,N_27907);
and U28188 (N_28188,N_27985,N_27841);
nor U28189 (N_28189,N_27889,N_27872);
and U28190 (N_28190,N_27909,N_27945);
xnor U28191 (N_28191,N_27801,N_27928);
nor U28192 (N_28192,N_27813,N_27823);
and U28193 (N_28193,N_27886,N_27828);
and U28194 (N_28194,N_27839,N_27993);
and U28195 (N_28195,N_27774,N_27758);
or U28196 (N_28196,N_27792,N_27966);
nor U28197 (N_28197,N_27791,N_27960);
xnor U28198 (N_28198,N_27809,N_27863);
nor U28199 (N_28199,N_27840,N_27885);
xnor U28200 (N_28200,N_27995,N_27987);
and U28201 (N_28201,N_27965,N_27973);
or U28202 (N_28202,N_27769,N_27852);
or U28203 (N_28203,N_27860,N_27925);
nand U28204 (N_28204,N_27896,N_27768);
and U28205 (N_28205,N_27800,N_27849);
and U28206 (N_28206,N_27965,N_27926);
or U28207 (N_28207,N_27850,N_27884);
or U28208 (N_28208,N_27928,N_27839);
and U28209 (N_28209,N_27816,N_27962);
and U28210 (N_28210,N_27927,N_27905);
nor U28211 (N_28211,N_27847,N_27957);
and U28212 (N_28212,N_27836,N_27924);
or U28213 (N_28213,N_27877,N_27858);
or U28214 (N_28214,N_27871,N_27867);
and U28215 (N_28215,N_27858,N_27911);
and U28216 (N_28216,N_27765,N_27973);
nand U28217 (N_28217,N_27816,N_27980);
and U28218 (N_28218,N_27854,N_27836);
nand U28219 (N_28219,N_27809,N_27975);
nand U28220 (N_28220,N_27925,N_27961);
nand U28221 (N_28221,N_27982,N_27845);
and U28222 (N_28222,N_27891,N_27763);
xor U28223 (N_28223,N_27840,N_27889);
nand U28224 (N_28224,N_27824,N_27931);
and U28225 (N_28225,N_27960,N_27916);
xnor U28226 (N_28226,N_27777,N_27934);
nor U28227 (N_28227,N_27797,N_27940);
nor U28228 (N_28228,N_27930,N_27840);
or U28229 (N_28229,N_27785,N_27946);
and U28230 (N_28230,N_27841,N_27760);
xnor U28231 (N_28231,N_27757,N_27988);
and U28232 (N_28232,N_27797,N_27956);
nor U28233 (N_28233,N_27802,N_27807);
nor U28234 (N_28234,N_27936,N_27850);
and U28235 (N_28235,N_27996,N_27998);
nand U28236 (N_28236,N_27905,N_27777);
nand U28237 (N_28237,N_27835,N_27865);
or U28238 (N_28238,N_27787,N_27789);
xor U28239 (N_28239,N_27965,N_27873);
and U28240 (N_28240,N_27879,N_27926);
or U28241 (N_28241,N_27906,N_27828);
nor U28242 (N_28242,N_27961,N_27959);
or U28243 (N_28243,N_27844,N_27817);
nand U28244 (N_28244,N_27902,N_27792);
and U28245 (N_28245,N_27755,N_27966);
or U28246 (N_28246,N_27907,N_27973);
nand U28247 (N_28247,N_27825,N_27792);
nand U28248 (N_28248,N_27940,N_27980);
nor U28249 (N_28249,N_27985,N_27863);
and U28250 (N_28250,N_28050,N_28216);
nand U28251 (N_28251,N_28037,N_28177);
and U28252 (N_28252,N_28209,N_28100);
nor U28253 (N_28253,N_28185,N_28132);
nor U28254 (N_28254,N_28093,N_28052);
or U28255 (N_28255,N_28241,N_28155);
and U28256 (N_28256,N_28181,N_28017);
nand U28257 (N_28257,N_28114,N_28152);
nand U28258 (N_28258,N_28023,N_28171);
nor U28259 (N_28259,N_28194,N_28053);
and U28260 (N_28260,N_28046,N_28073);
xnor U28261 (N_28261,N_28128,N_28071);
xnor U28262 (N_28262,N_28215,N_28163);
or U28263 (N_28263,N_28217,N_28158);
or U28264 (N_28264,N_28011,N_28248);
xor U28265 (N_28265,N_28089,N_28218);
or U28266 (N_28266,N_28153,N_28244);
or U28267 (N_28267,N_28124,N_28120);
xnor U28268 (N_28268,N_28129,N_28198);
and U28269 (N_28269,N_28015,N_28166);
xnor U28270 (N_28270,N_28201,N_28234);
or U28271 (N_28271,N_28055,N_28059);
or U28272 (N_28272,N_28227,N_28121);
nor U28273 (N_28273,N_28006,N_28139);
or U28274 (N_28274,N_28080,N_28156);
xnor U28275 (N_28275,N_28150,N_28001);
nand U28276 (N_28276,N_28200,N_28187);
and U28277 (N_28277,N_28178,N_28033);
xnor U28278 (N_28278,N_28056,N_28179);
nor U28279 (N_28279,N_28136,N_28028);
nor U28280 (N_28280,N_28126,N_28088);
xnor U28281 (N_28281,N_28009,N_28000);
and U28282 (N_28282,N_28054,N_28110);
and U28283 (N_28283,N_28151,N_28229);
xnor U28284 (N_28284,N_28210,N_28233);
nor U28285 (N_28285,N_28197,N_28096);
xor U28286 (N_28286,N_28008,N_28095);
and U28287 (N_28287,N_28122,N_28167);
or U28288 (N_28288,N_28098,N_28228);
nand U28289 (N_28289,N_28224,N_28208);
or U28290 (N_28290,N_28212,N_28221);
and U28291 (N_28291,N_28143,N_28131);
or U28292 (N_28292,N_28020,N_28076);
nor U28293 (N_28293,N_28002,N_28094);
nand U28294 (N_28294,N_28077,N_28026);
or U28295 (N_28295,N_28149,N_28063);
nor U28296 (N_28296,N_28174,N_28083);
or U28297 (N_28297,N_28070,N_28159);
xnor U28298 (N_28298,N_28051,N_28188);
nand U28299 (N_28299,N_28082,N_28106);
and U28300 (N_28300,N_28142,N_28115);
or U28301 (N_28301,N_28062,N_28160);
nor U28302 (N_28302,N_28192,N_28065);
nand U28303 (N_28303,N_28214,N_28117);
nor U28304 (N_28304,N_28084,N_28223);
nor U28305 (N_28305,N_28225,N_28048);
nand U28306 (N_28306,N_28213,N_28005);
nor U28307 (N_28307,N_28147,N_28134);
xnor U28308 (N_28308,N_28183,N_28058);
nor U28309 (N_28309,N_28034,N_28186);
xor U28310 (N_28310,N_28101,N_28220);
or U28311 (N_28311,N_28184,N_28113);
xor U28312 (N_28312,N_28003,N_28108);
or U28313 (N_28313,N_28014,N_28109);
or U28314 (N_28314,N_28049,N_28041);
and U28315 (N_28315,N_28067,N_28164);
nor U28316 (N_28316,N_28099,N_28104);
xnor U28317 (N_28317,N_28190,N_28045);
nand U28318 (N_28318,N_28086,N_28138);
nand U28319 (N_28319,N_28111,N_28107);
or U28320 (N_28320,N_28091,N_28146);
nor U28321 (N_28321,N_28105,N_28237);
nand U28322 (N_28322,N_28247,N_28127);
and U28323 (N_28323,N_28019,N_28075);
and U28324 (N_28324,N_28203,N_28024);
xor U28325 (N_28325,N_28144,N_28030);
and U28326 (N_28326,N_28137,N_28061);
xor U28327 (N_28327,N_28079,N_28066);
nor U28328 (N_28328,N_28141,N_28157);
nand U28329 (N_28329,N_28010,N_28012);
nor U28330 (N_28330,N_28044,N_28236);
nand U28331 (N_28331,N_28195,N_28118);
xor U28332 (N_28332,N_28211,N_28004);
nor U28333 (N_28333,N_28145,N_28140);
or U28334 (N_28334,N_28222,N_28205);
or U28335 (N_28335,N_28199,N_28087);
nor U28336 (N_28336,N_28074,N_28047);
nand U28337 (N_28337,N_28206,N_28173);
nor U28338 (N_28338,N_28246,N_28172);
or U28339 (N_28339,N_28018,N_28043);
nand U28340 (N_28340,N_28239,N_28112);
nand U28341 (N_28341,N_28240,N_28231);
nor U28342 (N_28342,N_28238,N_28007);
nand U28343 (N_28343,N_28175,N_28202);
nand U28344 (N_28344,N_28085,N_28021);
xor U28345 (N_28345,N_28170,N_28097);
and U28346 (N_28346,N_28090,N_28176);
nor U28347 (N_28347,N_28032,N_28013);
xnor U28348 (N_28348,N_28064,N_28092);
nand U28349 (N_28349,N_28249,N_28103);
or U28350 (N_28350,N_28072,N_28029);
or U28351 (N_28351,N_28207,N_28165);
nor U28352 (N_28352,N_28069,N_28035);
nand U28353 (N_28353,N_28230,N_28189);
and U28354 (N_28354,N_28161,N_28204);
or U28355 (N_28355,N_28042,N_28169);
nand U28356 (N_28356,N_28119,N_28022);
and U28357 (N_28357,N_28036,N_28027);
or U28358 (N_28358,N_28123,N_28078);
or U28359 (N_28359,N_28116,N_28040);
or U28360 (N_28360,N_28154,N_28245);
and U28361 (N_28361,N_28196,N_28219);
xnor U28362 (N_28362,N_28243,N_28060);
or U28363 (N_28363,N_28102,N_28016);
nand U28364 (N_28364,N_28135,N_28242);
or U28365 (N_28365,N_28232,N_28191);
xor U28366 (N_28366,N_28038,N_28193);
nand U28367 (N_28367,N_28133,N_28025);
xnor U28368 (N_28368,N_28125,N_28031);
and U28369 (N_28369,N_28130,N_28162);
and U28370 (N_28370,N_28057,N_28182);
and U28371 (N_28371,N_28180,N_28226);
and U28372 (N_28372,N_28235,N_28148);
nor U28373 (N_28373,N_28039,N_28168);
or U28374 (N_28374,N_28068,N_28081);
and U28375 (N_28375,N_28037,N_28179);
xnor U28376 (N_28376,N_28086,N_28007);
and U28377 (N_28377,N_28019,N_28170);
or U28378 (N_28378,N_28044,N_28056);
nand U28379 (N_28379,N_28164,N_28043);
nor U28380 (N_28380,N_28066,N_28170);
xor U28381 (N_28381,N_28100,N_28123);
and U28382 (N_28382,N_28150,N_28024);
nor U28383 (N_28383,N_28173,N_28005);
xor U28384 (N_28384,N_28150,N_28214);
xor U28385 (N_28385,N_28235,N_28073);
and U28386 (N_28386,N_28073,N_28237);
nor U28387 (N_28387,N_28067,N_28245);
nor U28388 (N_28388,N_28052,N_28115);
xnor U28389 (N_28389,N_28206,N_28001);
and U28390 (N_28390,N_28070,N_28077);
or U28391 (N_28391,N_28222,N_28085);
xnor U28392 (N_28392,N_28091,N_28180);
and U28393 (N_28393,N_28232,N_28097);
and U28394 (N_28394,N_28062,N_28059);
or U28395 (N_28395,N_28210,N_28020);
and U28396 (N_28396,N_28213,N_28113);
nand U28397 (N_28397,N_28037,N_28238);
and U28398 (N_28398,N_28197,N_28160);
nand U28399 (N_28399,N_28031,N_28190);
xor U28400 (N_28400,N_28072,N_28234);
nand U28401 (N_28401,N_28176,N_28198);
and U28402 (N_28402,N_28098,N_28064);
nand U28403 (N_28403,N_28223,N_28043);
xor U28404 (N_28404,N_28227,N_28129);
and U28405 (N_28405,N_28206,N_28035);
nand U28406 (N_28406,N_28212,N_28215);
and U28407 (N_28407,N_28244,N_28121);
nand U28408 (N_28408,N_28120,N_28212);
xnor U28409 (N_28409,N_28228,N_28172);
xor U28410 (N_28410,N_28033,N_28132);
nor U28411 (N_28411,N_28034,N_28233);
xnor U28412 (N_28412,N_28229,N_28209);
nor U28413 (N_28413,N_28144,N_28233);
nand U28414 (N_28414,N_28225,N_28129);
xnor U28415 (N_28415,N_28127,N_28182);
nor U28416 (N_28416,N_28201,N_28092);
nand U28417 (N_28417,N_28084,N_28218);
xor U28418 (N_28418,N_28217,N_28008);
nor U28419 (N_28419,N_28148,N_28193);
nor U28420 (N_28420,N_28094,N_28106);
xor U28421 (N_28421,N_28062,N_28091);
and U28422 (N_28422,N_28132,N_28190);
or U28423 (N_28423,N_28173,N_28000);
and U28424 (N_28424,N_28057,N_28213);
or U28425 (N_28425,N_28051,N_28169);
and U28426 (N_28426,N_28001,N_28088);
nand U28427 (N_28427,N_28091,N_28179);
nand U28428 (N_28428,N_28138,N_28081);
xor U28429 (N_28429,N_28071,N_28218);
nand U28430 (N_28430,N_28008,N_28110);
nand U28431 (N_28431,N_28113,N_28146);
xor U28432 (N_28432,N_28172,N_28155);
nand U28433 (N_28433,N_28146,N_28187);
nand U28434 (N_28434,N_28092,N_28169);
xnor U28435 (N_28435,N_28010,N_28044);
nand U28436 (N_28436,N_28167,N_28029);
xor U28437 (N_28437,N_28216,N_28188);
nand U28438 (N_28438,N_28239,N_28011);
xnor U28439 (N_28439,N_28120,N_28084);
nand U28440 (N_28440,N_28072,N_28023);
xor U28441 (N_28441,N_28139,N_28053);
nand U28442 (N_28442,N_28071,N_28092);
xor U28443 (N_28443,N_28072,N_28011);
or U28444 (N_28444,N_28187,N_28199);
nor U28445 (N_28445,N_28080,N_28228);
xnor U28446 (N_28446,N_28068,N_28138);
or U28447 (N_28447,N_28040,N_28218);
and U28448 (N_28448,N_28113,N_28207);
xnor U28449 (N_28449,N_28170,N_28036);
nand U28450 (N_28450,N_28148,N_28245);
and U28451 (N_28451,N_28092,N_28156);
xor U28452 (N_28452,N_28088,N_28219);
nor U28453 (N_28453,N_28144,N_28211);
nand U28454 (N_28454,N_28102,N_28066);
and U28455 (N_28455,N_28177,N_28058);
nand U28456 (N_28456,N_28214,N_28093);
and U28457 (N_28457,N_28206,N_28012);
xnor U28458 (N_28458,N_28080,N_28130);
xor U28459 (N_28459,N_28088,N_28182);
and U28460 (N_28460,N_28097,N_28191);
nand U28461 (N_28461,N_28091,N_28199);
xor U28462 (N_28462,N_28139,N_28197);
and U28463 (N_28463,N_28003,N_28016);
and U28464 (N_28464,N_28224,N_28171);
and U28465 (N_28465,N_28066,N_28237);
or U28466 (N_28466,N_28110,N_28103);
nand U28467 (N_28467,N_28167,N_28194);
xor U28468 (N_28468,N_28017,N_28061);
xnor U28469 (N_28469,N_28028,N_28044);
nor U28470 (N_28470,N_28082,N_28232);
xnor U28471 (N_28471,N_28134,N_28176);
nor U28472 (N_28472,N_28135,N_28131);
or U28473 (N_28473,N_28194,N_28026);
or U28474 (N_28474,N_28009,N_28125);
or U28475 (N_28475,N_28103,N_28140);
xor U28476 (N_28476,N_28155,N_28006);
nand U28477 (N_28477,N_28092,N_28004);
or U28478 (N_28478,N_28074,N_28214);
and U28479 (N_28479,N_28083,N_28227);
xor U28480 (N_28480,N_28194,N_28241);
or U28481 (N_28481,N_28061,N_28247);
and U28482 (N_28482,N_28210,N_28050);
nand U28483 (N_28483,N_28045,N_28080);
nor U28484 (N_28484,N_28064,N_28248);
nor U28485 (N_28485,N_28122,N_28163);
nor U28486 (N_28486,N_28044,N_28184);
and U28487 (N_28487,N_28100,N_28141);
or U28488 (N_28488,N_28042,N_28036);
xnor U28489 (N_28489,N_28168,N_28214);
or U28490 (N_28490,N_28239,N_28077);
or U28491 (N_28491,N_28098,N_28061);
nand U28492 (N_28492,N_28004,N_28064);
xor U28493 (N_28493,N_28109,N_28164);
nor U28494 (N_28494,N_28107,N_28031);
nand U28495 (N_28495,N_28025,N_28218);
nor U28496 (N_28496,N_28086,N_28201);
nor U28497 (N_28497,N_28030,N_28098);
or U28498 (N_28498,N_28133,N_28131);
nand U28499 (N_28499,N_28009,N_28146);
nand U28500 (N_28500,N_28315,N_28388);
or U28501 (N_28501,N_28371,N_28497);
nand U28502 (N_28502,N_28290,N_28333);
xnor U28503 (N_28503,N_28412,N_28307);
nand U28504 (N_28504,N_28498,N_28303);
or U28505 (N_28505,N_28357,N_28366);
xor U28506 (N_28506,N_28422,N_28443);
nand U28507 (N_28507,N_28255,N_28479);
or U28508 (N_28508,N_28386,N_28337);
nand U28509 (N_28509,N_28458,N_28400);
and U28510 (N_28510,N_28302,N_28346);
nand U28511 (N_28511,N_28253,N_28446);
nor U28512 (N_28512,N_28439,N_28477);
or U28513 (N_28513,N_28352,N_28392);
and U28514 (N_28514,N_28276,N_28384);
or U28515 (N_28515,N_28360,N_28490);
xor U28516 (N_28516,N_28430,N_28327);
xnor U28517 (N_28517,N_28285,N_28317);
and U28518 (N_28518,N_28372,N_28408);
and U28519 (N_28519,N_28274,N_28453);
or U28520 (N_28520,N_28311,N_28266);
and U28521 (N_28521,N_28326,N_28358);
and U28522 (N_28522,N_28454,N_28420);
nor U28523 (N_28523,N_28319,N_28341);
nand U28524 (N_28524,N_28278,N_28434);
nand U28525 (N_28525,N_28464,N_28322);
and U28526 (N_28526,N_28273,N_28316);
nand U28527 (N_28527,N_28272,N_28288);
or U28528 (N_28528,N_28297,N_28277);
or U28529 (N_28529,N_28336,N_28398);
nand U28530 (N_28530,N_28472,N_28414);
xnor U28531 (N_28531,N_28381,N_28335);
and U28532 (N_28532,N_28495,N_28413);
nor U28533 (N_28533,N_28283,N_28329);
nand U28534 (N_28534,N_28451,N_28361);
nor U28535 (N_28535,N_28262,N_28339);
xor U28536 (N_28536,N_28314,N_28416);
nor U28537 (N_28537,N_28362,N_28499);
nand U28538 (N_28538,N_28353,N_28407);
nand U28539 (N_28539,N_28456,N_28296);
or U28540 (N_28540,N_28305,N_28265);
xor U28541 (N_28541,N_28279,N_28258);
nand U28542 (N_28542,N_28375,N_28462);
or U28543 (N_28543,N_28435,N_28478);
and U28544 (N_28544,N_28496,N_28251);
and U28545 (N_28545,N_28461,N_28349);
xnor U28546 (N_28546,N_28468,N_28481);
or U28547 (N_28547,N_28440,N_28489);
or U28548 (N_28548,N_28394,N_28321);
xor U28549 (N_28549,N_28488,N_28356);
nor U28550 (N_28550,N_28399,N_28491);
and U28551 (N_28551,N_28294,N_28330);
nor U28552 (N_28552,N_28493,N_28484);
xnor U28553 (N_28553,N_28445,N_28494);
and U28554 (N_28554,N_28259,N_28318);
nor U28555 (N_28555,N_28291,N_28415);
nand U28556 (N_28556,N_28482,N_28402);
xnor U28557 (N_28557,N_28382,N_28355);
and U28558 (N_28558,N_28264,N_28368);
xnor U28559 (N_28559,N_28250,N_28448);
or U28560 (N_28560,N_28282,N_28338);
nand U28561 (N_28561,N_28359,N_28469);
xnor U28562 (N_28562,N_28260,N_28404);
nand U28563 (N_28563,N_28252,N_28310);
nand U28564 (N_28564,N_28347,N_28410);
xor U28565 (N_28565,N_28261,N_28483);
xnor U28566 (N_28566,N_28377,N_28292);
or U28567 (N_28567,N_28289,N_28401);
nand U28568 (N_28568,N_28450,N_28268);
or U28569 (N_28569,N_28431,N_28390);
or U28570 (N_28570,N_28396,N_28363);
or U28571 (N_28571,N_28423,N_28471);
or U28572 (N_28572,N_28345,N_28441);
xor U28573 (N_28573,N_28373,N_28295);
xor U28574 (N_28574,N_28269,N_28304);
xnor U28575 (N_28575,N_28470,N_28455);
and U28576 (N_28576,N_28286,N_28300);
and U28577 (N_28577,N_28417,N_28449);
nor U28578 (N_28578,N_28348,N_28328);
xnor U28579 (N_28579,N_28301,N_28391);
nand U28580 (N_28580,N_28320,N_28428);
and U28581 (N_28581,N_28308,N_28480);
nand U28582 (N_28582,N_28460,N_28473);
and U28583 (N_28583,N_28299,N_28267);
xor U28584 (N_28584,N_28343,N_28436);
xor U28585 (N_28585,N_28351,N_28485);
nand U28586 (N_28586,N_28406,N_28324);
and U28587 (N_28587,N_28452,N_28486);
nand U28588 (N_28588,N_28340,N_28271);
xor U28589 (N_28589,N_28447,N_28306);
and U28590 (N_28590,N_28444,N_28332);
nor U28591 (N_28591,N_28331,N_28395);
nor U28592 (N_28592,N_28393,N_28463);
xnor U28593 (N_28593,N_28312,N_28378);
xnor U28594 (N_28594,N_28442,N_28424);
and U28595 (N_28595,N_28379,N_28280);
or U28596 (N_28596,N_28437,N_28364);
or U28597 (N_28597,N_28284,N_28459);
or U28598 (N_28598,N_28344,N_28487);
xor U28599 (N_28599,N_28293,N_28387);
nor U28600 (N_28600,N_28342,N_28474);
nand U28601 (N_28601,N_28275,N_28403);
nor U28602 (N_28602,N_28257,N_28323);
xor U28603 (N_28603,N_28397,N_28425);
xnor U28604 (N_28604,N_28254,N_28438);
nor U28605 (N_28605,N_28256,N_28354);
and U28606 (N_28606,N_28476,N_28475);
or U28607 (N_28607,N_28365,N_28465);
xnor U28608 (N_28608,N_28457,N_28426);
and U28609 (N_28609,N_28287,N_28427);
nand U28610 (N_28610,N_28421,N_28263);
nor U28611 (N_28611,N_28405,N_28492);
or U28612 (N_28612,N_28369,N_28380);
or U28613 (N_28613,N_28411,N_28429);
nand U28614 (N_28614,N_28433,N_28298);
nand U28615 (N_28615,N_28409,N_28313);
nor U28616 (N_28616,N_28270,N_28350);
xor U28617 (N_28617,N_28367,N_28385);
nand U28618 (N_28618,N_28418,N_28467);
and U28619 (N_28619,N_28466,N_28389);
and U28620 (N_28620,N_28374,N_28419);
xor U28621 (N_28621,N_28383,N_28334);
nand U28622 (N_28622,N_28376,N_28281);
and U28623 (N_28623,N_28432,N_28370);
xor U28624 (N_28624,N_28325,N_28309);
xor U28625 (N_28625,N_28446,N_28250);
xnor U28626 (N_28626,N_28299,N_28284);
nand U28627 (N_28627,N_28283,N_28322);
nand U28628 (N_28628,N_28330,N_28469);
nor U28629 (N_28629,N_28323,N_28470);
xnor U28630 (N_28630,N_28420,N_28272);
and U28631 (N_28631,N_28397,N_28406);
xor U28632 (N_28632,N_28393,N_28441);
and U28633 (N_28633,N_28490,N_28334);
xor U28634 (N_28634,N_28274,N_28257);
and U28635 (N_28635,N_28468,N_28336);
xor U28636 (N_28636,N_28382,N_28493);
or U28637 (N_28637,N_28456,N_28313);
nor U28638 (N_28638,N_28491,N_28262);
xor U28639 (N_28639,N_28431,N_28391);
xor U28640 (N_28640,N_28492,N_28422);
nor U28641 (N_28641,N_28290,N_28252);
or U28642 (N_28642,N_28403,N_28470);
nor U28643 (N_28643,N_28402,N_28440);
and U28644 (N_28644,N_28349,N_28478);
xnor U28645 (N_28645,N_28450,N_28442);
nor U28646 (N_28646,N_28416,N_28343);
and U28647 (N_28647,N_28365,N_28415);
and U28648 (N_28648,N_28377,N_28403);
nand U28649 (N_28649,N_28482,N_28412);
nor U28650 (N_28650,N_28281,N_28480);
xnor U28651 (N_28651,N_28279,N_28401);
nand U28652 (N_28652,N_28438,N_28304);
nand U28653 (N_28653,N_28445,N_28427);
xor U28654 (N_28654,N_28383,N_28327);
or U28655 (N_28655,N_28462,N_28451);
or U28656 (N_28656,N_28374,N_28320);
nand U28657 (N_28657,N_28290,N_28374);
nor U28658 (N_28658,N_28254,N_28286);
nand U28659 (N_28659,N_28314,N_28350);
nand U28660 (N_28660,N_28473,N_28288);
and U28661 (N_28661,N_28279,N_28260);
xnor U28662 (N_28662,N_28413,N_28431);
nor U28663 (N_28663,N_28346,N_28392);
nand U28664 (N_28664,N_28426,N_28439);
xnor U28665 (N_28665,N_28470,N_28256);
nor U28666 (N_28666,N_28298,N_28326);
or U28667 (N_28667,N_28354,N_28317);
or U28668 (N_28668,N_28270,N_28308);
nor U28669 (N_28669,N_28322,N_28434);
or U28670 (N_28670,N_28424,N_28376);
and U28671 (N_28671,N_28446,N_28353);
nand U28672 (N_28672,N_28440,N_28459);
xor U28673 (N_28673,N_28294,N_28368);
and U28674 (N_28674,N_28270,N_28393);
xnor U28675 (N_28675,N_28287,N_28406);
xnor U28676 (N_28676,N_28360,N_28411);
and U28677 (N_28677,N_28379,N_28468);
and U28678 (N_28678,N_28410,N_28348);
or U28679 (N_28679,N_28250,N_28342);
xor U28680 (N_28680,N_28299,N_28318);
and U28681 (N_28681,N_28326,N_28340);
nand U28682 (N_28682,N_28444,N_28484);
nand U28683 (N_28683,N_28260,N_28345);
and U28684 (N_28684,N_28362,N_28318);
nor U28685 (N_28685,N_28489,N_28375);
nor U28686 (N_28686,N_28472,N_28356);
and U28687 (N_28687,N_28355,N_28346);
nor U28688 (N_28688,N_28393,N_28287);
or U28689 (N_28689,N_28487,N_28401);
and U28690 (N_28690,N_28359,N_28471);
nor U28691 (N_28691,N_28460,N_28435);
nor U28692 (N_28692,N_28417,N_28479);
xor U28693 (N_28693,N_28358,N_28376);
nor U28694 (N_28694,N_28291,N_28292);
nor U28695 (N_28695,N_28440,N_28447);
and U28696 (N_28696,N_28415,N_28417);
xor U28697 (N_28697,N_28394,N_28411);
xor U28698 (N_28698,N_28261,N_28495);
or U28699 (N_28699,N_28347,N_28358);
and U28700 (N_28700,N_28323,N_28284);
and U28701 (N_28701,N_28361,N_28298);
nand U28702 (N_28702,N_28397,N_28367);
nand U28703 (N_28703,N_28434,N_28255);
or U28704 (N_28704,N_28358,N_28252);
nand U28705 (N_28705,N_28361,N_28283);
nand U28706 (N_28706,N_28475,N_28421);
xnor U28707 (N_28707,N_28373,N_28329);
and U28708 (N_28708,N_28278,N_28369);
or U28709 (N_28709,N_28277,N_28348);
nor U28710 (N_28710,N_28355,N_28277);
or U28711 (N_28711,N_28329,N_28426);
and U28712 (N_28712,N_28456,N_28301);
nor U28713 (N_28713,N_28265,N_28269);
nor U28714 (N_28714,N_28389,N_28472);
or U28715 (N_28715,N_28444,N_28469);
and U28716 (N_28716,N_28288,N_28433);
or U28717 (N_28717,N_28324,N_28327);
and U28718 (N_28718,N_28447,N_28251);
xnor U28719 (N_28719,N_28434,N_28477);
nor U28720 (N_28720,N_28398,N_28328);
or U28721 (N_28721,N_28375,N_28365);
xnor U28722 (N_28722,N_28469,N_28273);
xnor U28723 (N_28723,N_28480,N_28425);
or U28724 (N_28724,N_28320,N_28471);
and U28725 (N_28725,N_28348,N_28301);
nand U28726 (N_28726,N_28267,N_28337);
or U28727 (N_28727,N_28446,N_28402);
and U28728 (N_28728,N_28276,N_28444);
nand U28729 (N_28729,N_28400,N_28392);
or U28730 (N_28730,N_28266,N_28356);
nand U28731 (N_28731,N_28461,N_28483);
and U28732 (N_28732,N_28265,N_28349);
nand U28733 (N_28733,N_28475,N_28268);
or U28734 (N_28734,N_28384,N_28436);
xor U28735 (N_28735,N_28323,N_28399);
nand U28736 (N_28736,N_28361,N_28413);
xor U28737 (N_28737,N_28285,N_28496);
or U28738 (N_28738,N_28275,N_28404);
and U28739 (N_28739,N_28286,N_28368);
nor U28740 (N_28740,N_28369,N_28305);
xor U28741 (N_28741,N_28355,N_28272);
nand U28742 (N_28742,N_28342,N_28324);
nand U28743 (N_28743,N_28316,N_28368);
xnor U28744 (N_28744,N_28465,N_28260);
and U28745 (N_28745,N_28422,N_28280);
or U28746 (N_28746,N_28422,N_28259);
xnor U28747 (N_28747,N_28330,N_28327);
nor U28748 (N_28748,N_28458,N_28387);
or U28749 (N_28749,N_28419,N_28384);
nand U28750 (N_28750,N_28540,N_28741);
xor U28751 (N_28751,N_28576,N_28570);
nand U28752 (N_28752,N_28569,N_28608);
xnor U28753 (N_28753,N_28738,N_28505);
and U28754 (N_28754,N_28676,N_28714);
nand U28755 (N_28755,N_28749,N_28597);
nor U28756 (N_28756,N_28709,N_28510);
xor U28757 (N_28757,N_28737,N_28643);
nand U28758 (N_28758,N_28698,N_28504);
and U28759 (N_28759,N_28582,N_28558);
nand U28760 (N_28760,N_28736,N_28673);
xor U28761 (N_28761,N_28630,N_28546);
or U28762 (N_28762,N_28583,N_28631);
and U28763 (N_28763,N_28634,N_28713);
nand U28764 (N_28764,N_28685,N_28694);
or U28765 (N_28765,N_28719,N_28571);
nor U28766 (N_28766,N_28620,N_28729);
or U28767 (N_28767,N_28657,N_28588);
nor U28768 (N_28768,N_28573,N_28579);
or U28769 (N_28769,N_28644,N_28521);
xor U28770 (N_28770,N_28642,N_28535);
nand U28771 (N_28771,N_28598,N_28735);
nand U28772 (N_28772,N_28740,N_28522);
nand U28773 (N_28773,N_28675,N_28525);
xnor U28774 (N_28774,N_28528,N_28635);
xor U28775 (N_28775,N_28523,N_28697);
xor U28776 (N_28776,N_28653,N_28515);
nand U28777 (N_28777,N_28672,N_28640);
or U28778 (N_28778,N_28671,N_28686);
nand U28779 (N_28779,N_28744,N_28746);
or U28780 (N_28780,N_28708,N_28556);
nor U28781 (N_28781,N_28734,N_28659);
and U28782 (N_28782,N_28724,N_28606);
nor U28783 (N_28783,N_28629,N_28661);
xor U28784 (N_28784,N_28649,N_28710);
nand U28785 (N_28785,N_28628,N_28706);
nor U28786 (N_28786,N_28575,N_28516);
xnor U28787 (N_28787,N_28555,N_28632);
or U28788 (N_28788,N_28539,N_28536);
or U28789 (N_28789,N_28548,N_28626);
nand U28790 (N_28790,N_28589,N_28615);
nor U28791 (N_28791,N_28503,N_28660);
nand U28792 (N_28792,N_28645,N_28586);
or U28793 (N_28793,N_28511,N_28502);
xnor U28794 (N_28794,N_28611,N_28532);
and U28795 (N_28795,N_28731,N_28529);
or U28796 (N_28796,N_28509,N_28739);
and U28797 (N_28797,N_28715,N_28531);
nor U28798 (N_28798,N_28607,N_28692);
nand U28799 (N_28799,N_28595,N_28552);
xor U28800 (N_28800,N_28633,N_28567);
nor U28801 (N_28801,N_28530,N_28553);
nand U28802 (N_28802,N_28602,N_28683);
nand U28803 (N_28803,N_28512,N_28604);
nor U28804 (N_28804,N_28679,N_28636);
and U28805 (N_28805,N_28517,N_28500);
and U28806 (N_28806,N_28674,N_28668);
and U28807 (N_28807,N_28725,N_28748);
xor U28808 (N_28808,N_28591,N_28616);
xor U28809 (N_28809,N_28614,N_28665);
and U28810 (N_28810,N_28732,N_28681);
nand U28811 (N_28811,N_28705,N_28701);
nor U28812 (N_28812,N_28652,N_28551);
nand U28813 (N_28813,N_28663,N_28609);
nor U28814 (N_28814,N_28689,N_28621);
nor U28815 (N_28815,N_28574,N_28585);
or U28816 (N_28816,N_28599,N_28596);
nand U28817 (N_28817,N_28541,N_28581);
nor U28818 (N_28818,N_28678,N_28742);
nor U28819 (N_28819,N_28610,N_28519);
xor U28820 (N_28820,N_28688,N_28712);
nor U28821 (N_28821,N_28584,N_28545);
or U28822 (N_28822,N_28594,N_28730);
nand U28823 (N_28823,N_28613,N_28533);
xor U28824 (N_28824,N_28508,N_28646);
and U28825 (N_28825,N_28538,N_28580);
and U28826 (N_28826,N_28721,N_28718);
nand U28827 (N_28827,N_28695,N_28703);
or U28828 (N_28828,N_28641,N_28702);
or U28829 (N_28829,N_28654,N_28572);
nor U28830 (N_28830,N_28560,N_28527);
xnor U28831 (N_28831,N_28648,N_28603);
and U28832 (N_28832,N_28664,N_28514);
nor U28833 (N_28833,N_28578,N_28524);
nor U28834 (N_28834,N_28720,N_28566);
xor U28835 (N_28835,N_28537,N_28650);
or U28836 (N_28836,N_28728,N_28534);
nor U28837 (N_28837,N_28651,N_28617);
nor U28838 (N_28838,N_28550,N_28690);
or U28839 (N_28839,N_28513,N_28745);
or U28840 (N_28840,N_28587,N_28726);
or U28841 (N_28841,N_28590,N_28623);
or U28842 (N_28842,N_28563,N_28704);
nor U28843 (N_28843,N_28562,N_28559);
nor U28844 (N_28844,N_28627,N_28677);
nand U28845 (N_28845,N_28707,N_28684);
and U28846 (N_28846,N_28600,N_28687);
and U28847 (N_28847,N_28662,N_28625);
xnor U28848 (N_28848,N_28542,N_28543);
or U28849 (N_28849,N_28693,N_28507);
nand U28850 (N_28850,N_28592,N_28544);
and U28851 (N_28851,N_28612,N_28547);
and U28852 (N_28852,N_28669,N_28624);
and U28853 (N_28853,N_28639,N_28743);
nor U28854 (N_28854,N_28622,N_28554);
nor U28855 (N_28855,N_28637,N_28501);
xor U28856 (N_28856,N_28722,N_28618);
or U28857 (N_28857,N_28518,N_28506);
nand U28858 (N_28858,N_28655,N_28717);
xor U28859 (N_28859,N_28747,N_28565);
nor U28860 (N_28860,N_28561,N_28619);
xor U28861 (N_28861,N_28733,N_28577);
xnor U28862 (N_28862,N_28670,N_28667);
or U28863 (N_28863,N_28716,N_28680);
and U28864 (N_28864,N_28557,N_28696);
xnor U28865 (N_28865,N_28605,N_28568);
nand U28866 (N_28866,N_28711,N_28601);
xor U28867 (N_28867,N_28666,N_28564);
and U28868 (N_28868,N_28658,N_28700);
and U28869 (N_28869,N_28656,N_28691);
nand U28870 (N_28870,N_28593,N_28638);
xor U28871 (N_28871,N_28727,N_28699);
nand U28872 (N_28872,N_28549,N_28647);
nand U28873 (N_28873,N_28520,N_28526);
or U28874 (N_28874,N_28723,N_28682);
and U28875 (N_28875,N_28555,N_28506);
nand U28876 (N_28876,N_28692,N_28621);
nor U28877 (N_28877,N_28690,N_28588);
and U28878 (N_28878,N_28678,N_28713);
xnor U28879 (N_28879,N_28749,N_28585);
or U28880 (N_28880,N_28529,N_28735);
xnor U28881 (N_28881,N_28548,N_28748);
or U28882 (N_28882,N_28725,N_28551);
or U28883 (N_28883,N_28529,N_28515);
or U28884 (N_28884,N_28623,N_28579);
nand U28885 (N_28885,N_28605,N_28502);
or U28886 (N_28886,N_28640,N_28528);
or U28887 (N_28887,N_28740,N_28729);
or U28888 (N_28888,N_28684,N_28714);
xnor U28889 (N_28889,N_28678,N_28515);
or U28890 (N_28890,N_28606,N_28575);
and U28891 (N_28891,N_28609,N_28707);
and U28892 (N_28892,N_28702,N_28579);
nor U28893 (N_28893,N_28663,N_28700);
nand U28894 (N_28894,N_28741,N_28743);
or U28895 (N_28895,N_28562,N_28613);
xor U28896 (N_28896,N_28647,N_28582);
and U28897 (N_28897,N_28714,N_28700);
or U28898 (N_28898,N_28726,N_28516);
or U28899 (N_28899,N_28670,N_28739);
and U28900 (N_28900,N_28629,N_28539);
or U28901 (N_28901,N_28645,N_28542);
nor U28902 (N_28902,N_28501,N_28524);
or U28903 (N_28903,N_28608,N_28739);
and U28904 (N_28904,N_28511,N_28701);
xnor U28905 (N_28905,N_28741,N_28688);
or U28906 (N_28906,N_28626,N_28672);
nand U28907 (N_28907,N_28736,N_28668);
nor U28908 (N_28908,N_28581,N_28719);
or U28909 (N_28909,N_28667,N_28591);
nand U28910 (N_28910,N_28694,N_28706);
nand U28911 (N_28911,N_28597,N_28576);
nand U28912 (N_28912,N_28526,N_28637);
and U28913 (N_28913,N_28634,N_28686);
or U28914 (N_28914,N_28730,N_28569);
nor U28915 (N_28915,N_28704,N_28728);
nand U28916 (N_28916,N_28567,N_28681);
nand U28917 (N_28917,N_28569,N_28524);
and U28918 (N_28918,N_28646,N_28681);
xor U28919 (N_28919,N_28665,N_28615);
nor U28920 (N_28920,N_28618,N_28620);
nand U28921 (N_28921,N_28665,N_28526);
nor U28922 (N_28922,N_28656,N_28693);
or U28923 (N_28923,N_28618,N_28666);
xnor U28924 (N_28924,N_28698,N_28640);
xnor U28925 (N_28925,N_28698,N_28599);
xor U28926 (N_28926,N_28506,N_28690);
or U28927 (N_28927,N_28743,N_28723);
or U28928 (N_28928,N_28646,N_28529);
or U28929 (N_28929,N_28581,N_28665);
nand U28930 (N_28930,N_28747,N_28667);
xor U28931 (N_28931,N_28512,N_28637);
xor U28932 (N_28932,N_28617,N_28729);
xnor U28933 (N_28933,N_28676,N_28740);
or U28934 (N_28934,N_28723,N_28627);
nand U28935 (N_28935,N_28511,N_28519);
xor U28936 (N_28936,N_28711,N_28511);
nor U28937 (N_28937,N_28711,N_28561);
xnor U28938 (N_28938,N_28569,N_28727);
or U28939 (N_28939,N_28575,N_28709);
and U28940 (N_28940,N_28732,N_28737);
xor U28941 (N_28941,N_28570,N_28543);
and U28942 (N_28942,N_28547,N_28669);
or U28943 (N_28943,N_28580,N_28570);
or U28944 (N_28944,N_28564,N_28575);
nor U28945 (N_28945,N_28572,N_28510);
or U28946 (N_28946,N_28512,N_28521);
xor U28947 (N_28947,N_28525,N_28732);
or U28948 (N_28948,N_28654,N_28664);
nand U28949 (N_28949,N_28668,N_28656);
nand U28950 (N_28950,N_28512,N_28695);
nand U28951 (N_28951,N_28571,N_28677);
nand U28952 (N_28952,N_28598,N_28714);
nor U28953 (N_28953,N_28606,N_28681);
or U28954 (N_28954,N_28641,N_28640);
xnor U28955 (N_28955,N_28639,N_28725);
and U28956 (N_28956,N_28703,N_28501);
nor U28957 (N_28957,N_28641,N_28569);
nand U28958 (N_28958,N_28724,N_28590);
nand U28959 (N_28959,N_28602,N_28676);
xor U28960 (N_28960,N_28697,N_28529);
nor U28961 (N_28961,N_28559,N_28663);
nor U28962 (N_28962,N_28598,N_28704);
or U28963 (N_28963,N_28540,N_28660);
or U28964 (N_28964,N_28729,N_28513);
and U28965 (N_28965,N_28603,N_28626);
and U28966 (N_28966,N_28554,N_28621);
nand U28967 (N_28967,N_28536,N_28724);
or U28968 (N_28968,N_28690,N_28606);
nor U28969 (N_28969,N_28606,N_28609);
or U28970 (N_28970,N_28562,N_28665);
and U28971 (N_28971,N_28628,N_28566);
and U28972 (N_28972,N_28601,N_28668);
xnor U28973 (N_28973,N_28541,N_28559);
nand U28974 (N_28974,N_28510,N_28670);
xor U28975 (N_28975,N_28580,N_28713);
nand U28976 (N_28976,N_28590,N_28663);
xor U28977 (N_28977,N_28671,N_28665);
xor U28978 (N_28978,N_28537,N_28665);
nand U28979 (N_28979,N_28509,N_28628);
and U28980 (N_28980,N_28567,N_28607);
or U28981 (N_28981,N_28686,N_28640);
and U28982 (N_28982,N_28542,N_28617);
or U28983 (N_28983,N_28654,N_28557);
nand U28984 (N_28984,N_28546,N_28573);
nand U28985 (N_28985,N_28699,N_28648);
nor U28986 (N_28986,N_28598,N_28662);
nand U28987 (N_28987,N_28616,N_28610);
and U28988 (N_28988,N_28649,N_28593);
nand U28989 (N_28989,N_28575,N_28661);
nor U28990 (N_28990,N_28661,N_28605);
or U28991 (N_28991,N_28591,N_28549);
or U28992 (N_28992,N_28662,N_28685);
nand U28993 (N_28993,N_28724,N_28624);
and U28994 (N_28994,N_28659,N_28504);
nand U28995 (N_28995,N_28505,N_28610);
nor U28996 (N_28996,N_28667,N_28598);
xnor U28997 (N_28997,N_28521,N_28643);
nand U28998 (N_28998,N_28674,N_28525);
nand U28999 (N_28999,N_28501,N_28533);
nor U29000 (N_29000,N_28936,N_28980);
or U29001 (N_29001,N_28792,N_28803);
and U29002 (N_29002,N_28893,N_28890);
and U29003 (N_29003,N_28884,N_28965);
xor U29004 (N_29004,N_28881,N_28998);
and U29005 (N_29005,N_28943,N_28789);
nor U29006 (N_29006,N_28925,N_28960);
nor U29007 (N_29007,N_28759,N_28798);
nor U29008 (N_29008,N_28904,N_28988);
xnor U29009 (N_29009,N_28915,N_28986);
nand U29010 (N_29010,N_28838,N_28973);
nor U29011 (N_29011,N_28877,N_28836);
nor U29012 (N_29012,N_28773,N_28996);
nand U29013 (N_29013,N_28945,N_28796);
nor U29014 (N_29014,N_28833,N_28958);
or U29015 (N_29015,N_28782,N_28847);
or U29016 (N_29016,N_28811,N_28897);
nor U29017 (N_29017,N_28829,N_28917);
xor U29018 (N_29018,N_28757,N_28860);
and U29019 (N_29019,N_28822,N_28856);
nor U29020 (N_29020,N_28933,N_28812);
or U29021 (N_29021,N_28935,N_28823);
and U29022 (N_29022,N_28774,N_28941);
nand U29023 (N_29023,N_28889,N_28862);
nand U29024 (N_29024,N_28837,N_28895);
or U29025 (N_29025,N_28871,N_28934);
and U29026 (N_29026,N_28835,N_28995);
and U29027 (N_29027,N_28850,N_28880);
or U29028 (N_29028,N_28928,N_28769);
xor U29029 (N_29029,N_28857,N_28826);
xor U29030 (N_29030,N_28954,N_28852);
xnor U29031 (N_29031,N_28962,N_28765);
and U29032 (N_29032,N_28808,N_28939);
nand U29033 (N_29033,N_28964,N_28882);
xnor U29034 (N_29034,N_28914,N_28911);
nand U29035 (N_29035,N_28899,N_28799);
and U29036 (N_29036,N_28907,N_28787);
and U29037 (N_29037,N_28987,N_28815);
and U29038 (N_29038,N_28931,N_28824);
and U29039 (N_29039,N_28976,N_28961);
xnor U29040 (N_29040,N_28758,N_28948);
or U29041 (N_29041,N_28763,N_28870);
and U29042 (N_29042,N_28989,N_28866);
nand U29043 (N_29043,N_28861,N_28818);
or U29044 (N_29044,N_28752,N_28817);
xor U29045 (N_29045,N_28992,N_28854);
nor U29046 (N_29046,N_28993,N_28896);
xnor U29047 (N_29047,N_28971,N_28806);
nand U29048 (N_29048,N_28977,N_28903);
and U29049 (N_29049,N_28937,N_28793);
nor U29050 (N_29050,N_28885,N_28924);
nor U29051 (N_29051,N_28950,N_28846);
or U29052 (N_29052,N_28766,N_28968);
nand U29053 (N_29053,N_28900,N_28839);
xnor U29054 (N_29054,N_28983,N_28804);
and U29055 (N_29055,N_28784,N_28786);
xor U29056 (N_29056,N_28938,N_28946);
nor U29057 (N_29057,N_28775,N_28865);
and U29058 (N_29058,N_28843,N_28827);
and U29059 (N_29059,N_28790,N_28832);
xnor U29060 (N_29060,N_28794,N_28819);
nand U29061 (N_29061,N_28791,N_28970);
or U29062 (N_29062,N_28929,N_28873);
nor U29063 (N_29063,N_28947,N_28779);
nand U29064 (N_29064,N_28898,N_28869);
nor U29065 (N_29065,N_28888,N_28825);
xor U29066 (N_29066,N_28920,N_28783);
xor U29067 (N_29067,N_28767,N_28919);
nand U29068 (N_29068,N_28800,N_28966);
or U29069 (N_29069,N_28830,N_28840);
nor U29070 (N_29070,N_28776,N_28875);
nand U29071 (N_29071,N_28864,N_28777);
or U29072 (N_29072,N_28756,N_28762);
xor U29073 (N_29073,N_28849,N_28879);
and U29074 (N_29074,N_28807,N_28994);
or U29075 (N_29075,N_28750,N_28778);
nor U29076 (N_29076,N_28878,N_28886);
xnor U29077 (N_29077,N_28760,N_28801);
and U29078 (N_29078,N_28972,N_28932);
xnor U29079 (N_29079,N_28788,N_28772);
or U29080 (N_29080,N_28926,N_28955);
and U29081 (N_29081,N_28809,N_28802);
and U29082 (N_29082,N_28816,N_28979);
or U29083 (N_29083,N_28883,N_28953);
or U29084 (N_29084,N_28867,N_28959);
or U29085 (N_29085,N_28909,N_28927);
xor U29086 (N_29086,N_28813,N_28906);
xnor U29087 (N_29087,N_28834,N_28785);
nand U29088 (N_29088,N_28753,N_28910);
or U29089 (N_29089,N_28751,N_28923);
and U29090 (N_29090,N_28863,N_28999);
xnor U29091 (N_29091,N_28894,N_28872);
or U29092 (N_29092,N_28952,N_28761);
or U29093 (N_29093,N_28975,N_28918);
or U29094 (N_29094,N_28805,N_28892);
and U29095 (N_29095,N_28951,N_28991);
nand U29096 (N_29096,N_28940,N_28902);
xnor U29097 (N_29097,N_28922,N_28853);
or U29098 (N_29098,N_28957,N_28795);
xnor U29099 (N_29099,N_28810,N_28944);
nor U29100 (N_29100,N_28990,N_28887);
nor U29101 (N_29101,N_28981,N_28985);
or U29102 (N_29102,N_28814,N_28755);
or U29103 (N_29103,N_28874,N_28912);
or U29104 (N_29104,N_28764,N_28754);
nand U29105 (N_29105,N_28967,N_28820);
nand U29106 (N_29106,N_28771,N_28916);
nand U29107 (N_29107,N_28891,N_28876);
and U29108 (N_29108,N_28770,N_28921);
xnor U29109 (N_29109,N_28913,N_28949);
nand U29110 (N_29110,N_28841,N_28831);
nand U29111 (N_29111,N_28978,N_28781);
or U29112 (N_29112,N_28768,N_28908);
nand U29113 (N_29113,N_28974,N_28797);
and U29114 (N_29114,N_28930,N_28901);
or U29115 (N_29115,N_28969,N_28868);
or U29116 (N_29116,N_28942,N_28821);
xnor U29117 (N_29117,N_28828,N_28844);
or U29118 (N_29118,N_28845,N_28997);
xor U29119 (N_29119,N_28963,N_28905);
and U29120 (N_29120,N_28859,N_28858);
nand U29121 (N_29121,N_28956,N_28851);
nor U29122 (N_29122,N_28982,N_28855);
and U29123 (N_29123,N_28848,N_28780);
or U29124 (N_29124,N_28984,N_28842);
xor U29125 (N_29125,N_28932,N_28923);
nand U29126 (N_29126,N_28852,N_28877);
nor U29127 (N_29127,N_28927,N_28888);
nand U29128 (N_29128,N_28932,N_28988);
or U29129 (N_29129,N_28816,N_28868);
nor U29130 (N_29130,N_28907,N_28784);
or U29131 (N_29131,N_28973,N_28850);
or U29132 (N_29132,N_28992,N_28760);
nor U29133 (N_29133,N_28799,N_28836);
nor U29134 (N_29134,N_28797,N_28968);
nor U29135 (N_29135,N_28917,N_28945);
nor U29136 (N_29136,N_28838,N_28763);
or U29137 (N_29137,N_28926,N_28944);
xnor U29138 (N_29138,N_28952,N_28905);
and U29139 (N_29139,N_28814,N_28771);
and U29140 (N_29140,N_28911,N_28868);
nand U29141 (N_29141,N_28916,N_28867);
and U29142 (N_29142,N_28931,N_28926);
nor U29143 (N_29143,N_28826,N_28765);
and U29144 (N_29144,N_28839,N_28952);
nor U29145 (N_29145,N_28774,N_28761);
and U29146 (N_29146,N_28786,N_28781);
xor U29147 (N_29147,N_28958,N_28935);
nor U29148 (N_29148,N_28860,N_28892);
nand U29149 (N_29149,N_28931,N_28850);
xnor U29150 (N_29150,N_28992,N_28890);
and U29151 (N_29151,N_28912,N_28779);
or U29152 (N_29152,N_28900,N_28966);
or U29153 (N_29153,N_28972,N_28951);
or U29154 (N_29154,N_28769,N_28796);
and U29155 (N_29155,N_28925,N_28951);
nand U29156 (N_29156,N_28832,N_28775);
xnor U29157 (N_29157,N_28998,N_28826);
or U29158 (N_29158,N_28865,N_28814);
xor U29159 (N_29159,N_28758,N_28786);
or U29160 (N_29160,N_28981,N_28957);
and U29161 (N_29161,N_28996,N_28827);
or U29162 (N_29162,N_28952,N_28825);
nand U29163 (N_29163,N_28811,N_28760);
nor U29164 (N_29164,N_28776,N_28924);
or U29165 (N_29165,N_28831,N_28805);
and U29166 (N_29166,N_28887,N_28807);
nor U29167 (N_29167,N_28844,N_28904);
nand U29168 (N_29168,N_28771,N_28887);
or U29169 (N_29169,N_28945,N_28944);
or U29170 (N_29170,N_28849,N_28810);
nor U29171 (N_29171,N_28815,N_28790);
xnor U29172 (N_29172,N_28822,N_28931);
or U29173 (N_29173,N_28892,N_28959);
nand U29174 (N_29174,N_28941,N_28844);
or U29175 (N_29175,N_28850,N_28758);
nor U29176 (N_29176,N_28964,N_28871);
or U29177 (N_29177,N_28989,N_28971);
and U29178 (N_29178,N_28941,N_28905);
or U29179 (N_29179,N_28937,N_28765);
xor U29180 (N_29180,N_28773,N_28876);
and U29181 (N_29181,N_28918,N_28951);
nor U29182 (N_29182,N_28778,N_28942);
xnor U29183 (N_29183,N_28861,N_28982);
nand U29184 (N_29184,N_28931,N_28984);
or U29185 (N_29185,N_28762,N_28974);
xor U29186 (N_29186,N_28942,N_28855);
and U29187 (N_29187,N_28828,N_28948);
xor U29188 (N_29188,N_28962,N_28763);
nand U29189 (N_29189,N_28987,N_28802);
xor U29190 (N_29190,N_28812,N_28940);
nor U29191 (N_29191,N_28839,N_28853);
nor U29192 (N_29192,N_28812,N_28885);
or U29193 (N_29193,N_28958,N_28760);
nor U29194 (N_29194,N_28925,N_28831);
and U29195 (N_29195,N_28803,N_28920);
nor U29196 (N_29196,N_28896,N_28980);
and U29197 (N_29197,N_28934,N_28760);
and U29198 (N_29198,N_28863,N_28948);
xor U29199 (N_29199,N_28758,N_28844);
or U29200 (N_29200,N_28989,N_28777);
or U29201 (N_29201,N_28768,N_28955);
and U29202 (N_29202,N_28957,N_28985);
nor U29203 (N_29203,N_28901,N_28762);
and U29204 (N_29204,N_28911,N_28989);
and U29205 (N_29205,N_28778,N_28931);
or U29206 (N_29206,N_28985,N_28838);
and U29207 (N_29207,N_28770,N_28806);
or U29208 (N_29208,N_28780,N_28930);
xnor U29209 (N_29209,N_28763,N_28939);
and U29210 (N_29210,N_28885,N_28856);
nor U29211 (N_29211,N_28947,N_28801);
nand U29212 (N_29212,N_28937,N_28956);
nor U29213 (N_29213,N_28760,N_28975);
nand U29214 (N_29214,N_28892,N_28936);
or U29215 (N_29215,N_28893,N_28771);
nand U29216 (N_29216,N_28754,N_28900);
nor U29217 (N_29217,N_28882,N_28927);
or U29218 (N_29218,N_28888,N_28850);
or U29219 (N_29219,N_28838,N_28847);
xor U29220 (N_29220,N_28771,N_28928);
nor U29221 (N_29221,N_28802,N_28856);
nand U29222 (N_29222,N_28790,N_28773);
nand U29223 (N_29223,N_28867,N_28951);
or U29224 (N_29224,N_28821,N_28983);
and U29225 (N_29225,N_28839,N_28942);
nor U29226 (N_29226,N_28993,N_28847);
or U29227 (N_29227,N_28832,N_28922);
nor U29228 (N_29228,N_28766,N_28833);
xnor U29229 (N_29229,N_28772,N_28952);
xor U29230 (N_29230,N_28820,N_28837);
nand U29231 (N_29231,N_28974,N_28914);
or U29232 (N_29232,N_28901,N_28861);
nor U29233 (N_29233,N_28780,N_28827);
xor U29234 (N_29234,N_28864,N_28964);
nand U29235 (N_29235,N_28874,N_28872);
nor U29236 (N_29236,N_28883,N_28826);
and U29237 (N_29237,N_28849,N_28861);
and U29238 (N_29238,N_28778,N_28910);
and U29239 (N_29239,N_28873,N_28920);
xnor U29240 (N_29240,N_28950,N_28753);
nor U29241 (N_29241,N_28950,N_28768);
and U29242 (N_29242,N_28950,N_28966);
xnor U29243 (N_29243,N_28775,N_28837);
xor U29244 (N_29244,N_28993,N_28967);
nor U29245 (N_29245,N_28780,N_28902);
or U29246 (N_29246,N_28760,N_28796);
nand U29247 (N_29247,N_28840,N_28957);
or U29248 (N_29248,N_28912,N_28908);
or U29249 (N_29249,N_28845,N_28913);
and U29250 (N_29250,N_29246,N_29089);
or U29251 (N_29251,N_29190,N_29195);
and U29252 (N_29252,N_29088,N_29124);
and U29253 (N_29253,N_29078,N_29063);
and U29254 (N_29254,N_29097,N_29093);
and U29255 (N_29255,N_29162,N_29056);
nand U29256 (N_29256,N_29073,N_29134);
xnor U29257 (N_29257,N_29053,N_29083);
xor U29258 (N_29258,N_29198,N_29248);
nor U29259 (N_29259,N_29171,N_29103);
nand U29260 (N_29260,N_29080,N_29173);
xor U29261 (N_29261,N_29081,N_29242);
nand U29262 (N_29262,N_29021,N_29002);
nor U29263 (N_29263,N_29033,N_29241);
xor U29264 (N_29264,N_29031,N_29028);
and U29265 (N_29265,N_29090,N_29102);
nand U29266 (N_29266,N_29163,N_29064);
nand U29267 (N_29267,N_29015,N_29219);
nor U29268 (N_29268,N_29147,N_29038);
or U29269 (N_29269,N_29127,N_29239);
xor U29270 (N_29270,N_29023,N_29245);
nand U29271 (N_29271,N_29112,N_29184);
and U29272 (N_29272,N_29186,N_29010);
nand U29273 (N_29273,N_29049,N_29019);
and U29274 (N_29274,N_29111,N_29125);
or U29275 (N_29275,N_29249,N_29065);
and U29276 (N_29276,N_29176,N_29243);
and U29277 (N_29277,N_29217,N_29116);
or U29278 (N_29278,N_29157,N_29223);
and U29279 (N_29279,N_29043,N_29143);
nor U29280 (N_29280,N_29183,N_29235);
nor U29281 (N_29281,N_29177,N_29085);
or U29282 (N_29282,N_29032,N_29206);
nand U29283 (N_29283,N_29213,N_29165);
or U29284 (N_29284,N_29231,N_29040);
or U29285 (N_29285,N_29120,N_29109);
and U29286 (N_29286,N_29188,N_29192);
nor U29287 (N_29287,N_29168,N_29045);
nand U29288 (N_29288,N_29185,N_29018);
and U29289 (N_29289,N_29092,N_29114);
xor U29290 (N_29290,N_29175,N_29204);
and U29291 (N_29291,N_29121,N_29167);
xor U29292 (N_29292,N_29054,N_29087);
nor U29293 (N_29293,N_29156,N_29164);
and U29294 (N_29294,N_29137,N_29237);
xor U29295 (N_29295,N_29196,N_29075);
xnor U29296 (N_29296,N_29071,N_29230);
nand U29297 (N_29297,N_29179,N_29142);
nor U29298 (N_29298,N_29225,N_29050);
xnor U29299 (N_29299,N_29158,N_29170);
nor U29300 (N_29300,N_29100,N_29036);
xnor U29301 (N_29301,N_29153,N_29210);
or U29302 (N_29302,N_29070,N_29013);
nand U29303 (N_29303,N_29079,N_29145);
and U29304 (N_29304,N_29154,N_29232);
xnor U29305 (N_29305,N_29006,N_29020);
or U29306 (N_29306,N_29069,N_29205);
or U29307 (N_29307,N_29151,N_29024);
or U29308 (N_29308,N_29214,N_29123);
xnor U29309 (N_29309,N_29039,N_29076);
or U29310 (N_29310,N_29193,N_29030);
xor U29311 (N_29311,N_29149,N_29110);
or U29312 (N_29312,N_29104,N_29060);
nand U29313 (N_29313,N_29201,N_29001);
nand U29314 (N_29314,N_29128,N_29048);
nand U29315 (N_29315,N_29209,N_29099);
and U29316 (N_29316,N_29191,N_29000);
or U29317 (N_29317,N_29215,N_29224);
nor U29318 (N_29318,N_29062,N_29199);
nor U29319 (N_29319,N_29055,N_29234);
nor U29320 (N_29320,N_29026,N_29159);
nand U29321 (N_29321,N_29052,N_29095);
and U29322 (N_29322,N_29057,N_29135);
nand U29323 (N_29323,N_29084,N_29150);
or U29324 (N_29324,N_29007,N_29059);
and U29325 (N_29325,N_29227,N_29203);
nand U29326 (N_29326,N_29220,N_29106);
or U29327 (N_29327,N_29148,N_29197);
xnor U29328 (N_29328,N_29037,N_29034);
xor U29329 (N_29329,N_29202,N_29136);
xnor U29330 (N_29330,N_29117,N_29161);
nor U29331 (N_29331,N_29025,N_29094);
xor U29332 (N_29332,N_29221,N_29181);
and U29333 (N_29333,N_29118,N_29035);
and U29334 (N_29334,N_29014,N_29132);
nor U29335 (N_29335,N_29126,N_29003);
nand U29336 (N_29336,N_29096,N_29009);
and U29337 (N_29337,N_29022,N_29077);
nand U29338 (N_29338,N_29155,N_29130);
nand U29339 (N_29339,N_29172,N_29194);
xnor U29340 (N_29340,N_29180,N_29067);
nor U29341 (N_29341,N_29041,N_29119);
or U29342 (N_29342,N_29140,N_29240);
xor U29343 (N_29343,N_29046,N_29228);
xnor U29344 (N_29344,N_29146,N_29011);
or U29345 (N_29345,N_29105,N_29004);
and U29346 (N_29346,N_29218,N_29101);
nand U29347 (N_29347,N_29017,N_29008);
or U29348 (N_29348,N_29016,N_29222);
or U29349 (N_29349,N_29012,N_29082);
nand U29350 (N_29350,N_29141,N_29061);
nor U29351 (N_29351,N_29027,N_29072);
nor U29352 (N_29352,N_29047,N_29216);
and U29353 (N_29353,N_29108,N_29233);
xor U29354 (N_29354,N_29236,N_29174);
or U29355 (N_29355,N_29166,N_29238);
nand U29356 (N_29356,N_29247,N_29229);
or U29357 (N_29357,N_29144,N_29091);
nor U29358 (N_29358,N_29139,N_29189);
or U29359 (N_29359,N_29044,N_29098);
or U29360 (N_29360,N_29122,N_29115);
or U29361 (N_29361,N_29244,N_29051);
and U29362 (N_29362,N_29029,N_29129);
nand U29363 (N_29363,N_29169,N_29178);
or U29364 (N_29364,N_29200,N_29066);
nand U29365 (N_29365,N_29182,N_29058);
nor U29366 (N_29366,N_29207,N_29212);
nand U29367 (N_29367,N_29138,N_29086);
and U29368 (N_29368,N_29133,N_29131);
nor U29369 (N_29369,N_29211,N_29074);
xor U29370 (N_29370,N_29226,N_29187);
or U29371 (N_29371,N_29160,N_29005);
xnor U29372 (N_29372,N_29208,N_29152);
nor U29373 (N_29373,N_29113,N_29068);
or U29374 (N_29374,N_29107,N_29042);
nand U29375 (N_29375,N_29237,N_29170);
nand U29376 (N_29376,N_29169,N_29092);
and U29377 (N_29377,N_29074,N_29197);
nor U29378 (N_29378,N_29174,N_29180);
xor U29379 (N_29379,N_29224,N_29159);
xnor U29380 (N_29380,N_29084,N_29217);
xnor U29381 (N_29381,N_29140,N_29148);
and U29382 (N_29382,N_29125,N_29216);
xnor U29383 (N_29383,N_29037,N_29096);
and U29384 (N_29384,N_29068,N_29209);
and U29385 (N_29385,N_29139,N_29018);
nand U29386 (N_29386,N_29213,N_29091);
and U29387 (N_29387,N_29164,N_29082);
nor U29388 (N_29388,N_29096,N_29042);
or U29389 (N_29389,N_29120,N_29209);
and U29390 (N_29390,N_29075,N_29025);
xor U29391 (N_29391,N_29036,N_29038);
nor U29392 (N_29392,N_29156,N_29122);
nand U29393 (N_29393,N_29208,N_29162);
nor U29394 (N_29394,N_29204,N_29097);
xnor U29395 (N_29395,N_29162,N_29003);
or U29396 (N_29396,N_29026,N_29043);
xnor U29397 (N_29397,N_29043,N_29102);
and U29398 (N_29398,N_29076,N_29065);
nand U29399 (N_29399,N_29176,N_29043);
nand U29400 (N_29400,N_29063,N_29183);
xor U29401 (N_29401,N_29246,N_29127);
nand U29402 (N_29402,N_29144,N_29131);
or U29403 (N_29403,N_29203,N_29001);
nor U29404 (N_29404,N_29002,N_29222);
xor U29405 (N_29405,N_29013,N_29208);
nand U29406 (N_29406,N_29027,N_29107);
or U29407 (N_29407,N_29150,N_29087);
and U29408 (N_29408,N_29208,N_29183);
nand U29409 (N_29409,N_29174,N_29022);
and U29410 (N_29410,N_29148,N_29082);
nor U29411 (N_29411,N_29240,N_29241);
nor U29412 (N_29412,N_29170,N_29142);
nor U29413 (N_29413,N_29208,N_29101);
nor U29414 (N_29414,N_29123,N_29117);
and U29415 (N_29415,N_29121,N_29036);
nand U29416 (N_29416,N_29024,N_29139);
xnor U29417 (N_29417,N_29018,N_29083);
and U29418 (N_29418,N_29110,N_29097);
and U29419 (N_29419,N_29203,N_29088);
nand U29420 (N_29420,N_29156,N_29036);
or U29421 (N_29421,N_29080,N_29153);
nor U29422 (N_29422,N_29089,N_29113);
nand U29423 (N_29423,N_29145,N_29141);
and U29424 (N_29424,N_29179,N_29089);
and U29425 (N_29425,N_29174,N_29028);
and U29426 (N_29426,N_29235,N_29245);
and U29427 (N_29427,N_29215,N_29130);
nand U29428 (N_29428,N_29096,N_29113);
nor U29429 (N_29429,N_29001,N_29174);
or U29430 (N_29430,N_29009,N_29166);
or U29431 (N_29431,N_29136,N_29161);
or U29432 (N_29432,N_29091,N_29182);
and U29433 (N_29433,N_29015,N_29242);
xnor U29434 (N_29434,N_29017,N_29083);
nand U29435 (N_29435,N_29032,N_29111);
nor U29436 (N_29436,N_29043,N_29220);
and U29437 (N_29437,N_29179,N_29203);
nand U29438 (N_29438,N_29218,N_29060);
xnor U29439 (N_29439,N_29158,N_29114);
nor U29440 (N_29440,N_29093,N_29199);
nand U29441 (N_29441,N_29205,N_29010);
xnor U29442 (N_29442,N_29231,N_29049);
or U29443 (N_29443,N_29102,N_29223);
nand U29444 (N_29444,N_29058,N_29242);
and U29445 (N_29445,N_29168,N_29136);
xnor U29446 (N_29446,N_29092,N_29059);
and U29447 (N_29447,N_29095,N_29042);
nor U29448 (N_29448,N_29171,N_29143);
nand U29449 (N_29449,N_29189,N_29025);
xnor U29450 (N_29450,N_29037,N_29212);
nand U29451 (N_29451,N_29196,N_29121);
xnor U29452 (N_29452,N_29081,N_29034);
or U29453 (N_29453,N_29114,N_29127);
or U29454 (N_29454,N_29206,N_29156);
nand U29455 (N_29455,N_29196,N_29067);
or U29456 (N_29456,N_29012,N_29245);
nor U29457 (N_29457,N_29143,N_29121);
xor U29458 (N_29458,N_29015,N_29052);
nor U29459 (N_29459,N_29128,N_29025);
nor U29460 (N_29460,N_29150,N_29060);
nand U29461 (N_29461,N_29042,N_29103);
xor U29462 (N_29462,N_29151,N_29128);
and U29463 (N_29463,N_29221,N_29025);
xor U29464 (N_29464,N_29225,N_29166);
nor U29465 (N_29465,N_29145,N_29089);
xnor U29466 (N_29466,N_29165,N_29061);
or U29467 (N_29467,N_29038,N_29215);
nand U29468 (N_29468,N_29205,N_29134);
and U29469 (N_29469,N_29109,N_29175);
xor U29470 (N_29470,N_29093,N_29000);
nand U29471 (N_29471,N_29040,N_29134);
nand U29472 (N_29472,N_29111,N_29147);
nor U29473 (N_29473,N_29241,N_29037);
nand U29474 (N_29474,N_29135,N_29036);
or U29475 (N_29475,N_29149,N_29014);
or U29476 (N_29476,N_29139,N_29247);
xnor U29477 (N_29477,N_29183,N_29135);
and U29478 (N_29478,N_29100,N_29227);
nand U29479 (N_29479,N_29178,N_29087);
or U29480 (N_29480,N_29030,N_29029);
xor U29481 (N_29481,N_29032,N_29216);
or U29482 (N_29482,N_29192,N_29114);
xnor U29483 (N_29483,N_29163,N_29188);
nor U29484 (N_29484,N_29062,N_29116);
and U29485 (N_29485,N_29143,N_29126);
nand U29486 (N_29486,N_29221,N_29047);
and U29487 (N_29487,N_29151,N_29045);
and U29488 (N_29488,N_29236,N_29068);
nor U29489 (N_29489,N_29163,N_29013);
and U29490 (N_29490,N_29209,N_29248);
or U29491 (N_29491,N_29225,N_29108);
xnor U29492 (N_29492,N_29226,N_29095);
and U29493 (N_29493,N_29153,N_29098);
and U29494 (N_29494,N_29015,N_29194);
nand U29495 (N_29495,N_29184,N_29247);
xor U29496 (N_29496,N_29166,N_29178);
nand U29497 (N_29497,N_29159,N_29109);
and U29498 (N_29498,N_29076,N_29212);
and U29499 (N_29499,N_29200,N_29059);
or U29500 (N_29500,N_29326,N_29405);
xnor U29501 (N_29501,N_29498,N_29265);
and U29502 (N_29502,N_29475,N_29434);
or U29503 (N_29503,N_29492,N_29357);
nand U29504 (N_29504,N_29483,N_29488);
nor U29505 (N_29505,N_29379,N_29419);
nor U29506 (N_29506,N_29378,N_29410);
nor U29507 (N_29507,N_29325,N_29283);
or U29508 (N_29508,N_29360,N_29340);
xor U29509 (N_29509,N_29396,N_29468);
xnor U29510 (N_29510,N_29438,N_29281);
nor U29511 (N_29511,N_29331,N_29383);
xnor U29512 (N_29512,N_29368,N_29342);
nor U29513 (N_29513,N_29384,N_29258);
and U29514 (N_29514,N_29344,N_29404);
or U29515 (N_29515,N_29428,N_29359);
xnor U29516 (N_29516,N_29278,N_29499);
and U29517 (N_29517,N_29358,N_29470);
nor U29518 (N_29518,N_29361,N_29348);
and U29519 (N_29519,N_29422,N_29469);
nor U29520 (N_29520,N_29286,N_29430);
and U29521 (N_29521,N_29260,N_29320);
nand U29522 (N_29522,N_29427,N_29456);
xor U29523 (N_29523,N_29295,N_29481);
and U29524 (N_29524,N_29352,N_29255);
nor U29525 (N_29525,N_29496,N_29349);
or U29526 (N_29526,N_29392,N_29400);
nand U29527 (N_29527,N_29429,N_29487);
nand U29528 (N_29528,N_29346,N_29312);
nand U29529 (N_29529,N_29339,N_29397);
or U29530 (N_29530,N_29453,N_29341);
nor U29531 (N_29531,N_29332,N_29343);
nor U29532 (N_29532,N_29403,N_29460);
or U29533 (N_29533,N_29280,N_29369);
nand U29534 (N_29534,N_29318,N_29333);
nand U29535 (N_29535,N_29464,N_29374);
nand U29536 (N_29536,N_29347,N_29465);
or U29537 (N_29537,N_29495,N_29304);
xor U29538 (N_29538,N_29375,N_29445);
or U29539 (N_29539,N_29293,N_29267);
nand U29540 (N_29540,N_29380,N_29484);
nand U29541 (N_29541,N_29459,N_29412);
or U29542 (N_29542,N_29313,N_29291);
or U29543 (N_29543,N_29305,N_29406);
nand U29544 (N_29544,N_29310,N_29424);
or U29545 (N_29545,N_29443,N_29376);
nand U29546 (N_29546,N_29282,N_29418);
or U29547 (N_29547,N_29268,N_29448);
xnor U29548 (N_29548,N_29411,N_29393);
or U29549 (N_29549,N_29337,N_29323);
or U29550 (N_29550,N_29275,N_29463);
or U29551 (N_29551,N_29257,N_29261);
xor U29552 (N_29552,N_29319,N_29390);
or U29553 (N_29553,N_29355,N_29446);
and U29554 (N_29554,N_29316,N_29262);
nor U29555 (N_29555,N_29420,N_29287);
nand U29556 (N_29556,N_29253,N_29381);
nand U29557 (N_29557,N_29303,N_29308);
nand U29558 (N_29558,N_29317,N_29285);
nand U29559 (N_29559,N_29284,N_29370);
and U29560 (N_29560,N_29364,N_29389);
xor U29561 (N_29561,N_29417,N_29345);
or U29562 (N_29562,N_29480,N_29299);
or U29563 (N_29563,N_29266,N_29270);
and U29564 (N_29564,N_29482,N_29387);
and U29565 (N_29565,N_29290,N_29415);
xor U29566 (N_29566,N_29479,N_29371);
and U29567 (N_29567,N_29450,N_29321);
xnor U29568 (N_29568,N_29407,N_29431);
xnor U29569 (N_29569,N_29425,N_29372);
xor U29570 (N_29570,N_29367,N_29473);
nand U29571 (N_29571,N_29497,N_29421);
xor U29572 (N_29572,N_29451,N_29276);
nand U29573 (N_29573,N_29489,N_29351);
xnor U29574 (N_29574,N_29277,N_29385);
nand U29575 (N_29575,N_29338,N_29288);
xnor U29576 (N_29576,N_29394,N_29273);
nand U29577 (N_29577,N_29413,N_29478);
nor U29578 (N_29578,N_29435,N_29433);
and U29579 (N_29579,N_29494,N_29442);
xor U29580 (N_29580,N_29272,N_29315);
xor U29581 (N_29581,N_29251,N_29335);
nand U29582 (N_29582,N_29362,N_29455);
and U29583 (N_29583,N_29382,N_29263);
nor U29584 (N_29584,N_29324,N_29327);
xnor U29585 (N_29585,N_29377,N_29329);
nor U29586 (N_29586,N_29426,N_29264);
or U29587 (N_29587,N_29409,N_29471);
xor U29588 (N_29588,N_29458,N_29354);
and U29589 (N_29589,N_29289,N_29423);
and U29590 (N_29590,N_29302,N_29490);
nand U29591 (N_29591,N_29491,N_29300);
or U29592 (N_29592,N_29449,N_29440);
or U29593 (N_29593,N_29356,N_29454);
nand U29594 (N_29594,N_29402,N_29259);
nand U29595 (N_29595,N_29472,N_29322);
and U29596 (N_29596,N_29373,N_29365);
and U29597 (N_29597,N_29269,N_29452);
or U29598 (N_29598,N_29314,N_29432);
nor U29599 (N_29599,N_29476,N_29386);
and U29600 (N_29600,N_29297,N_29467);
xnor U29601 (N_29601,N_29350,N_29493);
nor U29602 (N_29602,N_29466,N_29441);
or U29603 (N_29603,N_29334,N_29485);
or U29604 (N_29604,N_29294,N_29279);
nor U29605 (N_29605,N_29398,N_29296);
and U29606 (N_29606,N_29309,N_29477);
nor U29607 (N_29607,N_29437,N_29457);
nor U29608 (N_29608,N_29271,N_29363);
nand U29609 (N_29609,N_29444,N_29256);
nor U29610 (N_29610,N_29391,N_29395);
xnor U29611 (N_29611,N_29252,N_29462);
nand U29612 (N_29612,N_29292,N_29461);
nor U29613 (N_29613,N_29366,N_29274);
nand U29614 (N_29614,N_29474,N_29336);
xnor U29615 (N_29615,N_29401,N_29439);
and U29616 (N_29616,N_29399,N_29436);
nand U29617 (N_29617,N_29353,N_29328);
xnor U29618 (N_29618,N_29388,N_29298);
and U29619 (N_29619,N_29307,N_29306);
nand U29620 (N_29620,N_29486,N_29330);
nor U29621 (N_29621,N_29416,N_29301);
nand U29622 (N_29622,N_29447,N_29408);
or U29623 (N_29623,N_29311,N_29254);
and U29624 (N_29624,N_29250,N_29414);
or U29625 (N_29625,N_29459,N_29414);
nor U29626 (N_29626,N_29313,N_29318);
xor U29627 (N_29627,N_29364,N_29436);
xor U29628 (N_29628,N_29265,N_29369);
nand U29629 (N_29629,N_29283,N_29256);
nor U29630 (N_29630,N_29289,N_29266);
xor U29631 (N_29631,N_29447,N_29427);
and U29632 (N_29632,N_29425,N_29400);
nor U29633 (N_29633,N_29470,N_29268);
nand U29634 (N_29634,N_29445,N_29412);
xnor U29635 (N_29635,N_29476,N_29392);
and U29636 (N_29636,N_29327,N_29308);
nor U29637 (N_29637,N_29484,N_29279);
or U29638 (N_29638,N_29470,N_29304);
and U29639 (N_29639,N_29477,N_29461);
nand U29640 (N_29640,N_29313,N_29419);
nor U29641 (N_29641,N_29478,N_29358);
and U29642 (N_29642,N_29279,N_29477);
xor U29643 (N_29643,N_29456,N_29382);
nand U29644 (N_29644,N_29269,N_29299);
nor U29645 (N_29645,N_29451,N_29462);
and U29646 (N_29646,N_29375,N_29370);
xnor U29647 (N_29647,N_29293,N_29431);
nor U29648 (N_29648,N_29252,N_29374);
xnor U29649 (N_29649,N_29477,N_29311);
nor U29650 (N_29650,N_29387,N_29434);
nand U29651 (N_29651,N_29259,N_29440);
and U29652 (N_29652,N_29280,N_29467);
xnor U29653 (N_29653,N_29365,N_29343);
or U29654 (N_29654,N_29482,N_29481);
xnor U29655 (N_29655,N_29492,N_29298);
nor U29656 (N_29656,N_29496,N_29266);
nand U29657 (N_29657,N_29367,N_29321);
and U29658 (N_29658,N_29437,N_29471);
or U29659 (N_29659,N_29443,N_29311);
nor U29660 (N_29660,N_29342,N_29479);
xor U29661 (N_29661,N_29334,N_29272);
xor U29662 (N_29662,N_29347,N_29255);
xor U29663 (N_29663,N_29283,N_29445);
xor U29664 (N_29664,N_29421,N_29358);
nor U29665 (N_29665,N_29292,N_29413);
and U29666 (N_29666,N_29340,N_29299);
nor U29667 (N_29667,N_29445,N_29291);
nand U29668 (N_29668,N_29313,N_29255);
xnor U29669 (N_29669,N_29385,N_29284);
or U29670 (N_29670,N_29369,N_29445);
or U29671 (N_29671,N_29475,N_29476);
nand U29672 (N_29672,N_29429,N_29262);
nor U29673 (N_29673,N_29281,N_29428);
nor U29674 (N_29674,N_29374,N_29417);
or U29675 (N_29675,N_29453,N_29360);
xnor U29676 (N_29676,N_29394,N_29434);
and U29677 (N_29677,N_29358,N_29388);
xor U29678 (N_29678,N_29360,N_29467);
or U29679 (N_29679,N_29395,N_29373);
nand U29680 (N_29680,N_29379,N_29461);
nand U29681 (N_29681,N_29342,N_29319);
nand U29682 (N_29682,N_29338,N_29254);
nor U29683 (N_29683,N_29354,N_29391);
or U29684 (N_29684,N_29365,N_29472);
or U29685 (N_29685,N_29362,N_29460);
nor U29686 (N_29686,N_29398,N_29434);
and U29687 (N_29687,N_29403,N_29264);
nor U29688 (N_29688,N_29267,N_29283);
nand U29689 (N_29689,N_29340,N_29479);
nor U29690 (N_29690,N_29415,N_29408);
nor U29691 (N_29691,N_29392,N_29372);
or U29692 (N_29692,N_29432,N_29285);
xnor U29693 (N_29693,N_29368,N_29396);
nand U29694 (N_29694,N_29333,N_29272);
xor U29695 (N_29695,N_29435,N_29389);
nor U29696 (N_29696,N_29465,N_29419);
or U29697 (N_29697,N_29395,N_29433);
nor U29698 (N_29698,N_29378,N_29442);
xor U29699 (N_29699,N_29288,N_29388);
and U29700 (N_29700,N_29438,N_29485);
xnor U29701 (N_29701,N_29335,N_29383);
and U29702 (N_29702,N_29257,N_29305);
xor U29703 (N_29703,N_29335,N_29309);
nor U29704 (N_29704,N_29455,N_29409);
nor U29705 (N_29705,N_29412,N_29383);
nand U29706 (N_29706,N_29310,N_29329);
nor U29707 (N_29707,N_29444,N_29427);
nor U29708 (N_29708,N_29496,N_29396);
or U29709 (N_29709,N_29406,N_29486);
nor U29710 (N_29710,N_29347,N_29402);
nor U29711 (N_29711,N_29496,N_29493);
xor U29712 (N_29712,N_29328,N_29294);
nand U29713 (N_29713,N_29279,N_29296);
or U29714 (N_29714,N_29352,N_29359);
and U29715 (N_29715,N_29444,N_29493);
or U29716 (N_29716,N_29390,N_29432);
nand U29717 (N_29717,N_29455,N_29286);
and U29718 (N_29718,N_29350,N_29272);
nand U29719 (N_29719,N_29386,N_29334);
or U29720 (N_29720,N_29356,N_29416);
and U29721 (N_29721,N_29272,N_29464);
nor U29722 (N_29722,N_29365,N_29459);
nand U29723 (N_29723,N_29399,N_29282);
and U29724 (N_29724,N_29489,N_29445);
nand U29725 (N_29725,N_29374,N_29310);
and U29726 (N_29726,N_29448,N_29429);
and U29727 (N_29727,N_29468,N_29404);
nand U29728 (N_29728,N_29298,N_29255);
and U29729 (N_29729,N_29426,N_29495);
or U29730 (N_29730,N_29302,N_29308);
nand U29731 (N_29731,N_29493,N_29303);
and U29732 (N_29732,N_29356,N_29489);
or U29733 (N_29733,N_29441,N_29358);
or U29734 (N_29734,N_29493,N_29499);
xnor U29735 (N_29735,N_29298,N_29293);
xnor U29736 (N_29736,N_29455,N_29293);
xor U29737 (N_29737,N_29311,N_29434);
xnor U29738 (N_29738,N_29283,N_29379);
or U29739 (N_29739,N_29413,N_29357);
xor U29740 (N_29740,N_29424,N_29460);
nor U29741 (N_29741,N_29431,N_29378);
nor U29742 (N_29742,N_29308,N_29495);
nor U29743 (N_29743,N_29460,N_29377);
xor U29744 (N_29744,N_29348,N_29256);
nand U29745 (N_29745,N_29408,N_29432);
xnor U29746 (N_29746,N_29274,N_29268);
and U29747 (N_29747,N_29472,N_29306);
nand U29748 (N_29748,N_29426,N_29275);
or U29749 (N_29749,N_29380,N_29303);
xor U29750 (N_29750,N_29674,N_29727);
or U29751 (N_29751,N_29581,N_29715);
nand U29752 (N_29752,N_29708,N_29563);
or U29753 (N_29753,N_29723,N_29559);
xnor U29754 (N_29754,N_29749,N_29724);
or U29755 (N_29755,N_29738,N_29714);
xnor U29756 (N_29756,N_29619,N_29536);
nand U29757 (N_29757,N_29602,N_29571);
nand U29758 (N_29758,N_29503,N_29670);
or U29759 (N_29759,N_29606,N_29548);
nand U29760 (N_29760,N_29580,N_29520);
and U29761 (N_29761,N_29565,N_29644);
nand U29762 (N_29762,N_29583,N_29586);
nor U29763 (N_29763,N_29707,N_29717);
xnor U29764 (N_29764,N_29542,N_29656);
nor U29765 (N_29765,N_29729,N_29607);
or U29766 (N_29766,N_29667,N_29735);
nand U29767 (N_29767,N_29524,N_29595);
or U29768 (N_29768,N_29693,N_29544);
or U29769 (N_29769,N_29614,N_29545);
nor U29770 (N_29770,N_29584,N_29731);
xnor U29771 (N_29771,N_29637,N_29515);
nor U29772 (N_29772,N_29541,N_29730);
xnor U29773 (N_29773,N_29574,N_29537);
or U29774 (N_29774,N_29554,N_29745);
xnor U29775 (N_29775,N_29593,N_29538);
xnor U29776 (N_29776,N_29550,N_29576);
xor U29777 (N_29777,N_29500,N_29628);
nand U29778 (N_29778,N_29528,N_29603);
and U29779 (N_29779,N_29646,N_29533);
nand U29780 (N_29780,N_29675,N_29560);
nand U29781 (N_29781,N_29666,N_29720);
nand U29782 (N_29782,N_29673,N_29645);
xor U29783 (N_29783,N_29668,N_29592);
nor U29784 (N_29784,N_29712,N_29655);
or U29785 (N_29785,N_29549,N_29722);
and U29786 (N_29786,N_29513,N_29744);
nor U29787 (N_29787,N_29691,N_29716);
nor U29788 (N_29788,N_29532,N_29654);
xor U29789 (N_29789,N_29652,N_29534);
and U29790 (N_29790,N_29709,N_29695);
xor U29791 (N_29791,N_29599,N_29570);
nor U29792 (N_29792,N_29627,N_29507);
and U29793 (N_29793,N_29590,N_29526);
nand U29794 (N_29794,N_29687,N_29521);
and U29795 (N_29795,N_29684,N_29509);
nand U29796 (N_29796,N_29636,N_29582);
nand U29797 (N_29797,N_29683,N_29685);
or U29798 (N_29798,N_29643,N_29501);
nor U29799 (N_29799,N_29622,N_29615);
nand U29800 (N_29800,N_29625,N_29621);
and U29801 (N_29801,N_29694,N_29594);
or U29802 (N_29802,N_29530,N_29710);
or U29803 (N_29803,N_29728,N_29539);
and U29804 (N_29804,N_29510,N_29657);
and U29805 (N_29805,N_29523,N_29742);
nand U29806 (N_29806,N_29679,N_29671);
and U29807 (N_29807,N_29608,N_29697);
xnor U29808 (N_29808,N_29589,N_29527);
or U29809 (N_29809,N_29650,N_29686);
nor U29810 (N_29810,N_29511,N_29663);
and U29811 (N_29811,N_29651,N_29613);
nor U29812 (N_29812,N_29601,N_29699);
or U29813 (N_29813,N_29649,N_29564);
or U29814 (N_29814,N_29692,N_29543);
and U29815 (N_29815,N_29746,N_29566);
and U29816 (N_29816,N_29680,N_29702);
nor U29817 (N_29817,N_29626,N_29688);
xor U29818 (N_29818,N_29741,N_29502);
nor U29819 (N_29819,N_29557,N_29640);
nand U29820 (N_29820,N_29732,N_29681);
nand U29821 (N_29821,N_29623,N_29653);
nand U29822 (N_29822,N_29672,N_29711);
xor U29823 (N_29823,N_29642,N_29600);
xnor U29824 (N_29824,N_29618,N_29561);
nor U29825 (N_29825,N_29633,N_29573);
nor U29826 (N_29826,N_29555,N_29629);
nor U29827 (N_29827,N_29518,N_29661);
xnor U29828 (N_29828,N_29531,N_29588);
or U29829 (N_29829,N_29529,N_29556);
and U29830 (N_29830,N_29591,N_29577);
xor U29831 (N_29831,N_29682,N_29700);
nor U29832 (N_29832,N_29706,N_29748);
nor U29833 (N_29833,N_29665,N_29669);
and U29834 (N_29834,N_29739,N_29734);
nor U29835 (N_29835,N_29719,N_29690);
nand U29836 (N_29836,N_29662,N_29547);
xnor U29837 (N_29837,N_29726,N_29689);
nor U29838 (N_29838,N_29553,N_29517);
nand U29839 (N_29839,N_29508,N_29659);
nand U29840 (N_29840,N_29630,N_29609);
and U29841 (N_29841,N_29535,N_29612);
and U29842 (N_29842,N_29512,N_29567);
or U29843 (N_29843,N_29616,N_29743);
or U29844 (N_29844,N_29620,N_29604);
xnor U29845 (N_29845,N_29648,N_29579);
xor U29846 (N_29846,N_29525,N_29516);
nand U29847 (N_29847,N_29505,N_29737);
nor U29848 (N_29848,N_29558,N_29552);
nand U29849 (N_29849,N_29562,N_29721);
xnor U29850 (N_29850,N_29631,N_29660);
nand U29851 (N_29851,N_29736,N_29747);
nor U29852 (N_29852,N_29634,N_29598);
or U29853 (N_29853,N_29597,N_29572);
or U29854 (N_29854,N_29635,N_29522);
nand U29855 (N_29855,N_29568,N_29664);
or U29856 (N_29856,N_29677,N_29596);
and U29857 (N_29857,N_29725,N_29733);
or U29858 (N_29858,N_29504,N_29569);
nor U29859 (N_29859,N_29703,N_29696);
nand U29860 (N_29860,N_29639,N_29551);
nand U29861 (N_29861,N_29641,N_29701);
nor U29862 (N_29862,N_29638,N_29540);
and U29863 (N_29863,N_29632,N_29617);
and U29864 (N_29864,N_29519,N_29506);
nand U29865 (N_29865,N_29698,N_29587);
nor U29866 (N_29866,N_29575,N_29713);
and U29867 (N_29867,N_29740,N_29704);
or U29868 (N_29868,N_29610,N_29676);
nor U29869 (N_29869,N_29705,N_29658);
xnor U29870 (N_29870,N_29718,N_29585);
or U29871 (N_29871,N_29678,N_29647);
or U29872 (N_29872,N_29546,N_29611);
or U29873 (N_29873,N_29605,N_29514);
and U29874 (N_29874,N_29578,N_29624);
xnor U29875 (N_29875,N_29597,N_29728);
nor U29876 (N_29876,N_29621,N_29749);
nor U29877 (N_29877,N_29610,N_29656);
nand U29878 (N_29878,N_29506,N_29593);
nand U29879 (N_29879,N_29556,N_29590);
or U29880 (N_29880,N_29540,N_29534);
or U29881 (N_29881,N_29569,N_29645);
xor U29882 (N_29882,N_29544,N_29669);
nand U29883 (N_29883,N_29591,N_29558);
xnor U29884 (N_29884,N_29571,N_29735);
or U29885 (N_29885,N_29667,N_29654);
xnor U29886 (N_29886,N_29557,N_29568);
nand U29887 (N_29887,N_29537,N_29653);
nor U29888 (N_29888,N_29605,N_29675);
nor U29889 (N_29889,N_29748,N_29699);
or U29890 (N_29890,N_29586,N_29522);
xnor U29891 (N_29891,N_29599,N_29587);
nor U29892 (N_29892,N_29562,N_29520);
nor U29893 (N_29893,N_29588,N_29711);
or U29894 (N_29894,N_29574,N_29520);
nor U29895 (N_29895,N_29620,N_29635);
nor U29896 (N_29896,N_29715,N_29740);
xnor U29897 (N_29897,N_29743,N_29681);
nand U29898 (N_29898,N_29731,N_29612);
nand U29899 (N_29899,N_29599,N_29609);
or U29900 (N_29900,N_29582,N_29562);
and U29901 (N_29901,N_29640,N_29694);
or U29902 (N_29902,N_29628,N_29656);
or U29903 (N_29903,N_29509,N_29501);
or U29904 (N_29904,N_29586,N_29680);
or U29905 (N_29905,N_29526,N_29534);
and U29906 (N_29906,N_29638,N_29668);
nand U29907 (N_29907,N_29575,N_29539);
and U29908 (N_29908,N_29601,N_29506);
xor U29909 (N_29909,N_29662,N_29611);
or U29910 (N_29910,N_29602,N_29621);
nor U29911 (N_29911,N_29665,N_29505);
or U29912 (N_29912,N_29717,N_29637);
nand U29913 (N_29913,N_29572,N_29674);
nor U29914 (N_29914,N_29577,N_29641);
nand U29915 (N_29915,N_29613,N_29530);
nor U29916 (N_29916,N_29562,N_29587);
or U29917 (N_29917,N_29538,N_29596);
nor U29918 (N_29918,N_29530,N_29672);
or U29919 (N_29919,N_29645,N_29743);
xnor U29920 (N_29920,N_29743,N_29731);
nor U29921 (N_29921,N_29530,N_29508);
or U29922 (N_29922,N_29700,N_29501);
nand U29923 (N_29923,N_29651,N_29545);
nand U29924 (N_29924,N_29717,N_29691);
and U29925 (N_29925,N_29698,N_29669);
or U29926 (N_29926,N_29639,N_29719);
and U29927 (N_29927,N_29573,N_29638);
or U29928 (N_29928,N_29669,N_29657);
nor U29929 (N_29929,N_29539,N_29503);
and U29930 (N_29930,N_29688,N_29693);
nand U29931 (N_29931,N_29679,N_29711);
nand U29932 (N_29932,N_29599,N_29680);
or U29933 (N_29933,N_29642,N_29584);
and U29934 (N_29934,N_29658,N_29536);
nand U29935 (N_29935,N_29595,N_29708);
and U29936 (N_29936,N_29557,N_29536);
nor U29937 (N_29937,N_29658,N_29635);
and U29938 (N_29938,N_29582,N_29591);
and U29939 (N_29939,N_29617,N_29593);
nor U29940 (N_29940,N_29533,N_29628);
and U29941 (N_29941,N_29649,N_29586);
nor U29942 (N_29942,N_29602,N_29532);
or U29943 (N_29943,N_29590,N_29743);
nand U29944 (N_29944,N_29644,N_29571);
nand U29945 (N_29945,N_29575,N_29646);
nor U29946 (N_29946,N_29627,N_29730);
or U29947 (N_29947,N_29711,N_29736);
xnor U29948 (N_29948,N_29533,N_29521);
or U29949 (N_29949,N_29548,N_29649);
xor U29950 (N_29950,N_29734,N_29511);
xnor U29951 (N_29951,N_29664,N_29714);
and U29952 (N_29952,N_29676,N_29717);
or U29953 (N_29953,N_29691,N_29654);
nor U29954 (N_29954,N_29588,N_29538);
nor U29955 (N_29955,N_29504,N_29513);
or U29956 (N_29956,N_29621,N_29675);
nand U29957 (N_29957,N_29564,N_29735);
xor U29958 (N_29958,N_29693,N_29523);
nor U29959 (N_29959,N_29607,N_29662);
nor U29960 (N_29960,N_29549,N_29632);
nand U29961 (N_29961,N_29674,N_29577);
nand U29962 (N_29962,N_29623,N_29549);
and U29963 (N_29963,N_29748,N_29722);
nand U29964 (N_29964,N_29645,N_29572);
nor U29965 (N_29965,N_29540,N_29705);
nand U29966 (N_29966,N_29699,N_29735);
nand U29967 (N_29967,N_29671,N_29563);
nand U29968 (N_29968,N_29509,N_29743);
nor U29969 (N_29969,N_29535,N_29587);
nand U29970 (N_29970,N_29543,N_29578);
nand U29971 (N_29971,N_29530,N_29654);
or U29972 (N_29972,N_29694,N_29615);
xnor U29973 (N_29973,N_29629,N_29744);
or U29974 (N_29974,N_29629,N_29626);
or U29975 (N_29975,N_29512,N_29585);
or U29976 (N_29976,N_29534,N_29690);
nor U29977 (N_29977,N_29706,N_29670);
xnor U29978 (N_29978,N_29519,N_29662);
or U29979 (N_29979,N_29712,N_29720);
and U29980 (N_29980,N_29608,N_29509);
nand U29981 (N_29981,N_29604,N_29557);
and U29982 (N_29982,N_29739,N_29666);
or U29983 (N_29983,N_29658,N_29733);
nor U29984 (N_29984,N_29657,N_29539);
nand U29985 (N_29985,N_29622,N_29609);
xor U29986 (N_29986,N_29526,N_29561);
or U29987 (N_29987,N_29539,N_29644);
nand U29988 (N_29988,N_29716,N_29506);
and U29989 (N_29989,N_29740,N_29723);
nor U29990 (N_29990,N_29702,N_29735);
nand U29991 (N_29991,N_29595,N_29629);
or U29992 (N_29992,N_29627,N_29563);
xnor U29993 (N_29993,N_29736,N_29619);
and U29994 (N_29994,N_29530,N_29635);
and U29995 (N_29995,N_29715,N_29593);
nor U29996 (N_29996,N_29655,N_29748);
and U29997 (N_29997,N_29653,N_29611);
nor U29998 (N_29998,N_29612,N_29554);
nor U29999 (N_29999,N_29651,N_29729);
nor U30000 (N_30000,N_29922,N_29985);
xnor U30001 (N_30001,N_29822,N_29969);
nor U30002 (N_30002,N_29841,N_29973);
and U30003 (N_30003,N_29881,N_29975);
or U30004 (N_30004,N_29809,N_29825);
nand U30005 (N_30005,N_29959,N_29757);
nand U30006 (N_30006,N_29955,N_29824);
xnor U30007 (N_30007,N_29924,N_29782);
xor U30008 (N_30008,N_29788,N_29868);
nor U30009 (N_30009,N_29886,N_29986);
nor U30010 (N_30010,N_29902,N_29870);
or U30011 (N_30011,N_29843,N_29981);
xor U30012 (N_30012,N_29828,N_29764);
and U30013 (N_30013,N_29941,N_29767);
xor U30014 (N_30014,N_29854,N_29778);
nand U30015 (N_30015,N_29765,N_29996);
and U30016 (N_30016,N_29775,N_29948);
or U30017 (N_30017,N_29808,N_29939);
nand U30018 (N_30018,N_29839,N_29999);
or U30019 (N_30019,N_29880,N_29889);
nor U30020 (N_30020,N_29997,N_29750);
xnor U30021 (N_30021,N_29813,N_29908);
nor U30022 (N_30022,N_29925,N_29872);
or U30023 (N_30023,N_29848,N_29810);
nor U30024 (N_30024,N_29761,N_29840);
nor U30025 (N_30025,N_29927,N_29912);
xor U30026 (N_30026,N_29799,N_29937);
nor U30027 (N_30027,N_29784,N_29879);
nor U30028 (N_30028,N_29857,N_29911);
xnor U30029 (N_30029,N_29883,N_29835);
nand U30030 (N_30030,N_29935,N_29771);
nor U30031 (N_30031,N_29890,N_29792);
nand U30032 (N_30032,N_29984,N_29979);
and U30033 (N_30033,N_29861,N_29753);
nand U30034 (N_30034,N_29844,N_29992);
xor U30035 (N_30035,N_29966,N_29960);
nand U30036 (N_30036,N_29919,N_29884);
and U30037 (N_30037,N_29779,N_29863);
and U30038 (N_30038,N_29790,N_29789);
and U30039 (N_30039,N_29817,N_29993);
and U30040 (N_30040,N_29899,N_29953);
or U30041 (N_30041,N_29807,N_29932);
or U30042 (N_30042,N_29982,N_29988);
or U30043 (N_30043,N_29787,N_29791);
nand U30044 (N_30044,N_29850,N_29907);
or U30045 (N_30045,N_29929,N_29990);
and U30046 (N_30046,N_29849,N_29759);
nand U30047 (N_30047,N_29842,N_29876);
nand U30048 (N_30048,N_29887,N_29766);
or U30049 (N_30049,N_29751,N_29957);
or U30050 (N_30050,N_29991,N_29987);
or U30051 (N_30051,N_29962,N_29958);
xnor U30052 (N_30052,N_29972,N_29760);
and U30053 (N_30053,N_29977,N_29914);
or U30054 (N_30054,N_29819,N_29818);
nor U30055 (N_30055,N_29794,N_29917);
or U30056 (N_30056,N_29888,N_29777);
or U30057 (N_30057,N_29947,N_29971);
nand U30058 (N_30058,N_29785,N_29938);
nand U30059 (N_30059,N_29893,N_29823);
nand U30060 (N_30060,N_29877,N_29847);
or U30061 (N_30061,N_29949,N_29903);
or U30062 (N_30062,N_29866,N_29995);
or U30063 (N_30063,N_29834,N_29803);
nor U30064 (N_30064,N_29943,N_29853);
xnor U30065 (N_30065,N_29860,N_29951);
nand U30066 (N_30066,N_29798,N_29852);
and U30067 (N_30067,N_29950,N_29826);
nand U30068 (N_30068,N_29768,N_29773);
nor U30069 (N_30069,N_29815,N_29797);
xnor U30070 (N_30070,N_29913,N_29867);
nand U30071 (N_30071,N_29900,N_29805);
and U30072 (N_30072,N_29837,N_29871);
nand U30073 (N_30073,N_29930,N_29897);
nor U30074 (N_30074,N_29994,N_29864);
or U30075 (N_30075,N_29931,N_29856);
nor U30076 (N_30076,N_29940,N_29758);
or U30077 (N_30077,N_29967,N_29901);
nand U30078 (N_30078,N_29942,N_29769);
nand U30079 (N_30079,N_29795,N_29980);
or U30080 (N_30080,N_29933,N_29801);
or U30081 (N_30081,N_29974,N_29921);
nand U30082 (N_30082,N_29793,N_29838);
and U30083 (N_30083,N_29821,N_29816);
or U30084 (N_30084,N_29936,N_29800);
nor U30085 (N_30085,N_29865,N_29875);
and U30086 (N_30086,N_29970,N_29820);
and U30087 (N_30087,N_29963,N_29783);
xnor U30088 (N_30088,N_29926,N_29954);
nand U30089 (N_30089,N_29952,N_29906);
nor U30090 (N_30090,N_29796,N_29873);
xor U30091 (N_30091,N_29812,N_29916);
nand U30092 (N_30092,N_29989,N_29878);
nor U30093 (N_30093,N_29920,N_29858);
nor U30094 (N_30094,N_29832,N_29776);
nand U30095 (N_30095,N_29998,N_29786);
xor U30096 (N_30096,N_29811,N_29829);
nor U30097 (N_30097,N_29923,N_29869);
and U30098 (N_30098,N_29806,N_29885);
or U30099 (N_30099,N_29763,N_29896);
xor U30100 (N_30100,N_29814,N_29928);
or U30101 (N_30101,N_29946,N_29874);
or U30102 (N_30102,N_29895,N_29827);
nor U30103 (N_30103,N_29862,N_29846);
and U30104 (N_30104,N_29905,N_29915);
xnor U30105 (N_30105,N_29892,N_29904);
and U30106 (N_30106,N_29891,N_29918);
xnor U30107 (N_30107,N_29762,N_29934);
and U30108 (N_30108,N_29894,N_29976);
xor U30109 (N_30109,N_29978,N_29802);
xor U30110 (N_30110,N_29836,N_29833);
xnor U30111 (N_30111,N_29831,N_29830);
nor U30112 (N_30112,N_29983,N_29968);
or U30113 (N_30113,N_29752,N_29956);
and U30114 (N_30114,N_29772,N_29855);
or U30115 (N_30115,N_29859,N_29910);
or U30116 (N_30116,N_29804,N_29961);
nor U30117 (N_30117,N_29964,N_29781);
nand U30118 (N_30118,N_29845,N_29754);
and U30119 (N_30119,N_29756,N_29965);
and U30120 (N_30120,N_29780,N_29851);
nand U30121 (N_30121,N_29944,N_29945);
and U30122 (N_30122,N_29755,N_29882);
and U30123 (N_30123,N_29770,N_29898);
or U30124 (N_30124,N_29774,N_29909);
or U30125 (N_30125,N_29799,N_29956);
xnor U30126 (N_30126,N_29913,N_29860);
xnor U30127 (N_30127,N_29811,N_29975);
nor U30128 (N_30128,N_29784,N_29822);
or U30129 (N_30129,N_29793,N_29876);
nor U30130 (N_30130,N_29910,N_29863);
nand U30131 (N_30131,N_29788,N_29991);
nor U30132 (N_30132,N_29931,N_29997);
and U30133 (N_30133,N_29822,N_29773);
nand U30134 (N_30134,N_29920,N_29991);
and U30135 (N_30135,N_29867,N_29904);
nand U30136 (N_30136,N_29822,N_29849);
or U30137 (N_30137,N_29773,N_29911);
or U30138 (N_30138,N_29806,N_29888);
and U30139 (N_30139,N_29780,N_29862);
and U30140 (N_30140,N_29840,N_29767);
nor U30141 (N_30141,N_29781,N_29890);
xor U30142 (N_30142,N_29980,N_29859);
nor U30143 (N_30143,N_29839,N_29931);
or U30144 (N_30144,N_29752,N_29985);
or U30145 (N_30145,N_29768,N_29916);
or U30146 (N_30146,N_29788,N_29770);
nor U30147 (N_30147,N_29771,N_29869);
nor U30148 (N_30148,N_29979,N_29826);
or U30149 (N_30149,N_29913,N_29759);
or U30150 (N_30150,N_29788,N_29829);
nand U30151 (N_30151,N_29854,N_29870);
or U30152 (N_30152,N_29870,N_29890);
xor U30153 (N_30153,N_29832,N_29977);
nor U30154 (N_30154,N_29990,N_29923);
or U30155 (N_30155,N_29775,N_29930);
xnor U30156 (N_30156,N_29994,N_29761);
nand U30157 (N_30157,N_29892,N_29850);
and U30158 (N_30158,N_29927,N_29972);
or U30159 (N_30159,N_29990,N_29799);
nand U30160 (N_30160,N_29814,N_29917);
nor U30161 (N_30161,N_29758,N_29775);
and U30162 (N_30162,N_29970,N_29965);
xor U30163 (N_30163,N_29994,N_29960);
and U30164 (N_30164,N_29995,N_29884);
and U30165 (N_30165,N_29758,N_29961);
and U30166 (N_30166,N_29925,N_29842);
nor U30167 (N_30167,N_29901,N_29979);
xnor U30168 (N_30168,N_29920,N_29879);
nor U30169 (N_30169,N_29866,N_29824);
nor U30170 (N_30170,N_29878,N_29798);
and U30171 (N_30171,N_29932,N_29929);
xor U30172 (N_30172,N_29819,N_29947);
nand U30173 (N_30173,N_29815,N_29831);
and U30174 (N_30174,N_29931,N_29951);
nand U30175 (N_30175,N_29896,N_29826);
or U30176 (N_30176,N_29838,N_29794);
nand U30177 (N_30177,N_29909,N_29761);
and U30178 (N_30178,N_29822,N_29909);
or U30179 (N_30179,N_29875,N_29935);
or U30180 (N_30180,N_29768,N_29831);
nand U30181 (N_30181,N_29854,N_29904);
nor U30182 (N_30182,N_29786,N_29801);
nand U30183 (N_30183,N_29940,N_29952);
and U30184 (N_30184,N_29783,N_29946);
xnor U30185 (N_30185,N_29988,N_29987);
nor U30186 (N_30186,N_29873,N_29928);
and U30187 (N_30187,N_29860,N_29831);
and U30188 (N_30188,N_29961,N_29981);
nor U30189 (N_30189,N_29984,N_29858);
nand U30190 (N_30190,N_29933,N_29985);
nor U30191 (N_30191,N_29796,N_29957);
xnor U30192 (N_30192,N_29894,N_29783);
and U30193 (N_30193,N_29965,N_29771);
nor U30194 (N_30194,N_29776,N_29897);
nand U30195 (N_30195,N_29999,N_29836);
xnor U30196 (N_30196,N_29998,N_29857);
or U30197 (N_30197,N_29869,N_29912);
xor U30198 (N_30198,N_29919,N_29983);
and U30199 (N_30199,N_29874,N_29837);
or U30200 (N_30200,N_29986,N_29979);
xnor U30201 (N_30201,N_29879,N_29955);
nand U30202 (N_30202,N_29845,N_29930);
nand U30203 (N_30203,N_29752,N_29902);
nand U30204 (N_30204,N_29761,N_29866);
xnor U30205 (N_30205,N_29760,N_29982);
and U30206 (N_30206,N_29827,N_29926);
nor U30207 (N_30207,N_29887,N_29883);
xor U30208 (N_30208,N_29778,N_29876);
and U30209 (N_30209,N_29781,N_29916);
or U30210 (N_30210,N_29862,N_29901);
nand U30211 (N_30211,N_29793,N_29823);
nand U30212 (N_30212,N_29858,N_29886);
xor U30213 (N_30213,N_29907,N_29795);
or U30214 (N_30214,N_29755,N_29875);
and U30215 (N_30215,N_29963,N_29789);
nand U30216 (N_30216,N_29875,N_29806);
or U30217 (N_30217,N_29908,N_29998);
nor U30218 (N_30218,N_29906,N_29953);
nand U30219 (N_30219,N_29970,N_29994);
nor U30220 (N_30220,N_29848,N_29995);
nor U30221 (N_30221,N_29824,N_29932);
and U30222 (N_30222,N_29973,N_29916);
or U30223 (N_30223,N_29983,N_29878);
nand U30224 (N_30224,N_29803,N_29876);
or U30225 (N_30225,N_29875,N_29857);
and U30226 (N_30226,N_29822,N_29858);
or U30227 (N_30227,N_29771,N_29801);
nand U30228 (N_30228,N_29938,N_29936);
nand U30229 (N_30229,N_29894,N_29960);
or U30230 (N_30230,N_29873,N_29926);
and U30231 (N_30231,N_29962,N_29816);
nand U30232 (N_30232,N_29812,N_29965);
nor U30233 (N_30233,N_29866,N_29832);
and U30234 (N_30234,N_29794,N_29894);
nand U30235 (N_30235,N_29837,N_29886);
and U30236 (N_30236,N_29862,N_29784);
xnor U30237 (N_30237,N_29906,N_29909);
nand U30238 (N_30238,N_29990,N_29994);
nand U30239 (N_30239,N_29888,N_29982);
nor U30240 (N_30240,N_29944,N_29897);
xnor U30241 (N_30241,N_29887,N_29908);
nand U30242 (N_30242,N_29915,N_29954);
xor U30243 (N_30243,N_29993,N_29806);
and U30244 (N_30244,N_29956,N_29866);
xnor U30245 (N_30245,N_29864,N_29820);
nor U30246 (N_30246,N_29948,N_29941);
xnor U30247 (N_30247,N_29856,N_29799);
or U30248 (N_30248,N_29781,N_29841);
or U30249 (N_30249,N_29814,N_29875);
and U30250 (N_30250,N_30105,N_30177);
nor U30251 (N_30251,N_30079,N_30071);
or U30252 (N_30252,N_30035,N_30112);
nor U30253 (N_30253,N_30024,N_30104);
or U30254 (N_30254,N_30229,N_30041);
and U30255 (N_30255,N_30189,N_30069);
and U30256 (N_30256,N_30190,N_30039);
or U30257 (N_30257,N_30057,N_30012);
and U30258 (N_30258,N_30116,N_30222);
nor U30259 (N_30259,N_30201,N_30078);
nand U30260 (N_30260,N_30203,N_30233);
or U30261 (N_30261,N_30195,N_30234);
and U30262 (N_30262,N_30074,N_30220);
nor U30263 (N_30263,N_30036,N_30236);
nor U30264 (N_30264,N_30058,N_30180);
nor U30265 (N_30265,N_30099,N_30033);
or U30266 (N_30266,N_30188,N_30152);
or U30267 (N_30267,N_30157,N_30130);
nand U30268 (N_30268,N_30174,N_30055);
or U30269 (N_30269,N_30169,N_30230);
nor U30270 (N_30270,N_30240,N_30001);
nor U30271 (N_30271,N_30209,N_30198);
and U30272 (N_30272,N_30048,N_30026);
xnor U30273 (N_30273,N_30192,N_30211);
nand U30274 (N_30274,N_30046,N_30158);
nand U30275 (N_30275,N_30061,N_30227);
and U30276 (N_30276,N_30051,N_30159);
nand U30277 (N_30277,N_30129,N_30197);
or U30278 (N_30278,N_30175,N_30148);
or U30279 (N_30279,N_30094,N_30010);
and U30280 (N_30280,N_30005,N_30137);
nor U30281 (N_30281,N_30021,N_30185);
xor U30282 (N_30282,N_30030,N_30049);
nor U30283 (N_30283,N_30059,N_30204);
nor U30284 (N_30284,N_30173,N_30194);
or U30285 (N_30285,N_30066,N_30006);
nor U30286 (N_30286,N_30085,N_30163);
or U30287 (N_30287,N_30047,N_30062);
xnor U30288 (N_30288,N_30064,N_30031);
xnor U30289 (N_30289,N_30165,N_30239);
and U30290 (N_30290,N_30052,N_30170);
nor U30291 (N_30291,N_30214,N_30206);
nor U30292 (N_30292,N_30120,N_30145);
or U30293 (N_30293,N_30007,N_30097);
nor U30294 (N_30294,N_30076,N_30123);
xor U30295 (N_30295,N_30118,N_30176);
and U30296 (N_30296,N_30122,N_30155);
nor U30297 (N_30297,N_30045,N_30022);
xor U30298 (N_30298,N_30161,N_30065);
or U30299 (N_30299,N_30060,N_30136);
xor U30300 (N_30300,N_30027,N_30088);
xor U30301 (N_30301,N_30138,N_30092);
nor U30302 (N_30302,N_30207,N_30077);
xnor U30303 (N_30303,N_30011,N_30224);
xor U30304 (N_30304,N_30090,N_30015);
and U30305 (N_30305,N_30156,N_30098);
or U30306 (N_30306,N_30042,N_30100);
xnor U30307 (N_30307,N_30108,N_30162);
or U30308 (N_30308,N_30187,N_30023);
and U30309 (N_30309,N_30226,N_30243);
and U30310 (N_30310,N_30232,N_30133);
and U30311 (N_30311,N_30082,N_30218);
nand U30312 (N_30312,N_30181,N_30053);
and U30313 (N_30313,N_30183,N_30068);
and U30314 (N_30314,N_30111,N_30154);
or U30315 (N_30315,N_30200,N_30142);
xnor U30316 (N_30316,N_30109,N_30083);
or U30317 (N_30317,N_30225,N_30017);
or U30318 (N_30318,N_30144,N_30020);
nor U30319 (N_30319,N_30228,N_30089);
xnor U30320 (N_30320,N_30184,N_30249);
xor U30321 (N_30321,N_30205,N_30168);
and U30322 (N_30322,N_30219,N_30140);
xnor U30323 (N_30323,N_30160,N_30131);
and U30324 (N_30324,N_30210,N_30182);
and U30325 (N_30325,N_30241,N_30101);
xor U30326 (N_30326,N_30172,N_30106);
nand U30327 (N_30327,N_30143,N_30223);
nor U30328 (N_30328,N_30217,N_30215);
xor U30329 (N_30329,N_30019,N_30171);
nor U30330 (N_30330,N_30246,N_30032);
and U30331 (N_30331,N_30086,N_30153);
xor U30332 (N_30332,N_30000,N_30221);
and U30333 (N_30333,N_30102,N_30093);
xor U30334 (N_30334,N_30009,N_30212);
xor U30335 (N_30335,N_30084,N_30095);
xor U30336 (N_30336,N_30238,N_30124);
nand U30337 (N_30337,N_30166,N_30110);
xnor U30338 (N_30338,N_30151,N_30167);
and U30339 (N_30339,N_30147,N_30008);
and U30340 (N_30340,N_30128,N_30040);
or U30341 (N_30341,N_30034,N_30127);
nand U30342 (N_30342,N_30072,N_30056);
or U30343 (N_30343,N_30121,N_30038);
xor U30344 (N_30344,N_30146,N_30016);
and U30345 (N_30345,N_30196,N_30063);
nand U30346 (N_30346,N_30050,N_30018);
and U30347 (N_30347,N_30029,N_30025);
nand U30348 (N_30348,N_30004,N_30141);
or U30349 (N_30349,N_30037,N_30213);
or U30350 (N_30350,N_30149,N_30087);
or U30351 (N_30351,N_30135,N_30113);
nand U30352 (N_30352,N_30091,N_30075);
xnor U30353 (N_30353,N_30216,N_30028);
xor U30354 (N_30354,N_30242,N_30134);
nor U30355 (N_30355,N_30235,N_30244);
nor U30356 (N_30356,N_30179,N_30139);
nor U30357 (N_30357,N_30044,N_30070);
and U30358 (N_30358,N_30043,N_30115);
nor U30359 (N_30359,N_30248,N_30126);
xor U30360 (N_30360,N_30081,N_30013);
nor U30361 (N_30361,N_30103,N_30150);
or U30362 (N_30362,N_30107,N_30117);
xor U30363 (N_30363,N_30202,N_30247);
nand U30364 (N_30364,N_30054,N_30014);
xor U30365 (N_30365,N_30114,N_30002);
nand U30366 (N_30366,N_30073,N_30191);
nor U30367 (N_30367,N_30164,N_30186);
nor U30368 (N_30368,N_30231,N_30193);
or U30369 (N_30369,N_30080,N_30132);
and U30370 (N_30370,N_30245,N_30067);
nor U30371 (N_30371,N_30199,N_30208);
and U30372 (N_30372,N_30119,N_30178);
or U30373 (N_30373,N_30003,N_30237);
and U30374 (N_30374,N_30125,N_30096);
or U30375 (N_30375,N_30241,N_30136);
or U30376 (N_30376,N_30023,N_30177);
nand U30377 (N_30377,N_30076,N_30129);
and U30378 (N_30378,N_30034,N_30021);
xnor U30379 (N_30379,N_30014,N_30026);
nor U30380 (N_30380,N_30026,N_30032);
nor U30381 (N_30381,N_30193,N_30174);
nor U30382 (N_30382,N_30190,N_30003);
and U30383 (N_30383,N_30108,N_30093);
nand U30384 (N_30384,N_30194,N_30183);
nand U30385 (N_30385,N_30242,N_30199);
xor U30386 (N_30386,N_30198,N_30116);
nand U30387 (N_30387,N_30218,N_30118);
xor U30388 (N_30388,N_30145,N_30212);
and U30389 (N_30389,N_30146,N_30124);
xnor U30390 (N_30390,N_30044,N_30095);
xnor U30391 (N_30391,N_30167,N_30249);
and U30392 (N_30392,N_30204,N_30249);
xor U30393 (N_30393,N_30109,N_30031);
or U30394 (N_30394,N_30029,N_30189);
xor U30395 (N_30395,N_30234,N_30085);
or U30396 (N_30396,N_30053,N_30054);
or U30397 (N_30397,N_30149,N_30160);
and U30398 (N_30398,N_30162,N_30149);
xnor U30399 (N_30399,N_30032,N_30212);
nand U30400 (N_30400,N_30131,N_30141);
and U30401 (N_30401,N_30047,N_30006);
nand U30402 (N_30402,N_30022,N_30064);
or U30403 (N_30403,N_30118,N_30057);
nand U30404 (N_30404,N_30128,N_30163);
nor U30405 (N_30405,N_30161,N_30028);
or U30406 (N_30406,N_30045,N_30113);
nor U30407 (N_30407,N_30054,N_30122);
or U30408 (N_30408,N_30042,N_30182);
and U30409 (N_30409,N_30230,N_30165);
nor U30410 (N_30410,N_30112,N_30029);
or U30411 (N_30411,N_30145,N_30049);
and U30412 (N_30412,N_30107,N_30220);
nor U30413 (N_30413,N_30155,N_30003);
or U30414 (N_30414,N_30087,N_30035);
nor U30415 (N_30415,N_30188,N_30083);
xnor U30416 (N_30416,N_30161,N_30001);
and U30417 (N_30417,N_30207,N_30048);
and U30418 (N_30418,N_30244,N_30162);
and U30419 (N_30419,N_30109,N_30074);
nand U30420 (N_30420,N_30009,N_30144);
or U30421 (N_30421,N_30073,N_30169);
or U30422 (N_30422,N_30226,N_30060);
and U30423 (N_30423,N_30159,N_30147);
nand U30424 (N_30424,N_30063,N_30203);
and U30425 (N_30425,N_30123,N_30053);
nand U30426 (N_30426,N_30020,N_30148);
nor U30427 (N_30427,N_30210,N_30138);
nand U30428 (N_30428,N_30101,N_30023);
or U30429 (N_30429,N_30216,N_30233);
or U30430 (N_30430,N_30245,N_30221);
or U30431 (N_30431,N_30141,N_30088);
nand U30432 (N_30432,N_30088,N_30136);
nand U30433 (N_30433,N_30216,N_30224);
nand U30434 (N_30434,N_30049,N_30067);
nand U30435 (N_30435,N_30178,N_30235);
nand U30436 (N_30436,N_30080,N_30026);
nand U30437 (N_30437,N_30149,N_30161);
nand U30438 (N_30438,N_30231,N_30109);
xor U30439 (N_30439,N_30144,N_30129);
nor U30440 (N_30440,N_30194,N_30072);
nand U30441 (N_30441,N_30203,N_30152);
nand U30442 (N_30442,N_30234,N_30163);
nand U30443 (N_30443,N_30085,N_30214);
or U30444 (N_30444,N_30008,N_30192);
nand U30445 (N_30445,N_30204,N_30085);
or U30446 (N_30446,N_30216,N_30132);
xor U30447 (N_30447,N_30081,N_30244);
nand U30448 (N_30448,N_30107,N_30097);
nor U30449 (N_30449,N_30233,N_30021);
xor U30450 (N_30450,N_30043,N_30214);
nand U30451 (N_30451,N_30004,N_30075);
and U30452 (N_30452,N_30106,N_30156);
and U30453 (N_30453,N_30027,N_30092);
xor U30454 (N_30454,N_30224,N_30117);
and U30455 (N_30455,N_30082,N_30063);
nand U30456 (N_30456,N_30183,N_30022);
nand U30457 (N_30457,N_30000,N_30108);
nand U30458 (N_30458,N_30156,N_30005);
nor U30459 (N_30459,N_30109,N_30065);
xnor U30460 (N_30460,N_30007,N_30238);
nor U30461 (N_30461,N_30209,N_30093);
nor U30462 (N_30462,N_30202,N_30230);
nand U30463 (N_30463,N_30177,N_30065);
nand U30464 (N_30464,N_30169,N_30022);
nand U30465 (N_30465,N_30240,N_30028);
or U30466 (N_30466,N_30096,N_30147);
and U30467 (N_30467,N_30169,N_30049);
or U30468 (N_30468,N_30173,N_30053);
nor U30469 (N_30469,N_30011,N_30036);
nor U30470 (N_30470,N_30193,N_30084);
nor U30471 (N_30471,N_30203,N_30190);
nand U30472 (N_30472,N_30052,N_30196);
and U30473 (N_30473,N_30058,N_30089);
or U30474 (N_30474,N_30097,N_30085);
and U30475 (N_30475,N_30029,N_30045);
and U30476 (N_30476,N_30233,N_30087);
and U30477 (N_30477,N_30174,N_30056);
and U30478 (N_30478,N_30115,N_30062);
and U30479 (N_30479,N_30150,N_30052);
nand U30480 (N_30480,N_30119,N_30106);
nor U30481 (N_30481,N_30104,N_30148);
nand U30482 (N_30482,N_30053,N_30047);
xor U30483 (N_30483,N_30205,N_30085);
and U30484 (N_30484,N_30236,N_30219);
nand U30485 (N_30485,N_30165,N_30236);
or U30486 (N_30486,N_30174,N_30016);
nand U30487 (N_30487,N_30034,N_30049);
or U30488 (N_30488,N_30207,N_30164);
nor U30489 (N_30489,N_30141,N_30157);
xnor U30490 (N_30490,N_30127,N_30048);
nor U30491 (N_30491,N_30011,N_30051);
xor U30492 (N_30492,N_30236,N_30222);
xnor U30493 (N_30493,N_30023,N_30127);
and U30494 (N_30494,N_30176,N_30248);
nor U30495 (N_30495,N_30012,N_30027);
or U30496 (N_30496,N_30175,N_30156);
and U30497 (N_30497,N_30097,N_30233);
or U30498 (N_30498,N_30078,N_30066);
nor U30499 (N_30499,N_30043,N_30036);
nor U30500 (N_30500,N_30431,N_30473);
and U30501 (N_30501,N_30257,N_30321);
nand U30502 (N_30502,N_30487,N_30317);
nor U30503 (N_30503,N_30363,N_30447);
xor U30504 (N_30504,N_30357,N_30320);
or U30505 (N_30505,N_30377,N_30415);
nand U30506 (N_30506,N_30311,N_30366);
or U30507 (N_30507,N_30260,N_30337);
xor U30508 (N_30508,N_30486,N_30346);
nor U30509 (N_30509,N_30284,N_30325);
xnor U30510 (N_30510,N_30347,N_30448);
xor U30511 (N_30511,N_30371,N_30450);
nor U30512 (N_30512,N_30358,N_30334);
nand U30513 (N_30513,N_30414,N_30376);
xor U30514 (N_30514,N_30445,N_30453);
nor U30515 (N_30515,N_30352,N_30350);
and U30516 (N_30516,N_30250,N_30294);
nand U30517 (N_30517,N_30452,N_30485);
and U30518 (N_30518,N_30293,N_30396);
and U30519 (N_30519,N_30299,N_30307);
nor U30520 (N_30520,N_30411,N_30282);
nor U30521 (N_30521,N_30476,N_30316);
nand U30522 (N_30522,N_30392,N_30483);
or U30523 (N_30523,N_30412,N_30429);
or U30524 (N_30524,N_30289,N_30413);
nand U30525 (N_30525,N_30398,N_30298);
or U30526 (N_30526,N_30304,N_30460);
nor U30527 (N_30527,N_30335,N_30345);
or U30528 (N_30528,N_30281,N_30336);
xor U30529 (N_30529,N_30322,N_30467);
xnor U30530 (N_30530,N_30455,N_30261);
xnor U30531 (N_30531,N_30416,N_30446);
nand U30532 (N_30532,N_30463,N_30382);
and U30533 (N_30533,N_30339,N_30403);
and U30534 (N_30534,N_30305,N_30472);
or U30535 (N_30535,N_30441,N_30395);
nor U30536 (N_30536,N_30484,N_30297);
xor U30537 (N_30537,N_30433,N_30381);
nand U30538 (N_30538,N_30373,N_30349);
nand U30539 (N_30539,N_30313,N_30380);
and U30540 (N_30540,N_30418,N_30374);
and U30541 (N_30541,N_30389,N_30385);
nor U30542 (N_30542,N_30329,N_30259);
xnor U30543 (N_30543,N_30459,N_30405);
or U30544 (N_30544,N_30326,N_30456);
and U30545 (N_30545,N_30391,N_30400);
and U30546 (N_30546,N_30465,N_30383);
and U30547 (N_30547,N_30277,N_30470);
nand U30548 (N_30548,N_30399,N_30330);
and U30549 (N_30549,N_30471,N_30499);
nor U30550 (N_30550,N_30386,N_30296);
nor U30551 (N_30551,N_30478,N_30430);
and U30552 (N_30552,N_30319,N_30435);
xnor U30553 (N_30553,N_30360,N_30369);
or U30554 (N_30554,N_30475,N_30269);
xnor U30555 (N_30555,N_30268,N_30390);
or U30556 (N_30556,N_30401,N_30355);
and U30557 (N_30557,N_30315,N_30425);
xor U30558 (N_30558,N_30498,N_30362);
xnor U30559 (N_30559,N_30328,N_30312);
nand U30560 (N_30560,N_30443,N_30480);
nor U30561 (N_30561,N_30375,N_30440);
nor U30562 (N_30562,N_30341,N_30290);
or U30563 (N_30563,N_30333,N_30271);
nor U30564 (N_30564,N_30351,N_30353);
and U30565 (N_30565,N_30372,N_30303);
nand U30566 (N_30566,N_30370,N_30331);
or U30567 (N_30567,N_30428,N_30361);
nand U30568 (N_30568,N_30356,N_30457);
and U30569 (N_30569,N_30464,N_30344);
nor U30570 (N_30570,N_30496,N_30394);
xnor U30571 (N_30571,N_30327,N_30436);
xnor U30572 (N_30572,N_30340,N_30384);
nand U30573 (N_30573,N_30292,N_30492);
or U30574 (N_30574,N_30253,N_30488);
nor U30575 (N_30575,N_30308,N_30274);
or U30576 (N_30576,N_30302,N_30417);
or U30577 (N_30577,N_30388,N_30354);
and U30578 (N_30578,N_30427,N_30301);
nand U30579 (N_30579,N_30287,N_30423);
xnor U30580 (N_30580,N_30262,N_30309);
xnor U30581 (N_30581,N_30490,N_30468);
nor U30582 (N_30582,N_30367,N_30310);
and U30583 (N_30583,N_30404,N_30426);
nor U30584 (N_30584,N_30275,N_30266);
or U30585 (N_30585,N_30291,N_30458);
and U30586 (N_30586,N_30343,N_30379);
or U30587 (N_30587,N_30494,N_30397);
xnor U30588 (N_30588,N_30489,N_30437);
and U30589 (N_30589,N_30364,N_30306);
or U30590 (N_30590,N_30421,N_30466);
xnor U30591 (N_30591,N_30420,N_30348);
nor U30592 (N_30592,N_30407,N_30342);
or U30593 (N_30593,N_30479,N_30288);
nand U30594 (N_30594,N_30273,N_30387);
nand U30595 (N_30595,N_30264,N_30314);
xor U30596 (N_30596,N_30365,N_30497);
nand U30597 (N_30597,N_30267,N_30285);
nand U30598 (N_30598,N_30258,N_30481);
or U30599 (N_30599,N_30286,N_30451);
nor U30600 (N_30600,N_30477,N_30461);
nor U30601 (N_30601,N_30300,N_30359);
nor U30602 (N_30602,N_30434,N_30424);
nor U30603 (N_30603,N_30252,N_30255);
xor U30604 (N_30604,N_30402,N_30280);
nor U30605 (N_30605,N_30256,N_30263);
nand U30606 (N_30606,N_30491,N_30419);
and U30607 (N_30607,N_30368,N_30393);
nor U30608 (N_30608,N_30254,N_30283);
nand U30609 (N_30609,N_30332,N_30462);
xnor U30610 (N_30610,N_30265,N_30276);
nor U30611 (N_30611,N_30318,N_30409);
nor U30612 (N_30612,N_30449,N_30323);
nor U30613 (N_30613,N_30338,N_30439);
nand U30614 (N_30614,N_30270,N_30410);
nor U30615 (N_30615,N_30474,N_30378);
xor U30616 (N_30616,N_30422,N_30438);
or U30617 (N_30617,N_30272,N_30406);
xnor U30618 (N_30618,N_30279,N_30432);
and U30619 (N_30619,N_30251,N_30408);
or U30620 (N_30620,N_30444,N_30442);
nor U30621 (N_30621,N_30324,N_30482);
and U30622 (N_30622,N_30495,N_30278);
nor U30623 (N_30623,N_30295,N_30454);
nand U30624 (N_30624,N_30493,N_30469);
or U30625 (N_30625,N_30342,N_30352);
and U30626 (N_30626,N_30285,N_30409);
and U30627 (N_30627,N_30430,N_30290);
nor U30628 (N_30628,N_30403,N_30368);
nand U30629 (N_30629,N_30298,N_30358);
nand U30630 (N_30630,N_30372,N_30396);
and U30631 (N_30631,N_30364,N_30292);
xnor U30632 (N_30632,N_30300,N_30325);
nor U30633 (N_30633,N_30307,N_30466);
and U30634 (N_30634,N_30278,N_30447);
and U30635 (N_30635,N_30300,N_30458);
nor U30636 (N_30636,N_30484,N_30478);
and U30637 (N_30637,N_30338,N_30337);
nand U30638 (N_30638,N_30498,N_30393);
nand U30639 (N_30639,N_30278,N_30341);
nand U30640 (N_30640,N_30319,N_30499);
nor U30641 (N_30641,N_30384,N_30254);
nand U30642 (N_30642,N_30399,N_30467);
nand U30643 (N_30643,N_30413,N_30284);
nand U30644 (N_30644,N_30268,N_30393);
nor U30645 (N_30645,N_30474,N_30252);
nand U30646 (N_30646,N_30378,N_30414);
and U30647 (N_30647,N_30439,N_30457);
and U30648 (N_30648,N_30294,N_30386);
or U30649 (N_30649,N_30482,N_30466);
nand U30650 (N_30650,N_30391,N_30286);
xnor U30651 (N_30651,N_30339,N_30327);
or U30652 (N_30652,N_30426,N_30457);
xor U30653 (N_30653,N_30291,N_30444);
or U30654 (N_30654,N_30297,N_30250);
or U30655 (N_30655,N_30257,N_30263);
xnor U30656 (N_30656,N_30391,N_30498);
xor U30657 (N_30657,N_30267,N_30364);
nor U30658 (N_30658,N_30391,N_30469);
or U30659 (N_30659,N_30478,N_30485);
nand U30660 (N_30660,N_30404,N_30450);
and U30661 (N_30661,N_30407,N_30483);
nand U30662 (N_30662,N_30301,N_30496);
xor U30663 (N_30663,N_30452,N_30356);
xor U30664 (N_30664,N_30446,N_30324);
nor U30665 (N_30665,N_30324,N_30287);
or U30666 (N_30666,N_30457,N_30280);
nor U30667 (N_30667,N_30467,N_30282);
xnor U30668 (N_30668,N_30292,N_30407);
xor U30669 (N_30669,N_30264,N_30280);
xnor U30670 (N_30670,N_30397,N_30423);
nand U30671 (N_30671,N_30450,N_30437);
and U30672 (N_30672,N_30444,N_30445);
and U30673 (N_30673,N_30489,N_30346);
nand U30674 (N_30674,N_30367,N_30298);
nand U30675 (N_30675,N_30409,N_30469);
or U30676 (N_30676,N_30484,N_30360);
nand U30677 (N_30677,N_30406,N_30265);
and U30678 (N_30678,N_30488,N_30429);
or U30679 (N_30679,N_30343,N_30290);
nand U30680 (N_30680,N_30393,N_30485);
nor U30681 (N_30681,N_30307,N_30301);
or U30682 (N_30682,N_30374,N_30466);
nor U30683 (N_30683,N_30442,N_30279);
nand U30684 (N_30684,N_30393,N_30422);
or U30685 (N_30685,N_30443,N_30424);
xnor U30686 (N_30686,N_30364,N_30336);
nor U30687 (N_30687,N_30488,N_30355);
and U30688 (N_30688,N_30289,N_30449);
or U30689 (N_30689,N_30418,N_30465);
or U30690 (N_30690,N_30276,N_30355);
nand U30691 (N_30691,N_30417,N_30485);
xnor U30692 (N_30692,N_30275,N_30337);
nand U30693 (N_30693,N_30302,N_30328);
nor U30694 (N_30694,N_30332,N_30277);
nand U30695 (N_30695,N_30319,N_30321);
and U30696 (N_30696,N_30252,N_30342);
and U30697 (N_30697,N_30310,N_30279);
or U30698 (N_30698,N_30308,N_30303);
and U30699 (N_30699,N_30418,N_30296);
nor U30700 (N_30700,N_30352,N_30377);
or U30701 (N_30701,N_30306,N_30475);
or U30702 (N_30702,N_30475,N_30301);
and U30703 (N_30703,N_30265,N_30337);
nand U30704 (N_30704,N_30255,N_30286);
nor U30705 (N_30705,N_30352,N_30317);
nand U30706 (N_30706,N_30356,N_30443);
and U30707 (N_30707,N_30345,N_30456);
or U30708 (N_30708,N_30417,N_30449);
or U30709 (N_30709,N_30384,N_30430);
or U30710 (N_30710,N_30453,N_30409);
nand U30711 (N_30711,N_30393,N_30433);
xnor U30712 (N_30712,N_30273,N_30394);
and U30713 (N_30713,N_30414,N_30433);
nor U30714 (N_30714,N_30404,N_30491);
xor U30715 (N_30715,N_30485,N_30336);
xor U30716 (N_30716,N_30461,N_30462);
xnor U30717 (N_30717,N_30447,N_30330);
nor U30718 (N_30718,N_30425,N_30423);
nor U30719 (N_30719,N_30390,N_30273);
nor U30720 (N_30720,N_30362,N_30318);
xor U30721 (N_30721,N_30345,N_30479);
nor U30722 (N_30722,N_30481,N_30393);
xor U30723 (N_30723,N_30338,N_30266);
or U30724 (N_30724,N_30309,N_30441);
nor U30725 (N_30725,N_30281,N_30265);
xor U30726 (N_30726,N_30366,N_30457);
and U30727 (N_30727,N_30323,N_30398);
xor U30728 (N_30728,N_30307,N_30377);
nor U30729 (N_30729,N_30454,N_30471);
and U30730 (N_30730,N_30436,N_30281);
and U30731 (N_30731,N_30441,N_30450);
nor U30732 (N_30732,N_30439,N_30495);
nand U30733 (N_30733,N_30307,N_30298);
nor U30734 (N_30734,N_30346,N_30351);
nor U30735 (N_30735,N_30435,N_30410);
nor U30736 (N_30736,N_30286,N_30316);
and U30737 (N_30737,N_30258,N_30281);
nand U30738 (N_30738,N_30390,N_30497);
or U30739 (N_30739,N_30486,N_30260);
and U30740 (N_30740,N_30356,N_30431);
or U30741 (N_30741,N_30463,N_30283);
xor U30742 (N_30742,N_30368,N_30379);
and U30743 (N_30743,N_30434,N_30414);
nor U30744 (N_30744,N_30318,N_30413);
and U30745 (N_30745,N_30414,N_30349);
and U30746 (N_30746,N_30384,N_30320);
and U30747 (N_30747,N_30301,N_30290);
xnor U30748 (N_30748,N_30477,N_30356);
and U30749 (N_30749,N_30457,N_30272);
nor U30750 (N_30750,N_30660,N_30540);
and U30751 (N_30751,N_30694,N_30528);
and U30752 (N_30752,N_30560,N_30678);
xnor U30753 (N_30753,N_30650,N_30740);
nand U30754 (N_30754,N_30716,N_30556);
or U30755 (N_30755,N_30683,N_30729);
xnor U30756 (N_30756,N_30693,N_30685);
or U30757 (N_30757,N_30561,N_30669);
or U30758 (N_30758,N_30645,N_30712);
or U30759 (N_30759,N_30552,N_30646);
nor U30760 (N_30760,N_30732,N_30743);
or U30761 (N_30761,N_30546,N_30591);
nor U30762 (N_30762,N_30704,N_30526);
xnor U30763 (N_30763,N_30698,N_30737);
nand U30764 (N_30764,N_30639,N_30612);
or U30765 (N_30765,N_30534,N_30714);
or U30766 (N_30766,N_30619,N_30609);
and U30767 (N_30767,N_30731,N_30558);
nor U30768 (N_30768,N_30705,N_30511);
nand U30769 (N_30769,N_30575,N_30718);
nor U30770 (N_30770,N_30519,N_30583);
nand U30771 (N_30771,N_30506,N_30687);
nor U30772 (N_30772,N_30626,N_30539);
and U30773 (N_30773,N_30501,N_30670);
nand U30774 (N_30774,N_30588,N_30620);
nor U30775 (N_30775,N_30565,N_30621);
nor U30776 (N_30776,N_30702,N_30638);
or U30777 (N_30777,N_30636,N_30542);
xnor U30778 (N_30778,N_30708,N_30677);
or U30779 (N_30779,N_30628,N_30727);
nor U30780 (N_30780,N_30746,N_30610);
nor U30781 (N_30781,N_30742,N_30662);
and U30782 (N_30782,N_30553,N_30555);
or U30783 (N_30783,N_30520,N_30635);
nor U30784 (N_30784,N_30672,N_30548);
xnor U30785 (N_30785,N_30514,N_30541);
nand U30786 (N_30786,N_30507,N_30529);
nor U30787 (N_30787,N_30574,N_30533);
xnor U30788 (N_30788,N_30518,N_30577);
nand U30789 (N_30789,N_30625,N_30633);
and U30790 (N_30790,N_30689,N_30654);
nor U30791 (N_30791,N_30691,N_30631);
and U30792 (N_30792,N_30744,N_30713);
nand U30793 (N_30793,N_30584,N_30652);
nand U30794 (N_30794,N_30585,N_30594);
nand U30795 (N_30795,N_30724,N_30606);
and U30796 (N_30796,N_30728,N_30597);
or U30797 (N_30797,N_30655,N_30668);
nand U30798 (N_30798,N_30617,N_30525);
nor U30799 (N_30799,N_30527,N_30503);
nor U30800 (N_30800,N_30537,N_30564);
nor U30801 (N_30801,N_30675,N_30692);
or U30802 (N_30802,N_30578,N_30624);
nand U30803 (N_30803,N_30661,N_30706);
xnor U30804 (N_30804,N_30730,N_30695);
xnor U30805 (N_30805,N_30641,N_30523);
and U30806 (N_30806,N_30642,N_30616);
nor U30807 (N_30807,N_30604,N_30508);
and U30808 (N_30808,N_30592,N_30711);
or U30809 (N_30809,N_30632,N_30674);
xor U30810 (N_30810,N_30559,N_30657);
or U30811 (N_30811,N_30515,N_30627);
nor U30812 (N_30812,N_30573,N_30681);
nand U30813 (N_30813,N_30502,N_30690);
and U30814 (N_30814,N_30726,N_30747);
xor U30815 (N_30815,N_30658,N_30586);
nand U30816 (N_30816,N_30580,N_30505);
xnor U30817 (N_30817,N_30521,N_30673);
nand U30818 (N_30818,N_30739,N_30563);
and U30819 (N_30819,N_30719,N_30651);
xnor U30820 (N_30820,N_30733,N_30615);
xnor U30821 (N_30821,N_30500,N_30710);
nand U30822 (N_30822,N_30684,N_30579);
or U30823 (N_30823,N_30699,N_30667);
nor U30824 (N_30824,N_30554,N_30587);
nor U30825 (N_30825,N_30663,N_30545);
and U30826 (N_30826,N_30600,N_30601);
and U30827 (N_30827,N_30530,N_30649);
nor U30828 (N_30828,N_30735,N_30623);
or U30829 (N_30829,N_30504,N_30644);
and U30830 (N_30830,N_30640,N_30725);
or U30831 (N_30831,N_30572,N_30569);
xor U30832 (N_30832,N_30590,N_30630);
nor U30833 (N_30833,N_30602,N_30535);
xnor U30834 (N_30834,N_30679,N_30582);
or U30835 (N_30835,N_30571,N_30707);
or U30836 (N_30836,N_30656,N_30532);
nand U30837 (N_30837,N_30576,N_30614);
nor U30838 (N_30838,N_30538,N_30589);
nand U30839 (N_30839,N_30720,N_30688);
and U30840 (N_30840,N_30603,N_30509);
or U30841 (N_30841,N_30550,N_30664);
and U30842 (N_30842,N_30653,N_30647);
or U30843 (N_30843,N_30721,N_30516);
xnor U30844 (N_30844,N_30512,N_30596);
xnor U30845 (N_30845,N_30715,N_30531);
or U30846 (N_30846,N_30517,N_30749);
and U30847 (N_30847,N_30543,N_30593);
nand U30848 (N_30848,N_30723,N_30607);
nor U30849 (N_30849,N_30736,N_30709);
xor U30850 (N_30850,N_30637,N_30549);
nand U30851 (N_30851,N_30717,N_30557);
or U30852 (N_30852,N_30666,N_30547);
or U30853 (N_30853,N_30567,N_30700);
or U30854 (N_30854,N_30599,N_30513);
nor U30855 (N_30855,N_30738,N_30510);
xor U30856 (N_30856,N_30703,N_30665);
and U30857 (N_30857,N_30734,N_30611);
or U30858 (N_30858,N_30622,N_30659);
or U30859 (N_30859,N_30748,N_30568);
xor U30860 (N_30860,N_30595,N_30570);
and U30861 (N_30861,N_30686,N_30544);
and U30862 (N_30862,N_30745,N_30680);
or U30863 (N_30863,N_30741,N_30696);
nand U30864 (N_30864,N_30551,N_30618);
nand U30865 (N_30865,N_30671,N_30608);
nor U30866 (N_30866,N_30524,N_30581);
or U30867 (N_30867,N_30697,N_30629);
nor U30868 (N_30868,N_30722,N_30522);
and U30869 (N_30869,N_30566,N_30598);
and U30870 (N_30870,N_30648,N_30676);
xor U30871 (N_30871,N_30682,N_30634);
nand U30872 (N_30872,N_30701,N_30643);
xor U30873 (N_30873,N_30613,N_30605);
nor U30874 (N_30874,N_30536,N_30562);
or U30875 (N_30875,N_30574,N_30719);
or U30876 (N_30876,N_30594,N_30587);
and U30877 (N_30877,N_30679,N_30568);
and U30878 (N_30878,N_30687,N_30597);
and U30879 (N_30879,N_30524,N_30567);
nand U30880 (N_30880,N_30506,N_30615);
or U30881 (N_30881,N_30570,N_30583);
nand U30882 (N_30882,N_30675,N_30609);
nand U30883 (N_30883,N_30588,N_30708);
nand U30884 (N_30884,N_30552,N_30641);
and U30885 (N_30885,N_30505,N_30546);
or U30886 (N_30886,N_30550,N_30533);
and U30887 (N_30887,N_30653,N_30722);
nand U30888 (N_30888,N_30638,N_30579);
or U30889 (N_30889,N_30510,N_30528);
nand U30890 (N_30890,N_30552,N_30691);
nand U30891 (N_30891,N_30722,N_30611);
nor U30892 (N_30892,N_30647,N_30686);
and U30893 (N_30893,N_30524,N_30621);
or U30894 (N_30894,N_30574,N_30664);
nor U30895 (N_30895,N_30679,N_30589);
and U30896 (N_30896,N_30720,N_30629);
or U30897 (N_30897,N_30729,N_30560);
nor U30898 (N_30898,N_30565,N_30711);
or U30899 (N_30899,N_30503,N_30500);
nand U30900 (N_30900,N_30747,N_30569);
nand U30901 (N_30901,N_30704,N_30542);
nand U30902 (N_30902,N_30579,N_30692);
nand U30903 (N_30903,N_30715,N_30580);
or U30904 (N_30904,N_30585,N_30612);
and U30905 (N_30905,N_30674,N_30539);
xnor U30906 (N_30906,N_30566,N_30746);
and U30907 (N_30907,N_30630,N_30546);
or U30908 (N_30908,N_30506,N_30517);
and U30909 (N_30909,N_30629,N_30587);
xor U30910 (N_30910,N_30704,N_30743);
xnor U30911 (N_30911,N_30575,N_30561);
nand U30912 (N_30912,N_30556,N_30528);
or U30913 (N_30913,N_30585,N_30715);
nor U30914 (N_30914,N_30557,N_30701);
or U30915 (N_30915,N_30733,N_30663);
xnor U30916 (N_30916,N_30674,N_30604);
xor U30917 (N_30917,N_30632,N_30681);
nand U30918 (N_30918,N_30604,N_30568);
or U30919 (N_30919,N_30631,N_30552);
and U30920 (N_30920,N_30647,N_30680);
or U30921 (N_30921,N_30628,N_30670);
and U30922 (N_30922,N_30708,N_30574);
xnor U30923 (N_30923,N_30691,N_30528);
and U30924 (N_30924,N_30722,N_30714);
or U30925 (N_30925,N_30727,N_30718);
nor U30926 (N_30926,N_30514,N_30612);
and U30927 (N_30927,N_30735,N_30641);
nand U30928 (N_30928,N_30739,N_30576);
xor U30929 (N_30929,N_30528,N_30602);
nand U30930 (N_30930,N_30506,N_30519);
xnor U30931 (N_30931,N_30725,N_30650);
nand U30932 (N_30932,N_30599,N_30512);
xor U30933 (N_30933,N_30671,N_30740);
or U30934 (N_30934,N_30701,N_30566);
or U30935 (N_30935,N_30569,N_30563);
or U30936 (N_30936,N_30719,N_30606);
nand U30937 (N_30937,N_30567,N_30610);
or U30938 (N_30938,N_30633,N_30686);
nand U30939 (N_30939,N_30726,N_30578);
nor U30940 (N_30940,N_30739,N_30669);
nand U30941 (N_30941,N_30561,N_30505);
or U30942 (N_30942,N_30583,N_30613);
nor U30943 (N_30943,N_30700,N_30571);
nand U30944 (N_30944,N_30685,N_30692);
xor U30945 (N_30945,N_30556,N_30650);
nand U30946 (N_30946,N_30554,N_30676);
or U30947 (N_30947,N_30710,N_30575);
nor U30948 (N_30948,N_30542,N_30511);
nor U30949 (N_30949,N_30643,N_30683);
and U30950 (N_30950,N_30525,N_30532);
nand U30951 (N_30951,N_30749,N_30695);
nand U30952 (N_30952,N_30534,N_30573);
xnor U30953 (N_30953,N_30681,N_30605);
or U30954 (N_30954,N_30512,N_30586);
nor U30955 (N_30955,N_30625,N_30675);
xnor U30956 (N_30956,N_30529,N_30513);
xor U30957 (N_30957,N_30553,N_30738);
or U30958 (N_30958,N_30622,N_30639);
nand U30959 (N_30959,N_30733,N_30670);
and U30960 (N_30960,N_30667,N_30637);
nor U30961 (N_30961,N_30709,N_30609);
nand U30962 (N_30962,N_30566,N_30744);
xor U30963 (N_30963,N_30555,N_30515);
nand U30964 (N_30964,N_30746,N_30548);
nand U30965 (N_30965,N_30594,N_30632);
xor U30966 (N_30966,N_30554,N_30711);
nand U30967 (N_30967,N_30577,N_30633);
nor U30968 (N_30968,N_30544,N_30694);
or U30969 (N_30969,N_30651,N_30588);
and U30970 (N_30970,N_30540,N_30717);
nor U30971 (N_30971,N_30720,N_30656);
and U30972 (N_30972,N_30677,N_30740);
nand U30973 (N_30973,N_30563,N_30728);
nor U30974 (N_30974,N_30612,N_30542);
and U30975 (N_30975,N_30603,N_30545);
and U30976 (N_30976,N_30638,N_30710);
xnor U30977 (N_30977,N_30593,N_30659);
nand U30978 (N_30978,N_30507,N_30601);
or U30979 (N_30979,N_30728,N_30714);
nor U30980 (N_30980,N_30560,N_30697);
nand U30981 (N_30981,N_30636,N_30528);
nor U30982 (N_30982,N_30539,N_30722);
and U30983 (N_30983,N_30677,N_30597);
xnor U30984 (N_30984,N_30669,N_30733);
or U30985 (N_30985,N_30716,N_30746);
nor U30986 (N_30986,N_30577,N_30641);
xnor U30987 (N_30987,N_30554,N_30512);
or U30988 (N_30988,N_30638,N_30646);
nand U30989 (N_30989,N_30572,N_30539);
nand U30990 (N_30990,N_30572,N_30744);
xnor U30991 (N_30991,N_30610,N_30722);
or U30992 (N_30992,N_30514,N_30674);
nor U30993 (N_30993,N_30721,N_30555);
and U30994 (N_30994,N_30608,N_30595);
and U30995 (N_30995,N_30648,N_30528);
or U30996 (N_30996,N_30583,N_30573);
nand U30997 (N_30997,N_30634,N_30532);
or U30998 (N_30998,N_30544,N_30566);
nand U30999 (N_30999,N_30690,N_30560);
and U31000 (N_31000,N_30860,N_30834);
nand U31001 (N_31001,N_30854,N_30919);
xnor U31002 (N_31002,N_30873,N_30986);
xor U31003 (N_31003,N_30900,N_30908);
nand U31004 (N_31004,N_30903,N_30935);
nor U31005 (N_31005,N_30942,N_30819);
xnor U31006 (N_31006,N_30941,N_30815);
or U31007 (N_31007,N_30996,N_30766);
and U31008 (N_31008,N_30825,N_30969);
or U31009 (N_31009,N_30938,N_30852);
and U31010 (N_31010,N_30764,N_30929);
nor U31011 (N_31011,N_30803,N_30799);
or U31012 (N_31012,N_30896,N_30811);
or U31013 (N_31013,N_30875,N_30800);
and U31014 (N_31014,N_30792,N_30933);
xnor U31015 (N_31015,N_30756,N_30925);
xnor U31016 (N_31016,N_30865,N_30977);
nor U31017 (N_31017,N_30808,N_30951);
nor U31018 (N_31018,N_30840,N_30774);
nor U31019 (N_31019,N_30778,N_30769);
and U31020 (N_31020,N_30861,N_30892);
xor U31021 (N_31021,N_30971,N_30761);
nor U31022 (N_31022,N_30975,N_30985);
nand U31023 (N_31023,N_30777,N_30899);
nor U31024 (N_31024,N_30857,N_30856);
and U31025 (N_31025,N_30902,N_30968);
nand U31026 (N_31026,N_30979,N_30920);
and U31027 (N_31027,N_30895,N_30906);
and U31028 (N_31028,N_30832,N_30960);
nor U31029 (N_31029,N_30930,N_30783);
nand U31030 (N_31030,N_30984,N_30904);
nand U31031 (N_31031,N_30912,N_30788);
nor U31032 (N_31032,N_30995,N_30779);
xnor U31033 (N_31033,N_30916,N_30866);
nor U31034 (N_31034,N_30793,N_30915);
or U31035 (N_31035,N_30822,N_30926);
nor U31036 (N_31036,N_30901,N_30849);
nand U31037 (N_31037,N_30872,N_30956);
nor U31038 (N_31038,N_30970,N_30843);
and U31039 (N_31039,N_30999,N_30871);
and U31040 (N_31040,N_30889,N_30961);
or U31041 (N_31041,N_30982,N_30905);
or U31042 (N_31042,N_30824,N_30768);
nor U31043 (N_31043,N_30910,N_30772);
xnor U31044 (N_31044,N_30812,N_30967);
nand U31045 (N_31045,N_30785,N_30802);
or U31046 (N_31046,N_30964,N_30936);
xor U31047 (N_31047,N_30878,N_30787);
and U31048 (N_31048,N_30835,N_30923);
nor U31049 (N_31049,N_30810,N_30952);
nor U31050 (N_31050,N_30775,N_30953);
or U31051 (N_31051,N_30939,N_30876);
xnor U31052 (N_31052,N_30780,N_30751);
nor U31053 (N_31053,N_30750,N_30911);
xnor U31054 (N_31054,N_30789,N_30838);
and U31055 (N_31055,N_30944,N_30993);
nor U31056 (N_31056,N_30830,N_30868);
and U31057 (N_31057,N_30864,N_30885);
and U31058 (N_31058,N_30989,N_30886);
xor U31059 (N_31059,N_30781,N_30796);
nor U31060 (N_31060,N_30949,N_30874);
nor U31061 (N_31061,N_30859,N_30898);
xor U31062 (N_31062,N_30927,N_30757);
or U31063 (N_31063,N_30829,N_30945);
xor U31064 (N_31064,N_30882,N_30847);
and U31065 (N_31065,N_30786,N_30831);
or U31066 (N_31066,N_30821,N_30978);
xnor U31067 (N_31067,N_30758,N_30770);
nor U31068 (N_31068,N_30937,N_30817);
nor U31069 (N_31069,N_30963,N_30994);
xnor U31070 (N_31070,N_30828,N_30869);
nor U31071 (N_31071,N_30932,N_30890);
and U31072 (N_31072,N_30807,N_30752);
xor U31073 (N_31073,N_30947,N_30836);
nor U31074 (N_31074,N_30813,N_30897);
and U31075 (N_31075,N_30958,N_30790);
nor U31076 (N_31076,N_30797,N_30983);
and U31077 (N_31077,N_30974,N_30826);
xnor U31078 (N_31078,N_30981,N_30791);
or U31079 (N_31079,N_30921,N_30760);
nor U31080 (N_31080,N_30759,N_30998);
nand U31081 (N_31081,N_30881,N_30883);
nor U31082 (N_31082,N_30755,N_30842);
xor U31083 (N_31083,N_30798,N_30990);
and U31084 (N_31084,N_30833,N_30848);
or U31085 (N_31085,N_30863,N_30965);
or U31086 (N_31086,N_30907,N_30794);
nand U31087 (N_31087,N_30943,N_30893);
xor U31088 (N_31088,N_30820,N_30827);
nor U31089 (N_31089,N_30880,N_30959);
nor U31090 (N_31090,N_30851,N_30913);
xor U31091 (N_31091,N_30955,N_30972);
xnor U31092 (N_31092,N_30818,N_30934);
nand U31093 (N_31093,N_30784,N_30924);
nor U31094 (N_31094,N_30948,N_30773);
nand U31095 (N_31095,N_30877,N_30962);
nand U31096 (N_31096,N_30917,N_30884);
nor U31097 (N_31097,N_30853,N_30806);
xnor U31098 (N_31098,N_30763,N_30891);
nand U31099 (N_31099,N_30914,N_30894);
or U31100 (N_31100,N_30809,N_30862);
or U31101 (N_31101,N_30950,N_30858);
or U31102 (N_31102,N_30887,N_30795);
or U31103 (N_31103,N_30844,N_30816);
nand U31104 (N_31104,N_30957,N_30767);
xnor U31105 (N_31105,N_30992,N_30801);
or U31106 (N_31106,N_30771,N_30931);
nand U31107 (N_31107,N_30753,N_30867);
or U31108 (N_31108,N_30918,N_30946);
xor U31109 (N_31109,N_30855,N_30776);
nor U31110 (N_31110,N_30762,N_30870);
and U31111 (N_31111,N_30940,N_30754);
and U31112 (N_31112,N_30837,N_30805);
nor U31113 (N_31113,N_30888,N_30973);
nor U31114 (N_31114,N_30988,N_30928);
nor U31115 (N_31115,N_30954,N_30980);
xor U31116 (N_31116,N_30909,N_30839);
xnor U31117 (N_31117,N_30850,N_30823);
xnor U31118 (N_31118,N_30782,N_30922);
nand U31119 (N_31119,N_30879,N_30841);
and U31120 (N_31120,N_30997,N_30845);
xor U31121 (N_31121,N_30991,N_30976);
and U31122 (N_31122,N_30966,N_30765);
or U31123 (N_31123,N_30804,N_30846);
nand U31124 (N_31124,N_30814,N_30987);
nor U31125 (N_31125,N_30957,N_30928);
and U31126 (N_31126,N_30826,N_30838);
or U31127 (N_31127,N_30904,N_30923);
nand U31128 (N_31128,N_30812,N_30916);
or U31129 (N_31129,N_30859,N_30969);
and U31130 (N_31130,N_30787,N_30877);
and U31131 (N_31131,N_30924,N_30901);
nand U31132 (N_31132,N_30928,N_30841);
xnor U31133 (N_31133,N_30918,N_30818);
nand U31134 (N_31134,N_30896,N_30801);
nand U31135 (N_31135,N_30829,N_30999);
nor U31136 (N_31136,N_30772,N_30905);
xor U31137 (N_31137,N_30923,N_30764);
or U31138 (N_31138,N_30911,N_30846);
xor U31139 (N_31139,N_30924,N_30849);
nor U31140 (N_31140,N_30917,N_30765);
and U31141 (N_31141,N_30970,N_30924);
nor U31142 (N_31142,N_30914,N_30886);
nand U31143 (N_31143,N_30964,N_30951);
xor U31144 (N_31144,N_30866,N_30774);
nor U31145 (N_31145,N_30823,N_30954);
or U31146 (N_31146,N_30818,N_30823);
or U31147 (N_31147,N_30840,N_30865);
or U31148 (N_31148,N_30882,N_30824);
or U31149 (N_31149,N_30955,N_30937);
or U31150 (N_31150,N_30992,N_30851);
nor U31151 (N_31151,N_30944,N_30776);
nand U31152 (N_31152,N_30893,N_30808);
nand U31153 (N_31153,N_30776,N_30931);
or U31154 (N_31154,N_30750,N_30833);
xor U31155 (N_31155,N_30924,N_30889);
xnor U31156 (N_31156,N_30883,N_30901);
or U31157 (N_31157,N_30902,N_30807);
or U31158 (N_31158,N_30831,N_30951);
nand U31159 (N_31159,N_30898,N_30858);
xor U31160 (N_31160,N_30761,N_30967);
nand U31161 (N_31161,N_30855,N_30856);
or U31162 (N_31162,N_30850,N_30964);
or U31163 (N_31163,N_30760,N_30966);
nor U31164 (N_31164,N_30775,N_30926);
xor U31165 (N_31165,N_30834,N_30796);
and U31166 (N_31166,N_30853,N_30979);
nand U31167 (N_31167,N_30890,N_30999);
and U31168 (N_31168,N_30799,N_30928);
or U31169 (N_31169,N_30831,N_30888);
nand U31170 (N_31170,N_30956,N_30904);
and U31171 (N_31171,N_30831,N_30886);
nor U31172 (N_31172,N_30999,N_30959);
xnor U31173 (N_31173,N_30874,N_30779);
and U31174 (N_31174,N_30841,N_30970);
or U31175 (N_31175,N_30866,N_30815);
and U31176 (N_31176,N_30784,N_30869);
and U31177 (N_31177,N_30947,N_30883);
nand U31178 (N_31178,N_30827,N_30883);
nor U31179 (N_31179,N_30805,N_30868);
xnor U31180 (N_31180,N_30925,N_30880);
and U31181 (N_31181,N_30763,N_30995);
xnor U31182 (N_31182,N_30958,N_30859);
or U31183 (N_31183,N_30964,N_30891);
nand U31184 (N_31184,N_30869,N_30859);
nand U31185 (N_31185,N_30903,N_30989);
and U31186 (N_31186,N_30800,N_30855);
or U31187 (N_31187,N_30994,N_30890);
nand U31188 (N_31188,N_30906,N_30896);
nand U31189 (N_31189,N_30941,N_30816);
or U31190 (N_31190,N_30900,N_30755);
and U31191 (N_31191,N_30974,N_30861);
xnor U31192 (N_31192,N_30833,N_30905);
nor U31193 (N_31193,N_30886,N_30779);
and U31194 (N_31194,N_30872,N_30985);
xnor U31195 (N_31195,N_30787,N_30943);
nor U31196 (N_31196,N_30867,N_30889);
xnor U31197 (N_31197,N_30902,N_30831);
and U31198 (N_31198,N_30878,N_30984);
or U31199 (N_31199,N_30957,N_30992);
or U31200 (N_31200,N_30797,N_30796);
nand U31201 (N_31201,N_30999,N_30891);
nand U31202 (N_31202,N_30827,N_30859);
and U31203 (N_31203,N_30888,N_30754);
nor U31204 (N_31204,N_30892,N_30946);
or U31205 (N_31205,N_30991,N_30928);
and U31206 (N_31206,N_30881,N_30810);
or U31207 (N_31207,N_30990,N_30811);
xnor U31208 (N_31208,N_30875,N_30900);
nor U31209 (N_31209,N_30861,N_30995);
and U31210 (N_31210,N_30982,N_30854);
or U31211 (N_31211,N_30894,N_30997);
nand U31212 (N_31212,N_30908,N_30880);
nor U31213 (N_31213,N_30848,N_30759);
nor U31214 (N_31214,N_30893,N_30957);
and U31215 (N_31215,N_30766,N_30778);
and U31216 (N_31216,N_30889,N_30929);
and U31217 (N_31217,N_30886,N_30912);
nand U31218 (N_31218,N_30784,N_30757);
or U31219 (N_31219,N_30757,N_30891);
nand U31220 (N_31220,N_30771,N_30785);
or U31221 (N_31221,N_30987,N_30775);
nand U31222 (N_31222,N_30835,N_30818);
or U31223 (N_31223,N_30957,N_30801);
or U31224 (N_31224,N_30850,N_30998);
xnor U31225 (N_31225,N_30962,N_30846);
and U31226 (N_31226,N_30843,N_30775);
or U31227 (N_31227,N_30941,N_30782);
and U31228 (N_31228,N_30792,N_30780);
nand U31229 (N_31229,N_30778,N_30819);
nand U31230 (N_31230,N_30773,N_30969);
nand U31231 (N_31231,N_30943,N_30878);
nand U31232 (N_31232,N_30837,N_30798);
or U31233 (N_31233,N_30958,N_30781);
xor U31234 (N_31234,N_30804,N_30916);
or U31235 (N_31235,N_30782,N_30834);
or U31236 (N_31236,N_30941,N_30889);
xor U31237 (N_31237,N_30787,N_30751);
nor U31238 (N_31238,N_30925,N_30944);
nor U31239 (N_31239,N_30872,N_30838);
xor U31240 (N_31240,N_30844,N_30873);
nand U31241 (N_31241,N_30884,N_30835);
nand U31242 (N_31242,N_30778,N_30869);
and U31243 (N_31243,N_30994,N_30937);
and U31244 (N_31244,N_30821,N_30951);
or U31245 (N_31245,N_30930,N_30782);
xnor U31246 (N_31246,N_30900,N_30782);
and U31247 (N_31247,N_30795,N_30934);
or U31248 (N_31248,N_30990,N_30893);
or U31249 (N_31249,N_30965,N_30913);
nand U31250 (N_31250,N_31190,N_31113);
xnor U31251 (N_31251,N_31175,N_31046);
and U31252 (N_31252,N_31106,N_31216);
or U31253 (N_31253,N_31018,N_31017);
and U31254 (N_31254,N_31029,N_31158);
or U31255 (N_31255,N_31003,N_31191);
xnor U31256 (N_31256,N_31064,N_31015);
and U31257 (N_31257,N_31233,N_31164);
or U31258 (N_31258,N_31173,N_31187);
or U31259 (N_31259,N_31068,N_31119);
or U31260 (N_31260,N_31202,N_31193);
xnor U31261 (N_31261,N_31053,N_31041);
xor U31262 (N_31262,N_31085,N_31004);
nor U31263 (N_31263,N_31063,N_31033);
nor U31264 (N_31264,N_31122,N_31206);
xnor U31265 (N_31265,N_31146,N_31060);
nor U31266 (N_31266,N_31209,N_31066);
and U31267 (N_31267,N_31176,N_31139);
and U31268 (N_31268,N_31054,N_31249);
and U31269 (N_31269,N_31155,N_31081);
or U31270 (N_31270,N_31088,N_31099);
and U31271 (N_31271,N_31080,N_31042);
or U31272 (N_31272,N_31074,N_31138);
nand U31273 (N_31273,N_31096,N_31192);
xnor U31274 (N_31274,N_31133,N_31028);
or U31275 (N_31275,N_31157,N_31174);
nor U31276 (N_31276,N_31211,N_31087);
xnor U31277 (N_31277,N_31184,N_31023);
xnor U31278 (N_31278,N_31130,N_31245);
nand U31279 (N_31279,N_31210,N_31246);
or U31280 (N_31280,N_31230,N_31144);
or U31281 (N_31281,N_31071,N_31016);
nand U31282 (N_31282,N_31105,N_31201);
nor U31283 (N_31283,N_31057,N_31231);
nor U31284 (N_31284,N_31083,N_31020);
nor U31285 (N_31285,N_31218,N_31115);
or U31286 (N_31286,N_31142,N_31059);
xnor U31287 (N_31287,N_31019,N_31215);
or U31288 (N_31288,N_31076,N_31200);
nand U31289 (N_31289,N_31093,N_31135);
xor U31290 (N_31290,N_31150,N_31036);
or U31291 (N_31291,N_31167,N_31109);
nand U31292 (N_31292,N_31182,N_31049);
or U31293 (N_31293,N_31243,N_31108);
xnor U31294 (N_31294,N_31082,N_31116);
nand U31295 (N_31295,N_31025,N_31178);
and U31296 (N_31296,N_31011,N_31153);
nor U31297 (N_31297,N_31169,N_31128);
and U31298 (N_31298,N_31100,N_31072);
and U31299 (N_31299,N_31196,N_31168);
xnor U31300 (N_31300,N_31172,N_31156);
xor U31301 (N_31301,N_31125,N_31188);
nand U31302 (N_31302,N_31079,N_31183);
xor U31303 (N_31303,N_31037,N_31213);
and U31304 (N_31304,N_31091,N_31006);
and U31305 (N_31305,N_31204,N_31152);
xor U31306 (N_31306,N_31198,N_31160);
nand U31307 (N_31307,N_31131,N_31166);
or U31308 (N_31308,N_31217,N_31141);
nor U31309 (N_31309,N_31244,N_31110);
and U31310 (N_31310,N_31008,N_31061);
nand U31311 (N_31311,N_31161,N_31219);
xnor U31312 (N_31312,N_31043,N_31039);
nand U31313 (N_31313,N_31097,N_31239);
and U31314 (N_31314,N_31001,N_31228);
and U31315 (N_31315,N_31031,N_31225);
or U31316 (N_31316,N_31129,N_31002);
nor U31317 (N_31317,N_31189,N_31170);
and U31318 (N_31318,N_31095,N_31048);
nor U31319 (N_31319,N_31154,N_31073);
nand U31320 (N_31320,N_31009,N_31229);
or U31321 (N_31321,N_31112,N_31121);
and U31322 (N_31322,N_31226,N_31007);
nor U31323 (N_31323,N_31165,N_31247);
or U31324 (N_31324,N_31094,N_31092);
nand U31325 (N_31325,N_31140,N_31104);
xor U31326 (N_31326,N_31137,N_31021);
nand U31327 (N_31327,N_31207,N_31084);
nand U31328 (N_31328,N_31062,N_31223);
and U31329 (N_31329,N_31237,N_31050);
xor U31330 (N_31330,N_31222,N_31051);
xnor U31331 (N_31331,N_31038,N_31199);
or U31332 (N_31332,N_31220,N_31194);
or U31333 (N_31333,N_31055,N_31221);
nor U31334 (N_31334,N_31089,N_31040);
or U31335 (N_31335,N_31232,N_31123);
nand U31336 (N_31336,N_31058,N_31236);
or U31337 (N_31337,N_31102,N_31024);
nand U31338 (N_31338,N_31159,N_31056);
xor U31339 (N_31339,N_31124,N_31052);
nand U31340 (N_31340,N_31151,N_31235);
and U31341 (N_31341,N_31070,N_31208);
nor U31342 (N_31342,N_31238,N_31111);
nor U31343 (N_31343,N_31162,N_31047);
nand U31344 (N_31344,N_31134,N_31114);
nand U31345 (N_31345,N_31034,N_31045);
or U31346 (N_31346,N_31203,N_31101);
nand U31347 (N_31347,N_31242,N_31241);
nand U31348 (N_31348,N_31132,N_31013);
nand U31349 (N_31349,N_31148,N_31214);
or U31350 (N_31350,N_31143,N_31035);
nor U31351 (N_31351,N_31224,N_31149);
and U31352 (N_31352,N_31118,N_31012);
and U31353 (N_31353,N_31186,N_31117);
nand U31354 (N_31354,N_31147,N_31163);
nor U31355 (N_31355,N_31032,N_31090);
and U31356 (N_31356,N_31127,N_31044);
nor U31357 (N_31357,N_31179,N_31136);
nor U31358 (N_31358,N_31107,N_31069);
or U31359 (N_31359,N_31030,N_31212);
and U31360 (N_31360,N_31180,N_31065);
nand U31361 (N_31361,N_31077,N_31126);
and U31362 (N_31362,N_31075,N_31022);
and U31363 (N_31363,N_31205,N_31067);
xor U31364 (N_31364,N_31248,N_31185);
and U31365 (N_31365,N_31120,N_31234);
nor U31366 (N_31366,N_31098,N_31014);
nor U31367 (N_31367,N_31103,N_31197);
nor U31368 (N_31368,N_31010,N_31026);
and U31369 (N_31369,N_31027,N_31227);
xnor U31370 (N_31370,N_31000,N_31145);
and U31371 (N_31371,N_31195,N_31005);
or U31372 (N_31372,N_31171,N_31078);
nand U31373 (N_31373,N_31181,N_31086);
or U31374 (N_31374,N_31240,N_31177);
nand U31375 (N_31375,N_31129,N_31212);
xnor U31376 (N_31376,N_31017,N_31030);
or U31377 (N_31377,N_31097,N_31013);
nand U31378 (N_31378,N_31248,N_31191);
or U31379 (N_31379,N_31220,N_31004);
nand U31380 (N_31380,N_31235,N_31087);
or U31381 (N_31381,N_31028,N_31120);
nand U31382 (N_31382,N_31029,N_31123);
nand U31383 (N_31383,N_31221,N_31081);
nor U31384 (N_31384,N_31075,N_31063);
or U31385 (N_31385,N_31085,N_31133);
nand U31386 (N_31386,N_31139,N_31013);
nor U31387 (N_31387,N_31216,N_31033);
nand U31388 (N_31388,N_31038,N_31165);
or U31389 (N_31389,N_31072,N_31044);
nand U31390 (N_31390,N_31144,N_31193);
and U31391 (N_31391,N_31070,N_31249);
xor U31392 (N_31392,N_31014,N_31111);
and U31393 (N_31393,N_31095,N_31205);
or U31394 (N_31394,N_31003,N_31145);
or U31395 (N_31395,N_31103,N_31160);
or U31396 (N_31396,N_31134,N_31050);
and U31397 (N_31397,N_31229,N_31240);
nor U31398 (N_31398,N_31090,N_31112);
and U31399 (N_31399,N_31119,N_31157);
and U31400 (N_31400,N_31096,N_31107);
nand U31401 (N_31401,N_31053,N_31188);
nor U31402 (N_31402,N_31184,N_31026);
and U31403 (N_31403,N_31220,N_31114);
and U31404 (N_31404,N_31159,N_31179);
or U31405 (N_31405,N_31027,N_31059);
nor U31406 (N_31406,N_31016,N_31163);
xor U31407 (N_31407,N_31241,N_31083);
nand U31408 (N_31408,N_31234,N_31226);
and U31409 (N_31409,N_31230,N_31006);
xnor U31410 (N_31410,N_31246,N_31141);
or U31411 (N_31411,N_31072,N_31014);
and U31412 (N_31412,N_31143,N_31240);
and U31413 (N_31413,N_31043,N_31093);
or U31414 (N_31414,N_31100,N_31012);
or U31415 (N_31415,N_31078,N_31001);
nor U31416 (N_31416,N_31138,N_31166);
nor U31417 (N_31417,N_31170,N_31152);
or U31418 (N_31418,N_31198,N_31138);
and U31419 (N_31419,N_31128,N_31030);
and U31420 (N_31420,N_31148,N_31235);
nor U31421 (N_31421,N_31236,N_31119);
nor U31422 (N_31422,N_31155,N_31024);
xor U31423 (N_31423,N_31249,N_31115);
nor U31424 (N_31424,N_31061,N_31106);
and U31425 (N_31425,N_31014,N_31118);
or U31426 (N_31426,N_31083,N_31201);
nand U31427 (N_31427,N_31204,N_31018);
xor U31428 (N_31428,N_31051,N_31088);
and U31429 (N_31429,N_31050,N_31209);
nand U31430 (N_31430,N_31169,N_31201);
xor U31431 (N_31431,N_31023,N_31114);
nor U31432 (N_31432,N_31081,N_31079);
and U31433 (N_31433,N_31247,N_31178);
or U31434 (N_31434,N_31053,N_31244);
nor U31435 (N_31435,N_31159,N_31224);
or U31436 (N_31436,N_31215,N_31068);
and U31437 (N_31437,N_31127,N_31183);
nand U31438 (N_31438,N_31181,N_31206);
and U31439 (N_31439,N_31003,N_31017);
or U31440 (N_31440,N_31021,N_31010);
or U31441 (N_31441,N_31107,N_31126);
or U31442 (N_31442,N_31184,N_31040);
xnor U31443 (N_31443,N_31012,N_31149);
nand U31444 (N_31444,N_31244,N_31094);
or U31445 (N_31445,N_31159,N_31231);
xor U31446 (N_31446,N_31115,N_31016);
nor U31447 (N_31447,N_31211,N_31120);
nand U31448 (N_31448,N_31042,N_31032);
xnor U31449 (N_31449,N_31001,N_31221);
or U31450 (N_31450,N_31102,N_31109);
xor U31451 (N_31451,N_31089,N_31198);
nand U31452 (N_31452,N_31060,N_31140);
and U31453 (N_31453,N_31117,N_31171);
nor U31454 (N_31454,N_31232,N_31238);
or U31455 (N_31455,N_31205,N_31133);
nand U31456 (N_31456,N_31225,N_31102);
nand U31457 (N_31457,N_31134,N_31023);
xnor U31458 (N_31458,N_31155,N_31164);
and U31459 (N_31459,N_31091,N_31111);
nor U31460 (N_31460,N_31001,N_31105);
nor U31461 (N_31461,N_31117,N_31037);
nand U31462 (N_31462,N_31005,N_31092);
nand U31463 (N_31463,N_31210,N_31037);
xnor U31464 (N_31464,N_31236,N_31237);
or U31465 (N_31465,N_31138,N_31120);
nand U31466 (N_31466,N_31235,N_31013);
nor U31467 (N_31467,N_31233,N_31073);
or U31468 (N_31468,N_31077,N_31215);
or U31469 (N_31469,N_31034,N_31200);
xor U31470 (N_31470,N_31106,N_31062);
or U31471 (N_31471,N_31187,N_31014);
nor U31472 (N_31472,N_31210,N_31004);
nor U31473 (N_31473,N_31245,N_31062);
nor U31474 (N_31474,N_31120,N_31075);
nor U31475 (N_31475,N_31079,N_31171);
xnor U31476 (N_31476,N_31217,N_31205);
xor U31477 (N_31477,N_31175,N_31059);
or U31478 (N_31478,N_31072,N_31119);
nand U31479 (N_31479,N_31242,N_31210);
nor U31480 (N_31480,N_31160,N_31126);
nand U31481 (N_31481,N_31233,N_31153);
xor U31482 (N_31482,N_31158,N_31083);
nand U31483 (N_31483,N_31239,N_31198);
and U31484 (N_31484,N_31049,N_31095);
or U31485 (N_31485,N_31030,N_31228);
xnor U31486 (N_31486,N_31093,N_31086);
nor U31487 (N_31487,N_31067,N_31197);
nor U31488 (N_31488,N_31011,N_31127);
or U31489 (N_31489,N_31038,N_31236);
or U31490 (N_31490,N_31083,N_31006);
or U31491 (N_31491,N_31033,N_31244);
and U31492 (N_31492,N_31162,N_31022);
xnor U31493 (N_31493,N_31080,N_31093);
nor U31494 (N_31494,N_31112,N_31165);
or U31495 (N_31495,N_31098,N_31177);
and U31496 (N_31496,N_31033,N_31055);
nor U31497 (N_31497,N_31133,N_31196);
xor U31498 (N_31498,N_31055,N_31137);
or U31499 (N_31499,N_31231,N_31230);
or U31500 (N_31500,N_31350,N_31394);
nor U31501 (N_31501,N_31381,N_31438);
or U31502 (N_31502,N_31296,N_31316);
and U31503 (N_31503,N_31386,N_31494);
nand U31504 (N_31504,N_31369,N_31356);
nor U31505 (N_31505,N_31334,N_31304);
nand U31506 (N_31506,N_31366,N_31418);
and U31507 (N_31507,N_31377,N_31413);
xnor U31508 (N_31508,N_31362,N_31491);
or U31509 (N_31509,N_31330,N_31324);
nand U31510 (N_31510,N_31462,N_31393);
nor U31511 (N_31511,N_31463,N_31434);
nor U31512 (N_31512,N_31314,N_31274);
and U31513 (N_31513,N_31308,N_31480);
or U31514 (N_31514,N_31251,N_31301);
and U31515 (N_31515,N_31412,N_31273);
xor U31516 (N_31516,N_31283,N_31429);
and U31517 (N_31517,N_31286,N_31349);
or U31518 (N_31518,N_31470,N_31351);
and U31519 (N_31519,N_31344,N_31489);
nand U31520 (N_31520,N_31469,N_31495);
nand U31521 (N_31521,N_31307,N_31457);
nor U31522 (N_31522,N_31252,N_31257);
nand U31523 (N_31523,N_31454,N_31355);
and U31524 (N_31524,N_31477,N_31395);
or U31525 (N_31525,N_31315,N_31352);
nand U31526 (N_31526,N_31338,N_31289);
and U31527 (N_31527,N_31300,N_31364);
nor U31528 (N_31528,N_31467,N_31426);
nor U31529 (N_31529,N_31335,N_31375);
nor U31530 (N_31530,N_31340,N_31476);
xor U31531 (N_31531,N_31488,N_31253);
nand U31532 (N_31532,N_31409,N_31423);
xnor U31533 (N_31533,N_31416,N_31405);
and U31534 (N_31534,N_31450,N_31396);
or U31535 (N_31535,N_31347,N_31328);
nor U31536 (N_31536,N_31415,N_31460);
or U31537 (N_31537,N_31456,N_31407);
nand U31538 (N_31538,N_31404,N_31442);
nand U31539 (N_31539,N_31378,N_31472);
and U31540 (N_31540,N_31285,N_31400);
and U31541 (N_31541,N_31260,N_31342);
or U31542 (N_31542,N_31422,N_31379);
nor U31543 (N_31543,N_31449,N_31436);
xor U31544 (N_31544,N_31433,N_31365);
nor U31545 (N_31545,N_31266,N_31295);
xor U31546 (N_31546,N_31388,N_31337);
nand U31547 (N_31547,N_31325,N_31496);
or U31548 (N_31548,N_31261,N_31326);
nand U31549 (N_31549,N_31309,N_31398);
xor U31550 (N_31550,N_31411,N_31431);
or U31551 (N_31551,N_31403,N_31255);
and U31552 (N_31552,N_31485,N_31294);
xor U31553 (N_31553,N_31391,N_31414);
nand U31554 (N_31554,N_31376,N_31389);
nor U31555 (N_31555,N_31271,N_31357);
nor U31556 (N_31556,N_31372,N_31320);
nand U31557 (N_31557,N_31451,N_31367);
or U31558 (N_31558,N_31430,N_31440);
nand U31559 (N_31559,N_31331,N_31336);
nand U31560 (N_31560,N_31332,N_31432);
nand U31561 (N_31561,N_31392,N_31466);
nor U31562 (N_31562,N_31464,N_31258);
nand U31563 (N_31563,N_31250,N_31361);
nor U31564 (N_31564,N_31493,N_31427);
and U31565 (N_31565,N_31487,N_31303);
and U31566 (N_31566,N_31406,N_31397);
or U31567 (N_31567,N_31358,N_31475);
nand U31568 (N_31568,N_31482,N_31297);
nor U31569 (N_31569,N_31319,N_31348);
or U31570 (N_31570,N_31302,N_31270);
xor U31571 (N_31571,N_31368,N_31385);
nand U31572 (N_31572,N_31383,N_31390);
nor U31573 (N_31573,N_31317,N_31499);
xnor U31574 (N_31574,N_31321,N_31458);
xor U31575 (N_31575,N_31275,N_31322);
and U31576 (N_31576,N_31447,N_31401);
nand U31577 (N_31577,N_31498,N_31313);
nand U31578 (N_31578,N_31287,N_31473);
or U31579 (N_31579,N_31387,N_31497);
or U31580 (N_31580,N_31419,N_31276);
nor U31581 (N_31581,N_31268,N_31262);
and U31582 (N_31582,N_31323,N_31256);
xor U31583 (N_31583,N_31373,N_31265);
and U31584 (N_31584,N_31492,N_31259);
or U31585 (N_31585,N_31267,N_31382);
or U31586 (N_31586,N_31292,N_31448);
nor U31587 (N_31587,N_31402,N_31481);
nor U31588 (N_31588,N_31479,N_31346);
xnor U31589 (N_31589,N_31474,N_31468);
xor U31590 (N_31590,N_31264,N_31343);
or U31591 (N_31591,N_31465,N_31380);
nand U31592 (N_31592,N_31311,N_31374);
xnor U31593 (N_31593,N_31329,N_31278);
nor U31594 (N_31594,N_31299,N_31437);
and U31595 (N_31595,N_31312,N_31280);
nor U31596 (N_31596,N_31443,N_31439);
nand U31597 (N_31597,N_31370,N_31490);
xnor U31598 (N_31598,N_31445,N_31354);
nand U31599 (N_31599,N_31269,N_31310);
xor U31600 (N_31600,N_31363,N_31327);
nor U31601 (N_31601,N_31288,N_31384);
and U31602 (N_31602,N_31282,N_31399);
xnor U31603 (N_31603,N_31453,N_31444);
or U31604 (N_31604,N_31446,N_31408);
nand U31605 (N_31605,N_31441,N_31435);
or U31606 (N_31606,N_31410,N_31290);
or U31607 (N_31607,N_31371,N_31425);
xor U31608 (N_31608,N_31272,N_31281);
or U31609 (N_31609,N_31478,N_31305);
or U31610 (N_31610,N_31424,N_31291);
and U31611 (N_31611,N_31484,N_31421);
and U31612 (N_31612,N_31298,N_31417);
or U31613 (N_31613,N_31461,N_31345);
or U31614 (N_31614,N_31279,N_31254);
xor U31615 (N_31615,N_31452,N_31306);
or U31616 (N_31616,N_31341,N_31483);
and U31617 (N_31617,N_31359,N_31333);
nand U31618 (N_31618,N_31293,N_31420);
nor U31619 (N_31619,N_31277,N_31263);
nand U31620 (N_31620,N_31318,N_31428);
nor U31621 (N_31621,N_31486,N_31459);
or U31622 (N_31622,N_31471,N_31360);
or U31623 (N_31623,N_31353,N_31284);
and U31624 (N_31624,N_31455,N_31339);
nor U31625 (N_31625,N_31290,N_31430);
nor U31626 (N_31626,N_31498,N_31414);
nand U31627 (N_31627,N_31425,N_31355);
and U31628 (N_31628,N_31361,N_31364);
nand U31629 (N_31629,N_31330,N_31423);
xor U31630 (N_31630,N_31293,N_31274);
or U31631 (N_31631,N_31412,N_31307);
and U31632 (N_31632,N_31457,N_31264);
and U31633 (N_31633,N_31261,N_31256);
or U31634 (N_31634,N_31332,N_31301);
nor U31635 (N_31635,N_31393,N_31333);
or U31636 (N_31636,N_31266,N_31290);
xor U31637 (N_31637,N_31385,N_31459);
nand U31638 (N_31638,N_31415,N_31497);
xnor U31639 (N_31639,N_31385,N_31400);
nor U31640 (N_31640,N_31420,N_31465);
nand U31641 (N_31641,N_31375,N_31381);
nand U31642 (N_31642,N_31313,N_31492);
and U31643 (N_31643,N_31270,N_31463);
and U31644 (N_31644,N_31409,N_31379);
nand U31645 (N_31645,N_31309,N_31353);
nor U31646 (N_31646,N_31374,N_31456);
nand U31647 (N_31647,N_31259,N_31330);
nand U31648 (N_31648,N_31365,N_31477);
or U31649 (N_31649,N_31408,N_31347);
or U31650 (N_31650,N_31273,N_31283);
nand U31651 (N_31651,N_31306,N_31447);
or U31652 (N_31652,N_31295,N_31408);
or U31653 (N_31653,N_31336,N_31297);
nor U31654 (N_31654,N_31390,N_31290);
xnor U31655 (N_31655,N_31466,N_31475);
xnor U31656 (N_31656,N_31467,N_31410);
nand U31657 (N_31657,N_31414,N_31326);
xnor U31658 (N_31658,N_31251,N_31269);
or U31659 (N_31659,N_31426,N_31477);
or U31660 (N_31660,N_31259,N_31357);
nor U31661 (N_31661,N_31302,N_31348);
or U31662 (N_31662,N_31458,N_31491);
nor U31663 (N_31663,N_31265,N_31400);
xor U31664 (N_31664,N_31298,N_31472);
or U31665 (N_31665,N_31320,N_31384);
or U31666 (N_31666,N_31451,N_31492);
nand U31667 (N_31667,N_31269,N_31373);
nor U31668 (N_31668,N_31272,N_31441);
and U31669 (N_31669,N_31349,N_31424);
or U31670 (N_31670,N_31379,N_31493);
and U31671 (N_31671,N_31379,N_31405);
or U31672 (N_31672,N_31489,N_31390);
xnor U31673 (N_31673,N_31413,N_31454);
nand U31674 (N_31674,N_31347,N_31387);
and U31675 (N_31675,N_31378,N_31358);
and U31676 (N_31676,N_31347,N_31377);
or U31677 (N_31677,N_31455,N_31264);
and U31678 (N_31678,N_31452,N_31346);
nand U31679 (N_31679,N_31299,N_31387);
nor U31680 (N_31680,N_31399,N_31273);
and U31681 (N_31681,N_31476,N_31419);
or U31682 (N_31682,N_31285,N_31263);
or U31683 (N_31683,N_31378,N_31479);
xnor U31684 (N_31684,N_31363,N_31277);
nand U31685 (N_31685,N_31446,N_31485);
or U31686 (N_31686,N_31300,N_31317);
or U31687 (N_31687,N_31307,N_31376);
nand U31688 (N_31688,N_31275,N_31369);
nand U31689 (N_31689,N_31442,N_31358);
and U31690 (N_31690,N_31328,N_31318);
nor U31691 (N_31691,N_31251,N_31464);
nand U31692 (N_31692,N_31427,N_31436);
or U31693 (N_31693,N_31477,N_31330);
nor U31694 (N_31694,N_31275,N_31446);
nor U31695 (N_31695,N_31387,N_31394);
nor U31696 (N_31696,N_31314,N_31323);
or U31697 (N_31697,N_31454,N_31280);
nand U31698 (N_31698,N_31444,N_31477);
or U31699 (N_31699,N_31359,N_31433);
and U31700 (N_31700,N_31314,N_31418);
nand U31701 (N_31701,N_31473,N_31354);
nand U31702 (N_31702,N_31385,N_31407);
or U31703 (N_31703,N_31389,N_31407);
or U31704 (N_31704,N_31252,N_31301);
nor U31705 (N_31705,N_31267,N_31416);
xor U31706 (N_31706,N_31446,N_31290);
or U31707 (N_31707,N_31476,N_31472);
or U31708 (N_31708,N_31293,N_31387);
and U31709 (N_31709,N_31282,N_31468);
and U31710 (N_31710,N_31397,N_31282);
nand U31711 (N_31711,N_31455,N_31269);
nor U31712 (N_31712,N_31454,N_31472);
and U31713 (N_31713,N_31261,N_31462);
xnor U31714 (N_31714,N_31332,N_31250);
or U31715 (N_31715,N_31325,N_31386);
nand U31716 (N_31716,N_31467,N_31276);
xnor U31717 (N_31717,N_31326,N_31300);
xnor U31718 (N_31718,N_31368,N_31325);
xor U31719 (N_31719,N_31359,N_31369);
and U31720 (N_31720,N_31261,N_31362);
and U31721 (N_31721,N_31404,N_31371);
nor U31722 (N_31722,N_31355,N_31419);
or U31723 (N_31723,N_31390,N_31494);
and U31724 (N_31724,N_31309,N_31334);
nand U31725 (N_31725,N_31376,N_31354);
nor U31726 (N_31726,N_31255,N_31264);
and U31727 (N_31727,N_31371,N_31458);
nand U31728 (N_31728,N_31447,N_31403);
and U31729 (N_31729,N_31365,N_31383);
or U31730 (N_31730,N_31315,N_31455);
and U31731 (N_31731,N_31377,N_31322);
and U31732 (N_31732,N_31323,N_31456);
nand U31733 (N_31733,N_31277,N_31291);
nand U31734 (N_31734,N_31483,N_31401);
nand U31735 (N_31735,N_31333,N_31286);
nand U31736 (N_31736,N_31371,N_31359);
nor U31737 (N_31737,N_31284,N_31419);
nor U31738 (N_31738,N_31309,N_31451);
xor U31739 (N_31739,N_31408,N_31428);
nand U31740 (N_31740,N_31326,N_31349);
xnor U31741 (N_31741,N_31380,N_31488);
or U31742 (N_31742,N_31341,N_31419);
nand U31743 (N_31743,N_31328,N_31460);
nor U31744 (N_31744,N_31290,N_31419);
xnor U31745 (N_31745,N_31281,N_31313);
and U31746 (N_31746,N_31340,N_31293);
xnor U31747 (N_31747,N_31491,N_31447);
nand U31748 (N_31748,N_31276,N_31485);
or U31749 (N_31749,N_31439,N_31362);
nand U31750 (N_31750,N_31670,N_31687);
nand U31751 (N_31751,N_31700,N_31706);
nor U31752 (N_31752,N_31638,N_31748);
nand U31753 (N_31753,N_31526,N_31552);
nor U31754 (N_31754,N_31690,N_31529);
nor U31755 (N_31755,N_31749,N_31554);
and U31756 (N_31756,N_31738,N_31646);
or U31757 (N_31757,N_31719,N_31740);
xor U31758 (N_31758,N_31657,N_31515);
and U31759 (N_31759,N_31722,N_31715);
or U31760 (N_31760,N_31698,N_31709);
and U31761 (N_31761,N_31602,N_31573);
nor U31762 (N_31762,N_31581,N_31513);
xor U31763 (N_31763,N_31590,N_31630);
nand U31764 (N_31764,N_31626,N_31625);
nand U31765 (N_31765,N_31579,N_31665);
and U31766 (N_31766,N_31596,N_31696);
or U31767 (N_31767,N_31644,N_31619);
or U31768 (N_31768,N_31627,N_31724);
or U31769 (N_31769,N_31673,N_31500);
nor U31770 (N_31770,N_31651,N_31647);
and U31771 (N_31771,N_31659,N_31697);
nor U31772 (N_31772,N_31585,N_31539);
or U31773 (N_31773,N_31588,N_31679);
xor U31774 (N_31774,N_31576,N_31747);
nand U31775 (N_31775,N_31561,N_31654);
and U31776 (N_31776,N_31624,N_31571);
and U31777 (N_31777,N_31595,N_31612);
nor U31778 (N_31778,N_31604,N_31660);
or U31779 (N_31779,N_31721,N_31613);
xnor U31780 (N_31780,N_31556,N_31746);
nor U31781 (N_31781,N_31664,N_31666);
xnor U31782 (N_31782,N_31682,N_31507);
and U31783 (N_31783,N_31582,N_31621);
or U31784 (N_31784,N_31591,N_31508);
nor U31785 (N_31785,N_31531,N_31663);
xnor U31786 (N_31786,N_31536,N_31530);
xnor U31787 (N_31787,N_31684,N_31546);
nor U31788 (N_31788,N_31712,N_31685);
nand U31789 (N_31789,N_31533,N_31667);
nor U31790 (N_31790,N_31708,N_31577);
xnor U31791 (N_31791,N_31528,N_31688);
and U31792 (N_31792,N_31734,N_31723);
nand U31793 (N_31793,N_31538,N_31661);
or U31794 (N_31794,N_31710,N_31523);
or U31795 (N_31795,N_31575,N_31564);
and U31796 (N_31796,N_31689,N_31681);
xor U31797 (N_31797,N_31742,N_31672);
nand U31798 (N_31798,N_31540,N_31695);
nor U31799 (N_31799,N_31677,N_31691);
xnor U31800 (N_31800,N_31675,N_31509);
nand U31801 (N_31801,N_31631,N_31683);
nor U31802 (N_31802,N_31648,N_31645);
xnor U31803 (N_31803,N_31720,N_31519);
or U31804 (N_31804,N_31615,N_31547);
nand U31805 (N_31805,N_31586,N_31545);
or U31806 (N_31806,N_31551,N_31725);
nand U31807 (N_31807,N_31628,N_31521);
nand U31808 (N_31808,N_31518,N_31583);
and U31809 (N_31809,N_31548,N_31668);
and U31810 (N_31810,N_31597,N_31739);
nor U31811 (N_31811,N_31578,N_31587);
xor U31812 (N_31812,N_31732,N_31680);
and U31813 (N_31813,N_31568,N_31733);
xnor U31814 (N_31814,N_31601,N_31557);
xnor U31815 (N_31815,N_31671,N_31729);
or U31816 (N_31816,N_31505,N_31555);
nor U31817 (N_31817,N_31520,N_31705);
nand U31818 (N_31818,N_31510,N_31653);
nor U31819 (N_31819,N_31730,N_31674);
xnor U31820 (N_31820,N_31650,N_31598);
and U31821 (N_31821,N_31504,N_31516);
and U31822 (N_31822,N_31514,N_31714);
nor U31823 (N_31823,N_31692,N_31711);
nor U31824 (N_31824,N_31565,N_31512);
nor U31825 (N_31825,N_31678,N_31594);
or U31826 (N_31826,N_31542,N_31707);
nand U31827 (N_31827,N_31603,N_31580);
or U31828 (N_31828,N_31629,N_31617);
nand U31829 (N_31829,N_31703,N_31537);
or U31830 (N_31830,N_31641,N_31544);
nand U31831 (N_31831,N_31634,N_31570);
and U31832 (N_31832,N_31559,N_31716);
or U31833 (N_31833,N_31676,N_31693);
nand U31834 (N_31834,N_31502,N_31636);
nor U31835 (N_31835,N_31567,N_31614);
and U31836 (N_31836,N_31637,N_31609);
xnor U31837 (N_31837,N_31642,N_31726);
xnor U31838 (N_31838,N_31541,N_31643);
nor U31839 (N_31839,N_31517,N_31592);
xor U31840 (N_31840,N_31702,N_31699);
nor U31841 (N_31841,N_31635,N_31616);
xor U31842 (N_31842,N_31704,N_31600);
nand U31843 (N_31843,N_31735,N_31550);
or U31844 (N_31844,N_31572,N_31607);
and U31845 (N_31845,N_31605,N_31524);
nor U31846 (N_31846,N_31741,N_31562);
and U31847 (N_31847,N_31611,N_31501);
nor U31848 (N_31848,N_31649,N_31543);
nor U31849 (N_31849,N_31569,N_31511);
and U31850 (N_31850,N_31608,N_31694);
xnor U31851 (N_31851,N_31632,N_31652);
xor U31852 (N_31852,N_31610,N_31686);
nand U31853 (N_31853,N_31662,N_31525);
or U31854 (N_31854,N_31633,N_31618);
and U31855 (N_31855,N_31589,N_31655);
nor U31856 (N_31856,N_31745,N_31713);
or U31857 (N_31857,N_31503,N_31669);
nor U31858 (N_31858,N_31506,N_31553);
xor U31859 (N_31859,N_31640,N_31606);
xnor U31860 (N_31860,N_31532,N_31731);
and U31861 (N_31861,N_31743,N_31593);
or U31862 (N_31862,N_31639,N_31584);
nand U31863 (N_31863,N_31737,N_31535);
nand U31864 (N_31864,N_31717,N_31549);
nand U31865 (N_31865,N_31560,N_31522);
and U31866 (N_31866,N_31622,N_31563);
and U31867 (N_31867,N_31566,N_31574);
nand U31868 (N_31868,N_31718,N_31728);
nand U31869 (N_31869,N_31658,N_31527);
nor U31870 (N_31870,N_31744,N_31656);
or U31871 (N_31871,N_31534,N_31736);
and U31872 (N_31872,N_31558,N_31623);
xnor U31873 (N_31873,N_31727,N_31701);
and U31874 (N_31874,N_31620,N_31599);
and U31875 (N_31875,N_31747,N_31676);
nand U31876 (N_31876,N_31609,N_31648);
or U31877 (N_31877,N_31716,N_31686);
and U31878 (N_31878,N_31560,N_31746);
and U31879 (N_31879,N_31742,N_31602);
or U31880 (N_31880,N_31714,N_31737);
nand U31881 (N_31881,N_31670,N_31620);
nor U31882 (N_31882,N_31550,N_31719);
and U31883 (N_31883,N_31680,N_31658);
nand U31884 (N_31884,N_31727,N_31590);
xnor U31885 (N_31885,N_31556,N_31605);
nor U31886 (N_31886,N_31521,N_31676);
or U31887 (N_31887,N_31624,N_31671);
and U31888 (N_31888,N_31513,N_31636);
and U31889 (N_31889,N_31626,N_31662);
nand U31890 (N_31890,N_31669,N_31566);
xnor U31891 (N_31891,N_31745,N_31731);
nand U31892 (N_31892,N_31684,N_31704);
or U31893 (N_31893,N_31703,N_31724);
nor U31894 (N_31894,N_31572,N_31645);
and U31895 (N_31895,N_31515,N_31740);
xnor U31896 (N_31896,N_31563,N_31670);
and U31897 (N_31897,N_31544,N_31601);
nand U31898 (N_31898,N_31669,N_31731);
nor U31899 (N_31899,N_31667,N_31674);
xnor U31900 (N_31900,N_31639,N_31731);
xnor U31901 (N_31901,N_31539,N_31619);
and U31902 (N_31902,N_31676,N_31617);
xor U31903 (N_31903,N_31518,N_31679);
and U31904 (N_31904,N_31668,N_31739);
and U31905 (N_31905,N_31653,N_31575);
nand U31906 (N_31906,N_31638,N_31608);
and U31907 (N_31907,N_31547,N_31599);
and U31908 (N_31908,N_31523,N_31698);
or U31909 (N_31909,N_31702,N_31600);
nand U31910 (N_31910,N_31673,N_31558);
nor U31911 (N_31911,N_31552,N_31744);
nor U31912 (N_31912,N_31628,N_31652);
or U31913 (N_31913,N_31728,N_31687);
and U31914 (N_31914,N_31542,N_31649);
or U31915 (N_31915,N_31536,N_31525);
and U31916 (N_31916,N_31578,N_31696);
xnor U31917 (N_31917,N_31721,N_31740);
xor U31918 (N_31918,N_31645,N_31721);
nor U31919 (N_31919,N_31670,N_31528);
nor U31920 (N_31920,N_31639,N_31628);
and U31921 (N_31921,N_31562,N_31596);
or U31922 (N_31922,N_31644,N_31620);
or U31923 (N_31923,N_31559,N_31604);
or U31924 (N_31924,N_31503,N_31585);
xor U31925 (N_31925,N_31676,N_31551);
xnor U31926 (N_31926,N_31705,N_31669);
and U31927 (N_31927,N_31749,N_31516);
and U31928 (N_31928,N_31580,N_31632);
xor U31929 (N_31929,N_31732,N_31681);
or U31930 (N_31930,N_31688,N_31591);
or U31931 (N_31931,N_31525,N_31694);
and U31932 (N_31932,N_31517,N_31568);
nor U31933 (N_31933,N_31546,N_31703);
xnor U31934 (N_31934,N_31541,N_31581);
xor U31935 (N_31935,N_31534,N_31566);
or U31936 (N_31936,N_31713,N_31663);
nor U31937 (N_31937,N_31652,N_31575);
nor U31938 (N_31938,N_31697,N_31555);
nor U31939 (N_31939,N_31744,N_31714);
nor U31940 (N_31940,N_31514,N_31603);
or U31941 (N_31941,N_31509,N_31590);
nor U31942 (N_31942,N_31643,N_31513);
or U31943 (N_31943,N_31583,N_31635);
xnor U31944 (N_31944,N_31711,N_31559);
nor U31945 (N_31945,N_31660,N_31615);
or U31946 (N_31946,N_31654,N_31707);
or U31947 (N_31947,N_31541,N_31660);
nand U31948 (N_31948,N_31566,N_31594);
nor U31949 (N_31949,N_31561,N_31634);
nor U31950 (N_31950,N_31611,N_31632);
xnor U31951 (N_31951,N_31697,N_31692);
xor U31952 (N_31952,N_31598,N_31728);
and U31953 (N_31953,N_31732,N_31584);
or U31954 (N_31954,N_31534,N_31618);
or U31955 (N_31955,N_31652,N_31570);
nor U31956 (N_31956,N_31555,N_31680);
or U31957 (N_31957,N_31687,N_31550);
xnor U31958 (N_31958,N_31583,N_31500);
nor U31959 (N_31959,N_31719,N_31690);
nand U31960 (N_31960,N_31617,N_31684);
and U31961 (N_31961,N_31559,N_31588);
nor U31962 (N_31962,N_31748,N_31682);
and U31963 (N_31963,N_31652,N_31694);
nor U31964 (N_31964,N_31747,N_31584);
nand U31965 (N_31965,N_31668,N_31552);
nor U31966 (N_31966,N_31608,N_31542);
nand U31967 (N_31967,N_31694,N_31576);
nand U31968 (N_31968,N_31689,N_31647);
nor U31969 (N_31969,N_31713,N_31623);
xnor U31970 (N_31970,N_31629,N_31711);
nand U31971 (N_31971,N_31648,N_31604);
or U31972 (N_31972,N_31742,N_31705);
nor U31973 (N_31973,N_31732,N_31729);
nor U31974 (N_31974,N_31542,N_31505);
nand U31975 (N_31975,N_31672,N_31598);
or U31976 (N_31976,N_31556,N_31747);
nand U31977 (N_31977,N_31527,N_31585);
or U31978 (N_31978,N_31555,N_31514);
and U31979 (N_31979,N_31735,N_31522);
nand U31980 (N_31980,N_31707,N_31680);
or U31981 (N_31981,N_31674,N_31573);
nand U31982 (N_31982,N_31552,N_31698);
nor U31983 (N_31983,N_31589,N_31717);
nor U31984 (N_31984,N_31628,N_31728);
nand U31985 (N_31985,N_31727,N_31711);
or U31986 (N_31986,N_31521,N_31612);
nand U31987 (N_31987,N_31704,N_31691);
or U31988 (N_31988,N_31747,N_31535);
and U31989 (N_31989,N_31713,N_31513);
nand U31990 (N_31990,N_31584,N_31692);
nor U31991 (N_31991,N_31735,N_31630);
or U31992 (N_31992,N_31706,N_31671);
or U31993 (N_31993,N_31749,N_31644);
or U31994 (N_31994,N_31636,N_31647);
nand U31995 (N_31995,N_31673,N_31697);
xor U31996 (N_31996,N_31597,N_31674);
and U31997 (N_31997,N_31652,N_31503);
and U31998 (N_31998,N_31668,N_31625);
or U31999 (N_31999,N_31516,N_31667);
nand U32000 (N_32000,N_31925,N_31883);
or U32001 (N_32001,N_31967,N_31923);
or U32002 (N_32002,N_31830,N_31957);
or U32003 (N_32003,N_31871,N_31993);
and U32004 (N_32004,N_31998,N_31778);
and U32005 (N_32005,N_31906,N_31915);
nor U32006 (N_32006,N_31912,N_31950);
or U32007 (N_32007,N_31935,N_31836);
and U32008 (N_32008,N_31876,N_31838);
xor U32009 (N_32009,N_31844,N_31983);
nand U32010 (N_32010,N_31793,N_31920);
nand U32011 (N_32011,N_31849,N_31779);
nor U32012 (N_32012,N_31914,N_31986);
nand U32013 (N_32013,N_31994,N_31865);
xnor U32014 (N_32014,N_31867,N_31898);
xnor U32015 (N_32015,N_31858,N_31921);
nor U32016 (N_32016,N_31841,N_31803);
nor U32017 (N_32017,N_31929,N_31862);
or U32018 (N_32018,N_31976,N_31826);
and U32019 (N_32019,N_31825,N_31888);
xnor U32020 (N_32020,N_31786,N_31901);
nor U32021 (N_32021,N_31918,N_31872);
nand U32022 (N_32022,N_31981,N_31954);
nand U32023 (N_32023,N_31909,N_31820);
nand U32024 (N_32024,N_31910,N_31751);
and U32025 (N_32025,N_31943,N_31772);
nor U32026 (N_32026,N_31848,N_31958);
and U32027 (N_32027,N_31795,N_31856);
nand U32028 (N_32028,N_31816,N_31972);
xnor U32029 (N_32029,N_31989,N_31752);
nor U32030 (N_32030,N_31970,N_31886);
and U32031 (N_32031,N_31762,N_31866);
nand U32032 (N_32032,N_31938,N_31829);
nand U32033 (N_32033,N_31911,N_31904);
xor U32034 (N_32034,N_31859,N_31975);
nor U32035 (N_32035,N_31968,N_31945);
xor U32036 (N_32036,N_31894,N_31895);
nand U32037 (N_32037,N_31817,N_31837);
and U32038 (N_32038,N_31870,N_31878);
nand U32039 (N_32039,N_31979,N_31831);
and U32040 (N_32040,N_31775,N_31771);
and U32041 (N_32041,N_31790,N_31916);
xnor U32042 (N_32042,N_31939,N_31833);
and U32043 (N_32043,N_31812,N_31947);
or U32044 (N_32044,N_31889,N_31763);
xnor U32045 (N_32045,N_31982,N_31757);
nand U32046 (N_32046,N_31917,N_31791);
xor U32047 (N_32047,N_31965,N_31990);
xor U32048 (N_32048,N_31861,N_31864);
or U32049 (N_32049,N_31783,N_31900);
xor U32050 (N_32050,N_31884,N_31896);
nand U32051 (N_32051,N_31755,N_31835);
and U32052 (N_32052,N_31818,N_31934);
nor U32053 (N_32053,N_31960,N_31801);
nor U32054 (N_32054,N_31953,N_31873);
nand U32055 (N_32055,N_31810,N_31774);
nor U32056 (N_32056,N_31773,N_31956);
nor U32057 (N_32057,N_31897,N_31766);
and U32058 (N_32058,N_31842,N_31987);
and U32059 (N_32059,N_31787,N_31794);
or U32060 (N_32060,N_31834,N_31991);
nor U32061 (N_32061,N_31776,N_31941);
xor U32062 (N_32062,N_31902,N_31819);
nor U32063 (N_32063,N_31931,N_31892);
nor U32064 (N_32064,N_31875,N_31891);
xor U32065 (N_32065,N_31937,N_31824);
nor U32066 (N_32066,N_31952,N_31913);
nor U32067 (N_32067,N_31797,N_31928);
nand U32068 (N_32068,N_31893,N_31823);
xnor U32069 (N_32069,N_31759,N_31764);
xor U32070 (N_32070,N_31985,N_31854);
xor U32071 (N_32071,N_31940,N_31782);
xor U32072 (N_32072,N_31851,N_31868);
nor U32073 (N_32073,N_31890,N_31846);
and U32074 (N_32074,N_31805,N_31959);
or U32075 (N_32075,N_31997,N_31984);
xnor U32076 (N_32076,N_31908,N_31814);
and U32077 (N_32077,N_31857,N_31996);
nand U32078 (N_32078,N_31758,N_31840);
and U32079 (N_32079,N_31977,N_31880);
and U32080 (N_32080,N_31750,N_31944);
or U32081 (N_32081,N_31964,N_31753);
nor U32082 (N_32082,N_31922,N_31808);
nand U32083 (N_32083,N_31788,N_31770);
and U32084 (N_32084,N_31999,N_31877);
xor U32085 (N_32085,N_31863,N_31926);
nand U32086 (N_32086,N_31980,N_31828);
or U32087 (N_32087,N_31827,N_31806);
xor U32088 (N_32088,N_31882,N_31881);
and U32089 (N_32089,N_31885,N_31804);
nand U32090 (N_32090,N_31860,N_31955);
and U32091 (N_32091,N_31839,N_31936);
or U32092 (N_32092,N_31754,N_31978);
xnor U32093 (N_32093,N_31815,N_31777);
xor U32094 (N_32094,N_31781,N_31949);
nand U32095 (N_32095,N_31822,N_31948);
nand U32096 (N_32096,N_31850,N_31927);
and U32097 (N_32097,N_31756,N_31799);
nor U32098 (N_32098,N_31951,N_31887);
nor U32099 (N_32099,N_31800,N_31852);
xnor U32100 (N_32100,N_31899,N_31855);
and U32101 (N_32101,N_31761,N_31768);
nor U32102 (N_32102,N_31845,N_31907);
nand U32103 (N_32103,N_31802,N_31813);
and U32104 (N_32104,N_31946,N_31847);
nand U32105 (N_32105,N_31853,N_31780);
or U32106 (N_32106,N_31821,N_31843);
xnor U32107 (N_32107,N_31789,N_31879);
or U32108 (N_32108,N_31785,N_31760);
nor U32109 (N_32109,N_31942,N_31807);
nor U32110 (N_32110,N_31903,N_31796);
and U32111 (N_32111,N_31784,N_31930);
or U32112 (N_32112,N_31905,N_31966);
xor U32113 (N_32113,N_31963,N_31962);
nor U32114 (N_32114,N_31995,N_31961);
or U32115 (N_32115,N_31874,N_31932);
or U32116 (N_32116,N_31924,N_31767);
xor U32117 (N_32117,N_31992,N_31809);
nand U32118 (N_32118,N_31974,N_31919);
and U32119 (N_32119,N_31969,N_31988);
nor U32120 (N_32120,N_31973,N_31769);
or U32121 (N_32121,N_31933,N_31792);
nor U32122 (N_32122,N_31798,N_31832);
nor U32123 (N_32123,N_31765,N_31811);
xor U32124 (N_32124,N_31971,N_31869);
and U32125 (N_32125,N_31869,N_31801);
nand U32126 (N_32126,N_31957,N_31867);
nor U32127 (N_32127,N_31751,N_31761);
or U32128 (N_32128,N_31904,N_31898);
nor U32129 (N_32129,N_31773,N_31867);
nor U32130 (N_32130,N_31992,N_31781);
xor U32131 (N_32131,N_31841,N_31926);
or U32132 (N_32132,N_31882,N_31924);
and U32133 (N_32133,N_31858,N_31909);
or U32134 (N_32134,N_31966,N_31798);
nand U32135 (N_32135,N_31929,N_31964);
and U32136 (N_32136,N_31972,N_31770);
nand U32137 (N_32137,N_31972,N_31771);
and U32138 (N_32138,N_31992,N_31824);
and U32139 (N_32139,N_31870,N_31993);
nor U32140 (N_32140,N_31869,N_31929);
nand U32141 (N_32141,N_31759,N_31951);
or U32142 (N_32142,N_31768,N_31931);
nand U32143 (N_32143,N_31866,N_31950);
nor U32144 (N_32144,N_31881,N_31801);
xnor U32145 (N_32145,N_31806,N_31894);
nor U32146 (N_32146,N_31828,N_31998);
and U32147 (N_32147,N_31931,N_31928);
nand U32148 (N_32148,N_31866,N_31862);
and U32149 (N_32149,N_31994,N_31812);
and U32150 (N_32150,N_31773,N_31975);
and U32151 (N_32151,N_31785,N_31995);
nor U32152 (N_32152,N_31808,N_31952);
and U32153 (N_32153,N_31928,N_31872);
nand U32154 (N_32154,N_31754,N_31993);
or U32155 (N_32155,N_31760,N_31987);
nand U32156 (N_32156,N_31959,N_31750);
xnor U32157 (N_32157,N_31811,N_31809);
and U32158 (N_32158,N_31932,N_31860);
nor U32159 (N_32159,N_31811,N_31980);
xnor U32160 (N_32160,N_31840,N_31989);
and U32161 (N_32161,N_31930,N_31926);
nor U32162 (N_32162,N_31808,N_31836);
xor U32163 (N_32163,N_31991,N_31762);
nor U32164 (N_32164,N_31881,N_31789);
nand U32165 (N_32165,N_31856,N_31814);
xnor U32166 (N_32166,N_31815,N_31837);
xor U32167 (N_32167,N_31885,N_31925);
xnor U32168 (N_32168,N_31826,N_31919);
nand U32169 (N_32169,N_31884,N_31961);
nor U32170 (N_32170,N_31914,N_31765);
nand U32171 (N_32171,N_31819,N_31876);
and U32172 (N_32172,N_31989,N_31803);
or U32173 (N_32173,N_31980,N_31943);
xnor U32174 (N_32174,N_31811,N_31986);
nor U32175 (N_32175,N_31994,N_31953);
nand U32176 (N_32176,N_31872,N_31884);
and U32177 (N_32177,N_31776,N_31841);
or U32178 (N_32178,N_31880,N_31960);
xnor U32179 (N_32179,N_31866,N_31996);
xnor U32180 (N_32180,N_31956,N_31913);
nand U32181 (N_32181,N_31968,N_31985);
nand U32182 (N_32182,N_31914,N_31853);
nand U32183 (N_32183,N_31916,N_31922);
and U32184 (N_32184,N_31904,N_31774);
nand U32185 (N_32185,N_31931,N_31866);
nor U32186 (N_32186,N_31971,N_31834);
nand U32187 (N_32187,N_31907,N_31840);
and U32188 (N_32188,N_31988,N_31853);
and U32189 (N_32189,N_31851,N_31908);
or U32190 (N_32190,N_31815,N_31981);
or U32191 (N_32191,N_31779,N_31851);
nor U32192 (N_32192,N_31792,N_31784);
xnor U32193 (N_32193,N_31778,N_31812);
xor U32194 (N_32194,N_31982,N_31961);
nor U32195 (N_32195,N_31845,N_31750);
or U32196 (N_32196,N_31966,N_31984);
xnor U32197 (N_32197,N_31992,N_31880);
and U32198 (N_32198,N_31813,N_31757);
or U32199 (N_32199,N_31904,N_31978);
nand U32200 (N_32200,N_31765,N_31918);
xnor U32201 (N_32201,N_31884,N_31873);
nor U32202 (N_32202,N_31966,N_31982);
and U32203 (N_32203,N_31786,N_31915);
nand U32204 (N_32204,N_31827,N_31905);
or U32205 (N_32205,N_31840,N_31902);
or U32206 (N_32206,N_31985,N_31976);
nor U32207 (N_32207,N_31907,N_31966);
nor U32208 (N_32208,N_31879,N_31880);
xor U32209 (N_32209,N_31966,N_31954);
nand U32210 (N_32210,N_31929,N_31791);
nand U32211 (N_32211,N_31988,N_31881);
or U32212 (N_32212,N_31846,N_31896);
nand U32213 (N_32213,N_31830,N_31780);
nand U32214 (N_32214,N_31979,N_31937);
xnor U32215 (N_32215,N_31967,N_31997);
nand U32216 (N_32216,N_31877,N_31931);
and U32217 (N_32217,N_31959,N_31865);
xor U32218 (N_32218,N_31869,N_31757);
and U32219 (N_32219,N_31970,N_31878);
or U32220 (N_32220,N_31849,N_31981);
nor U32221 (N_32221,N_31937,N_31968);
xnor U32222 (N_32222,N_31845,N_31935);
xor U32223 (N_32223,N_31936,N_31762);
or U32224 (N_32224,N_31792,N_31929);
or U32225 (N_32225,N_31971,N_31863);
or U32226 (N_32226,N_31899,N_31883);
or U32227 (N_32227,N_31815,N_31798);
nor U32228 (N_32228,N_31906,N_31952);
xnor U32229 (N_32229,N_31821,N_31872);
xor U32230 (N_32230,N_31760,N_31850);
and U32231 (N_32231,N_31796,N_31794);
and U32232 (N_32232,N_31994,N_31974);
and U32233 (N_32233,N_31826,N_31892);
or U32234 (N_32234,N_31762,N_31893);
xor U32235 (N_32235,N_31751,N_31898);
or U32236 (N_32236,N_31990,N_31830);
or U32237 (N_32237,N_31979,N_31847);
or U32238 (N_32238,N_31762,N_31945);
nor U32239 (N_32239,N_31772,N_31917);
xor U32240 (N_32240,N_31841,N_31851);
xnor U32241 (N_32241,N_31915,N_31789);
or U32242 (N_32242,N_31903,N_31832);
and U32243 (N_32243,N_31849,N_31830);
nand U32244 (N_32244,N_31809,N_31947);
nor U32245 (N_32245,N_31943,N_31782);
or U32246 (N_32246,N_31907,N_31922);
nand U32247 (N_32247,N_31924,N_31929);
and U32248 (N_32248,N_31828,N_31899);
nand U32249 (N_32249,N_31765,N_31857);
and U32250 (N_32250,N_32076,N_32113);
nand U32251 (N_32251,N_32009,N_32146);
xor U32252 (N_32252,N_32137,N_32246);
and U32253 (N_32253,N_32139,N_32169);
or U32254 (N_32254,N_32235,N_32188);
xor U32255 (N_32255,N_32104,N_32056);
xnor U32256 (N_32256,N_32021,N_32239);
xnor U32257 (N_32257,N_32058,N_32130);
or U32258 (N_32258,N_32236,N_32230);
xor U32259 (N_32259,N_32055,N_32197);
nor U32260 (N_32260,N_32196,N_32073);
or U32261 (N_32261,N_32211,N_32098);
xor U32262 (N_32262,N_32013,N_32042);
nand U32263 (N_32263,N_32161,N_32063);
or U32264 (N_32264,N_32031,N_32008);
or U32265 (N_32265,N_32208,N_32233);
and U32266 (N_32266,N_32140,N_32005);
nand U32267 (N_32267,N_32043,N_32052);
or U32268 (N_32268,N_32238,N_32154);
nor U32269 (N_32269,N_32229,N_32074);
xor U32270 (N_32270,N_32184,N_32177);
or U32271 (N_32271,N_32114,N_32051);
nor U32272 (N_32272,N_32214,N_32151);
nor U32273 (N_32273,N_32090,N_32062);
nor U32274 (N_32274,N_32147,N_32125);
or U32275 (N_32275,N_32133,N_32115);
xor U32276 (N_32276,N_32038,N_32200);
nor U32277 (N_32277,N_32245,N_32007);
xor U32278 (N_32278,N_32057,N_32045);
or U32279 (N_32279,N_32105,N_32195);
and U32280 (N_32280,N_32120,N_32150);
nand U32281 (N_32281,N_32136,N_32217);
or U32282 (N_32282,N_32095,N_32143);
or U32283 (N_32283,N_32092,N_32180);
nand U32284 (N_32284,N_32059,N_32163);
or U32285 (N_32285,N_32141,N_32039);
xor U32286 (N_32286,N_32025,N_32019);
xnor U32287 (N_32287,N_32131,N_32102);
or U32288 (N_32288,N_32036,N_32249);
and U32289 (N_32289,N_32152,N_32018);
or U32290 (N_32290,N_32165,N_32089);
xor U32291 (N_32291,N_32030,N_32190);
xor U32292 (N_32292,N_32004,N_32168);
nor U32293 (N_32293,N_32223,N_32127);
and U32294 (N_32294,N_32047,N_32103);
nand U32295 (N_32295,N_32212,N_32119);
and U32296 (N_32296,N_32162,N_32198);
or U32297 (N_32297,N_32240,N_32170);
nor U32298 (N_32298,N_32017,N_32040);
or U32299 (N_32299,N_32110,N_32189);
and U32300 (N_32300,N_32209,N_32087);
nor U32301 (N_32301,N_32012,N_32156);
xnor U32302 (N_32302,N_32153,N_32122);
nand U32303 (N_32303,N_32175,N_32194);
nor U32304 (N_32304,N_32167,N_32086);
nand U32305 (N_32305,N_32145,N_32160);
or U32306 (N_32306,N_32015,N_32049);
and U32307 (N_32307,N_32024,N_32046);
nand U32308 (N_32308,N_32106,N_32203);
xor U32309 (N_32309,N_32075,N_32080);
and U32310 (N_32310,N_32226,N_32243);
xor U32311 (N_32311,N_32002,N_32044);
nor U32312 (N_32312,N_32069,N_32037);
and U32313 (N_32313,N_32020,N_32187);
nand U32314 (N_32314,N_32201,N_32096);
nor U32315 (N_32315,N_32222,N_32082);
nor U32316 (N_32316,N_32224,N_32183);
and U32317 (N_32317,N_32228,N_32128);
or U32318 (N_32318,N_32091,N_32001);
and U32319 (N_32319,N_32084,N_32027);
and U32320 (N_32320,N_32132,N_32033);
and U32321 (N_32321,N_32023,N_32181);
nor U32322 (N_32322,N_32179,N_32094);
or U32323 (N_32323,N_32107,N_32078);
nor U32324 (N_32324,N_32101,N_32210);
and U32325 (N_32325,N_32144,N_32193);
and U32326 (N_32326,N_32158,N_32121);
nand U32327 (N_32327,N_32173,N_32010);
or U32328 (N_32328,N_32241,N_32157);
or U32329 (N_32329,N_32166,N_32220);
nand U32330 (N_32330,N_32244,N_32232);
xor U32331 (N_32331,N_32081,N_32029);
nand U32332 (N_32332,N_32138,N_32108);
and U32333 (N_32333,N_32206,N_32050);
xnor U32334 (N_32334,N_32109,N_32221);
or U32335 (N_32335,N_32186,N_32202);
nand U32336 (N_32336,N_32159,N_32155);
and U32337 (N_32337,N_32142,N_32085);
or U32338 (N_32338,N_32060,N_32213);
nand U32339 (N_32339,N_32053,N_32248);
nor U32340 (N_32340,N_32215,N_32124);
nand U32341 (N_32341,N_32216,N_32117);
and U32342 (N_32342,N_32192,N_32099);
xor U32343 (N_32343,N_32247,N_32205);
or U32344 (N_32344,N_32219,N_32032);
xor U32345 (N_32345,N_32067,N_32207);
nand U32346 (N_32346,N_32199,N_32176);
nor U32347 (N_32347,N_32185,N_32225);
nor U32348 (N_32348,N_32077,N_32171);
nor U32349 (N_32349,N_32148,N_32054);
and U32350 (N_32350,N_32227,N_32000);
xor U32351 (N_32351,N_32079,N_32164);
nand U32352 (N_32352,N_32234,N_32178);
and U32353 (N_32353,N_32231,N_32118);
xor U32354 (N_32354,N_32237,N_32068);
xnor U32355 (N_32355,N_32026,N_32061);
xnor U32356 (N_32356,N_32172,N_32116);
xor U32357 (N_32357,N_32071,N_32126);
or U32358 (N_32358,N_32135,N_32097);
or U32359 (N_32359,N_32011,N_32112);
or U32360 (N_32360,N_32083,N_32093);
and U32361 (N_32361,N_32048,N_32072);
nand U32362 (N_32362,N_32100,N_32066);
nor U32363 (N_32363,N_32204,N_32123);
nand U32364 (N_32364,N_32014,N_32003);
or U32365 (N_32365,N_32028,N_32088);
or U32366 (N_32366,N_32035,N_32022);
nand U32367 (N_32367,N_32191,N_32129);
nand U32368 (N_32368,N_32218,N_32182);
nand U32369 (N_32369,N_32065,N_32006);
nor U32370 (N_32370,N_32041,N_32149);
nand U32371 (N_32371,N_32174,N_32070);
nor U32372 (N_32372,N_32016,N_32034);
nor U32373 (N_32373,N_32111,N_32134);
nand U32374 (N_32374,N_32242,N_32064);
xnor U32375 (N_32375,N_32001,N_32079);
xor U32376 (N_32376,N_32176,N_32107);
or U32377 (N_32377,N_32189,N_32206);
and U32378 (N_32378,N_32165,N_32144);
or U32379 (N_32379,N_32243,N_32115);
nor U32380 (N_32380,N_32171,N_32154);
nor U32381 (N_32381,N_32046,N_32136);
nor U32382 (N_32382,N_32010,N_32136);
or U32383 (N_32383,N_32144,N_32099);
and U32384 (N_32384,N_32074,N_32039);
nand U32385 (N_32385,N_32225,N_32017);
and U32386 (N_32386,N_32057,N_32085);
xor U32387 (N_32387,N_32098,N_32014);
and U32388 (N_32388,N_32082,N_32181);
and U32389 (N_32389,N_32002,N_32109);
xnor U32390 (N_32390,N_32107,N_32123);
xor U32391 (N_32391,N_32174,N_32020);
nand U32392 (N_32392,N_32043,N_32139);
xnor U32393 (N_32393,N_32121,N_32084);
and U32394 (N_32394,N_32155,N_32072);
nor U32395 (N_32395,N_32028,N_32084);
and U32396 (N_32396,N_32004,N_32011);
nor U32397 (N_32397,N_32186,N_32114);
nor U32398 (N_32398,N_32140,N_32063);
and U32399 (N_32399,N_32215,N_32052);
and U32400 (N_32400,N_32059,N_32151);
nand U32401 (N_32401,N_32005,N_32046);
nand U32402 (N_32402,N_32114,N_32011);
and U32403 (N_32403,N_32065,N_32191);
and U32404 (N_32404,N_32086,N_32087);
or U32405 (N_32405,N_32146,N_32134);
nand U32406 (N_32406,N_32077,N_32225);
nand U32407 (N_32407,N_32070,N_32045);
or U32408 (N_32408,N_32023,N_32006);
and U32409 (N_32409,N_32188,N_32093);
nand U32410 (N_32410,N_32175,N_32243);
or U32411 (N_32411,N_32048,N_32028);
nand U32412 (N_32412,N_32225,N_32164);
nand U32413 (N_32413,N_32200,N_32176);
nor U32414 (N_32414,N_32065,N_32098);
nor U32415 (N_32415,N_32103,N_32089);
or U32416 (N_32416,N_32105,N_32055);
nor U32417 (N_32417,N_32081,N_32200);
xnor U32418 (N_32418,N_32083,N_32022);
nor U32419 (N_32419,N_32034,N_32174);
xor U32420 (N_32420,N_32244,N_32201);
and U32421 (N_32421,N_32034,N_32131);
nand U32422 (N_32422,N_32196,N_32229);
and U32423 (N_32423,N_32136,N_32224);
or U32424 (N_32424,N_32079,N_32152);
and U32425 (N_32425,N_32046,N_32249);
or U32426 (N_32426,N_32091,N_32179);
nand U32427 (N_32427,N_32008,N_32073);
xor U32428 (N_32428,N_32239,N_32174);
xor U32429 (N_32429,N_32097,N_32022);
and U32430 (N_32430,N_32041,N_32179);
nor U32431 (N_32431,N_32183,N_32082);
and U32432 (N_32432,N_32050,N_32019);
nor U32433 (N_32433,N_32003,N_32157);
or U32434 (N_32434,N_32098,N_32125);
and U32435 (N_32435,N_32100,N_32009);
xor U32436 (N_32436,N_32070,N_32098);
and U32437 (N_32437,N_32142,N_32239);
xor U32438 (N_32438,N_32071,N_32244);
nor U32439 (N_32439,N_32155,N_32065);
nand U32440 (N_32440,N_32184,N_32161);
nand U32441 (N_32441,N_32096,N_32237);
xor U32442 (N_32442,N_32222,N_32149);
or U32443 (N_32443,N_32062,N_32068);
nand U32444 (N_32444,N_32082,N_32000);
nand U32445 (N_32445,N_32043,N_32058);
nor U32446 (N_32446,N_32039,N_32138);
xnor U32447 (N_32447,N_32166,N_32198);
or U32448 (N_32448,N_32220,N_32202);
nor U32449 (N_32449,N_32222,N_32189);
or U32450 (N_32450,N_32183,N_32213);
xnor U32451 (N_32451,N_32063,N_32164);
xnor U32452 (N_32452,N_32098,N_32081);
nor U32453 (N_32453,N_32182,N_32206);
nand U32454 (N_32454,N_32009,N_32139);
nand U32455 (N_32455,N_32247,N_32075);
and U32456 (N_32456,N_32127,N_32035);
nand U32457 (N_32457,N_32230,N_32118);
nor U32458 (N_32458,N_32107,N_32040);
nor U32459 (N_32459,N_32007,N_32071);
xnor U32460 (N_32460,N_32074,N_32214);
and U32461 (N_32461,N_32242,N_32067);
or U32462 (N_32462,N_32185,N_32028);
xnor U32463 (N_32463,N_32132,N_32240);
or U32464 (N_32464,N_32141,N_32208);
xnor U32465 (N_32465,N_32105,N_32109);
or U32466 (N_32466,N_32228,N_32206);
nand U32467 (N_32467,N_32028,N_32068);
nand U32468 (N_32468,N_32049,N_32119);
nand U32469 (N_32469,N_32053,N_32127);
nor U32470 (N_32470,N_32167,N_32229);
or U32471 (N_32471,N_32133,N_32101);
or U32472 (N_32472,N_32223,N_32154);
nand U32473 (N_32473,N_32106,N_32082);
xor U32474 (N_32474,N_32162,N_32201);
nand U32475 (N_32475,N_32242,N_32205);
xor U32476 (N_32476,N_32199,N_32003);
nand U32477 (N_32477,N_32032,N_32221);
xor U32478 (N_32478,N_32095,N_32038);
and U32479 (N_32479,N_32014,N_32234);
nand U32480 (N_32480,N_32169,N_32231);
and U32481 (N_32481,N_32004,N_32083);
nor U32482 (N_32482,N_32044,N_32049);
nand U32483 (N_32483,N_32015,N_32120);
xnor U32484 (N_32484,N_32168,N_32244);
or U32485 (N_32485,N_32093,N_32068);
nand U32486 (N_32486,N_32242,N_32211);
and U32487 (N_32487,N_32198,N_32183);
xnor U32488 (N_32488,N_32142,N_32039);
or U32489 (N_32489,N_32145,N_32030);
nor U32490 (N_32490,N_32073,N_32149);
and U32491 (N_32491,N_32214,N_32179);
xor U32492 (N_32492,N_32033,N_32239);
or U32493 (N_32493,N_32116,N_32058);
and U32494 (N_32494,N_32093,N_32131);
and U32495 (N_32495,N_32135,N_32224);
xnor U32496 (N_32496,N_32213,N_32021);
nand U32497 (N_32497,N_32107,N_32243);
and U32498 (N_32498,N_32113,N_32152);
xnor U32499 (N_32499,N_32016,N_32133);
or U32500 (N_32500,N_32430,N_32445);
and U32501 (N_32501,N_32400,N_32362);
xnor U32502 (N_32502,N_32332,N_32357);
and U32503 (N_32503,N_32365,N_32410);
xor U32504 (N_32504,N_32315,N_32294);
or U32505 (N_32505,N_32419,N_32301);
nor U32506 (N_32506,N_32428,N_32311);
nand U32507 (N_32507,N_32436,N_32469);
or U32508 (N_32508,N_32392,N_32429);
nor U32509 (N_32509,N_32285,N_32406);
xor U32510 (N_32510,N_32342,N_32283);
and U32511 (N_32511,N_32328,N_32461);
xnor U32512 (N_32512,N_32325,N_32456);
and U32513 (N_32513,N_32355,N_32420);
and U32514 (N_32514,N_32390,N_32281);
nand U32515 (N_32515,N_32286,N_32309);
and U32516 (N_32516,N_32348,N_32273);
nand U32517 (N_32517,N_32438,N_32297);
nand U32518 (N_32518,N_32450,N_32389);
xnor U32519 (N_32519,N_32405,N_32466);
nand U32520 (N_32520,N_32270,N_32495);
nor U32521 (N_32521,N_32434,N_32326);
and U32522 (N_32522,N_32352,N_32278);
xor U32523 (N_32523,N_32289,N_32319);
nor U32524 (N_32524,N_32486,N_32378);
or U32525 (N_32525,N_32475,N_32300);
and U32526 (N_32526,N_32255,N_32314);
nor U32527 (N_32527,N_32320,N_32358);
or U32528 (N_32528,N_32498,N_32393);
nor U32529 (N_32529,N_32418,N_32427);
xor U32530 (N_32530,N_32367,N_32318);
xor U32531 (N_32531,N_32472,N_32423);
or U32532 (N_32532,N_32383,N_32499);
nor U32533 (N_32533,N_32312,N_32329);
xor U32534 (N_32534,N_32492,N_32464);
or U32535 (N_32535,N_32402,N_32449);
and U32536 (N_32536,N_32261,N_32265);
xor U32537 (N_32537,N_32432,N_32408);
xor U32538 (N_32538,N_32396,N_32287);
xor U32539 (N_32539,N_32439,N_32368);
xor U32540 (N_32540,N_32340,N_32424);
xor U32541 (N_32541,N_32480,N_32431);
nand U32542 (N_32542,N_32394,N_32307);
or U32543 (N_32543,N_32447,N_32382);
and U32544 (N_32544,N_32391,N_32381);
or U32545 (N_32545,N_32483,N_32361);
xor U32546 (N_32546,N_32359,N_32440);
and U32547 (N_32547,N_32284,N_32413);
and U32548 (N_32548,N_32275,N_32346);
nor U32549 (N_32549,N_32337,N_32462);
or U32550 (N_32550,N_32448,N_32298);
and U32551 (N_32551,N_32372,N_32327);
nor U32552 (N_32552,N_32330,N_32454);
and U32553 (N_32553,N_32259,N_32268);
and U32554 (N_32554,N_32334,N_32313);
or U32555 (N_32555,N_32292,N_32351);
xnor U32556 (N_32556,N_32282,N_32258);
or U32557 (N_32557,N_32338,N_32460);
or U32558 (N_32558,N_32415,N_32349);
and U32559 (N_32559,N_32433,N_32344);
or U32560 (N_32560,N_32291,N_32366);
xor U32561 (N_32561,N_32435,N_32279);
and U32562 (N_32562,N_32478,N_32463);
and U32563 (N_32563,N_32306,N_32474);
or U32564 (N_32564,N_32395,N_32290);
xnor U32565 (N_32565,N_32274,N_32266);
xnor U32566 (N_32566,N_32250,N_32253);
and U32567 (N_32567,N_32323,N_32467);
nand U32568 (N_32568,N_32386,N_32437);
or U32569 (N_32569,N_32263,N_32387);
nor U32570 (N_32570,N_32335,N_32321);
and U32571 (N_32571,N_32267,N_32451);
nor U32572 (N_32572,N_32452,N_32401);
nand U32573 (N_32573,N_32426,N_32444);
nor U32574 (N_32574,N_32488,N_32399);
nand U32575 (N_32575,N_32299,N_32446);
xor U32576 (N_32576,N_32494,N_32497);
or U32577 (N_32577,N_32404,N_32331);
or U32578 (N_32578,N_32341,N_32468);
and U32579 (N_32579,N_32479,N_32398);
xnor U32580 (N_32580,N_32354,N_32345);
nand U32581 (N_32581,N_32373,N_32257);
xor U32582 (N_32582,N_32407,N_32384);
or U32583 (N_32583,N_32293,N_32316);
nand U32584 (N_32584,N_32322,N_32484);
and U32585 (N_32585,N_32277,N_32455);
nor U32586 (N_32586,N_32397,N_32379);
or U32587 (N_32587,N_32443,N_32371);
xor U32588 (N_32588,N_32347,N_32416);
nor U32589 (N_32589,N_32324,N_32271);
and U32590 (N_32590,N_32276,N_32308);
or U32591 (N_32591,N_32376,N_32262);
nand U32592 (N_32592,N_32411,N_32356);
nor U32593 (N_32593,N_32256,N_32487);
and U32594 (N_32594,N_32491,N_32490);
nor U32595 (N_32595,N_32333,N_32305);
and U32596 (N_32596,N_32377,N_32441);
nand U32597 (N_32597,N_32473,N_32374);
and U32598 (N_32598,N_32370,N_32272);
nor U32599 (N_32599,N_32388,N_32310);
nand U32600 (N_32600,N_32482,N_32425);
or U32601 (N_32601,N_32254,N_32459);
or U32602 (N_32602,N_32422,N_32295);
or U32603 (N_32603,N_32360,N_32264);
nor U32604 (N_32604,N_32412,N_32260);
or U32605 (N_32605,N_32252,N_32477);
and U32606 (N_32606,N_32414,N_32403);
nor U32607 (N_32607,N_32476,N_32269);
nor U32608 (N_32608,N_32465,N_32288);
or U32609 (N_32609,N_32303,N_32280);
nor U32610 (N_32610,N_32363,N_32409);
nor U32611 (N_32611,N_32302,N_32489);
or U32612 (N_32612,N_32481,N_32421);
and U32613 (N_32613,N_32317,N_32417);
and U32614 (N_32614,N_32485,N_32458);
xnor U32615 (N_32615,N_32493,N_32380);
nand U32616 (N_32616,N_32350,N_32369);
nand U32617 (N_32617,N_32457,N_32470);
and U32618 (N_32618,N_32251,N_32385);
xor U32619 (N_32619,N_32336,N_32375);
xnor U32620 (N_32620,N_32364,N_32343);
nor U32621 (N_32621,N_32296,N_32339);
nand U32622 (N_32622,N_32471,N_32453);
and U32623 (N_32623,N_32442,N_32496);
xnor U32624 (N_32624,N_32304,N_32353);
or U32625 (N_32625,N_32491,N_32416);
nand U32626 (N_32626,N_32333,N_32440);
nand U32627 (N_32627,N_32375,N_32382);
nand U32628 (N_32628,N_32438,N_32349);
or U32629 (N_32629,N_32271,N_32274);
xnor U32630 (N_32630,N_32360,N_32280);
nand U32631 (N_32631,N_32484,N_32381);
or U32632 (N_32632,N_32254,N_32347);
nor U32633 (N_32633,N_32418,N_32470);
nand U32634 (N_32634,N_32367,N_32415);
or U32635 (N_32635,N_32485,N_32347);
nand U32636 (N_32636,N_32341,N_32302);
and U32637 (N_32637,N_32318,N_32317);
xor U32638 (N_32638,N_32320,N_32428);
or U32639 (N_32639,N_32343,N_32290);
nand U32640 (N_32640,N_32287,N_32353);
nor U32641 (N_32641,N_32391,N_32267);
nor U32642 (N_32642,N_32495,N_32367);
nor U32643 (N_32643,N_32492,N_32393);
and U32644 (N_32644,N_32483,N_32323);
nor U32645 (N_32645,N_32466,N_32302);
xnor U32646 (N_32646,N_32448,N_32369);
and U32647 (N_32647,N_32420,N_32252);
or U32648 (N_32648,N_32440,N_32413);
nand U32649 (N_32649,N_32325,N_32471);
or U32650 (N_32650,N_32360,N_32294);
and U32651 (N_32651,N_32397,N_32304);
nor U32652 (N_32652,N_32383,N_32355);
or U32653 (N_32653,N_32454,N_32489);
xnor U32654 (N_32654,N_32269,N_32468);
xor U32655 (N_32655,N_32364,N_32369);
xor U32656 (N_32656,N_32299,N_32413);
and U32657 (N_32657,N_32278,N_32339);
nand U32658 (N_32658,N_32285,N_32379);
or U32659 (N_32659,N_32309,N_32352);
xor U32660 (N_32660,N_32488,N_32428);
nand U32661 (N_32661,N_32319,N_32392);
and U32662 (N_32662,N_32285,N_32443);
nand U32663 (N_32663,N_32492,N_32426);
xor U32664 (N_32664,N_32321,N_32428);
nand U32665 (N_32665,N_32365,N_32272);
and U32666 (N_32666,N_32289,N_32436);
or U32667 (N_32667,N_32457,N_32402);
nand U32668 (N_32668,N_32312,N_32499);
xnor U32669 (N_32669,N_32297,N_32262);
nor U32670 (N_32670,N_32459,N_32408);
and U32671 (N_32671,N_32282,N_32325);
nor U32672 (N_32672,N_32312,N_32291);
or U32673 (N_32673,N_32497,N_32327);
and U32674 (N_32674,N_32383,N_32428);
xor U32675 (N_32675,N_32405,N_32336);
nor U32676 (N_32676,N_32321,N_32368);
and U32677 (N_32677,N_32288,N_32260);
xnor U32678 (N_32678,N_32312,N_32471);
and U32679 (N_32679,N_32301,N_32395);
and U32680 (N_32680,N_32483,N_32286);
and U32681 (N_32681,N_32402,N_32498);
nor U32682 (N_32682,N_32433,N_32332);
nand U32683 (N_32683,N_32281,N_32395);
and U32684 (N_32684,N_32434,N_32419);
nor U32685 (N_32685,N_32293,N_32345);
and U32686 (N_32686,N_32404,N_32464);
or U32687 (N_32687,N_32317,N_32442);
nor U32688 (N_32688,N_32343,N_32381);
and U32689 (N_32689,N_32474,N_32268);
and U32690 (N_32690,N_32335,N_32487);
nand U32691 (N_32691,N_32474,N_32426);
nand U32692 (N_32692,N_32452,N_32286);
nand U32693 (N_32693,N_32432,N_32435);
or U32694 (N_32694,N_32361,N_32308);
nand U32695 (N_32695,N_32440,N_32326);
or U32696 (N_32696,N_32335,N_32280);
nand U32697 (N_32697,N_32456,N_32434);
or U32698 (N_32698,N_32396,N_32427);
xnor U32699 (N_32699,N_32405,N_32362);
or U32700 (N_32700,N_32383,N_32480);
and U32701 (N_32701,N_32388,N_32322);
and U32702 (N_32702,N_32372,N_32269);
nand U32703 (N_32703,N_32466,N_32290);
xnor U32704 (N_32704,N_32438,N_32494);
nor U32705 (N_32705,N_32331,N_32374);
xor U32706 (N_32706,N_32360,N_32475);
xor U32707 (N_32707,N_32456,N_32358);
or U32708 (N_32708,N_32297,N_32425);
or U32709 (N_32709,N_32479,N_32349);
and U32710 (N_32710,N_32442,N_32320);
nor U32711 (N_32711,N_32313,N_32436);
nand U32712 (N_32712,N_32299,N_32395);
xnor U32713 (N_32713,N_32283,N_32257);
or U32714 (N_32714,N_32401,N_32341);
or U32715 (N_32715,N_32388,N_32491);
xnor U32716 (N_32716,N_32384,N_32423);
and U32717 (N_32717,N_32436,N_32405);
or U32718 (N_32718,N_32274,N_32316);
nand U32719 (N_32719,N_32283,N_32354);
nor U32720 (N_32720,N_32466,N_32428);
xnor U32721 (N_32721,N_32409,N_32366);
xor U32722 (N_32722,N_32432,N_32292);
or U32723 (N_32723,N_32316,N_32265);
nand U32724 (N_32724,N_32372,N_32431);
and U32725 (N_32725,N_32489,N_32418);
xor U32726 (N_32726,N_32309,N_32258);
xnor U32727 (N_32727,N_32390,N_32335);
xnor U32728 (N_32728,N_32399,N_32270);
and U32729 (N_32729,N_32303,N_32334);
nand U32730 (N_32730,N_32378,N_32494);
nor U32731 (N_32731,N_32281,N_32492);
xor U32732 (N_32732,N_32320,N_32483);
and U32733 (N_32733,N_32396,N_32492);
or U32734 (N_32734,N_32494,N_32482);
xnor U32735 (N_32735,N_32253,N_32414);
nand U32736 (N_32736,N_32417,N_32259);
nor U32737 (N_32737,N_32375,N_32348);
nor U32738 (N_32738,N_32397,N_32467);
or U32739 (N_32739,N_32372,N_32344);
nor U32740 (N_32740,N_32319,N_32368);
or U32741 (N_32741,N_32484,N_32461);
and U32742 (N_32742,N_32407,N_32454);
or U32743 (N_32743,N_32347,N_32274);
nand U32744 (N_32744,N_32393,N_32428);
or U32745 (N_32745,N_32297,N_32329);
or U32746 (N_32746,N_32349,N_32414);
and U32747 (N_32747,N_32380,N_32466);
or U32748 (N_32748,N_32329,N_32360);
xor U32749 (N_32749,N_32488,N_32426);
or U32750 (N_32750,N_32623,N_32635);
nand U32751 (N_32751,N_32558,N_32641);
nor U32752 (N_32752,N_32663,N_32527);
nor U32753 (N_32753,N_32538,N_32520);
and U32754 (N_32754,N_32511,N_32578);
nand U32755 (N_32755,N_32540,N_32512);
or U32756 (N_32756,N_32725,N_32572);
or U32757 (N_32757,N_32655,N_32592);
and U32758 (N_32758,N_32565,N_32660);
nand U32759 (N_32759,N_32616,N_32588);
and U32760 (N_32760,N_32691,N_32508);
or U32761 (N_32761,N_32646,N_32638);
xor U32762 (N_32762,N_32502,N_32639);
and U32763 (N_32763,N_32524,N_32513);
and U32764 (N_32764,N_32571,N_32585);
nand U32765 (N_32765,N_32703,N_32740);
and U32766 (N_32766,N_32554,N_32579);
nor U32767 (N_32767,N_32622,N_32701);
or U32768 (N_32768,N_32667,N_32574);
and U32769 (N_32769,N_32710,N_32704);
and U32770 (N_32770,N_32723,N_32545);
nand U32771 (N_32771,N_32687,N_32728);
xnor U32772 (N_32772,N_32620,N_32659);
or U32773 (N_32773,N_32549,N_32500);
nand U32774 (N_32774,N_32619,N_32727);
nand U32775 (N_32775,N_32741,N_32544);
nor U32776 (N_32776,N_32736,N_32665);
nand U32777 (N_32777,N_32570,N_32734);
and U32778 (N_32778,N_32539,N_32542);
nand U32779 (N_32779,N_32607,N_32680);
or U32780 (N_32780,N_32551,N_32673);
xnor U32781 (N_32781,N_32681,N_32747);
xor U32782 (N_32782,N_32706,N_32608);
or U32783 (N_32783,N_32679,N_32514);
nand U32784 (N_32784,N_32716,N_32525);
nor U32785 (N_32785,N_32521,N_32656);
xnor U32786 (N_32786,N_32529,N_32614);
or U32787 (N_32787,N_32552,N_32519);
xor U32788 (N_32788,N_32564,N_32684);
and U32789 (N_32789,N_32606,N_32501);
and U32790 (N_32790,N_32748,N_32702);
nor U32791 (N_32791,N_32628,N_32737);
nand U32792 (N_32792,N_32683,N_32651);
nor U32793 (N_32793,N_32615,N_32590);
and U32794 (N_32794,N_32749,N_32694);
nand U32795 (N_32795,N_32535,N_32528);
xnor U32796 (N_32796,N_32582,N_32658);
or U32797 (N_32797,N_32686,N_32647);
nor U32798 (N_32798,N_32746,N_32605);
and U32799 (N_32799,N_32739,N_32547);
nand U32800 (N_32800,N_32721,N_32504);
xnor U32801 (N_32801,N_32555,N_32503);
nand U32802 (N_32802,N_32629,N_32726);
nor U32803 (N_32803,N_32583,N_32642);
nand U32804 (N_32804,N_32695,N_32643);
and U32805 (N_32805,N_32589,N_32711);
and U32806 (N_32806,N_32580,N_32515);
nor U32807 (N_32807,N_32617,N_32560);
and U32808 (N_32808,N_32530,N_32719);
or U32809 (N_32809,N_32633,N_32612);
xor U32810 (N_32810,N_32644,N_32613);
and U32811 (N_32811,N_32671,N_32581);
nor U32812 (N_32812,N_32598,N_32682);
nand U32813 (N_32813,N_32626,N_32696);
nand U32814 (N_32814,N_32599,N_32556);
or U32815 (N_32815,N_32604,N_32713);
xor U32816 (N_32816,N_32591,N_32689);
and U32817 (N_32817,N_32627,N_32705);
or U32818 (N_32818,N_32596,N_32670);
nor U32819 (N_32819,N_32699,N_32603);
or U32820 (N_32820,N_32559,N_32649);
and U32821 (N_32821,N_32692,N_32505);
and U32822 (N_32822,N_32573,N_32700);
or U32823 (N_32823,N_32742,N_32637);
nand U32824 (N_32824,N_32664,N_32715);
or U32825 (N_32825,N_32611,N_32677);
or U32826 (N_32826,N_32553,N_32669);
nand U32827 (N_32827,N_32523,N_32506);
nand U32828 (N_32828,N_32609,N_32575);
and U32829 (N_32829,N_32546,N_32593);
and U32830 (N_32830,N_32730,N_32640);
and U32831 (N_32831,N_32654,N_32733);
or U32832 (N_32832,N_32724,N_32586);
nand U32833 (N_32833,N_32557,N_32532);
nor U32834 (N_32834,N_32708,N_32632);
and U32835 (N_32835,N_32662,N_32714);
nand U32836 (N_32836,N_32517,N_32735);
or U32837 (N_32837,N_32631,N_32709);
nor U32838 (N_32838,N_32566,N_32674);
nor U32839 (N_32839,N_32732,N_32536);
nand U32840 (N_32840,N_32743,N_32533);
nand U32841 (N_32841,N_32685,N_32738);
and U32842 (N_32842,N_32518,N_32698);
xor U32843 (N_32843,N_32645,N_32722);
or U32844 (N_32844,N_32634,N_32595);
nand U32845 (N_32845,N_32569,N_32526);
nand U32846 (N_32846,N_32657,N_32576);
nand U32847 (N_32847,N_32676,N_32668);
or U32848 (N_32848,N_32744,N_32618);
and U32849 (N_32849,N_32510,N_32688);
xor U32850 (N_32850,N_32534,N_32597);
xor U32851 (N_32851,N_32666,N_32567);
nor U32852 (N_32852,N_32672,N_32577);
and U32853 (N_32853,N_32652,N_32675);
or U32854 (N_32854,N_32636,N_32601);
nor U32855 (N_32855,N_32712,N_32624);
nor U32856 (N_32856,N_32522,N_32717);
or U32857 (N_32857,N_32625,N_32548);
and U32858 (N_32858,N_32720,N_32690);
xor U32859 (N_32859,N_32563,N_32509);
xnor U32860 (N_32860,N_32600,N_32587);
nand U32861 (N_32861,N_32621,N_32693);
nand U32862 (N_32862,N_32653,N_32507);
xnor U32863 (N_32863,N_32543,N_32550);
or U32864 (N_32864,N_32697,N_32610);
nand U32865 (N_32865,N_32707,N_32630);
nand U32866 (N_32866,N_32568,N_32650);
and U32867 (N_32867,N_32584,N_32745);
nor U32868 (N_32868,N_32594,N_32718);
nand U32869 (N_32869,N_32531,N_32731);
and U32870 (N_32870,N_32562,N_32561);
nand U32871 (N_32871,N_32541,N_32602);
nand U32872 (N_32872,N_32678,N_32648);
xor U32873 (N_32873,N_32516,N_32729);
and U32874 (N_32874,N_32661,N_32537);
xor U32875 (N_32875,N_32507,N_32541);
and U32876 (N_32876,N_32641,N_32662);
and U32877 (N_32877,N_32642,N_32590);
nand U32878 (N_32878,N_32559,N_32601);
nor U32879 (N_32879,N_32726,N_32655);
or U32880 (N_32880,N_32554,N_32521);
xnor U32881 (N_32881,N_32533,N_32728);
and U32882 (N_32882,N_32655,N_32606);
nand U32883 (N_32883,N_32597,N_32576);
nand U32884 (N_32884,N_32546,N_32544);
or U32885 (N_32885,N_32735,N_32612);
or U32886 (N_32886,N_32567,N_32556);
or U32887 (N_32887,N_32603,N_32648);
and U32888 (N_32888,N_32502,N_32598);
xor U32889 (N_32889,N_32531,N_32636);
or U32890 (N_32890,N_32673,N_32731);
nand U32891 (N_32891,N_32607,N_32593);
nand U32892 (N_32892,N_32638,N_32589);
and U32893 (N_32893,N_32680,N_32683);
xnor U32894 (N_32894,N_32652,N_32695);
nand U32895 (N_32895,N_32597,N_32706);
nor U32896 (N_32896,N_32639,N_32647);
or U32897 (N_32897,N_32592,N_32518);
xor U32898 (N_32898,N_32573,N_32606);
xor U32899 (N_32899,N_32557,N_32694);
nor U32900 (N_32900,N_32535,N_32652);
nand U32901 (N_32901,N_32586,N_32557);
xnor U32902 (N_32902,N_32590,N_32563);
nor U32903 (N_32903,N_32629,N_32724);
or U32904 (N_32904,N_32637,N_32628);
or U32905 (N_32905,N_32582,N_32624);
nand U32906 (N_32906,N_32683,N_32539);
or U32907 (N_32907,N_32614,N_32636);
nor U32908 (N_32908,N_32565,N_32599);
nor U32909 (N_32909,N_32654,N_32540);
xnor U32910 (N_32910,N_32580,N_32727);
nand U32911 (N_32911,N_32577,N_32620);
nand U32912 (N_32912,N_32575,N_32541);
or U32913 (N_32913,N_32630,N_32646);
xor U32914 (N_32914,N_32733,N_32642);
xnor U32915 (N_32915,N_32546,N_32642);
nand U32916 (N_32916,N_32676,N_32741);
and U32917 (N_32917,N_32549,N_32714);
and U32918 (N_32918,N_32711,N_32536);
nor U32919 (N_32919,N_32681,N_32601);
and U32920 (N_32920,N_32532,N_32583);
nor U32921 (N_32921,N_32544,N_32737);
nor U32922 (N_32922,N_32697,N_32702);
or U32923 (N_32923,N_32508,N_32725);
nand U32924 (N_32924,N_32706,N_32701);
and U32925 (N_32925,N_32708,N_32623);
nor U32926 (N_32926,N_32653,N_32577);
xnor U32927 (N_32927,N_32669,N_32580);
nor U32928 (N_32928,N_32639,N_32528);
and U32929 (N_32929,N_32663,N_32596);
xnor U32930 (N_32930,N_32689,N_32680);
xnor U32931 (N_32931,N_32579,N_32529);
nand U32932 (N_32932,N_32648,N_32653);
nand U32933 (N_32933,N_32612,N_32725);
nor U32934 (N_32934,N_32592,N_32623);
xnor U32935 (N_32935,N_32596,N_32623);
nor U32936 (N_32936,N_32666,N_32677);
nor U32937 (N_32937,N_32673,N_32681);
nor U32938 (N_32938,N_32603,N_32638);
and U32939 (N_32939,N_32553,N_32585);
or U32940 (N_32940,N_32670,N_32681);
or U32941 (N_32941,N_32688,N_32587);
or U32942 (N_32942,N_32578,N_32639);
nor U32943 (N_32943,N_32513,N_32743);
xor U32944 (N_32944,N_32594,N_32627);
nand U32945 (N_32945,N_32507,N_32676);
or U32946 (N_32946,N_32628,N_32642);
or U32947 (N_32947,N_32615,N_32707);
xnor U32948 (N_32948,N_32590,N_32604);
nor U32949 (N_32949,N_32700,N_32609);
nand U32950 (N_32950,N_32630,N_32541);
and U32951 (N_32951,N_32536,N_32717);
and U32952 (N_32952,N_32599,N_32543);
or U32953 (N_32953,N_32596,N_32508);
or U32954 (N_32954,N_32713,N_32652);
and U32955 (N_32955,N_32525,N_32674);
and U32956 (N_32956,N_32632,N_32618);
or U32957 (N_32957,N_32651,N_32502);
or U32958 (N_32958,N_32630,N_32654);
or U32959 (N_32959,N_32663,N_32648);
and U32960 (N_32960,N_32558,N_32706);
nand U32961 (N_32961,N_32646,N_32743);
nand U32962 (N_32962,N_32679,N_32658);
nor U32963 (N_32963,N_32549,N_32744);
nor U32964 (N_32964,N_32719,N_32584);
xnor U32965 (N_32965,N_32655,N_32611);
or U32966 (N_32966,N_32611,N_32718);
nor U32967 (N_32967,N_32638,N_32573);
and U32968 (N_32968,N_32746,N_32747);
xor U32969 (N_32969,N_32564,N_32565);
nor U32970 (N_32970,N_32559,N_32588);
nand U32971 (N_32971,N_32683,N_32654);
xor U32972 (N_32972,N_32745,N_32563);
nand U32973 (N_32973,N_32641,N_32546);
nand U32974 (N_32974,N_32507,N_32667);
xor U32975 (N_32975,N_32636,N_32666);
or U32976 (N_32976,N_32741,N_32646);
or U32977 (N_32977,N_32508,N_32698);
nor U32978 (N_32978,N_32646,N_32566);
or U32979 (N_32979,N_32644,N_32749);
nor U32980 (N_32980,N_32602,N_32525);
xor U32981 (N_32981,N_32525,N_32530);
xnor U32982 (N_32982,N_32730,N_32524);
nor U32983 (N_32983,N_32682,N_32511);
nand U32984 (N_32984,N_32520,N_32689);
and U32985 (N_32985,N_32624,N_32620);
or U32986 (N_32986,N_32590,N_32706);
and U32987 (N_32987,N_32602,N_32612);
xnor U32988 (N_32988,N_32676,N_32717);
or U32989 (N_32989,N_32519,N_32583);
nand U32990 (N_32990,N_32504,N_32512);
nand U32991 (N_32991,N_32641,N_32682);
or U32992 (N_32992,N_32563,N_32669);
or U32993 (N_32993,N_32731,N_32618);
or U32994 (N_32994,N_32691,N_32637);
nor U32995 (N_32995,N_32564,N_32569);
nand U32996 (N_32996,N_32726,N_32588);
or U32997 (N_32997,N_32658,N_32707);
nor U32998 (N_32998,N_32708,N_32597);
and U32999 (N_32999,N_32500,N_32621);
nor U33000 (N_33000,N_32815,N_32903);
or U33001 (N_33001,N_32847,N_32914);
nor U33002 (N_33002,N_32832,N_32809);
or U33003 (N_33003,N_32759,N_32766);
nand U33004 (N_33004,N_32896,N_32968);
xnor U33005 (N_33005,N_32886,N_32774);
nand U33006 (N_33006,N_32854,N_32934);
and U33007 (N_33007,N_32825,N_32911);
or U33008 (N_33008,N_32818,N_32959);
nand U33009 (N_33009,N_32865,N_32802);
or U33010 (N_33010,N_32816,N_32840);
xor U33011 (N_33011,N_32789,N_32933);
and U33012 (N_33012,N_32915,N_32790);
nand U33013 (N_33013,N_32960,N_32850);
nand U33014 (N_33014,N_32918,N_32885);
nor U33015 (N_33015,N_32770,N_32877);
or U33016 (N_33016,N_32967,N_32970);
nor U33017 (N_33017,N_32921,N_32949);
and U33018 (N_33018,N_32930,N_32812);
or U33019 (N_33019,N_32834,N_32971);
nor U33020 (N_33020,N_32807,N_32909);
nor U33021 (N_33021,N_32999,N_32983);
xor U33022 (N_33022,N_32820,N_32767);
xnor U33023 (N_33023,N_32758,N_32898);
nand U33024 (N_33024,N_32778,N_32799);
xor U33025 (N_33025,N_32926,N_32943);
nand U33026 (N_33026,N_32768,N_32964);
and U33027 (N_33027,N_32864,N_32821);
nand U33028 (N_33028,N_32756,N_32856);
nor U33029 (N_33029,N_32878,N_32845);
or U33030 (N_33030,N_32777,N_32861);
nor U33031 (N_33031,N_32848,N_32793);
nand U33032 (N_33032,N_32876,N_32763);
nand U33033 (N_33033,N_32944,N_32953);
and U33034 (N_33034,N_32884,N_32986);
and U33035 (N_33035,N_32773,N_32843);
nand U33036 (N_33036,N_32753,N_32868);
or U33037 (N_33037,N_32761,N_32795);
or U33038 (N_33038,N_32754,N_32811);
and U33039 (N_33039,N_32955,N_32800);
xor U33040 (N_33040,N_32844,N_32829);
nand U33041 (N_33041,N_32855,N_32880);
and U33042 (N_33042,N_32905,N_32931);
xor U33043 (N_33043,N_32846,N_32836);
nand U33044 (N_33044,N_32912,N_32833);
nor U33045 (N_33045,N_32966,N_32819);
nand U33046 (N_33046,N_32991,N_32988);
and U33047 (N_33047,N_32920,N_32980);
or U33048 (N_33048,N_32797,N_32922);
nor U33049 (N_33049,N_32941,N_32917);
or U33050 (N_33050,N_32958,N_32869);
nor U33051 (N_33051,N_32830,N_32948);
xnor U33052 (N_33052,N_32978,N_32977);
or U33053 (N_33053,N_32791,N_32938);
and U33054 (N_33054,N_32858,N_32798);
and U33055 (N_33055,N_32989,N_32751);
or U33056 (N_33056,N_32952,N_32822);
or U33057 (N_33057,N_32862,N_32769);
nor U33058 (N_33058,N_32881,N_32838);
nor U33059 (N_33059,N_32771,N_32801);
xnor U33060 (N_33060,N_32965,N_32806);
nor U33061 (N_33061,N_32932,N_32784);
and U33062 (N_33062,N_32853,N_32923);
nor U33063 (N_33063,N_32987,N_32985);
xor U33064 (N_33064,N_32904,N_32908);
xor U33065 (N_33065,N_32835,N_32849);
or U33066 (N_33066,N_32870,N_32940);
nor U33067 (N_33067,N_32863,N_32924);
or U33068 (N_33068,N_32919,N_32950);
nor U33069 (N_33069,N_32872,N_32956);
and U33070 (N_33070,N_32982,N_32814);
xnor U33071 (N_33071,N_32936,N_32975);
xnor U33072 (N_33072,N_32851,N_32894);
nand U33073 (N_33073,N_32782,N_32757);
and U33074 (N_33074,N_32939,N_32901);
and U33075 (N_33075,N_32883,N_32997);
nand U33076 (N_33076,N_32906,N_32852);
and U33077 (N_33077,N_32826,N_32925);
xnor U33078 (N_33078,N_32857,N_32962);
nand U33079 (N_33079,N_32951,N_32786);
xnor U33080 (N_33080,N_32867,N_32947);
nand U33081 (N_33081,N_32895,N_32890);
and U33082 (N_33082,N_32875,N_32866);
and U33083 (N_33083,N_32963,N_32837);
xnor U33084 (N_33084,N_32892,N_32755);
xor U33085 (N_33085,N_32992,N_32887);
xor U33086 (N_33086,N_32805,N_32860);
or U33087 (N_33087,N_32961,N_32808);
and U33088 (N_33088,N_32817,N_32957);
nor U33089 (N_33089,N_32927,N_32760);
xnor U33090 (N_33090,N_32996,N_32796);
or U33091 (N_33091,N_32882,N_32841);
and U33092 (N_33092,N_32879,N_32910);
nor U33093 (N_33093,N_32973,N_32780);
xor U33094 (N_33094,N_32827,N_32781);
nor U33095 (N_33095,N_32998,N_32913);
nor U33096 (N_33096,N_32981,N_32979);
or U33097 (N_33097,N_32937,N_32750);
and U33098 (N_33098,N_32976,N_32889);
nand U33099 (N_33099,N_32893,N_32810);
xor U33100 (N_33100,N_32765,N_32839);
nor U33101 (N_33101,N_32779,N_32942);
xor U33102 (N_33102,N_32762,N_32974);
and U33103 (N_33103,N_32928,N_32929);
xor U33104 (N_33104,N_32907,N_32823);
nor U33105 (N_33105,N_32803,N_32935);
and U33106 (N_33106,N_32787,N_32804);
and U33107 (N_33107,N_32946,N_32871);
and U33108 (N_33108,N_32954,N_32900);
xor U33109 (N_33109,N_32764,N_32994);
nand U33110 (N_33110,N_32828,N_32776);
xnor U33111 (N_33111,N_32772,N_32899);
nand U33112 (N_33112,N_32831,N_32995);
and U33113 (N_33113,N_32972,N_32824);
nand U33114 (N_33114,N_32897,N_32873);
xnor U33115 (N_33115,N_32916,N_32785);
or U33116 (N_33116,N_32891,N_32842);
and U33117 (N_33117,N_32792,N_32775);
nand U33118 (N_33118,N_32752,N_32945);
or U33119 (N_33119,N_32783,N_32813);
nand U33120 (N_33120,N_32969,N_32859);
xnor U33121 (N_33121,N_32984,N_32788);
xor U33122 (N_33122,N_32993,N_32874);
xor U33123 (N_33123,N_32794,N_32888);
xor U33124 (N_33124,N_32902,N_32990);
and U33125 (N_33125,N_32917,N_32808);
xnor U33126 (N_33126,N_32776,N_32935);
and U33127 (N_33127,N_32862,N_32835);
and U33128 (N_33128,N_32913,N_32816);
nor U33129 (N_33129,N_32994,N_32993);
nor U33130 (N_33130,N_32768,N_32937);
or U33131 (N_33131,N_32855,N_32970);
and U33132 (N_33132,N_32865,N_32751);
and U33133 (N_33133,N_32908,N_32877);
nor U33134 (N_33134,N_32771,N_32870);
and U33135 (N_33135,N_32918,N_32824);
nand U33136 (N_33136,N_32753,N_32791);
xnor U33137 (N_33137,N_32972,N_32815);
nand U33138 (N_33138,N_32766,N_32921);
and U33139 (N_33139,N_32778,N_32890);
or U33140 (N_33140,N_32774,N_32879);
and U33141 (N_33141,N_32795,N_32937);
and U33142 (N_33142,N_32762,N_32918);
xnor U33143 (N_33143,N_32997,N_32786);
and U33144 (N_33144,N_32845,N_32897);
xnor U33145 (N_33145,N_32978,N_32825);
and U33146 (N_33146,N_32950,N_32763);
nor U33147 (N_33147,N_32765,N_32893);
nand U33148 (N_33148,N_32761,N_32896);
or U33149 (N_33149,N_32797,N_32806);
or U33150 (N_33150,N_32926,N_32921);
nor U33151 (N_33151,N_32867,N_32750);
or U33152 (N_33152,N_32759,N_32817);
and U33153 (N_33153,N_32845,N_32791);
xor U33154 (N_33154,N_32853,N_32956);
nor U33155 (N_33155,N_32892,N_32974);
nand U33156 (N_33156,N_32907,N_32824);
xnor U33157 (N_33157,N_32776,N_32763);
or U33158 (N_33158,N_32894,N_32890);
or U33159 (N_33159,N_32825,N_32956);
and U33160 (N_33160,N_32896,N_32879);
xor U33161 (N_33161,N_32900,N_32827);
or U33162 (N_33162,N_32890,N_32945);
and U33163 (N_33163,N_32777,N_32915);
or U33164 (N_33164,N_32770,N_32784);
nand U33165 (N_33165,N_32890,N_32878);
or U33166 (N_33166,N_32910,N_32940);
xnor U33167 (N_33167,N_32776,N_32967);
nor U33168 (N_33168,N_32840,N_32998);
nand U33169 (N_33169,N_32944,N_32782);
or U33170 (N_33170,N_32869,N_32854);
or U33171 (N_33171,N_32994,N_32959);
xor U33172 (N_33172,N_32835,N_32931);
and U33173 (N_33173,N_32988,N_32985);
nand U33174 (N_33174,N_32792,N_32924);
xnor U33175 (N_33175,N_32991,N_32752);
and U33176 (N_33176,N_32754,N_32823);
or U33177 (N_33177,N_32776,N_32851);
and U33178 (N_33178,N_32897,N_32804);
nor U33179 (N_33179,N_32875,N_32879);
xor U33180 (N_33180,N_32784,N_32750);
and U33181 (N_33181,N_32863,N_32876);
xnor U33182 (N_33182,N_32789,N_32773);
xor U33183 (N_33183,N_32926,N_32816);
nand U33184 (N_33184,N_32863,N_32778);
or U33185 (N_33185,N_32842,N_32950);
xnor U33186 (N_33186,N_32924,N_32968);
or U33187 (N_33187,N_32951,N_32828);
nor U33188 (N_33188,N_32917,N_32910);
xnor U33189 (N_33189,N_32857,N_32839);
xnor U33190 (N_33190,N_32877,N_32944);
or U33191 (N_33191,N_32754,N_32964);
xor U33192 (N_33192,N_32751,N_32798);
and U33193 (N_33193,N_32990,N_32917);
or U33194 (N_33194,N_32762,N_32767);
nor U33195 (N_33195,N_32884,N_32827);
xor U33196 (N_33196,N_32773,N_32924);
nor U33197 (N_33197,N_32916,N_32982);
or U33198 (N_33198,N_32803,N_32930);
nor U33199 (N_33199,N_32807,N_32759);
and U33200 (N_33200,N_32829,N_32891);
xor U33201 (N_33201,N_32911,N_32963);
and U33202 (N_33202,N_32995,N_32789);
or U33203 (N_33203,N_32862,N_32893);
or U33204 (N_33204,N_32768,N_32976);
xnor U33205 (N_33205,N_32918,N_32835);
and U33206 (N_33206,N_32780,N_32925);
xor U33207 (N_33207,N_32957,N_32807);
xor U33208 (N_33208,N_32916,N_32786);
nor U33209 (N_33209,N_32913,N_32902);
nor U33210 (N_33210,N_32980,N_32953);
xnor U33211 (N_33211,N_32771,N_32975);
and U33212 (N_33212,N_32839,N_32817);
and U33213 (N_33213,N_32937,N_32935);
or U33214 (N_33214,N_32952,N_32998);
nand U33215 (N_33215,N_32891,N_32892);
nor U33216 (N_33216,N_32912,N_32826);
nor U33217 (N_33217,N_32801,N_32911);
nor U33218 (N_33218,N_32882,N_32863);
and U33219 (N_33219,N_32925,N_32975);
nand U33220 (N_33220,N_32891,N_32880);
and U33221 (N_33221,N_32815,N_32875);
and U33222 (N_33222,N_32986,N_32895);
and U33223 (N_33223,N_32860,N_32991);
and U33224 (N_33224,N_32798,N_32776);
or U33225 (N_33225,N_32980,N_32961);
or U33226 (N_33226,N_32867,N_32890);
xnor U33227 (N_33227,N_32761,N_32827);
xnor U33228 (N_33228,N_32914,N_32978);
and U33229 (N_33229,N_32912,N_32823);
and U33230 (N_33230,N_32899,N_32902);
nand U33231 (N_33231,N_32874,N_32814);
nand U33232 (N_33232,N_32829,N_32902);
and U33233 (N_33233,N_32937,N_32832);
nor U33234 (N_33234,N_32979,N_32751);
nand U33235 (N_33235,N_32938,N_32778);
nor U33236 (N_33236,N_32852,N_32973);
and U33237 (N_33237,N_32789,N_32870);
or U33238 (N_33238,N_32969,N_32820);
or U33239 (N_33239,N_32948,N_32930);
xnor U33240 (N_33240,N_32978,N_32830);
xnor U33241 (N_33241,N_32798,N_32907);
nand U33242 (N_33242,N_32757,N_32896);
nor U33243 (N_33243,N_32967,N_32863);
xor U33244 (N_33244,N_32879,N_32937);
and U33245 (N_33245,N_32887,N_32883);
nor U33246 (N_33246,N_32760,N_32817);
and U33247 (N_33247,N_32964,N_32784);
and U33248 (N_33248,N_32941,N_32858);
and U33249 (N_33249,N_32898,N_32775);
and U33250 (N_33250,N_33221,N_33199);
xor U33251 (N_33251,N_33149,N_33182);
xor U33252 (N_33252,N_33083,N_33205);
nand U33253 (N_33253,N_33102,N_33174);
nor U33254 (N_33254,N_33235,N_33016);
or U33255 (N_33255,N_33151,N_33075);
nor U33256 (N_33256,N_33076,N_33132);
xnor U33257 (N_33257,N_33040,N_33024);
xor U33258 (N_33258,N_33012,N_33164);
xnor U33259 (N_33259,N_33120,N_33062);
xor U33260 (N_33260,N_33082,N_33013);
and U33261 (N_33261,N_33190,N_33006);
xor U33262 (N_33262,N_33050,N_33162);
nand U33263 (N_33263,N_33131,N_33070);
xor U33264 (N_33264,N_33063,N_33193);
and U33265 (N_33265,N_33072,N_33121);
or U33266 (N_33266,N_33023,N_33157);
or U33267 (N_33267,N_33052,N_33169);
xnor U33268 (N_33268,N_33002,N_33033);
or U33269 (N_33269,N_33030,N_33163);
and U33270 (N_33270,N_33233,N_33108);
nor U33271 (N_33271,N_33191,N_33207);
nand U33272 (N_33272,N_33056,N_33154);
xnor U33273 (N_33273,N_33046,N_33137);
and U33274 (N_33274,N_33077,N_33009);
nand U33275 (N_33275,N_33015,N_33194);
and U33276 (N_33276,N_33152,N_33029);
or U33277 (N_33277,N_33085,N_33160);
and U33278 (N_33278,N_33247,N_33051);
nor U33279 (N_33279,N_33088,N_33228);
or U33280 (N_33280,N_33113,N_33143);
or U33281 (N_33281,N_33204,N_33220);
nand U33282 (N_33282,N_33064,N_33045);
and U33283 (N_33283,N_33008,N_33166);
or U33284 (N_33284,N_33101,N_33014);
and U33285 (N_33285,N_33249,N_33058);
and U33286 (N_33286,N_33195,N_33216);
and U33287 (N_33287,N_33021,N_33031);
nor U33288 (N_33288,N_33068,N_33153);
xnor U33289 (N_33289,N_33211,N_33104);
and U33290 (N_33290,N_33073,N_33186);
nand U33291 (N_33291,N_33087,N_33141);
and U33292 (N_33292,N_33133,N_33219);
and U33293 (N_33293,N_33043,N_33167);
xor U33294 (N_33294,N_33078,N_33231);
nor U33295 (N_33295,N_33042,N_33138);
or U33296 (N_33296,N_33244,N_33148);
nor U33297 (N_33297,N_33208,N_33209);
xnor U33298 (N_33298,N_33242,N_33177);
or U33299 (N_33299,N_33094,N_33188);
or U33300 (N_33300,N_33055,N_33217);
nand U33301 (N_33301,N_33005,N_33239);
or U33302 (N_33302,N_33202,N_33041);
nand U33303 (N_33303,N_33060,N_33245);
or U33304 (N_33304,N_33097,N_33053);
nand U33305 (N_33305,N_33067,N_33165);
xnor U33306 (N_33306,N_33238,N_33059);
or U33307 (N_33307,N_33183,N_33147);
or U33308 (N_33308,N_33081,N_33025);
and U33309 (N_33309,N_33236,N_33019);
and U33310 (N_33310,N_33126,N_33084);
or U33311 (N_33311,N_33028,N_33139);
and U33312 (N_33312,N_33173,N_33071);
xor U33313 (N_33313,N_33079,N_33069);
xor U33314 (N_33314,N_33004,N_33170);
and U33315 (N_33315,N_33035,N_33196);
nand U33316 (N_33316,N_33061,N_33054);
nor U33317 (N_33317,N_33158,N_33232);
or U33318 (N_33318,N_33122,N_33037);
nand U33319 (N_33319,N_33017,N_33145);
xnor U33320 (N_33320,N_33189,N_33192);
nor U33321 (N_33321,N_33038,N_33213);
nor U33322 (N_33322,N_33119,N_33246);
or U33323 (N_33323,N_33091,N_33155);
nand U33324 (N_33324,N_33111,N_33210);
or U33325 (N_33325,N_33020,N_33107);
xor U33326 (N_33326,N_33034,N_33048);
and U33327 (N_33327,N_33206,N_33144);
and U33328 (N_33328,N_33156,N_33172);
and U33329 (N_33329,N_33112,N_33047);
nor U33330 (N_33330,N_33110,N_33098);
xor U33331 (N_33331,N_33032,N_33080);
or U33332 (N_33332,N_33197,N_33136);
and U33333 (N_33333,N_33168,N_33036);
nor U33334 (N_33334,N_33116,N_33212);
nor U33335 (N_33335,N_33099,N_33114);
or U33336 (N_33336,N_33134,N_33175);
nor U33337 (N_33337,N_33100,N_33001);
xnor U33338 (N_33338,N_33003,N_33011);
and U33339 (N_33339,N_33117,N_33184);
and U33340 (N_33340,N_33142,N_33198);
or U33341 (N_33341,N_33159,N_33105);
nand U33342 (N_33342,N_33089,N_33225);
and U33343 (N_33343,N_33027,N_33127);
xor U33344 (N_33344,N_33171,N_33026);
nor U33345 (N_33345,N_33074,N_33000);
or U33346 (N_33346,N_33092,N_33044);
xor U33347 (N_33347,N_33185,N_33125);
xnor U33348 (N_33348,N_33123,N_33178);
nor U33349 (N_33349,N_33103,N_33203);
or U33350 (N_33350,N_33234,N_33227);
and U33351 (N_33351,N_33229,N_33241);
and U33352 (N_33352,N_33022,N_33201);
or U33353 (N_33353,N_33129,N_33214);
nand U33354 (N_33354,N_33049,N_33200);
and U33355 (N_33355,N_33140,N_33230);
xor U33356 (N_33356,N_33187,N_33215);
xor U33357 (N_33357,N_33240,N_33130);
and U33358 (N_33358,N_33124,N_33109);
nor U33359 (N_33359,N_33181,N_33010);
and U33360 (N_33360,N_33161,N_33218);
nand U33361 (N_33361,N_33150,N_33090);
nand U33362 (N_33362,N_33179,N_33248);
xor U33363 (N_33363,N_33237,N_33066);
xor U33364 (N_33364,N_33243,N_33095);
and U33365 (N_33365,N_33146,N_33118);
and U33366 (N_33366,N_33176,N_33128);
nand U33367 (N_33367,N_33224,N_33096);
xnor U33368 (N_33368,N_33086,N_33222);
nand U33369 (N_33369,N_33039,N_33223);
and U33370 (N_33370,N_33180,N_33065);
and U33371 (N_33371,N_33093,N_33106);
or U33372 (N_33372,N_33007,N_33226);
xor U33373 (N_33373,N_33135,N_33018);
nor U33374 (N_33374,N_33057,N_33115);
xnor U33375 (N_33375,N_33118,N_33209);
nor U33376 (N_33376,N_33219,N_33175);
or U33377 (N_33377,N_33160,N_33244);
nand U33378 (N_33378,N_33083,N_33102);
and U33379 (N_33379,N_33118,N_33074);
nor U33380 (N_33380,N_33122,N_33113);
and U33381 (N_33381,N_33240,N_33090);
nor U33382 (N_33382,N_33050,N_33146);
nor U33383 (N_33383,N_33041,N_33063);
or U33384 (N_33384,N_33187,N_33118);
xnor U33385 (N_33385,N_33222,N_33108);
and U33386 (N_33386,N_33099,N_33142);
nand U33387 (N_33387,N_33020,N_33206);
nand U33388 (N_33388,N_33156,N_33114);
xnor U33389 (N_33389,N_33161,N_33129);
xnor U33390 (N_33390,N_33153,N_33128);
nor U33391 (N_33391,N_33056,N_33211);
nand U33392 (N_33392,N_33046,N_33094);
or U33393 (N_33393,N_33172,N_33104);
nor U33394 (N_33394,N_33004,N_33190);
and U33395 (N_33395,N_33235,N_33211);
and U33396 (N_33396,N_33084,N_33059);
nand U33397 (N_33397,N_33149,N_33104);
xor U33398 (N_33398,N_33238,N_33155);
and U33399 (N_33399,N_33100,N_33112);
nand U33400 (N_33400,N_33199,N_33061);
nor U33401 (N_33401,N_33031,N_33234);
or U33402 (N_33402,N_33176,N_33016);
xor U33403 (N_33403,N_33054,N_33176);
xor U33404 (N_33404,N_33000,N_33173);
or U33405 (N_33405,N_33233,N_33214);
nand U33406 (N_33406,N_33130,N_33235);
or U33407 (N_33407,N_33240,N_33233);
xnor U33408 (N_33408,N_33152,N_33010);
xor U33409 (N_33409,N_33000,N_33234);
and U33410 (N_33410,N_33145,N_33072);
xor U33411 (N_33411,N_33022,N_33007);
xor U33412 (N_33412,N_33211,N_33024);
nand U33413 (N_33413,N_33004,N_33084);
nand U33414 (N_33414,N_33151,N_33113);
nand U33415 (N_33415,N_33174,N_33088);
nand U33416 (N_33416,N_33243,N_33200);
xnor U33417 (N_33417,N_33165,N_33190);
nand U33418 (N_33418,N_33179,N_33052);
nor U33419 (N_33419,N_33079,N_33167);
nor U33420 (N_33420,N_33149,N_33076);
xor U33421 (N_33421,N_33228,N_33234);
or U33422 (N_33422,N_33035,N_33063);
nor U33423 (N_33423,N_33184,N_33065);
xnor U33424 (N_33424,N_33045,N_33238);
or U33425 (N_33425,N_33185,N_33228);
and U33426 (N_33426,N_33165,N_33086);
and U33427 (N_33427,N_33168,N_33113);
nor U33428 (N_33428,N_33209,N_33131);
or U33429 (N_33429,N_33222,N_33197);
or U33430 (N_33430,N_33193,N_33104);
nor U33431 (N_33431,N_33004,N_33223);
xor U33432 (N_33432,N_33200,N_33207);
and U33433 (N_33433,N_33009,N_33015);
nand U33434 (N_33434,N_33236,N_33072);
xnor U33435 (N_33435,N_33101,N_33134);
xor U33436 (N_33436,N_33109,N_33003);
nand U33437 (N_33437,N_33231,N_33051);
nor U33438 (N_33438,N_33111,N_33102);
xnor U33439 (N_33439,N_33018,N_33075);
nand U33440 (N_33440,N_33201,N_33230);
nand U33441 (N_33441,N_33113,N_33046);
nand U33442 (N_33442,N_33146,N_33226);
nor U33443 (N_33443,N_33138,N_33097);
and U33444 (N_33444,N_33141,N_33041);
nor U33445 (N_33445,N_33162,N_33115);
nor U33446 (N_33446,N_33207,N_33097);
and U33447 (N_33447,N_33245,N_33145);
and U33448 (N_33448,N_33217,N_33205);
nand U33449 (N_33449,N_33016,N_33047);
or U33450 (N_33450,N_33094,N_33196);
xor U33451 (N_33451,N_33231,N_33137);
and U33452 (N_33452,N_33002,N_33134);
nor U33453 (N_33453,N_33084,N_33028);
or U33454 (N_33454,N_33033,N_33017);
nor U33455 (N_33455,N_33236,N_33003);
nor U33456 (N_33456,N_33128,N_33006);
nand U33457 (N_33457,N_33097,N_33176);
and U33458 (N_33458,N_33187,N_33026);
nor U33459 (N_33459,N_33002,N_33099);
nand U33460 (N_33460,N_33015,N_33100);
xor U33461 (N_33461,N_33194,N_33235);
xor U33462 (N_33462,N_33003,N_33141);
or U33463 (N_33463,N_33181,N_33065);
or U33464 (N_33464,N_33167,N_33045);
nand U33465 (N_33465,N_33067,N_33227);
nand U33466 (N_33466,N_33014,N_33229);
or U33467 (N_33467,N_33002,N_33057);
nand U33468 (N_33468,N_33083,N_33064);
and U33469 (N_33469,N_33133,N_33085);
nor U33470 (N_33470,N_33022,N_33103);
and U33471 (N_33471,N_33077,N_33033);
xor U33472 (N_33472,N_33152,N_33115);
nand U33473 (N_33473,N_33229,N_33177);
nand U33474 (N_33474,N_33087,N_33227);
nor U33475 (N_33475,N_33077,N_33097);
nand U33476 (N_33476,N_33174,N_33076);
and U33477 (N_33477,N_33187,N_33070);
nand U33478 (N_33478,N_33114,N_33178);
or U33479 (N_33479,N_33157,N_33040);
nor U33480 (N_33480,N_33182,N_33086);
or U33481 (N_33481,N_33073,N_33065);
nand U33482 (N_33482,N_33031,N_33003);
nand U33483 (N_33483,N_33068,N_33182);
xor U33484 (N_33484,N_33212,N_33051);
nand U33485 (N_33485,N_33209,N_33048);
or U33486 (N_33486,N_33101,N_33039);
and U33487 (N_33487,N_33007,N_33078);
nor U33488 (N_33488,N_33204,N_33010);
nand U33489 (N_33489,N_33222,N_33232);
nand U33490 (N_33490,N_33130,N_33085);
or U33491 (N_33491,N_33159,N_33183);
nand U33492 (N_33492,N_33213,N_33067);
nor U33493 (N_33493,N_33027,N_33044);
nor U33494 (N_33494,N_33074,N_33046);
or U33495 (N_33495,N_33004,N_33146);
and U33496 (N_33496,N_33147,N_33012);
xor U33497 (N_33497,N_33177,N_33157);
xor U33498 (N_33498,N_33103,N_33036);
or U33499 (N_33499,N_33185,N_33236);
nor U33500 (N_33500,N_33262,N_33474);
nand U33501 (N_33501,N_33299,N_33455);
nor U33502 (N_33502,N_33380,N_33288);
nor U33503 (N_33503,N_33497,N_33267);
or U33504 (N_33504,N_33289,N_33470);
or U33505 (N_33505,N_33291,N_33420);
xnor U33506 (N_33506,N_33373,N_33406);
nand U33507 (N_33507,N_33416,N_33303);
xnor U33508 (N_33508,N_33361,N_33413);
nand U33509 (N_33509,N_33486,N_33426);
nand U33510 (N_33510,N_33346,N_33254);
or U33511 (N_33511,N_33448,N_33278);
or U33512 (N_33512,N_33264,N_33394);
and U33513 (N_33513,N_33489,N_33384);
and U33514 (N_33514,N_33461,N_33472);
nand U33515 (N_33515,N_33386,N_33396);
and U33516 (N_33516,N_33319,N_33429);
xor U33517 (N_33517,N_33250,N_33438);
and U33518 (N_33518,N_33366,N_33395);
nand U33519 (N_33519,N_33315,N_33403);
nor U33520 (N_33520,N_33374,N_33440);
and U33521 (N_33521,N_33463,N_33375);
or U33522 (N_33522,N_33333,N_33404);
or U33523 (N_33523,N_33270,N_33482);
nor U33524 (N_33524,N_33391,N_33478);
nand U33525 (N_33525,N_33454,N_33359);
nor U33526 (N_33526,N_33281,N_33480);
and U33527 (N_33527,N_33444,N_33377);
or U33528 (N_33528,N_33447,N_33269);
xor U33529 (N_33529,N_33357,N_33422);
nand U33530 (N_33530,N_33390,N_33485);
nor U33531 (N_33531,N_33276,N_33496);
and U33532 (N_33532,N_33335,N_33273);
nor U33533 (N_33533,N_33378,N_33256);
nand U33534 (N_33534,N_33369,N_33473);
xnor U33535 (N_33535,N_33251,N_33467);
nor U33536 (N_33536,N_33353,N_33477);
nand U33537 (N_33537,N_33405,N_33293);
and U33538 (N_33538,N_33283,N_33450);
nor U33539 (N_33539,N_33253,N_33457);
xnor U33540 (N_33540,N_33311,N_33327);
nand U33541 (N_33541,N_33399,N_33261);
xnor U33542 (N_33542,N_33268,N_33339);
xnor U33543 (N_33543,N_33314,N_33313);
or U33544 (N_33544,N_33487,N_33318);
and U33545 (N_33545,N_33362,N_33322);
nor U33546 (N_33546,N_33295,N_33383);
nor U33547 (N_33547,N_33342,N_33317);
nand U33548 (N_33548,N_33490,N_33464);
and U33549 (N_33549,N_33427,N_33436);
or U33550 (N_33550,N_33257,N_33338);
nand U33551 (N_33551,N_33302,N_33286);
nor U33552 (N_33552,N_33451,N_33398);
nand U33553 (N_33553,N_33458,N_33300);
and U33554 (N_33554,N_33370,N_33259);
nor U33555 (N_33555,N_33441,N_33381);
or U33556 (N_33556,N_33494,N_33323);
nand U33557 (N_33557,N_33424,N_33312);
and U33558 (N_33558,N_33400,N_33280);
nor U33559 (N_33559,N_33471,N_33347);
or U33560 (N_33560,N_33498,N_33354);
nand U33561 (N_33561,N_33428,N_33397);
nor U33562 (N_33562,N_33445,N_33433);
or U33563 (N_33563,N_33414,N_33358);
xnor U33564 (N_33564,N_33456,N_33421);
nand U33565 (N_33565,N_33307,N_33355);
xor U33566 (N_33566,N_33439,N_33479);
nand U33567 (N_33567,N_33304,N_33310);
or U33568 (N_33568,N_33266,N_33402);
xor U33569 (N_33569,N_33349,N_33407);
xor U33570 (N_33570,N_33481,N_33356);
nor U33571 (N_33571,N_33410,N_33385);
nor U33572 (N_33572,N_33483,N_33435);
xnor U33573 (N_33573,N_33459,N_33419);
or U33574 (N_33574,N_33351,N_33341);
nand U33575 (N_33575,N_33475,N_33305);
xnor U33576 (N_33576,N_33308,N_33279);
or U33577 (N_33577,N_33408,N_33326);
and U33578 (N_33578,N_33417,N_33469);
nor U33579 (N_33579,N_33389,N_33282);
or U33580 (N_33580,N_33430,N_33292);
nor U33581 (N_33581,N_33465,N_33336);
xnor U33582 (N_33582,N_33368,N_33484);
nand U33583 (N_33583,N_33392,N_33294);
xnor U33584 (N_33584,N_33255,N_33343);
and U33585 (N_33585,N_33274,N_33320);
nand U33586 (N_33586,N_33443,N_33263);
nand U33587 (N_33587,N_33285,N_33379);
xnor U33588 (N_33588,N_33388,N_33442);
nor U33589 (N_33589,N_33334,N_33409);
nand U33590 (N_33590,N_33446,N_33382);
nor U33591 (N_33591,N_33350,N_33344);
nor U33592 (N_33592,N_33423,N_33431);
or U33593 (N_33593,N_33296,N_33331);
nor U33594 (N_33594,N_33434,N_33258);
or U33595 (N_33595,N_33411,N_33488);
or U33596 (N_33596,N_33321,N_33297);
xor U33597 (N_33597,N_33332,N_33337);
and U33598 (N_33598,N_33372,N_33460);
or U33599 (N_33599,N_33298,N_33328);
nor U33600 (N_33600,N_33376,N_33287);
nor U33601 (N_33601,N_33437,N_33365);
nand U33602 (N_33602,N_33348,N_33387);
or U33603 (N_33603,N_33284,N_33275);
xor U33604 (N_33604,N_33272,N_33316);
nor U33605 (N_33605,N_33345,N_33393);
or U33606 (N_33606,N_33371,N_33360);
nor U33607 (N_33607,N_33493,N_33401);
nor U33608 (N_33608,N_33265,N_33329);
or U33609 (N_33609,N_33301,N_33277);
nor U33610 (N_33610,N_33364,N_33340);
xnor U33611 (N_33611,N_33415,N_33499);
nand U33612 (N_33612,N_33412,N_33432);
xnor U33613 (N_33613,N_33367,N_33260);
nor U33614 (N_33614,N_33466,N_33271);
nor U33615 (N_33615,N_33492,N_33363);
nor U33616 (N_33616,N_33462,N_33491);
or U33617 (N_33617,N_33495,N_33452);
nand U33618 (N_33618,N_33468,N_33290);
nand U33619 (N_33619,N_33352,N_33453);
nor U33620 (N_33620,N_33418,N_33330);
or U33621 (N_33621,N_33425,N_33325);
and U33622 (N_33622,N_33309,N_33252);
or U33623 (N_33623,N_33476,N_33449);
nand U33624 (N_33624,N_33306,N_33324);
xnor U33625 (N_33625,N_33382,N_33379);
xor U33626 (N_33626,N_33458,N_33306);
or U33627 (N_33627,N_33452,N_33367);
and U33628 (N_33628,N_33354,N_33415);
xnor U33629 (N_33629,N_33255,N_33316);
nor U33630 (N_33630,N_33293,N_33455);
and U33631 (N_33631,N_33458,N_33367);
xor U33632 (N_33632,N_33463,N_33250);
nor U33633 (N_33633,N_33409,N_33468);
xnor U33634 (N_33634,N_33415,N_33352);
nor U33635 (N_33635,N_33429,N_33386);
nand U33636 (N_33636,N_33387,N_33491);
and U33637 (N_33637,N_33445,N_33450);
or U33638 (N_33638,N_33450,N_33497);
or U33639 (N_33639,N_33264,N_33465);
and U33640 (N_33640,N_33390,N_33304);
nor U33641 (N_33641,N_33498,N_33321);
nor U33642 (N_33642,N_33385,N_33432);
nand U33643 (N_33643,N_33473,N_33390);
nand U33644 (N_33644,N_33430,N_33406);
nand U33645 (N_33645,N_33287,N_33272);
xnor U33646 (N_33646,N_33275,N_33466);
nand U33647 (N_33647,N_33464,N_33412);
xor U33648 (N_33648,N_33362,N_33472);
and U33649 (N_33649,N_33437,N_33475);
xor U33650 (N_33650,N_33351,N_33377);
nor U33651 (N_33651,N_33391,N_33328);
nor U33652 (N_33652,N_33471,N_33286);
or U33653 (N_33653,N_33255,N_33464);
or U33654 (N_33654,N_33365,N_33409);
nand U33655 (N_33655,N_33349,N_33323);
xor U33656 (N_33656,N_33344,N_33454);
nor U33657 (N_33657,N_33454,N_33367);
or U33658 (N_33658,N_33254,N_33281);
nor U33659 (N_33659,N_33494,N_33460);
or U33660 (N_33660,N_33370,N_33317);
and U33661 (N_33661,N_33381,N_33327);
xnor U33662 (N_33662,N_33326,N_33324);
nand U33663 (N_33663,N_33362,N_33269);
nor U33664 (N_33664,N_33458,N_33396);
xor U33665 (N_33665,N_33467,N_33445);
or U33666 (N_33666,N_33441,N_33319);
nand U33667 (N_33667,N_33307,N_33338);
xnor U33668 (N_33668,N_33296,N_33473);
xor U33669 (N_33669,N_33318,N_33324);
xnor U33670 (N_33670,N_33384,N_33423);
xor U33671 (N_33671,N_33447,N_33324);
xor U33672 (N_33672,N_33303,N_33344);
or U33673 (N_33673,N_33453,N_33254);
xnor U33674 (N_33674,N_33361,N_33440);
nor U33675 (N_33675,N_33287,N_33263);
or U33676 (N_33676,N_33338,N_33340);
nor U33677 (N_33677,N_33345,N_33264);
xor U33678 (N_33678,N_33394,N_33283);
nand U33679 (N_33679,N_33297,N_33410);
nor U33680 (N_33680,N_33286,N_33443);
nand U33681 (N_33681,N_33434,N_33366);
or U33682 (N_33682,N_33300,N_33445);
xor U33683 (N_33683,N_33473,N_33458);
nor U33684 (N_33684,N_33382,N_33334);
and U33685 (N_33685,N_33296,N_33320);
nor U33686 (N_33686,N_33455,N_33334);
and U33687 (N_33687,N_33313,N_33297);
nand U33688 (N_33688,N_33380,N_33479);
or U33689 (N_33689,N_33427,N_33291);
and U33690 (N_33690,N_33298,N_33424);
nor U33691 (N_33691,N_33326,N_33407);
nor U33692 (N_33692,N_33333,N_33260);
and U33693 (N_33693,N_33395,N_33250);
xor U33694 (N_33694,N_33372,N_33484);
nor U33695 (N_33695,N_33354,N_33256);
and U33696 (N_33696,N_33471,N_33456);
or U33697 (N_33697,N_33393,N_33412);
nor U33698 (N_33698,N_33385,N_33394);
xor U33699 (N_33699,N_33452,N_33393);
and U33700 (N_33700,N_33469,N_33323);
nand U33701 (N_33701,N_33266,N_33416);
xor U33702 (N_33702,N_33250,N_33485);
nand U33703 (N_33703,N_33311,N_33286);
and U33704 (N_33704,N_33321,N_33356);
xnor U33705 (N_33705,N_33467,N_33415);
xnor U33706 (N_33706,N_33458,N_33291);
and U33707 (N_33707,N_33337,N_33424);
xnor U33708 (N_33708,N_33404,N_33297);
nand U33709 (N_33709,N_33368,N_33327);
nand U33710 (N_33710,N_33315,N_33473);
or U33711 (N_33711,N_33291,N_33475);
or U33712 (N_33712,N_33436,N_33284);
and U33713 (N_33713,N_33400,N_33300);
and U33714 (N_33714,N_33294,N_33338);
or U33715 (N_33715,N_33272,N_33338);
or U33716 (N_33716,N_33255,N_33285);
and U33717 (N_33717,N_33386,N_33418);
nand U33718 (N_33718,N_33414,N_33276);
nand U33719 (N_33719,N_33425,N_33259);
or U33720 (N_33720,N_33357,N_33293);
and U33721 (N_33721,N_33286,N_33483);
xnor U33722 (N_33722,N_33351,N_33472);
nand U33723 (N_33723,N_33433,N_33280);
or U33724 (N_33724,N_33498,N_33451);
or U33725 (N_33725,N_33383,N_33271);
nor U33726 (N_33726,N_33287,N_33265);
xnor U33727 (N_33727,N_33259,N_33392);
xor U33728 (N_33728,N_33265,N_33268);
and U33729 (N_33729,N_33464,N_33465);
xor U33730 (N_33730,N_33355,N_33489);
or U33731 (N_33731,N_33313,N_33312);
nand U33732 (N_33732,N_33485,N_33338);
nand U33733 (N_33733,N_33281,N_33424);
nor U33734 (N_33734,N_33467,N_33272);
xor U33735 (N_33735,N_33421,N_33409);
nand U33736 (N_33736,N_33271,N_33417);
xnor U33737 (N_33737,N_33392,N_33312);
nor U33738 (N_33738,N_33416,N_33358);
nor U33739 (N_33739,N_33448,N_33394);
xnor U33740 (N_33740,N_33454,N_33403);
and U33741 (N_33741,N_33323,N_33300);
or U33742 (N_33742,N_33336,N_33258);
nor U33743 (N_33743,N_33328,N_33392);
nor U33744 (N_33744,N_33265,N_33324);
and U33745 (N_33745,N_33428,N_33344);
or U33746 (N_33746,N_33334,N_33389);
nand U33747 (N_33747,N_33422,N_33390);
nand U33748 (N_33748,N_33410,N_33406);
and U33749 (N_33749,N_33379,N_33489);
or U33750 (N_33750,N_33578,N_33699);
nor U33751 (N_33751,N_33554,N_33706);
nor U33752 (N_33752,N_33672,N_33619);
xnor U33753 (N_33753,N_33610,N_33624);
xnor U33754 (N_33754,N_33673,N_33580);
nand U33755 (N_33755,N_33703,N_33723);
and U33756 (N_33756,N_33719,N_33535);
nor U33757 (N_33757,N_33568,N_33641);
and U33758 (N_33758,N_33717,N_33542);
nand U33759 (N_33759,N_33654,N_33518);
nor U33760 (N_33760,N_33689,N_33504);
xnor U33761 (N_33761,N_33503,N_33726);
and U33762 (N_33762,N_33537,N_33541);
xnor U33763 (N_33763,N_33708,N_33727);
nor U33764 (N_33764,N_33538,N_33634);
nand U33765 (N_33765,N_33638,N_33546);
nand U33766 (N_33766,N_33704,N_33735);
nor U33767 (N_33767,N_33661,N_33651);
nand U33768 (N_33768,N_33631,N_33682);
nand U33769 (N_33769,N_33599,N_33628);
and U33770 (N_33770,N_33591,N_33570);
and U33771 (N_33771,N_33680,N_33512);
xnor U33772 (N_33772,N_33569,N_33553);
and U33773 (N_33773,N_33574,N_33604);
and U33774 (N_33774,N_33677,N_33687);
xor U33775 (N_33775,N_33564,N_33743);
nor U33776 (N_33776,N_33584,N_33501);
nor U33777 (N_33777,N_33620,N_33738);
and U33778 (N_33778,N_33525,N_33557);
xnor U33779 (N_33779,N_33647,N_33626);
xor U33780 (N_33780,N_33532,N_33595);
nor U33781 (N_33781,N_33614,N_33592);
or U33782 (N_33782,N_33739,N_33508);
and U33783 (N_33783,N_33649,N_33730);
nor U33784 (N_33784,N_33572,N_33731);
nor U33785 (N_33785,N_33734,N_33520);
xor U33786 (N_33786,N_33623,N_33566);
and U33787 (N_33787,N_33548,N_33733);
nand U33788 (N_33788,N_33526,N_33674);
nor U33789 (N_33789,N_33664,N_33729);
xnor U33790 (N_33790,N_33665,N_33539);
or U33791 (N_33791,N_33593,N_33600);
nor U33792 (N_33792,N_33709,N_33728);
nor U33793 (N_33793,N_33506,N_33573);
and U33794 (N_33794,N_33582,N_33710);
or U33795 (N_33795,N_33653,N_33556);
nor U33796 (N_33796,N_33724,N_33702);
nand U33797 (N_33797,N_33605,N_33579);
or U33798 (N_33798,N_33720,N_33581);
or U33799 (N_33799,N_33606,N_33552);
and U33800 (N_33800,N_33718,N_33561);
xnor U33801 (N_33801,N_33607,N_33712);
xnor U33802 (N_33802,N_33521,N_33558);
nand U33803 (N_33803,N_33722,N_33523);
nand U33804 (N_33804,N_33583,N_33744);
or U33805 (N_33805,N_33669,N_33594);
nand U33806 (N_33806,N_33589,N_33666);
xor U33807 (N_33807,N_33622,N_33510);
or U33808 (N_33808,N_33560,N_33602);
xnor U33809 (N_33809,N_33658,N_33650);
xnor U33810 (N_33810,N_33652,N_33696);
and U33811 (N_33811,N_33711,N_33505);
xnor U33812 (N_33812,N_33637,N_33517);
nand U33813 (N_33813,N_33642,N_33567);
nor U33814 (N_33814,N_33611,N_33616);
nor U33815 (N_33815,N_33587,N_33742);
and U33816 (N_33816,N_33714,N_33676);
xor U33817 (N_33817,N_33563,N_33571);
nand U33818 (N_33818,N_33635,N_33697);
nor U33819 (N_33819,N_33576,N_33640);
xnor U33820 (N_33820,N_33547,N_33615);
xor U33821 (N_33821,N_33534,N_33705);
xnor U33822 (N_33822,N_33588,N_33543);
nor U33823 (N_33823,N_33540,N_33522);
nand U33824 (N_33824,N_33528,N_33693);
xor U33825 (N_33825,N_33740,N_33630);
xnor U33826 (N_33826,N_33684,N_33559);
nand U33827 (N_33827,N_33700,N_33617);
and U33828 (N_33828,N_33660,N_33685);
and U33829 (N_33829,N_33681,N_33633);
xor U33830 (N_33830,N_33713,N_33632);
nand U33831 (N_33831,N_33545,N_33695);
and U33832 (N_33832,N_33646,N_33678);
or U33833 (N_33833,N_33663,N_33648);
xor U33834 (N_33834,N_33721,N_33612);
and U33835 (N_33835,N_33577,N_33745);
xor U33836 (N_33836,N_33618,N_33550);
xnor U33837 (N_33837,N_33645,N_33502);
xnor U33838 (N_33838,N_33668,N_33597);
nand U33839 (N_33839,N_33688,N_33690);
xor U33840 (N_33840,N_33500,N_33629);
or U33841 (N_33841,N_33749,N_33657);
nand U33842 (N_33842,N_33675,N_33701);
or U33843 (N_33843,N_33686,N_33530);
nand U33844 (N_33844,N_33746,N_33509);
nand U33845 (N_33845,N_33516,N_33585);
or U33846 (N_33846,N_33544,N_33515);
and U33847 (N_33847,N_33698,N_33643);
or U33848 (N_33848,N_33621,N_33694);
and U33849 (N_33849,N_33636,N_33529);
and U33850 (N_33850,N_33608,N_33609);
or U33851 (N_33851,N_33562,N_33565);
and U33852 (N_33852,N_33639,N_33601);
or U33853 (N_33853,N_33692,N_33656);
nor U33854 (N_33854,N_33670,N_33511);
nand U33855 (N_33855,N_33716,N_33555);
nor U33856 (N_33856,N_33575,N_33737);
or U33857 (N_33857,N_33613,N_33549);
nor U33858 (N_33858,N_33736,N_33667);
and U33859 (N_33859,N_33747,N_33644);
and U33860 (N_33860,N_33514,N_33691);
and U33861 (N_33861,N_33551,N_33524);
and U33862 (N_33862,N_33662,N_33625);
nor U33863 (N_33863,N_33596,N_33732);
or U33864 (N_33864,N_33536,N_33725);
xor U33865 (N_33865,N_33627,N_33741);
or U33866 (N_33866,N_33655,N_33748);
nand U33867 (N_33867,N_33679,N_33715);
xor U33868 (N_33868,N_33513,N_33598);
nand U33869 (N_33869,N_33533,N_33659);
and U33870 (N_33870,N_33707,N_33507);
nor U33871 (N_33871,N_33519,N_33527);
and U33872 (N_33872,N_33586,N_33683);
nand U33873 (N_33873,N_33531,N_33671);
nand U33874 (N_33874,N_33590,N_33603);
and U33875 (N_33875,N_33532,N_33735);
or U33876 (N_33876,N_33647,N_33619);
xor U33877 (N_33877,N_33540,N_33700);
and U33878 (N_33878,N_33556,N_33668);
and U33879 (N_33879,N_33644,N_33553);
and U33880 (N_33880,N_33507,N_33524);
or U33881 (N_33881,N_33599,N_33524);
nand U33882 (N_33882,N_33618,N_33615);
or U33883 (N_33883,N_33724,N_33568);
xor U33884 (N_33884,N_33575,N_33705);
xnor U33885 (N_33885,N_33667,N_33593);
nor U33886 (N_33886,N_33507,N_33529);
and U33887 (N_33887,N_33594,N_33698);
nand U33888 (N_33888,N_33590,N_33564);
nand U33889 (N_33889,N_33543,N_33664);
nor U33890 (N_33890,N_33618,N_33518);
or U33891 (N_33891,N_33585,N_33656);
or U33892 (N_33892,N_33708,N_33517);
or U33893 (N_33893,N_33747,N_33643);
xor U33894 (N_33894,N_33690,N_33717);
xor U33895 (N_33895,N_33607,N_33719);
or U33896 (N_33896,N_33593,N_33607);
or U33897 (N_33897,N_33566,N_33667);
xor U33898 (N_33898,N_33505,N_33624);
nor U33899 (N_33899,N_33740,N_33532);
and U33900 (N_33900,N_33642,N_33574);
nand U33901 (N_33901,N_33728,N_33584);
or U33902 (N_33902,N_33585,N_33749);
or U33903 (N_33903,N_33697,N_33705);
and U33904 (N_33904,N_33613,N_33659);
xnor U33905 (N_33905,N_33649,N_33642);
xor U33906 (N_33906,N_33647,N_33670);
or U33907 (N_33907,N_33529,N_33587);
nand U33908 (N_33908,N_33654,N_33642);
or U33909 (N_33909,N_33701,N_33685);
nand U33910 (N_33910,N_33509,N_33733);
nor U33911 (N_33911,N_33539,N_33513);
or U33912 (N_33912,N_33715,N_33560);
or U33913 (N_33913,N_33518,N_33672);
nand U33914 (N_33914,N_33738,N_33560);
or U33915 (N_33915,N_33697,N_33622);
or U33916 (N_33916,N_33549,N_33709);
nor U33917 (N_33917,N_33606,N_33526);
nor U33918 (N_33918,N_33620,N_33529);
nor U33919 (N_33919,N_33605,N_33666);
and U33920 (N_33920,N_33570,N_33732);
nand U33921 (N_33921,N_33647,N_33709);
nand U33922 (N_33922,N_33525,N_33624);
xor U33923 (N_33923,N_33643,N_33584);
nand U33924 (N_33924,N_33747,N_33549);
and U33925 (N_33925,N_33573,N_33610);
nand U33926 (N_33926,N_33531,N_33685);
or U33927 (N_33927,N_33522,N_33525);
and U33928 (N_33928,N_33699,N_33704);
xnor U33929 (N_33929,N_33567,N_33651);
or U33930 (N_33930,N_33530,N_33544);
xor U33931 (N_33931,N_33723,N_33535);
nor U33932 (N_33932,N_33507,N_33604);
nor U33933 (N_33933,N_33596,N_33644);
nand U33934 (N_33934,N_33673,N_33590);
nor U33935 (N_33935,N_33694,N_33592);
nand U33936 (N_33936,N_33737,N_33506);
or U33937 (N_33937,N_33746,N_33675);
nand U33938 (N_33938,N_33542,N_33606);
or U33939 (N_33939,N_33657,N_33641);
nand U33940 (N_33940,N_33658,N_33719);
and U33941 (N_33941,N_33746,N_33719);
nand U33942 (N_33942,N_33630,N_33729);
or U33943 (N_33943,N_33659,N_33569);
nand U33944 (N_33944,N_33677,N_33579);
nand U33945 (N_33945,N_33714,N_33501);
nor U33946 (N_33946,N_33667,N_33604);
nor U33947 (N_33947,N_33628,N_33705);
and U33948 (N_33948,N_33561,N_33544);
nor U33949 (N_33949,N_33693,N_33602);
or U33950 (N_33950,N_33596,N_33605);
nor U33951 (N_33951,N_33657,N_33720);
nor U33952 (N_33952,N_33722,N_33636);
nor U33953 (N_33953,N_33554,N_33582);
nand U33954 (N_33954,N_33729,N_33529);
or U33955 (N_33955,N_33672,N_33542);
nand U33956 (N_33956,N_33625,N_33600);
nor U33957 (N_33957,N_33547,N_33591);
or U33958 (N_33958,N_33717,N_33722);
nor U33959 (N_33959,N_33529,N_33678);
and U33960 (N_33960,N_33551,N_33703);
and U33961 (N_33961,N_33548,N_33528);
xor U33962 (N_33962,N_33654,N_33623);
nor U33963 (N_33963,N_33609,N_33552);
nor U33964 (N_33964,N_33543,N_33684);
and U33965 (N_33965,N_33569,N_33584);
nor U33966 (N_33966,N_33674,N_33616);
and U33967 (N_33967,N_33743,N_33503);
nor U33968 (N_33968,N_33728,N_33666);
or U33969 (N_33969,N_33545,N_33700);
nor U33970 (N_33970,N_33608,N_33574);
nor U33971 (N_33971,N_33514,N_33729);
nor U33972 (N_33972,N_33682,N_33743);
and U33973 (N_33973,N_33612,N_33707);
xor U33974 (N_33974,N_33705,N_33679);
nor U33975 (N_33975,N_33601,N_33504);
nand U33976 (N_33976,N_33628,N_33586);
nand U33977 (N_33977,N_33666,N_33580);
or U33978 (N_33978,N_33686,N_33723);
or U33979 (N_33979,N_33627,N_33551);
xnor U33980 (N_33980,N_33553,N_33533);
nor U33981 (N_33981,N_33677,N_33578);
or U33982 (N_33982,N_33596,N_33638);
nor U33983 (N_33983,N_33522,N_33621);
and U33984 (N_33984,N_33644,N_33574);
nor U33985 (N_33985,N_33650,N_33588);
nor U33986 (N_33986,N_33730,N_33635);
or U33987 (N_33987,N_33676,N_33721);
nor U33988 (N_33988,N_33538,N_33686);
nand U33989 (N_33989,N_33717,N_33739);
and U33990 (N_33990,N_33699,N_33695);
or U33991 (N_33991,N_33595,N_33604);
nor U33992 (N_33992,N_33575,N_33697);
nor U33993 (N_33993,N_33596,N_33608);
nor U33994 (N_33994,N_33663,N_33724);
xor U33995 (N_33995,N_33732,N_33601);
nand U33996 (N_33996,N_33714,N_33513);
nand U33997 (N_33997,N_33603,N_33660);
nor U33998 (N_33998,N_33629,N_33620);
xor U33999 (N_33999,N_33598,N_33698);
or U34000 (N_34000,N_33904,N_33877);
and U34001 (N_34001,N_33860,N_33823);
xnor U34002 (N_34002,N_33826,N_33899);
nor U34003 (N_34003,N_33893,N_33954);
or U34004 (N_34004,N_33952,N_33998);
and U34005 (N_34005,N_33829,N_33945);
nor U34006 (N_34006,N_33857,N_33780);
nand U34007 (N_34007,N_33787,N_33891);
nand U34008 (N_34008,N_33918,N_33966);
or U34009 (N_34009,N_33870,N_33751);
or U34010 (N_34010,N_33781,N_33789);
nor U34011 (N_34011,N_33873,N_33775);
xnor U34012 (N_34012,N_33889,N_33943);
nor U34013 (N_34013,N_33764,N_33782);
nand U34014 (N_34014,N_33793,N_33853);
and U34015 (N_34015,N_33810,N_33797);
or U34016 (N_34016,N_33993,N_33763);
nor U34017 (N_34017,N_33987,N_33822);
nor U34018 (N_34018,N_33800,N_33811);
xnor U34019 (N_34019,N_33921,N_33944);
and U34020 (N_34020,N_33843,N_33972);
or U34021 (N_34021,N_33957,N_33771);
xnor U34022 (N_34022,N_33942,N_33928);
or U34023 (N_34023,N_33869,N_33785);
or U34024 (N_34024,N_33828,N_33985);
nor U34025 (N_34025,N_33794,N_33802);
or U34026 (N_34026,N_33948,N_33849);
nor U34027 (N_34027,N_33755,N_33908);
xor U34028 (N_34028,N_33990,N_33871);
and U34029 (N_34029,N_33827,N_33799);
xor U34030 (N_34030,N_33769,N_33933);
xnor U34031 (N_34031,N_33892,N_33819);
or U34032 (N_34032,N_33890,N_33913);
xor U34033 (N_34033,N_33753,N_33880);
nor U34034 (N_34034,N_33754,N_33956);
xor U34035 (N_34035,N_33760,N_33920);
xnor U34036 (N_34036,N_33975,N_33861);
and U34037 (N_34037,N_33981,N_33852);
nor U34038 (N_34038,N_33984,N_33814);
or U34039 (N_34039,N_33784,N_33982);
nor U34040 (N_34040,N_33844,N_33919);
xnor U34041 (N_34041,N_33858,N_33806);
nand U34042 (N_34042,N_33922,N_33971);
or U34043 (N_34043,N_33974,N_33836);
and U34044 (N_34044,N_33947,N_33911);
nand U34045 (N_34045,N_33901,N_33856);
xor U34046 (N_34046,N_33900,N_33803);
nor U34047 (N_34047,N_33773,N_33986);
or U34048 (N_34048,N_33905,N_33847);
or U34049 (N_34049,N_33838,N_33850);
xnor U34050 (N_34050,N_33906,N_33968);
xor U34051 (N_34051,N_33996,N_33970);
or U34052 (N_34052,N_33995,N_33865);
or U34053 (N_34053,N_33795,N_33876);
nand U34054 (N_34054,N_33978,N_33770);
nand U34055 (N_34055,N_33756,N_33798);
nor U34056 (N_34056,N_33950,N_33766);
and U34057 (N_34057,N_33897,N_33909);
or U34058 (N_34058,N_33941,N_33851);
or U34059 (N_34059,N_33961,N_33896);
nand U34060 (N_34060,N_33834,N_33768);
or U34061 (N_34061,N_33772,N_33807);
nor U34062 (N_34062,N_33969,N_33820);
xor U34063 (N_34063,N_33809,N_33872);
and U34064 (N_34064,N_33959,N_33761);
or U34065 (N_34065,N_33832,N_33994);
or U34066 (N_34066,N_33779,N_33831);
xor U34067 (N_34067,N_33992,N_33980);
and U34068 (N_34068,N_33778,N_33878);
nor U34069 (N_34069,N_33859,N_33940);
and U34070 (N_34070,N_33946,N_33774);
or U34071 (N_34071,N_33884,N_33817);
nand U34072 (N_34072,N_33816,N_33841);
nand U34073 (N_34073,N_33818,N_33930);
or U34074 (N_34074,N_33805,N_33937);
or U34075 (N_34075,N_33757,N_33885);
xnor U34076 (N_34076,N_33791,N_33963);
xor U34077 (N_34077,N_33830,N_33962);
and U34078 (N_34078,N_33977,N_33912);
and U34079 (N_34079,N_33926,N_33935);
nor U34080 (N_34080,N_33997,N_33840);
nand U34081 (N_34081,N_33953,N_33855);
nand U34082 (N_34082,N_33894,N_33765);
nor U34083 (N_34083,N_33874,N_33750);
and U34084 (N_34084,N_33882,N_33932);
xnor U34085 (N_34085,N_33837,N_33898);
xor U34086 (N_34086,N_33783,N_33923);
or U34087 (N_34087,N_33936,N_33801);
nor U34088 (N_34088,N_33938,N_33999);
xor U34089 (N_34089,N_33910,N_33862);
and U34090 (N_34090,N_33960,N_33796);
or U34091 (N_34091,N_33839,N_33758);
xnor U34092 (N_34092,N_33907,N_33788);
xor U34093 (N_34093,N_33863,N_33914);
or U34094 (N_34094,N_33989,N_33752);
nand U34095 (N_34095,N_33762,N_33866);
nor U34096 (N_34096,N_33854,N_33888);
nand U34097 (N_34097,N_33777,N_33915);
nor U34098 (N_34098,N_33903,N_33845);
xor U34099 (N_34099,N_33808,N_33875);
and U34100 (N_34100,N_33902,N_33879);
nand U34101 (N_34101,N_33976,N_33759);
or U34102 (N_34102,N_33883,N_33867);
nand U34103 (N_34103,N_33934,N_33842);
xor U34104 (N_34104,N_33949,N_33886);
and U34105 (N_34105,N_33812,N_33917);
nor U34106 (N_34106,N_33835,N_33887);
xnor U34107 (N_34107,N_33821,N_33776);
or U34108 (N_34108,N_33881,N_33786);
or U34109 (N_34109,N_33958,N_33813);
xor U34110 (N_34110,N_33824,N_33815);
nand U34111 (N_34111,N_33925,N_33833);
nand U34112 (N_34112,N_33965,N_33973);
nor U34113 (N_34113,N_33964,N_33927);
nand U34114 (N_34114,N_33895,N_33955);
xor U34115 (N_34115,N_33951,N_33931);
xnor U34116 (N_34116,N_33967,N_33991);
xnor U34117 (N_34117,N_33804,N_33924);
nor U34118 (N_34118,N_33790,N_33825);
nand U34119 (N_34119,N_33916,N_33846);
nor U34120 (N_34120,N_33929,N_33983);
nor U34121 (N_34121,N_33868,N_33767);
or U34122 (N_34122,N_33792,N_33864);
nand U34123 (N_34123,N_33848,N_33988);
nand U34124 (N_34124,N_33939,N_33979);
nand U34125 (N_34125,N_33776,N_33797);
nand U34126 (N_34126,N_33810,N_33766);
and U34127 (N_34127,N_33996,N_33769);
and U34128 (N_34128,N_33789,N_33920);
xnor U34129 (N_34129,N_33919,N_33754);
nor U34130 (N_34130,N_33887,N_33994);
or U34131 (N_34131,N_33844,N_33965);
or U34132 (N_34132,N_33900,N_33972);
and U34133 (N_34133,N_33920,N_33772);
xor U34134 (N_34134,N_33952,N_33876);
nor U34135 (N_34135,N_33988,N_33928);
and U34136 (N_34136,N_33808,N_33864);
and U34137 (N_34137,N_33992,N_33775);
or U34138 (N_34138,N_33805,N_33902);
or U34139 (N_34139,N_33971,N_33972);
or U34140 (N_34140,N_33987,N_33957);
and U34141 (N_34141,N_33797,N_33878);
xor U34142 (N_34142,N_33940,N_33785);
xnor U34143 (N_34143,N_33764,N_33789);
xor U34144 (N_34144,N_33919,N_33895);
and U34145 (N_34145,N_33933,N_33785);
xor U34146 (N_34146,N_33845,N_33909);
or U34147 (N_34147,N_33794,N_33934);
and U34148 (N_34148,N_33920,N_33992);
nand U34149 (N_34149,N_33792,N_33775);
nor U34150 (N_34150,N_33847,N_33779);
and U34151 (N_34151,N_33947,N_33753);
xnor U34152 (N_34152,N_33856,N_33896);
nand U34153 (N_34153,N_33825,N_33787);
nor U34154 (N_34154,N_33837,N_33897);
or U34155 (N_34155,N_33939,N_33935);
and U34156 (N_34156,N_33765,N_33946);
nor U34157 (N_34157,N_33917,N_33753);
or U34158 (N_34158,N_33788,N_33831);
or U34159 (N_34159,N_33992,N_33753);
xnor U34160 (N_34160,N_33901,N_33923);
nor U34161 (N_34161,N_33968,N_33788);
xor U34162 (N_34162,N_33945,N_33751);
and U34163 (N_34163,N_33957,N_33895);
and U34164 (N_34164,N_33774,N_33892);
nand U34165 (N_34165,N_33803,N_33801);
xor U34166 (N_34166,N_33910,N_33909);
xor U34167 (N_34167,N_33764,N_33856);
nor U34168 (N_34168,N_33882,N_33858);
nand U34169 (N_34169,N_33772,N_33777);
xnor U34170 (N_34170,N_33805,N_33888);
nor U34171 (N_34171,N_33812,N_33753);
xor U34172 (N_34172,N_33852,N_33833);
and U34173 (N_34173,N_33793,N_33804);
nand U34174 (N_34174,N_33832,N_33778);
xor U34175 (N_34175,N_33820,N_33781);
xor U34176 (N_34176,N_33881,N_33860);
nand U34177 (N_34177,N_33788,N_33954);
or U34178 (N_34178,N_33834,N_33892);
nand U34179 (N_34179,N_33756,N_33831);
nand U34180 (N_34180,N_33789,N_33802);
or U34181 (N_34181,N_33966,N_33828);
xor U34182 (N_34182,N_33889,N_33891);
xor U34183 (N_34183,N_33759,N_33894);
nand U34184 (N_34184,N_33962,N_33898);
xor U34185 (N_34185,N_33822,N_33826);
or U34186 (N_34186,N_33921,N_33869);
nor U34187 (N_34187,N_33936,N_33816);
xnor U34188 (N_34188,N_33972,N_33799);
or U34189 (N_34189,N_33839,N_33885);
nand U34190 (N_34190,N_33984,N_33777);
nor U34191 (N_34191,N_33777,N_33798);
and U34192 (N_34192,N_33818,N_33778);
xnor U34193 (N_34193,N_33880,N_33815);
nor U34194 (N_34194,N_33829,N_33762);
nor U34195 (N_34195,N_33801,N_33921);
xnor U34196 (N_34196,N_33807,N_33858);
nand U34197 (N_34197,N_33753,N_33816);
nor U34198 (N_34198,N_33987,N_33960);
nand U34199 (N_34199,N_33772,N_33798);
nor U34200 (N_34200,N_33760,N_33874);
and U34201 (N_34201,N_33984,N_33857);
xor U34202 (N_34202,N_33762,N_33803);
or U34203 (N_34203,N_33810,N_33867);
and U34204 (N_34204,N_33831,N_33968);
nand U34205 (N_34205,N_33787,N_33813);
or U34206 (N_34206,N_33923,N_33773);
nand U34207 (N_34207,N_33781,N_33901);
nand U34208 (N_34208,N_33818,N_33884);
xnor U34209 (N_34209,N_33879,N_33952);
and U34210 (N_34210,N_33897,N_33980);
nand U34211 (N_34211,N_33933,N_33937);
nor U34212 (N_34212,N_33761,N_33914);
or U34213 (N_34213,N_33956,N_33821);
xnor U34214 (N_34214,N_33900,N_33949);
nor U34215 (N_34215,N_33753,N_33863);
nand U34216 (N_34216,N_33997,N_33832);
nor U34217 (N_34217,N_33972,N_33845);
nor U34218 (N_34218,N_33883,N_33835);
xor U34219 (N_34219,N_33842,N_33828);
xnor U34220 (N_34220,N_33876,N_33789);
nand U34221 (N_34221,N_33987,N_33770);
nand U34222 (N_34222,N_33963,N_33971);
and U34223 (N_34223,N_33973,N_33976);
and U34224 (N_34224,N_33808,N_33859);
nor U34225 (N_34225,N_33899,N_33841);
nor U34226 (N_34226,N_33793,N_33861);
and U34227 (N_34227,N_33870,N_33803);
nand U34228 (N_34228,N_33865,N_33855);
xor U34229 (N_34229,N_33806,N_33881);
nand U34230 (N_34230,N_33962,N_33802);
nor U34231 (N_34231,N_33848,N_33882);
nand U34232 (N_34232,N_33940,N_33769);
xor U34233 (N_34233,N_33965,N_33934);
xnor U34234 (N_34234,N_33978,N_33936);
xnor U34235 (N_34235,N_33927,N_33947);
nand U34236 (N_34236,N_33874,N_33895);
xnor U34237 (N_34237,N_33761,N_33872);
or U34238 (N_34238,N_33991,N_33989);
nor U34239 (N_34239,N_33970,N_33968);
nor U34240 (N_34240,N_33752,N_33955);
or U34241 (N_34241,N_33990,N_33914);
nand U34242 (N_34242,N_33759,N_33971);
or U34243 (N_34243,N_33759,N_33852);
xor U34244 (N_34244,N_33860,N_33825);
and U34245 (N_34245,N_33889,N_33772);
and U34246 (N_34246,N_33974,N_33782);
and U34247 (N_34247,N_33921,N_33772);
nand U34248 (N_34248,N_33856,N_33889);
xnor U34249 (N_34249,N_33778,N_33875);
xnor U34250 (N_34250,N_34005,N_34197);
nor U34251 (N_34251,N_34095,N_34156);
and U34252 (N_34252,N_34002,N_34089);
xnor U34253 (N_34253,N_34239,N_34078);
or U34254 (N_34254,N_34063,N_34111);
nor U34255 (N_34255,N_34218,N_34171);
or U34256 (N_34256,N_34195,N_34150);
nor U34257 (N_34257,N_34069,N_34140);
and U34258 (N_34258,N_34240,N_34099);
nand U34259 (N_34259,N_34247,N_34014);
nor U34260 (N_34260,N_34176,N_34248);
and U34261 (N_34261,N_34153,N_34003);
nor U34262 (N_34262,N_34203,N_34055);
and U34263 (N_34263,N_34161,N_34104);
nand U34264 (N_34264,N_34193,N_34225);
nor U34265 (N_34265,N_34024,N_34145);
or U34266 (N_34266,N_34213,N_34096);
and U34267 (N_34267,N_34148,N_34141);
or U34268 (N_34268,N_34102,N_34072);
xnor U34269 (N_34269,N_34129,N_34058);
and U34270 (N_34270,N_34092,N_34091);
or U34271 (N_34271,N_34036,N_34128);
or U34272 (N_34272,N_34194,N_34186);
xnor U34273 (N_34273,N_34031,N_34086);
nor U34274 (N_34274,N_34043,N_34184);
nor U34275 (N_34275,N_34162,N_34059);
or U34276 (N_34276,N_34076,N_34136);
nand U34277 (N_34277,N_34135,N_34023);
or U34278 (N_34278,N_34124,N_34066);
or U34279 (N_34279,N_34202,N_34125);
xor U34280 (N_34280,N_34115,N_34019);
nand U34281 (N_34281,N_34147,N_34052);
nand U34282 (N_34282,N_34109,N_34177);
nand U34283 (N_34283,N_34048,N_34214);
and U34284 (N_34284,N_34015,N_34167);
or U34285 (N_34285,N_34191,N_34057);
and U34286 (N_34286,N_34179,N_34042);
nand U34287 (N_34287,N_34119,N_34212);
or U34288 (N_34288,N_34082,N_34236);
xnor U34289 (N_34289,N_34081,N_34016);
xor U34290 (N_34290,N_34118,N_34073);
or U34291 (N_34291,N_34241,N_34209);
or U34292 (N_34292,N_34246,N_34056);
or U34293 (N_34293,N_34190,N_34219);
or U34294 (N_34294,N_34068,N_34245);
xnor U34295 (N_34295,N_34224,N_34093);
xor U34296 (N_34296,N_34106,N_34100);
xnor U34297 (N_34297,N_34229,N_34178);
and U34298 (N_34298,N_34210,N_34062);
nor U34299 (N_34299,N_34044,N_34080);
nand U34300 (N_34300,N_34130,N_34143);
or U34301 (N_34301,N_34011,N_34127);
or U34302 (N_34302,N_34030,N_34013);
nand U34303 (N_34303,N_34230,N_34049);
nand U34304 (N_34304,N_34039,N_34032);
nor U34305 (N_34305,N_34110,N_34154);
xnor U34306 (N_34306,N_34004,N_34198);
nor U34307 (N_34307,N_34164,N_34227);
nor U34308 (N_34308,N_34243,N_34001);
xnor U34309 (N_34309,N_34208,N_34009);
or U34310 (N_34310,N_34220,N_34216);
or U34311 (N_34311,N_34105,N_34211);
and U34312 (N_34312,N_34217,N_34025);
or U34313 (N_34313,N_34064,N_34079);
nand U34314 (N_34314,N_34183,N_34000);
and U34315 (N_34315,N_34007,N_34157);
xor U34316 (N_34316,N_34189,N_34114);
nor U34317 (N_34317,N_34122,N_34146);
and U34318 (N_34318,N_34235,N_34022);
xor U34319 (N_34319,N_34199,N_34149);
and U34320 (N_34320,N_34249,N_34181);
nor U34321 (N_34321,N_34006,N_34027);
or U34322 (N_34322,N_34012,N_34221);
nand U34323 (N_34323,N_34020,N_34166);
and U34324 (N_34324,N_34094,N_34170);
nand U34325 (N_34325,N_34168,N_34201);
nor U34326 (N_34326,N_34206,N_34126);
xnor U34327 (N_34327,N_34174,N_34173);
xnor U34328 (N_34328,N_34021,N_34101);
and U34329 (N_34329,N_34097,N_34215);
or U34330 (N_34330,N_34121,N_34008);
or U34331 (N_34331,N_34192,N_34165);
nand U34332 (N_34332,N_34244,N_34175);
and U34333 (N_34333,N_34108,N_34232);
or U34334 (N_34334,N_34222,N_34144);
nor U34335 (N_34335,N_34083,N_34163);
and U34336 (N_34336,N_34131,N_34137);
and U34337 (N_34337,N_34142,N_34053);
nand U34338 (N_34338,N_34017,N_34160);
or U34339 (N_34339,N_34234,N_34077);
or U34340 (N_34340,N_34204,N_34050);
xor U34341 (N_34341,N_34085,N_34098);
or U34342 (N_34342,N_34158,N_34026);
xor U34343 (N_34343,N_34196,N_34172);
nor U34344 (N_34344,N_34117,N_34112);
and U34345 (N_34345,N_34067,N_34065);
or U34346 (N_34346,N_34084,N_34238);
nor U34347 (N_34347,N_34038,N_34113);
and U34348 (N_34348,N_34226,N_34074);
or U34349 (N_34349,N_34034,N_34070);
and U34350 (N_34350,N_34123,N_34159);
nor U34351 (N_34351,N_34028,N_34120);
xor U34352 (N_34352,N_34046,N_34116);
xor U34353 (N_34353,N_34040,N_34187);
nor U34354 (N_34354,N_34205,N_34200);
xor U34355 (N_34355,N_34151,N_34045);
xnor U34356 (N_34356,N_34223,N_34075);
and U34357 (N_34357,N_34182,N_34061);
xor U34358 (N_34358,N_34233,N_34041);
or U34359 (N_34359,N_34231,N_34035);
xor U34360 (N_34360,N_34087,N_34010);
xnor U34361 (N_34361,N_34169,N_34037);
nand U34362 (N_34362,N_34155,N_34132);
nand U34363 (N_34363,N_34103,N_34188);
or U34364 (N_34364,N_34228,N_34185);
nand U34365 (N_34365,N_34051,N_34139);
nand U34366 (N_34366,N_34107,N_34138);
nand U34367 (N_34367,N_34134,N_34088);
xnor U34368 (N_34368,N_34152,N_34047);
xor U34369 (N_34369,N_34018,N_34242);
xor U34370 (N_34370,N_34133,N_34207);
and U34371 (N_34371,N_34054,N_34029);
and U34372 (N_34372,N_34071,N_34237);
nor U34373 (N_34373,N_34090,N_34060);
xnor U34374 (N_34374,N_34033,N_34180);
xnor U34375 (N_34375,N_34095,N_34215);
or U34376 (N_34376,N_34045,N_34098);
nor U34377 (N_34377,N_34209,N_34076);
nand U34378 (N_34378,N_34171,N_34197);
or U34379 (N_34379,N_34245,N_34005);
xnor U34380 (N_34380,N_34049,N_34235);
nand U34381 (N_34381,N_34050,N_34177);
or U34382 (N_34382,N_34150,N_34160);
or U34383 (N_34383,N_34240,N_34091);
xnor U34384 (N_34384,N_34084,N_34068);
xor U34385 (N_34385,N_34225,N_34207);
nor U34386 (N_34386,N_34051,N_34241);
xor U34387 (N_34387,N_34240,N_34102);
nor U34388 (N_34388,N_34063,N_34031);
nor U34389 (N_34389,N_34177,N_34111);
nor U34390 (N_34390,N_34022,N_34151);
or U34391 (N_34391,N_34147,N_34152);
or U34392 (N_34392,N_34239,N_34014);
and U34393 (N_34393,N_34087,N_34205);
and U34394 (N_34394,N_34160,N_34120);
nor U34395 (N_34395,N_34086,N_34112);
or U34396 (N_34396,N_34227,N_34221);
xnor U34397 (N_34397,N_34113,N_34058);
or U34398 (N_34398,N_34002,N_34056);
and U34399 (N_34399,N_34122,N_34104);
and U34400 (N_34400,N_34008,N_34142);
nor U34401 (N_34401,N_34168,N_34118);
nand U34402 (N_34402,N_34153,N_34050);
nand U34403 (N_34403,N_34229,N_34056);
nand U34404 (N_34404,N_34070,N_34011);
xor U34405 (N_34405,N_34127,N_34172);
and U34406 (N_34406,N_34153,N_34084);
or U34407 (N_34407,N_34078,N_34131);
nand U34408 (N_34408,N_34154,N_34043);
nand U34409 (N_34409,N_34011,N_34081);
or U34410 (N_34410,N_34114,N_34133);
nor U34411 (N_34411,N_34027,N_34075);
nor U34412 (N_34412,N_34142,N_34106);
xor U34413 (N_34413,N_34240,N_34113);
nor U34414 (N_34414,N_34089,N_34059);
or U34415 (N_34415,N_34208,N_34010);
or U34416 (N_34416,N_34181,N_34221);
nand U34417 (N_34417,N_34247,N_34060);
and U34418 (N_34418,N_34033,N_34249);
nor U34419 (N_34419,N_34148,N_34190);
xnor U34420 (N_34420,N_34031,N_34011);
nor U34421 (N_34421,N_34040,N_34103);
nand U34422 (N_34422,N_34224,N_34136);
and U34423 (N_34423,N_34057,N_34004);
nand U34424 (N_34424,N_34085,N_34062);
or U34425 (N_34425,N_34087,N_34069);
and U34426 (N_34426,N_34068,N_34022);
or U34427 (N_34427,N_34094,N_34205);
nor U34428 (N_34428,N_34173,N_34231);
nor U34429 (N_34429,N_34052,N_34005);
nor U34430 (N_34430,N_34157,N_34242);
nand U34431 (N_34431,N_34196,N_34074);
nand U34432 (N_34432,N_34000,N_34248);
xnor U34433 (N_34433,N_34026,N_34024);
xnor U34434 (N_34434,N_34226,N_34021);
nor U34435 (N_34435,N_34147,N_34011);
xnor U34436 (N_34436,N_34124,N_34228);
or U34437 (N_34437,N_34213,N_34116);
nor U34438 (N_34438,N_34196,N_34211);
and U34439 (N_34439,N_34193,N_34204);
xor U34440 (N_34440,N_34147,N_34234);
or U34441 (N_34441,N_34085,N_34232);
xor U34442 (N_34442,N_34056,N_34102);
nand U34443 (N_34443,N_34076,N_34096);
nor U34444 (N_34444,N_34145,N_34130);
nor U34445 (N_34445,N_34021,N_34081);
xnor U34446 (N_34446,N_34171,N_34240);
nand U34447 (N_34447,N_34160,N_34168);
xor U34448 (N_34448,N_34194,N_34035);
nor U34449 (N_34449,N_34038,N_34107);
nor U34450 (N_34450,N_34174,N_34212);
xnor U34451 (N_34451,N_34207,N_34148);
xnor U34452 (N_34452,N_34133,N_34091);
nor U34453 (N_34453,N_34100,N_34131);
and U34454 (N_34454,N_34168,N_34078);
and U34455 (N_34455,N_34027,N_34009);
nand U34456 (N_34456,N_34036,N_34108);
nand U34457 (N_34457,N_34132,N_34033);
nand U34458 (N_34458,N_34170,N_34070);
and U34459 (N_34459,N_34036,N_34065);
xnor U34460 (N_34460,N_34004,N_34026);
nand U34461 (N_34461,N_34012,N_34204);
nor U34462 (N_34462,N_34160,N_34095);
nor U34463 (N_34463,N_34191,N_34072);
nor U34464 (N_34464,N_34132,N_34240);
nor U34465 (N_34465,N_34167,N_34120);
or U34466 (N_34466,N_34012,N_34062);
nand U34467 (N_34467,N_34226,N_34071);
and U34468 (N_34468,N_34171,N_34228);
and U34469 (N_34469,N_34036,N_34056);
nand U34470 (N_34470,N_34235,N_34155);
or U34471 (N_34471,N_34067,N_34095);
and U34472 (N_34472,N_34156,N_34122);
xnor U34473 (N_34473,N_34054,N_34163);
nand U34474 (N_34474,N_34110,N_34239);
xor U34475 (N_34475,N_34241,N_34136);
or U34476 (N_34476,N_34239,N_34217);
and U34477 (N_34477,N_34088,N_34116);
nor U34478 (N_34478,N_34149,N_34140);
nor U34479 (N_34479,N_34100,N_34013);
nand U34480 (N_34480,N_34133,N_34198);
xnor U34481 (N_34481,N_34248,N_34170);
xnor U34482 (N_34482,N_34238,N_34043);
nand U34483 (N_34483,N_34083,N_34069);
and U34484 (N_34484,N_34186,N_34119);
and U34485 (N_34485,N_34121,N_34142);
nor U34486 (N_34486,N_34146,N_34226);
xor U34487 (N_34487,N_34183,N_34234);
and U34488 (N_34488,N_34033,N_34005);
nor U34489 (N_34489,N_34054,N_34189);
nand U34490 (N_34490,N_34009,N_34017);
xor U34491 (N_34491,N_34211,N_34054);
or U34492 (N_34492,N_34154,N_34217);
or U34493 (N_34493,N_34098,N_34166);
nand U34494 (N_34494,N_34054,N_34102);
nor U34495 (N_34495,N_34041,N_34091);
xnor U34496 (N_34496,N_34165,N_34137);
and U34497 (N_34497,N_34202,N_34222);
nor U34498 (N_34498,N_34059,N_34078);
xnor U34499 (N_34499,N_34149,N_34222);
xor U34500 (N_34500,N_34269,N_34487);
nor U34501 (N_34501,N_34424,N_34484);
xor U34502 (N_34502,N_34427,N_34360);
and U34503 (N_34503,N_34476,N_34290);
nor U34504 (N_34504,N_34363,N_34276);
nand U34505 (N_34505,N_34389,N_34382);
xnor U34506 (N_34506,N_34444,N_34282);
nor U34507 (N_34507,N_34456,N_34332);
and U34508 (N_34508,N_34357,N_34293);
nand U34509 (N_34509,N_34384,N_34458);
nand U34510 (N_34510,N_34469,N_34258);
xnor U34511 (N_34511,N_34305,N_34435);
xnor U34512 (N_34512,N_34297,N_34467);
nor U34513 (N_34513,N_34265,N_34472);
nand U34514 (N_34514,N_34474,N_34488);
or U34515 (N_34515,N_34272,N_34473);
and U34516 (N_34516,N_34404,N_34370);
and U34517 (N_34517,N_34314,N_34278);
nand U34518 (N_34518,N_34431,N_34356);
or U34519 (N_34519,N_34354,N_34273);
nand U34520 (N_34520,N_34257,N_34291);
nor U34521 (N_34521,N_34364,N_34387);
xnor U34522 (N_34522,N_34287,N_34274);
and U34523 (N_34523,N_34414,N_34288);
nand U34524 (N_34524,N_34317,N_34439);
or U34525 (N_34525,N_34409,N_34405);
xnor U34526 (N_34526,N_34490,N_34468);
xnor U34527 (N_34527,N_34253,N_34448);
or U34528 (N_34528,N_34461,N_34335);
nor U34529 (N_34529,N_34397,N_34412);
and U34530 (N_34530,N_34316,N_34355);
or U34531 (N_34531,N_34422,N_34496);
nor U34532 (N_34532,N_34313,N_34377);
nor U34533 (N_34533,N_34386,N_34462);
xor U34534 (N_34534,N_34491,N_34268);
xnor U34535 (N_34535,N_34263,N_34483);
and U34536 (N_34536,N_34307,N_34270);
xor U34537 (N_34537,N_34479,N_34441);
xnor U34538 (N_34538,N_34267,N_34380);
xor U34539 (N_34539,N_34406,N_34396);
nand U34540 (N_34540,N_34326,N_34275);
xnor U34541 (N_34541,N_34298,N_34450);
or U34542 (N_34542,N_34436,N_34336);
or U34543 (N_34543,N_34259,N_34320);
nand U34544 (N_34544,N_34499,N_34327);
or U34545 (N_34545,N_34334,N_34271);
nand U34546 (N_34546,N_34452,N_34383);
xor U34547 (N_34547,N_34369,N_34361);
nand U34548 (N_34548,N_34465,N_34433);
nand U34549 (N_34549,N_34296,N_34333);
nand U34550 (N_34550,N_34366,N_34261);
and U34551 (N_34551,N_34310,N_34493);
or U34552 (N_34552,N_34459,N_34300);
and U34553 (N_34553,N_34455,N_34285);
xor U34554 (N_34554,N_34342,N_34480);
xor U34555 (N_34555,N_34315,N_34475);
or U34556 (N_34556,N_34368,N_34250);
and U34557 (N_34557,N_34385,N_34277);
and U34558 (N_34558,N_34260,N_34324);
nand U34559 (N_34559,N_34308,N_34289);
nor U34560 (N_34560,N_34351,N_34413);
nand U34561 (N_34561,N_34379,N_34255);
nor U34562 (N_34562,N_34375,N_34466);
nand U34563 (N_34563,N_34254,N_34264);
xnor U34564 (N_34564,N_34348,N_34304);
or U34565 (N_34565,N_34292,N_34301);
nor U34566 (N_34566,N_34251,N_34295);
nor U34567 (N_34567,N_34319,N_34393);
and U34568 (N_34568,N_34343,N_34378);
or U34569 (N_34569,N_34279,N_34395);
nor U34570 (N_34570,N_34451,N_34376);
and U34571 (N_34571,N_34339,N_34399);
and U34572 (N_34572,N_34374,N_34373);
nor U34573 (N_34573,N_34391,N_34471);
xnor U34574 (N_34574,N_34392,N_34464);
or U34575 (N_34575,N_34495,N_34252);
nor U34576 (N_34576,N_34485,N_34447);
nor U34577 (N_34577,N_34437,N_34494);
xor U34578 (N_34578,N_34489,N_34421);
nor U34579 (N_34579,N_34434,N_34286);
and U34580 (N_34580,N_34284,N_34345);
nor U34581 (N_34581,N_34331,N_34478);
nor U34582 (N_34582,N_34438,N_34430);
nand U34583 (N_34583,N_34470,N_34415);
nand U34584 (N_34584,N_34417,N_34486);
xnor U34585 (N_34585,N_34394,N_34429);
nand U34586 (N_34586,N_34381,N_34463);
xor U34587 (N_34587,N_34482,N_34453);
and U34588 (N_34588,N_34322,N_34410);
and U34589 (N_34589,N_34403,N_34426);
xnor U34590 (N_34590,N_34311,N_34371);
or U34591 (N_34591,N_34408,N_34325);
and U34592 (N_34592,N_34323,N_34498);
or U34593 (N_34593,N_34388,N_34497);
nor U34594 (N_34594,N_34338,N_34349);
nand U34595 (N_34595,N_34347,N_34367);
and U34596 (N_34596,N_34362,N_34337);
and U34597 (N_34597,N_34280,N_34477);
nor U34598 (N_34598,N_34318,N_34390);
or U34599 (N_34599,N_34423,N_34442);
xnor U34600 (N_34600,N_34402,N_34481);
nand U34601 (N_34601,N_34341,N_34346);
nor U34602 (N_34602,N_34359,N_34294);
nand U34603 (N_34603,N_34266,N_34330);
or U34604 (N_34604,N_34365,N_34401);
and U34605 (N_34605,N_34328,N_34353);
and U34606 (N_34606,N_34309,N_34350);
and U34607 (N_34607,N_34321,N_34457);
nand U34608 (N_34608,N_34418,N_34440);
or U34609 (N_34609,N_34398,N_34358);
xor U34610 (N_34610,N_34419,N_34446);
or U34611 (N_34611,N_34256,N_34449);
and U34612 (N_34612,N_34428,N_34262);
xnor U34613 (N_34613,N_34416,N_34340);
or U34614 (N_34614,N_34460,N_34411);
and U34615 (N_34615,N_34400,N_34432);
or U34616 (N_34616,N_34372,N_34407);
nor U34617 (N_34617,N_34302,N_34344);
or U34618 (N_34618,N_34306,N_34454);
and U34619 (N_34619,N_34303,N_34283);
nor U34620 (N_34620,N_34299,N_34425);
xor U34621 (N_34621,N_34443,N_34329);
xnor U34622 (N_34622,N_34420,N_34492);
and U34623 (N_34623,N_34445,N_34352);
and U34624 (N_34624,N_34312,N_34281);
and U34625 (N_34625,N_34488,N_34290);
nand U34626 (N_34626,N_34349,N_34321);
or U34627 (N_34627,N_34334,N_34466);
xor U34628 (N_34628,N_34302,N_34294);
nand U34629 (N_34629,N_34322,N_34285);
and U34630 (N_34630,N_34296,N_34287);
or U34631 (N_34631,N_34459,N_34411);
or U34632 (N_34632,N_34325,N_34328);
and U34633 (N_34633,N_34386,N_34436);
or U34634 (N_34634,N_34336,N_34306);
nor U34635 (N_34635,N_34359,N_34415);
nor U34636 (N_34636,N_34360,N_34291);
nand U34637 (N_34637,N_34433,N_34280);
nor U34638 (N_34638,N_34347,N_34366);
nor U34639 (N_34639,N_34402,N_34413);
and U34640 (N_34640,N_34419,N_34327);
xor U34641 (N_34641,N_34267,N_34426);
xnor U34642 (N_34642,N_34479,N_34355);
and U34643 (N_34643,N_34382,N_34278);
or U34644 (N_34644,N_34305,N_34370);
nor U34645 (N_34645,N_34299,N_34484);
and U34646 (N_34646,N_34358,N_34282);
and U34647 (N_34647,N_34289,N_34390);
nor U34648 (N_34648,N_34418,N_34454);
or U34649 (N_34649,N_34403,N_34437);
nor U34650 (N_34650,N_34287,N_34279);
or U34651 (N_34651,N_34431,N_34273);
xor U34652 (N_34652,N_34488,N_34417);
xor U34653 (N_34653,N_34290,N_34397);
nor U34654 (N_34654,N_34454,N_34489);
or U34655 (N_34655,N_34356,N_34415);
xnor U34656 (N_34656,N_34362,N_34360);
nand U34657 (N_34657,N_34390,N_34401);
or U34658 (N_34658,N_34427,N_34391);
nor U34659 (N_34659,N_34422,N_34275);
or U34660 (N_34660,N_34364,N_34488);
and U34661 (N_34661,N_34295,N_34276);
nor U34662 (N_34662,N_34406,N_34479);
nor U34663 (N_34663,N_34309,N_34472);
or U34664 (N_34664,N_34488,N_34399);
nor U34665 (N_34665,N_34476,N_34307);
xnor U34666 (N_34666,N_34263,N_34352);
and U34667 (N_34667,N_34396,N_34262);
nand U34668 (N_34668,N_34476,N_34423);
nand U34669 (N_34669,N_34490,N_34345);
nand U34670 (N_34670,N_34390,N_34443);
and U34671 (N_34671,N_34316,N_34363);
xnor U34672 (N_34672,N_34301,N_34465);
and U34673 (N_34673,N_34328,N_34484);
nor U34674 (N_34674,N_34393,N_34453);
nor U34675 (N_34675,N_34419,N_34401);
nand U34676 (N_34676,N_34324,N_34286);
or U34677 (N_34677,N_34362,N_34487);
nand U34678 (N_34678,N_34314,N_34268);
nor U34679 (N_34679,N_34295,N_34339);
and U34680 (N_34680,N_34275,N_34269);
or U34681 (N_34681,N_34389,N_34359);
or U34682 (N_34682,N_34468,N_34434);
xnor U34683 (N_34683,N_34261,N_34316);
nor U34684 (N_34684,N_34456,N_34434);
nor U34685 (N_34685,N_34499,N_34390);
or U34686 (N_34686,N_34417,N_34362);
nor U34687 (N_34687,N_34316,N_34351);
nor U34688 (N_34688,N_34387,N_34360);
and U34689 (N_34689,N_34379,N_34498);
or U34690 (N_34690,N_34463,N_34404);
and U34691 (N_34691,N_34387,N_34282);
xnor U34692 (N_34692,N_34260,N_34342);
nand U34693 (N_34693,N_34336,N_34450);
nor U34694 (N_34694,N_34317,N_34354);
nor U34695 (N_34695,N_34487,N_34364);
nand U34696 (N_34696,N_34387,N_34482);
nor U34697 (N_34697,N_34372,N_34411);
xnor U34698 (N_34698,N_34456,N_34489);
nand U34699 (N_34699,N_34346,N_34355);
nor U34700 (N_34700,N_34365,N_34371);
and U34701 (N_34701,N_34458,N_34427);
nand U34702 (N_34702,N_34437,N_34295);
nor U34703 (N_34703,N_34299,N_34373);
nand U34704 (N_34704,N_34467,N_34295);
nor U34705 (N_34705,N_34407,N_34468);
and U34706 (N_34706,N_34450,N_34473);
or U34707 (N_34707,N_34314,N_34370);
nor U34708 (N_34708,N_34432,N_34433);
and U34709 (N_34709,N_34499,N_34368);
nand U34710 (N_34710,N_34353,N_34417);
xor U34711 (N_34711,N_34355,N_34487);
nand U34712 (N_34712,N_34296,N_34423);
nor U34713 (N_34713,N_34434,N_34264);
nand U34714 (N_34714,N_34466,N_34474);
nand U34715 (N_34715,N_34477,N_34490);
or U34716 (N_34716,N_34475,N_34456);
nor U34717 (N_34717,N_34387,N_34278);
or U34718 (N_34718,N_34403,N_34417);
xor U34719 (N_34719,N_34284,N_34266);
nand U34720 (N_34720,N_34312,N_34280);
nor U34721 (N_34721,N_34295,N_34454);
or U34722 (N_34722,N_34494,N_34473);
and U34723 (N_34723,N_34259,N_34458);
nand U34724 (N_34724,N_34429,N_34452);
and U34725 (N_34725,N_34459,N_34305);
xnor U34726 (N_34726,N_34388,N_34465);
and U34727 (N_34727,N_34447,N_34369);
or U34728 (N_34728,N_34393,N_34448);
or U34729 (N_34729,N_34329,N_34435);
nor U34730 (N_34730,N_34369,N_34434);
and U34731 (N_34731,N_34271,N_34437);
and U34732 (N_34732,N_34453,N_34399);
xor U34733 (N_34733,N_34279,N_34344);
nor U34734 (N_34734,N_34411,N_34497);
and U34735 (N_34735,N_34259,N_34416);
xor U34736 (N_34736,N_34357,N_34274);
nand U34737 (N_34737,N_34420,N_34491);
xor U34738 (N_34738,N_34358,N_34423);
nand U34739 (N_34739,N_34255,N_34455);
nor U34740 (N_34740,N_34439,N_34466);
and U34741 (N_34741,N_34405,N_34343);
nor U34742 (N_34742,N_34314,N_34495);
and U34743 (N_34743,N_34452,N_34409);
nor U34744 (N_34744,N_34409,N_34475);
xor U34745 (N_34745,N_34335,N_34312);
nor U34746 (N_34746,N_34476,N_34455);
nor U34747 (N_34747,N_34424,N_34402);
nand U34748 (N_34748,N_34257,N_34477);
or U34749 (N_34749,N_34336,N_34317);
xor U34750 (N_34750,N_34648,N_34518);
xnor U34751 (N_34751,N_34535,N_34561);
nor U34752 (N_34752,N_34671,N_34724);
nor U34753 (N_34753,N_34629,N_34602);
and U34754 (N_34754,N_34734,N_34720);
nor U34755 (N_34755,N_34547,N_34745);
xor U34756 (N_34756,N_34549,N_34557);
xor U34757 (N_34757,N_34637,N_34598);
or U34758 (N_34758,N_34626,N_34636);
or U34759 (N_34759,N_34522,N_34566);
nor U34760 (N_34760,N_34688,N_34613);
nand U34761 (N_34761,N_34612,N_34558);
nand U34762 (N_34762,N_34645,N_34502);
nor U34763 (N_34763,N_34619,N_34701);
xnor U34764 (N_34764,N_34530,N_34615);
and U34765 (N_34765,N_34593,N_34512);
and U34766 (N_34766,N_34507,N_34742);
nor U34767 (N_34767,N_34555,N_34526);
nand U34768 (N_34768,N_34737,N_34616);
nand U34769 (N_34769,N_34610,N_34622);
nor U34770 (N_34770,N_34633,N_34659);
xnor U34771 (N_34771,N_34591,N_34652);
nand U34772 (N_34772,N_34592,N_34571);
xnor U34773 (N_34773,N_34679,N_34509);
nand U34774 (N_34774,N_34513,N_34623);
xor U34775 (N_34775,N_34542,N_34572);
and U34776 (N_34776,N_34657,N_34505);
nor U34777 (N_34777,N_34560,N_34698);
xnor U34778 (N_34778,N_34503,N_34638);
nand U34779 (N_34779,N_34641,N_34736);
nor U34780 (N_34780,N_34672,N_34706);
or U34781 (N_34781,N_34600,N_34650);
nand U34782 (N_34782,N_34697,N_34634);
nor U34783 (N_34783,N_34563,N_34614);
nor U34784 (N_34784,N_34670,N_34725);
xnor U34785 (N_34785,N_34527,N_34709);
xnor U34786 (N_34786,N_34677,N_34694);
and U34787 (N_34787,N_34746,N_34573);
xor U34788 (N_34788,N_34531,N_34544);
nand U34789 (N_34789,N_34601,N_34730);
and U34790 (N_34790,N_34689,N_34747);
or U34791 (N_34791,N_34727,N_34577);
nor U34792 (N_34792,N_34569,N_34665);
nand U34793 (N_34793,N_34738,N_34647);
nand U34794 (N_34794,N_34556,N_34643);
xnor U34795 (N_34795,N_34667,N_34539);
or U34796 (N_34796,N_34704,N_34587);
and U34797 (N_34797,N_34562,N_34553);
xnor U34798 (N_34798,N_34675,N_34682);
nor U34799 (N_34799,N_34673,N_34708);
nand U34800 (N_34800,N_34597,N_34695);
nor U34801 (N_34801,N_34590,N_34584);
and U34802 (N_34802,N_34570,N_34550);
or U34803 (N_34803,N_34632,N_34525);
and U34804 (N_34804,N_34664,N_34705);
nor U34805 (N_34805,N_34683,N_34583);
nand U34806 (N_34806,N_34674,N_34735);
or U34807 (N_34807,N_34702,N_34565);
xnor U34808 (N_34808,N_34710,N_34718);
and U34809 (N_34809,N_34743,N_34656);
xor U34810 (N_34810,N_34548,N_34536);
or U34811 (N_34811,N_34580,N_34511);
and U34812 (N_34812,N_34715,N_34608);
xor U34813 (N_34813,N_34521,N_34520);
nand U34814 (N_34814,N_34681,N_34533);
nor U34815 (N_34815,N_34690,N_34582);
or U34816 (N_34816,N_34728,N_34546);
nand U34817 (N_34817,N_34635,N_34604);
and U34818 (N_34818,N_34740,N_34581);
nand U34819 (N_34819,N_34739,N_34712);
xnor U34820 (N_34820,N_34621,N_34524);
or U34821 (N_34821,N_34574,N_34567);
nand U34822 (N_34822,N_34551,N_34676);
and U34823 (N_34823,N_34501,N_34646);
nand U34824 (N_34824,N_34504,N_34627);
nand U34825 (N_34825,N_34661,N_34532);
nor U34826 (N_34826,N_34585,N_34660);
nand U34827 (N_34827,N_34651,N_34552);
nand U34828 (N_34828,N_34721,N_34628);
and U34829 (N_34829,N_34700,N_34617);
xnor U34830 (N_34830,N_34696,N_34655);
nand U34831 (N_34831,N_34537,N_34625);
or U34832 (N_34832,N_34603,N_34576);
and U34833 (N_34833,N_34639,N_34516);
and U34834 (N_34834,N_34642,N_34618);
and U34835 (N_34835,N_34506,N_34631);
or U34836 (N_34836,N_34515,N_34540);
nor U34837 (N_34837,N_34510,N_34594);
or U34838 (N_34838,N_34579,N_34686);
nand U34839 (N_34839,N_34630,N_34719);
or U34840 (N_34840,N_34691,N_34749);
xnor U34841 (N_34841,N_34589,N_34620);
or U34842 (N_34842,N_34568,N_34529);
nor U34843 (N_34843,N_34519,N_34722);
nor U34844 (N_34844,N_34692,N_34733);
nor U34845 (N_34845,N_34599,N_34644);
or U34846 (N_34846,N_34663,N_34731);
nor U34847 (N_34847,N_34523,N_34609);
or U34848 (N_34848,N_34554,N_34596);
nor U34849 (N_34849,N_34559,N_34748);
and U34850 (N_34850,N_34564,N_34543);
xnor U34851 (N_34851,N_34726,N_34732);
and U34852 (N_34852,N_34541,N_34624);
or U34853 (N_34853,N_34528,N_34680);
and U34854 (N_34854,N_34666,N_34703);
and U34855 (N_34855,N_34741,N_34668);
nor U34856 (N_34856,N_34729,N_34693);
nor U34857 (N_34857,N_34606,N_34699);
or U34858 (N_34858,N_34713,N_34744);
and U34859 (N_34859,N_34687,N_34716);
or U34860 (N_34860,N_34723,N_34611);
nor U34861 (N_34861,N_34654,N_34607);
nand U34862 (N_34862,N_34707,N_34500);
nor U34863 (N_34863,N_34640,N_34595);
and U34864 (N_34864,N_34649,N_34714);
nor U34865 (N_34865,N_34534,N_34578);
nand U34866 (N_34866,N_34517,N_34586);
nor U34867 (N_34867,N_34658,N_34514);
or U34868 (N_34868,N_34662,N_34711);
xnor U34869 (N_34869,N_34508,N_34575);
and U34870 (N_34870,N_34669,N_34588);
nand U34871 (N_34871,N_34685,N_34717);
nand U34872 (N_34872,N_34678,N_34538);
nor U34873 (N_34873,N_34605,N_34653);
nor U34874 (N_34874,N_34684,N_34545);
or U34875 (N_34875,N_34650,N_34715);
and U34876 (N_34876,N_34687,N_34724);
or U34877 (N_34877,N_34729,N_34684);
nand U34878 (N_34878,N_34566,N_34651);
nor U34879 (N_34879,N_34608,N_34618);
and U34880 (N_34880,N_34605,N_34641);
nand U34881 (N_34881,N_34671,N_34638);
nor U34882 (N_34882,N_34663,N_34630);
nand U34883 (N_34883,N_34634,N_34616);
nor U34884 (N_34884,N_34608,N_34695);
nand U34885 (N_34885,N_34613,N_34719);
xor U34886 (N_34886,N_34664,N_34639);
nand U34887 (N_34887,N_34511,N_34521);
xor U34888 (N_34888,N_34749,N_34505);
and U34889 (N_34889,N_34704,N_34674);
nor U34890 (N_34890,N_34554,N_34581);
and U34891 (N_34891,N_34569,N_34593);
and U34892 (N_34892,N_34649,N_34531);
xor U34893 (N_34893,N_34691,N_34747);
or U34894 (N_34894,N_34505,N_34695);
or U34895 (N_34895,N_34533,N_34514);
and U34896 (N_34896,N_34637,N_34557);
or U34897 (N_34897,N_34739,N_34741);
nor U34898 (N_34898,N_34663,N_34714);
or U34899 (N_34899,N_34527,N_34661);
and U34900 (N_34900,N_34641,N_34572);
nor U34901 (N_34901,N_34541,N_34583);
or U34902 (N_34902,N_34524,N_34737);
xnor U34903 (N_34903,N_34694,N_34637);
nor U34904 (N_34904,N_34552,N_34657);
or U34905 (N_34905,N_34597,N_34738);
and U34906 (N_34906,N_34686,N_34615);
xnor U34907 (N_34907,N_34619,N_34722);
and U34908 (N_34908,N_34643,N_34617);
and U34909 (N_34909,N_34731,N_34510);
or U34910 (N_34910,N_34647,N_34603);
nand U34911 (N_34911,N_34724,N_34563);
and U34912 (N_34912,N_34718,N_34682);
and U34913 (N_34913,N_34570,N_34574);
xnor U34914 (N_34914,N_34723,N_34733);
or U34915 (N_34915,N_34736,N_34659);
nand U34916 (N_34916,N_34619,N_34628);
and U34917 (N_34917,N_34728,N_34731);
nor U34918 (N_34918,N_34502,N_34651);
nor U34919 (N_34919,N_34529,N_34717);
xnor U34920 (N_34920,N_34560,N_34574);
xnor U34921 (N_34921,N_34732,N_34645);
nor U34922 (N_34922,N_34685,N_34714);
and U34923 (N_34923,N_34616,N_34524);
nand U34924 (N_34924,N_34524,N_34665);
or U34925 (N_34925,N_34549,N_34511);
xnor U34926 (N_34926,N_34664,N_34523);
nand U34927 (N_34927,N_34723,N_34688);
nand U34928 (N_34928,N_34604,N_34520);
nor U34929 (N_34929,N_34524,N_34710);
nor U34930 (N_34930,N_34714,N_34743);
nand U34931 (N_34931,N_34631,N_34733);
nand U34932 (N_34932,N_34610,N_34690);
or U34933 (N_34933,N_34576,N_34640);
or U34934 (N_34934,N_34603,N_34542);
xnor U34935 (N_34935,N_34621,N_34668);
xor U34936 (N_34936,N_34537,N_34575);
xnor U34937 (N_34937,N_34534,N_34543);
nor U34938 (N_34938,N_34551,N_34682);
or U34939 (N_34939,N_34546,N_34705);
and U34940 (N_34940,N_34668,N_34697);
nand U34941 (N_34941,N_34559,N_34727);
or U34942 (N_34942,N_34701,N_34682);
or U34943 (N_34943,N_34526,N_34603);
xor U34944 (N_34944,N_34706,N_34598);
xnor U34945 (N_34945,N_34670,N_34612);
or U34946 (N_34946,N_34609,N_34531);
nand U34947 (N_34947,N_34628,N_34625);
and U34948 (N_34948,N_34510,N_34635);
or U34949 (N_34949,N_34693,N_34556);
nand U34950 (N_34950,N_34731,N_34532);
and U34951 (N_34951,N_34675,N_34522);
and U34952 (N_34952,N_34702,N_34632);
nor U34953 (N_34953,N_34550,N_34691);
and U34954 (N_34954,N_34688,N_34712);
nor U34955 (N_34955,N_34642,N_34698);
and U34956 (N_34956,N_34728,N_34634);
or U34957 (N_34957,N_34723,N_34555);
nor U34958 (N_34958,N_34692,N_34517);
or U34959 (N_34959,N_34605,N_34527);
or U34960 (N_34960,N_34660,N_34561);
or U34961 (N_34961,N_34552,N_34532);
nand U34962 (N_34962,N_34596,N_34744);
xnor U34963 (N_34963,N_34725,N_34642);
or U34964 (N_34964,N_34717,N_34522);
and U34965 (N_34965,N_34584,N_34610);
or U34966 (N_34966,N_34628,N_34678);
and U34967 (N_34967,N_34591,N_34678);
or U34968 (N_34968,N_34557,N_34517);
and U34969 (N_34969,N_34578,N_34709);
nor U34970 (N_34970,N_34584,N_34536);
xnor U34971 (N_34971,N_34743,N_34612);
or U34972 (N_34972,N_34620,N_34608);
nand U34973 (N_34973,N_34501,N_34564);
xor U34974 (N_34974,N_34674,N_34649);
xnor U34975 (N_34975,N_34580,N_34659);
xnor U34976 (N_34976,N_34680,N_34685);
xor U34977 (N_34977,N_34672,N_34722);
or U34978 (N_34978,N_34563,N_34645);
or U34979 (N_34979,N_34705,N_34736);
nand U34980 (N_34980,N_34696,N_34737);
nor U34981 (N_34981,N_34515,N_34587);
and U34982 (N_34982,N_34743,N_34690);
or U34983 (N_34983,N_34669,N_34571);
nor U34984 (N_34984,N_34733,N_34725);
or U34985 (N_34985,N_34583,N_34657);
or U34986 (N_34986,N_34588,N_34665);
nand U34987 (N_34987,N_34548,N_34745);
or U34988 (N_34988,N_34602,N_34700);
xor U34989 (N_34989,N_34550,N_34552);
and U34990 (N_34990,N_34663,N_34547);
xnor U34991 (N_34991,N_34647,N_34601);
nand U34992 (N_34992,N_34672,N_34619);
and U34993 (N_34993,N_34627,N_34611);
xor U34994 (N_34994,N_34511,N_34612);
nor U34995 (N_34995,N_34501,N_34507);
nand U34996 (N_34996,N_34633,N_34668);
nor U34997 (N_34997,N_34746,N_34602);
or U34998 (N_34998,N_34625,N_34585);
nor U34999 (N_34999,N_34715,N_34691);
xnor U35000 (N_35000,N_34803,N_34955);
and U35001 (N_35001,N_34976,N_34995);
xor U35002 (N_35002,N_34936,N_34792);
or U35003 (N_35003,N_34941,N_34895);
nand U35004 (N_35004,N_34877,N_34813);
nor U35005 (N_35005,N_34844,N_34853);
nor U35006 (N_35006,N_34908,N_34916);
nand U35007 (N_35007,N_34885,N_34979);
xor U35008 (N_35008,N_34759,N_34760);
and U35009 (N_35009,N_34915,N_34876);
or U35010 (N_35010,N_34870,N_34778);
nand U35011 (N_35011,N_34871,N_34882);
nand U35012 (N_35012,N_34851,N_34774);
xor U35013 (N_35013,N_34761,N_34904);
nor U35014 (N_35014,N_34926,N_34999);
or U35015 (N_35015,N_34994,N_34951);
or U35016 (N_35016,N_34767,N_34900);
xnor U35017 (N_35017,N_34850,N_34873);
nor U35018 (N_35018,N_34776,N_34939);
and U35019 (N_35019,N_34790,N_34791);
xnor U35020 (N_35020,N_34865,N_34913);
or U35021 (N_35021,N_34785,N_34883);
nor U35022 (N_35022,N_34835,N_34808);
or U35023 (N_35023,N_34780,N_34875);
or U35024 (N_35024,N_34831,N_34910);
xor U35025 (N_35025,N_34897,N_34920);
xnor U35026 (N_35026,N_34912,N_34830);
nand U35027 (N_35027,N_34923,N_34846);
xnor U35028 (N_35028,N_34942,N_34860);
and U35029 (N_35029,N_34927,N_34931);
xnor U35030 (N_35030,N_34948,N_34845);
xor U35031 (N_35031,N_34949,N_34932);
nand U35032 (N_35032,N_34985,N_34903);
nand U35033 (N_35033,N_34751,N_34818);
xnor U35034 (N_35034,N_34811,N_34757);
and U35035 (N_35035,N_34919,N_34809);
xor U35036 (N_35036,N_34820,N_34991);
or U35037 (N_35037,N_34821,N_34967);
nand U35038 (N_35038,N_34977,N_34914);
and U35039 (N_35039,N_34950,N_34905);
nand U35040 (N_35040,N_34944,N_34802);
nor U35041 (N_35041,N_34956,N_34772);
nand U35042 (N_35042,N_34928,N_34793);
xnor U35043 (N_35043,N_34962,N_34963);
and U35044 (N_35044,N_34783,N_34843);
xnor U35045 (N_35045,N_34828,N_34922);
nor U35046 (N_35046,N_34887,N_34837);
nor U35047 (N_35047,N_34989,N_34960);
nor U35048 (N_35048,N_34798,N_34833);
nor U35049 (N_35049,N_34947,N_34959);
xor U35050 (N_35050,N_34954,N_34771);
nor U35051 (N_35051,N_34825,N_34917);
and U35052 (N_35052,N_34909,N_34864);
nand U35053 (N_35053,N_34766,N_34874);
xnor U35054 (N_35054,N_34840,N_34980);
or U35055 (N_35055,N_34769,N_34834);
xnor U35056 (N_35056,N_34801,N_34805);
and U35057 (N_35057,N_34894,N_34987);
or U35058 (N_35058,N_34911,N_34896);
or U35059 (N_35059,N_34964,N_34898);
or U35060 (N_35060,N_34770,N_34777);
xnor U35061 (N_35061,N_34943,N_34918);
nor U35062 (N_35062,N_34815,N_34849);
xnor U35063 (N_35063,N_34861,N_34969);
nor U35064 (N_35064,N_34878,N_34879);
nand U35065 (N_35065,N_34762,N_34816);
and U35066 (N_35066,N_34988,N_34930);
or U35067 (N_35067,N_34938,N_34996);
nor U35068 (N_35068,N_34775,N_34993);
xnor U35069 (N_35069,N_34836,N_34997);
nor U35070 (N_35070,N_34990,N_34856);
or U35071 (N_35071,N_34984,N_34901);
xor U35072 (N_35072,N_34992,N_34817);
xor U35073 (N_35073,N_34839,N_34953);
or U35074 (N_35074,N_34924,N_34972);
and U35075 (N_35075,N_34807,N_34786);
or U35076 (N_35076,N_34841,N_34934);
nor U35077 (N_35077,N_34812,N_34892);
xor U35078 (N_35078,N_34804,N_34750);
nand U35079 (N_35079,N_34952,N_34797);
nor U35080 (N_35080,N_34862,N_34970);
or U35081 (N_35081,N_34796,N_34899);
nor U35082 (N_35082,N_34753,N_34935);
nor U35083 (N_35083,N_34819,N_34961);
nor U35084 (N_35084,N_34787,N_34906);
nor U35085 (N_35085,N_34966,N_34789);
nor U35086 (N_35086,N_34857,N_34978);
and U35087 (N_35087,N_34823,N_34784);
nand U35088 (N_35088,N_34758,N_34756);
and U35089 (N_35089,N_34824,N_34880);
or U35090 (N_35090,N_34814,N_34854);
or U35091 (N_35091,N_34763,N_34795);
nor U35092 (N_35092,N_34869,N_34794);
or U35093 (N_35093,N_34902,N_34937);
xnor U35094 (N_35094,N_34881,N_34838);
or U35095 (N_35095,N_34889,N_34781);
or U35096 (N_35096,N_34884,N_34982);
xor U35097 (N_35097,N_34921,N_34764);
and U35098 (N_35098,N_34810,N_34755);
nand U35099 (N_35099,N_34765,N_34933);
nand U35100 (N_35100,N_34940,N_34806);
nor U35101 (N_35101,N_34852,N_34858);
xor U35102 (N_35102,N_34773,N_34973);
and U35103 (N_35103,N_34829,N_34832);
xor U35104 (N_35104,N_34888,N_34891);
nor U35105 (N_35105,N_34957,N_34975);
xnor U35106 (N_35106,N_34752,N_34863);
or U35107 (N_35107,N_34800,N_34827);
nor U35108 (N_35108,N_34946,N_34782);
nor U35109 (N_35109,N_34998,N_34907);
nand U35110 (N_35110,N_34754,N_34981);
nor U35111 (N_35111,N_34866,N_34855);
nor U35112 (N_35112,N_34868,N_34822);
and U35113 (N_35113,N_34826,N_34890);
or U35114 (N_35114,N_34799,N_34886);
nand U35115 (N_35115,N_34965,N_34925);
xor U35116 (N_35116,N_34842,N_34929);
and U35117 (N_35117,N_34945,N_34788);
and U35118 (N_35118,N_34968,N_34872);
xor U35119 (N_35119,N_34779,N_34867);
and U35120 (N_35120,N_34983,N_34958);
nand U35121 (N_35121,N_34848,N_34859);
xor U35122 (N_35122,N_34986,N_34971);
or U35123 (N_35123,N_34974,N_34768);
nor U35124 (N_35124,N_34893,N_34847);
and U35125 (N_35125,N_34902,N_34914);
or U35126 (N_35126,N_34978,N_34967);
nor U35127 (N_35127,N_34938,N_34966);
nand U35128 (N_35128,N_34865,N_34751);
nand U35129 (N_35129,N_34997,N_34894);
nand U35130 (N_35130,N_34790,N_34946);
or U35131 (N_35131,N_34952,N_34884);
xor U35132 (N_35132,N_34947,N_34890);
and U35133 (N_35133,N_34970,N_34930);
or U35134 (N_35134,N_34855,N_34979);
or U35135 (N_35135,N_34922,N_34822);
or U35136 (N_35136,N_34750,N_34908);
and U35137 (N_35137,N_34973,N_34946);
nand U35138 (N_35138,N_34989,N_34967);
and U35139 (N_35139,N_34963,N_34922);
nand U35140 (N_35140,N_34801,N_34808);
nand U35141 (N_35141,N_34779,N_34810);
and U35142 (N_35142,N_34943,N_34751);
and U35143 (N_35143,N_34885,N_34890);
or U35144 (N_35144,N_34861,N_34847);
xnor U35145 (N_35145,N_34925,N_34957);
nand U35146 (N_35146,N_34792,N_34966);
nor U35147 (N_35147,N_34942,N_34906);
xnor U35148 (N_35148,N_34916,N_34859);
or U35149 (N_35149,N_34793,N_34764);
and U35150 (N_35150,N_34949,N_34833);
nor U35151 (N_35151,N_34905,N_34814);
and U35152 (N_35152,N_34829,N_34827);
nand U35153 (N_35153,N_34762,N_34984);
and U35154 (N_35154,N_34849,N_34937);
nor U35155 (N_35155,N_34875,N_34983);
and U35156 (N_35156,N_34987,N_34770);
nor U35157 (N_35157,N_34824,N_34982);
nand U35158 (N_35158,N_34793,N_34783);
and U35159 (N_35159,N_34892,N_34750);
and U35160 (N_35160,N_34757,N_34828);
xor U35161 (N_35161,N_34753,N_34842);
or U35162 (N_35162,N_34855,N_34861);
nand U35163 (N_35163,N_34844,N_34751);
xnor U35164 (N_35164,N_34908,N_34985);
nor U35165 (N_35165,N_34922,N_34823);
nand U35166 (N_35166,N_34841,N_34918);
xor U35167 (N_35167,N_34872,N_34938);
and U35168 (N_35168,N_34865,N_34782);
xor U35169 (N_35169,N_34764,N_34905);
xnor U35170 (N_35170,N_34777,N_34932);
or U35171 (N_35171,N_34853,N_34925);
or U35172 (N_35172,N_34977,N_34928);
and U35173 (N_35173,N_34847,N_34999);
xor U35174 (N_35174,N_34960,N_34950);
and U35175 (N_35175,N_34979,N_34933);
nand U35176 (N_35176,N_34948,N_34867);
nand U35177 (N_35177,N_34878,N_34917);
nand U35178 (N_35178,N_34876,N_34773);
and U35179 (N_35179,N_34979,N_34951);
and U35180 (N_35180,N_34808,N_34798);
and U35181 (N_35181,N_34771,N_34941);
nor U35182 (N_35182,N_34881,N_34849);
or U35183 (N_35183,N_34913,N_34812);
nand U35184 (N_35184,N_34849,N_34864);
xnor U35185 (N_35185,N_34909,N_34954);
and U35186 (N_35186,N_34833,N_34876);
and U35187 (N_35187,N_34889,N_34816);
nor U35188 (N_35188,N_34914,N_34751);
nand U35189 (N_35189,N_34770,N_34996);
and U35190 (N_35190,N_34934,N_34782);
nor U35191 (N_35191,N_34951,N_34944);
nand U35192 (N_35192,N_34959,N_34914);
xnor U35193 (N_35193,N_34957,N_34899);
and U35194 (N_35194,N_34841,N_34876);
or U35195 (N_35195,N_34813,N_34995);
and U35196 (N_35196,N_34766,N_34822);
nand U35197 (N_35197,N_34936,N_34756);
xnor U35198 (N_35198,N_34980,N_34978);
nor U35199 (N_35199,N_34882,N_34994);
nor U35200 (N_35200,N_34831,N_34755);
nor U35201 (N_35201,N_34912,N_34873);
xnor U35202 (N_35202,N_34862,N_34770);
nor U35203 (N_35203,N_34910,N_34890);
nand U35204 (N_35204,N_34823,N_34820);
xor U35205 (N_35205,N_34857,N_34891);
nand U35206 (N_35206,N_34799,N_34934);
xnor U35207 (N_35207,N_34924,N_34760);
and U35208 (N_35208,N_34852,N_34918);
xnor U35209 (N_35209,N_34983,N_34908);
or U35210 (N_35210,N_34983,N_34922);
nor U35211 (N_35211,N_34824,N_34873);
nand U35212 (N_35212,N_34894,N_34934);
xnor U35213 (N_35213,N_34884,N_34968);
or U35214 (N_35214,N_34803,N_34941);
and U35215 (N_35215,N_34840,N_34949);
xnor U35216 (N_35216,N_34850,N_34968);
xor U35217 (N_35217,N_34887,N_34770);
nand U35218 (N_35218,N_34782,N_34916);
nor U35219 (N_35219,N_34860,N_34935);
or U35220 (N_35220,N_34932,N_34826);
or U35221 (N_35221,N_34831,N_34851);
xnor U35222 (N_35222,N_34947,N_34833);
nor U35223 (N_35223,N_34862,N_34865);
or U35224 (N_35224,N_34818,N_34796);
nor U35225 (N_35225,N_34828,N_34763);
or U35226 (N_35226,N_34922,N_34818);
nor U35227 (N_35227,N_34919,N_34854);
nand U35228 (N_35228,N_34885,N_34985);
and U35229 (N_35229,N_34902,N_34922);
and U35230 (N_35230,N_34768,N_34985);
or U35231 (N_35231,N_34939,N_34773);
nand U35232 (N_35232,N_34966,N_34992);
or U35233 (N_35233,N_34811,N_34855);
nor U35234 (N_35234,N_34990,N_34928);
nand U35235 (N_35235,N_34809,N_34950);
xor U35236 (N_35236,N_34963,N_34800);
and U35237 (N_35237,N_34835,N_34905);
xnor U35238 (N_35238,N_34842,N_34989);
xnor U35239 (N_35239,N_34767,N_34802);
nand U35240 (N_35240,N_34788,N_34910);
nand U35241 (N_35241,N_34969,N_34947);
or U35242 (N_35242,N_34761,N_34826);
or U35243 (N_35243,N_34978,N_34937);
and U35244 (N_35244,N_34780,N_34845);
nor U35245 (N_35245,N_34767,N_34893);
nand U35246 (N_35246,N_34939,N_34917);
xnor U35247 (N_35247,N_34891,N_34802);
and U35248 (N_35248,N_34844,N_34861);
nand U35249 (N_35249,N_34977,N_34902);
xor U35250 (N_35250,N_35239,N_35247);
or U35251 (N_35251,N_35154,N_35014);
xor U35252 (N_35252,N_35196,N_35182);
or U35253 (N_35253,N_35229,N_35051);
or U35254 (N_35254,N_35195,N_35115);
xnor U35255 (N_35255,N_35123,N_35158);
or U35256 (N_35256,N_35000,N_35220);
nor U35257 (N_35257,N_35032,N_35075);
and U35258 (N_35258,N_35160,N_35070);
or U35259 (N_35259,N_35230,N_35164);
nand U35260 (N_35260,N_35235,N_35117);
nand U35261 (N_35261,N_35095,N_35097);
xor U35262 (N_35262,N_35168,N_35128);
xnor U35263 (N_35263,N_35024,N_35145);
and U35264 (N_35264,N_35137,N_35105);
nand U35265 (N_35265,N_35039,N_35236);
nor U35266 (N_35266,N_35143,N_35172);
or U35267 (N_35267,N_35203,N_35042);
and U35268 (N_35268,N_35101,N_35170);
xnor U35269 (N_35269,N_35006,N_35028);
xnor U35270 (N_35270,N_35085,N_35036);
xor U35271 (N_35271,N_35017,N_35161);
and U35272 (N_35272,N_35033,N_35233);
or U35273 (N_35273,N_35073,N_35237);
and U35274 (N_35274,N_35001,N_35022);
xnor U35275 (N_35275,N_35029,N_35193);
nor U35276 (N_35276,N_35133,N_35003);
xnor U35277 (N_35277,N_35238,N_35165);
or U35278 (N_35278,N_35059,N_35119);
or U35279 (N_35279,N_35194,N_35149);
nand U35280 (N_35280,N_35118,N_35088);
nand U35281 (N_35281,N_35197,N_35210);
nand U35282 (N_35282,N_35030,N_35010);
and U35283 (N_35283,N_35108,N_35183);
and U35284 (N_35284,N_35249,N_35111);
nand U35285 (N_35285,N_35018,N_35023);
or U35286 (N_35286,N_35005,N_35192);
and U35287 (N_35287,N_35110,N_35140);
and U35288 (N_35288,N_35175,N_35081);
xor U35289 (N_35289,N_35144,N_35217);
xnor U35290 (N_35290,N_35087,N_35082);
and U35291 (N_35291,N_35157,N_35050);
or U35292 (N_35292,N_35178,N_35244);
and U35293 (N_35293,N_35212,N_35112);
or U35294 (N_35294,N_35216,N_35248);
xnor U35295 (N_35295,N_35027,N_35054);
nor U35296 (N_35296,N_35132,N_35093);
or U35297 (N_35297,N_35113,N_35222);
nand U35298 (N_35298,N_35114,N_35211);
nand U35299 (N_35299,N_35246,N_35231);
and U35300 (N_35300,N_35184,N_35130);
nor U35301 (N_35301,N_35067,N_35065);
or U35302 (N_35302,N_35173,N_35189);
and U35303 (N_35303,N_35138,N_35198);
nand U35304 (N_35304,N_35103,N_35146);
nor U35305 (N_35305,N_35046,N_35076);
nand U35306 (N_35306,N_35031,N_35156);
and U35307 (N_35307,N_35100,N_35056);
nor U35308 (N_35308,N_35241,N_35190);
and U35309 (N_35309,N_35135,N_35092);
xnor U35310 (N_35310,N_35007,N_35038);
or U35311 (N_35311,N_35109,N_35226);
xor U35312 (N_35312,N_35185,N_35011);
nand U35313 (N_35313,N_35209,N_35136);
and U35314 (N_35314,N_35129,N_35052);
nand U35315 (N_35315,N_35060,N_35094);
and U35316 (N_35316,N_35064,N_35057);
xnor U35317 (N_35317,N_35163,N_35245);
nand U35318 (N_35318,N_35047,N_35131);
nand U35319 (N_35319,N_35171,N_35008);
nand U35320 (N_35320,N_35240,N_35019);
nor U35321 (N_35321,N_35035,N_35228);
nor U35322 (N_35322,N_35116,N_35043);
nand U35323 (N_35323,N_35134,N_35208);
xnor U35324 (N_35324,N_35013,N_35021);
or U35325 (N_35325,N_35166,N_35126);
xor U35326 (N_35326,N_35063,N_35139);
nor U35327 (N_35327,N_35049,N_35153);
and U35328 (N_35328,N_35053,N_35004);
nor U35329 (N_35329,N_35147,N_35242);
xnor U35330 (N_35330,N_35181,N_35096);
nor U35331 (N_35331,N_35077,N_35176);
or U35332 (N_35332,N_35159,N_35012);
nor U35333 (N_35333,N_35102,N_35083);
and U35334 (N_35334,N_35232,N_35151);
nand U35335 (N_35335,N_35214,N_35098);
or U35336 (N_35336,N_35150,N_35125);
nand U35337 (N_35337,N_35058,N_35169);
or U35338 (N_35338,N_35104,N_35223);
nand U35339 (N_35339,N_35219,N_35078);
xnor U35340 (N_35340,N_35068,N_35048);
xor U35341 (N_35341,N_35200,N_35188);
or U35342 (N_35342,N_35084,N_35199);
and U35343 (N_35343,N_35080,N_35148);
or U35344 (N_35344,N_35155,N_35234);
xor U35345 (N_35345,N_35162,N_35243);
and U35346 (N_35346,N_35089,N_35121);
or U35347 (N_35347,N_35090,N_35215);
nand U35348 (N_35348,N_35191,N_35086);
xnor U35349 (N_35349,N_35205,N_35227);
and U35350 (N_35350,N_35072,N_35179);
xnor U35351 (N_35351,N_35106,N_35091);
nor U35352 (N_35352,N_35218,N_35122);
and U35353 (N_35353,N_35061,N_35120);
xnor U35354 (N_35354,N_35002,N_35177);
xnor U35355 (N_35355,N_35201,N_35041);
xnor U35356 (N_35356,N_35204,N_35016);
nor U35357 (N_35357,N_35045,N_35079);
and U35358 (N_35358,N_35055,N_35074);
or U35359 (N_35359,N_35167,N_35009);
xor U35360 (N_35360,N_35213,N_35025);
nor U35361 (N_35361,N_35099,N_35066);
or U35362 (N_35362,N_35186,N_35026);
and U35363 (N_35363,N_35221,N_35127);
xnor U35364 (N_35364,N_35040,N_35207);
nand U35365 (N_35365,N_35062,N_35071);
or U35366 (N_35366,N_35044,N_35037);
xnor U35367 (N_35367,N_35224,N_35225);
nand U35368 (N_35368,N_35020,N_35141);
xor U35369 (N_35369,N_35174,N_35152);
xor U35370 (N_35370,N_35180,N_35034);
nor U35371 (N_35371,N_35142,N_35202);
xor U35372 (N_35372,N_35015,N_35069);
and U35373 (N_35373,N_35187,N_35107);
and U35374 (N_35374,N_35124,N_35206);
xor U35375 (N_35375,N_35177,N_35133);
and U35376 (N_35376,N_35147,N_35087);
and U35377 (N_35377,N_35070,N_35006);
nand U35378 (N_35378,N_35231,N_35166);
and U35379 (N_35379,N_35139,N_35037);
nor U35380 (N_35380,N_35247,N_35000);
nand U35381 (N_35381,N_35060,N_35180);
or U35382 (N_35382,N_35082,N_35106);
or U35383 (N_35383,N_35068,N_35118);
or U35384 (N_35384,N_35136,N_35153);
xnor U35385 (N_35385,N_35102,N_35234);
nor U35386 (N_35386,N_35067,N_35127);
and U35387 (N_35387,N_35052,N_35211);
and U35388 (N_35388,N_35177,N_35171);
and U35389 (N_35389,N_35015,N_35112);
or U35390 (N_35390,N_35107,N_35091);
xor U35391 (N_35391,N_35009,N_35069);
nor U35392 (N_35392,N_35123,N_35172);
or U35393 (N_35393,N_35138,N_35209);
nor U35394 (N_35394,N_35031,N_35008);
or U35395 (N_35395,N_35137,N_35083);
and U35396 (N_35396,N_35229,N_35122);
or U35397 (N_35397,N_35041,N_35143);
nand U35398 (N_35398,N_35195,N_35178);
or U35399 (N_35399,N_35184,N_35188);
nand U35400 (N_35400,N_35196,N_35016);
and U35401 (N_35401,N_35125,N_35094);
xor U35402 (N_35402,N_35162,N_35102);
nor U35403 (N_35403,N_35174,N_35020);
and U35404 (N_35404,N_35073,N_35065);
or U35405 (N_35405,N_35044,N_35147);
nor U35406 (N_35406,N_35072,N_35051);
nand U35407 (N_35407,N_35005,N_35056);
or U35408 (N_35408,N_35106,N_35151);
or U35409 (N_35409,N_35201,N_35011);
or U35410 (N_35410,N_35155,N_35056);
xnor U35411 (N_35411,N_35156,N_35120);
nand U35412 (N_35412,N_35110,N_35037);
nand U35413 (N_35413,N_35208,N_35063);
nor U35414 (N_35414,N_35208,N_35062);
nand U35415 (N_35415,N_35187,N_35224);
xor U35416 (N_35416,N_35099,N_35174);
nor U35417 (N_35417,N_35247,N_35180);
nor U35418 (N_35418,N_35112,N_35104);
xor U35419 (N_35419,N_35178,N_35130);
or U35420 (N_35420,N_35170,N_35119);
and U35421 (N_35421,N_35249,N_35044);
xor U35422 (N_35422,N_35003,N_35113);
xnor U35423 (N_35423,N_35224,N_35007);
or U35424 (N_35424,N_35161,N_35133);
xnor U35425 (N_35425,N_35015,N_35155);
nor U35426 (N_35426,N_35139,N_35105);
nor U35427 (N_35427,N_35140,N_35242);
and U35428 (N_35428,N_35028,N_35238);
or U35429 (N_35429,N_35068,N_35100);
nor U35430 (N_35430,N_35125,N_35015);
and U35431 (N_35431,N_35164,N_35042);
nor U35432 (N_35432,N_35203,N_35087);
xnor U35433 (N_35433,N_35004,N_35019);
and U35434 (N_35434,N_35112,N_35239);
or U35435 (N_35435,N_35207,N_35076);
nand U35436 (N_35436,N_35074,N_35048);
and U35437 (N_35437,N_35103,N_35134);
nor U35438 (N_35438,N_35034,N_35051);
nor U35439 (N_35439,N_35069,N_35093);
xnor U35440 (N_35440,N_35109,N_35212);
and U35441 (N_35441,N_35221,N_35145);
nand U35442 (N_35442,N_35165,N_35150);
or U35443 (N_35443,N_35024,N_35128);
or U35444 (N_35444,N_35191,N_35164);
nor U35445 (N_35445,N_35186,N_35241);
nor U35446 (N_35446,N_35120,N_35149);
nor U35447 (N_35447,N_35244,N_35069);
or U35448 (N_35448,N_35163,N_35226);
nand U35449 (N_35449,N_35125,N_35237);
and U35450 (N_35450,N_35176,N_35136);
nor U35451 (N_35451,N_35016,N_35102);
nor U35452 (N_35452,N_35154,N_35161);
xor U35453 (N_35453,N_35097,N_35099);
or U35454 (N_35454,N_35133,N_35106);
xor U35455 (N_35455,N_35086,N_35025);
nor U35456 (N_35456,N_35167,N_35059);
and U35457 (N_35457,N_35228,N_35082);
xnor U35458 (N_35458,N_35231,N_35079);
or U35459 (N_35459,N_35023,N_35084);
nor U35460 (N_35460,N_35074,N_35172);
or U35461 (N_35461,N_35230,N_35177);
xor U35462 (N_35462,N_35124,N_35023);
or U35463 (N_35463,N_35008,N_35065);
xor U35464 (N_35464,N_35112,N_35226);
nand U35465 (N_35465,N_35103,N_35242);
or U35466 (N_35466,N_35214,N_35068);
and U35467 (N_35467,N_35025,N_35160);
or U35468 (N_35468,N_35187,N_35180);
xnor U35469 (N_35469,N_35226,N_35074);
or U35470 (N_35470,N_35102,N_35048);
nor U35471 (N_35471,N_35037,N_35122);
nand U35472 (N_35472,N_35099,N_35052);
and U35473 (N_35473,N_35052,N_35245);
or U35474 (N_35474,N_35235,N_35000);
and U35475 (N_35475,N_35242,N_35122);
nor U35476 (N_35476,N_35088,N_35203);
or U35477 (N_35477,N_35070,N_35080);
xor U35478 (N_35478,N_35134,N_35146);
or U35479 (N_35479,N_35098,N_35210);
nand U35480 (N_35480,N_35149,N_35060);
and U35481 (N_35481,N_35071,N_35035);
nand U35482 (N_35482,N_35093,N_35249);
nand U35483 (N_35483,N_35227,N_35132);
xnor U35484 (N_35484,N_35101,N_35175);
xor U35485 (N_35485,N_35132,N_35236);
xnor U35486 (N_35486,N_35010,N_35072);
nor U35487 (N_35487,N_35115,N_35142);
xnor U35488 (N_35488,N_35094,N_35150);
or U35489 (N_35489,N_35079,N_35226);
xnor U35490 (N_35490,N_35037,N_35003);
xor U35491 (N_35491,N_35173,N_35238);
and U35492 (N_35492,N_35249,N_35092);
and U35493 (N_35493,N_35238,N_35139);
nor U35494 (N_35494,N_35043,N_35235);
nand U35495 (N_35495,N_35090,N_35196);
nor U35496 (N_35496,N_35081,N_35117);
xnor U35497 (N_35497,N_35175,N_35217);
nor U35498 (N_35498,N_35048,N_35135);
nor U35499 (N_35499,N_35133,N_35004);
and U35500 (N_35500,N_35353,N_35273);
and U35501 (N_35501,N_35440,N_35411);
nand U35502 (N_35502,N_35336,N_35345);
nor U35503 (N_35503,N_35361,N_35334);
nor U35504 (N_35504,N_35298,N_35370);
and U35505 (N_35505,N_35275,N_35299);
nor U35506 (N_35506,N_35465,N_35392);
or U35507 (N_35507,N_35255,N_35481);
nor U35508 (N_35508,N_35486,N_35401);
nand U35509 (N_35509,N_35406,N_35423);
or U35510 (N_35510,N_35258,N_35412);
xnor U35511 (N_35511,N_35252,N_35407);
and U35512 (N_35512,N_35438,N_35292);
or U35513 (N_35513,N_35377,N_35359);
and U35514 (N_35514,N_35363,N_35385);
nor U35515 (N_35515,N_35270,N_35371);
nor U35516 (N_35516,N_35400,N_35290);
nand U35517 (N_35517,N_35383,N_35282);
or U35518 (N_35518,N_35435,N_35442);
xor U35519 (N_35519,N_35351,N_35264);
nand U35520 (N_35520,N_35356,N_35259);
xor U35521 (N_35521,N_35338,N_35414);
xnor U35522 (N_35522,N_35410,N_35395);
nand U35523 (N_35523,N_35462,N_35434);
xor U35524 (N_35524,N_35297,N_35253);
nor U35525 (N_35525,N_35478,N_35350);
nor U35526 (N_35526,N_35380,N_35289);
nor U35527 (N_35527,N_35376,N_35330);
and U35528 (N_35528,N_35307,N_35452);
nor U35529 (N_35529,N_35287,N_35387);
nand U35530 (N_35530,N_35327,N_35293);
nand U35531 (N_35531,N_35313,N_35367);
and U35532 (N_35532,N_35357,N_35429);
or U35533 (N_35533,N_35384,N_35453);
nand U35534 (N_35534,N_35403,N_35381);
and U35535 (N_35535,N_35346,N_35267);
nor U35536 (N_35536,N_35262,N_35343);
xor U35537 (N_35537,N_35458,N_35467);
or U35538 (N_35538,N_35416,N_35421);
xnor U35539 (N_35539,N_35487,N_35301);
nor U35540 (N_35540,N_35328,N_35344);
xor U35541 (N_35541,N_35348,N_35433);
xnor U35542 (N_35542,N_35399,N_35316);
xor U35543 (N_35543,N_35254,N_35446);
nor U35544 (N_35544,N_35490,N_35482);
or U35545 (N_35545,N_35324,N_35422);
nand U35546 (N_35546,N_35447,N_35499);
nand U35547 (N_35547,N_35358,N_35477);
and U35548 (N_35548,N_35280,N_35460);
nand U35549 (N_35549,N_35302,N_35450);
nand U35550 (N_35550,N_35455,N_35360);
and U35551 (N_35551,N_35374,N_35314);
and U35552 (N_35552,N_35451,N_35300);
xor U35553 (N_35553,N_35295,N_35492);
nand U35554 (N_35554,N_35496,N_35261);
xor U35555 (N_35555,N_35271,N_35272);
or U35556 (N_35556,N_35266,N_35340);
xnor U35557 (N_35557,N_35257,N_35472);
or U35558 (N_35558,N_35473,N_35480);
nand U35559 (N_35559,N_35366,N_35365);
or U35560 (N_35560,N_35484,N_35488);
nor U35561 (N_35561,N_35250,N_35296);
or U35562 (N_35562,N_35339,N_35483);
or U35563 (N_35563,N_35388,N_35493);
nand U35564 (N_35564,N_35305,N_35286);
xnor U35565 (N_35565,N_35448,N_35386);
xnor U35566 (N_35566,N_35362,N_35394);
xnor U35567 (N_35567,N_35441,N_35278);
nand U35568 (N_35568,N_35449,N_35456);
nor U35569 (N_35569,N_35437,N_35439);
nand U35570 (N_35570,N_35319,N_35475);
and U35571 (N_35571,N_35428,N_35479);
xor U35572 (N_35572,N_35379,N_35393);
nand U35573 (N_35573,N_35333,N_35276);
xnor U35574 (N_35574,N_35418,N_35329);
or U35575 (N_35575,N_35463,N_35445);
xor U35576 (N_35576,N_35268,N_35265);
nand U35577 (N_35577,N_35405,N_35409);
xnor U35578 (N_35578,N_35263,N_35331);
nor U35579 (N_35579,N_35341,N_35323);
or U35580 (N_35580,N_35373,N_35495);
and U35581 (N_35581,N_35485,N_35432);
nor U35582 (N_35582,N_35498,N_35491);
and U35583 (N_35583,N_35260,N_35279);
nand U35584 (N_35584,N_35332,N_35378);
xor U35585 (N_35585,N_35466,N_35284);
xnor U35586 (N_35586,N_35459,N_35326);
and U35587 (N_35587,N_35454,N_35337);
and U35588 (N_35588,N_35396,N_35431);
nor U35589 (N_35589,N_35303,N_35390);
xor U35590 (N_35590,N_35369,N_35281);
or U35591 (N_35591,N_35494,N_35309);
and U35592 (N_35592,N_35355,N_35352);
nor U35593 (N_35593,N_35294,N_35408);
nand U35594 (N_35594,N_35285,N_35425);
or U35595 (N_35595,N_35468,N_35469);
and U35596 (N_35596,N_35404,N_35322);
and U35597 (N_35597,N_35424,N_35426);
nand U35598 (N_35598,N_35402,N_35443);
nand U35599 (N_35599,N_35372,N_35335);
nand U35600 (N_35600,N_35375,N_35283);
and U35601 (N_35601,N_35389,N_35342);
or U35602 (N_35602,N_35415,N_35420);
nor U35603 (N_35603,N_35457,N_35274);
and U35604 (N_35604,N_35288,N_35306);
nand U35605 (N_35605,N_35347,N_35497);
nand U35606 (N_35606,N_35269,N_35320);
xnor U35607 (N_35607,N_35427,N_35308);
nor U35608 (N_35608,N_35304,N_35251);
nand U35609 (N_35609,N_35419,N_35382);
xor U35610 (N_35610,N_35398,N_35413);
or U35611 (N_35611,N_35397,N_35318);
nor U35612 (N_35612,N_35430,N_35464);
xor U35613 (N_35613,N_35354,N_35317);
xor U35614 (N_35614,N_35315,N_35277);
or U35615 (N_35615,N_35291,N_35310);
or U35616 (N_35616,N_35256,N_35461);
nand U35617 (N_35617,N_35368,N_35364);
and U35618 (N_35618,N_35311,N_35312);
and U35619 (N_35619,N_35474,N_35349);
and U35620 (N_35620,N_35471,N_35417);
or U35621 (N_35621,N_35444,N_35321);
nand U35622 (N_35622,N_35470,N_35476);
and U35623 (N_35623,N_35489,N_35436);
xnor U35624 (N_35624,N_35391,N_35325);
nand U35625 (N_35625,N_35355,N_35488);
nand U35626 (N_35626,N_35260,N_35349);
xor U35627 (N_35627,N_35498,N_35397);
nor U35628 (N_35628,N_35440,N_35369);
or U35629 (N_35629,N_35446,N_35452);
nand U35630 (N_35630,N_35433,N_35488);
nand U35631 (N_35631,N_35273,N_35458);
nand U35632 (N_35632,N_35368,N_35388);
xnor U35633 (N_35633,N_35379,N_35387);
nand U35634 (N_35634,N_35431,N_35294);
nor U35635 (N_35635,N_35348,N_35280);
nand U35636 (N_35636,N_35368,N_35379);
nand U35637 (N_35637,N_35346,N_35375);
xnor U35638 (N_35638,N_35271,N_35263);
nand U35639 (N_35639,N_35446,N_35431);
xor U35640 (N_35640,N_35294,N_35385);
or U35641 (N_35641,N_35401,N_35392);
and U35642 (N_35642,N_35431,N_35384);
nor U35643 (N_35643,N_35353,N_35476);
or U35644 (N_35644,N_35356,N_35405);
xnor U35645 (N_35645,N_35322,N_35355);
or U35646 (N_35646,N_35405,N_35392);
nor U35647 (N_35647,N_35446,N_35372);
xnor U35648 (N_35648,N_35257,N_35481);
nor U35649 (N_35649,N_35417,N_35367);
nor U35650 (N_35650,N_35263,N_35276);
nand U35651 (N_35651,N_35332,N_35334);
xnor U35652 (N_35652,N_35292,N_35356);
nor U35653 (N_35653,N_35338,N_35430);
nand U35654 (N_35654,N_35467,N_35328);
or U35655 (N_35655,N_35346,N_35270);
nor U35656 (N_35656,N_35374,N_35475);
and U35657 (N_35657,N_35328,N_35427);
or U35658 (N_35658,N_35481,N_35279);
nand U35659 (N_35659,N_35345,N_35398);
and U35660 (N_35660,N_35344,N_35405);
and U35661 (N_35661,N_35442,N_35476);
nor U35662 (N_35662,N_35488,N_35350);
nand U35663 (N_35663,N_35292,N_35315);
and U35664 (N_35664,N_35260,N_35417);
or U35665 (N_35665,N_35332,N_35286);
nand U35666 (N_35666,N_35344,N_35490);
or U35667 (N_35667,N_35497,N_35450);
xor U35668 (N_35668,N_35437,N_35486);
and U35669 (N_35669,N_35297,N_35316);
nand U35670 (N_35670,N_35332,N_35424);
nand U35671 (N_35671,N_35286,N_35344);
nor U35672 (N_35672,N_35348,N_35271);
or U35673 (N_35673,N_35312,N_35371);
nor U35674 (N_35674,N_35252,N_35441);
nand U35675 (N_35675,N_35373,N_35428);
nand U35676 (N_35676,N_35424,N_35397);
nand U35677 (N_35677,N_35405,N_35305);
or U35678 (N_35678,N_35460,N_35433);
and U35679 (N_35679,N_35298,N_35272);
nor U35680 (N_35680,N_35343,N_35393);
nand U35681 (N_35681,N_35263,N_35264);
and U35682 (N_35682,N_35382,N_35365);
xor U35683 (N_35683,N_35305,N_35298);
and U35684 (N_35684,N_35324,N_35480);
and U35685 (N_35685,N_35395,N_35411);
or U35686 (N_35686,N_35438,N_35388);
or U35687 (N_35687,N_35290,N_35335);
xor U35688 (N_35688,N_35371,N_35311);
or U35689 (N_35689,N_35398,N_35310);
nor U35690 (N_35690,N_35385,N_35404);
nand U35691 (N_35691,N_35467,N_35271);
nand U35692 (N_35692,N_35375,N_35318);
xnor U35693 (N_35693,N_35426,N_35286);
nand U35694 (N_35694,N_35471,N_35384);
or U35695 (N_35695,N_35477,N_35320);
nor U35696 (N_35696,N_35451,N_35321);
nand U35697 (N_35697,N_35344,N_35327);
or U35698 (N_35698,N_35468,N_35399);
nor U35699 (N_35699,N_35366,N_35444);
or U35700 (N_35700,N_35499,N_35277);
xnor U35701 (N_35701,N_35317,N_35298);
or U35702 (N_35702,N_35319,N_35290);
nand U35703 (N_35703,N_35367,N_35380);
nor U35704 (N_35704,N_35282,N_35303);
or U35705 (N_35705,N_35328,N_35317);
and U35706 (N_35706,N_35355,N_35481);
xnor U35707 (N_35707,N_35259,N_35275);
nand U35708 (N_35708,N_35430,N_35397);
and U35709 (N_35709,N_35485,N_35253);
xnor U35710 (N_35710,N_35349,N_35398);
nand U35711 (N_35711,N_35431,N_35357);
xnor U35712 (N_35712,N_35334,N_35313);
nand U35713 (N_35713,N_35446,N_35259);
nor U35714 (N_35714,N_35307,N_35270);
and U35715 (N_35715,N_35330,N_35314);
nor U35716 (N_35716,N_35486,N_35360);
nand U35717 (N_35717,N_35353,N_35468);
nand U35718 (N_35718,N_35462,N_35386);
nor U35719 (N_35719,N_35406,N_35421);
or U35720 (N_35720,N_35328,N_35460);
or U35721 (N_35721,N_35416,N_35314);
or U35722 (N_35722,N_35490,N_35353);
or U35723 (N_35723,N_35486,N_35310);
xnor U35724 (N_35724,N_35335,N_35461);
nand U35725 (N_35725,N_35484,N_35343);
and U35726 (N_35726,N_35484,N_35287);
nand U35727 (N_35727,N_35282,N_35430);
or U35728 (N_35728,N_35338,N_35366);
nand U35729 (N_35729,N_35270,N_35400);
xnor U35730 (N_35730,N_35486,N_35473);
nand U35731 (N_35731,N_35327,N_35352);
xnor U35732 (N_35732,N_35371,N_35343);
nand U35733 (N_35733,N_35389,N_35479);
xnor U35734 (N_35734,N_35349,N_35492);
nand U35735 (N_35735,N_35277,N_35371);
xor U35736 (N_35736,N_35361,N_35480);
and U35737 (N_35737,N_35356,N_35390);
or U35738 (N_35738,N_35359,N_35314);
nand U35739 (N_35739,N_35279,N_35311);
and U35740 (N_35740,N_35272,N_35461);
nand U35741 (N_35741,N_35395,N_35351);
nand U35742 (N_35742,N_35363,N_35481);
nor U35743 (N_35743,N_35413,N_35314);
and U35744 (N_35744,N_35250,N_35428);
nor U35745 (N_35745,N_35483,N_35488);
or U35746 (N_35746,N_35444,N_35425);
or U35747 (N_35747,N_35412,N_35416);
nand U35748 (N_35748,N_35403,N_35356);
nor U35749 (N_35749,N_35361,N_35463);
nand U35750 (N_35750,N_35719,N_35554);
or U35751 (N_35751,N_35679,N_35715);
nand U35752 (N_35752,N_35546,N_35542);
or U35753 (N_35753,N_35512,N_35670);
or U35754 (N_35754,N_35585,N_35571);
xor U35755 (N_35755,N_35532,N_35710);
nand U35756 (N_35756,N_35541,N_35613);
or U35757 (N_35757,N_35620,N_35608);
nor U35758 (N_35758,N_35616,N_35568);
xor U35759 (N_35759,N_35527,N_35652);
nand U35760 (N_35760,N_35696,N_35517);
and U35761 (N_35761,N_35632,N_35572);
or U35762 (N_35762,N_35737,N_35666);
nor U35763 (N_35763,N_35721,N_35627);
or U35764 (N_35764,N_35558,N_35686);
nand U35765 (N_35765,N_35544,N_35559);
nand U35766 (N_35766,N_35680,N_35665);
or U35767 (N_35767,N_35619,N_35743);
and U35768 (N_35768,N_35535,N_35557);
or U35769 (N_35769,N_35553,N_35582);
nor U35770 (N_35770,N_35712,N_35525);
xor U35771 (N_35771,N_35511,N_35706);
or U35772 (N_35772,N_35579,N_35731);
nor U35773 (N_35773,N_35503,N_35614);
nor U35774 (N_35774,N_35515,N_35725);
nand U35775 (N_35775,N_35707,N_35703);
nor U35776 (N_35776,N_35672,N_35508);
and U35777 (N_35777,N_35700,N_35705);
nand U35778 (N_35778,N_35726,N_35714);
or U35779 (N_35779,N_35640,N_35528);
or U35780 (N_35780,N_35661,N_35513);
nor U35781 (N_35781,N_35501,N_35556);
nand U35782 (N_35782,N_35656,N_35734);
nor U35783 (N_35783,N_35746,N_35685);
nor U35784 (N_35784,N_35654,N_35575);
and U35785 (N_35785,N_35645,N_35567);
nor U35786 (N_35786,N_35713,N_35641);
nand U35787 (N_35787,N_35624,N_35583);
nand U35788 (N_35788,N_35650,N_35735);
and U35789 (N_35789,N_35601,N_35736);
or U35790 (N_35790,N_35637,N_35563);
and U35791 (N_35791,N_35742,N_35574);
nand U35792 (N_35792,N_35524,N_35610);
nand U35793 (N_35793,N_35519,N_35674);
nor U35794 (N_35794,N_35642,N_35505);
or U35795 (N_35795,N_35662,N_35718);
xor U35796 (N_35796,N_35593,N_35590);
nand U35797 (N_35797,N_35653,N_35693);
and U35798 (N_35798,N_35521,N_35600);
nand U35799 (N_35799,N_35671,N_35548);
nor U35800 (N_35800,N_35588,N_35540);
or U35801 (N_35801,N_35595,N_35529);
and U35802 (N_35802,N_35561,N_35691);
xor U35803 (N_35803,N_35668,N_35500);
and U35804 (N_35804,N_35722,N_35678);
xor U35805 (N_35805,N_35748,N_35516);
and U35806 (N_35806,N_35741,N_35584);
nor U35807 (N_35807,N_35651,N_35720);
xor U35808 (N_35808,N_35599,N_35667);
or U35809 (N_35809,N_35676,N_35536);
xor U35810 (N_35810,N_35522,N_35682);
nand U35811 (N_35811,N_35638,N_35580);
nor U35812 (N_35812,N_35581,N_35659);
xor U35813 (N_35813,N_35576,N_35539);
xnor U35814 (N_35814,N_35586,N_35695);
or U35815 (N_35815,N_35514,N_35739);
or U35816 (N_35816,N_35749,N_35628);
nand U35817 (N_35817,N_35533,N_35502);
or U35818 (N_35818,N_35745,N_35692);
xor U35819 (N_35819,N_35607,N_35708);
nor U35820 (N_35820,N_35688,N_35740);
and U35821 (N_35821,N_35675,N_35534);
or U35822 (N_35822,N_35663,N_35604);
nor U35823 (N_35823,N_35611,N_35550);
nor U35824 (N_35824,N_35606,N_35698);
and U35825 (N_35825,N_35643,N_35615);
xnor U35826 (N_35826,N_35697,N_35597);
nor U35827 (N_35827,N_35612,N_35509);
nor U35828 (N_35828,N_35635,N_35587);
or U35829 (N_35829,N_35626,N_35657);
nand U35830 (N_35830,N_35646,N_35658);
or U35831 (N_35831,N_35631,N_35647);
nor U35832 (N_35832,N_35565,N_35636);
nand U35833 (N_35833,N_35738,N_35723);
xnor U35834 (N_35834,N_35603,N_35547);
or U35835 (N_35835,N_35598,N_35727);
and U35836 (N_35836,N_35555,N_35520);
nor U35837 (N_35837,N_35560,N_35562);
or U35838 (N_35838,N_35744,N_35605);
nor U35839 (N_35839,N_35702,N_35621);
nor U35840 (N_35840,N_35523,N_35673);
xor U35841 (N_35841,N_35617,N_35596);
nor U35842 (N_35842,N_35537,N_35629);
xor U35843 (N_35843,N_35681,N_35578);
or U35844 (N_35844,N_35618,N_35526);
or U35845 (N_35845,N_35709,N_35538);
nor U35846 (N_35846,N_35644,N_35570);
nand U35847 (N_35847,N_35699,N_35602);
nor U35848 (N_35848,N_35591,N_35716);
and U35849 (N_35849,N_35552,N_35639);
xnor U35850 (N_35850,N_35649,N_35711);
or U35851 (N_35851,N_35623,N_35594);
xor U35852 (N_35852,N_35577,N_35566);
or U35853 (N_35853,N_35687,N_35733);
and U35854 (N_35854,N_35689,N_35747);
and U35855 (N_35855,N_35728,N_35683);
and U35856 (N_35856,N_35530,N_35622);
and U35857 (N_35857,N_35684,N_35543);
nor U35858 (N_35858,N_35704,N_35655);
nand U35859 (N_35859,N_35732,N_35625);
nor U35860 (N_35860,N_35504,N_35592);
and U35861 (N_35861,N_35630,N_35660);
nand U35862 (N_35862,N_35694,N_35730);
nand U35863 (N_35863,N_35589,N_35549);
nand U35864 (N_35864,N_35545,N_35677);
nand U35865 (N_35865,N_35573,N_35609);
or U35866 (N_35866,N_35648,N_35690);
xor U35867 (N_35867,N_35664,N_35507);
nand U35868 (N_35868,N_35701,N_35724);
or U35869 (N_35869,N_35717,N_35564);
nor U35870 (N_35870,N_35634,N_35569);
and U35871 (N_35871,N_35669,N_35551);
xnor U35872 (N_35872,N_35510,N_35633);
or U35873 (N_35873,N_35531,N_35729);
and U35874 (N_35874,N_35518,N_35506);
xor U35875 (N_35875,N_35569,N_35530);
and U35876 (N_35876,N_35701,N_35714);
nor U35877 (N_35877,N_35581,N_35619);
xnor U35878 (N_35878,N_35631,N_35659);
xor U35879 (N_35879,N_35604,N_35698);
nand U35880 (N_35880,N_35621,N_35672);
xor U35881 (N_35881,N_35619,N_35676);
xor U35882 (N_35882,N_35619,N_35515);
nand U35883 (N_35883,N_35547,N_35709);
and U35884 (N_35884,N_35622,N_35706);
or U35885 (N_35885,N_35593,N_35559);
xor U35886 (N_35886,N_35514,N_35541);
nand U35887 (N_35887,N_35713,N_35656);
nor U35888 (N_35888,N_35506,N_35731);
nor U35889 (N_35889,N_35645,N_35723);
and U35890 (N_35890,N_35504,N_35610);
and U35891 (N_35891,N_35593,N_35654);
or U35892 (N_35892,N_35619,N_35559);
and U35893 (N_35893,N_35531,N_35748);
and U35894 (N_35894,N_35644,N_35638);
nand U35895 (N_35895,N_35742,N_35711);
or U35896 (N_35896,N_35733,N_35664);
xnor U35897 (N_35897,N_35740,N_35554);
or U35898 (N_35898,N_35733,N_35632);
nand U35899 (N_35899,N_35706,N_35680);
nor U35900 (N_35900,N_35605,N_35529);
nor U35901 (N_35901,N_35718,N_35601);
and U35902 (N_35902,N_35686,N_35689);
xor U35903 (N_35903,N_35585,N_35507);
and U35904 (N_35904,N_35511,N_35503);
or U35905 (N_35905,N_35550,N_35620);
xnor U35906 (N_35906,N_35647,N_35517);
or U35907 (N_35907,N_35518,N_35708);
or U35908 (N_35908,N_35565,N_35697);
xnor U35909 (N_35909,N_35642,N_35624);
and U35910 (N_35910,N_35668,N_35556);
xnor U35911 (N_35911,N_35740,N_35615);
and U35912 (N_35912,N_35572,N_35719);
nor U35913 (N_35913,N_35548,N_35667);
and U35914 (N_35914,N_35744,N_35701);
and U35915 (N_35915,N_35608,N_35601);
nor U35916 (N_35916,N_35622,N_35514);
xor U35917 (N_35917,N_35571,N_35664);
nor U35918 (N_35918,N_35559,N_35671);
and U35919 (N_35919,N_35603,N_35618);
or U35920 (N_35920,N_35549,N_35511);
and U35921 (N_35921,N_35601,N_35533);
and U35922 (N_35922,N_35697,N_35715);
and U35923 (N_35923,N_35712,N_35576);
and U35924 (N_35924,N_35701,N_35666);
and U35925 (N_35925,N_35735,N_35606);
nor U35926 (N_35926,N_35726,N_35718);
xor U35927 (N_35927,N_35500,N_35589);
nor U35928 (N_35928,N_35726,N_35658);
xor U35929 (N_35929,N_35509,N_35623);
xnor U35930 (N_35930,N_35720,N_35606);
xor U35931 (N_35931,N_35654,N_35613);
and U35932 (N_35932,N_35662,N_35614);
nor U35933 (N_35933,N_35616,N_35685);
xnor U35934 (N_35934,N_35565,N_35689);
and U35935 (N_35935,N_35515,N_35610);
nor U35936 (N_35936,N_35540,N_35547);
or U35937 (N_35937,N_35632,N_35542);
xnor U35938 (N_35938,N_35618,N_35719);
nand U35939 (N_35939,N_35660,N_35743);
or U35940 (N_35940,N_35741,N_35715);
xnor U35941 (N_35941,N_35594,N_35626);
nand U35942 (N_35942,N_35517,N_35737);
nor U35943 (N_35943,N_35521,N_35559);
nand U35944 (N_35944,N_35626,N_35508);
nand U35945 (N_35945,N_35625,N_35579);
or U35946 (N_35946,N_35656,N_35636);
or U35947 (N_35947,N_35600,N_35557);
or U35948 (N_35948,N_35647,N_35659);
xor U35949 (N_35949,N_35627,N_35659);
or U35950 (N_35950,N_35567,N_35661);
nand U35951 (N_35951,N_35699,N_35576);
xor U35952 (N_35952,N_35556,N_35640);
xor U35953 (N_35953,N_35562,N_35582);
and U35954 (N_35954,N_35728,N_35722);
and U35955 (N_35955,N_35649,N_35655);
nand U35956 (N_35956,N_35658,N_35599);
xnor U35957 (N_35957,N_35507,N_35620);
xor U35958 (N_35958,N_35691,N_35738);
nand U35959 (N_35959,N_35698,N_35600);
nor U35960 (N_35960,N_35701,N_35505);
or U35961 (N_35961,N_35715,N_35720);
nor U35962 (N_35962,N_35660,N_35736);
or U35963 (N_35963,N_35721,N_35622);
xor U35964 (N_35964,N_35583,N_35747);
and U35965 (N_35965,N_35511,N_35591);
nor U35966 (N_35966,N_35504,N_35540);
or U35967 (N_35967,N_35617,N_35592);
nand U35968 (N_35968,N_35547,N_35505);
or U35969 (N_35969,N_35694,N_35601);
or U35970 (N_35970,N_35702,N_35561);
nand U35971 (N_35971,N_35602,N_35594);
and U35972 (N_35972,N_35749,N_35644);
and U35973 (N_35973,N_35550,N_35680);
and U35974 (N_35974,N_35697,N_35589);
or U35975 (N_35975,N_35715,N_35588);
nand U35976 (N_35976,N_35523,N_35518);
nor U35977 (N_35977,N_35740,N_35566);
nand U35978 (N_35978,N_35568,N_35592);
xnor U35979 (N_35979,N_35628,N_35681);
nor U35980 (N_35980,N_35738,N_35684);
and U35981 (N_35981,N_35629,N_35586);
nor U35982 (N_35982,N_35676,N_35543);
nor U35983 (N_35983,N_35703,N_35518);
nor U35984 (N_35984,N_35670,N_35596);
nor U35985 (N_35985,N_35644,N_35672);
nor U35986 (N_35986,N_35629,N_35689);
nor U35987 (N_35987,N_35663,N_35744);
or U35988 (N_35988,N_35502,N_35590);
nor U35989 (N_35989,N_35548,N_35559);
or U35990 (N_35990,N_35679,N_35675);
xnor U35991 (N_35991,N_35691,N_35592);
or U35992 (N_35992,N_35571,N_35565);
or U35993 (N_35993,N_35722,N_35735);
xnor U35994 (N_35994,N_35698,N_35541);
nand U35995 (N_35995,N_35741,N_35731);
nand U35996 (N_35996,N_35683,N_35584);
and U35997 (N_35997,N_35578,N_35674);
and U35998 (N_35998,N_35696,N_35697);
nand U35999 (N_35999,N_35640,N_35736);
xnor U36000 (N_36000,N_35850,N_35792);
and U36001 (N_36001,N_35891,N_35818);
or U36002 (N_36002,N_35914,N_35965);
xor U36003 (N_36003,N_35861,N_35892);
and U36004 (N_36004,N_35781,N_35790);
xnor U36005 (N_36005,N_35811,N_35981);
or U36006 (N_36006,N_35798,N_35779);
nor U36007 (N_36007,N_35785,N_35973);
xnor U36008 (N_36008,N_35899,N_35947);
nor U36009 (N_36009,N_35900,N_35826);
nor U36010 (N_36010,N_35888,N_35925);
nand U36011 (N_36011,N_35800,N_35944);
nand U36012 (N_36012,N_35830,N_35956);
nor U36013 (N_36013,N_35897,N_35889);
and U36014 (N_36014,N_35905,N_35776);
nand U36015 (N_36015,N_35955,N_35774);
nand U36016 (N_36016,N_35822,N_35838);
nor U36017 (N_36017,N_35812,N_35927);
nand U36018 (N_36018,N_35751,N_35863);
nand U36019 (N_36019,N_35866,N_35986);
or U36020 (N_36020,N_35877,N_35991);
nor U36021 (N_36021,N_35964,N_35980);
or U36022 (N_36022,N_35805,N_35951);
xor U36023 (N_36023,N_35881,N_35756);
xor U36024 (N_36024,N_35894,N_35911);
or U36025 (N_36025,N_35856,N_35876);
and U36026 (N_36026,N_35921,N_35929);
nor U36027 (N_36027,N_35848,N_35868);
nor U36028 (N_36028,N_35815,N_35940);
and U36029 (N_36029,N_35988,N_35860);
nor U36030 (N_36030,N_35928,N_35936);
xor U36031 (N_36031,N_35972,N_35755);
xor U36032 (N_36032,N_35954,N_35898);
nor U36033 (N_36033,N_35885,N_35757);
nand U36034 (N_36034,N_35982,N_35858);
and U36035 (N_36035,N_35807,N_35804);
and U36036 (N_36036,N_35990,N_35904);
and U36037 (N_36037,N_35942,N_35813);
xnor U36038 (N_36038,N_35864,N_35821);
and U36039 (N_36039,N_35976,N_35962);
nor U36040 (N_36040,N_35884,N_35840);
xor U36041 (N_36041,N_35966,N_35855);
and U36042 (N_36042,N_35832,N_35946);
nor U36043 (N_36043,N_35970,N_35880);
or U36044 (N_36044,N_35780,N_35799);
nor U36045 (N_36045,N_35913,N_35852);
xnor U36046 (N_36046,N_35949,N_35907);
or U36047 (N_36047,N_35901,N_35761);
nand U36048 (N_36048,N_35920,N_35854);
and U36049 (N_36049,N_35923,N_35987);
nor U36050 (N_36050,N_35797,N_35778);
and U36051 (N_36051,N_35809,N_35789);
xnor U36052 (N_36052,N_35843,N_35869);
xnor U36053 (N_36053,N_35788,N_35853);
nand U36054 (N_36054,N_35930,N_35859);
xor U36055 (N_36055,N_35924,N_35872);
or U36056 (N_36056,N_35862,N_35837);
nor U36057 (N_36057,N_35933,N_35874);
or U36058 (N_36058,N_35819,N_35752);
nor U36059 (N_36059,N_35817,N_35828);
nor U36060 (N_36060,N_35794,N_35814);
or U36061 (N_36061,N_35934,N_35831);
xnor U36062 (N_36062,N_35918,N_35750);
nand U36063 (N_36063,N_35791,N_35847);
nand U36064 (N_36064,N_35762,N_35820);
xor U36065 (N_36065,N_35753,N_35796);
nand U36066 (N_36066,N_35903,N_35915);
nand U36067 (N_36067,N_35984,N_35922);
nor U36068 (N_36068,N_35997,N_35938);
nand U36069 (N_36069,N_35878,N_35824);
or U36070 (N_36070,N_35948,N_35836);
nand U36071 (N_36071,N_35764,N_35769);
or U36072 (N_36072,N_35953,N_35959);
xnor U36073 (N_36073,N_35795,N_35857);
nor U36074 (N_36074,N_35871,N_35909);
nor U36075 (N_36075,N_35810,N_35802);
or U36076 (N_36076,N_35967,N_35834);
nor U36077 (N_36077,N_35782,N_35787);
or U36078 (N_36078,N_35971,N_35926);
nand U36079 (N_36079,N_35974,N_35775);
nor U36080 (N_36080,N_35935,N_35879);
nor U36081 (N_36081,N_35994,N_35945);
nand U36082 (N_36082,N_35978,N_35768);
nor U36083 (N_36083,N_35963,N_35952);
xnor U36084 (N_36084,N_35765,N_35902);
nand U36085 (N_36085,N_35844,N_35867);
xnor U36086 (N_36086,N_35958,N_35816);
and U36087 (N_36087,N_35882,N_35985);
or U36088 (N_36088,N_35968,N_35849);
or U36089 (N_36089,N_35960,N_35771);
nand U36090 (N_36090,N_35808,N_35989);
nand U36091 (N_36091,N_35941,N_35767);
and U36092 (N_36092,N_35754,N_35931);
nand U36093 (N_36093,N_35841,N_35996);
nand U36094 (N_36094,N_35937,N_35845);
and U36095 (N_36095,N_35995,N_35763);
xor U36096 (N_36096,N_35887,N_35992);
nor U36097 (N_36097,N_35950,N_35783);
and U36098 (N_36098,N_35895,N_35806);
nor U36099 (N_36099,N_35916,N_35893);
and U36100 (N_36100,N_35772,N_35793);
nor U36101 (N_36101,N_35998,N_35993);
nand U36102 (N_36102,N_35870,N_35896);
or U36103 (N_36103,N_35833,N_35786);
nor U36104 (N_36104,N_35865,N_35827);
and U36105 (N_36105,N_35890,N_35908);
nand U36106 (N_36106,N_35883,N_35875);
nand U36107 (N_36107,N_35829,N_35766);
nor U36108 (N_36108,N_35823,N_35851);
nor U36109 (N_36109,N_35873,N_35803);
and U36110 (N_36110,N_35912,N_35759);
nand U36111 (N_36111,N_35969,N_35939);
nand U36112 (N_36112,N_35835,N_35777);
and U36113 (N_36113,N_35773,N_35983);
nand U36114 (N_36114,N_35975,N_35760);
nor U36115 (N_36115,N_35979,N_35957);
nand U36116 (N_36116,N_35961,N_35943);
nor U36117 (N_36117,N_35886,N_35977);
xnor U36118 (N_36118,N_35770,N_35801);
nor U36119 (N_36119,N_35932,N_35842);
or U36120 (N_36120,N_35999,N_35825);
xnor U36121 (N_36121,N_35839,N_35784);
and U36122 (N_36122,N_35758,N_35846);
nor U36123 (N_36123,N_35917,N_35919);
nand U36124 (N_36124,N_35910,N_35906);
and U36125 (N_36125,N_35850,N_35982);
xnor U36126 (N_36126,N_35961,N_35787);
and U36127 (N_36127,N_35954,N_35924);
nand U36128 (N_36128,N_35974,N_35807);
nand U36129 (N_36129,N_35763,N_35825);
xor U36130 (N_36130,N_35987,N_35806);
xnor U36131 (N_36131,N_35849,N_35965);
nor U36132 (N_36132,N_35869,N_35752);
or U36133 (N_36133,N_35910,N_35923);
or U36134 (N_36134,N_35984,N_35811);
nor U36135 (N_36135,N_35888,N_35899);
or U36136 (N_36136,N_35916,N_35816);
xnor U36137 (N_36137,N_35924,N_35815);
xor U36138 (N_36138,N_35930,N_35804);
nor U36139 (N_36139,N_35750,N_35841);
or U36140 (N_36140,N_35934,N_35962);
nand U36141 (N_36141,N_35783,N_35963);
nand U36142 (N_36142,N_35829,N_35756);
nor U36143 (N_36143,N_35919,N_35920);
nand U36144 (N_36144,N_35835,N_35941);
nand U36145 (N_36145,N_35844,N_35951);
nor U36146 (N_36146,N_35886,N_35965);
xor U36147 (N_36147,N_35953,N_35839);
xnor U36148 (N_36148,N_35926,N_35752);
nor U36149 (N_36149,N_35881,N_35878);
nor U36150 (N_36150,N_35943,N_35826);
xnor U36151 (N_36151,N_35784,N_35835);
nor U36152 (N_36152,N_35781,N_35971);
and U36153 (N_36153,N_35757,N_35785);
or U36154 (N_36154,N_35771,N_35835);
xnor U36155 (N_36155,N_35979,N_35842);
nand U36156 (N_36156,N_35998,N_35757);
nand U36157 (N_36157,N_35938,N_35964);
or U36158 (N_36158,N_35955,N_35806);
or U36159 (N_36159,N_35904,N_35911);
or U36160 (N_36160,N_35956,N_35969);
xor U36161 (N_36161,N_35818,N_35877);
or U36162 (N_36162,N_35761,N_35908);
xnor U36163 (N_36163,N_35950,N_35785);
nor U36164 (N_36164,N_35802,N_35792);
or U36165 (N_36165,N_35949,N_35805);
xnor U36166 (N_36166,N_35812,N_35887);
nor U36167 (N_36167,N_35975,N_35808);
and U36168 (N_36168,N_35846,N_35934);
nand U36169 (N_36169,N_35757,N_35793);
and U36170 (N_36170,N_35842,N_35841);
nor U36171 (N_36171,N_35971,N_35875);
nand U36172 (N_36172,N_35892,N_35787);
and U36173 (N_36173,N_35805,N_35877);
xor U36174 (N_36174,N_35910,N_35853);
xor U36175 (N_36175,N_35954,N_35775);
or U36176 (N_36176,N_35883,N_35914);
nand U36177 (N_36177,N_35816,N_35753);
and U36178 (N_36178,N_35915,N_35884);
nor U36179 (N_36179,N_35826,N_35762);
nor U36180 (N_36180,N_35975,N_35943);
and U36181 (N_36181,N_35990,N_35783);
or U36182 (N_36182,N_35999,N_35927);
xor U36183 (N_36183,N_35955,N_35973);
or U36184 (N_36184,N_35908,N_35944);
xnor U36185 (N_36185,N_35774,N_35867);
nand U36186 (N_36186,N_35783,N_35928);
and U36187 (N_36187,N_35934,N_35810);
xor U36188 (N_36188,N_35953,N_35895);
xnor U36189 (N_36189,N_35808,N_35782);
nor U36190 (N_36190,N_35937,N_35791);
xor U36191 (N_36191,N_35955,N_35991);
nor U36192 (N_36192,N_35783,N_35828);
or U36193 (N_36193,N_35850,N_35834);
nand U36194 (N_36194,N_35830,N_35817);
and U36195 (N_36195,N_35900,N_35922);
nor U36196 (N_36196,N_35864,N_35792);
nor U36197 (N_36197,N_35799,N_35977);
xor U36198 (N_36198,N_35974,N_35898);
nand U36199 (N_36199,N_35828,N_35797);
or U36200 (N_36200,N_35904,N_35913);
or U36201 (N_36201,N_35835,N_35955);
and U36202 (N_36202,N_35837,N_35942);
xnor U36203 (N_36203,N_35816,N_35812);
or U36204 (N_36204,N_35973,N_35799);
or U36205 (N_36205,N_35817,N_35791);
xor U36206 (N_36206,N_35995,N_35923);
xnor U36207 (N_36207,N_35865,N_35916);
xnor U36208 (N_36208,N_35918,N_35839);
nor U36209 (N_36209,N_35892,N_35859);
and U36210 (N_36210,N_35762,N_35836);
nand U36211 (N_36211,N_35910,N_35843);
xnor U36212 (N_36212,N_35991,N_35806);
nand U36213 (N_36213,N_35792,N_35829);
nand U36214 (N_36214,N_35865,N_35783);
or U36215 (N_36215,N_35857,N_35751);
and U36216 (N_36216,N_35778,N_35841);
nand U36217 (N_36217,N_35802,N_35982);
nor U36218 (N_36218,N_35972,N_35765);
nand U36219 (N_36219,N_35997,N_35911);
and U36220 (N_36220,N_35829,N_35901);
and U36221 (N_36221,N_35976,N_35947);
or U36222 (N_36222,N_35987,N_35788);
or U36223 (N_36223,N_35979,N_35889);
nor U36224 (N_36224,N_35869,N_35924);
nand U36225 (N_36225,N_35999,N_35852);
and U36226 (N_36226,N_35812,N_35796);
or U36227 (N_36227,N_35832,N_35757);
xnor U36228 (N_36228,N_35883,N_35789);
xnor U36229 (N_36229,N_35836,N_35871);
xnor U36230 (N_36230,N_35989,N_35930);
xor U36231 (N_36231,N_35940,N_35884);
xor U36232 (N_36232,N_35803,N_35846);
xor U36233 (N_36233,N_35939,N_35971);
nand U36234 (N_36234,N_35777,N_35817);
and U36235 (N_36235,N_35776,N_35974);
and U36236 (N_36236,N_35990,N_35813);
and U36237 (N_36237,N_35812,N_35896);
and U36238 (N_36238,N_35902,N_35868);
nor U36239 (N_36239,N_35914,N_35768);
xor U36240 (N_36240,N_35896,N_35920);
nor U36241 (N_36241,N_35779,N_35860);
nor U36242 (N_36242,N_35999,N_35861);
and U36243 (N_36243,N_35945,N_35977);
nand U36244 (N_36244,N_35939,N_35774);
nand U36245 (N_36245,N_35987,N_35815);
nor U36246 (N_36246,N_35889,N_35846);
or U36247 (N_36247,N_35966,N_35968);
or U36248 (N_36248,N_35766,N_35867);
nand U36249 (N_36249,N_35829,N_35972);
or U36250 (N_36250,N_36146,N_36185);
nand U36251 (N_36251,N_36232,N_36019);
and U36252 (N_36252,N_36095,N_36199);
and U36253 (N_36253,N_36130,N_36048);
xnor U36254 (N_36254,N_36083,N_36025);
and U36255 (N_36255,N_36222,N_36170);
or U36256 (N_36256,N_36110,N_36078);
or U36257 (N_36257,N_36047,N_36072);
or U36258 (N_36258,N_36040,N_36049);
xor U36259 (N_36259,N_36147,N_36060);
xnor U36260 (N_36260,N_36059,N_36108);
nor U36261 (N_36261,N_36073,N_36247);
or U36262 (N_36262,N_36217,N_36223);
or U36263 (N_36263,N_36057,N_36114);
or U36264 (N_36264,N_36155,N_36142);
or U36265 (N_36265,N_36200,N_36208);
or U36266 (N_36266,N_36165,N_36103);
nand U36267 (N_36267,N_36211,N_36125);
or U36268 (N_36268,N_36192,N_36236);
or U36269 (N_36269,N_36240,N_36031);
nand U36270 (N_36270,N_36190,N_36241);
nor U36271 (N_36271,N_36037,N_36050);
nor U36272 (N_36272,N_36084,N_36118);
or U36273 (N_36273,N_36100,N_36004);
and U36274 (N_36274,N_36041,N_36184);
xnor U36275 (N_36275,N_36024,N_36226);
nand U36276 (N_36276,N_36051,N_36087);
nand U36277 (N_36277,N_36163,N_36010);
nand U36278 (N_36278,N_36138,N_36067);
or U36279 (N_36279,N_36015,N_36137);
and U36280 (N_36280,N_36066,N_36206);
and U36281 (N_36281,N_36121,N_36213);
or U36282 (N_36282,N_36055,N_36153);
nand U36283 (N_36283,N_36166,N_36180);
nor U36284 (N_36284,N_36209,N_36196);
nor U36285 (N_36285,N_36054,N_36034);
nor U36286 (N_36286,N_36104,N_36126);
and U36287 (N_36287,N_36149,N_36134);
nand U36288 (N_36288,N_36098,N_36145);
and U36289 (N_36289,N_36133,N_36000);
or U36290 (N_36290,N_36178,N_36141);
and U36291 (N_36291,N_36122,N_36007);
and U36292 (N_36292,N_36242,N_36127);
xor U36293 (N_36293,N_36008,N_36152);
and U36294 (N_36294,N_36197,N_36003);
nor U36295 (N_36295,N_36109,N_36111);
xor U36296 (N_36296,N_36071,N_36020);
or U36297 (N_36297,N_36044,N_36102);
xor U36298 (N_36298,N_36099,N_36091);
nand U36299 (N_36299,N_36002,N_36156);
and U36300 (N_36300,N_36220,N_36062);
or U36301 (N_36301,N_36117,N_36143);
or U36302 (N_36302,N_36045,N_36172);
and U36303 (N_36303,N_36245,N_36092);
nand U36304 (N_36304,N_36239,N_36177);
and U36305 (N_36305,N_36225,N_36203);
nand U36306 (N_36306,N_36173,N_36227);
xnor U36307 (N_36307,N_36120,N_36077);
and U36308 (N_36308,N_36082,N_36079);
or U36309 (N_36309,N_36248,N_36063);
xnor U36310 (N_36310,N_36161,N_36081);
nand U36311 (N_36311,N_36159,N_36115);
nor U36312 (N_36312,N_36032,N_36148);
nand U36313 (N_36313,N_36016,N_36001);
or U36314 (N_36314,N_36017,N_36097);
or U36315 (N_36315,N_36075,N_36154);
nor U36316 (N_36316,N_36119,N_36086);
or U36317 (N_36317,N_36021,N_36191);
or U36318 (N_36318,N_36135,N_36036);
and U36319 (N_36319,N_36068,N_36246);
and U36320 (N_36320,N_36136,N_36204);
xnor U36321 (N_36321,N_36090,N_36249);
xor U36322 (N_36322,N_36027,N_36006);
xor U36323 (N_36323,N_36175,N_36128);
nor U36324 (N_36324,N_36116,N_36219);
and U36325 (N_36325,N_36043,N_36129);
and U36326 (N_36326,N_36198,N_36089);
nor U36327 (N_36327,N_36131,N_36238);
or U36328 (N_36328,N_36244,N_36065);
and U36329 (N_36329,N_36224,N_36235);
and U36330 (N_36330,N_36005,N_36018);
and U36331 (N_36331,N_36076,N_36113);
nor U36332 (N_36332,N_36169,N_36174);
and U36333 (N_36333,N_36124,N_36101);
or U36334 (N_36334,N_36107,N_36088);
or U36335 (N_36335,N_36207,N_36009);
nand U36336 (N_36336,N_36061,N_36064);
nand U36337 (N_36337,N_36243,N_36053);
nand U36338 (N_36338,N_36167,N_36218);
or U36339 (N_36339,N_36123,N_36234);
xnor U36340 (N_36340,N_36038,N_36033);
nand U36341 (N_36341,N_36014,N_36189);
nor U36342 (N_36342,N_36210,N_36164);
nor U36343 (N_36343,N_36183,N_36106);
nor U36344 (N_36344,N_36158,N_36039);
or U36345 (N_36345,N_36215,N_36112);
or U36346 (N_36346,N_36212,N_36056);
xnor U36347 (N_36347,N_36221,N_36150);
nand U36348 (N_36348,N_36216,N_36080);
nor U36349 (N_36349,N_36012,N_36139);
nand U36350 (N_36350,N_36013,N_36023);
nor U36351 (N_36351,N_36035,N_36201);
nand U36352 (N_36352,N_36162,N_36214);
xor U36353 (N_36353,N_36085,N_36140);
nor U36354 (N_36354,N_36230,N_36160);
and U36355 (N_36355,N_36030,N_36029);
xnor U36356 (N_36356,N_36231,N_36193);
nand U36357 (N_36357,N_36229,N_36181);
nand U36358 (N_36358,N_36187,N_36151);
or U36359 (N_36359,N_36070,N_36093);
nand U36360 (N_36360,N_36182,N_36096);
and U36361 (N_36361,N_36074,N_36228);
xor U36362 (N_36362,N_36195,N_36011);
xor U36363 (N_36363,N_36233,N_36186);
nor U36364 (N_36364,N_36132,N_36157);
nand U36365 (N_36365,N_36026,N_36105);
xnor U36366 (N_36366,N_36179,N_36168);
and U36367 (N_36367,N_36144,N_36171);
nand U36368 (N_36368,N_36205,N_36052);
and U36369 (N_36369,N_36237,N_36094);
or U36370 (N_36370,N_36194,N_36042);
nor U36371 (N_36371,N_36069,N_36058);
nor U36372 (N_36372,N_36046,N_36028);
nand U36373 (N_36373,N_36022,N_36202);
nor U36374 (N_36374,N_36176,N_36188);
nor U36375 (N_36375,N_36150,N_36222);
xnor U36376 (N_36376,N_36088,N_36119);
and U36377 (N_36377,N_36096,N_36083);
or U36378 (N_36378,N_36117,N_36080);
xnor U36379 (N_36379,N_36072,N_36220);
nand U36380 (N_36380,N_36017,N_36018);
nor U36381 (N_36381,N_36116,N_36012);
nor U36382 (N_36382,N_36191,N_36063);
or U36383 (N_36383,N_36125,N_36068);
or U36384 (N_36384,N_36180,N_36110);
and U36385 (N_36385,N_36207,N_36150);
nand U36386 (N_36386,N_36199,N_36248);
nor U36387 (N_36387,N_36145,N_36015);
and U36388 (N_36388,N_36183,N_36203);
xor U36389 (N_36389,N_36092,N_36143);
xor U36390 (N_36390,N_36060,N_36057);
xnor U36391 (N_36391,N_36053,N_36157);
xnor U36392 (N_36392,N_36213,N_36040);
xnor U36393 (N_36393,N_36091,N_36056);
and U36394 (N_36394,N_36194,N_36033);
or U36395 (N_36395,N_36172,N_36166);
nor U36396 (N_36396,N_36226,N_36189);
nor U36397 (N_36397,N_36197,N_36049);
nor U36398 (N_36398,N_36224,N_36241);
nand U36399 (N_36399,N_36169,N_36205);
and U36400 (N_36400,N_36165,N_36076);
nand U36401 (N_36401,N_36003,N_36240);
nand U36402 (N_36402,N_36092,N_36178);
nand U36403 (N_36403,N_36067,N_36189);
xor U36404 (N_36404,N_36007,N_36045);
nor U36405 (N_36405,N_36070,N_36120);
and U36406 (N_36406,N_36047,N_36125);
nor U36407 (N_36407,N_36132,N_36092);
nand U36408 (N_36408,N_36156,N_36179);
xor U36409 (N_36409,N_36204,N_36242);
nand U36410 (N_36410,N_36101,N_36174);
nor U36411 (N_36411,N_36009,N_36119);
xor U36412 (N_36412,N_36179,N_36005);
xnor U36413 (N_36413,N_36065,N_36082);
or U36414 (N_36414,N_36153,N_36170);
xnor U36415 (N_36415,N_36090,N_36080);
xnor U36416 (N_36416,N_36242,N_36082);
nand U36417 (N_36417,N_36150,N_36188);
or U36418 (N_36418,N_36046,N_36116);
and U36419 (N_36419,N_36196,N_36178);
xor U36420 (N_36420,N_36036,N_36046);
and U36421 (N_36421,N_36117,N_36224);
nand U36422 (N_36422,N_36010,N_36204);
xnor U36423 (N_36423,N_36213,N_36131);
or U36424 (N_36424,N_36027,N_36242);
and U36425 (N_36425,N_36120,N_36018);
nand U36426 (N_36426,N_36009,N_36228);
nor U36427 (N_36427,N_36133,N_36205);
nand U36428 (N_36428,N_36142,N_36215);
or U36429 (N_36429,N_36185,N_36066);
xor U36430 (N_36430,N_36213,N_36196);
xnor U36431 (N_36431,N_36160,N_36196);
xor U36432 (N_36432,N_36094,N_36143);
nor U36433 (N_36433,N_36131,N_36230);
xnor U36434 (N_36434,N_36076,N_36121);
nand U36435 (N_36435,N_36119,N_36186);
nor U36436 (N_36436,N_36211,N_36192);
nor U36437 (N_36437,N_36069,N_36090);
xor U36438 (N_36438,N_36190,N_36145);
nor U36439 (N_36439,N_36236,N_36180);
and U36440 (N_36440,N_36062,N_36219);
xor U36441 (N_36441,N_36076,N_36018);
and U36442 (N_36442,N_36219,N_36242);
xor U36443 (N_36443,N_36005,N_36171);
xnor U36444 (N_36444,N_36190,N_36142);
nand U36445 (N_36445,N_36190,N_36132);
nand U36446 (N_36446,N_36001,N_36137);
xnor U36447 (N_36447,N_36030,N_36101);
nor U36448 (N_36448,N_36126,N_36071);
nand U36449 (N_36449,N_36014,N_36084);
nand U36450 (N_36450,N_36027,N_36020);
nand U36451 (N_36451,N_36218,N_36247);
and U36452 (N_36452,N_36161,N_36128);
xnor U36453 (N_36453,N_36017,N_36014);
nor U36454 (N_36454,N_36030,N_36110);
or U36455 (N_36455,N_36245,N_36065);
nand U36456 (N_36456,N_36034,N_36081);
nor U36457 (N_36457,N_36229,N_36199);
xor U36458 (N_36458,N_36110,N_36233);
xnor U36459 (N_36459,N_36195,N_36022);
and U36460 (N_36460,N_36055,N_36120);
xor U36461 (N_36461,N_36070,N_36150);
nand U36462 (N_36462,N_36014,N_36201);
and U36463 (N_36463,N_36246,N_36154);
and U36464 (N_36464,N_36039,N_36012);
nand U36465 (N_36465,N_36104,N_36206);
nor U36466 (N_36466,N_36169,N_36170);
nand U36467 (N_36467,N_36145,N_36076);
nor U36468 (N_36468,N_36045,N_36204);
nor U36469 (N_36469,N_36197,N_36227);
nand U36470 (N_36470,N_36245,N_36190);
or U36471 (N_36471,N_36074,N_36243);
xor U36472 (N_36472,N_36223,N_36103);
nand U36473 (N_36473,N_36144,N_36088);
nand U36474 (N_36474,N_36187,N_36144);
nand U36475 (N_36475,N_36198,N_36032);
xnor U36476 (N_36476,N_36001,N_36167);
and U36477 (N_36477,N_36007,N_36247);
and U36478 (N_36478,N_36041,N_36238);
nor U36479 (N_36479,N_36163,N_36162);
xnor U36480 (N_36480,N_36141,N_36173);
or U36481 (N_36481,N_36162,N_36068);
or U36482 (N_36482,N_36048,N_36001);
nor U36483 (N_36483,N_36237,N_36178);
or U36484 (N_36484,N_36197,N_36050);
or U36485 (N_36485,N_36205,N_36114);
or U36486 (N_36486,N_36239,N_36058);
nor U36487 (N_36487,N_36121,N_36102);
nor U36488 (N_36488,N_36020,N_36073);
xnor U36489 (N_36489,N_36197,N_36092);
or U36490 (N_36490,N_36157,N_36052);
nand U36491 (N_36491,N_36096,N_36068);
nand U36492 (N_36492,N_36176,N_36107);
nand U36493 (N_36493,N_36199,N_36194);
nand U36494 (N_36494,N_36017,N_36243);
nand U36495 (N_36495,N_36089,N_36077);
xor U36496 (N_36496,N_36100,N_36115);
nor U36497 (N_36497,N_36205,N_36187);
nand U36498 (N_36498,N_36137,N_36019);
nor U36499 (N_36499,N_36027,N_36120);
xnor U36500 (N_36500,N_36488,N_36429);
nor U36501 (N_36501,N_36331,N_36321);
or U36502 (N_36502,N_36337,N_36317);
and U36503 (N_36503,N_36348,N_36436);
nand U36504 (N_36504,N_36487,N_36334);
nor U36505 (N_36505,N_36485,N_36373);
nor U36506 (N_36506,N_36264,N_36390);
and U36507 (N_36507,N_36423,N_36292);
or U36508 (N_36508,N_36343,N_36335);
xor U36509 (N_36509,N_36405,N_36428);
xnor U36510 (N_36510,N_36283,N_36445);
nor U36511 (N_36511,N_36290,N_36346);
nor U36512 (N_36512,N_36320,N_36288);
and U36513 (N_36513,N_36456,N_36457);
nand U36514 (N_36514,N_36276,N_36257);
nor U36515 (N_36515,N_36496,N_36359);
nand U36516 (N_36516,N_36322,N_36280);
nand U36517 (N_36517,N_36284,N_36260);
xnor U36518 (N_36518,N_36493,N_36427);
xnor U36519 (N_36519,N_36294,N_36384);
nand U36520 (N_36520,N_36286,N_36449);
xor U36521 (N_36521,N_36266,N_36250);
xor U36522 (N_36522,N_36259,N_36267);
nand U36523 (N_36523,N_36459,N_36497);
nand U36524 (N_36524,N_36389,N_36361);
xor U36525 (N_36525,N_36467,N_36351);
nor U36526 (N_36526,N_36491,N_36375);
and U36527 (N_36527,N_36347,N_36352);
nand U36528 (N_36528,N_36304,N_36470);
and U36529 (N_36529,N_36480,N_36499);
and U36530 (N_36530,N_36476,N_36446);
or U36531 (N_36531,N_36377,N_36272);
and U36532 (N_36532,N_36430,N_36297);
nand U36533 (N_36533,N_36291,N_36270);
and U36534 (N_36534,N_36329,N_36438);
xor U36535 (N_36535,N_36349,N_36385);
or U36536 (N_36536,N_36313,N_36439);
and U36537 (N_36537,N_36401,N_36357);
xor U36538 (N_36538,N_36412,N_36444);
and U36539 (N_36539,N_36269,N_36400);
and U36540 (N_36540,N_36353,N_36378);
or U36541 (N_36541,N_36471,N_36342);
nor U36542 (N_36542,N_36364,N_36255);
or U36543 (N_36543,N_36299,N_36425);
xnor U36544 (N_36544,N_36447,N_36277);
and U36545 (N_36545,N_36475,N_36302);
or U36546 (N_36546,N_36417,N_36363);
and U36547 (N_36547,N_36473,N_36376);
or U36548 (N_36548,N_36323,N_36479);
nor U36549 (N_36549,N_36455,N_36381);
nor U36550 (N_36550,N_36422,N_36298);
nand U36551 (N_36551,N_36490,N_36339);
nand U36552 (N_36552,N_36413,N_36311);
nor U36553 (N_36553,N_36395,N_36251);
or U36554 (N_36554,N_36486,N_36345);
nor U36555 (N_36555,N_36482,N_36397);
or U36556 (N_36556,N_36319,N_36281);
xor U36557 (N_36557,N_36415,N_36484);
xnor U36558 (N_36558,N_36492,N_36388);
and U36559 (N_36559,N_36426,N_36287);
or U36560 (N_36560,N_36399,N_36443);
and U36561 (N_36561,N_36461,N_36409);
or U36562 (N_36562,N_36263,N_36418);
xor U36563 (N_36563,N_36495,N_36282);
xnor U36564 (N_36564,N_36396,N_36458);
nor U36565 (N_36565,N_36421,N_36442);
nand U36566 (N_36566,N_36453,N_36391);
or U36567 (N_36567,N_36408,N_36498);
nor U36568 (N_36568,N_36474,N_36275);
nand U36569 (N_36569,N_36296,N_36465);
or U36570 (N_36570,N_36338,N_36424);
and U36571 (N_36571,N_36316,N_36410);
or U36572 (N_36572,N_36318,N_36340);
nor U36573 (N_36573,N_36308,N_36472);
and U36574 (N_36574,N_36365,N_36289);
nor U36575 (N_36575,N_36411,N_36440);
xor U36576 (N_36576,N_36301,N_36354);
nor U36577 (N_36577,N_36450,N_36402);
xor U36578 (N_36578,N_36326,N_36285);
xor U36579 (N_36579,N_36256,N_36307);
or U36580 (N_36580,N_36360,N_36383);
or U36581 (N_36581,N_36435,N_36262);
or U36582 (N_36582,N_36494,N_36483);
and U36583 (N_36583,N_36466,N_36481);
and U36584 (N_36584,N_36303,N_36437);
nand U36585 (N_36585,N_36394,N_36478);
and U36586 (N_36586,N_36477,N_36252);
nor U36587 (N_36587,N_36367,N_36268);
or U36588 (N_36588,N_36419,N_36464);
and U36589 (N_36589,N_36382,N_36452);
or U36590 (N_36590,N_36404,N_36386);
or U36591 (N_36591,N_36300,N_36392);
xnor U36592 (N_36592,N_36315,N_36431);
and U36593 (N_36593,N_36274,N_36258);
nand U36594 (N_36594,N_36306,N_36432);
xnor U36595 (N_36595,N_36253,N_36489);
nor U36596 (N_36596,N_36309,N_36368);
nor U36597 (N_36597,N_36310,N_36324);
and U36598 (N_36598,N_36393,N_36279);
and U36599 (N_36599,N_36332,N_36398);
xnor U36600 (N_36600,N_36463,N_36403);
nand U36601 (N_36601,N_36407,N_36325);
nand U36602 (N_36602,N_36460,N_36265);
and U36603 (N_36603,N_36333,N_36341);
and U36604 (N_36604,N_36305,N_36271);
xnor U36605 (N_36605,N_36330,N_36350);
xnor U36606 (N_36606,N_36261,N_36416);
and U36607 (N_36607,N_36420,N_36356);
and U36608 (N_36608,N_36358,N_36468);
and U36609 (N_36609,N_36355,N_36387);
xnor U36610 (N_36610,N_36374,N_36293);
nor U36611 (N_36611,N_36314,N_36278);
xor U36612 (N_36612,N_36344,N_36254);
nand U36613 (N_36613,N_36362,N_36406);
and U36614 (N_36614,N_36380,N_36414);
and U36615 (N_36615,N_36312,N_36372);
and U36616 (N_36616,N_36328,N_36273);
and U36617 (N_36617,N_36371,N_36454);
and U36618 (N_36618,N_36469,N_36369);
and U36619 (N_36619,N_36336,N_36379);
and U36620 (N_36620,N_36433,N_36370);
xnor U36621 (N_36621,N_36434,N_36441);
nor U36622 (N_36622,N_36327,N_36448);
or U36623 (N_36623,N_36462,N_36295);
nand U36624 (N_36624,N_36451,N_36366);
nand U36625 (N_36625,N_36447,N_36436);
nor U36626 (N_36626,N_36470,N_36474);
and U36627 (N_36627,N_36282,N_36468);
or U36628 (N_36628,N_36388,N_36339);
nor U36629 (N_36629,N_36475,N_36466);
or U36630 (N_36630,N_36394,N_36286);
xnor U36631 (N_36631,N_36476,N_36338);
nand U36632 (N_36632,N_36339,N_36314);
nand U36633 (N_36633,N_36452,N_36294);
and U36634 (N_36634,N_36253,N_36306);
nand U36635 (N_36635,N_36367,N_36390);
nor U36636 (N_36636,N_36324,N_36422);
or U36637 (N_36637,N_36293,N_36260);
nor U36638 (N_36638,N_36315,N_36460);
xor U36639 (N_36639,N_36432,N_36267);
and U36640 (N_36640,N_36315,N_36262);
nor U36641 (N_36641,N_36360,N_36460);
nor U36642 (N_36642,N_36350,N_36412);
and U36643 (N_36643,N_36300,N_36388);
nor U36644 (N_36644,N_36316,N_36446);
xor U36645 (N_36645,N_36342,N_36475);
nand U36646 (N_36646,N_36311,N_36315);
nand U36647 (N_36647,N_36360,N_36364);
nor U36648 (N_36648,N_36481,N_36499);
nand U36649 (N_36649,N_36481,N_36280);
nor U36650 (N_36650,N_36357,N_36303);
or U36651 (N_36651,N_36322,N_36458);
and U36652 (N_36652,N_36459,N_36275);
nand U36653 (N_36653,N_36404,N_36409);
xor U36654 (N_36654,N_36490,N_36485);
xor U36655 (N_36655,N_36393,N_36443);
and U36656 (N_36656,N_36389,N_36458);
nand U36657 (N_36657,N_36470,N_36334);
and U36658 (N_36658,N_36461,N_36275);
or U36659 (N_36659,N_36410,N_36280);
and U36660 (N_36660,N_36390,N_36323);
xor U36661 (N_36661,N_36481,N_36378);
nand U36662 (N_36662,N_36270,N_36456);
nor U36663 (N_36663,N_36343,N_36488);
or U36664 (N_36664,N_36273,N_36373);
nand U36665 (N_36665,N_36270,N_36442);
nand U36666 (N_36666,N_36343,N_36301);
nor U36667 (N_36667,N_36315,N_36285);
or U36668 (N_36668,N_36339,N_36387);
nor U36669 (N_36669,N_36328,N_36416);
and U36670 (N_36670,N_36469,N_36418);
nand U36671 (N_36671,N_36335,N_36471);
xor U36672 (N_36672,N_36279,N_36484);
and U36673 (N_36673,N_36289,N_36390);
nor U36674 (N_36674,N_36305,N_36413);
and U36675 (N_36675,N_36449,N_36279);
nor U36676 (N_36676,N_36328,N_36381);
and U36677 (N_36677,N_36480,N_36346);
nand U36678 (N_36678,N_36372,N_36378);
nand U36679 (N_36679,N_36250,N_36297);
and U36680 (N_36680,N_36289,N_36386);
or U36681 (N_36681,N_36463,N_36408);
and U36682 (N_36682,N_36316,N_36406);
xor U36683 (N_36683,N_36320,N_36310);
nor U36684 (N_36684,N_36448,N_36259);
nand U36685 (N_36685,N_36492,N_36436);
xnor U36686 (N_36686,N_36344,N_36495);
and U36687 (N_36687,N_36297,N_36434);
nor U36688 (N_36688,N_36263,N_36432);
and U36689 (N_36689,N_36287,N_36433);
or U36690 (N_36690,N_36455,N_36427);
and U36691 (N_36691,N_36375,N_36449);
xor U36692 (N_36692,N_36256,N_36352);
or U36693 (N_36693,N_36313,N_36422);
nand U36694 (N_36694,N_36447,N_36433);
xor U36695 (N_36695,N_36439,N_36362);
xnor U36696 (N_36696,N_36387,N_36299);
and U36697 (N_36697,N_36338,N_36418);
xor U36698 (N_36698,N_36438,N_36422);
xnor U36699 (N_36699,N_36289,N_36297);
nand U36700 (N_36700,N_36294,N_36293);
nor U36701 (N_36701,N_36474,N_36342);
nor U36702 (N_36702,N_36482,N_36342);
nand U36703 (N_36703,N_36455,N_36474);
nor U36704 (N_36704,N_36259,N_36282);
nand U36705 (N_36705,N_36394,N_36354);
nor U36706 (N_36706,N_36362,N_36496);
or U36707 (N_36707,N_36377,N_36267);
nor U36708 (N_36708,N_36281,N_36469);
nor U36709 (N_36709,N_36374,N_36305);
nand U36710 (N_36710,N_36412,N_36328);
nor U36711 (N_36711,N_36433,N_36489);
nor U36712 (N_36712,N_36345,N_36413);
and U36713 (N_36713,N_36388,N_36499);
nand U36714 (N_36714,N_36494,N_36291);
and U36715 (N_36715,N_36498,N_36475);
and U36716 (N_36716,N_36330,N_36406);
or U36717 (N_36717,N_36466,N_36293);
and U36718 (N_36718,N_36305,N_36294);
nand U36719 (N_36719,N_36338,N_36299);
nand U36720 (N_36720,N_36414,N_36353);
xor U36721 (N_36721,N_36415,N_36436);
and U36722 (N_36722,N_36410,N_36412);
nor U36723 (N_36723,N_36374,N_36465);
and U36724 (N_36724,N_36342,N_36279);
nand U36725 (N_36725,N_36295,N_36250);
nand U36726 (N_36726,N_36465,N_36308);
nand U36727 (N_36727,N_36336,N_36296);
or U36728 (N_36728,N_36358,N_36280);
xor U36729 (N_36729,N_36352,N_36426);
and U36730 (N_36730,N_36374,N_36277);
or U36731 (N_36731,N_36393,N_36330);
xnor U36732 (N_36732,N_36479,N_36351);
nand U36733 (N_36733,N_36499,N_36493);
xor U36734 (N_36734,N_36419,N_36272);
or U36735 (N_36735,N_36282,N_36313);
or U36736 (N_36736,N_36427,N_36439);
xor U36737 (N_36737,N_36375,N_36310);
and U36738 (N_36738,N_36449,N_36327);
and U36739 (N_36739,N_36272,N_36381);
nor U36740 (N_36740,N_36349,N_36451);
xnor U36741 (N_36741,N_36372,N_36259);
and U36742 (N_36742,N_36385,N_36443);
xnor U36743 (N_36743,N_36469,N_36288);
and U36744 (N_36744,N_36381,N_36441);
and U36745 (N_36745,N_36381,N_36386);
and U36746 (N_36746,N_36472,N_36442);
nor U36747 (N_36747,N_36308,N_36257);
nor U36748 (N_36748,N_36447,N_36253);
nand U36749 (N_36749,N_36327,N_36275);
nand U36750 (N_36750,N_36639,N_36584);
nand U36751 (N_36751,N_36730,N_36708);
and U36752 (N_36752,N_36644,N_36632);
nand U36753 (N_36753,N_36676,N_36692);
nand U36754 (N_36754,N_36694,N_36622);
and U36755 (N_36755,N_36670,N_36574);
nand U36756 (N_36756,N_36569,N_36606);
xnor U36757 (N_36757,N_36556,N_36681);
nand U36758 (N_36758,N_36700,N_36502);
nand U36759 (N_36759,N_36686,N_36646);
nand U36760 (N_36760,N_36733,N_36528);
or U36761 (N_36761,N_36548,N_36665);
and U36762 (N_36762,N_36673,N_36567);
or U36763 (N_36763,N_36672,N_36721);
or U36764 (N_36764,N_36626,N_36614);
nand U36765 (N_36765,N_36546,N_36650);
nor U36766 (N_36766,N_36581,N_36624);
nand U36767 (N_36767,N_36542,N_36679);
nand U36768 (N_36768,N_36643,N_36653);
nand U36769 (N_36769,N_36738,N_36648);
nand U36770 (N_36770,N_36531,N_36613);
and U36771 (N_36771,N_36664,N_36545);
nand U36772 (N_36772,N_36607,N_36675);
or U36773 (N_36773,N_36507,N_36683);
and U36774 (N_36774,N_36520,N_36602);
or U36775 (N_36775,N_36645,N_36580);
xor U36776 (N_36776,N_36662,N_36704);
or U36777 (N_36777,N_36635,N_36501);
nand U36778 (N_36778,N_36695,N_36717);
nor U36779 (N_36779,N_36526,N_36511);
nand U36780 (N_36780,N_36585,N_36504);
xor U36781 (N_36781,N_36699,N_36609);
nor U36782 (N_36782,N_36727,N_36718);
nand U36783 (N_36783,N_36663,N_36518);
and U36784 (N_36784,N_36570,N_36596);
and U36785 (N_36785,N_36552,N_36657);
or U36786 (N_36786,N_36568,N_36598);
nor U36787 (N_36787,N_36680,N_36521);
nand U36788 (N_36788,N_36611,N_36661);
and U36789 (N_36789,N_36538,N_36541);
xnor U36790 (N_36790,N_36740,N_36677);
and U36791 (N_36791,N_36748,N_36658);
nand U36792 (N_36792,N_36578,N_36656);
or U36793 (N_36793,N_36515,N_36642);
or U36794 (N_36794,N_36522,N_36517);
and U36795 (N_36795,N_36678,N_36557);
nor U36796 (N_36796,N_36610,N_36603);
nand U36797 (N_36797,N_36714,N_36513);
nand U36798 (N_36798,N_36636,N_36563);
nor U36799 (N_36799,N_36629,N_36737);
nand U36800 (N_36800,N_36595,N_36617);
nor U36801 (N_36801,N_36591,N_36641);
nand U36802 (N_36802,N_36638,N_36691);
nand U36803 (N_36803,N_36735,N_36640);
nor U36804 (N_36804,N_36747,N_36597);
nand U36805 (N_36805,N_36566,N_36600);
and U36806 (N_36806,N_36628,N_36734);
nor U36807 (N_36807,N_36558,N_36573);
or U36808 (N_36808,N_36529,N_36561);
and U36809 (N_36809,N_36512,N_36623);
xnor U36810 (N_36810,N_36741,N_36516);
or U36811 (N_36811,N_36729,N_36723);
and U36812 (N_36812,N_36536,N_36589);
nand U36813 (N_36813,N_36712,N_36559);
and U36814 (N_36814,N_36685,N_36533);
nand U36815 (N_36815,N_36716,N_36668);
nor U36816 (N_36816,N_36583,N_36711);
nand U36817 (N_36817,N_36746,N_36593);
or U36818 (N_36818,N_36582,N_36509);
nand U36819 (N_36819,N_36550,N_36713);
nand U36820 (N_36820,N_36621,N_36523);
nor U36821 (N_36821,N_36689,N_36633);
or U36822 (N_36822,N_36654,N_36627);
or U36823 (N_36823,N_36728,N_36722);
xnor U36824 (N_36824,N_36690,N_36736);
nor U36825 (N_36825,N_36535,N_36693);
nor U36826 (N_36826,N_36510,N_36667);
nor U36827 (N_36827,N_36587,N_36553);
or U36828 (N_36828,N_36705,N_36506);
nor U36829 (N_36829,N_36508,N_36709);
nor U36830 (N_36830,N_36549,N_36537);
or U36831 (N_36831,N_36555,N_36710);
xor U36832 (N_36832,N_36500,N_36625);
xnor U36833 (N_36833,N_36744,N_36706);
nand U36834 (N_36834,N_36575,N_36749);
nand U36835 (N_36835,N_36649,N_36539);
xnor U36836 (N_36836,N_36742,N_36588);
nand U36837 (N_36837,N_36660,N_36540);
nand U36838 (N_36838,N_36599,N_36666);
and U36839 (N_36839,N_36586,N_36590);
or U36840 (N_36840,N_36564,N_36659);
nand U36841 (N_36841,N_36696,N_36674);
and U36842 (N_36842,N_36608,N_36731);
or U36843 (N_36843,N_36620,N_36503);
xnor U36844 (N_36844,N_36572,N_36684);
or U36845 (N_36845,N_36707,N_36577);
and U36846 (N_36846,N_36701,N_36618);
nand U36847 (N_36847,N_36605,N_36615);
xor U36848 (N_36848,N_36671,N_36579);
xor U36849 (N_36849,N_36631,N_36724);
xnor U36850 (N_36850,N_36719,N_36687);
nor U36851 (N_36851,N_36519,N_36630);
xnor U36852 (N_36852,N_36505,N_36576);
and U36853 (N_36853,N_36562,N_36715);
or U36854 (N_36854,N_36698,N_36688);
or U36855 (N_36855,N_36726,N_36697);
or U36856 (N_36856,N_36612,N_36530);
nand U36857 (N_36857,N_36544,N_36652);
nand U36858 (N_36858,N_36571,N_36682);
nand U36859 (N_36859,N_36554,N_36725);
nor U36860 (N_36860,N_36702,N_36651);
and U36861 (N_36861,N_36527,N_36619);
or U36862 (N_36862,N_36547,N_36745);
or U36863 (N_36863,N_36560,N_36594);
xor U36864 (N_36864,N_36551,N_36655);
nor U36865 (N_36865,N_36592,N_36604);
nand U36866 (N_36866,N_36647,N_36732);
or U36867 (N_36867,N_36532,N_36514);
xnor U36868 (N_36868,N_36669,N_36703);
or U36869 (N_36869,N_36601,N_36743);
or U36870 (N_36870,N_36534,N_36637);
and U36871 (N_36871,N_36525,N_36616);
nor U36872 (N_36872,N_36739,N_36543);
xor U36873 (N_36873,N_36565,N_36720);
nor U36874 (N_36874,N_36524,N_36634);
and U36875 (N_36875,N_36640,N_36655);
nand U36876 (N_36876,N_36622,N_36741);
or U36877 (N_36877,N_36569,N_36675);
nor U36878 (N_36878,N_36749,N_36660);
and U36879 (N_36879,N_36520,N_36670);
or U36880 (N_36880,N_36632,N_36650);
nor U36881 (N_36881,N_36696,N_36545);
nor U36882 (N_36882,N_36631,N_36568);
xnor U36883 (N_36883,N_36712,N_36729);
nand U36884 (N_36884,N_36501,N_36748);
xnor U36885 (N_36885,N_36580,N_36563);
nand U36886 (N_36886,N_36542,N_36557);
and U36887 (N_36887,N_36675,N_36542);
xnor U36888 (N_36888,N_36646,N_36738);
nor U36889 (N_36889,N_36516,N_36655);
nor U36890 (N_36890,N_36577,N_36527);
nand U36891 (N_36891,N_36746,N_36528);
and U36892 (N_36892,N_36587,N_36571);
and U36893 (N_36893,N_36651,N_36705);
xor U36894 (N_36894,N_36734,N_36736);
nor U36895 (N_36895,N_36608,N_36712);
nor U36896 (N_36896,N_36701,N_36539);
xor U36897 (N_36897,N_36683,N_36616);
nor U36898 (N_36898,N_36728,N_36688);
nor U36899 (N_36899,N_36553,N_36564);
nor U36900 (N_36900,N_36702,N_36574);
nor U36901 (N_36901,N_36636,N_36523);
nand U36902 (N_36902,N_36690,N_36710);
nand U36903 (N_36903,N_36615,N_36684);
xor U36904 (N_36904,N_36505,N_36629);
or U36905 (N_36905,N_36579,N_36620);
nor U36906 (N_36906,N_36678,N_36577);
xnor U36907 (N_36907,N_36643,N_36567);
nor U36908 (N_36908,N_36633,N_36570);
and U36909 (N_36909,N_36583,N_36577);
or U36910 (N_36910,N_36623,N_36542);
nand U36911 (N_36911,N_36540,N_36685);
nor U36912 (N_36912,N_36645,N_36732);
nor U36913 (N_36913,N_36643,N_36556);
nor U36914 (N_36914,N_36620,N_36582);
and U36915 (N_36915,N_36561,N_36716);
nand U36916 (N_36916,N_36712,N_36604);
or U36917 (N_36917,N_36532,N_36665);
nand U36918 (N_36918,N_36586,N_36703);
and U36919 (N_36919,N_36581,N_36530);
xor U36920 (N_36920,N_36638,N_36557);
nor U36921 (N_36921,N_36570,N_36711);
or U36922 (N_36922,N_36545,N_36630);
nor U36923 (N_36923,N_36590,N_36615);
and U36924 (N_36924,N_36593,N_36596);
xnor U36925 (N_36925,N_36628,N_36540);
or U36926 (N_36926,N_36734,N_36684);
and U36927 (N_36927,N_36614,N_36576);
and U36928 (N_36928,N_36717,N_36536);
or U36929 (N_36929,N_36669,N_36625);
or U36930 (N_36930,N_36708,N_36707);
or U36931 (N_36931,N_36614,N_36567);
and U36932 (N_36932,N_36701,N_36534);
xor U36933 (N_36933,N_36580,N_36577);
xor U36934 (N_36934,N_36671,N_36728);
xnor U36935 (N_36935,N_36653,N_36682);
or U36936 (N_36936,N_36543,N_36519);
and U36937 (N_36937,N_36622,N_36527);
nor U36938 (N_36938,N_36740,N_36539);
and U36939 (N_36939,N_36550,N_36571);
or U36940 (N_36940,N_36685,N_36743);
nand U36941 (N_36941,N_36591,N_36565);
nor U36942 (N_36942,N_36741,N_36596);
or U36943 (N_36943,N_36686,N_36521);
nand U36944 (N_36944,N_36527,N_36606);
or U36945 (N_36945,N_36676,N_36746);
or U36946 (N_36946,N_36602,N_36575);
nand U36947 (N_36947,N_36589,N_36550);
and U36948 (N_36948,N_36705,N_36522);
or U36949 (N_36949,N_36565,N_36713);
nand U36950 (N_36950,N_36722,N_36537);
xnor U36951 (N_36951,N_36722,N_36686);
and U36952 (N_36952,N_36731,N_36655);
nand U36953 (N_36953,N_36663,N_36747);
nand U36954 (N_36954,N_36653,N_36734);
xor U36955 (N_36955,N_36543,N_36504);
and U36956 (N_36956,N_36672,N_36644);
nor U36957 (N_36957,N_36573,N_36692);
or U36958 (N_36958,N_36593,N_36697);
or U36959 (N_36959,N_36658,N_36540);
and U36960 (N_36960,N_36558,N_36621);
and U36961 (N_36961,N_36734,N_36703);
or U36962 (N_36962,N_36623,N_36565);
nand U36963 (N_36963,N_36646,N_36637);
and U36964 (N_36964,N_36676,N_36542);
xor U36965 (N_36965,N_36619,N_36522);
nor U36966 (N_36966,N_36610,N_36561);
or U36967 (N_36967,N_36616,N_36520);
and U36968 (N_36968,N_36587,N_36716);
or U36969 (N_36969,N_36716,N_36672);
and U36970 (N_36970,N_36626,N_36509);
xnor U36971 (N_36971,N_36522,N_36512);
nand U36972 (N_36972,N_36637,N_36689);
nor U36973 (N_36973,N_36536,N_36570);
xnor U36974 (N_36974,N_36634,N_36660);
xor U36975 (N_36975,N_36574,N_36647);
nand U36976 (N_36976,N_36710,N_36512);
xor U36977 (N_36977,N_36714,N_36607);
xor U36978 (N_36978,N_36688,N_36638);
or U36979 (N_36979,N_36558,N_36574);
xnor U36980 (N_36980,N_36501,N_36721);
and U36981 (N_36981,N_36742,N_36620);
xnor U36982 (N_36982,N_36532,N_36686);
and U36983 (N_36983,N_36733,N_36605);
and U36984 (N_36984,N_36737,N_36693);
nand U36985 (N_36985,N_36676,N_36575);
nor U36986 (N_36986,N_36741,N_36545);
nand U36987 (N_36987,N_36585,N_36712);
nand U36988 (N_36988,N_36554,N_36565);
or U36989 (N_36989,N_36629,N_36583);
nand U36990 (N_36990,N_36570,N_36589);
xnor U36991 (N_36991,N_36725,N_36687);
and U36992 (N_36992,N_36666,N_36603);
and U36993 (N_36993,N_36606,N_36728);
and U36994 (N_36994,N_36544,N_36545);
xnor U36995 (N_36995,N_36739,N_36701);
or U36996 (N_36996,N_36620,N_36585);
xnor U36997 (N_36997,N_36604,N_36662);
nand U36998 (N_36998,N_36633,N_36726);
xnor U36999 (N_36999,N_36578,N_36681);
nor U37000 (N_37000,N_36875,N_36815);
xnor U37001 (N_37001,N_36823,N_36996);
xor U37002 (N_37002,N_36844,N_36828);
xnor U37003 (N_37003,N_36765,N_36910);
nor U37004 (N_37004,N_36973,N_36798);
nand U37005 (N_37005,N_36860,N_36892);
or U37006 (N_37006,N_36976,N_36997);
nor U37007 (N_37007,N_36877,N_36781);
xor U37008 (N_37008,N_36836,N_36893);
xnor U37009 (N_37009,N_36943,N_36852);
and U37010 (N_37010,N_36822,N_36995);
nand U37011 (N_37011,N_36988,N_36948);
or U37012 (N_37012,N_36794,N_36767);
nand U37013 (N_37013,N_36946,N_36944);
nor U37014 (N_37014,N_36920,N_36945);
nand U37015 (N_37015,N_36799,N_36842);
or U37016 (N_37016,N_36766,N_36957);
xor U37017 (N_37017,N_36806,N_36797);
nor U37018 (N_37018,N_36991,N_36887);
nor U37019 (N_37019,N_36950,N_36763);
nor U37020 (N_37020,N_36753,N_36812);
nand U37021 (N_37021,N_36999,N_36856);
nand U37022 (N_37022,N_36888,N_36963);
or U37023 (N_37023,N_36977,N_36863);
nor U37024 (N_37024,N_36845,N_36961);
and U37025 (N_37025,N_36974,N_36898);
and U37026 (N_37026,N_36838,N_36847);
or U37027 (N_37027,N_36962,N_36850);
and U37028 (N_37028,N_36903,N_36855);
or U37029 (N_37029,N_36992,N_36938);
and U37030 (N_37030,N_36866,N_36993);
or U37031 (N_37031,N_36909,N_36921);
xor U37032 (N_37032,N_36897,N_36879);
and U37033 (N_37033,N_36861,N_36759);
xnor U37034 (N_37034,N_36762,N_36810);
nand U37035 (N_37035,N_36800,N_36784);
nor U37036 (N_37036,N_36965,N_36779);
or U37037 (N_37037,N_36785,N_36830);
or U37038 (N_37038,N_36827,N_36918);
or U37039 (N_37039,N_36883,N_36956);
and U37040 (N_37040,N_36876,N_36777);
and U37041 (N_37041,N_36834,N_36872);
nor U37042 (N_37042,N_36839,N_36813);
nor U37043 (N_37043,N_36843,N_36979);
nor U37044 (N_37044,N_36841,N_36791);
nand U37045 (N_37045,N_36966,N_36868);
and U37046 (N_37046,N_36922,N_36801);
xnor U37047 (N_37047,N_36899,N_36953);
nor U37048 (N_37048,N_36930,N_36871);
nand U37049 (N_37049,N_36831,N_36934);
nor U37050 (N_37050,N_36951,N_36870);
nor U37051 (N_37051,N_36837,N_36833);
nor U37052 (N_37052,N_36981,N_36771);
or U37053 (N_37053,N_36895,N_36983);
and U37054 (N_37054,N_36817,N_36774);
xnor U37055 (N_37055,N_36886,N_36751);
xnor U37056 (N_37056,N_36756,N_36885);
xor U37057 (N_37057,N_36890,N_36937);
nand U37058 (N_37058,N_36928,N_36964);
nand U37059 (N_37059,N_36873,N_36780);
and U37060 (N_37060,N_36939,N_36755);
nand U37061 (N_37061,N_36935,N_36805);
or U37062 (N_37062,N_36969,N_36959);
nand U37063 (N_37063,N_36859,N_36757);
nand U37064 (N_37064,N_36835,N_36960);
or U37065 (N_37065,N_36804,N_36936);
xnor U37066 (N_37066,N_36840,N_36915);
xnor U37067 (N_37067,N_36750,N_36994);
xnor U37068 (N_37068,N_36891,N_36929);
nand U37069 (N_37069,N_36792,N_36754);
xor U37070 (N_37070,N_36923,N_36807);
nor U37071 (N_37071,N_36772,N_36987);
nand U37072 (N_37072,N_36821,N_36958);
nand U37073 (N_37073,N_36865,N_36814);
and U37074 (N_37074,N_36896,N_36914);
nor U37075 (N_37075,N_36968,N_36954);
nand U37076 (N_37076,N_36940,N_36990);
and U37077 (N_37077,N_36829,N_36917);
nand U37078 (N_37078,N_36808,N_36776);
nand U37079 (N_37079,N_36913,N_36760);
nor U37080 (N_37080,N_36971,N_36816);
nor U37081 (N_37081,N_36911,N_36846);
and U37082 (N_37082,N_36789,N_36884);
or U37083 (N_37083,N_36775,N_36933);
and U37084 (N_37084,N_36878,N_36819);
or U37085 (N_37085,N_36824,N_36985);
nor U37086 (N_37086,N_36849,N_36809);
nor U37087 (N_37087,N_36924,N_36952);
nand U37088 (N_37088,N_36802,N_36906);
nor U37089 (N_37089,N_36787,N_36980);
and U37090 (N_37090,N_36818,N_36978);
and U37091 (N_37091,N_36778,N_36881);
nor U37092 (N_37092,N_36848,N_36882);
nand U37093 (N_37093,N_36874,N_36826);
xor U37094 (N_37094,N_36925,N_36773);
xnor U37095 (N_37095,N_36904,N_36908);
xor U37096 (N_37096,N_36768,N_36912);
xor U37097 (N_37097,N_36786,N_36867);
nand U37098 (N_37098,N_36752,N_36782);
xor U37099 (N_37099,N_36982,N_36864);
and U37100 (N_37100,N_36955,N_36947);
or U37101 (N_37101,N_36931,N_36770);
or U37102 (N_37102,N_36790,N_36764);
nand U37103 (N_37103,N_36967,N_36862);
or U37104 (N_37104,N_36907,N_36793);
and U37105 (N_37105,N_36894,N_36820);
nor U37106 (N_37106,N_36942,N_36927);
nor U37107 (N_37107,N_36975,N_36880);
nor U37108 (N_37108,N_36783,N_36796);
and U37109 (N_37109,N_36832,N_36788);
and U37110 (N_37110,N_36949,N_36854);
xnor U37111 (N_37111,N_36919,N_36916);
nor U37112 (N_37112,N_36905,N_36972);
nor U37113 (N_37113,N_36984,N_36857);
nor U37114 (N_37114,N_36758,N_36803);
or U37115 (N_37115,N_36986,N_36795);
or U37116 (N_37116,N_36941,N_36970);
xor U37117 (N_37117,N_36900,N_36998);
nand U37118 (N_37118,N_36858,N_36902);
and U37119 (N_37119,N_36889,N_36769);
nor U37120 (N_37120,N_36989,N_36869);
xnor U37121 (N_37121,N_36932,N_36901);
nor U37122 (N_37122,N_36811,N_36761);
nand U37123 (N_37123,N_36926,N_36853);
nor U37124 (N_37124,N_36851,N_36825);
xor U37125 (N_37125,N_36894,N_36760);
nor U37126 (N_37126,N_36859,N_36872);
nor U37127 (N_37127,N_36842,N_36988);
or U37128 (N_37128,N_36833,N_36901);
nand U37129 (N_37129,N_36809,N_36784);
or U37130 (N_37130,N_36985,N_36907);
and U37131 (N_37131,N_36885,N_36922);
or U37132 (N_37132,N_36989,N_36921);
and U37133 (N_37133,N_36767,N_36753);
xor U37134 (N_37134,N_36968,N_36823);
nor U37135 (N_37135,N_36951,N_36871);
nand U37136 (N_37136,N_36905,N_36899);
nor U37137 (N_37137,N_36773,N_36838);
nand U37138 (N_37138,N_36965,N_36901);
and U37139 (N_37139,N_36965,N_36767);
nand U37140 (N_37140,N_36850,N_36941);
nor U37141 (N_37141,N_36937,N_36761);
and U37142 (N_37142,N_36762,N_36882);
and U37143 (N_37143,N_36980,N_36969);
nand U37144 (N_37144,N_36777,N_36909);
or U37145 (N_37145,N_36996,N_36750);
nand U37146 (N_37146,N_36872,N_36758);
and U37147 (N_37147,N_36859,N_36940);
xnor U37148 (N_37148,N_36821,N_36893);
xnor U37149 (N_37149,N_36969,N_36861);
xor U37150 (N_37150,N_36953,N_36981);
or U37151 (N_37151,N_36902,N_36918);
xnor U37152 (N_37152,N_36798,N_36861);
nand U37153 (N_37153,N_36976,N_36864);
or U37154 (N_37154,N_36904,N_36832);
nand U37155 (N_37155,N_36851,N_36801);
xnor U37156 (N_37156,N_36915,N_36864);
and U37157 (N_37157,N_36902,N_36974);
or U37158 (N_37158,N_36992,N_36828);
and U37159 (N_37159,N_36859,N_36765);
xnor U37160 (N_37160,N_36887,N_36809);
and U37161 (N_37161,N_36858,N_36815);
nor U37162 (N_37162,N_36808,N_36908);
and U37163 (N_37163,N_36888,N_36779);
nor U37164 (N_37164,N_36753,N_36947);
nor U37165 (N_37165,N_36928,N_36820);
nand U37166 (N_37166,N_36912,N_36951);
nor U37167 (N_37167,N_36962,N_36976);
nand U37168 (N_37168,N_36882,N_36969);
nor U37169 (N_37169,N_36875,N_36896);
nor U37170 (N_37170,N_36950,N_36937);
nor U37171 (N_37171,N_36831,N_36834);
nand U37172 (N_37172,N_36791,N_36777);
xnor U37173 (N_37173,N_36903,N_36864);
and U37174 (N_37174,N_36953,N_36753);
and U37175 (N_37175,N_36803,N_36785);
xnor U37176 (N_37176,N_36772,N_36810);
xnor U37177 (N_37177,N_36990,N_36899);
nor U37178 (N_37178,N_36853,N_36829);
nor U37179 (N_37179,N_36759,N_36842);
xor U37180 (N_37180,N_36768,N_36828);
and U37181 (N_37181,N_36888,N_36948);
nand U37182 (N_37182,N_36954,N_36946);
and U37183 (N_37183,N_36915,N_36830);
and U37184 (N_37184,N_36986,N_36758);
nor U37185 (N_37185,N_36826,N_36864);
xnor U37186 (N_37186,N_36815,N_36965);
xor U37187 (N_37187,N_36841,N_36854);
xor U37188 (N_37188,N_36779,N_36985);
or U37189 (N_37189,N_36970,N_36813);
and U37190 (N_37190,N_36979,N_36898);
or U37191 (N_37191,N_36947,N_36993);
nor U37192 (N_37192,N_36961,N_36830);
xor U37193 (N_37193,N_36978,N_36927);
nor U37194 (N_37194,N_36997,N_36807);
nor U37195 (N_37195,N_36909,N_36831);
or U37196 (N_37196,N_36762,N_36930);
xor U37197 (N_37197,N_36924,N_36856);
or U37198 (N_37198,N_36920,N_36891);
xnor U37199 (N_37199,N_36877,N_36837);
xor U37200 (N_37200,N_36911,N_36782);
nand U37201 (N_37201,N_36980,N_36943);
or U37202 (N_37202,N_36992,N_36876);
xor U37203 (N_37203,N_36940,N_36773);
or U37204 (N_37204,N_36833,N_36836);
nand U37205 (N_37205,N_36986,N_36806);
xnor U37206 (N_37206,N_36975,N_36836);
nor U37207 (N_37207,N_36999,N_36851);
nor U37208 (N_37208,N_36827,N_36968);
and U37209 (N_37209,N_36868,N_36795);
xor U37210 (N_37210,N_36832,N_36839);
nor U37211 (N_37211,N_36916,N_36840);
nand U37212 (N_37212,N_36852,N_36942);
nor U37213 (N_37213,N_36780,N_36968);
and U37214 (N_37214,N_36867,N_36953);
or U37215 (N_37215,N_36757,N_36968);
nor U37216 (N_37216,N_36963,N_36786);
nor U37217 (N_37217,N_36793,N_36909);
nand U37218 (N_37218,N_36764,N_36763);
or U37219 (N_37219,N_36762,N_36897);
xor U37220 (N_37220,N_36823,N_36870);
and U37221 (N_37221,N_36817,N_36819);
nor U37222 (N_37222,N_36874,N_36919);
xor U37223 (N_37223,N_36776,N_36904);
nand U37224 (N_37224,N_36907,N_36903);
xnor U37225 (N_37225,N_36768,N_36856);
xor U37226 (N_37226,N_36846,N_36840);
nor U37227 (N_37227,N_36869,N_36935);
nor U37228 (N_37228,N_36842,N_36916);
nor U37229 (N_37229,N_36969,N_36847);
or U37230 (N_37230,N_36892,N_36763);
nor U37231 (N_37231,N_36764,N_36880);
xnor U37232 (N_37232,N_36829,N_36905);
nor U37233 (N_37233,N_36937,N_36906);
or U37234 (N_37234,N_36909,N_36769);
nor U37235 (N_37235,N_36752,N_36755);
and U37236 (N_37236,N_36818,N_36808);
or U37237 (N_37237,N_36968,N_36751);
and U37238 (N_37238,N_36900,N_36863);
nor U37239 (N_37239,N_36974,N_36892);
xor U37240 (N_37240,N_36929,N_36967);
or U37241 (N_37241,N_36917,N_36927);
and U37242 (N_37242,N_36779,N_36979);
xnor U37243 (N_37243,N_36795,N_36809);
or U37244 (N_37244,N_36835,N_36887);
xnor U37245 (N_37245,N_36945,N_36921);
xnor U37246 (N_37246,N_36797,N_36792);
xnor U37247 (N_37247,N_36960,N_36787);
xor U37248 (N_37248,N_36750,N_36919);
nor U37249 (N_37249,N_36872,N_36922);
nand U37250 (N_37250,N_37122,N_37178);
or U37251 (N_37251,N_37221,N_37154);
nor U37252 (N_37252,N_37160,N_37225);
or U37253 (N_37253,N_37132,N_37170);
nor U37254 (N_37254,N_37049,N_37103);
xnor U37255 (N_37255,N_37097,N_37030);
xor U37256 (N_37256,N_37055,N_37077);
and U37257 (N_37257,N_37022,N_37151);
and U37258 (N_37258,N_37102,N_37156);
xnor U37259 (N_37259,N_37084,N_37241);
xor U37260 (N_37260,N_37012,N_37153);
xor U37261 (N_37261,N_37107,N_37139);
and U37262 (N_37262,N_37075,N_37138);
nor U37263 (N_37263,N_37167,N_37215);
or U37264 (N_37264,N_37029,N_37050);
xnor U37265 (N_37265,N_37141,N_37010);
nor U37266 (N_37266,N_37190,N_37105);
xor U37267 (N_37267,N_37112,N_37203);
and U37268 (N_37268,N_37155,N_37180);
nor U37269 (N_37269,N_37004,N_37024);
xnor U37270 (N_37270,N_37230,N_37109);
or U37271 (N_37271,N_37043,N_37249);
nor U37272 (N_37272,N_37080,N_37071);
nand U37273 (N_37273,N_37235,N_37015);
nand U37274 (N_37274,N_37014,N_37161);
or U37275 (N_37275,N_37066,N_37032);
nand U37276 (N_37276,N_37159,N_37150);
and U37277 (N_37277,N_37248,N_37130);
nand U37278 (N_37278,N_37128,N_37088);
and U37279 (N_37279,N_37117,N_37184);
and U37280 (N_37280,N_37006,N_37200);
or U37281 (N_37281,N_37134,N_37183);
nor U37282 (N_37282,N_37202,N_37121);
and U37283 (N_37283,N_37100,N_37091);
nor U37284 (N_37284,N_37101,N_37174);
nand U37285 (N_37285,N_37229,N_37042);
or U37286 (N_37286,N_37137,N_37094);
or U37287 (N_37287,N_37240,N_37162);
xor U37288 (N_37288,N_37168,N_37228);
or U37289 (N_37289,N_37211,N_37172);
and U37290 (N_37290,N_37152,N_37069);
or U37291 (N_37291,N_37096,N_37163);
nor U37292 (N_37292,N_37058,N_37036);
xor U37293 (N_37293,N_37019,N_37199);
xnor U37294 (N_37294,N_37243,N_37237);
nand U37295 (N_37295,N_37089,N_37166);
xnor U37296 (N_37296,N_37081,N_37171);
and U37297 (N_37297,N_37108,N_37233);
nand U37298 (N_37298,N_37035,N_37148);
or U37299 (N_37299,N_37198,N_37245);
xnor U37300 (N_37300,N_37057,N_37149);
nand U37301 (N_37301,N_37104,N_37223);
nand U37302 (N_37302,N_37064,N_37095);
and U37303 (N_37303,N_37113,N_37188);
xnor U37304 (N_37304,N_37186,N_37169);
or U37305 (N_37305,N_37244,N_37195);
and U37306 (N_37306,N_37085,N_37083);
and U37307 (N_37307,N_37191,N_37118);
nor U37308 (N_37308,N_37142,N_37189);
xor U37309 (N_37309,N_37158,N_37079);
or U37310 (N_37310,N_37187,N_37067);
xnor U37311 (N_37311,N_37034,N_37060);
or U37312 (N_37312,N_37226,N_37125);
xnor U37313 (N_37313,N_37143,N_37236);
or U37314 (N_37314,N_37216,N_37000);
nand U37315 (N_37315,N_37037,N_37059);
nor U37316 (N_37316,N_37051,N_37246);
and U37317 (N_37317,N_37056,N_37192);
nand U37318 (N_37318,N_37007,N_37013);
and U37319 (N_37319,N_37129,N_37041);
xnor U37320 (N_37320,N_37238,N_37214);
nor U37321 (N_37321,N_37026,N_37011);
and U37322 (N_37322,N_37193,N_37028);
nor U37323 (N_37323,N_37205,N_37092);
nor U37324 (N_37324,N_37082,N_37005);
nand U37325 (N_37325,N_37086,N_37123);
or U37326 (N_37326,N_37234,N_37023);
and U37327 (N_37327,N_37027,N_37076);
nand U37328 (N_37328,N_37115,N_37207);
and U37329 (N_37329,N_37213,N_37073);
nand U37330 (N_37330,N_37197,N_37031);
or U37331 (N_37331,N_37247,N_37093);
nor U37332 (N_37332,N_37218,N_37144);
nand U37333 (N_37333,N_37220,N_37106);
nand U37334 (N_37334,N_37176,N_37116);
xnor U37335 (N_37335,N_37018,N_37127);
nand U37336 (N_37336,N_37099,N_37146);
and U37337 (N_37337,N_37133,N_37157);
xor U37338 (N_37338,N_37124,N_37061);
nand U37339 (N_37339,N_37017,N_37074);
xnor U37340 (N_37340,N_37140,N_37111);
or U37341 (N_37341,N_37078,N_37208);
xor U37342 (N_37342,N_37063,N_37048);
nand U37343 (N_37343,N_37204,N_37131);
or U37344 (N_37344,N_37212,N_37025);
or U37345 (N_37345,N_37185,N_37045);
nor U37346 (N_37346,N_37072,N_37239);
nor U37347 (N_37347,N_37219,N_37009);
and U37348 (N_37348,N_37175,N_37016);
or U37349 (N_37349,N_37054,N_37165);
nand U37350 (N_37350,N_37177,N_37065);
xnor U37351 (N_37351,N_37206,N_37003);
and U37352 (N_37352,N_37053,N_37222);
xor U37353 (N_37353,N_37052,N_37098);
nand U37354 (N_37354,N_37232,N_37145);
and U37355 (N_37355,N_37194,N_37090);
or U37356 (N_37356,N_37068,N_37008);
nand U37357 (N_37357,N_37040,N_37001);
nand U37358 (N_37358,N_37181,N_37047);
or U37359 (N_37359,N_37173,N_37209);
xor U37360 (N_37360,N_37119,N_37217);
xnor U37361 (N_37361,N_37002,N_37044);
and U37362 (N_37362,N_37136,N_37224);
and U37363 (N_37363,N_37114,N_37062);
nor U37364 (N_37364,N_37164,N_37242);
nor U37365 (N_37365,N_37126,N_37120);
or U37366 (N_37366,N_37033,N_37210);
nor U37367 (N_37367,N_37231,N_37021);
or U37368 (N_37368,N_37201,N_37147);
nand U37369 (N_37369,N_37135,N_37038);
or U37370 (N_37370,N_37110,N_37179);
and U37371 (N_37371,N_37196,N_37046);
xnor U37372 (N_37372,N_37087,N_37070);
xor U37373 (N_37373,N_37020,N_37182);
and U37374 (N_37374,N_37227,N_37039);
or U37375 (N_37375,N_37212,N_37190);
xor U37376 (N_37376,N_37074,N_37093);
or U37377 (N_37377,N_37031,N_37223);
or U37378 (N_37378,N_37040,N_37083);
nor U37379 (N_37379,N_37053,N_37156);
xor U37380 (N_37380,N_37154,N_37128);
nand U37381 (N_37381,N_37060,N_37132);
and U37382 (N_37382,N_37191,N_37116);
nor U37383 (N_37383,N_37047,N_37112);
nor U37384 (N_37384,N_37052,N_37229);
nand U37385 (N_37385,N_37124,N_37008);
nor U37386 (N_37386,N_37078,N_37032);
xor U37387 (N_37387,N_37128,N_37062);
nand U37388 (N_37388,N_37028,N_37002);
xnor U37389 (N_37389,N_37123,N_37026);
nand U37390 (N_37390,N_37211,N_37225);
and U37391 (N_37391,N_37233,N_37069);
nand U37392 (N_37392,N_37112,N_37027);
xnor U37393 (N_37393,N_37195,N_37191);
nor U37394 (N_37394,N_37108,N_37193);
nor U37395 (N_37395,N_37082,N_37170);
xor U37396 (N_37396,N_37243,N_37151);
or U37397 (N_37397,N_37043,N_37041);
nand U37398 (N_37398,N_37178,N_37040);
or U37399 (N_37399,N_37169,N_37106);
and U37400 (N_37400,N_37237,N_37226);
nand U37401 (N_37401,N_37061,N_37050);
or U37402 (N_37402,N_37174,N_37031);
xor U37403 (N_37403,N_37113,N_37121);
and U37404 (N_37404,N_37069,N_37146);
and U37405 (N_37405,N_37167,N_37041);
and U37406 (N_37406,N_37211,N_37049);
or U37407 (N_37407,N_37247,N_37207);
or U37408 (N_37408,N_37043,N_37108);
and U37409 (N_37409,N_37036,N_37056);
nor U37410 (N_37410,N_37055,N_37047);
nor U37411 (N_37411,N_37097,N_37035);
nand U37412 (N_37412,N_37132,N_37162);
xor U37413 (N_37413,N_37084,N_37190);
nor U37414 (N_37414,N_37170,N_37055);
xnor U37415 (N_37415,N_37202,N_37072);
xor U37416 (N_37416,N_37026,N_37146);
or U37417 (N_37417,N_37104,N_37076);
nand U37418 (N_37418,N_37094,N_37030);
and U37419 (N_37419,N_37049,N_37091);
nor U37420 (N_37420,N_37052,N_37191);
or U37421 (N_37421,N_37113,N_37124);
or U37422 (N_37422,N_37187,N_37229);
nor U37423 (N_37423,N_37214,N_37075);
xnor U37424 (N_37424,N_37092,N_37085);
and U37425 (N_37425,N_37133,N_37229);
xnor U37426 (N_37426,N_37219,N_37132);
or U37427 (N_37427,N_37202,N_37214);
xnor U37428 (N_37428,N_37062,N_37232);
and U37429 (N_37429,N_37016,N_37232);
nor U37430 (N_37430,N_37233,N_37073);
nor U37431 (N_37431,N_37027,N_37171);
xnor U37432 (N_37432,N_37172,N_37133);
and U37433 (N_37433,N_37086,N_37140);
or U37434 (N_37434,N_37125,N_37019);
or U37435 (N_37435,N_37166,N_37105);
or U37436 (N_37436,N_37202,N_37110);
nand U37437 (N_37437,N_37074,N_37068);
and U37438 (N_37438,N_37093,N_37148);
or U37439 (N_37439,N_37050,N_37191);
nand U37440 (N_37440,N_37223,N_37158);
or U37441 (N_37441,N_37144,N_37031);
and U37442 (N_37442,N_37198,N_37193);
xor U37443 (N_37443,N_37151,N_37140);
and U37444 (N_37444,N_37167,N_37242);
nor U37445 (N_37445,N_37004,N_37063);
or U37446 (N_37446,N_37178,N_37132);
and U37447 (N_37447,N_37006,N_37067);
nor U37448 (N_37448,N_37042,N_37129);
nand U37449 (N_37449,N_37194,N_37190);
and U37450 (N_37450,N_37122,N_37233);
xor U37451 (N_37451,N_37139,N_37167);
xnor U37452 (N_37452,N_37058,N_37115);
or U37453 (N_37453,N_37122,N_37039);
or U37454 (N_37454,N_37121,N_37153);
nand U37455 (N_37455,N_37109,N_37217);
nand U37456 (N_37456,N_37056,N_37133);
and U37457 (N_37457,N_37247,N_37233);
or U37458 (N_37458,N_37123,N_37032);
nand U37459 (N_37459,N_37233,N_37248);
xor U37460 (N_37460,N_37068,N_37217);
xnor U37461 (N_37461,N_37173,N_37034);
nand U37462 (N_37462,N_37183,N_37061);
or U37463 (N_37463,N_37223,N_37148);
nor U37464 (N_37464,N_37184,N_37002);
nor U37465 (N_37465,N_37083,N_37231);
nand U37466 (N_37466,N_37194,N_37139);
nand U37467 (N_37467,N_37210,N_37135);
and U37468 (N_37468,N_37047,N_37105);
nand U37469 (N_37469,N_37192,N_37183);
xor U37470 (N_37470,N_37014,N_37024);
or U37471 (N_37471,N_37228,N_37144);
xnor U37472 (N_37472,N_37120,N_37055);
xnor U37473 (N_37473,N_37058,N_37094);
and U37474 (N_37474,N_37233,N_37049);
xor U37475 (N_37475,N_37240,N_37137);
xnor U37476 (N_37476,N_37084,N_37202);
and U37477 (N_37477,N_37022,N_37009);
and U37478 (N_37478,N_37201,N_37235);
nand U37479 (N_37479,N_37182,N_37243);
xor U37480 (N_37480,N_37235,N_37192);
or U37481 (N_37481,N_37002,N_37227);
or U37482 (N_37482,N_37168,N_37045);
and U37483 (N_37483,N_37075,N_37197);
and U37484 (N_37484,N_37151,N_37213);
and U37485 (N_37485,N_37241,N_37015);
nor U37486 (N_37486,N_37186,N_37200);
or U37487 (N_37487,N_37075,N_37141);
nand U37488 (N_37488,N_37048,N_37180);
nand U37489 (N_37489,N_37034,N_37002);
nand U37490 (N_37490,N_37140,N_37090);
nor U37491 (N_37491,N_37139,N_37205);
nand U37492 (N_37492,N_37232,N_37214);
or U37493 (N_37493,N_37231,N_37098);
xor U37494 (N_37494,N_37162,N_37113);
nand U37495 (N_37495,N_37054,N_37173);
nand U37496 (N_37496,N_37174,N_37218);
xnor U37497 (N_37497,N_37128,N_37019);
and U37498 (N_37498,N_37210,N_37118);
nor U37499 (N_37499,N_37140,N_37236);
or U37500 (N_37500,N_37430,N_37392);
and U37501 (N_37501,N_37417,N_37299);
nand U37502 (N_37502,N_37489,N_37293);
and U37503 (N_37503,N_37446,N_37463);
xor U37504 (N_37504,N_37422,N_37384);
xnor U37505 (N_37505,N_37393,N_37331);
or U37506 (N_37506,N_37376,N_37379);
nor U37507 (N_37507,N_37498,N_37314);
xor U37508 (N_37508,N_37418,N_37334);
nor U37509 (N_37509,N_37277,N_37354);
or U37510 (N_37510,N_37265,N_37321);
nor U37511 (N_37511,N_37264,N_37263);
or U37512 (N_37512,N_37282,N_37385);
xor U37513 (N_37513,N_37359,N_37316);
or U37514 (N_37514,N_37473,N_37391);
and U37515 (N_37515,N_37464,N_37344);
nor U37516 (N_37516,N_37395,N_37477);
and U37517 (N_37517,N_37257,N_37343);
and U37518 (N_37518,N_37411,N_37375);
nor U37519 (N_37519,N_37357,N_37353);
nand U37520 (N_37520,N_37472,N_37400);
nor U37521 (N_37521,N_37338,N_37499);
xor U37522 (N_37522,N_37371,N_37300);
xnor U37523 (N_37523,N_37423,N_37479);
or U37524 (N_37524,N_37459,N_37483);
nand U37525 (N_37525,N_37284,N_37429);
nand U37526 (N_37526,N_37268,N_37267);
nor U37527 (N_37527,N_37481,N_37348);
and U37528 (N_37528,N_37485,N_37408);
xnor U37529 (N_37529,N_37413,N_37466);
and U37530 (N_37530,N_37435,N_37358);
and U37531 (N_37531,N_37296,N_37258);
nand U37532 (N_37532,N_37449,N_37490);
and U37533 (N_37533,N_37336,N_37323);
xnor U37534 (N_37534,N_37251,N_37330);
nor U37535 (N_37535,N_37401,N_37420);
and U37536 (N_37536,N_37351,N_37329);
and U37537 (N_37537,N_37261,N_37283);
nor U37538 (N_37538,N_37310,N_37339);
and U37539 (N_37539,N_37428,N_37365);
nor U37540 (N_37540,N_37362,N_37455);
and U37541 (N_37541,N_37325,N_37432);
or U37542 (N_37542,N_37469,N_37346);
nor U37543 (N_37543,N_37404,N_37315);
and U37544 (N_37544,N_37292,N_37288);
or U37545 (N_37545,N_37274,N_37445);
nand U37546 (N_37546,N_37317,N_37494);
or U37547 (N_37547,N_37443,N_37286);
nand U37548 (N_37548,N_37378,N_37252);
nor U37549 (N_37549,N_37409,N_37306);
nand U37550 (N_37550,N_37403,N_37397);
xor U37551 (N_37551,N_37335,N_37301);
nor U37552 (N_37552,N_37295,N_37437);
nor U37553 (N_37553,N_37298,N_37345);
xor U37554 (N_37554,N_37297,N_37434);
and U37555 (N_37555,N_37386,N_37438);
xnor U37556 (N_37556,N_37496,N_37281);
nand U37557 (N_37557,N_37394,N_37308);
xor U37558 (N_37558,N_37426,N_37484);
xnor U37559 (N_37559,N_37279,N_37349);
xor U37560 (N_37560,N_37419,N_37414);
xor U37561 (N_37561,N_37280,N_37340);
or U37562 (N_37562,N_37382,N_37327);
or U37563 (N_37563,N_37398,N_37273);
nand U37564 (N_37564,N_37337,N_37328);
nor U37565 (N_37565,N_37361,N_37250);
xnor U37566 (N_37566,N_37368,N_37369);
and U37567 (N_37567,N_37360,N_37387);
xor U37568 (N_37568,N_37461,N_37352);
xor U37569 (N_37569,N_37342,N_37441);
or U37570 (N_37570,N_37374,N_37470);
xnor U37571 (N_37571,N_37474,N_37383);
and U37572 (N_37572,N_37302,N_37276);
nor U37573 (N_37573,N_37407,N_37377);
nor U37574 (N_37574,N_37272,N_37253);
or U37575 (N_37575,N_37410,N_37424);
xor U37576 (N_37576,N_37256,N_37322);
nand U37577 (N_37577,N_37366,N_37255);
or U37578 (N_37578,N_37373,N_37491);
nor U37579 (N_37579,N_37467,N_37259);
xor U37580 (N_37580,N_37260,N_37486);
xor U37581 (N_37581,N_37431,N_37380);
and U37582 (N_37582,N_37451,N_37465);
xnor U37583 (N_37583,N_37311,N_37309);
nand U37584 (N_37584,N_37313,N_37275);
and U37585 (N_37585,N_37381,N_37433);
nor U37586 (N_37586,N_37287,N_37402);
nand U37587 (N_37587,N_37495,N_37271);
xor U37588 (N_37588,N_37350,N_37318);
nand U37589 (N_37589,N_37370,N_37436);
nor U37590 (N_37590,N_37452,N_37440);
xor U37591 (N_37591,N_37497,N_37460);
xor U37592 (N_37592,N_37269,N_37388);
nand U37593 (N_37593,N_37475,N_37290);
or U37594 (N_37594,N_37456,N_37305);
and U37595 (N_37595,N_37478,N_37307);
nand U37596 (N_37596,N_37262,N_37326);
or U37597 (N_37597,N_37448,N_37493);
xor U37598 (N_37598,N_37487,N_37303);
or U37599 (N_37599,N_37444,N_37364);
or U37600 (N_37600,N_37396,N_37285);
nand U37601 (N_37601,N_37324,N_37320);
nand U37602 (N_37602,N_37390,N_37488);
nor U37603 (N_37603,N_37492,N_37447);
nand U37604 (N_37604,N_37399,N_37304);
and U37605 (N_37605,N_37356,N_37372);
xor U37606 (N_37606,N_37389,N_37458);
nand U37607 (N_37607,N_37355,N_37427);
and U37608 (N_37608,N_37406,N_37416);
and U37609 (N_37609,N_37450,N_37439);
nor U37610 (N_37610,N_37333,N_37482);
and U37611 (N_37611,N_37270,N_37254);
xnor U37612 (N_37612,N_37405,N_37341);
nor U37613 (N_37613,N_37367,N_37347);
nand U37614 (N_37614,N_37291,N_37421);
or U37615 (N_37615,N_37415,N_37480);
and U37616 (N_37616,N_37294,N_37442);
or U37617 (N_37617,N_37319,N_37278);
nor U37618 (N_37618,N_37457,N_37289);
xor U37619 (N_37619,N_37312,N_37471);
nand U37620 (N_37620,N_37454,N_37468);
nand U37621 (N_37621,N_37425,N_37476);
nand U37622 (N_37622,N_37412,N_37266);
nand U37623 (N_37623,N_37453,N_37363);
xor U37624 (N_37624,N_37332,N_37462);
nor U37625 (N_37625,N_37392,N_37324);
nor U37626 (N_37626,N_37413,N_37394);
and U37627 (N_37627,N_37363,N_37349);
or U37628 (N_37628,N_37281,N_37336);
nor U37629 (N_37629,N_37388,N_37332);
nor U37630 (N_37630,N_37322,N_37270);
or U37631 (N_37631,N_37462,N_37302);
xnor U37632 (N_37632,N_37292,N_37297);
xor U37633 (N_37633,N_37472,N_37296);
nand U37634 (N_37634,N_37492,N_37397);
nor U37635 (N_37635,N_37259,N_37443);
or U37636 (N_37636,N_37414,N_37429);
and U37637 (N_37637,N_37440,N_37394);
or U37638 (N_37638,N_37325,N_37463);
or U37639 (N_37639,N_37437,N_37453);
xor U37640 (N_37640,N_37394,N_37388);
nand U37641 (N_37641,N_37460,N_37445);
xor U37642 (N_37642,N_37303,N_37379);
xor U37643 (N_37643,N_37445,N_37288);
and U37644 (N_37644,N_37411,N_37382);
or U37645 (N_37645,N_37370,N_37441);
xor U37646 (N_37646,N_37301,N_37482);
nand U37647 (N_37647,N_37449,N_37382);
and U37648 (N_37648,N_37361,N_37279);
xor U37649 (N_37649,N_37269,N_37453);
nor U37650 (N_37650,N_37461,N_37258);
or U37651 (N_37651,N_37387,N_37439);
or U37652 (N_37652,N_37353,N_37279);
or U37653 (N_37653,N_37333,N_37254);
nor U37654 (N_37654,N_37338,N_37480);
nand U37655 (N_37655,N_37328,N_37345);
and U37656 (N_37656,N_37361,N_37324);
xor U37657 (N_37657,N_37368,N_37473);
and U37658 (N_37658,N_37487,N_37416);
nor U37659 (N_37659,N_37336,N_37485);
nand U37660 (N_37660,N_37254,N_37454);
or U37661 (N_37661,N_37285,N_37468);
nand U37662 (N_37662,N_37258,N_37453);
nand U37663 (N_37663,N_37294,N_37298);
and U37664 (N_37664,N_37386,N_37494);
xor U37665 (N_37665,N_37467,N_37427);
nand U37666 (N_37666,N_37488,N_37405);
xnor U37667 (N_37667,N_37355,N_37409);
or U37668 (N_37668,N_37265,N_37492);
or U37669 (N_37669,N_37425,N_37363);
nor U37670 (N_37670,N_37438,N_37352);
and U37671 (N_37671,N_37304,N_37300);
nand U37672 (N_37672,N_37365,N_37279);
and U37673 (N_37673,N_37393,N_37383);
xnor U37674 (N_37674,N_37448,N_37300);
nor U37675 (N_37675,N_37324,N_37330);
nand U37676 (N_37676,N_37397,N_37300);
nand U37677 (N_37677,N_37295,N_37360);
and U37678 (N_37678,N_37431,N_37349);
and U37679 (N_37679,N_37469,N_37273);
and U37680 (N_37680,N_37433,N_37427);
and U37681 (N_37681,N_37372,N_37359);
or U37682 (N_37682,N_37263,N_37410);
or U37683 (N_37683,N_37325,N_37439);
nand U37684 (N_37684,N_37264,N_37288);
nor U37685 (N_37685,N_37346,N_37458);
and U37686 (N_37686,N_37372,N_37322);
and U37687 (N_37687,N_37254,N_37430);
xnor U37688 (N_37688,N_37345,N_37369);
or U37689 (N_37689,N_37395,N_37432);
and U37690 (N_37690,N_37440,N_37427);
nand U37691 (N_37691,N_37408,N_37357);
nand U37692 (N_37692,N_37309,N_37369);
nand U37693 (N_37693,N_37376,N_37485);
nand U37694 (N_37694,N_37259,N_37318);
and U37695 (N_37695,N_37288,N_37389);
or U37696 (N_37696,N_37378,N_37480);
nand U37697 (N_37697,N_37456,N_37272);
or U37698 (N_37698,N_37279,N_37482);
xor U37699 (N_37699,N_37483,N_37374);
nand U37700 (N_37700,N_37389,N_37319);
xor U37701 (N_37701,N_37284,N_37382);
xnor U37702 (N_37702,N_37374,N_37356);
and U37703 (N_37703,N_37430,N_37474);
and U37704 (N_37704,N_37335,N_37268);
nor U37705 (N_37705,N_37436,N_37470);
or U37706 (N_37706,N_37315,N_37260);
and U37707 (N_37707,N_37348,N_37288);
and U37708 (N_37708,N_37299,N_37260);
and U37709 (N_37709,N_37438,N_37469);
nand U37710 (N_37710,N_37398,N_37441);
xor U37711 (N_37711,N_37374,N_37282);
nand U37712 (N_37712,N_37379,N_37422);
nor U37713 (N_37713,N_37475,N_37461);
xnor U37714 (N_37714,N_37485,N_37494);
or U37715 (N_37715,N_37346,N_37439);
or U37716 (N_37716,N_37419,N_37435);
xnor U37717 (N_37717,N_37303,N_37461);
nor U37718 (N_37718,N_37266,N_37298);
nand U37719 (N_37719,N_37421,N_37316);
nand U37720 (N_37720,N_37489,N_37420);
or U37721 (N_37721,N_37413,N_37362);
and U37722 (N_37722,N_37433,N_37405);
xnor U37723 (N_37723,N_37357,N_37266);
or U37724 (N_37724,N_37464,N_37367);
and U37725 (N_37725,N_37277,N_37454);
xor U37726 (N_37726,N_37260,N_37337);
nand U37727 (N_37727,N_37465,N_37329);
xnor U37728 (N_37728,N_37275,N_37456);
or U37729 (N_37729,N_37422,N_37329);
nand U37730 (N_37730,N_37284,N_37428);
nor U37731 (N_37731,N_37335,N_37381);
xnor U37732 (N_37732,N_37369,N_37430);
nor U37733 (N_37733,N_37281,N_37335);
nor U37734 (N_37734,N_37409,N_37379);
nor U37735 (N_37735,N_37414,N_37497);
nand U37736 (N_37736,N_37396,N_37391);
and U37737 (N_37737,N_37376,N_37377);
nand U37738 (N_37738,N_37309,N_37427);
nand U37739 (N_37739,N_37313,N_37368);
nor U37740 (N_37740,N_37393,N_37379);
or U37741 (N_37741,N_37416,N_37339);
nand U37742 (N_37742,N_37459,N_37481);
nor U37743 (N_37743,N_37304,N_37452);
xnor U37744 (N_37744,N_37298,N_37332);
and U37745 (N_37745,N_37338,N_37265);
nor U37746 (N_37746,N_37496,N_37291);
or U37747 (N_37747,N_37320,N_37473);
and U37748 (N_37748,N_37319,N_37291);
and U37749 (N_37749,N_37268,N_37337);
xor U37750 (N_37750,N_37665,N_37699);
or U37751 (N_37751,N_37746,N_37747);
xor U37752 (N_37752,N_37614,N_37598);
nand U37753 (N_37753,N_37654,N_37647);
and U37754 (N_37754,N_37670,N_37696);
and U37755 (N_37755,N_37588,N_37677);
nor U37756 (N_37756,N_37657,N_37674);
nor U37757 (N_37757,N_37728,N_37623);
xor U37758 (N_37758,N_37527,N_37611);
xnor U37759 (N_37759,N_37649,N_37564);
and U37760 (N_37760,N_37544,N_37620);
and U37761 (N_37761,N_37703,N_37679);
xor U37762 (N_37762,N_37547,N_37740);
and U37763 (N_37763,N_37624,N_37700);
xnor U37764 (N_37764,N_37744,N_37538);
xor U37765 (N_37765,N_37736,N_37511);
xnor U37766 (N_37766,N_37621,N_37526);
xnor U37767 (N_37767,N_37570,N_37590);
nand U37768 (N_37768,N_37643,N_37635);
nand U37769 (N_37769,N_37726,N_37594);
nand U37770 (N_37770,N_37537,N_37519);
nand U37771 (N_37771,N_37622,N_37552);
or U37772 (N_37772,N_37539,N_37713);
nand U37773 (N_37773,N_37546,N_37615);
and U37774 (N_37774,N_37716,N_37613);
xnor U37775 (N_37775,N_37609,N_37507);
and U37776 (N_37776,N_37673,N_37708);
nor U37777 (N_37777,N_37516,N_37535);
xnor U37778 (N_37778,N_37645,N_37691);
and U37779 (N_37779,N_37510,N_37693);
nor U37780 (N_37780,N_37671,N_37541);
xor U37781 (N_37781,N_37604,N_37733);
and U37782 (N_37782,N_37596,N_37737);
nor U37783 (N_37783,N_37722,N_37509);
nand U37784 (N_37784,N_37707,N_37548);
nand U37785 (N_37785,N_37543,N_37506);
and U37786 (N_37786,N_37682,N_37639);
and U37787 (N_37787,N_37636,N_37618);
nand U37788 (N_37788,N_37721,N_37606);
xor U37789 (N_37789,N_37686,N_37522);
xnor U37790 (N_37790,N_37640,N_37698);
or U37791 (N_37791,N_37638,N_37560);
nand U37792 (N_37792,N_37616,N_37669);
xor U37793 (N_37793,N_37702,N_37508);
nand U37794 (N_37794,N_37581,N_37617);
nor U37795 (N_37795,N_37748,N_37578);
and U37796 (N_37796,N_37550,N_37629);
xor U37797 (N_37797,N_37556,N_37666);
xnor U37798 (N_37798,N_37569,N_37530);
nand U37799 (N_37799,N_37563,N_37658);
nor U37800 (N_37800,N_37675,N_37549);
xor U37801 (N_37801,N_37601,N_37749);
and U37802 (N_37802,N_37690,N_37553);
or U37803 (N_37803,N_37571,N_37630);
or U37804 (N_37804,N_37694,N_37582);
nor U37805 (N_37805,N_37641,N_37695);
nand U37806 (N_37806,N_37644,N_37566);
or U37807 (N_37807,N_37687,N_37719);
xor U37808 (N_37808,N_37559,N_37661);
nand U37809 (N_37809,N_37685,N_37576);
nand U37810 (N_37810,N_37642,N_37727);
or U37811 (N_37811,N_37592,N_37612);
xor U37812 (N_37812,N_37723,N_37524);
and U37813 (N_37813,N_37701,N_37709);
and U37814 (N_37814,N_37741,N_37579);
and U37815 (N_37815,N_37589,N_37565);
or U37816 (N_37816,N_37531,N_37520);
xor U37817 (N_37817,N_37575,N_37529);
and U37818 (N_37818,N_37706,N_37512);
and U37819 (N_37819,N_37729,N_37653);
xnor U37820 (N_37820,N_37634,N_37731);
nand U37821 (N_37821,N_37646,N_37659);
or U37822 (N_37822,N_37577,N_37584);
and U37823 (N_37823,N_37540,N_37562);
or U37824 (N_37824,N_37625,N_37710);
nand U37825 (N_37825,N_37632,N_37554);
or U37826 (N_37826,N_37678,N_37514);
nand U37827 (N_37827,N_37501,N_37610);
xor U37828 (N_37828,N_37568,N_37626);
nor U37829 (N_37829,N_37504,N_37715);
nand U37830 (N_37830,N_37650,N_37697);
xor U37831 (N_37831,N_37724,N_37689);
or U37832 (N_37832,N_37717,N_37718);
nor U37833 (N_37833,N_37743,N_37593);
nand U37834 (N_37834,N_37502,N_37664);
or U37835 (N_37835,N_37534,N_37681);
nand U37836 (N_37836,N_37655,N_37599);
xor U37837 (N_37837,N_37652,N_37608);
or U37838 (N_37838,N_37725,N_37521);
nor U37839 (N_37839,N_37631,N_37574);
or U37840 (N_37840,N_37518,N_37734);
and U37841 (N_37841,N_37633,N_37533);
or U37842 (N_37842,N_37500,N_37503);
nand U37843 (N_37843,N_37745,N_37603);
nor U37844 (N_37844,N_37667,N_37648);
or U37845 (N_37845,N_37513,N_37662);
nand U37846 (N_37846,N_37739,N_37551);
nor U37847 (N_37847,N_37567,N_37711);
nor U37848 (N_37848,N_37672,N_37525);
and U37849 (N_37849,N_37732,N_37668);
nor U37850 (N_37850,N_37676,N_37742);
nand U37851 (N_37851,N_37712,N_37558);
xor U37852 (N_37852,N_37714,N_37627);
or U37853 (N_37853,N_37705,N_37607);
nor U37854 (N_37854,N_37542,N_37557);
nand U37855 (N_37855,N_37684,N_37688);
and U37856 (N_37856,N_37683,N_37580);
nor U37857 (N_37857,N_37663,N_37704);
xor U37858 (N_37858,N_37720,N_37532);
xor U37859 (N_37859,N_37515,N_37517);
nand U37860 (N_37860,N_37730,N_37572);
nand U37861 (N_37861,N_37597,N_37619);
xor U37862 (N_37862,N_37735,N_37585);
and U37863 (N_37863,N_37536,N_37505);
and U37864 (N_37864,N_37680,N_37656);
or U37865 (N_37865,N_37605,N_37651);
nor U37866 (N_37866,N_37573,N_37561);
nor U37867 (N_37867,N_37738,N_37583);
nor U37868 (N_37868,N_37545,N_37591);
xor U37869 (N_37869,N_37602,N_37555);
xor U37870 (N_37870,N_37692,N_37600);
xor U37871 (N_37871,N_37660,N_37528);
xnor U37872 (N_37872,N_37637,N_37587);
and U37873 (N_37873,N_37523,N_37595);
xnor U37874 (N_37874,N_37586,N_37628);
or U37875 (N_37875,N_37669,N_37619);
nor U37876 (N_37876,N_37508,N_37696);
nand U37877 (N_37877,N_37592,N_37609);
xnor U37878 (N_37878,N_37690,N_37669);
xnor U37879 (N_37879,N_37649,N_37724);
and U37880 (N_37880,N_37687,N_37501);
or U37881 (N_37881,N_37700,N_37717);
or U37882 (N_37882,N_37582,N_37638);
xnor U37883 (N_37883,N_37652,N_37567);
nor U37884 (N_37884,N_37690,N_37582);
xnor U37885 (N_37885,N_37707,N_37684);
or U37886 (N_37886,N_37739,N_37713);
and U37887 (N_37887,N_37685,N_37589);
and U37888 (N_37888,N_37718,N_37581);
nor U37889 (N_37889,N_37550,N_37742);
nand U37890 (N_37890,N_37737,N_37684);
nand U37891 (N_37891,N_37517,N_37511);
nand U37892 (N_37892,N_37724,N_37721);
xnor U37893 (N_37893,N_37607,N_37677);
nand U37894 (N_37894,N_37589,N_37716);
nand U37895 (N_37895,N_37555,N_37739);
and U37896 (N_37896,N_37536,N_37558);
nand U37897 (N_37897,N_37522,N_37549);
or U37898 (N_37898,N_37503,N_37667);
xor U37899 (N_37899,N_37735,N_37667);
nand U37900 (N_37900,N_37511,N_37503);
nor U37901 (N_37901,N_37747,N_37608);
nor U37902 (N_37902,N_37549,N_37570);
nand U37903 (N_37903,N_37613,N_37701);
nor U37904 (N_37904,N_37538,N_37734);
and U37905 (N_37905,N_37691,N_37621);
nor U37906 (N_37906,N_37539,N_37564);
or U37907 (N_37907,N_37576,N_37730);
nand U37908 (N_37908,N_37531,N_37749);
and U37909 (N_37909,N_37723,N_37717);
xor U37910 (N_37910,N_37516,N_37684);
xnor U37911 (N_37911,N_37502,N_37661);
or U37912 (N_37912,N_37670,N_37525);
nand U37913 (N_37913,N_37647,N_37644);
or U37914 (N_37914,N_37559,N_37543);
or U37915 (N_37915,N_37555,N_37623);
or U37916 (N_37916,N_37508,N_37530);
and U37917 (N_37917,N_37562,N_37653);
and U37918 (N_37918,N_37709,N_37629);
and U37919 (N_37919,N_37598,N_37557);
or U37920 (N_37920,N_37643,N_37680);
nor U37921 (N_37921,N_37605,N_37706);
nand U37922 (N_37922,N_37718,N_37713);
xor U37923 (N_37923,N_37622,N_37687);
and U37924 (N_37924,N_37677,N_37739);
nand U37925 (N_37925,N_37647,N_37541);
nor U37926 (N_37926,N_37744,N_37519);
nand U37927 (N_37927,N_37710,N_37661);
or U37928 (N_37928,N_37745,N_37570);
or U37929 (N_37929,N_37632,N_37676);
nor U37930 (N_37930,N_37682,N_37697);
or U37931 (N_37931,N_37608,N_37500);
or U37932 (N_37932,N_37521,N_37507);
and U37933 (N_37933,N_37725,N_37721);
nand U37934 (N_37934,N_37599,N_37684);
nand U37935 (N_37935,N_37746,N_37697);
nand U37936 (N_37936,N_37542,N_37646);
nor U37937 (N_37937,N_37697,N_37701);
nand U37938 (N_37938,N_37685,N_37620);
and U37939 (N_37939,N_37689,N_37723);
nor U37940 (N_37940,N_37556,N_37603);
and U37941 (N_37941,N_37653,N_37553);
nor U37942 (N_37942,N_37579,N_37677);
nand U37943 (N_37943,N_37678,N_37723);
nand U37944 (N_37944,N_37739,N_37710);
nand U37945 (N_37945,N_37528,N_37560);
nand U37946 (N_37946,N_37702,N_37674);
xnor U37947 (N_37947,N_37593,N_37673);
nor U37948 (N_37948,N_37683,N_37748);
xnor U37949 (N_37949,N_37522,N_37654);
or U37950 (N_37950,N_37558,N_37656);
nor U37951 (N_37951,N_37558,N_37653);
xnor U37952 (N_37952,N_37727,N_37690);
nor U37953 (N_37953,N_37509,N_37533);
nand U37954 (N_37954,N_37565,N_37539);
and U37955 (N_37955,N_37580,N_37611);
xor U37956 (N_37956,N_37576,N_37640);
and U37957 (N_37957,N_37642,N_37695);
and U37958 (N_37958,N_37593,N_37590);
nand U37959 (N_37959,N_37568,N_37677);
or U37960 (N_37960,N_37659,N_37530);
and U37961 (N_37961,N_37695,N_37535);
or U37962 (N_37962,N_37573,N_37607);
or U37963 (N_37963,N_37685,N_37548);
nor U37964 (N_37964,N_37620,N_37622);
nand U37965 (N_37965,N_37588,N_37583);
and U37966 (N_37966,N_37564,N_37549);
xor U37967 (N_37967,N_37532,N_37536);
and U37968 (N_37968,N_37542,N_37551);
xnor U37969 (N_37969,N_37628,N_37517);
nor U37970 (N_37970,N_37566,N_37564);
and U37971 (N_37971,N_37630,N_37679);
nor U37972 (N_37972,N_37619,N_37565);
nor U37973 (N_37973,N_37550,N_37612);
and U37974 (N_37974,N_37720,N_37645);
or U37975 (N_37975,N_37714,N_37523);
nand U37976 (N_37976,N_37729,N_37500);
and U37977 (N_37977,N_37721,N_37716);
or U37978 (N_37978,N_37624,N_37579);
nand U37979 (N_37979,N_37659,N_37742);
or U37980 (N_37980,N_37610,N_37592);
xor U37981 (N_37981,N_37581,N_37558);
xor U37982 (N_37982,N_37534,N_37710);
nor U37983 (N_37983,N_37740,N_37597);
and U37984 (N_37984,N_37649,N_37692);
and U37985 (N_37985,N_37647,N_37530);
nand U37986 (N_37986,N_37541,N_37500);
and U37987 (N_37987,N_37566,N_37513);
nor U37988 (N_37988,N_37714,N_37660);
xor U37989 (N_37989,N_37524,N_37734);
and U37990 (N_37990,N_37600,N_37515);
nor U37991 (N_37991,N_37711,N_37671);
nor U37992 (N_37992,N_37576,N_37699);
and U37993 (N_37993,N_37704,N_37668);
nor U37994 (N_37994,N_37539,N_37679);
nand U37995 (N_37995,N_37638,N_37737);
or U37996 (N_37996,N_37608,N_37551);
and U37997 (N_37997,N_37572,N_37589);
or U37998 (N_37998,N_37587,N_37636);
nand U37999 (N_37999,N_37554,N_37586);
and U38000 (N_38000,N_37824,N_37968);
and U38001 (N_38001,N_37954,N_37854);
or U38002 (N_38002,N_37802,N_37997);
or U38003 (N_38003,N_37805,N_37832);
and U38004 (N_38004,N_37781,N_37962);
and U38005 (N_38005,N_37931,N_37933);
and U38006 (N_38006,N_37856,N_37953);
xor U38007 (N_38007,N_37794,N_37889);
xnor U38008 (N_38008,N_37766,N_37967);
xnor U38009 (N_38009,N_37771,N_37846);
or U38010 (N_38010,N_37974,N_37810);
and U38011 (N_38011,N_37793,N_37911);
or U38012 (N_38012,N_37892,N_37993);
xor U38013 (N_38013,N_37948,N_37878);
nand U38014 (N_38014,N_37891,N_37995);
xor U38015 (N_38015,N_37830,N_37982);
nor U38016 (N_38016,N_37775,N_37866);
or U38017 (N_38017,N_37849,N_37867);
and U38018 (N_38018,N_37760,N_37937);
or U38019 (N_38019,N_37976,N_37940);
or U38020 (N_38020,N_37780,N_37880);
nor U38021 (N_38021,N_37768,N_37938);
or U38022 (N_38022,N_37779,N_37978);
xnor U38023 (N_38023,N_37828,N_37947);
xor U38024 (N_38024,N_37876,N_37848);
nor U38025 (N_38025,N_37888,N_37847);
nor U38026 (N_38026,N_37773,N_37902);
and U38027 (N_38027,N_37970,N_37965);
nor U38028 (N_38028,N_37899,N_37914);
nor U38029 (N_38029,N_37986,N_37930);
or U38030 (N_38030,N_37945,N_37894);
and U38031 (N_38031,N_37851,N_37922);
and U38032 (N_38032,N_37842,N_37898);
nand U38033 (N_38033,N_37753,N_37835);
and U38034 (N_38034,N_37815,N_37798);
nor U38035 (N_38035,N_37977,N_37836);
or U38036 (N_38036,N_37797,N_37785);
nand U38037 (N_38037,N_37936,N_37778);
nand U38038 (N_38038,N_37865,N_37907);
and U38039 (N_38039,N_37784,N_37825);
xor U38040 (N_38040,N_37811,N_37819);
xnor U38041 (N_38041,N_37783,N_37958);
and U38042 (N_38042,N_37883,N_37770);
or U38043 (N_38043,N_37998,N_37951);
or U38044 (N_38044,N_37840,N_37864);
nor U38045 (N_38045,N_37893,N_37787);
nand U38046 (N_38046,N_37764,N_37909);
and U38047 (N_38047,N_37837,N_37971);
and U38048 (N_38048,N_37926,N_37814);
and U38049 (N_38049,N_37859,N_37843);
xor U38050 (N_38050,N_37791,N_37756);
nor U38051 (N_38051,N_37942,N_37944);
xnor U38052 (N_38052,N_37872,N_37941);
nor U38053 (N_38053,N_37799,N_37786);
or U38054 (N_38054,N_37973,N_37757);
nand U38055 (N_38055,N_37987,N_37855);
and U38056 (N_38056,N_37873,N_37887);
xor U38057 (N_38057,N_37919,N_37917);
xnor U38058 (N_38058,N_37762,N_37890);
and U38059 (N_38059,N_37964,N_37761);
nor U38060 (N_38060,N_37896,N_37833);
nand U38061 (N_38061,N_37776,N_37874);
and U38062 (N_38062,N_37925,N_37981);
nand U38063 (N_38063,N_37861,N_37790);
and U38064 (N_38064,N_37817,N_37969);
or U38065 (N_38065,N_37881,N_37871);
nor U38066 (N_38066,N_37939,N_37895);
nand U38067 (N_38067,N_37765,N_37857);
nand U38068 (N_38068,N_37816,N_37863);
nor U38069 (N_38069,N_37988,N_37908);
nand U38070 (N_38070,N_37901,N_37803);
and U38071 (N_38071,N_37996,N_37956);
and U38072 (N_38072,N_37834,N_37915);
or U38073 (N_38073,N_37763,N_37991);
or U38074 (N_38074,N_37950,N_37852);
and U38075 (N_38075,N_37959,N_37979);
nor U38076 (N_38076,N_37961,N_37906);
or U38077 (N_38077,N_37809,N_37935);
nand U38078 (N_38078,N_37966,N_37860);
xnor U38079 (N_38079,N_37807,N_37980);
or U38080 (N_38080,N_37792,N_37868);
nor U38081 (N_38081,N_37806,N_37813);
nor U38082 (N_38082,N_37796,N_37989);
or U38083 (N_38083,N_37882,N_37920);
nor U38084 (N_38084,N_37788,N_37812);
xor U38085 (N_38085,N_37800,N_37820);
nand U38086 (N_38086,N_37990,N_37905);
nand U38087 (N_38087,N_37877,N_37910);
and U38088 (N_38088,N_37831,N_37759);
nor U38089 (N_38089,N_37772,N_37904);
and U38090 (N_38090,N_37829,N_37752);
and U38091 (N_38091,N_37769,N_37912);
and U38092 (N_38092,N_37818,N_37822);
and U38093 (N_38093,N_37853,N_37879);
xnor U38094 (N_38094,N_37924,N_37777);
and U38095 (N_38095,N_37900,N_37839);
or U38096 (N_38096,N_37929,N_37767);
and U38097 (N_38097,N_37827,N_37758);
and U38098 (N_38098,N_37949,N_37841);
nor U38099 (N_38099,N_37844,N_37903);
nand U38100 (N_38100,N_37913,N_37774);
nand U38101 (N_38101,N_37750,N_37808);
and U38102 (N_38102,N_37838,N_37823);
nor U38103 (N_38103,N_37886,N_37862);
or U38104 (N_38104,N_37985,N_37934);
or U38105 (N_38105,N_37923,N_37960);
nor U38106 (N_38106,N_37983,N_37845);
xnor U38107 (N_38107,N_37943,N_37804);
nand U38108 (N_38108,N_37932,N_37795);
xor U38109 (N_38109,N_37789,N_37850);
nand U38110 (N_38110,N_37801,N_37972);
xnor U38111 (N_38111,N_37918,N_37751);
nor U38112 (N_38112,N_37946,N_37921);
nor U38113 (N_38113,N_37826,N_37885);
nor U38114 (N_38114,N_37957,N_37884);
xnor U38115 (N_38115,N_37858,N_37955);
or U38116 (N_38116,N_37992,N_37963);
and U38117 (N_38117,N_37754,N_37999);
or U38118 (N_38118,N_37821,N_37782);
or U38119 (N_38119,N_37984,N_37875);
and U38120 (N_38120,N_37952,N_37927);
and U38121 (N_38121,N_37870,N_37916);
and U38122 (N_38122,N_37928,N_37869);
or U38123 (N_38123,N_37897,N_37755);
nand U38124 (N_38124,N_37975,N_37994);
nor U38125 (N_38125,N_37923,N_37928);
nor U38126 (N_38126,N_37770,N_37840);
nor U38127 (N_38127,N_37808,N_37926);
nand U38128 (N_38128,N_37946,N_37913);
and U38129 (N_38129,N_37921,N_37873);
and U38130 (N_38130,N_37774,N_37968);
nor U38131 (N_38131,N_37759,N_37779);
xnor U38132 (N_38132,N_37985,N_37892);
nor U38133 (N_38133,N_37921,N_37977);
or U38134 (N_38134,N_37991,N_37950);
or U38135 (N_38135,N_37927,N_37886);
or U38136 (N_38136,N_37881,N_37858);
or U38137 (N_38137,N_37839,N_37927);
nand U38138 (N_38138,N_37972,N_37793);
nand U38139 (N_38139,N_37806,N_37829);
nor U38140 (N_38140,N_37774,N_37953);
xor U38141 (N_38141,N_37868,N_37833);
or U38142 (N_38142,N_37820,N_37933);
xor U38143 (N_38143,N_37920,N_37898);
and U38144 (N_38144,N_37874,N_37953);
xnor U38145 (N_38145,N_37911,N_37874);
nand U38146 (N_38146,N_37756,N_37814);
and U38147 (N_38147,N_37933,N_37828);
and U38148 (N_38148,N_37968,N_37881);
nor U38149 (N_38149,N_37855,N_37793);
nor U38150 (N_38150,N_37750,N_37766);
nand U38151 (N_38151,N_37991,N_37755);
xnor U38152 (N_38152,N_37940,N_37993);
nand U38153 (N_38153,N_37979,N_37857);
and U38154 (N_38154,N_37858,N_37869);
nand U38155 (N_38155,N_37857,N_37858);
or U38156 (N_38156,N_37984,N_37965);
or U38157 (N_38157,N_37941,N_37798);
xnor U38158 (N_38158,N_37962,N_37915);
and U38159 (N_38159,N_37857,N_37833);
xnor U38160 (N_38160,N_37920,N_37949);
nand U38161 (N_38161,N_37979,N_37773);
or U38162 (N_38162,N_37754,N_37925);
or U38163 (N_38163,N_37855,N_37992);
nand U38164 (N_38164,N_37850,N_37898);
and U38165 (N_38165,N_37930,N_37839);
and U38166 (N_38166,N_37770,N_37908);
nand U38167 (N_38167,N_37803,N_37859);
and U38168 (N_38168,N_37959,N_37956);
nand U38169 (N_38169,N_37804,N_37879);
xor U38170 (N_38170,N_37981,N_37995);
nand U38171 (N_38171,N_37751,N_37941);
nor U38172 (N_38172,N_37968,N_37823);
or U38173 (N_38173,N_37782,N_37989);
or U38174 (N_38174,N_37993,N_37937);
or U38175 (N_38175,N_37962,N_37872);
nor U38176 (N_38176,N_37994,N_37864);
and U38177 (N_38177,N_37803,N_37969);
and U38178 (N_38178,N_37815,N_37769);
nand U38179 (N_38179,N_37870,N_37758);
nor U38180 (N_38180,N_37864,N_37762);
or U38181 (N_38181,N_37853,N_37787);
and U38182 (N_38182,N_37929,N_37813);
xor U38183 (N_38183,N_37777,N_37862);
nand U38184 (N_38184,N_37962,N_37857);
and U38185 (N_38185,N_37999,N_37793);
or U38186 (N_38186,N_37908,N_37921);
nor U38187 (N_38187,N_37898,N_37976);
and U38188 (N_38188,N_37859,N_37990);
nor U38189 (N_38189,N_37982,N_37990);
or U38190 (N_38190,N_37893,N_37806);
or U38191 (N_38191,N_37927,N_37815);
nand U38192 (N_38192,N_37782,N_37768);
nor U38193 (N_38193,N_37800,N_37850);
xor U38194 (N_38194,N_37755,N_37875);
nand U38195 (N_38195,N_37878,N_37850);
or U38196 (N_38196,N_37889,N_37995);
or U38197 (N_38197,N_37955,N_37965);
nor U38198 (N_38198,N_37958,N_37984);
nand U38199 (N_38199,N_37994,N_37836);
nor U38200 (N_38200,N_37786,N_37972);
or U38201 (N_38201,N_37801,N_37786);
xor U38202 (N_38202,N_37974,N_37762);
xor U38203 (N_38203,N_37847,N_37766);
or U38204 (N_38204,N_37783,N_37878);
nor U38205 (N_38205,N_37785,N_37752);
and U38206 (N_38206,N_37937,N_37824);
nor U38207 (N_38207,N_37844,N_37938);
or U38208 (N_38208,N_37915,N_37879);
and U38209 (N_38209,N_37948,N_37962);
and U38210 (N_38210,N_37867,N_37843);
xnor U38211 (N_38211,N_37804,N_37930);
nor U38212 (N_38212,N_37870,N_37850);
and U38213 (N_38213,N_37932,N_37783);
and U38214 (N_38214,N_37834,N_37800);
and U38215 (N_38215,N_37876,N_37777);
nor U38216 (N_38216,N_37825,N_37882);
or U38217 (N_38217,N_37770,N_37828);
and U38218 (N_38218,N_37992,N_37902);
or U38219 (N_38219,N_37799,N_37933);
or U38220 (N_38220,N_37949,N_37779);
nor U38221 (N_38221,N_37875,N_37819);
nand U38222 (N_38222,N_37795,N_37950);
nor U38223 (N_38223,N_37929,N_37990);
and U38224 (N_38224,N_37934,N_37852);
nand U38225 (N_38225,N_37863,N_37958);
nor U38226 (N_38226,N_37824,N_37799);
xor U38227 (N_38227,N_37854,N_37862);
or U38228 (N_38228,N_37784,N_37996);
nand U38229 (N_38229,N_37942,N_37922);
and U38230 (N_38230,N_37787,N_37931);
or U38231 (N_38231,N_37874,N_37976);
and U38232 (N_38232,N_37818,N_37870);
and U38233 (N_38233,N_37909,N_37816);
nor U38234 (N_38234,N_37865,N_37766);
xnor U38235 (N_38235,N_37963,N_37904);
and U38236 (N_38236,N_37990,N_37956);
nand U38237 (N_38237,N_37817,N_37857);
nand U38238 (N_38238,N_37857,N_37905);
xor U38239 (N_38239,N_37900,N_37811);
nor U38240 (N_38240,N_37864,N_37775);
nor U38241 (N_38241,N_37931,N_37908);
and U38242 (N_38242,N_37993,N_37958);
and U38243 (N_38243,N_37988,N_37811);
xnor U38244 (N_38244,N_37904,N_37908);
nand U38245 (N_38245,N_37819,N_37964);
xor U38246 (N_38246,N_37871,N_37805);
nand U38247 (N_38247,N_37993,N_37931);
nand U38248 (N_38248,N_37772,N_37879);
nor U38249 (N_38249,N_37911,N_37903);
nand U38250 (N_38250,N_38148,N_38197);
or U38251 (N_38251,N_38119,N_38139);
xor U38252 (N_38252,N_38134,N_38063);
nor U38253 (N_38253,N_38121,N_38126);
or U38254 (N_38254,N_38072,N_38048);
and U38255 (N_38255,N_38242,N_38075);
nor U38256 (N_38256,N_38183,N_38137);
nor U38257 (N_38257,N_38237,N_38098);
xor U38258 (N_38258,N_38171,N_38232);
nand U38259 (N_38259,N_38004,N_38114);
and U38260 (N_38260,N_38026,N_38194);
nor U38261 (N_38261,N_38052,N_38185);
nor U38262 (N_38262,N_38084,N_38046);
nand U38263 (N_38263,N_38078,N_38245);
xnor U38264 (N_38264,N_38211,N_38175);
nand U38265 (N_38265,N_38039,N_38249);
or U38266 (N_38266,N_38047,N_38125);
or U38267 (N_38267,N_38091,N_38213);
nor U38268 (N_38268,N_38243,N_38229);
nand U38269 (N_38269,N_38058,N_38124);
or U38270 (N_38270,N_38116,N_38246);
or U38271 (N_38271,N_38220,N_38135);
xor U38272 (N_38272,N_38132,N_38112);
or U38273 (N_38273,N_38085,N_38234);
xnor U38274 (N_38274,N_38081,N_38167);
or U38275 (N_38275,N_38044,N_38079);
or U38276 (N_38276,N_38147,N_38195);
nor U38277 (N_38277,N_38031,N_38153);
nor U38278 (N_38278,N_38199,N_38154);
and U38279 (N_38279,N_38160,N_38221);
xor U38280 (N_38280,N_38248,N_38188);
nand U38281 (N_38281,N_38163,N_38041);
xor U38282 (N_38282,N_38042,N_38035);
nand U38283 (N_38283,N_38028,N_38010);
nor U38284 (N_38284,N_38017,N_38182);
xnor U38285 (N_38285,N_38025,N_38051);
and U38286 (N_38286,N_38021,N_38166);
and U38287 (N_38287,N_38179,N_38128);
and U38288 (N_38288,N_38203,N_38009);
nand U38289 (N_38289,N_38108,N_38105);
or U38290 (N_38290,N_38155,N_38113);
nor U38291 (N_38291,N_38140,N_38193);
nand U38292 (N_38292,N_38145,N_38239);
nor U38293 (N_38293,N_38130,N_38002);
nor U38294 (N_38294,N_38169,N_38205);
nor U38295 (N_38295,N_38082,N_38056);
nand U38296 (N_38296,N_38136,N_38003);
nor U38297 (N_38297,N_38032,N_38177);
nor U38298 (N_38298,N_38170,N_38102);
and U38299 (N_38299,N_38208,N_38138);
nand U38300 (N_38300,N_38146,N_38071);
nand U38301 (N_38301,N_38012,N_38172);
or U38302 (N_38302,N_38219,N_38055);
nor U38303 (N_38303,N_38173,N_38149);
nor U38304 (N_38304,N_38038,N_38057);
nor U38305 (N_38305,N_38068,N_38049);
nor U38306 (N_38306,N_38162,N_38103);
xor U38307 (N_38307,N_38202,N_38088);
and U38308 (N_38308,N_38150,N_38164);
or U38309 (N_38309,N_38217,N_38216);
and U38310 (N_38310,N_38020,N_38090);
and U38311 (N_38311,N_38067,N_38120);
or U38312 (N_38312,N_38061,N_38151);
nand U38313 (N_38313,N_38196,N_38206);
or U38314 (N_38314,N_38238,N_38142);
and U38315 (N_38315,N_38062,N_38212);
nor U38316 (N_38316,N_38040,N_38089);
or U38317 (N_38317,N_38107,N_38198);
xor U38318 (N_38318,N_38027,N_38083);
or U38319 (N_38319,N_38099,N_38161);
nor U38320 (N_38320,N_38096,N_38227);
xor U38321 (N_38321,N_38122,N_38241);
nor U38322 (N_38322,N_38200,N_38118);
nand U38323 (N_38323,N_38129,N_38015);
nand U38324 (N_38324,N_38030,N_38192);
xnor U38325 (N_38325,N_38156,N_38022);
nand U38326 (N_38326,N_38152,N_38157);
nand U38327 (N_38327,N_38024,N_38000);
or U38328 (N_38328,N_38133,N_38244);
nor U38329 (N_38329,N_38008,N_38005);
xor U38330 (N_38330,N_38123,N_38180);
nor U38331 (N_38331,N_38168,N_38190);
and U38332 (N_38332,N_38235,N_38143);
nor U38333 (N_38333,N_38228,N_38247);
nand U38334 (N_38334,N_38225,N_38037);
xnor U38335 (N_38335,N_38034,N_38100);
nor U38336 (N_38336,N_38109,N_38097);
and U38337 (N_38337,N_38076,N_38236);
or U38338 (N_38338,N_38191,N_38018);
or U38339 (N_38339,N_38210,N_38001);
and U38340 (N_38340,N_38043,N_38053);
nand U38341 (N_38341,N_38158,N_38033);
xnor U38342 (N_38342,N_38060,N_38178);
nor U38343 (N_38343,N_38117,N_38189);
nor U38344 (N_38344,N_38054,N_38074);
and U38345 (N_38345,N_38087,N_38016);
xor U38346 (N_38346,N_38110,N_38080);
nor U38347 (N_38347,N_38230,N_38104);
xnor U38348 (N_38348,N_38214,N_38070);
and U38349 (N_38349,N_38240,N_38013);
xor U38350 (N_38350,N_38141,N_38111);
and U38351 (N_38351,N_38218,N_38207);
or U38352 (N_38352,N_38184,N_38014);
or U38353 (N_38353,N_38069,N_38181);
and U38354 (N_38354,N_38019,N_38159);
and U38355 (N_38355,N_38036,N_38215);
or U38356 (N_38356,N_38209,N_38201);
and U38357 (N_38357,N_38059,N_38144);
nand U38358 (N_38358,N_38092,N_38073);
nand U38359 (N_38359,N_38065,N_38115);
nor U38360 (N_38360,N_38064,N_38224);
and U38361 (N_38361,N_38231,N_38187);
nor U38362 (N_38362,N_38127,N_38077);
nor U38363 (N_38363,N_38101,N_38086);
nand U38364 (N_38364,N_38106,N_38094);
xor U38365 (N_38365,N_38045,N_38226);
nor U38366 (N_38366,N_38093,N_38095);
nand U38367 (N_38367,N_38165,N_38131);
or U38368 (N_38368,N_38233,N_38222);
nand U38369 (N_38369,N_38204,N_38066);
or U38370 (N_38370,N_38006,N_38029);
xor U38371 (N_38371,N_38186,N_38176);
and U38372 (N_38372,N_38007,N_38223);
xor U38373 (N_38373,N_38174,N_38011);
nor U38374 (N_38374,N_38050,N_38023);
and U38375 (N_38375,N_38135,N_38152);
and U38376 (N_38376,N_38215,N_38085);
and U38377 (N_38377,N_38214,N_38185);
nand U38378 (N_38378,N_38245,N_38075);
and U38379 (N_38379,N_38179,N_38235);
nand U38380 (N_38380,N_38024,N_38204);
nand U38381 (N_38381,N_38126,N_38122);
nor U38382 (N_38382,N_38230,N_38082);
nor U38383 (N_38383,N_38009,N_38198);
xnor U38384 (N_38384,N_38158,N_38191);
and U38385 (N_38385,N_38097,N_38009);
xor U38386 (N_38386,N_38052,N_38234);
nor U38387 (N_38387,N_38168,N_38136);
and U38388 (N_38388,N_38087,N_38006);
or U38389 (N_38389,N_38119,N_38039);
nand U38390 (N_38390,N_38174,N_38049);
nand U38391 (N_38391,N_38078,N_38123);
and U38392 (N_38392,N_38092,N_38080);
and U38393 (N_38393,N_38121,N_38244);
xor U38394 (N_38394,N_38142,N_38247);
nor U38395 (N_38395,N_38074,N_38097);
and U38396 (N_38396,N_38178,N_38157);
and U38397 (N_38397,N_38106,N_38122);
nand U38398 (N_38398,N_38189,N_38044);
nor U38399 (N_38399,N_38018,N_38228);
or U38400 (N_38400,N_38015,N_38092);
nor U38401 (N_38401,N_38005,N_38184);
and U38402 (N_38402,N_38167,N_38073);
nand U38403 (N_38403,N_38126,N_38040);
nand U38404 (N_38404,N_38083,N_38127);
nor U38405 (N_38405,N_38054,N_38040);
and U38406 (N_38406,N_38088,N_38232);
and U38407 (N_38407,N_38133,N_38027);
and U38408 (N_38408,N_38165,N_38112);
nand U38409 (N_38409,N_38136,N_38247);
xor U38410 (N_38410,N_38143,N_38231);
or U38411 (N_38411,N_38140,N_38206);
or U38412 (N_38412,N_38201,N_38038);
nor U38413 (N_38413,N_38212,N_38153);
xor U38414 (N_38414,N_38121,N_38115);
nor U38415 (N_38415,N_38023,N_38055);
nor U38416 (N_38416,N_38082,N_38115);
nor U38417 (N_38417,N_38103,N_38056);
and U38418 (N_38418,N_38215,N_38244);
xor U38419 (N_38419,N_38071,N_38031);
nand U38420 (N_38420,N_38096,N_38071);
and U38421 (N_38421,N_38044,N_38142);
xor U38422 (N_38422,N_38186,N_38010);
or U38423 (N_38423,N_38119,N_38059);
xor U38424 (N_38424,N_38116,N_38174);
nor U38425 (N_38425,N_38154,N_38059);
or U38426 (N_38426,N_38002,N_38171);
xor U38427 (N_38427,N_38221,N_38113);
nor U38428 (N_38428,N_38003,N_38022);
nor U38429 (N_38429,N_38249,N_38092);
nor U38430 (N_38430,N_38115,N_38027);
nor U38431 (N_38431,N_38143,N_38157);
and U38432 (N_38432,N_38195,N_38162);
or U38433 (N_38433,N_38239,N_38213);
and U38434 (N_38434,N_38001,N_38096);
nor U38435 (N_38435,N_38249,N_38200);
and U38436 (N_38436,N_38053,N_38026);
xor U38437 (N_38437,N_38248,N_38125);
nand U38438 (N_38438,N_38091,N_38172);
or U38439 (N_38439,N_38135,N_38081);
or U38440 (N_38440,N_38185,N_38042);
or U38441 (N_38441,N_38100,N_38157);
nor U38442 (N_38442,N_38219,N_38025);
or U38443 (N_38443,N_38187,N_38197);
or U38444 (N_38444,N_38080,N_38182);
xnor U38445 (N_38445,N_38017,N_38207);
nand U38446 (N_38446,N_38129,N_38000);
and U38447 (N_38447,N_38140,N_38065);
and U38448 (N_38448,N_38172,N_38063);
and U38449 (N_38449,N_38037,N_38035);
xnor U38450 (N_38450,N_38075,N_38142);
nand U38451 (N_38451,N_38116,N_38015);
or U38452 (N_38452,N_38084,N_38226);
nor U38453 (N_38453,N_38182,N_38178);
nand U38454 (N_38454,N_38059,N_38026);
xor U38455 (N_38455,N_38090,N_38222);
nand U38456 (N_38456,N_38086,N_38115);
xor U38457 (N_38457,N_38108,N_38003);
xor U38458 (N_38458,N_38225,N_38007);
nand U38459 (N_38459,N_38057,N_38055);
xor U38460 (N_38460,N_38101,N_38162);
xnor U38461 (N_38461,N_38236,N_38103);
or U38462 (N_38462,N_38010,N_38079);
or U38463 (N_38463,N_38031,N_38129);
nand U38464 (N_38464,N_38044,N_38001);
and U38465 (N_38465,N_38061,N_38072);
and U38466 (N_38466,N_38241,N_38203);
xnor U38467 (N_38467,N_38070,N_38012);
and U38468 (N_38468,N_38130,N_38178);
nor U38469 (N_38469,N_38149,N_38247);
and U38470 (N_38470,N_38084,N_38047);
xnor U38471 (N_38471,N_38203,N_38081);
and U38472 (N_38472,N_38005,N_38168);
or U38473 (N_38473,N_38228,N_38237);
or U38474 (N_38474,N_38231,N_38052);
and U38475 (N_38475,N_38164,N_38109);
and U38476 (N_38476,N_38024,N_38049);
and U38477 (N_38477,N_38004,N_38067);
xor U38478 (N_38478,N_38044,N_38152);
and U38479 (N_38479,N_38206,N_38057);
and U38480 (N_38480,N_38223,N_38248);
nand U38481 (N_38481,N_38219,N_38229);
and U38482 (N_38482,N_38234,N_38080);
and U38483 (N_38483,N_38233,N_38048);
nor U38484 (N_38484,N_38113,N_38187);
nor U38485 (N_38485,N_38241,N_38038);
or U38486 (N_38486,N_38018,N_38038);
nand U38487 (N_38487,N_38123,N_38102);
or U38488 (N_38488,N_38005,N_38014);
or U38489 (N_38489,N_38122,N_38045);
and U38490 (N_38490,N_38107,N_38064);
nor U38491 (N_38491,N_38075,N_38012);
xor U38492 (N_38492,N_38212,N_38026);
nor U38493 (N_38493,N_38226,N_38059);
nor U38494 (N_38494,N_38193,N_38241);
and U38495 (N_38495,N_38092,N_38205);
nand U38496 (N_38496,N_38008,N_38091);
or U38497 (N_38497,N_38020,N_38048);
or U38498 (N_38498,N_38085,N_38151);
or U38499 (N_38499,N_38182,N_38203);
xnor U38500 (N_38500,N_38435,N_38441);
nand U38501 (N_38501,N_38298,N_38389);
nand U38502 (N_38502,N_38343,N_38271);
nand U38503 (N_38503,N_38407,N_38348);
nand U38504 (N_38504,N_38466,N_38377);
xor U38505 (N_38505,N_38293,N_38374);
and U38506 (N_38506,N_38302,N_38439);
nand U38507 (N_38507,N_38290,N_38498);
xnor U38508 (N_38508,N_38264,N_38474);
nor U38509 (N_38509,N_38419,N_38438);
nor U38510 (N_38510,N_38266,N_38433);
nor U38511 (N_38511,N_38468,N_38454);
nor U38512 (N_38512,N_38379,N_38285);
and U38513 (N_38513,N_38375,N_38345);
xnor U38514 (N_38514,N_38294,N_38309);
nor U38515 (N_38515,N_38323,N_38284);
or U38516 (N_38516,N_38486,N_38333);
or U38517 (N_38517,N_38299,N_38459);
nor U38518 (N_38518,N_38378,N_38443);
and U38519 (N_38519,N_38316,N_38395);
nand U38520 (N_38520,N_38364,N_38278);
and U38521 (N_38521,N_38337,N_38499);
nor U38522 (N_38522,N_38366,N_38250);
or U38523 (N_38523,N_38444,N_38445);
nand U38524 (N_38524,N_38352,N_38307);
xor U38525 (N_38525,N_38400,N_38431);
or U38526 (N_38526,N_38350,N_38256);
nand U38527 (N_38527,N_38465,N_38283);
and U38528 (N_38528,N_38257,N_38406);
xnor U38529 (N_38529,N_38403,N_38413);
nor U38530 (N_38530,N_38399,N_38252);
xnor U38531 (N_38531,N_38341,N_38417);
nand U38532 (N_38532,N_38280,N_38460);
xnor U38533 (N_38533,N_38429,N_38321);
xor U38534 (N_38534,N_38416,N_38281);
or U38535 (N_38535,N_38484,N_38367);
xor U38536 (N_38536,N_38488,N_38356);
nand U38537 (N_38537,N_38329,N_38408);
nand U38538 (N_38538,N_38472,N_38275);
xnor U38539 (N_38539,N_38286,N_38267);
nand U38540 (N_38540,N_38258,N_38423);
and U38541 (N_38541,N_38317,N_38482);
nor U38542 (N_38542,N_38402,N_38253);
xnor U38543 (N_38543,N_38360,N_38453);
or U38544 (N_38544,N_38430,N_38291);
nor U38545 (N_38545,N_38344,N_38462);
or U38546 (N_38546,N_38437,N_38397);
nor U38547 (N_38547,N_38411,N_38491);
nor U38548 (N_38548,N_38426,N_38305);
and U38549 (N_38549,N_38268,N_38369);
nand U38550 (N_38550,N_38479,N_38464);
and U38551 (N_38551,N_38440,N_38306);
xor U38552 (N_38552,N_38361,N_38476);
and U38553 (N_38553,N_38382,N_38392);
or U38554 (N_38554,N_38446,N_38383);
nand U38555 (N_38555,N_38262,N_38292);
and U38556 (N_38556,N_38372,N_38297);
and U38557 (N_38557,N_38398,N_38418);
and U38558 (N_38558,N_38296,N_38477);
nand U38559 (N_38559,N_38370,N_38363);
or U38560 (N_38560,N_38422,N_38480);
xnor U38561 (N_38561,N_38319,N_38492);
nand U38562 (N_38562,N_38475,N_38269);
nand U38563 (N_38563,N_38357,N_38457);
xnor U38564 (N_38564,N_38282,N_38434);
nand U38565 (N_38565,N_38261,N_38469);
or U38566 (N_38566,N_38331,N_38335);
and U38567 (N_38567,N_38303,N_38270);
xor U38568 (N_38568,N_38428,N_38390);
xnor U38569 (N_38569,N_38421,N_38458);
nand U38570 (N_38570,N_38455,N_38481);
nand U38571 (N_38571,N_38373,N_38355);
nor U38572 (N_38572,N_38489,N_38362);
or U38573 (N_38573,N_38387,N_38495);
xor U38574 (N_38574,N_38409,N_38386);
nor U38575 (N_38575,N_38388,N_38276);
xnor U38576 (N_38576,N_38322,N_38315);
xor U38577 (N_38577,N_38277,N_38424);
xor U38578 (N_38578,N_38336,N_38456);
and U38579 (N_38579,N_38328,N_38354);
nor U38580 (N_38580,N_38427,N_38394);
nand U38581 (N_38581,N_38461,N_38471);
and U38582 (N_38582,N_38371,N_38310);
nand U38583 (N_38583,N_38405,N_38334);
xnor U38584 (N_38584,N_38380,N_38442);
nand U38585 (N_38585,N_38254,N_38393);
nor U38586 (N_38586,N_38436,N_38308);
or U38587 (N_38587,N_38487,N_38263);
nand U38588 (N_38588,N_38287,N_38396);
and U38589 (N_38589,N_38485,N_38314);
xor U38590 (N_38590,N_38324,N_38415);
or U38591 (N_38591,N_38432,N_38320);
nand U38592 (N_38592,N_38449,N_38300);
nor U38593 (N_38593,N_38295,N_38385);
or U38594 (N_38594,N_38412,N_38391);
nor U38595 (N_38595,N_38255,N_38332);
or U38596 (N_38596,N_38312,N_38326);
or U38597 (N_38597,N_38493,N_38497);
nand U38598 (N_38598,N_38410,N_38483);
nor U38599 (N_38599,N_38384,N_38447);
nand U38600 (N_38600,N_38289,N_38414);
nand U38601 (N_38601,N_38274,N_38470);
or U38602 (N_38602,N_38401,N_38490);
or U38603 (N_38603,N_38451,N_38381);
or U38604 (N_38604,N_38342,N_38376);
xnor U38605 (N_38605,N_38318,N_38325);
or U38606 (N_38606,N_38368,N_38313);
and U38607 (N_38607,N_38494,N_38330);
or U38608 (N_38608,N_38279,N_38478);
nand U38609 (N_38609,N_38359,N_38288);
and U38610 (N_38610,N_38346,N_38273);
nand U38611 (N_38611,N_38340,N_38450);
xor U38612 (N_38612,N_38452,N_38358);
nor U38613 (N_38613,N_38351,N_38311);
or U38614 (N_38614,N_38304,N_38347);
or U38615 (N_38615,N_38265,N_38272);
xnor U38616 (N_38616,N_38448,N_38463);
nor U38617 (N_38617,N_38338,N_38404);
nand U38618 (N_38618,N_38259,N_38496);
nor U38619 (N_38619,N_38349,N_38301);
or U38620 (N_38620,N_38420,N_38473);
nor U38621 (N_38621,N_38260,N_38251);
or U38622 (N_38622,N_38365,N_38425);
or U38623 (N_38623,N_38339,N_38327);
nor U38624 (N_38624,N_38467,N_38353);
nor U38625 (N_38625,N_38431,N_38363);
and U38626 (N_38626,N_38450,N_38375);
nor U38627 (N_38627,N_38264,N_38407);
nor U38628 (N_38628,N_38348,N_38489);
nor U38629 (N_38629,N_38319,N_38350);
nand U38630 (N_38630,N_38320,N_38428);
and U38631 (N_38631,N_38287,N_38406);
nand U38632 (N_38632,N_38470,N_38492);
or U38633 (N_38633,N_38293,N_38340);
nor U38634 (N_38634,N_38334,N_38363);
xor U38635 (N_38635,N_38432,N_38343);
nor U38636 (N_38636,N_38431,N_38373);
and U38637 (N_38637,N_38497,N_38471);
xnor U38638 (N_38638,N_38340,N_38392);
or U38639 (N_38639,N_38482,N_38393);
and U38640 (N_38640,N_38306,N_38358);
and U38641 (N_38641,N_38300,N_38290);
xnor U38642 (N_38642,N_38306,N_38330);
or U38643 (N_38643,N_38338,N_38378);
nand U38644 (N_38644,N_38480,N_38371);
nor U38645 (N_38645,N_38293,N_38368);
xnor U38646 (N_38646,N_38340,N_38461);
nand U38647 (N_38647,N_38479,N_38355);
nand U38648 (N_38648,N_38453,N_38444);
or U38649 (N_38649,N_38324,N_38438);
nand U38650 (N_38650,N_38443,N_38430);
or U38651 (N_38651,N_38469,N_38439);
nor U38652 (N_38652,N_38383,N_38265);
xnor U38653 (N_38653,N_38457,N_38363);
nor U38654 (N_38654,N_38370,N_38387);
or U38655 (N_38655,N_38270,N_38447);
or U38656 (N_38656,N_38348,N_38302);
or U38657 (N_38657,N_38338,N_38363);
and U38658 (N_38658,N_38403,N_38389);
nand U38659 (N_38659,N_38435,N_38313);
nand U38660 (N_38660,N_38275,N_38395);
nand U38661 (N_38661,N_38461,N_38372);
or U38662 (N_38662,N_38296,N_38470);
nand U38663 (N_38663,N_38436,N_38344);
xnor U38664 (N_38664,N_38339,N_38253);
or U38665 (N_38665,N_38356,N_38281);
nor U38666 (N_38666,N_38457,N_38390);
or U38667 (N_38667,N_38259,N_38360);
or U38668 (N_38668,N_38372,N_38251);
nand U38669 (N_38669,N_38387,N_38335);
xor U38670 (N_38670,N_38499,N_38455);
and U38671 (N_38671,N_38318,N_38450);
nor U38672 (N_38672,N_38282,N_38423);
and U38673 (N_38673,N_38464,N_38256);
nor U38674 (N_38674,N_38292,N_38405);
and U38675 (N_38675,N_38314,N_38374);
nand U38676 (N_38676,N_38257,N_38290);
xnor U38677 (N_38677,N_38465,N_38289);
or U38678 (N_38678,N_38337,N_38302);
and U38679 (N_38679,N_38291,N_38391);
xor U38680 (N_38680,N_38272,N_38317);
nand U38681 (N_38681,N_38272,N_38435);
nand U38682 (N_38682,N_38296,N_38402);
nor U38683 (N_38683,N_38304,N_38415);
nor U38684 (N_38684,N_38265,N_38371);
xor U38685 (N_38685,N_38329,N_38326);
xnor U38686 (N_38686,N_38267,N_38341);
xnor U38687 (N_38687,N_38253,N_38374);
and U38688 (N_38688,N_38277,N_38406);
xor U38689 (N_38689,N_38453,N_38274);
or U38690 (N_38690,N_38291,N_38348);
nand U38691 (N_38691,N_38449,N_38438);
nand U38692 (N_38692,N_38475,N_38413);
xnor U38693 (N_38693,N_38387,N_38379);
nor U38694 (N_38694,N_38481,N_38386);
nand U38695 (N_38695,N_38357,N_38430);
or U38696 (N_38696,N_38354,N_38266);
nand U38697 (N_38697,N_38361,N_38294);
or U38698 (N_38698,N_38382,N_38296);
nand U38699 (N_38699,N_38465,N_38303);
or U38700 (N_38700,N_38458,N_38399);
xor U38701 (N_38701,N_38452,N_38306);
or U38702 (N_38702,N_38491,N_38271);
nand U38703 (N_38703,N_38286,N_38317);
or U38704 (N_38704,N_38377,N_38472);
or U38705 (N_38705,N_38394,N_38280);
and U38706 (N_38706,N_38373,N_38415);
nand U38707 (N_38707,N_38444,N_38408);
xor U38708 (N_38708,N_38363,N_38299);
and U38709 (N_38709,N_38383,N_38287);
or U38710 (N_38710,N_38323,N_38348);
nand U38711 (N_38711,N_38304,N_38398);
nor U38712 (N_38712,N_38465,N_38372);
nand U38713 (N_38713,N_38434,N_38302);
nor U38714 (N_38714,N_38459,N_38372);
xnor U38715 (N_38715,N_38353,N_38391);
or U38716 (N_38716,N_38342,N_38263);
nor U38717 (N_38717,N_38305,N_38491);
nor U38718 (N_38718,N_38447,N_38345);
nand U38719 (N_38719,N_38326,N_38330);
and U38720 (N_38720,N_38347,N_38400);
nor U38721 (N_38721,N_38308,N_38263);
and U38722 (N_38722,N_38420,N_38354);
xnor U38723 (N_38723,N_38406,N_38261);
or U38724 (N_38724,N_38444,N_38376);
or U38725 (N_38725,N_38406,N_38485);
nor U38726 (N_38726,N_38383,N_38308);
or U38727 (N_38727,N_38473,N_38306);
nor U38728 (N_38728,N_38424,N_38472);
nor U38729 (N_38729,N_38399,N_38358);
or U38730 (N_38730,N_38469,N_38488);
nand U38731 (N_38731,N_38337,N_38341);
xor U38732 (N_38732,N_38339,N_38303);
nor U38733 (N_38733,N_38389,N_38478);
nor U38734 (N_38734,N_38414,N_38296);
and U38735 (N_38735,N_38346,N_38364);
nor U38736 (N_38736,N_38459,N_38321);
xor U38737 (N_38737,N_38275,N_38311);
nand U38738 (N_38738,N_38477,N_38412);
or U38739 (N_38739,N_38390,N_38279);
xor U38740 (N_38740,N_38393,N_38291);
nor U38741 (N_38741,N_38271,N_38496);
and U38742 (N_38742,N_38370,N_38284);
nand U38743 (N_38743,N_38475,N_38453);
xor U38744 (N_38744,N_38446,N_38409);
nand U38745 (N_38745,N_38316,N_38373);
or U38746 (N_38746,N_38359,N_38352);
or U38747 (N_38747,N_38459,N_38312);
and U38748 (N_38748,N_38360,N_38408);
nor U38749 (N_38749,N_38463,N_38334);
or U38750 (N_38750,N_38640,N_38623);
xnor U38751 (N_38751,N_38677,N_38680);
and U38752 (N_38752,N_38575,N_38657);
nor U38753 (N_38753,N_38667,N_38707);
xnor U38754 (N_38754,N_38741,N_38565);
xnor U38755 (N_38755,N_38549,N_38654);
or U38756 (N_38756,N_38560,N_38647);
nand U38757 (N_38757,N_38544,N_38691);
nand U38758 (N_38758,N_38642,N_38532);
nand U38759 (N_38759,N_38679,N_38606);
nand U38760 (N_38760,N_38619,N_38632);
nand U38761 (N_38761,N_38607,N_38730);
nand U38762 (N_38762,N_38625,N_38537);
xor U38763 (N_38763,N_38701,N_38683);
nand U38764 (N_38764,N_38681,N_38569);
or U38765 (N_38765,N_38540,N_38535);
or U38766 (N_38766,N_38543,N_38704);
nand U38767 (N_38767,N_38500,N_38586);
nand U38768 (N_38768,N_38558,N_38744);
or U38769 (N_38769,N_38655,N_38736);
or U38770 (N_38770,N_38637,N_38551);
or U38771 (N_38771,N_38723,N_38644);
nor U38772 (N_38772,N_38676,N_38511);
xnor U38773 (N_38773,N_38627,N_38717);
nand U38774 (N_38774,N_38584,N_38663);
nor U38775 (N_38775,N_38574,N_38539);
nand U38776 (N_38776,N_38698,N_38616);
nor U38777 (N_38777,N_38692,N_38602);
and U38778 (N_38778,N_38664,N_38641);
or U38779 (N_38779,N_38635,N_38579);
nor U38780 (N_38780,N_38588,N_38656);
nand U38781 (N_38781,N_38702,N_38621);
nor U38782 (N_38782,N_38706,N_38738);
nor U38783 (N_38783,N_38518,N_38709);
nand U38784 (N_38784,N_38572,N_38562);
and U38785 (N_38785,N_38697,N_38556);
xor U38786 (N_38786,N_38720,N_38716);
or U38787 (N_38787,N_38733,N_38514);
or U38788 (N_38788,N_38576,N_38638);
xor U38789 (N_38789,N_38665,N_38604);
or U38790 (N_38790,N_38531,N_38649);
xor U38791 (N_38791,N_38520,N_38687);
nand U38792 (N_38792,N_38748,N_38675);
and U38793 (N_38793,N_38737,N_38506);
nand U38794 (N_38794,N_38587,N_38591);
nand U38795 (N_38795,N_38609,N_38601);
xnor U38796 (N_38796,N_38521,N_38739);
xnor U38797 (N_38797,N_38600,N_38710);
or U38798 (N_38798,N_38512,N_38583);
and U38799 (N_38799,N_38618,N_38745);
nor U38800 (N_38800,N_38645,N_38548);
xor U38801 (N_38801,N_38564,N_38527);
or U38802 (N_38802,N_38732,N_38617);
xnor U38803 (N_38803,N_38554,N_38525);
and U38804 (N_38804,N_38747,N_38613);
xnor U38805 (N_38805,N_38594,N_38711);
or U38806 (N_38806,N_38721,N_38507);
nand U38807 (N_38807,N_38712,N_38626);
or U38808 (N_38808,N_38630,N_38529);
nor U38809 (N_38809,N_38533,N_38568);
or U38810 (N_38810,N_38666,N_38705);
or U38811 (N_38811,N_38610,N_38678);
xor U38812 (N_38812,N_38651,N_38605);
or U38813 (N_38813,N_38689,N_38585);
nor U38814 (N_38814,N_38582,N_38684);
xor U38815 (N_38815,N_38559,N_38530);
and U38816 (N_38816,N_38633,N_38573);
xnor U38817 (N_38817,N_38524,N_38714);
nor U38818 (N_38818,N_38670,N_38749);
nand U38819 (N_38819,N_38690,N_38567);
nor U38820 (N_38820,N_38546,N_38501);
nand U38821 (N_38821,N_38740,N_38636);
xnor U38822 (N_38822,N_38552,N_38693);
nor U38823 (N_38823,N_38671,N_38713);
nor U38824 (N_38824,N_38597,N_38728);
and U38825 (N_38825,N_38515,N_38603);
xor U38826 (N_38826,N_38542,N_38608);
xnor U38827 (N_38827,N_38615,N_38550);
nor U38828 (N_38828,N_38528,N_38646);
or U38829 (N_38829,N_38503,N_38522);
nand U38830 (N_38830,N_38699,N_38650);
xnor U38831 (N_38831,N_38547,N_38624);
nand U38832 (N_38832,N_38726,N_38545);
nand U38833 (N_38833,N_38566,N_38611);
xor U38834 (N_38834,N_38660,N_38599);
and U38835 (N_38835,N_38502,N_38508);
or U38836 (N_38836,N_38553,N_38735);
nand U38837 (N_38837,N_38563,N_38534);
or U38838 (N_38838,N_38622,N_38561);
xor U38839 (N_38839,N_38504,N_38694);
nand U38840 (N_38840,N_38703,N_38648);
and U38841 (N_38841,N_38672,N_38571);
xor U38842 (N_38842,N_38743,N_38513);
nand U38843 (N_38843,N_38653,N_38589);
nand U38844 (N_38844,N_38580,N_38727);
and U38845 (N_38845,N_38592,N_38612);
or U38846 (N_38846,N_38538,N_38541);
nor U38847 (N_38847,N_38696,N_38746);
nand U38848 (N_38848,N_38517,N_38685);
or U38849 (N_38849,N_38628,N_38700);
and U38850 (N_38850,N_38629,N_38510);
nand U38851 (N_38851,N_38634,N_38590);
xnor U38852 (N_38852,N_38724,N_38570);
xor U38853 (N_38853,N_38719,N_38742);
and U38854 (N_38854,N_38686,N_38526);
nand U38855 (N_38855,N_38734,N_38523);
or U38856 (N_38856,N_38639,N_38668);
and U38857 (N_38857,N_38652,N_38536);
nor U38858 (N_38858,N_38595,N_38620);
nand U38859 (N_38859,N_38643,N_38722);
or U38860 (N_38860,N_38673,N_38516);
nor U38861 (N_38861,N_38674,N_38658);
nand U38862 (N_38862,N_38661,N_38669);
or U38863 (N_38863,N_38659,N_38577);
or U38864 (N_38864,N_38688,N_38578);
and U38865 (N_38865,N_38718,N_38581);
or U38866 (N_38866,N_38725,N_38731);
or U38867 (N_38867,N_38631,N_38614);
nor U38868 (N_38868,N_38509,N_38593);
or U38869 (N_38869,N_38557,N_38596);
xnor U38870 (N_38870,N_38505,N_38715);
nor U38871 (N_38871,N_38729,N_38708);
nor U38872 (N_38872,N_38555,N_38662);
or U38873 (N_38873,N_38682,N_38519);
nand U38874 (N_38874,N_38598,N_38695);
nand U38875 (N_38875,N_38680,N_38739);
or U38876 (N_38876,N_38577,N_38616);
nor U38877 (N_38877,N_38691,N_38583);
nor U38878 (N_38878,N_38748,N_38649);
or U38879 (N_38879,N_38565,N_38564);
xnor U38880 (N_38880,N_38749,N_38688);
nor U38881 (N_38881,N_38603,N_38672);
nor U38882 (N_38882,N_38545,N_38664);
xor U38883 (N_38883,N_38520,N_38747);
nand U38884 (N_38884,N_38701,N_38661);
nor U38885 (N_38885,N_38693,N_38641);
nor U38886 (N_38886,N_38721,N_38644);
nand U38887 (N_38887,N_38704,N_38731);
xor U38888 (N_38888,N_38653,N_38538);
or U38889 (N_38889,N_38726,N_38583);
xor U38890 (N_38890,N_38534,N_38512);
nor U38891 (N_38891,N_38720,N_38596);
xnor U38892 (N_38892,N_38658,N_38501);
nand U38893 (N_38893,N_38553,N_38619);
and U38894 (N_38894,N_38561,N_38669);
nand U38895 (N_38895,N_38648,N_38746);
or U38896 (N_38896,N_38662,N_38627);
nor U38897 (N_38897,N_38521,N_38505);
nor U38898 (N_38898,N_38661,N_38686);
xnor U38899 (N_38899,N_38743,N_38655);
xor U38900 (N_38900,N_38739,N_38590);
or U38901 (N_38901,N_38680,N_38601);
or U38902 (N_38902,N_38688,N_38590);
nor U38903 (N_38903,N_38722,N_38705);
nor U38904 (N_38904,N_38515,N_38531);
xnor U38905 (N_38905,N_38675,N_38677);
and U38906 (N_38906,N_38627,N_38570);
and U38907 (N_38907,N_38630,N_38564);
nand U38908 (N_38908,N_38683,N_38618);
and U38909 (N_38909,N_38618,N_38735);
and U38910 (N_38910,N_38526,N_38707);
xnor U38911 (N_38911,N_38700,N_38512);
or U38912 (N_38912,N_38726,N_38560);
or U38913 (N_38913,N_38596,N_38671);
or U38914 (N_38914,N_38539,N_38679);
nand U38915 (N_38915,N_38589,N_38567);
nand U38916 (N_38916,N_38511,N_38541);
nand U38917 (N_38917,N_38680,N_38670);
nand U38918 (N_38918,N_38732,N_38612);
nand U38919 (N_38919,N_38536,N_38551);
and U38920 (N_38920,N_38721,N_38698);
xor U38921 (N_38921,N_38710,N_38713);
or U38922 (N_38922,N_38568,N_38618);
or U38923 (N_38923,N_38743,N_38588);
or U38924 (N_38924,N_38716,N_38725);
and U38925 (N_38925,N_38531,N_38623);
nand U38926 (N_38926,N_38598,N_38682);
or U38927 (N_38927,N_38501,N_38543);
xnor U38928 (N_38928,N_38582,N_38541);
or U38929 (N_38929,N_38733,N_38728);
nand U38930 (N_38930,N_38611,N_38642);
nand U38931 (N_38931,N_38619,N_38616);
nor U38932 (N_38932,N_38746,N_38713);
or U38933 (N_38933,N_38622,N_38650);
and U38934 (N_38934,N_38654,N_38657);
nand U38935 (N_38935,N_38629,N_38558);
nor U38936 (N_38936,N_38658,N_38600);
and U38937 (N_38937,N_38639,N_38729);
or U38938 (N_38938,N_38621,N_38540);
or U38939 (N_38939,N_38576,N_38676);
or U38940 (N_38940,N_38708,N_38553);
or U38941 (N_38941,N_38645,N_38522);
nor U38942 (N_38942,N_38557,N_38654);
and U38943 (N_38943,N_38621,N_38513);
and U38944 (N_38944,N_38652,N_38506);
or U38945 (N_38945,N_38705,N_38650);
or U38946 (N_38946,N_38507,N_38512);
or U38947 (N_38947,N_38733,N_38719);
nand U38948 (N_38948,N_38519,N_38567);
nor U38949 (N_38949,N_38609,N_38566);
xor U38950 (N_38950,N_38712,N_38572);
nand U38951 (N_38951,N_38642,N_38578);
nor U38952 (N_38952,N_38525,N_38679);
or U38953 (N_38953,N_38745,N_38559);
or U38954 (N_38954,N_38567,N_38640);
or U38955 (N_38955,N_38537,N_38551);
or U38956 (N_38956,N_38524,N_38672);
or U38957 (N_38957,N_38552,N_38703);
or U38958 (N_38958,N_38545,N_38659);
xor U38959 (N_38959,N_38703,N_38510);
xor U38960 (N_38960,N_38671,N_38670);
and U38961 (N_38961,N_38701,N_38705);
xor U38962 (N_38962,N_38644,N_38694);
or U38963 (N_38963,N_38574,N_38623);
nor U38964 (N_38964,N_38693,N_38662);
or U38965 (N_38965,N_38658,N_38739);
nor U38966 (N_38966,N_38657,N_38604);
or U38967 (N_38967,N_38509,N_38677);
or U38968 (N_38968,N_38689,N_38591);
xnor U38969 (N_38969,N_38657,N_38595);
or U38970 (N_38970,N_38704,N_38565);
nand U38971 (N_38971,N_38591,N_38548);
nor U38972 (N_38972,N_38516,N_38670);
nor U38973 (N_38973,N_38536,N_38719);
nand U38974 (N_38974,N_38659,N_38618);
or U38975 (N_38975,N_38558,N_38521);
and U38976 (N_38976,N_38612,N_38580);
and U38977 (N_38977,N_38605,N_38500);
or U38978 (N_38978,N_38657,N_38659);
nor U38979 (N_38979,N_38576,N_38683);
or U38980 (N_38980,N_38554,N_38667);
nand U38981 (N_38981,N_38637,N_38561);
nand U38982 (N_38982,N_38501,N_38706);
and U38983 (N_38983,N_38571,N_38703);
nand U38984 (N_38984,N_38664,N_38553);
and U38985 (N_38985,N_38654,N_38608);
and U38986 (N_38986,N_38697,N_38596);
nand U38987 (N_38987,N_38582,N_38667);
and U38988 (N_38988,N_38698,N_38737);
nor U38989 (N_38989,N_38668,N_38592);
and U38990 (N_38990,N_38531,N_38734);
nand U38991 (N_38991,N_38594,N_38520);
or U38992 (N_38992,N_38585,N_38730);
and U38993 (N_38993,N_38638,N_38560);
nand U38994 (N_38994,N_38701,N_38557);
or U38995 (N_38995,N_38513,N_38664);
and U38996 (N_38996,N_38584,N_38675);
and U38997 (N_38997,N_38645,N_38666);
nor U38998 (N_38998,N_38692,N_38619);
nor U38999 (N_38999,N_38609,N_38689);
and U39000 (N_39000,N_38786,N_38939);
and U39001 (N_39001,N_38992,N_38836);
and U39002 (N_39002,N_38973,N_38822);
nand U39003 (N_39003,N_38809,N_38837);
nand U39004 (N_39004,N_38814,N_38932);
nor U39005 (N_39005,N_38793,N_38885);
nor U39006 (N_39006,N_38870,N_38859);
nor U39007 (N_39007,N_38785,N_38926);
nand U39008 (N_39008,N_38883,N_38869);
or U39009 (N_39009,N_38994,N_38899);
or U39010 (N_39010,N_38964,N_38878);
and U39011 (N_39011,N_38820,N_38982);
xor U39012 (N_39012,N_38828,N_38882);
nor U39013 (N_39013,N_38936,N_38852);
and U39014 (N_39014,N_38796,N_38849);
nor U39015 (N_39015,N_38950,N_38933);
nand U39016 (N_39016,N_38881,N_38753);
nand U39017 (N_39017,N_38774,N_38951);
and U39018 (N_39018,N_38832,N_38845);
xor U39019 (N_39019,N_38897,N_38799);
xnor U39020 (N_39020,N_38771,N_38759);
nor U39021 (N_39021,N_38958,N_38967);
nor U39022 (N_39022,N_38857,N_38977);
and U39023 (N_39023,N_38969,N_38942);
xor U39024 (N_39024,N_38756,N_38829);
nor U39025 (N_39025,N_38779,N_38839);
nand U39026 (N_39026,N_38993,N_38998);
nor U39027 (N_39027,N_38776,N_38990);
or U39028 (N_39028,N_38818,N_38811);
nor U39029 (N_39029,N_38780,N_38900);
and U39030 (N_39030,N_38815,N_38928);
and U39031 (N_39031,N_38821,N_38914);
xnor U39032 (N_39032,N_38971,N_38922);
xnor U39033 (N_39033,N_38854,N_38850);
nor U39034 (N_39034,N_38924,N_38980);
nand U39035 (N_39035,N_38807,N_38901);
and U39036 (N_39036,N_38961,N_38787);
and U39037 (N_39037,N_38941,N_38817);
or U39038 (N_39038,N_38840,N_38848);
xnor U39039 (N_39039,N_38763,N_38920);
nand U39040 (N_39040,N_38898,N_38947);
or U39041 (N_39041,N_38868,N_38910);
nand U39042 (N_39042,N_38887,N_38810);
nand U39043 (N_39043,N_38877,N_38937);
and U39044 (N_39044,N_38988,N_38794);
and U39045 (N_39045,N_38875,N_38798);
or U39046 (N_39046,N_38767,N_38955);
nor U39047 (N_39047,N_38792,N_38931);
or U39048 (N_39048,N_38880,N_38865);
xnor U39049 (N_39049,N_38795,N_38975);
or U39050 (N_39050,N_38803,N_38952);
and U39051 (N_39051,N_38874,N_38861);
nand U39052 (N_39052,N_38921,N_38758);
or U39053 (N_39053,N_38761,N_38907);
nand U39054 (N_39054,N_38890,N_38813);
nor U39055 (N_39055,N_38866,N_38835);
nor U39056 (N_39056,N_38824,N_38927);
nand U39057 (N_39057,N_38784,N_38972);
xor U39058 (N_39058,N_38764,N_38903);
and U39059 (N_39059,N_38996,N_38935);
or U39060 (N_39060,N_38986,N_38984);
xnor U39061 (N_39061,N_38770,N_38826);
or U39062 (N_39062,N_38871,N_38889);
and U39063 (N_39063,N_38773,N_38884);
nor U39064 (N_39064,N_38790,N_38915);
and U39065 (N_39065,N_38772,N_38905);
and U39066 (N_39066,N_38844,N_38760);
nand U39067 (N_39067,N_38917,N_38954);
or U39068 (N_39068,N_38909,N_38768);
nand U39069 (N_39069,N_38962,N_38976);
and U39070 (N_39070,N_38804,N_38755);
xnor U39071 (N_39071,N_38892,N_38919);
nand U39072 (N_39072,N_38830,N_38775);
or U39073 (N_39073,N_38991,N_38841);
or U39074 (N_39074,N_38904,N_38968);
xor U39075 (N_39075,N_38953,N_38938);
xnor U39076 (N_39076,N_38987,N_38965);
xnor U39077 (N_39077,N_38856,N_38800);
xnor U39078 (N_39078,N_38978,N_38782);
or U39079 (N_39079,N_38985,N_38929);
nand U39080 (N_39080,N_38806,N_38959);
nand U39081 (N_39081,N_38940,N_38970);
nand U39082 (N_39082,N_38918,N_38823);
nand U39083 (N_39083,N_38974,N_38778);
or U39084 (N_39084,N_38966,N_38944);
nand U39085 (N_39085,N_38949,N_38834);
or U39086 (N_39086,N_38888,N_38989);
nand U39087 (N_39087,N_38934,N_38956);
or U39088 (N_39088,N_38825,N_38960);
nand U39089 (N_39089,N_38957,N_38902);
xnor U39090 (N_39090,N_38802,N_38752);
nand U39091 (N_39091,N_38851,N_38943);
and U39092 (N_39092,N_38963,N_38801);
and U39093 (N_39093,N_38831,N_38913);
xor U39094 (N_39094,N_38896,N_38911);
or U39095 (N_39095,N_38846,N_38999);
or U39096 (N_39096,N_38766,N_38751);
nand U39097 (N_39097,N_38946,N_38750);
or U39098 (N_39098,N_38789,N_38908);
nor U39099 (N_39099,N_38981,N_38879);
xnor U39100 (N_39100,N_38847,N_38769);
or U39101 (N_39101,N_38791,N_38906);
or U39102 (N_39102,N_38827,N_38762);
xnor U39103 (N_39103,N_38873,N_38808);
nand U39104 (N_39104,N_38872,N_38816);
nand U39105 (N_39105,N_38945,N_38788);
nand U39106 (N_39106,N_38916,N_38777);
or U39107 (N_39107,N_38860,N_38855);
nand U39108 (N_39108,N_38925,N_38765);
nand U39109 (N_39109,N_38754,N_38833);
and U39110 (N_39110,N_38862,N_38864);
nand U39111 (N_39111,N_38812,N_38781);
nand U39112 (N_39112,N_38783,N_38819);
nor U39113 (N_39113,N_38983,N_38853);
xnor U39114 (N_39114,N_38995,N_38979);
xnor U39115 (N_39115,N_38858,N_38805);
xnor U39116 (N_39116,N_38886,N_38797);
and U39117 (N_39117,N_38838,N_38912);
or U39118 (N_39118,N_38876,N_38923);
nand U39119 (N_39119,N_38948,N_38895);
xnor U39120 (N_39120,N_38930,N_38867);
or U39121 (N_39121,N_38757,N_38843);
and U39122 (N_39122,N_38891,N_38894);
and U39123 (N_39123,N_38863,N_38997);
and U39124 (N_39124,N_38893,N_38842);
nand U39125 (N_39125,N_38758,N_38836);
or U39126 (N_39126,N_38985,N_38998);
xnor U39127 (N_39127,N_38988,N_38861);
xnor U39128 (N_39128,N_38908,N_38861);
xnor U39129 (N_39129,N_38832,N_38791);
xnor U39130 (N_39130,N_38919,N_38939);
and U39131 (N_39131,N_38866,N_38771);
or U39132 (N_39132,N_38994,N_38969);
nand U39133 (N_39133,N_38956,N_38986);
nand U39134 (N_39134,N_38965,N_38809);
and U39135 (N_39135,N_38804,N_38752);
nor U39136 (N_39136,N_38887,N_38814);
nand U39137 (N_39137,N_38786,N_38798);
or U39138 (N_39138,N_38822,N_38944);
xnor U39139 (N_39139,N_38922,N_38802);
or U39140 (N_39140,N_38753,N_38958);
nor U39141 (N_39141,N_38881,N_38901);
xor U39142 (N_39142,N_38878,N_38807);
and U39143 (N_39143,N_38981,N_38916);
nand U39144 (N_39144,N_38906,N_38763);
nand U39145 (N_39145,N_38947,N_38900);
nand U39146 (N_39146,N_38955,N_38892);
nand U39147 (N_39147,N_38753,N_38979);
and U39148 (N_39148,N_38868,N_38810);
and U39149 (N_39149,N_38816,N_38758);
xnor U39150 (N_39150,N_38984,N_38909);
nand U39151 (N_39151,N_38899,N_38828);
nor U39152 (N_39152,N_38953,N_38754);
or U39153 (N_39153,N_38994,N_38809);
or U39154 (N_39154,N_38898,N_38905);
or U39155 (N_39155,N_38923,N_38883);
nand U39156 (N_39156,N_38906,N_38925);
nand U39157 (N_39157,N_38938,N_38778);
xnor U39158 (N_39158,N_38881,N_38895);
nand U39159 (N_39159,N_38844,N_38984);
nor U39160 (N_39160,N_38754,N_38962);
nand U39161 (N_39161,N_38980,N_38818);
xor U39162 (N_39162,N_38827,N_38954);
xnor U39163 (N_39163,N_38756,N_38914);
or U39164 (N_39164,N_38856,N_38770);
and U39165 (N_39165,N_38845,N_38776);
xnor U39166 (N_39166,N_38986,N_38884);
and U39167 (N_39167,N_38801,N_38797);
nor U39168 (N_39168,N_38814,N_38752);
and U39169 (N_39169,N_38799,N_38911);
or U39170 (N_39170,N_38873,N_38903);
xor U39171 (N_39171,N_38963,N_38920);
xor U39172 (N_39172,N_38902,N_38911);
and U39173 (N_39173,N_38979,N_38960);
nor U39174 (N_39174,N_38905,N_38973);
nor U39175 (N_39175,N_38906,N_38801);
or U39176 (N_39176,N_38825,N_38785);
or U39177 (N_39177,N_38858,N_38882);
and U39178 (N_39178,N_38859,N_38838);
xor U39179 (N_39179,N_38925,N_38929);
and U39180 (N_39180,N_38776,N_38853);
nor U39181 (N_39181,N_38967,N_38852);
nor U39182 (N_39182,N_38938,N_38865);
and U39183 (N_39183,N_38857,N_38774);
and U39184 (N_39184,N_38983,N_38982);
nand U39185 (N_39185,N_38807,N_38893);
xor U39186 (N_39186,N_38784,N_38975);
and U39187 (N_39187,N_38858,N_38928);
nand U39188 (N_39188,N_38946,N_38945);
and U39189 (N_39189,N_38928,N_38860);
or U39190 (N_39190,N_38894,N_38895);
or U39191 (N_39191,N_38849,N_38879);
nor U39192 (N_39192,N_38866,N_38931);
xor U39193 (N_39193,N_38954,N_38903);
or U39194 (N_39194,N_38769,N_38843);
and U39195 (N_39195,N_38966,N_38856);
and U39196 (N_39196,N_38762,N_38798);
or U39197 (N_39197,N_38887,N_38812);
xnor U39198 (N_39198,N_38764,N_38931);
and U39199 (N_39199,N_38804,N_38800);
and U39200 (N_39200,N_38828,N_38929);
and U39201 (N_39201,N_38881,N_38769);
and U39202 (N_39202,N_38989,N_38762);
nor U39203 (N_39203,N_38990,N_38808);
or U39204 (N_39204,N_38900,N_38865);
xor U39205 (N_39205,N_38823,N_38912);
or U39206 (N_39206,N_38806,N_38852);
nand U39207 (N_39207,N_38990,N_38912);
nor U39208 (N_39208,N_38942,N_38861);
or U39209 (N_39209,N_38915,N_38907);
and U39210 (N_39210,N_38781,N_38960);
and U39211 (N_39211,N_38821,N_38874);
xor U39212 (N_39212,N_38917,N_38769);
xnor U39213 (N_39213,N_38836,N_38948);
nor U39214 (N_39214,N_38919,N_38795);
nor U39215 (N_39215,N_38868,N_38808);
xor U39216 (N_39216,N_38768,N_38810);
or U39217 (N_39217,N_38837,N_38817);
and U39218 (N_39218,N_38799,N_38808);
nand U39219 (N_39219,N_38815,N_38763);
nand U39220 (N_39220,N_38963,N_38765);
or U39221 (N_39221,N_38897,N_38878);
nor U39222 (N_39222,N_38996,N_38937);
xor U39223 (N_39223,N_38784,N_38934);
nand U39224 (N_39224,N_38996,N_38906);
and U39225 (N_39225,N_38972,N_38980);
xnor U39226 (N_39226,N_38903,N_38830);
nand U39227 (N_39227,N_38969,N_38770);
nand U39228 (N_39228,N_38758,N_38974);
xnor U39229 (N_39229,N_38789,N_38826);
or U39230 (N_39230,N_38851,N_38868);
xor U39231 (N_39231,N_38848,N_38958);
nand U39232 (N_39232,N_38940,N_38857);
and U39233 (N_39233,N_38819,N_38915);
xnor U39234 (N_39234,N_38803,N_38752);
nor U39235 (N_39235,N_38821,N_38868);
and U39236 (N_39236,N_38782,N_38805);
nor U39237 (N_39237,N_38752,N_38957);
nor U39238 (N_39238,N_38893,N_38924);
or U39239 (N_39239,N_38957,N_38781);
and U39240 (N_39240,N_38980,N_38756);
nand U39241 (N_39241,N_38897,N_38894);
xnor U39242 (N_39242,N_38776,N_38870);
xnor U39243 (N_39243,N_38767,N_38878);
nand U39244 (N_39244,N_38808,N_38923);
or U39245 (N_39245,N_38877,N_38842);
and U39246 (N_39246,N_38822,N_38804);
nor U39247 (N_39247,N_38763,N_38898);
and U39248 (N_39248,N_38821,N_38824);
and U39249 (N_39249,N_38874,N_38993);
or U39250 (N_39250,N_39243,N_39032);
nand U39251 (N_39251,N_39008,N_39169);
nand U39252 (N_39252,N_39121,N_39213);
and U39253 (N_39253,N_39176,N_39071);
xor U39254 (N_39254,N_39134,N_39181);
and U39255 (N_39255,N_39240,N_39068);
and U39256 (N_39256,N_39045,N_39137);
or U39257 (N_39257,N_39086,N_39233);
or U39258 (N_39258,N_39157,N_39160);
xor U39259 (N_39259,N_39234,N_39222);
nor U39260 (N_39260,N_39153,N_39190);
nor U39261 (N_39261,N_39195,N_39168);
nor U39262 (N_39262,N_39117,N_39067);
nor U39263 (N_39263,N_39170,N_39131);
or U39264 (N_39264,N_39080,N_39038);
xnor U39265 (N_39265,N_39029,N_39120);
and U39266 (N_39266,N_39196,N_39209);
nand U39267 (N_39267,N_39145,N_39217);
nand U39268 (N_39268,N_39013,N_39184);
nand U39269 (N_39269,N_39161,N_39207);
or U39270 (N_39270,N_39092,N_39057);
and U39271 (N_39271,N_39191,N_39167);
or U39272 (N_39272,N_39107,N_39185);
nor U39273 (N_39273,N_39087,N_39237);
or U39274 (N_39274,N_39159,N_39204);
and U39275 (N_39275,N_39065,N_39174);
nor U39276 (N_39276,N_39044,N_39116);
xnor U39277 (N_39277,N_39102,N_39178);
nor U39278 (N_39278,N_39151,N_39074);
xnor U39279 (N_39279,N_39199,N_39079);
nor U39280 (N_39280,N_39024,N_39113);
or U39281 (N_39281,N_39218,N_39039);
or U39282 (N_39282,N_39000,N_39111);
nand U39283 (N_39283,N_39123,N_39027);
and U39284 (N_39284,N_39022,N_39056);
or U39285 (N_39285,N_39104,N_39173);
and U39286 (N_39286,N_39136,N_39096);
or U39287 (N_39287,N_39011,N_39200);
xnor U39288 (N_39288,N_39081,N_39155);
nor U39289 (N_39289,N_39069,N_39221);
xnor U39290 (N_39290,N_39122,N_39227);
nand U39291 (N_39291,N_39208,N_39232);
and U39292 (N_39292,N_39015,N_39009);
xor U39293 (N_39293,N_39202,N_39051);
or U39294 (N_39294,N_39070,N_39211);
nor U39295 (N_39295,N_39100,N_39103);
and U39296 (N_39296,N_39165,N_39231);
nor U39297 (N_39297,N_39110,N_39006);
nand U39298 (N_39298,N_39140,N_39150);
or U39299 (N_39299,N_39099,N_39130);
nor U39300 (N_39300,N_39052,N_39028);
and U39301 (N_39301,N_39025,N_39152);
xor U39302 (N_39302,N_39050,N_39084);
xnor U39303 (N_39303,N_39215,N_39192);
or U39304 (N_39304,N_39047,N_39062);
xor U39305 (N_39305,N_39125,N_39246);
and U39306 (N_39306,N_39072,N_39059);
xor U39307 (N_39307,N_39097,N_39216);
nand U39308 (N_39308,N_39220,N_39203);
xnor U39309 (N_39309,N_39049,N_39054);
nor U39310 (N_39310,N_39205,N_39249);
nor U39311 (N_39311,N_39118,N_39172);
or U39312 (N_39312,N_39127,N_39020);
and U39313 (N_39313,N_39148,N_39033);
and U39314 (N_39314,N_39230,N_39193);
and U39315 (N_39315,N_39187,N_39035);
nor U39316 (N_39316,N_39241,N_39064);
and U39317 (N_39317,N_39010,N_39083);
nor U39318 (N_39318,N_39019,N_39034);
and U39319 (N_39319,N_39094,N_39177);
or U39320 (N_39320,N_39078,N_39154);
nor U39321 (N_39321,N_39139,N_39112);
xnor U39322 (N_39322,N_39090,N_39016);
xor U39323 (N_39323,N_39158,N_39183);
and U39324 (N_39324,N_39046,N_39194);
xor U39325 (N_39325,N_39077,N_39214);
nor U39326 (N_39326,N_39189,N_39001);
and U39327 (N_39327,N_39180,N_39138);
nor U39328 (N_39328,N_39023,N_39114);
xnor U39329 (N_39329,N_39229,N_39055);
nand U39330 (N_39330,N_39085,N_39095);
nand U39331 (N_39331,N_39042,N_39166);
xnor U39332 (N_39332,N_39223,N_39101);
or U39333 (N_39333,N_39026,N_39239);
or U39334 (N_39334,N_39012,N_39063);
and U39335 (N_39335,N_39030,N_39021);
and U39336 (N_39336,N_39198,N_39115);
or U39337 (N_39337,N_39133,N_39197);
or U39338 (N_39338,N_39048,N_39060);
xnor U39339 (N_39339,N_39212,N_39007);
nand U39340 (N_39340,N_39066,N_39201);
or U39341 (N_39341,N_39058,N_39129);
xnor U39342 (N_39342,N_39040,N_39098);
nand U39343 (N_39343,N_39242,N_39082);
or U39344 (N_39344,N_39163,N_39018);
or U39345 (N_39345,N_39002,N_39017);
xnor U39346 (N_39346,N_39108,N_39119);
nand U39347 (N_39347,N_39061,N_39142);
nand U39348 (N_39348,N_39188,N_39132);
and U39349 (N_39349,N_39124,N_39004);
or U39350 (N_39350,N_39126,N_39236);
xor U39351 (N_39351,N_39089,N_39244);
and U39352 (N_39352,N_39149,N_39106);
nand U39353 (N_39353,N_39031,N_39238);
nand U39354 (N_39354,N_39146,N_39135);
nand U39355 (N_39355,N_39093,N_39219);
xnor U39356 (N_39356,N_39105,N_39144);
xor U39357 (N_39357,N_39041,N_39186);
nand U39358 (N_39358,N_39206,N_39235);
or U39359 (N_39359,N_39224,N_39143);
nor U39360 (N_39360,N_39037,N_39141);
nand U39361 (N_39361,N_39171,N_39005);
nand U39362 (N_39362,N_39225,N_39014);
nand U39363 (N_39363,N_39091,N_39075);
nand U39364 (N_39364,N_39248,N_39073);
nor U39365 (N_39365,N_39228,N_39076);
nor U39366 (N_39366,N_39156,N_39179);
and U39367 (N_39367,N_39053,N_39164);
nand U39368 (N_39368,N_39088,N_39162);
or U39369 (N_39369,N_39210,N_39175);
xnor U39370 (N_39370,N_39109,N_39247);
and U39371 (N_39371,N_39003,N_39226);
or U39372 (N_39372,N_39128,N_39182);
or U39373 (N_39373,N_39147,N_39043);
and U39374 (N_39374,N_39245,N_39036);
or U39375 (N_39375,N_39184,N_39206);
xor U39376 (N_39376,N_39162,N_39157);
nor U39377 (N_39377,N_39151,N_39000);
and U39378 (N_39378,N_39199,N_39049);
xor U39379 (N_39379,N_39083,N_39077);
xor U39380 (N_39380,N_39144,N_39098);
nand U39381 (N_39381,N_39065,N_39144);
nor U39382 (N_39382,N_39131,N_39035);
nand U39383 (N_39383,N_39217,N_39123);
or U39384 (N_39384,N_39236,N_39157);
xnor U39385 (N_39385,N_39082,N_39117);
or U39386 (N_39386,N_39117,N_39087);
nand U39387 (N_39387,N_39155,N_39136);
nor U39388 (N_39388,N_39084,N_39077);
xnor U39389 (N_39389,N_39183,N_39071);
xnor U39390 (N_39390,N_39018,N_39017);
or U39391 (N_39391,N_39115,N_39223);
and U39392 (N_39392,N_39094,N_39114);
nor U39393 (N_39393,N_39063,N_39013);
and U39394 (N_39394,N_39044,N_39036);
nand U39395 (N_39395,N_39002,N_39125);
nand U39396 (N_39396,N_39206,N_39123);
or U39397 (N_39397,N_39140,N_39142);
nand U39398 (N_39398,N_39149,N_39089);
nand U39399 (N_39399,N_39114,N_39061);
or U39400 (N_39400,N_39132,N_39171);
or U39401 (N_39401,N_39245,N_39028);
nor U39402 (N_39402,N_39185,N_39032);
or U39403 (N_39403,N_39177,N_39021);
nor U39404 (N_39404,N_39106,N_39222);
or U39405 (N_39405,N_39022,N_39162);
and U39406 (N_39406,N_39192,N_39222);
and U39407 (N_39407,N_39052,N_39209);
nand U39408 (N_39408,N_39196,N_39087);
nor U39409 (N_39409,N_39157,N_39061);
xnor U39410 (N_39410,N_39115,N_39082);
or U39411 (N_39411,N_39081,N_39077);
xor U39412 (N_39412,N_39116,N_39049);
xor U39413 (N_39413,N_39178,N_39019);
and U39414 (N_39414,N_39242,N_39156);
and U39415 (N_39415,N_39089,N_39020);
and U39416 (N_39416,N_39194,N_39165);
xnor U39417 (N_39417,N_39012,N_39234);
or U39418 (N_39418,N_39218,N_39156);
and U39419 (N_39419,N_39220,N_39148);
nor U39420 (N_39420,N_39223,N_39084);
xnor U39421 (N_39421,N_39087,N_39241);
nor U39422 (N_39422,N_39228,N_39085);
or U39423 (N_39423,N_39009,N_39078);
or U39424 (N_39424,N_39211,N_39053);
or U39425 (N_39425,N_39076,N_39095);
and U39426 (N_39426,N_39001,N_39096);
and U39427 (N_39427,N_39249,N_39189);
or U39428 (N_39428,N_39204,N_39011);
nor U39429 (N_39429,N_39150,N_39148);
nor U39430 (N_39430,N_39006,N_39184);
or U39431 (N_39431,N_39045,N_39000);
nor U39432 (N_39432,N_39153,N_39019);
or U39433 (N_39433,N_39112,N_39079);
and U39434 (N_39434,N_39055,N_39184);
nand U39435 (N_39435,N_39188,N_39047);
or U39436 (N_39436,N_39018,N_39088);
or U39437 (N_39437,N_39208,N_39239);
nand U39438 (N_39438,N_39068,N_39033);
xor U39439 (N_39439,N_39002,N_39130);
nor U39440 (N_39440,N_39179,N_39182);
xor U39441 (N_39441,N_39076,N_39107);
or U39442 (N_39442,N_39234,N_39037);
xor U39443 (N_39443,N_39030,N_39196);
nand U39444 (N_39444,N_39150,N_39009);
nand U39445 (N_39445,N_39002,N_39105);
nor U39446 (N_39446,N_39148,N_39089);
or U39447 (N_39447,N_39224,N_39025);
nand U39448 (N_39448,N_39097,N_39213);
nor U39449 (N_39449,N_39172,N_39080);
or U39450 (N_39450,N_39138,N_39243);
and U39451 (N_39451,N_39035,N_39249);
nor U39452 (N_39452,N_39164,N_39166);
nand U39453 (N_39453,N_39073,N_39068);
nand U39454 (N_39454,N_39052,N_39082);
and U39455 (N_39455,N_39187,N_39050);
and U39456 (N_39456,N_39092,N_39132);
and U39457 (N_39457,N_39113,N_39116);
nand U39458 (N_39458,N_39172,N_39109);
and U39459 (N_39459,N_39036,N_39150);
and U39460 (N_39460,N_39134,N_39126);
nor U39461 (N_39461,N_39150,N_39054);
and U39462 (N_39462,N_39087,N_39027);
xor U39463 (N_39463,N_39242,N_39137);
or U39464 (N_39464,N_39182,N_39228);
xnor U39465 (N_39465,N_39020,N_39180);
nand U39466 (N_39466,N_39079,N_39151);
nor U39467 (N_39467,N_39225,N_39001);
xnor U39468 (N_39468,N_39158,N_39133);
or U39469 (N_39469,N_39188,N_39203);
nand U39470 (N_39470,N_39194,N_39014);
and U39471 (N_39471,N_39069,N_39167);
nor U39472 (N_39472,N_39131,N_39200);
or U39473 (N_39473,N_39123,N_39009);
or U39474 (N_39474,N_39043,N_39146);
xor U39475 (N_39475,N_39160,N_39107);
xor U39476 (N_39476,N_39218,N_39134);
nor U39477 (N_39477,N_39155,N_39051);
nand U39478 (N_39478,N_39036,N_39016);
nand U39479 (N_39479,N_39098,N_39245);
or U39480 (N_39480,N_39006,N_39249);
nand U39481 (N_39481,N_39114,N_39055);
or U39482 (N_39482,N_39183,N_39101);
nand U39483 (N_39483,N_39131,N_39030);
nor U39484 (N_39484,N_39088,N_39203);
xor U39485 (N_39485,N_39237,N_39027);
and U39486 (N_39486,N_39003,N_39217);
and U39487 (N_39487,N_39031,N_39158);
xnor U39488 (N_39488,N_39210,N_39211);
xnor U39489 (N_39489,N_39051,N_39027);
xor U39490 (N_39490,N_39072,N_39050);
and U39491 (N_39491,N_39212,N_39220);
nand U39492 (N_39492,N_39213,N_39132);
xor U39493 (N_39493,N_39214,N_39236);
nor U39494 (N_39494,N_39027,N_39164);
or U39495 (N_39495,N_39077,N_39212);
nor U39496 (N_39496,N_39085,N_39020);
nand U39497 (N_39497,N_39170,N_39099);
nand U39498 (N_39498,N_39240,N_39214);
xor U39499 (N_39499,N_39019,N_39010);
and U39500 (N_39500,N_39445,N_39350);
and U39501 (N_39501,N_39357,N_39296);
nand U39502 (N_39502,N_39390,N_39433);
xnor U39503 (N_39503,N_39345,N_39325);
xnor U39504 (N_39504,N_39275,N_39414);
and U39505 (N_39505,N_39475,N_39283);
xor U39506 (N_39506,N_39257,N_39294);
nand U39507 (N_39507,N_39463,N_39338);
and U39508 (N_39508,N_39467,N_39438);
or U39509 (N_39509,N_39457,N_39251);
or U39510 (N_39510,N_39453,N_39281);
or U39511 (N_39511,N_39388,N_39340);
nor U39512 (N_39512,N_39455,N_39363);
or U39513 (N_39513,N_39370,N_39497);
nor U39514 (N_39514,N_39479,N_39344);
nor U39515 (N_39515,N_39343,N_39323);
xnor U39516 (N_39516,N_39452,N_39304);
xnor U39517 (N_39517,N_39347,N_39321);
nand U39518 (N_39518,N_39472,N_39373);
xnor U39519 (N_39519,N_39368,N_39400);
xor U39520 (N_39520,N_39422,N_39282);
xor U39521 (N_39521,N_39466,N_39402);
nand U39522 (N_39522,N_39495,N_39428);
and U39523 (N_39523,N_39427,N_39425);
xor U39524 (N_39524,N_39393,N_39426);
xor U39525 (N_39525,N_39330,N_39374);
or U39526 (N_39526,N_39488,N_39332);
xnor U39527 (N_39527,N_39253,N_39461);
nand U39528 (N_39528,N_39310,N_39268);
or U39529 (N_39529,N_39386,N_39396);
nand U39530 (N_39530,N_39486,N_39334);
nand U39531 (N_39531,N_39287,N_39314);
xnor U39532 (N_39532,N_39348,N_39276);
xnor U39533 (N_39533,N_39311,N_39417);
nor U39534 (N_39534,N_39277,N_39489);
nor U39535 (N_39535,N_39420,N_39369);
nand U39536 (N_39536,N_39473,N_39492);
xor U39537 (N_39537,N_39476,N_39423);
nor U39538 (N_39538,N_39435,N_39270);
or U39539 (N_39539,N_39405,N_39432);
xor U39540 (N_39540,N_39273,N_39421);
xnor U39541 (N_39541,N_39477,N_39415);
and U39542 (N_39542,N_39434,N_39354);
or U39543 (N_39543,N_39447,N_39364);
nand U39544 (N_39544,N_39329,N_39383);
xnor U39545 (N_39545,N_39362,N_39441);
and U39546 (N_39546,N_39490,N_39485);
nor U39547 (N_39547,N_39279,N_39286);
nor U39548 (N_39548,N_39288,N_39301);
and U39549 (N_39549,N_39449,N_39424);
xor U39550 (N_39550,N_39436,N_39465);
nand U39551 (N_39551,N_39456,N_39250);
or U39552 (N_39552,N_39356,N_39307);
and U39553 (N_39553,N_39291,N_39265);
nand U39554 (N_39554,N_39437,N_39469);
and U39555 (N_39555,N_39316,N_39297);
or U39556 (N_39556,N_39353,N_39493);
or U39557 (N_39557,N_39439,N_39289);
nand U39558 (N_39558,N_39444,N_39255);
nor U39559 (N_39559,N_39322,N_39342);
nor U39560 (N_39560,N_39292,N_39351);
nor U39561 (N_39561,N_39413,N_39442);
xor U39562 (N_39562,N_39418,N_39339);
or U39563 (N_39563,N_39487,N_39318);
xor U39564 (N_39564,N_39337,N_39303);
xnor U39565 (N_39565,N_39254,N_39317);
nand U39566 (N_39566,N_39252,N_39468);
and U39567 (N_39567,N_39411,N_39355);
xnor U39568 (N_39568,N_39382,N_39459);
nand U39569 (N_39569,N_39358,N_39406);
nor U39570 (N_39570,N_39419,N_39407);
and U39571 (N_39571,N_39326,N_39259);
or U39572 (N_39572,N_39328,N_39494);
and U39573 (N_39573,N_39480,N_39284);
nand U39574 (N_39574,N_39462,N_39387);
and U39575 (N_39575,N_39367,N_39352);
and U39576 (N_39576,N_39446,N_39416);
nor U39577 (N_39577,N_39460,N_39258);
xnor U39578 (N_39578,N_39377,N_39450);
xor U39579 (N_39579,N_39482,N_39299);
xnor U39580 (N_39580,N_39272,N_39379);
and U39581 (N_39581,N_39371,N_39331);
and U39582 (N_39582,N_39431,N_39346);
or U39583 (N_39583,N_39341,N_39274);
and U39584 (N_39584,N_39359,N_39404);
xor U39585 (N_39585,N_39260,N_39305);
and U39586 (N_39586,N_39399,N_39327);
nor U39587 (N_39587,N_39380,N_39440);
or U39588 (N_39588,N_39271,N_39430);
nor U39589 (N_39589,N_39499,N_39483);
nor U39590 (N_39590,N_39484,N_39384);
nand U39591 (N_39591,N_39319,N_39448);
or U39592 (N_39592,N_39306,N_39451);
nand U39593 (N_39593,N_39464,N_39394);
nand U39594 (N_39594,N_39376,N_39295);
nor U39595 (N_39595,N_39333,N_39458);
nand U39596 (N_39596,N_39491,N_39410);
or U39597 (N_39597,N_39381,N_39408);
xnor U39598 (N_39598,N_39366,N_39269);
nand U39599 (N_39599,N_39349,N_39471);
or U39600 (N_39600,N_39290,N_39302);
nor U39601 (N_39601,N_39443,N_39267);
and U39602 (N_39602,N_39264,N_39365);
xnor U39603 (N_39603,N_39478,N_39256);
nand U39604 (N_39604,N_39395,N_39320);
xor U39605 (N_39605,N_39375,N_39263);
and U39606 (N_39606,N_39280,N_39498);
xnor U39607 (N_39607,N_39309,N_39285);
and U39608 (N_39608,N_39398,N_39315);
nand U39609 (N_39609,N_39403,N_39360);
nor U39610 (N_39610,N_39308,N_39361);
or U39611 (N_39611,N_39261,N_39481);
or U39612 (N_39612,N_39312,N_39324);
or U39613 (N_39613,N_39385,N_39454);
nand U39614 (N_39614,N_39300,N_39389);
or U39615 (N_39615,N_39266,N_39313);
and U39616 (N_39616,N_39298,N_39397);
nand U39617 (N_39617,N_39262,N_39372);
or U39618 (N_39618,N_39412,N_39392);
nand U39619 (N_39619,N_39429,N_39378);
and U39620 (N_39620,N_39391,N_39474);
and U39621 (N_39621,N_39336,N_39278);
and U39622 (N_39622,N_39401,N_39470);
nor U39623 (N_39623,N_39335,N_39293);
xnor U39624 (N_39624,N_39409,N_39496);
or U39625 (N_39625,N_39448,N_39280);
xnor U39626 (N_39626,N_39364,N_39288);
or U39627 (N_39627,N_39349,N_39467);
nand U39628 (N_39628,N_39464,N_39393);
and U39629 (N_39629,N_39400,N_39364);
nand U39630 (N_39630,N_39278,N_39326);
and U39631 (N_39631,N_39257,N_39277);
and U39632 (N_39632,N_39301,N_39487);
and U39633 (N_39633,N_39410,N_39483);
nand U39634 (N_39634,N_39321,N_39365);
or U39635 (N_39635,N_39460,N_39334);
and U39636 (N_39636,N_39327,N_39304);
xnor U39637 (N_39637,N_39493,N_39331);
and U39638 (N_39638,N_39277,N_39497);
or U39639 (N_39639,N_39428,N_39440);
nand U39640 (N_39640,N_39356,N_39349);
and U39641 (N_39641,N_39443,N_39318);
nor U39642 (N_39642,N_39414,N_39299);
or U39643 (N_39643,N_39261,N_39283);
nand U39644 (N_39644,N_39282,N_39379);
and U39645 (N_39645,N_39253,N_39459);
and U39646 (N_39646,N_39419,N_39441);
nand U39647 (N_39647,N_39280,N_39397);
nor U39648 (N_39648,N_39427,N_39435);
xor U39649 (N_39649,N_39438,N_39344);
and U39650 (N_39650,N_39297,N_39386);
xor U39651 (N_39651,N_39421,N_39451);
or U39652 (N_39652,N_39324,N_39351);
and U39653 (N_39653,N_39353,N_39377);
and U39654 (N_39654,N_39367,N_39385);
nand U39655 (N_39655,N_39467,N_39477);
or U39656 (N_39656,N_39397,N_39262);
and U39657 (N_39657,N_39379,N_39403);
nand U39658 (N_39658,N_39490,N_39372);
or U39659 (N_39659,N_39460,N_39359);
or U39660 (N_39660,N_39325,N_39327);
or U39661 (N_39661,N_39281,N_39377);
nand U39662 (N_39662,N_39416,N_39268);
nand U39663 (N_39663,N_39312,N_39286);
xor U39664 (N_39664,N_39482,N_39348);
nor U39665 (N_39665,N_39318,N_39305);
xnor U39666 (N_39666,N_39490,N_39332);
and U39667 (N_39667,N_39481,N_39412);
xnor U39668 (N_39668,N_39471,N_39436);
nand U39669 (N_39669,N_39415,N_39431);
xor U39670 (N_39670,N_39451,N_39477);
nor U39671 (N_39671,N_39387,N_39392);
nand U39672 (N_39672,N_39426,N_39407);
or U39673 (N_39673,N_39422,N_39440);
xor U39674 (N_39674,N_39454,N_39448);
or U39675 (N_39675,N_39270,N_39496);
and U39676 (N_39676,N_39404,N_39482);
nand U39677 (N_39677,N_39460,N_39325);
and U39678 (N_39678,N_39452,N_39360);
and U39679 (N_39679,N_39456,N_39367);
nand U39680 (N_39680,N_39257,N_39493);
xor U39681 (N_39681,N_39250,N_39288);
xor U39682 (N_39682,N_39427,N_39344);
or U39683 (N_39683,N_39390,N_39404);
nor U39684 (N_39684,N_39434,N_39461);
and U39685 (N_39685,N_39344,N_39290);
xnor U39686 (N_39686,N_39465,N_39264);
or U39687 (N_39687,N_39332,N_39442);
nand U39688 (N_39688,N_39402,N_39304);
nand U39689 (N_39689,N_39472,N_39490);
nor U39690 (N_39690,N_39480,N_39297);
xor U39691 (N_39691,N_39485,N_39489);
nand U39692 (N_39692,N_39479,N_39451);
nand U39693 (N_39693,N_39278,N_39311);
or U39694 (N_39694,N_39262,N_39277);
xnor U39695 (N_39695,N_39335,N_39295);
nand U39696 (N_39696,N_39490,N_39253);
nand U39697 (N_39697,N_39322,N_39471);
and U39698 (N_39698,N_39282,N_39294);
and U39699 (N_39699,N_39485,N_39310);
nand U39700 (N_39700,N_39478,N_39292);
xnor U39701 (N_39701,N_39425,N_39302);
or U39702 (N_39702,N_39279,N_39312);
nand U39703 (N_39703,N_39398,N_39261);
and U39704 (N_39704,N_39422,N_39345);
nand U39705 (N_39705,N_39452,N_39488);
nor U39706 (N_39706,N_39489,N_39346);
and U39707 (N_39707,N_39327,N_39494);
nor U39708 (N_39708,N_39259,N_39352);
nand U39709 (N_39709,N_39284,N_39285);
nor U39710 (N_39710,N_39269,N_39270);
nand U39711 (N_39711,N_39346,N_39268);
nor U39712 (N_39712,N_39270,N_39258);
and U39713 (N_39713,N_39370,N_39277);
and U39714 (N_39714,N_39494,N_39297);
nand U39715 (N_39715,N_39272,N_39382);
nor U39716 (N_39716,N_39335,N_39296);
nor U39717 (N_39717,N_39378,N_39358);
nand U39718 (N_39718,N_39492,N_39477);
xnor U39719 (N_39719,N_39360,N_39250);
and U39720 (N_39720,N_39250,N_39493);
nand U39721 (N_39721,N_39282,N_39341);
nand U39722 (N_39722,N_39485,N_39402);
nand U39723 (N_39723,N_39457,N_39288);
xnor U39724 (N_39724,N_39353,N_39375);
nor U39725 (N_39725,N_39284,N_39389);
xor U39726 (N_39726,N_39395,N_39411);
nand U39727 (N_39727,N_39387,N_39468);
nand U39728 (N_39728,N_39332,N_39328);
nand U39729 (N_39729,N_39410,N_39437);
nor U39730 (N_39730,N_39302,N_39376);
xnor U39731 (N_39731,N_39252,N_39284);
and U39732 (N_39732,N_39384,N_39366);
and U39733 (N_39733,N_39317,N_39379);
xor U39734 (N_39734,N_39346,N_39342);
xnor U39735 (N_39735,N_39451,N_39355);
nor U39736 (N_39736,N_39392,N_39360);
nor U39737 (N_39737,N_39424,N_39257);
or U39738 (N_39738,N_39474,N_39493);
and U39739 (N_39739,N_39443,N_39478);
xor U39740 (N_39740,N_39478,N_39277);
or U39741 (N_39741,N_39290,N_39365);
nand U39742 (N_39742,N_39465,N_39296);
nand U39743 (N_39743,N_39280,N_39493);
or U39744 (N_39744,N_39357,N_39495);
and U39745 (N_39745,N_39409,N_39292);
nor U39746 (N_39746,N_39460,N_39371);
xnor U39747 (N_39747,N_39354,N_39387);
nor U39748 (N_39748,N_39258,N_39404);
or U39749 (N_39749,N_39441,N_39313);
or U39750 (N_39750,N_39664,N_39687);
nand U39751 (N_39751,N_39584,N_39728);
and U39752 (N_39752,N_39669,N_39749);
nand U39753 (N_39753,N_39685,N_39707);
or U39754 (N_39754,N_39681,N_39671);
and U39755 (N_39755,N_39635,N_39550);
and U39756 (N_39756,N_39587,N_39535);
nor U39757 (N_39757,N_39553,N_39693);
nand U39758 (N_39758,N_39588,N_39565);
nand U39759 (N_39759,N_39708,N_39609);
nand U39760 (N_39760,N_39725,N_39744);
nand U39761 (N_39761,N_39627,N_39651);
or U39762 (N_39762,N_39697,N_39520);
nand U39763 (N_39763,N_39726,N_39604);
and U39764 (N_39764,N_39714,N_39544);
and U39765 (N_39765,N_39735,N_39607);
or U39766 (N_39766,N_39619,N_39505);
and U39767 (N_39767,N_39716,N_39524);
nor U39768 (N_39768,N_39721,N_39519);
xor U39769 (N_39769,N_39545,N_39736);
and U39770 (N_39770,N_39624,N_39642);
and U39771 (N_39771,N_39608,N_39733);
or U39772 (N_39772,N_39576,N_39741);
or U39773 (N_39773,N_39622,N_39577);
nor U39774 (N_39774,N_39591,N_39515);
nand U39775 (N_39775,N_39719,N_39711);
and U39776 (N_39776,N_39720,N_39652);
nor U39777 (N_39777,N_39746,N_39675);
or U39778 (N_39778,N_39504,N_39743);
or U39779 (N_39779,N_39617,N_39657);
and U39780 (N_39780,N_39580,N_39598);
nand U39781 (N_39781,N_39512,N_39648);
or U39782 (N_39782,N_39632,N_39602);
xnor U39783 (N_39783,N_39742,N_39713);
and U39784 (N_39784,N_39636,N_39562);
nor U39785 (N_39785,N_39674,N_39528);
nor U39786 (N_39786,N_39601,N_39501);
or U39787 (N_39787,N_39715,N_39666);
nor U39788 (N_39788,N_39586,N_39611);
xnor U39789 (N_39789,N_39639,N_39668);
nor U39790 (N_39790,N_39731,N_39696);
nor U39791 (N_39791,N_39730,N_39634);
nand U39792 (N_39792,N_39556,N_39626);
or U39793 (N_39793,N_39558,N_39594);
nor U39794 (N_39794,N_39667,N_39575);
and U39795 (N_39795,N_39738,N_39518);
and U39796 (N_39796,N_39637,N_39739);
xnor U39797 (N_39797,N_39747,N_39542);
nand U39798 (N_39798,N_39699,N_39691);
and U39799 (N_39799,N_39514,N_39623);
nor U39800 (N_39800,N_39507,N_39698);
nor U39801 (N_39801,N_39682,N_39557);
or U39802 (N_39802,N_39672,N_39539);
or U39803 (N_39803,N_39676,N_39548);
and U39804 (N_39804,N_39621,N_39703);
nor U39805 (N_39805,N_39571,N_39560);
nand U39806 (N_39806,N_39543,N_39678);
or U39807 (N_39807,N_39516,N_39748);
or U39808 (N_39808,N_39702,N_39585);
or U39809 (N_39809,N_39701,N_39597);
xor U39810 (N_39810,N_39649,N_39547);
or U39811 (N_39811,N_39663,N_39660);
xnor U39812 (N_39812,N_39517,N_39616);
or U39813 (N_39813,N_39551,N_39723);
or U39814 (N_39814,N_39554,N_39628);
xor U39815 (N_39815,N_39724,N_39521);
nor U39816 (N_39816,N_39559,N_39629);
xor U39817 (N_39817,N_39700,N_39717);
or U39818 (N_39818,N_39612,N_39508);
xor U39819 (N_39819,N_39658,N_39677);
xor U39820 (N_39820,N_39643,N_39683);
or U39821 (N_39821,N_39572,N_39710);
and U39822 (N_39822,N_39606,N_39527);
nand U39823 (N_39823,N_39536,N_39570);
or U39824 (N_39824,N_39523,N_39582);
and U39825 (N_39825,N_39613,N_39509);
and U39826 (N_39826,N_39589,N_39537);
or U39827 (N_39827,N_39541,N_39618);
xnor U39828 (N_39828,N_39670,N_39532);
xor U39829 (N_39829,N_39630,N_39500);
and U39830 (N_39830,N_39625,N_39530);
nand U39831 (N_39831,N_39689,N_39640);
nand U39832 (N_39832,N_39641,N_39593);
xor U39833 (N_39833,N_39680,N_39727);
nand U39834 (N_39834,N_39647,N_39511);
or U39835 (N_39835,N_39526,N_39561);
nor U39836 (N_39836,N_39583,N_39600);
nand U39837 (N_39837,N_39605,N_39734);
nor U39838 (N_39838,N_39656,N_39610);
nand U39839 (N_39839,N_39704,N_39581);
nand U39840 (N_39840,N_39705,N_39638);
or U39841 (N_39841,N_39568,N_39614);
and U39842 (N_39842,N_39662,N_39534);
nor U39843 (N_39843,N_39540,N_39603);
and U39844 (N_39844,N_39574,N_39522);
or U39845 (N_39845,N_39695,N_39592);
nor U39846 (N_39846,N_39549,N_39564);
xnor U39847 (N_39847,N_39688,N_39538);
xnor U39848 (N_39848,N_39665,N_39631);
nand U39849 (N_39849,N_39555,N_39737);
nor U39850 (N_39850,N_39654,N_39531);
nor U39851 (N_39851,N_39567,N_39694);
nor U39852 (N_39852,N_39645,N_39513);
nor U39853 (N_39853,N_39644,N_39633);
or U39854 (N_39854,N_39740,N_39563);
xnor U39855 (N_39855,N_39653,N_39546);
xnor U39856 (N_39856,N_39690,N_39732);
nand U39857 (N_39857,N_39533,N_39525);
nand U39858 (N_39858,N_39599,N_39659);
xor U39859 (N_39859,N_39679,N_39590);
xor U39860 (N_39860,N_39569,N_39729);
xor U39861 (N_39861,N_39646,N_39673);
xnor U39862 (N_39862,N_39661,N_39718);
or U39863 (N_39863,N_39502,N_39706);
xor U39864 (N_39864,N_39579,N_39709);
nor U39865 (N_39865,N_39620,N_39595);
nand U39866 (N_39866,N_39722,N_39684);
or U39867 (N_39867,N_39552,N_39655);
xor U39868 (N_39868,N_39573,N_39578);
xor U39869 (N_39869,N_39745,N_39650);
nor U39870 (N_39870,N_39566,N_39686);
xnor U39871 (N_39871,N_39529,N_39692);
and U39872 (N_39872,N_39615,N_39596);
xor U39873 (N_39873,N_39712,N_39503);
xor U39874 (N_39874,N_39506,N_39510);
nor U39875 (N_39875,N_39689,N_39712);
or U39876 (N_39876,N_39729,N_39657);
nand U39877 (N_39877,N_39734,N_39728);
xnor U39878 (N_39878,N_39692,N_39696);
or U39879 (N_39879,N_39584,N_39689);
nor U39880 (N_39880,N_39666,N_39559);
xnor U39881 (N_39881,N_39621,N_39570);
nor U39882 (N_39882,N_39541,N_39652);
or U39883 (N_39883,N_39606,N_39737);
or U39884 (N_39884,N_39570,N_39644);
nand U39885 (N_39885,N_39692,N_39590);
or U39886 (N_39886,N_39592,N_39655);
nand U39887 (N_39887,N_39555,N_39512);
nor U39888 (N_39888,N_39651,N_39719);
xor U39889 (N_39889,N_39688,N_39506);
and U39890 (N_39890,N_39727,N_39521);
or U39891 (N_39891,N_39580,N_39689);
nand U39892 (N_39892,N_39717,N_39632);
xnor U39893 (N_39893,N_39676,N_39537);
xor U39894 (N_39894,N_39539,N_39724);
nand U39895 (N_39895,N_39547,N_39521);
and U39896 (N_39896,N_39696,N_39740);
nor U39897 (N_39897,N_39700,N_39716);
and U39898 (N_39898,N_39603,N_39502);
or U39899 (N_39899,N_39512,N_39504);
and U39900 (N_39900,N_39575,N_39694);
nor U39901 (N_39901,N_39651,N_39559);
or U39902 (N_39902,N_39713,N_39725);
nor U39903 (N_39903,N_39558,N_39658);
xor U39904 (N_39904,N_39600,N_39640);
nor U39905 (N_39905,N_39703,N_39513);
nor U39906 (N_39906,N_39558,N_39571);
and U39907 (N_39907,N_39697,N_39555);
nand U39908 (N_39908,N_39602,N_39742);
nor U39909 (N_39909,N_39669,N_39746);
and U39910 (N_39910,N_39536,N_39595);
or U39911 (N_39911,N_39658,N_39552);
nand U39912 (N_39912,N_39555,N_39746);
xnor U39913 (N_39913,N_39742,N_39518);
or U39914 (N_39914,N_39686,N_39606);
nand U39915 (N_39915,N_39654,N_39745);
or U39916 (N_39916,N_39526,N_39618);
or U39917 (N_39917,N_39667,N_39587);
nor U39918 (N_39918,N_39700,N_39696);
xor U39919 (N_39919,N_39529,N_39654);
and U39920 (N_39920,N_39513,N_39619);
and U39921 (N_39921,N_39677,N_39514);
or U39922 (N_39922,N_39515,N_39520);
nand U39923 (N_39923,N_39603,N_39710);
or U39924 (N_39924,N_39706,N_39505);
nor U39925 (N_39925,N_39617,N_39547);
nand U39926 (N_39926,N_39665,N_39709);
nand U39927 (N_39927,N_39503,N_39551);
xnor U39928 (N_39928,N_39725,N_39508);
xor U39929 (N_39929,N_39721,N_39528);
or U39930 (N_39930,N_39734,N_39706);
nand U39931 (N_39931,N_39619,N_39727);
xor U39932 (N_39932,N_39553,N_39624);
and U39933 (N_39933,N_39720,N_39602);
nand U39934 (N_39934,N_39572,N_39590);
nor U39935 (N_39935,N_39570,N_39529);
nor U39936 (N_39936,N_39552,N_39585);
nor U39937 (N_39937,N_39697,N_39613);
nand U39938 (N_39938,N_39522,N_39575);
and U39939 (N_39939,N_39684,N_39674);
and U39940 (N_39940,N_39721,N_39736);
or U39941 (N_39941,N_39648,N_39641);
and U39942 (N_39942,N_39725,N_39685);
nand U39943 (N_39943,N_39688,N_39711);
nor U39944 (N_39944,N_39722,N_39635);
or U39945 (N_39945,N_39669,N_39595);
xnor U39946 (N_39946,N_39618,N_39581);
nor U39947 (N_39947,N_39610,N_39712);
nand U39948 (N_39948,N_39674,N_39630);
or U39949 (N_39949,N_39612,N_39685);
xnor U39950 (N_39950,N_39629,N_39596);
and U39951 (N_39951,N_39576,N_39626);
or U39952 (N_39952,N_39729,N_39627);
nand U39953 (N_39953,N_39740,N_39581);
nor U39954 (N_39954,N_39699,N_39578);
nand U39955 (N_39955,N_39612,N_39515);
xor U39956 (N_39956,N_39623,N_39642);
nor U39957 (N_39957,N_39715,N_39649);
nand U39958 (N_39958,N_39527,N_39607);
or U39959 (N_39959,N_39745,N_39707);
nor U39960 (N_39960,N_39534,N_39626);
nand U39961 (N_39961,N_39530,N_39687);
nand U39962 (N_39962,N_39683,N_39730);
nor U39963 (N_39963,N_39516,N_39624);
xnor U39964 (N_39964,N_39508,N_39668);
nor U39965 (N_39965,N_39700,N_39582);
nand U39966 (N_39966,N_39613,N_39601);
and U39967 (N_39967,N_39609,N_39748);
nor U39968 (N_39968,N_39698,N_39702);
xor U39969 (N_39969,N_39727,N_39621);
xnor U39970 (N_39970,N_39502,N_39730);
or U39971 (N_39971,N_39544,N_39561);
and U39972 (N_39972,N_39612,N_39577);
xor U39973 (N_39973,N_39580,N_39538);
nand U39974 (N_39974,N_39510,N_39748);
or U39975 (N_39975,N_39524,N_39661);
nor U39976 (N_39976,N_39693,N_39580);
nor U39977 (N_39977,N_39587,N_39743);
nor U39978 (N_39978,N_39632,N_39572);
nand U39979 (N_39979,N_39513,N_39734);
nand U39980 (N_39980,N_39647,N_39702);
and U39981 (N_39981,N_39523,N_39718);
and U39982 (N_39982,N_39615,N_39716);
nand U39983 (N_39983,N_39749,N_39525);
nand U39984 (N_39984,N_39604,N_39639);
or U39985 (N_39985,N_39510,N_39708);
nand U39986 (N_39986,N_39560,N_39610);
nor U39987 (N_39987,N_39707,N_39662);
or U39988 (N_39988,N_39672,N_39635);
nor U39989 (N_39989,N_39630,N_39513);
or U39990 (N_39990,N_39664,N_39720);
or U39991 (N_39991,N_39539,N_39679);
xor U39992 (N_39992,N_39555,N_39690);
and U39993 (N_39993,N_39737,N_39543);
nand U39994 (N_39994,N_39637,N_39581);
xnor U39995 (N_39995,N_39740,N_39710);
xor U39996 (N_39996,N_39707,N_39666);
nor U39997 (N_39997,N_39577,N_39566);
nor U39998 (N_39998,N_39636,N_39717);
and U39999 (N_39999,N_39729,N_39572);
nor U40000 (N_40000,N_39804,N_39998);
or U40001 (N_40001,N_39858,N_39863);
nor U40002 (N_40002,N_39835,N_39794);
xnor U40003 (N_40003,N_39938,N_39844);
or U40004 (N_40004,N_39876,N_39812);
or U40005 (N_40005,N_39781,N_39855);
nand U40006 (N_40006,N_39929,N_39920);
xor U40007 (N_40007,N_39934,N_39931);
nor U40008 (N_40008,N_39915,N_39923);
xnor U40009 (N_40009,N_39788,N_39853);
nand U40010 (N_40010,N_39902,N_39914);
or U40011 (N_40011,N_39895,N_39912);
nand U40012 (N_40012,N_39966,N_39972);
and U40013 (N_40013,N_39963,N_39901);
xnor U40014 (N_40014,N_39764,N_39766);
nand U40015 (N_40015,N_39899,N_39866);
or U40016 (N_40016,N_39954,N_39905);
nor U40017 (N_40017,N_39860,N_39988);
and U40018 (N_40018,N_39878,N_39843);
nor U40019 (N_40019,N_39841,N_39758);
and U40020 (N_40020,N_39879,N_39810);
nand U40021 (N_40021,N_39777,N_39933);
and U40022 (N_40022,N_39943,N_39785);
nand U40023 (N_40023,N_39979,N_39936);
nand U40024 (N_40024,N_39891,N_39778);
nor U40025 (N_40025,N_39942,N_39865);
or U40026 (N_40026,N_39977,N_39859);
xnor U40027 (N_40027,N_39753,N_39969);
xor U40028 (N_40028,N_39884,N_39754);
nand U40029 (N_40029,N_39842,N_39837);
nor U40030 (N_40030,N_39997,N_39930);
or U40031 (N_40031,N_39981,N_39751);
or U40032 (N_40032,N_39992,N_39763);
or U40033 (N_40033,N_39984,N_39965);
nor U40034 (N_40034,N_39824,N_39765);
xor U40035 (N_40035,N_39845,N_39802);
or U40036 (N_40036,N_39761,N_39838);
nor U40037 (N_40037,N_39820,N_39769);
or U40038 (N_40038,N_39839,N_39791);
nor U40039 (N_40039,N_39955,N_39871);
and U40040 (N_40040,N_39830,N_39919);
nor U40041 (N_40041,N_39803,N_39913);
and U40042 (N_40042,N_39953,N_39962);
or U40043 (N_40043,N_39868,N_39896);
xor U40044 (N_40044,N_39944,N_39909);
nor U40045 (N_40045,N_39989,N_39809);
or U40046 (N_40046,N_39872,N_39806);
nor U40047 (N_40047,N_39925,N_39922);
xnor U40048 (N_40048,N_39819,N_39946);
and U40049 (N_40049,N_39889,N_39873);
nand U40050 (N_40050,N_39772,N_39993);
nor U40051 (N_40051,N_39924,N_39883);
nor U40052 (N_40052,N_39957,N_39921);
and U40053 (N_40053,N_39789,N_39795);
nand U40054 (N_40054,N_39894,N_39950);
and U40055 (N_40055,N_39826,N_39770);
and U40056 (N_40056,N_39910,N_39831);
or U40057 (N_40057,N_39877,N_39976);
and U40058 (N_40058,N_39825,N_39968);
xnor U40059 (N_40059,N_39864,N_39857);
nor U40060 (N_40060,N_39980,N_39932);
xnor U40061 (N_40061,N_39983,N_39828);
nor U40062 (N_40062,N_39827,N_39780);
or U40063 (N_40063,N_39900,N_39911);
nor U40064 (N_40064,N_39834,N_39974);
nor U40065 (N_40065,N_39886,N_39869);
nand U40066 (N_40066,N_39773,N_39898);
nor U40067 (N_40067,N_39903,N_39790);
nand U40068 (N_40068,N_39948,N_39862);
and U40069 (N_40069,N_39850,N_39750);
or U40070 (N_40070,N_39767,N_39907);
nand U40071 (N_40071,N_39951,N_39964);
and U40072 (N_40072,N_39796,N_39818);
nand U40073 (N_40073,N_39973,N_39755);
and U40074 (N_40074,N_39756,N_39823);
nand U40075 (N_40075,N_39958,N_39771);
or U40076 (N_40076,N_39822,N_39851);
xor U40077 (N_40077,N_39945,N_39959);
nor U40078 (N_40078,N_39941,N_39840);
or U40079 (N_40079,N_39996,N_39890);
and U40080 (N_40080,N_39787,N_39779);
and U40081 (N_40081,N_39971,N_39757);
and U40082 (N_40082,N_39885,N_39939);
or U40083 (N_40083,N_39817,N_39990);
or U40084 (N_40084,N_39978,N_39892);
xor U40085 (N_40085,N_39800,N_39882);
nor U40086 (N_40086,N_39982,N_39906);
or U40087 (N_40087,N_39897,N_39881);
nand U40088 (N_40088,N_39816,N_39867);
or U40089 (N_40089,N_39861,N_39782);
nor U40090 (N_40090,N_39995,N_39798);
xor U40091 (N_40091,N_39813,N_39784);
nand U40092 (N_40092,N_39847,N_39887);
and U40093 (N_40093,N_39832,N_39870);
nor U40094 (N_40094,N_39893,N_39985);
or U40095 (N_40095,N_39852,N_39807);
xor U40096 (N_40096,N_39760,N_39854);
xor U40097 (N_40097,N_39792,N_39952);
and U40098 (N_40098,N_39829,N_39799);
and U40099 (N_40099,N_39947,N_39833);
nand U40100 (N_40100,N_39940,N_39811);
xor U40101 (N_40101,N_39975,N_39797);
or U40102 (N_40102,N_39918,N_39880);
nor U40103 (N_40103,N_39991,N_39875);
or U40104 (N_40104,N_39908,N_39849);
nand U40105 (N_40105,N_39956,N_39916);
nor U40106 (N_40106,N_39821,N_39949);
and U40107 (N_40107,N_39848,N_39994);
nor U40108 (N_40108,N_39776,N_39762);
nand U40109 (N_40109,N_39752,N_39935);
nand U40110 (N_40110,N_39986,N_39856);
xor U40111 (N_40111,N_39814,N_39846);
nand U40112 (N_40112,N_39888,N_39774);
and U40113 (N_40113,N_39960,N_39793);
nor U40114 (N_40114,N_39815,N_39927);
nand U40115 (N_40115,N_39928,N_39801);
nand U40116 (N_40116,N_39926,N_39961);
nand U40117 (N_40117,N_39874,N_39970);
xnor U40118 (N_40118,N_39783,N_39808);
nor U40119 (N_40119,N_39768,N_39967);
or U40120 (N_40120,N_39805,N_39775);
nor U40121 (N_40121,N_39999,N_39987);
xor U40122 (N_40122,N_39836,N_39937);
or U40123 (N_40123,N_39786,N_39917);
nor U40124 (N_40124,N_39904,N_39759);
nand U40125 (N_40125,N_39842,N_39947);
xor U40126 (N_40126,N_39955,N_39999);
nor U40127 (N_40127,N_39936,N_39992);
nand U40128 (N_40128,N_39794,N_39879);
and U40129 (N_40129,N_39830,N_39778);
or U40130 (N_40130,N_39761,N_39867);
xor U40131 (N_40131,N_39897,N_39977);
xnor U40132 (N_40132,N_39922,N_39980);
xor U40133 (N_40133,N_39927,N_39990);
nand U40134 (N_40134,N_39802,N_39868);
or U40135 (N_40135,N_39857,N_39768);
nor U40136 (N_40136,N_39817,N_39759);
nand U40137 (N_40137,N_39877,N_39766);
nand U40138 (N_40138,N_39890,N_39821);
xnor U40139 (N_40139,N_39900,N_39886);
or U40140 (N_40140,N_39805,N_39833);
xnor U40141 (N_40141,N_39750,N_39949);
nor U40142 (N_40142,N_39883,N_39753);
nor U40143 (N_40143,N_39974,N_39804);
or U40144 (N_40144,N_39981,N_39788);
and U40145 (N_40145,N_39798,N_39998);
or U40146 (N_40146,N_39864,N_39899);
or U40147 (N_40147,N_39944,N_39769);
nand U40148 (N_40148,N_39986,N_39793);
and U40149 (N_40149,N_39753,N_39889);
nand U40150 (N_40150,N_39904,N_39779);
nand U40151 (N_40151,N_39845,N_39877);
nand U40152 (N_40152,N_39914,N_39887);
nand U40153 (N_40153,N_39954,N_39800);
xor U40154 (N_40154,N_39924,N_39818);
nand U40155 (N_40155,N_39981,N_39807);
or U40156 (N_40156,N_39768,N_39953);
or U40157 (N_40157,N_39768,N_39987);
or U40158 (N_40158,N_39912,N_39928);
nor U40159 (N_40159,N_39951,N_39807);
xnor U40160 (N_40160,N_39813,N_39824);
nand U40161 (N_40161,N_39798,N_39793);
nor U40162 (N_40162,N_39842,N_39927);
nor U40163 (N_40163,N_39891,N_39957);
nand U40164 (N_40164,N_39884,N_39848);
nor U40165 (N_40165,N_39750,N_39871);
xnor U40166 (N_40166,N_39973,N_39838);
and U40167 (N_40167,N_39848,N_39926);
or U40168 (N_40168,N_39979,N_39993);
or U40169 (N_40169,N_39878,N_39918);
nand U40170 (N_40170,N_39807,N_39763);
xor U40171 (N_40171,N_39844,N_39949);
or U40172 (N_40172,N_39998,N_39758);
nand U40173 (N_40173,N_39961,N_39908);
nor U40174 (N_40174,N_39908,N_39958);
nand U40175 (N_40175,N_39981,N_39841);
nor U40176 (N_40176,N_39917,N_39999);
nand U40177 (N_40177,N_39981,N_39845);
xor U40178 (N_40178,N_39785,N_39895);
or U40179 (N_40179,N_39844,N_39941);
or U40180 (N_40180,N_39980,N_39850);
and U40181 (N_40181,N_39881,N_39997);
or U40182 (N_40182,N_39870,N_39858);
nand U40183 (N_40183,N_39973,N_39952);
nand U40184 (N_40184,N_39803,N_39958);
xnor U40185 (N_40185,N_39909,N_39987);
or U40186 (N_40186,N_39772,N_39765);
xor U40187 (N_40187,N_39858,N_39894);
and U40188 (N_40188,N_39930,N_39769);
and U40189 (N_40189,N_39795,N_39956);
or U40190 (N_40190,N_39885,N_39919);
xnor U40191 (N_40191,N_39775,N_39830);
xor U40192 (N_40192,N_39922,N_39942);
and U40193 (N_40193,N_39935,N_39805);
or U40194 (N_40194,N_39981,N_39934);
nor U40195 (N_40195,N_39893,N_39814);
nand U40196 (N_40196,N_39764,N_39933);
and U40197 (N_40197,N_39944,N_39752);
xnor U40198 (N_40198,N_39855,N_39751);
xor U40199 (N_40199,N_39984,N_39859);
or U40200 (N_40200,N_39888,N_39921);
nand U40201 (N_40201,N_39958,N_39918);
or U40202 (N_40202,N_39790,N_39820);
nor U40203 (N_40203,N_39884,N_39951);
and U40204 (N_40204,N_39811,N_39893);
or U40205 (N_40205,N_39923,N_39860);
and U40206 (N_40206,N_39945,N_39855);
or U40207 (N_40207,N_39795,N_39751);
nand U40208 (N_40208,N_39969,N_39909);
nand U40209 (N_40209,N_39915,N_39841);
xnor U40210 (N_40210,N_39908,N_39970);
nand U40211 (N_40211,N_39877,N_39811);
xor U40212 (N_40212,N_39937,N_39979);
nand U40213 (N_40213,N_39919,N_39921);
nor U40214 (N_40214,N_39890,N_39880);
nor U40215 (N_40215,N_39951,N_39799);
or U40216 (N_40216,N_39796,N_39879);
nand U40217 (N_40217,N_39946,N_39906);
nor U40218 (N_40218,N_39935,N_39914);
xor U40219 (N_40219,N_39964,N_39992);
xnor U40220 (N_40220,N_39993,N_39880);
nand U40221 (N_40221,N_39866,N_39799);
nor U40222 (N_40222,N_39997,N_39956);
nor U40223 (N_40223,N_39839,N_39956);
nor U40224 (N_40224,N_39814,N_39972);
or U40225 (N_40225,N_39956,N_39954);
nor U40226 (N_40226,N_39829,N_39866);
nand U40227 (N_40227,N_39835,N_39864);
nor U40228 (N_40228,N_39885,N_39865);
nor U40229 (N_40229,N_39752,N_39821);
and U40230 (N_40230,N_39859,N_39781);
nand U40231 (N_40231,N_39853,N_39753);
xor U40232 (N_40232,N_39753,N_39780);
and U40233 (N_40233,N_39779,N_39913);
and U40234 (N_40234,N_39944,N_39816);
xnor U40235 (N_40235,N_39904,N_39946);
xnor U40236 (N_40236,N_39995,N_39858);
nor U40237 (N_40237,N_39924,N_39911);
nor U40238 (N_40238,N_39951,N_39809);
or U40239 (N_40239,N_39785,N_39992);
nor U40240 (N_40240,N_39867,N_39750);
xnor U40241 (N_40241,N_39790,N_39772);
and U40242 (N_40242,N_39885,N_39813);
nand U40243 (N_40243,N_39983,N_39980);
or U40244 (N_40244,N_39906,N_39847);
xor U40245 (N_40245,N_39819,N_39771);
nand U40246 (N_40246,N_39890,N_39820);
or U40247 (N_40247,N_39916,N_39919);
xnor U40248 (N_40248,N_39921,N_39807);
or U40249 (N_40249,N_39940,N_39981);
nor U40250 (N_40250,N_40110,N_40223);
or U40251 (N_40251,N_40021,N_40192);
and U40252 (N_40252,N_40219,N_40133);
nor U40253 (N_40253,N_40126,N_40097);
xnor U40254 (N_40254,N_40202,N_40165);
nor U40255 (N_40255,N_40161,N_40213);
xor U40256 (N_40256,N_40002,N_40237);
or U40257 (N_40257,N_40047,N_40184);
xor U40258 (N_40258,N_40150,N_40052);
or U40259 (N_40259,N_40107,N_40131);
and U40260 (N_40260,N_40101,N_40123);
xor U40261 (N_40261,N_40030,N_40036);
and U40262 (N_40262,N_40244,N_40146);
nor U40263 (N_40263,N_40095,N_40092);
nor U40264 (N_40264,N_40201,N_40157);
nand U40265 (N_40265,N_40164,N_40182);
xnor U40266 (N_40266,N_40240,N_40027);
nor U40267 (N_40267,N_40194,N_40087);
xor U40268 (N_40268,N_40246,N_40198);
and U40269 (N_40269,N_40100,N_40112);
or U40270 (N_40270,N_40230,N_40153);
or U40271 (N_40271,N_40159,N_40069);
nand U40272 (N_40272,N_40111,N_40050);
xnor U40273 (N_40273,N_40235,N_40233);
nand U40274 (N_40274,N_40227,N_40022);
nand U40275 (N_40275,N_40175,N_40135);
and U40276 (N_40276,N_40200,N_40248);
and U40277 (N_40277,N_40044,N_40168);
xor U40278 (N_40278,N_40177,N_40073);
nand U40279 (N_40279,N_40071,N_40207);
and U40280 (N_40280,N_40006,N_40234);
or U40281 (N_40281,N_40221,N_40118);
xor U40282 (N_40282,N_40004,N_40013);
xor U40283 (N_40283,N_40063,N_40141);
xnor U40284 (N_40284,N_40224,N_40045);
and U40285 (N_40285,N_40080,N_40122);
xnor U40286 (N_40286,N_40205,N_40025);
or U40287 (N_40287,N_40190,N_40086);
xnor U40288 (N_40288,N_40149,N_40232);
nor U40289 (N_40289,N_40003,N_40243);
or U40290 (N_40290,N_40059,N_40019);
xor U40291 (N_40291,N_40132,N_40093);
nor U40292 (N_40292,N_40226,N_40145);
nor U40293 (N_40293,N_40186,N_40139);
xor U40294 (N_40294,N_40204,N_40058);
nand U40295 (N_40295,N_40225,N_40179);
nor U40296 (N_40296,N_40077,N_40053);
and U40297 (N_40297,N_40136,N_40166);
nand U40298 (N_40298,N_40148,N_40178);
nor U40299 (N_40299,N_40151,N_40117);
xnor U40300 (N_40300,N_40172,N_40064);
and U40301 (N_40301,N_40158,N_40040);
or U40302 (N_40302,N_40137,N_40075);
or U40303 (N_40303,N_40090,N_40127);
nor U40304 (N_40304,N_40031,N_40241);
nand U40305 (N_40305,N_40079,N_40147);
nand U40306 (N_40306,N_40191,N_40152);
nand U40307 (N_40307,N_40067,N_40007);
nor U40308 (N_40308,N_40009,N_40169);
nand U40309 (N_40309,N_40104,N_40188);
nand U40310 (N_40310,N_40099,N_40010);
and U40311 (N_40311,N_40035,N_40160);
nand U40312 (N_40312,N_40109,N_40038);
and U40313 (N_40313,N_40231,N_40162);
nor U40314 (N_40314,N_40245,N_40054);
nand U40315 (N_40315,N_40134,N_40084);
xor U40316 (N_40316,N_40039,N_40018);
xor U40317 (N_40317,N_40026,N_40222);
and U40318 (N_40318,N_40094,N_40051);
nand U40319 (N_40319,N_40041,N_40074);
nor U40320 (N_40320,N_40203,N_40116);
nor U40321 (N_40321,N_40218,N_40196);
nand U40322 (N_40322,N_40056,N_40142);
nand U40323 (N_40323,N_40242,N_40048);
xnor U40324 (N_40324,N_40171,N_40032);
and U40325 (N_40325,N_40042,N_40174);
nand U40326 (N_40326,N_40208,N_40144);
nor U40327 (N_40327,N_40091,N_40114);
or U40328 (N_40328,N_40115,N_40215);
xnor U40329 (N_40329,N_40065,N_40055);
or U40330 (N_40330,N_40034,N_40217);
and U40331 (N_40331,N_40239,N_40062);
nor U40332 (N_40332,N_40096,N_40125);
xor U40333 (N_40333,N_40089,N_40037);
or U40334 (N_40334,N_40081,N_40216);
nand U40335 (N_40335,N_40119,N_40057);
or U40336 (N_40336,N_40085,N_40066);
nand U40337 (N_40337,N_40113,N_40236);
or U40338 (N_40338,N_40249,N_40143);
and U40339 (N_40339,N_40105,N_40170);
xor U40340 (N_40340,N_40049,N_40209);
or U40341 (N_40341,N_40156,N_40076);
nor U40342 (N_40342,N_40211,N_40088);
xnor U40343 (N_40343,N_40012,N_40212);
and U40344 (N_40344,N_40197,N_40140);
nand U40345 (N_40345,N_40189,N_40214);
and U40346 (N_40346,N_40017,N_40183);
xnor U40347 (N_40347,N_40078,N_40121);
and U40348 (N_40348,N_40228,N_40001);
and U40349 (N_40349,N_40108,N_40128);
nand U40350 (N_40350,N_40023,N_40180);
and U40351 (N_40351,N_40124,N_40033);
and U40352 (N_40352,N_40015,N_40068);
and U40353 (N_40353,N_40072,N_40020);
or U40354 (N_40354,N_40199,N_40060);
nor U40355 (N_40355,N_40193,N_40028);
or U40356 (N_40356,N_40195,N_40102);
and U40357 (N_40357,N_40206,N_40220);
xnor U40358 (N_40358,N_40098,N_40024);
and U40359 (N_40359,N_40247,N_40016);
nand U40360 (N_40360,N_40238,N_40046);
nor U40361 (N_40361,N_40061,N_40163);
or U40362 (N_40362,N_40014,N_40070);
nor U40363 (N_40363,N_40130,N_40229);
nand U40364 (N_40364,N_40106,N_40185);
and U40365 (N_40365,N_40176,N_40187);
nor U40366 (N_40366,N_40029,N_40120);
nor U40367 (N_40367,N_40155,N_40000);
or U40368 (N_40368,N_40083,N_40129);
and U40369 (N_40369,N_40138,N_40173);
and U40370 (N_40370,N_40210,N_40103);
or U40371 (N_40371,N_40082,N_40011);
nand U40372 (N_40372,N_40154,N_40005);
nor U40373 (N_40373,N_40008,N_40167);
xnor U40374 (N_40374,N_40181,N_40043);
or U40375 (N_40375,N_40193,N_40180);
and U40376 (N_40376,N_40060,N_40234);
and U40377 (N_40377,N_40246,N_40216);
and U40378 (N_40378,N_40235,N_40114);
nand U40379 (N_40379,N_40239,N_40218);
xor U40380 (N_40380,N_40089,N_40040);
xnor U40381 (N_40381,N_40205,N_40046);
nand U40382 (N_40382,N_40223,N_40229);
or U40383 (N_40383,N_40241,N_40092);
and U40384 (N_40384,N_40178,N_40149);
xor U40385 (N_40385,N_40030,N_40188);
or U40386 (N_40386,N_40003,N_40205);
nand U40387 (N_40387,N_40202,N_40000);
or U40388 (N_40388,N_40071,N_40194);
nor U40389 (N_40389,N_40183,N_40145);
xnor U40390 (N_40390,N_40124,N_40144);
or U40391 (N_40391,N_40242,N_40101);
nand U40392 (N_40392,N_40123,N_40010);
nand U40393 (N_40393,N_40035,N_40224);
nor U40394 (N_40394,N_40089,N_40105);
nor U40395 (N_40395,N_40044,N_40128);
or U40396 (N_40396,N_40126,N_40137);
and U40397 (N_40397,N_40006,N_40160);
or U40398 (N_40398,N_40191,N_40026);
nor U40399 (N_40399,N_40228,N_40154);
and U40400 (N_40400,N_40042,N_40073);
xnor U40401 (N_40401,N_40092,N_40089);
xnor U40402 (N_40402,N_40003,N_40227);
and U40403 (N_40403,N_40241,N_40122);
nand U40404 (N_40404,N_40192,N_40151);
xor U40405 (N_40405,N_40242,N_40211);
nand U40406 (N_40406,N_40039,N_40067);
nor U40407 (N_40407,N_40104,N_40119);
xor U40408 (N_40408,N_40109,N_40040);
nor U40409 (N_40409,N_40117,N_40112);
xnor U40410 (N_40410,N_40193,N_40072);
xnor U40411 (N_40411,N_40177,N_40062);
nand U40412 (N_40412,N_40025,N_40074);
or U40413 (N_40413,N_40064,N_40015);
nand U40414 (N_40414,N_40169,N_40030);
or U40415 (N_40415,N_40095,N_40028);
and U40416 (N_40416,N_40175,N_40232);
nor U40417 (N_40417,N_40047,N_40215);
nor U40418 (N_40418,N_40009,N_40006);
and U40419 (N_40419,N_40153,N_40243);
and U40420 (N_40420,N_40230,N_40196);
nor U40421 (N_40421,N_40023,N_40081);
xnor U40422 (N_40422,N_40046,N_40057);
and U40423 (N_40423,N_40040,N_40179);
or U40424 (N_40424,N_40062,N_40155);
nand U40425 (N_40425,N_40107,N_40183);
nor U40426 (N_40426,N_40240,N_40223);
nand U40427 (N_40427,N_40181,N_40163);
and U40428 (N_40428,N_40198,N_40127);
nand U40429 (N_40429,N_40191,N_40186);
nand U40430 (N_40430,N_40022,N_40124);
and U40431 (N_40431,N_40102,N_40037);
xnor U40432 (N_40432,N_40050,N_40223);
nor U40433 (N_40433,N_40207,N_40056);
and U40434 (N_40434,N_40032,N_40089);
nand U40435 (N_40435,N_40171,N_40024);
nor U40436 (N_40436,N_40026,N_40040);
nor U40437 (N_40437,N_40198,N_40154);
nor U40438 (N_40438,N_40244,N_40050);
or U40439 (N_40439,N_40095,N_40103);
xnor U40440 (N_40440,N_40239,N_40057);
or U40441 (N_40441,N_40087,N_40042);
or U40442 (N_40442,N_40221,N_40242);
nand U40443 (N_40443,N_40128,N_40143);
or U40444 (N_40444,N_40183,N_40196);
and U40445 (N_40445,N_40206,N_40047);
xnor U40446 (N_40446,N_40146,N_40163);
nand U40447 (N_40447,N_40197,N_40078);
and U40448 (N_40448,N_40046,N_40248);
xor U40449 (N_40449,N_40008,N_40032);
or U40450 (N_40450,N_40214,N_40097);
and U40451 (N_40451,N_40207,N_40036);
and U40452 (N_40452,N_40168,N_40049);
and U40453 (N_40453,N_40071,N_40225);
nor U40454 (N_40454,N_40220,N_40158);
nor U40455 (N_40455,N_40048,N_40161);
and U40456 (N_40456,N_40123,N_40049);
and U40457 (N_40457,N_40189,N_40149);
nor U40458 (N_40458,N_40078,N_40123);
nor U40459 (N_40459,N_40247,N_40211);
or U40460 (N_40460,N_40025,N_40230);
nand U40461 (N_40461,N_40016,N_40087);
nor U40462 (N_40462,N_40035,N_40083);
or U40463 (N_40463,N_40171,N_40085);
nor U40464 (N_40464,N_40127,N_40118);
nor U40465 (N_40465,N_40149,N_40236);
nand U40466 (N_40466,N_40072,N_40057);
and U40467 (N_40467,N_40224,N_40167);
nand U40468 (N_40468,N_40120,N_40166);
nand U40469 (N_40469,N_40095,N_40201);
or U40470 (N_40470,N_40152,N_40003);
xor U40471 (N_40471,N_40136,N_40147);
xnor U40472 (N_40472,N_40229,N_40010);
and U40473 (N_40473,N_40206,N_40119);
xnor U40474 (N_40474,N_40188,N_40155);
nand U40475 (N_40475,N_40007,N_40132);
and U40476 (N_40476,N_40227,N_40174);
or U40477 (N_40477,N_40059,N_40068);
xor U40478 (N_40478,N_40189,N_40009);
xnor U40479 (N_40479,N_40102,N_40019);
or U40480 (N_40480,N_40090,N_40139);
or U40481 (N_40481,N_40043,N_40210);
nand U40482 (N_40482,N_40213,N_40049);
nor U40483 (N_40483,N_40191,N_40163);
nand U40484 (N_40484,N_40038,N_40212);
or U40485 (N_40485,N_40210,N_40153);
nand U40486 (N_40486,N_40116,N_40067);
or U40487 (N_40487,N_40189,N_40231);
and U40488 (N_40488,N_40186,N_40014);
nor U40489 (N_40489,N_40096,N_40139);
and U40490 (N_40490,N_40068,N_40099);
nand U40491 (N_40491,N_40036,N_40016);
nand U40492 (N_40492,N_40061,N_40165);
xnor U40493 (N_40493,N_40162,N_40229);
and U40494 (N_40494,N_40150,N_40117);
and U40495 (N_40495,N_40115,N_40164);
nand U40496 (N_40496,N_40072,N_40190);
xor U40497 (N_40497,N_40015,N_40029);
nand U40498 (N_40498,N_40097,N_40008);
nand U40499 (N_40499,N_40141,N_40151);
nand U40500 (N_40500,N_40361,N_40389);
nor U40501 (N_40501,N_40267,N_40402);
nand U40502 (N_40502,N_40297,N_40376);
nand U40503 (N_40503,N_40476,N_40286);
or U40504 (N_40504,N_40463,N_40473);
or U40505 (N_40505,N_40282,N_40265);
xnor U40506 (N_40506,N_40264,N_40342);
nand U40507 (N_40507,N_40340,N_40377);
or U40508 (N_40508,N_40479,N_40273);
or U40509 (N_40509,N_40366,N_40441);
nand U40510 (N_40510,N_40390,N_40397);
or U40511 (N_40511,N_40437,N_40275);
xnor U40512 (N_40512,N_40354,N_40445);
nand U40513 (N_40513,N_40334,N_40499);
xor U40514 (N_40514,N_40438,N_40348);
nand U40515 (N_40515,N_40324,N_40337);
xnor U40516 (N_40516,N_40276,N_40492);
and U40517 (N_40517,N_40448,N_40381);
nand U40518 (N_40518,N_40363,N_40401);
or U40519 (N_40519,N_40280,N_40458);
and U40520 (N_40520,N_40316,N_40420);
xor U40521 (N_40521,N_40422,N_40289);
or U40522 (N_40522,N_40292,N_40318);
xnor U40523 (N_40523,N_40386,N_40255);
nand U40524 (N_40524,N_40315,N_40433);
nor U40525 (N_40525,N_40452,N_40455);
and U40526 (N_40526,N_40489,N_40410);
and U40527 (N_40527,N_40460,N_40364);
and U40528 (N_40528,N_40299,N_40303);
and U40529 (N_40529,N_40278,N_40439);
nand U40530 (N_40530,N_40494,N_40260);
and U40531 (N_40531,N_40263,N_40269);
or U40532 (N_40532,N_40344,N_40317);
xnor U40533 (N_40533,N_40442,N_40333);
nor U40534 (N_40534,N_40427,N_40332);
xnor U40535 (N_40535,N_40414,N_40398);
nor U40536 (N_40536,N_40411,N_40262);
or U40537 (N_40537,N_40434,N_40314);
and U40538 (N_40538,N_40415,N_40336);
or U40539 (N_40539,N_40496,N_40321);
xor U40540 (N_40540,N_40485,N_40309);
xor U40541 (N_40541,N_40481,N_40312);
nor U40542 (N_40542,N_40279,N_40253);
or U40543 (N_40543,N_40335,N_40486);
nand U40544 (N_40544,N_40284,N_40413);
nor U40545 (N_40545,N_40406,N_40367);
xnor U40546 (N_40546,N_40394,N_40274);
nor U40547 (N_40547,N_40319,N_40369);
xor U40548 (N_40548,N_40421,N_40399);
nor U40549 (N_40549,N_40444,N_40349);
and U40550 (N_40550,N_40480,N_40283);
nor U40551 (N_40551,N_40268,N_40368);
or U40552 (N_40552,N_40302,N_40483);
and U40553 (N_40553,N_40350,N_40478);
and U40554 (N_40554,N_40290,N_40423);
nor U40555 (N_40555,N_40346,N_40287);
nand U40556 (N_40556,N_40326,N_40261);
nor U40557 (N_40557,N_40491,N_40468);
nand U40558 (N_40558,N_40374,N_40392);
xor U40559 (N_40559,N_40471,N_40428);
and U40560 (N_40560,N_40493,N_40443);
xor U40561 (N_40561,N_40484,N_40416);
or U40562 (N_40562,N_40447,N_40424);
or U40563 (N_40563,N_40372,N_40432);
xor U40564 (N_40564,N_40482,N_40327);
xor U40565 (N_40565,N_40353,N_40488);
xor U40566 (N_40566,N_40304,N_40339);
nand U40567 (N_40567,N_40288,N_40412);
and U40568 (N_40568,N_40257,N_40469);
and U40569 (N_40569,N_40379,N_40300);
and U40570 (N_40570,N_40325,N_40281);
and U40571 (N_40571,N_40251,N_40474);
and U40572 (N_40572,N_40495,N_40453);
nor U40573 (N_40573,N_40396,N_40322);
xnor U40574 (N_40574,N_40407,N_40360);
and U40575 (N_40575,N_40450,N_40409);
nand U40576 (N_40576,N_40456,N_40436);
nand U40577 (N_40577,N_40403,N_40380);
and U40578 (N_40578,N_40378,N_40250);
nor U40579 (N_40579,N_40431,N_40446);
or U40580 (N_40580,N_40295,N_40266);
or U40581 (N_40581,N_40375,N_40388);
nand U40582 (N_40582,N_40291,N_40462);
nand U40583 (N_40583,N_40254,N_40408);
xnor U40584 (N_40584,N_40311,N_40355);
and U40585 (N_40585,N_40296,N_40466);
and U40586 (N_40586,N_40341,N_40429);
or U40587 (N_40587,N_40301,N_40454);
or U40588 (N_40588,N_40293,N_40395);
or U40589 (N_40589,N_40425,N_40271);
nand U40590 (N_40590,N_40345,N_40338);
xnor U40591 (N_40591,N_40384,N_40277);
or U40592 (N_40592,N_40256,N_40457);
nand U40593 (N_40593,N_40449,N_40467);
xor U40594 (N_40594,N_40465,N_40294);
or U40595 (N_40595,N_40418,N_40298);
or U40596 (N_40596,N_40270,N_40417);
and U40597 (N_40597,N_40383,N_40459);
nor U40598 (N_40598,N_40385,N_40490);
nor U40599 (N_40599,N_40357,N_40435);
and U40600 (N_40600,N_40472,N_40464);
or U40601 (N_40601,N_40430,N_40252);
nor U40602 (N_40602,N_40373,N_40343);
and U40603 (N_40603,N_40387,N_40498);
nor U40604 (N_40604,N_40306,N_40371);
nor U40605 (N_40605,N_40331,N_40330);
and U40606 (N_40606,N_40320,N_40461);
and U40607 (N_40607,N_40358,N_40258);
or U40608 (N_40608,N_40272,N_40365);
nor U40609 (N_40609,N_40487,N_40307);
nand U40610 (N_40610,N_40352,N_40351);
and U40611 (N_40611,N_40356,N_40259);
and U40612 (N_40612,N_40305,N_40347);
xor U40613 (N_40613,N_40451,N_40382);
nand U40614 (N_40614,N_40393,N_40359);
nor U40615 (N_40615,N_40328,N_40470);
or U40616 (N_40616,N_40310,N_40370);
and U40617 (N_40617,N_40405,N_40475);
xor U40618 (N_40618,N_40440,N_40329);
and U40619 (N_40619,N_40362,N_40391);
and U40620 (N_40620,N_40426,N_40285);
nor U40621 (N_40621,N_40419,N_40404);
and U40622 (N_40622,N_40308,N_40400);
and U40623 (N_40623,N_40323,N_40477);
nor U40624 (N_40624,N_40313,N_40497);
nor U40625 (N_40625,N_40393,N_40434);
nor U40626 (N_40626,N_40392,N_40466);
nor U40627 (N_40627,N_40279,N_40423);
nor U40628 (N_40628,N_40373,N_40356);
and U40629 (N_40629,N_40403,N_40432);
and U40630 (N_40630,N_40297,N_40380);
and U40631 (N_40631,N_40419,N_40280);
or U40632 (N_40632,N_40253,N_40359);
and U40633 (N_40633,N_40406,N_40464);
nor U40634 (N_40634,N_40281,N_40447);
nand U40635 (N_40635,N_40491,N_40443);
or U40636 (N_40636,N_40464,N_40443);
nand U40637 (N_40637,N_40416,N_40402);
xnor U40638 (N_40638,N_40458,N_40459);
xor U40639 (N_40639,N_40296,N_40292);
and U40640 (N_40640,N_40252,N_40257);
nor U40641 (N_40641,N_40291,N_40348);
xor U40642 (N_40642,N_40464,N_40396);
or U40643 (N_40643,N_40300,N_40251);
and U40644 (N_40644,N_40303,N_40342);
nor U40645 (N_40645,N_40256,N_40432);
nor U40646 (N_40646,N_40316,N_40455);
nor U40647 (N_40647,N_40302,N_40296);
or U40648 (N_40648,N_40270,N_40367);
and U40649 (N_40649,N_40428,N_40366);
or U40650 (N_40650,N_40499,N_40251);
xnor U40651 (N_40651,N_40449,N_40373);
or U40652 (N_40652,N_40466,N_40361);
nand U40653 (N_40653,N_40439,N_40399);
and U40654 (N_40654,N_40300,N_40410);
or U40655 (N_40655,N_40428,N_40467);
xor U40656 (N_40656,N_40311,N_40280);
or U40657 (N_40657,N_40355,N_40400);
or U40658 (N_40658,N_40494,N_40367);
and U40659 (N_40659,N_40290,N_40437);
nor U40660 (N_40660,N_40315,N_40495);
xnor U40661 (N_40661,N_40491,N_40359);
xor U40662 (N_40662,N_40378,N_40436);
or U40663 (N_40663,N_40272,N_40366);
nand U40664 (N_40664,N_40354,N_40296);
or U40665 (N_40665,N_40338,N_40452);
nor U40666 (N_40666,N_40272,N_40330);
xnor U40667 (N_40667,N_40295,N_40495);
or U40668 (N_40668,N_40350,N_40254);
nand U40669 (N_40669,N_40361,N_40259);
xnor U40670 (N_40670,N_40323,N_40432);
or U40671 (N_40671,N_40487,N_40396);
or U40672 (N_40672,N_40336,N_40455);
nand U40673 (N_40673,N_40359,N_40274);
or U40674 (N_40674,N_40267,N_40396);
and U40675 (N_40675,N_40484,N_40469);
nor U40676 (N_40676,N_40346,N_40309);
or U40677 (N_40677,N_40370,N_40491);
and U40678 (N_40678,N_40330,N_40352);
nand U40679 (N_40679,N_40300,N_40264);
and U40680 (N_40680,N_40433,N_40435);
and U40681 (N_40681,N_40405,N_40268);
and U40682 (N_40682,N_40313,N_40370);
nand U40683 (N_40683,N_40296,N_40297);
nor U40684 (N_40684,N_40478,N_40464);
nor U40685 (N_40685,N_40446,N_40429);
or U40686 (N_40686,N_40389,N_40376);
xnor U40687 (N_40687,N_40329,N_40265);
and U40688 (N_40688,N_40260,N_40252);
or U40689 (N_40689,N_40306,N_40464);
and U40690 (N_40690,N_40432,N_40449);
nand U40691 (N_40691,N_40319,N_40371);
and U40692 (N_40692,N_40250,N_40287);
or U40693 (N_40693,N_40448,N_40286);
xor U40694 (N_40694,N_40457,N_40292);
or U40695 (N_40695,N_40322,N_40398);
and U40696 (N_40696,N_40299,N_40347);
xor U40697 (N_40697,N_40349,N_40432);
nand U40698 (N_40698,N_40419,N_40493);
and U40699 (N_40699,N_40349,N_40278);
nand U40700 (N_40700,N_40272,N_40426);
nor U40701 (N_40701,N_40357,N_40484);
nand U40702 (N_40702,N_40409,N_40481);
nand U40703 (N_40703,N_40452,N_40391);
and U40704 (N_40704,N_40324,N_40488);
nor U40705 (N_40705,N_40437,N_40488);
xor U40706 (N_40706,N_40298,N_40389);
and U40707 (N_40707,N_40337,N_40284);
nor U40708 (N_40708,N_40339,N_40315);
nor U40709 (N_40709,N_40457,N_40372);
or U40710 (N_40710,N_40331,N_40383);
nor U40711 (N_40711,N_40254,N_40436);
nor U40712 (N_40712,N_40345,N_40420);
or U40713 (N_40713,N_40380,N_40382);
nand U40714 (N_40714,N_40264,N_40316);
or U40715 (N_40715,N_40397,N_40261);
and U40716 (N_40716,N_40260,N_40311);
nor U40717 (N_40717,N_40250,N_40480);
or U40718 (N_40718,N_40461,N_40474);
and U40719 (N_40719,N_40421,N_40282);
nor U40720 (N_40720,N_40414,N_40308);
xnor U40721 (N_40721,N_40266,N_40282);
nand U40722 (N_40722,N_40386,N_40337);
nand U40723 (N_40723,N_40479,N_40376);
xor U40724 (N_40724,N_40423,N_40343);
nand U40725 (N_40725,N_40305,N_40468);
nand U40726 (N_40726,N_40375,N_40327);
nand U40727 (N_40727,N_40366,N_40398);
xor U40728 (N_40728,N_40374,N_40395);
nor U40729 (N_40729,N_40405,N_40481);
xor U40730 (N_40730,N_40310,N_40410);
or U40731 (N_40731,N_40255,N_40354);
nor U40732 (N_40732,N_40358,N_40473);
nor U40733 (N_40733,N_40322,N_40382);
and U40734 (N_40734,N_40496,N_40358);
and U40735 (N_40735,N_40367,N_40317);
or U40736 (N_40736,N_40446,N_40493);
or U40737 (N_40737,N_40406,N_40309);
nor U40738 (N_40738,N_40330,N_40306);
nor U40739 (N_40739,N_40293,N_40352);
or U40740 (N_40740,N_40404,N_40488);
nand U40741 (N_40741,N_40441,N_40293);
nor U40742 (N_40742,N_40470,N_40360);
and U40743 (N_40743,N_40456,N_40429);
xnor U40744 (N_40744,N_40252,N_40356);
and U40745 (N_40745,N_40445,N_40448);
xor U40746 (N_40746,N_40315,N_40271);
xor U40747 (N_40747,N_40253,N_40496);
or U40748 (N_40748,N_40378,N_40251);
and U40749 (N_40749,N_40339,N_40293);
and U40750 (N_40750,N_40688,N_40714);
nor U40751 (N_40751,N_40730,N_40508);
nor U40752 (N_40752,N_40536,N_40746);
and U40753 (N_40753,N_40718,N_40622);
xor U40754 (N_40754,N_40669,N_40612);
or U40755 (N_40755,N_40582,N_40571);
xnor U40756 (N_40756,N_40556,N_40701);
nor U40757 (N_40757,N_40570,N_40717);
and U40758 (N_40758,N_40545,N_40640);
or U40759 (N_40759,N_40569,N_40677);
or U40760 (N_40760,N_40560,N_40651);
or U40761 (N_40761,N_40690,N_40632);
or U40762 (N_40762,N_40599,N_40647);
nand U40763 (N_40763,N_40505,N_40627);
and U40764 (N_40764,N_40650,N_40696);
and U40765 (N_40765,N_40520,N_40748);
or U40766 (N_40766,N_40521,N_40631);
or U40767 (N_40767,N_40658,N_40512);
nor U40768 (N_40768,N_40597,N_40601);
xor U40769 (N_40769,N_40674,N_40595);
or U40770 (N_40770,N_40618,N_40643);
xnor U40771 (N_40771,N_40518,N_40742);
and U40772 (N_40772,N_40608,N_40678);
nand U40773 (N_40773,N_40708,N_40524);
and U40774 (N_40774,N_40741,N_40574);
nand U40775 (N_40775,N_40633,N_40588);
nand U40776 (N_40776,N_40619,N_40725);
nor U40777 (N_40777,N_40507,N_40541);
or U40778 (N_40778,N_40620,N_40638);
nor U40779 (N_40779,N_40724,N_40702);
xnor U40780 (N_40780,N_40728,N_40504);
nor U40781 (N_40781,N_40605,N_40698);
nor U40782 (N_40782,N_40581,N_40609);
or U40783 (N_40783,N_40692,N_40733);
nand U40784 (N_40784,N_40729,N_40707);
and U40785 (N_40785,N_40589,N_40723);
nor U40786 (N_40786,N_40598,N_40513);
nand U40787 (N_40787,N_40652,N_40747);
or U40788 (N_40788,N_40558,N_40565);
nor U40789 (N_40789,N_40517,N_40537);
and U40790 (N_40790,N_40568,N_40712);
and U40791 (N_40791,N_40555,N_40519);
nor U40792 (N_40792,N_40680,N_40639);
nand U40793 (N_40793,N_40575,N_40740);
xor U40794 (N_40794,N_40550,N_40576);
or U40795 (N_40795,N_40584,N_40745);
or U40796 (N_40796,N_40596,N_40580);
nor U40797 (N_40797,N_40654,N_40563);
and U40798 (N_40798,N_40593,N_40557);
xnor U40799 (N_40799,N_40675,N_40559);
or U40800 (N_40800,N_40511,N_40616);
xor U40801 (N_40801,N_40653,N_40590);
nand U40802 (N_40802,N_40510,N_40539);
and U40803 (N_40803,N_40611,N_40682);
nand U40804 (N_40804,N_40585,N_40749);
and U40805 (N_40805,N_40624,N_40722);
or U40806 (N_40806,N_40710,N_40657);
and U40807 (N_40807,N_40637,N_40695);
nor U40808 (N_40808,N_40679,N_40744);
or U40809 (N_40809,N_40655,N_40607);
xor U40810 (N_40810,N_40530,N_40592);
nor U40811 (N_40811,N_40705,N_40543);
and U40812 (N_40812,N_40704,N_40737);
xor U40813 (N_40813,N_40734,N_40623);
and U40814 (N_40814,N_40672,N_40703);
nand U40815 (N_40815,N_40676,N_40579);
or U40816 (N_40816,N_40661,N_40685);
and U40817 (N_40817,N_40629,N_40673);
nand U40818 (N_40818,N_40583,N_40525);
or U40819 (N_40819,N_40625,N_40529);
nor U40820 (N_40820,N_40671,N_40626);
nor U40821 (N_40821,N_40660,N_40735);
nor U40822 (N_40822,N_40614,N_40538);
or U40823 (N_40823,N_40615,N_40526);
xnor U40824 (N_40824,N_40564,N_40533);
or U40825 (N_40825,N_40630,N_40720);
and U40826 (N_40826,N_40736,N_40665);
and U40827 (N_40827,N_40726,N_40621);
and U40828 (N_40828,N_40578,N_40602);
and U40829 (N_40829,N_40683,N_40635);
nand U40830 (N_40830,N_40659,N_40523);
nand U40831 (N_40831,N_40514,N_40648);
or U40832 (N_40832,N_40547,N_40689);
xor U40833 (N_40833,N_40663,N_40561);
nor U40834 (N_40834,N_40551,N_40693);
xnor U40835 (N_40835,N_40604,N_40641);
or U40836 (N_40836,N_40515,N_40670);
or U40837 (N_40837,N_40739,N_40642);
or U40838 (N_40838,N_40540,N_40668);
or U40839 (N_40839,N_40554,N_40743);
and U40840 (N_40840,N_40586,N_40573);
nand U40841 (N_40841,N_40634,N_40534);
or U40842 (N_40842,N_40546,N_40527);
nor U40843 (N_40843,N_40681,N_40587);
or U40844 (N_40844,N_40716,N_40577);
nor U40845 (N_40845,N_40552,N_40719);
or U40846 (N_40846,N_40644,N_40732);
nor U40847 (N_40847,N_40687,N_40594);
nand U40848 (N_40848,N_40501,N_40697);
nor U40849 (N_40849,N_40553,N_40617);
or U40850 (N_40850,N_40709,N_40591);
xnor U40851 (N_40851,N_40684,N_40711);
or U40852 (N_40852,N_40699,N_40566);
or U40853 (N_40853,N_40572,N_40603);
xor U40854 (N_40854,N_40664,N_40694);
nor U40855 (N_40855,N_40613,N_40567);
and U40856 (N_40856,N_40649,N_40531);
and U40857 (N_40857,N_40610,N_40721);
or U40858 (N_40858,N_40636,N_40549);
nor U40859 (N_40859,N_40503,N_40500);
nand U40860 (N_40860,N_40516,N_40548);
or U40861 (N_40861,N_40606,N_40528);
and U40862 (N_40862,N_40509,N_40522);
and U40863 (N_40863,N_40646,N_40731);
or U40864 (N_40864,N_40535,N_40544);
or U40865 (N_40865,N_40727,N_40738);
xnor U40866 (N_40866,N_40715,N_40667);
or U40867 (N_40867,N_40686,N_40542);
nor U40868 (N_40868,N_40628,N_40656);
nor U40869 (N_40869,N_40600,N_40691);
xor U40870 (N_40870,N_40713,N_40645);
and U40871 (N_40871,N_40506,N_40532);
xnor U40872 (N_40872,N_40562,N_40700);
and U40873 (N_40873,N_40502,N_40662);
xor U40874 (N_40874,N_40706,N_40666);
nor U40875 (N_40875,N_40673,N_40559);
nand U40876 (N_40876,N_40735,N_40563);
nor U40877 (N_40877,N_40706,N_40694);
nor U40878 (N_40878,N_40667,N_40651);
or U40879 (N_40879,N_40688,N_40735);
nor U40880 (N_40880,N_40594,N_40588);
nand U40881 (N_40881,N_40509,N_40693);
xnor U40882 (N_40882,N_40737,N_40507);
nand U40883 (N_40883,N_40624,N_40709);
nor U40884 (N_40884,N_40567,N_40720);
or U40885 (N_40885,N_40640,N_40728);
nor U40886 (N_40886,N_40698,N_40513);
xor U40887 (N_40887,N_40594,N_40523);
and U40888 (N_40888,N_40697,N_40593);
and U40889 (N_40889,N_40645,N_40695);
nor U40890 (N_40890,N_40628,N_40582);
xor U40891 (N_40891,N_40596,N_40585);
and U40892 (N_40892,N_40616,N_40568);
nand U40893 (N_40893,N_40550,N_40558);
nand U40894 (N_40894,N_40662,N_40576);
xor U40895 (N_40895,N_40627,N_40658);
and U40896 (N_40896,N_40510,N_40729);
nand U40897 (N_40897,N_40596,N_40577);
and U40898 (N_40898,N_40540,N_40512);
nand U40899 (N_40899,N_40646,N_40611);
nand U40900 (N_40900,N_40545,N_40582);
xnor U40901 (N_40901,N_40578,N_40749);
nor U40902 (N_40902,N_40537,N_40669);
and U40903 (N_40903,N_40579,N_40597);
xor U40904 (N_40904,N_40558,N_40685);
or U40905 (N_40905,N_40547,N_40530);
nor U40906 (N_40906,N_40546,N_40558);
and U40907 (N_40907,N_40516,N_40643);
xor U40908 (N_40908,N_40591,N_40729);
nor U40909 (N_40909,N_40553,N_40645);
nor U40910 (N_40910,N_40523,N_40696);
and U40911 (N_40911,N_40583,N_40554);
xnor U40912 (N_40912,N_40723,N_40540);
xor U40913 (N_40913,N_40500,N_40506);
nor U40914 (N_40914,N_40556,N_40606);
xnor U40915 (N_40915,N_40611,N_40679);
xnor U40916 (N_40916,N_40632,N_40696);
and U40917 (N_40917,N_40700,N_40609);
nor U40918 (N_40918,N_40536,N_40544);
xnor U40919 (N_40919,N_40696,N_40684);
and U40920 (N_40920,N_40611,N_40675);
nand U40921 (N_40921,N_40740,N_40513);
nor U40922 (N_40922,N_40515,N_40522);
nand U40923 (N_40923,N_40572,N_40589);
nand U40924 (N_40924,N_40659,N_40504);
or U40925 (N_40925,N_40525,N_40529);
nor U40926 (N_40926,N_40562,N_40580);
nand U40927 (N_40927,N_40521,N_40625);
nor U40928 (N_40928,N_40647,N_40637);
nor U40929 (N_40929,N_40656,N_40679);
or U40930 (N_40930,N_40528,N_40669);
xnor U40931 (N_40931,N_40635,N_40636);
nor U40932 (N_40932,N_40647,N_40706);
nand U40933 (N_40933,N_40660,N_40672);
xor U40934 (N_40934,N_40612,N_40677);
and U40935 (N_40935,N_40738,N_40636);
and U40936 (N_40936,N_40663,N_40655);
or U40937 (N_40937,N_40501,N_40679);
xor U40938 (N_40938,N_40721,N_40667);
or U40939 (N_40939,N_40665,N_40629);
nor U40940 (N_40940,N_40720,N_40531);
nand U40941 (N_40941,N_40554,N_40668);
or U40942 (N_40942,N_40708,N_40652);
xnor U40943 (N_40943,N_40551,N_40748);
xnor U40944 (N_40944,N_40514,N_40670);
or U40945 (N_40945,N_40701,N_40655);
nor U40946 (N_40946,N_40682,N_40591);
nand U40947 (N_40947,N_40747,N_40673);
nor U40948 (N_40948,N_40724,N_40625);
nor U40949 (N_40949,N_40708,N_40585);
xor U40950 (N_40950,N_40574,N_40732);
nor U40951 (N_40951,N_40610,N_40649);
nand U40952 (N_40952,N_40681,N_40610);
or U40953 (N_40953,N_40529,N_40719);
nor U40954 (N_40954,N_40624,N_40679);
and U40955 (N_40955,N_40550,N_40534);
and U40956 (N_40956,N_40608,N_40558);
xnor U40957 (N_40957,N_40547,N_40706);
nand U40958 (N_40958,N_40740,N_40687);
and U40959 (N_40959,N_40560,N_40647);
or U40960 (N_40960,N_40611,N_40551);
or U40961 (N_40961,N_40690,N_40685);
or U40962 (N_40962,N_40650,N_40519);
nor U40963 (N_40963,N_40627,N_40532);
nand U40964 (N_40964,N_40517,N_40693);
nand U40965 (N_40965,N_40639,N_40529);
or U40966 (N_40966,N_40548,N_40660);
xor U40967 (N_40967,N_40589,N_40665);
or U40968 (N_40968,N_40513,N_40683);
xnor U40969 (N_40969,N_40540,N_40621);
or U40970 (N_40970,N_40526,N_40679);
and U40971 (N_40971,N_40565,N_40729);
nor U40972 (N_40972,N_40540,N_40631);
and U40973 (N_40973,N_40710,N_40543);
nor U40974 (N_40974,N_40706,N_40531);
nand U40975 (N_40975,N_40608,N_40734);
nand U40976 (N_40976,N_40502,N_40639);
and U40977 (N_40977,N_40537,N_40604);
xor U40978 (N_40978,N_40595,N_40690);
nand U40979 (N_40979,N_40605,N_40653);
or U40980 (N_40980,N_40523,N_40589);
nand U40981 (N_40981,N_40720,N_40729);
or U40982 (N_40982,N_40530,N_40697);
nand U40983 (N_40983,N_40612,N_40678);
nand U40984 (N_40984,N_40740,N_40553);
xnor U40985 (N_40985,N_40564,N_40504);
or U40986 (N_40986,N_40587,N_40666);
or U40987 (N_40987,N_40562,N_40530);
nor U40988 (N_40988,N_40555,N_40741);
or U40989 (N_40989,N_40536,N_40624);
or U40990 (N_40990,N_40722,N_40658);
nor U40991 (N_40991,N_40648,N_40524);
nand U40992 (N_40992,N_40748,N_40694);
or U40993 (N_40993,N_40538,N_40575);
nand U40994 (N_40994,N_40731,N_40673);
nor U40995 (N_40995,N_40732,N_40560);
or U40996 (N_40996,N_40630,N_40551);
nor U40997 (N_40997,N_40520,N_40567);
or U40998 (N_40998,N_40661,N_40749);
or U40999 (N_40999,N_40523,N_40634);
nor U41000 (N_41000,N_40934,N_40854);
and U41001 (N_41001,N_40856,N_40946);
and U41002 (N_41002,N_40750,N_40905);
nand U41003 (N_41003,N_40892,N_40768);
xor U41004 (N_41004,N_40834,N_40790);
xnor U41005 (N_41005,N_40929,N_40815);
nor U41006 (N_41006,N_40864,N_40766);
nor U41007 (N_41007,N_40992,N_40969);
xor U41008 (N_41008,N_40894,N_40788);
nor U41009 (N_41009,N_40852,N_40923);
xor U41010 (N_41010,N_40846,N_40812);
and U41011 (N_41011,N_40830,N_40898);
xnor U41012 (N_41012,N_40811,N_40961);
nand U41013 (N_41013,N_40887,N_40993);
nand U41014 (N_41014,N_40867,N_40770);
nand U41015 (N_41015,N_40786,N_40882);
nand U41016 (N_41016,N_40798,N_40753);
nand U41017 (N_41017,N_40782,N_40848);
or U41018 (N_41018,N_40963,N_40860);
nand U41019 (N_41019,N_40955,N_40829);
nor U41020 (N_41020,N_40941,N_40914);
xor U41021 (N_41021,N_40945,N_40986);
nand U41022 (N_41022,N_40861,N_40962);
nor U41023 (N_41023,N_40783,N_40776);
and U41024 (N_41024,N_40779,N_40775);
nor U41025 (N_41025,N_40944,N_40859);
nor U41026 (N_41026,N_40756,N_40896);
or U41027 (N_41027,N_40876,N_40889);
or U41028 (N_41028,N_40833,N_40922);
and U41029 (N_41029,N_40924,N_40937);
xor U41030 (N_41030,N_40900,N_40839);
nor U41031 (N_41031,N_40930,N_40995);
nand U41032 (N_41032,N_40762,N_40821);
or U41033 (N_41033,N_40869,N_40967);
or U41034 (N_41034,N_40844,N_40931);
nand U41035 (N_41035,N_40773,N_40857);
xor U41036 (N_41036,N_40888,N_40949);
and U41037 (N_41037,N_40990,N_40881);
xor U41038 (N_41038,N_40810,N_40965);
and U41039 (N_41039,N_40910,N_40849);
and U41040 (N_41040,N_40939,N_40917);
nand U41041 (N_41041,N_40843,N_40904);
xor U41042 (N_41042,N_40865,N_40933);
and U41043 (N_41043,N_40928,N_40960);
xor U41044 (N_41044,N_40806,N_40774);
and U41045 (N_41045,N_40801,N_40845);
or U41046 (N_41046,N_40757,N_40912);
xnor U41047 (N_41047,N_40772,N_40883);
or U41048 (N_41048,N_40789,N_40897);
or U41049 (N_41049,N_40942,N_40982);
nor U41050 (N_41050,N_40901,N_40877);
or U41051 (N_41051,N_40862,N_40855);
nor U41052 (N_41052,N_40778,N_40759);
nand U41053 (N_41053,N_40863,N_40947);
or U41054 (N_41054,N_40777,N_40909);
or U41055 (N_41055,N_40974,N_40767);
and U41056 (N_41056,N_40771,N_40755);
or U41057 (N_41057,N_40813,N_40853);
or U41058 (N_41058,N_40987,N_40765);
nand U41059 (N_41059,N_40826,N_40754);
or U41060 (N_41060,N_40875,N_40822);
nand U41061 (N_41061,N_40840,N_40948);
nor U41062 (N_41062,N_40828,N_40927);
and U41063 (N_41063,N_40906,N_40998);
xnor U41064 (N_41064,N_40968,N_40994);
nor U41065 (N_41065,N_40973,N_40915);
xnor U41066 (N_41066,N_40784,N_40884);
and U41067 (N_41067,N_40985,N_40976);
nor U41068 (N_41068,N_40919,N_40842);
nor U41069 (N_41069,N_40950,N_40886);
xnor U41070 (N_41070,N_40820,N_40911);
nand U41071 (N_41071,N_40913,N_40885);
xor U41072 (N_41072,N_40851,N_40964);
or U41073 (N_41073,N_40835,N_40925);
or U41074 (N_41074,N_40797,N_40827);
and U41075 (N_41075,N_40841,N_40999);
or U41076 (N_41076,N_40940,N_40787);
nand U41077 (N_41077,N_40796,N_40804);
or U41078 (N_41078,N_40858,N_40921);
or U41079 (N_41079,N_40758,N_40825);
nand U41080 (N_41080,N_40872,N_40805);
nand U41081 (N_41081,N_40847,N_40997);
or U41082 (N_41082,N_40763,N_40803);
nand U41083 (N_41083,N_40954,N_40808);
nand U41084 (N_41084,N_40970,N_40957);
nand U41085 (N_41085,N_40817,N_40823);
nor U41086 (N_41086,N_40926,N_40868);
nor U41087 (N_41087,N_40938,N_40819);
nor U41088 (N_41088,N_40794,N_40932);
and U41089 (N_41089,N_40959,N_40751);
nor U41090 (N_41090,N_40837,N_40907);
and U41091 (N_41091,N_40793,N_40951);
or U41092 (N_41092,N_40935,N_40781);
nand U41093 (N_41093,N_40980,N_40890);
nand U41094 (N_41094,N_40870,N_40983);
nor U41095 (N_41095,N_40989,N_40977);
or U41096 (N_41096,N_40903,N_40936);
xnor U41097 (N_41097,N_40866,N_40832);
nand U41098 (N_41098,N_40943,N_40891);
nand U41099 (N_41099,N_40952,N_40879);
nand U41100 (N_41100,N_40752,N_40908);
or U41101 (N_41101,N_40769,N_40780);
nor U41102 (N_41102,N_40984,N_40958);
or U41103 (N_41103,N_40873,N_40918);
and U41104 (N_41104,N_40972,N_40814);
xor U41105 (N_41105,N_40978,N_40996);
nor U41106 (N_41106,N_40895,N_40979);
nand U41107 (N_41107,N_40764,N_40966);
xor U41108 (N_41108,N_40893,N_40981);
nand U41109 (N_41109,N_40761,N_40807);
and U41110 (N_41110,N_40988,N_40791);
or U41111 (N_41111,N_40799,N_40874);
nand U41112 (N_41112,N_40800,N_40871);
or U41113 (N_41113,N_40956,N_40785);
nand U41114 (N_41114,N_40902,N_40809);
nand U41115 (N_41115,N_40878,N_40792);
xnor U41116 (N_41116,N_40991,N_40850);
nand U41117 (N_41117,N_40971,N_40802);
nor U41118 (N_41118,N_40831,N_40760);
xor U41119 (N_41119,N_40920,N_40953);
nand U41120 (N_41120,N_40975,N_40899);
nand U41121 (N_41121,N_40880,N_40836);
or U41122 (N_41122,N_40795,N_40816);
or U41123 (N_41123,N_40916,N_40818);
or U41124 (N_41124,N_40824,N_40838);
nor U41125 (N_41125,N_40909,N_40801);
nor U41126 (N_41126,N_40948,N_40941);
xor U41127 (N_41127,N_40793,N_40819);
nand U41128 (N_41128,N_40909,N_40798);
or U41129 (N_41129,N_40874,N_40954);
xnor U41130 (N_41130,N_40994,N_40911);
xnor U41131 (N_41131,N_40989,N_40766);
nand U41132 (N_41132,N_40888,N_40805);
nor U41133 (N_41133,N_40939,N_40823);
or U41134 (N_41134,N_40801,N_40873);
nand U41135 (N_41135,N_40936,N_40809);
nor U41136 (N_41136,N_40770,N_40932);
nor U41137 (N_41137,N_40750,N_40878);
xor U41138 (N_41138,N_40828,N_40975);
and U41139 (N_41139,N_40909,N_40948);
or U41140 (N_41140,N_40975,N_40959);
nor U41141 (N_41141,N_40944,N_40934);
nand U41142 (N_41142,N_40990,N_40791);
nor U41143 (N_41143,N_40983,N_40866);
and U41144 (N_41144,N_40979,N_40935);
xnor U41145 (N_41145,N_40889,N_40850);
xor U41146 (N_41146,N_40996,N_40845);
nor U41147 (N_41147,N_40995,N_40837);
and U41148 (N_41148,N_40992,N_40956);
nand U41149 (N_41149,N_40937,N_40839);
nand U41150 (N_41150,N_40823,N_40937);
xnor U41151 (N_41151,N_40767,N_40915);
nand U41152 (N_41152,N_40824,N_40936);
xor U41153 (N_41153,N_40847,N_40901);
nor U41154 (N_41154,N_40759,N_40942);
nor U41155 (N_41155,N_40815,N_40861);
or U41156 (N_41156,N_40990,N_40979);
nand U41157 (N_41157,N_40776,N_40850);
or U41158 (N_41158,N_40801,N_40855);
or U41159 (N_41159,N_40765,N_40960);
nor U41160 (N_41160,N_40893,N_40991);
nand U41161 (N_41161,N_40850,N_40945);
and U41162 (N_41162,N_40879,N_40941);
nor U41163 (N_41163,N_40985,N_40872);
or U41164 (N_41164,N_40813,N_40788);
or U41165 (N_41165,N_40959,N_40869);
xor U41166 (N_41166,N_40781,N_40986);
xor U41167 (N_41167,N_40954,N_40929);
nor U41168 (N_41168,N_40940,N_40783);
nor U41169 (N_41169,N_40991,N_40914);
or U41170 (N_41170,N_40898,N_40803);
or U41171 (N_41171,N_40774,N_40832);
or U41172 (N_41172,N_40765,N_40818);
nor U41173 (N_41173,N_40859,N_40868);
nand U41174 (N_41174,N_40813,N_40884);
or U41175 (N_41175,N_40993,N_40961);
xor U41176 (N_41176,N_40955,N_40919);
and U41177 (N_41177,N_40891,N_40981);
or U41178 (N_41178,N_40873,N_40756);
nand U41179 (N_41179,N_40994,N_40914);
or U41180 (N_41180,N_40757,N_40819);
and U41181 (N_41181,N_40885,N_40899);
xnor U41182 (N_41182,N_40916,N_40808);
and U41183 (N_41183,N_40926,N_40760);
xor U41184 (N_41184,N_40920,N_40858);
nand U41185 (N_41185,N_40973,N_40809);
or U41186 (N_41186,N_40951,N_40825);
nand U41187 (N_41187,N_40926,N_40988);
nand U41188 (N_41188,N_40888,N_40852);
nand U41189 (N_41189,N_40977,N_40985);
or U41190 (N_41190,N_40834,N_40825);
xnor U41191 (N_41191,N_40750,N_40846);
or U41192 (N_41192,N_40917,N_40908);
nor U41193 (N_41193,N_40910,N_40843);
or U41194 (N_41194,N_40754,N_40897);
nand U41195 (N_41195,N_40758,N_40902);
nand U41196 (N_41196,N_40961,N_40783);
and U41197 (N_41197,N_40911,N_40867);
and U41198 (N_41198,N_40826,N_40833);
or U41199 (N_41199,N_40802,N_40935);
nand U41200 (N_41200,N_40900,N_40767);
or U41201 (N_41201,N_40922,N_40999);
xor U41202 (N_41202,N_40952,N_40841);
xor U41203 (N_41203,N_40920,N_40928);
and U41204 (N_41204,N_40763,N_40920);
nor U41205 (N_41205,N_40988,N_40863);
nor U41206 (N_41206,N_40933,N_40771);
and U41207 (N_41207,N_40985,N_40992);
or U41208 (N_41208,N_40905,N_40771);
or U41209 (N_41209,N_40801,N_40826);
or U41210 (N_41210,N_40992,N_40800);
xor U41211 (N_41211,N_40809,N_40956);
nand U41212 (N_41212,N_40868,N_40954);
xnor U41213 (N_41213,N_40914,N_40770);
or U41214 (N_41214,N_40813,N_40818);
nand U41215 (N_41215,N_40862,N_40916);
nor U41216 (N_41216,N_40838,N_40928);
xor U41217 (N_41217,N_40879,N_40936);
nand U41218 (N_41218,N_40863,N_40815);
nand U41219 (N_41219,N_40905,N_40778);
xor U41220 (N_41220,N_40882,N_40865);
or U41221 (N_41221,N_40841,N_40961);
and U41222 (N_41222,N_40828,N_40913);
nor U41223 (N_41223,N_40791,N_40927);
or U41224 (N_41224,N_40966,N_40750);
nand U41225 (N_41225,N_40911,N_40876);
nor U41226 (N_41226,N_40834,N_40912);
nor U41227 (N_41227,N_40907,N_40818);
and U41228 (N_41228,N_40913,N_40943);
or U41229 (N_41229,N_40905,N_40772);
or U41230 (N_41230,N_40815,N_40915);
xnor U41231 (N_41231,N_40875,N_40796);
xnor U41232 (N_41232,N_40846,N_40809);
nand U41233 (N_41233,N_40825,N_40925);
nor U41234 (N_41234,N_40802,N_40762);
nor U41235 (N_41235,N_40954,N_40940);
and U41236 (N_41236,N_40939,N_40871);
xor U41237 (N_41237,N_40807,N_40784);
xor U41238 (N_41238,N_40896,N_40955);
nand U41239 (N_41239,N_40950,N_40782);
nor U41240 (N_41240,N_40770,N_40951);
or U41241 (N_41241,N_40767,N_40967);
and U41242 (N_41242,N_40873,N_40786);
nand U41243 (N_41243,N_40915,N_40861);
and U41244 (N_41244,N_40785,N_40840);
or U41245 (N_41245,N_40912,N_40983);
and U41246 (N_41246,N_40955,N_40810);
or U41247 (N_41247,N_40962,N_40872);
xor U41248 (N_41248,N_40947,N_40753);
xnor U41249 (N_41249,N_40828,N_40862);
and U41250 (N_41250,N_41107,N_41225);
nand U41251 (N_41251,N_41111,N_41104);
nor U41252 (N_41252,N_41005,N_41139);
or U41253 (N_41253,N_41098,N_41212);
or U41254 (N_41254,N_41035,N_41190);
and U41255 (N_41255,N_41119,N_41061);
nand U41256 (N_41256,N_41090,N_41142);
and U41257 (N_41257,N_41100,N_41122);
and U41258 (N_41258,N_41203,N_41196);
and U41259 (N_41259,N_41125,N_41024);
and U41260 (N_41260,N_41221,N_41112);
nor U41261 (N_41261,N_41143,N_41219);
nand U41262 (N_41262,N_41017,N_41235);
nor U41263 (N_41263,N_41071,N_41237);
or U41264 (N_41264,N_41247,N_41106);
nand U41265 (N_41265,N_41145,N_41049);
and U41266 (N_41266,N_41186,N_41070);
or U41267 (N_41267,N_41141,N_41078);
nand U41268 (N_41268,N_41080,N_41168);
nor U41269 (N_41269,N_41191,N_41040);
nor U41270 (N_41270,N_41195,N_41204);
nand U41271 (N_41271,N_41217,N_41057);
nor U41272 (N_41272,N_41130,N_41223);
xor U41273 (N_41273,N_41041,N_41023);
and U41274 (N_41274,N_41224,N_41150);
or U41275 (N_41275,N_41129,N_41194);
and U41276 (N_41276,N_41092,N_41038);
and U41277 (N_41277,N_41158,N_41164);
nor U41278 (N_41278,N_41004,N_41079);
nand U41279 (N_41279,N_41007,N_41026);
xor U41280 (N_41280,N_41124,N_41064);
or U41281 (N_41281,N_41175,N_41137);
nor U41282 (N_41282,N_41188,N_41095);
nand U41283 (N_41283,N_41031,N_41131);
or U41284 (N_41284,N_41058,N_41116);
nor U41285 (N_41285,N_41135,N_41206);
xnor U41286 (N_41286,N_41138,N_41181);
nand U41287 (N_41287,N_41110,N_41063);
nor U41288 (N_41288,N_41220,N_41033);
nor U41289 (N_41289,N_41075,N_41170);
or U41290 (N_41290,N_41011,N_41010);
nand U41291 (N_41291,N_41218,N_41214);
xnor U41292 (N_41292,N_41000,N_41019);
nand U41293 (N_41293,N_41121,N_41236);
and U41294 (N_41294,N_41085,N_41020);
and U41295 (N_41295,N_41199,N_41157);
and U41296 (N_41296,N_41229,N_41179);
nand U41297 (N_41297,N_41249,N_41151);
xor U41298 (N_41298,N_41184,N_41113);
or U41299 (N_41299,N_41054,N_41183);
and U41300 (N_41300,N_41097,N_41123);
nand U41301 (N_41301,N_41128,N_41083);
xor U41302 (N_41302,N_41115,N_41166);
or U41303 (N_41303,N_41034,N_41159);
and U41304 (N_41304,N_41109,N_41144);
xnor U41305 (N_41305,N_41029,N_41248);
xnor U41306 (N_41306,N_41208,N_41173);
and U41307 (N_41307,N_41072,N_41198);
and U41308 (N_41308,N_41009,N_41082);
or U41309 (N_41309,N_41044,N_41146);
or U41310 (N_41310,N_41051,N_41185);
or U41311 (N_41311,N_41055,N_41230);
or U41312 (N_41312,N_41153,N_41001);
and U41313 (N_41313,N_41155,N_41102);
xor U41314 (N_41314,N_41013,N_41227);
or U41315 (N_41315,N_41239,N_41205);
or U41316 (N_41316,N_41241,N_41028);
nand U41317 (N_41317,N_41210,N_41209);
or U41318 (N_41318,N_41134,N_41012);
nand U41319 (N_41319,N_41233,N_41118);
or U41320 (N_41320,N_41120,N_41039);
and U41321 (N_41321,N_41032,N_41086);
or U41322 (N_41322,N_41114,N_41238);
nor U41323 (N_41323,N_41231,N_41169);
and U41324 (N_41324,N_41099,N_41021);
or U41325 (N_41325,N_41165,N_41172);
nor U41326 (N_41326,N_41093,N_41003);
nor U41327 (N_41327,N_41180,N_41067);
and U41328 (N_41328,N_41088,N_41096);
or U41329 (N_41329,N_41108,N_41008);
xnor U41330 (N_41330,N_41117,N_41043);
xor U41331 (N_41331,N_41060,N_41152);
nor U41332 (N_41332,N_41066,N_41215);
and U41333 (N_41333,N_41243,N_41046);
and U41334 (N_41334,N_41213,N_41176);
or U41335 (N_41335,N_41062,N_41234);
nor U41336 (N_41336,N_41177,N_41132);
or U41337 (N_41337,N_41059,N_41201);
nor U41338 (N_41338,N_41193,N_41167);
nand U41339 (N_41339,N_41202,N_41073);
xor U41340 (N_41340,N_41014,N_41094);
nor U41341 (N_41341,N_41171,N_41045);
or U41342 (N_41342,N_41016,N_41042);
nand U41343 (N_41343,N_41018,N_41147);
nor U41344 (N_41344,N_41047,N_41052);
xor U41345 (N_41345,N_41192,N_41228);
and U41346 (N_41346,N_41222,N_41101);
nor U41347 (N_41347,N_41160,N_41189);
and U41348 (N_41348,N_41140,N_41207);
and U41349 (N_41349,N_41068,N_41050);
nor U41350 (N_41350,N_41069,N_41077);
nor U41351 (N_41351,N_41226,N_41216);
or U41352 (N_41352,N_41065,N_41126);
nand U41353 (N_41353,N_41156,N_41161);
xnor U41354 (N_41354,N_41162,N_41036);
nor U41355 (N_41355,N_41149,N_41187);
nand U41356 (N_41356,N_41197,N_41240);
nand U41357 (N_41357,N_41048,N_41002);
and U41358 (N_41358,N_41154,N_41022);
and U41359 (N_41359,N_41174,N_41245);
xor U41360 (N_41360,N_41244,N_41027);
xor U41361 (N_41361,N_41006,N_41015);
nand U41362 (N_41362,N_41163,N_41084);
nand U41363 (N_41363,N_41056,N_41127);
nor U41364 (N_41364,N_41053,N_41211);
nor U41365 (N_41365,N_41025,N_41087);
or U41366 (N_41366,N_41037,N_41089);
or U41367 (N_41367,N_41076,N_41148);
xor U41368 (N_41368,N_41200,N_41182);
nand U41369 (N_41369,N_41246,N_41136);
and U41370 (N_41370,N_41133,N_41103);
or U41371 (N_41371,N_41242,N_41232);
nand U41372 (N_41372,N_41178,N_41091);
or U41373 (N_41373,N_41030,N_41105);
nand U41374 (N_41374,N_41074,N_41081);
nand U41375 (N_41375,N_41011,N_41130);
nor U41376 (N_41376,N_41109,N_41052);
nand U41377 (N_41377,N_41055,N_41246);
and U41378 (N_41378,N_41067,N_41081);
nand U41379 (N_41379,N_41123,N_41007);
nor U41380 (N_41380,N_41086,N_41157);
xnor U41381 (N_41381,N_41039,N_41228);
nor U41382 (N_41382,N_41067,N_41247);
and U41383 (N_41383,N_41095,N_41211);
or U41384 (N_41384,N_41120,N_41125);
or U41385 (N_41385,N_41223,N_41110);
or U41386 (N_41386,N_41080,N_41181);
xor U41387 (N_41387,N_41148,N_41122);
and U41388 (N_41388,N_41088,N_41113);
nor U41389 (N_41389,N_41009,N_41216);
xor U41390 (N_41390,N_41152,N_41091);
nand U41391 (N_41391,N_41232,N_41135);
and U41392 (N_41392,N_41170,N_41093);
nand U41393 (N_41393,N_41037,N_41013);
nor U41394 (N_41394,N_41155,N_41081);
nand U41395 (N_41395,N_41241,N_41090);
xor U41396 (N_41396,N_41065,N_41100);
or U41397 (N_41397,N_41215,N_41069);
and U41398 (N_41398,N_41121,N_41117);
nand U41399 (N_41399,N_41070,N_41127);
nand U41400 (N_41400,N_41182,N_41226);
or U41401 (N_41401,N_41074,N_41159);
and U41402 (N_41402,N_41088,N_41067);
nand U41403 (N_41403,N_41246,N_41186);
and U41404 (N_41404,N_41057,N_41174);
nor U41405 (N_41405,N_41206,N_41071);
nor U41406 (N_41406,N_41190,N_41056);
nor U41407 (N_41407,N_41051,N_41170);
nor U41408 (N_41408,N_41111,N_41160);
and U41409 (N_41409,N_41055,N_41158);
nor U41410 (N_41410,N_41059,N_41190);
xnor U41411 (N_41411,N_41228,N_41135);
and U41412 (N_41412,N_41068,N_41211);
or U41413 (N_41413,N_41045,N_41096);
and U41414 (N_41414,N_41131,N_41063);
nand U41415 (N_41415,N_41194,N_41012);
or U41416 (N_41416,N_41029,N_41244);
xnor U41417 (N_41417,N_41015,N_41030);
or U41418 (N_41418,N_41105,N_41026);
xor U41419 (N_41419,N_41093,N_41113);
and U41420 (N_41420,N_41061,N_41110);
or U41421 (N_41421,N_41041,N_41038);
nand U41422 (N_41422,N_41032,N_41079);
and U41423 (N_41423,N_41149,N_41172);
and U41424 (N_41424,N_41105,N_41001);
or U41425 (N_41425,N_41244,N_41207);
xnor U41426 (N_41426,N_41049,N_41215);
nand U41427 (N_41427,N_41219,N_41043);
or U41428 (N_41428,N_41001,N_41231);
or U41429 (N_41429,N_41104,N_41086);
and U41430 (N_41430,N_41076,N_41143);
and U41431 (N_41431,N_41181,N_41232);
and U41432 (N_41432,N_41105,N_41003);
nor U41433 (N_41433,N_41045,N_41004);
nand U41434 (N_41434,N_41035,N_41130);
nand U41435 (N_41435,N_41012,N_41074);
and U41436 (N_41436,N_41086,N_41108);
nand U41437 (N_41437,N_41155,N_41208);
xnor U41438 (N_41438,N_41151,N_41147);
or U41439 (N_41439,N_41025,N_41013);
or U41440 (N_41440,N_41056,N_41071);
and U41441 (N_41441,N_41217,N_41118);
nor U41442 (N_41442,N_41085,N_41163);
nand U41443 (N_41443,N_41005,N_41115);
nand U41444 (N_41444,N_41247,N_41179);
xnor U41445 (N_41445,N_41065,N_41096);
nor U41446 (N_41446,N_41027,N_41154);
nand U41447 (N_41447,N_41082,N_41092);
or U41448 (N_41448,N_41122,N_41018);
nand U41449 (N_41449,N_41070,N_41142);
nand U41450 (N_41450,N_41041,N_41161);
nand U41451 (N_41451,N_41148,N_41025);
nand U41452 (N_41452,N_41098,N_41132);
nand U41453 (N_41453,N_41197,N_41009);
nor U41454 (N_41454,N_41023,N_41092);
and U41455 (N_41455,N_41228,N_41072);
nand U41456 (N_41456,N_41103,N_41093);
and U41457 (N_41457,N_41189,N_41113);
nor U41458 (N_41458,N_41227,N_41229);
and U41459 (N_41459,N_41172,N_41099);
or U41460 (N_41460,N_41069,N_41248);
and U41461 (N_41461,N_41109,N_41005);
and U41462 (N_41462,N_41176,N_41059);
nor U41463 (N_41463,N_41092,N_41244);
or U41464 (N_41464,N_41225,N_41076);
xor U41465 (N_41465,N_41131,N_41040);
nor U41466 (N_41466,N_41095,N_41070);
and U41467 (N_41467,N_41116,N_41219);
and U41468 (N_41468,N_41181,N_41132);
nand U41469 (N_41469,N_41122,N_41195);
and U41470 (N_41470,N_41237,N_41106);
xor U41471 (N_41471,N_41075,N_41122);
nand U41472 (N_41472,N_41086,N_41042);
or U41473 (N_41473,N_41108,N_41085);
nor U41474 (N_41474,N_41155,N_41241);
nor U41475 (N_41475,N_41149,N_41095);
nand U41476 (N_41476,N_41007,N_41104);
and U41477 (N_41477,N_41125,N_41235);
nand U41478 (N_41478,N_41133,N_41155);
nand U41479 (N_41479,N_41026,N_41014);
and U41480 (N_41480,N_41096,N_41174);
and U41481 (N_41481,N_41104,N_41097);
nand U41482 (N_41482,N_41057,N_41220);
nor U41483 (N_41483,N_41052,N_41182);
xnor U41484 (N_41484,N_41077,N_41113);
xnor U41485 (N_41485,N_41087,N_41147);
or U41486 (N_41486,N_41145,N_41159);
xor U41487 (N_41487,N_41089,N_41209);
xnor U41488 (N_41488,N_41170,N_41030);
nand U41489 (N_41489,N_41194,N_41068);
nor U41490 (N_41490,N_41095,N_41028);
and U41491 (N_41491,N_41070,N_41214);
and U41492 (N_41492,N_41094,N_41059);
or U41493 (N_41493,N_41186,N_41124);
and U41494 (N_41494,N_41160,N_41013);
and U41495 (N_41495,N_41023,N_41031);
nor U41496 (N_41496,N_41106,N_41217);
and U41497 (N_41497,N_41188,N_41147);
xnor U41498 (N_41498,N_41136,N_41009);
and U41499 (N_41499,N_41035,N_41183);
and U41500 (N_41500,N_41265,N_41287);
xor U41501 (N_41501,N_41307,N_41254);
nand U41502 (N_41502,N_41489,N_41370);
and U41503 (N_41503,N_41279,N_41253);
xnor U41504 (N_41504,N_41405,N_41469);
nor U41505 (N_41505,N_41461,N_41331);
or U41506 (N_41506,N_41406,N_41393);
nor U41507 (N_41507,N_41472,N_41388);
or U41508 (N_41508,N_41484,N_41366);
or U41509 (N_41509,N_41264,N_41398);
or U41510 (N_41510,N_41262,N_41414);
nor U41511 (N_41511,N_41493,N_41435);
xnor U41512 (N_41512,N_41453,N_41288);
nor U41513 (N_41513,N_41436,N_41334);
or U41514 (N_41514,N_41263,N_41460);
and U41515 (N_41515,N_41261,N_41467);
nor U41516 (N_41516,N_41434,N_41286);
and U41517 (N_41517,N_41457,N_41409);
and U41518 (N_41518,N_41458,N_41323);
or U41519 (N_41519,N_41297,N_41449);
or U41520 (N_41520,N_41252,N_41289);
nor U41521 (N_41521,N_41255,N_41306);
xor U41522 (N_41522,N_41296,N_41421);
or U41523 (N_41523,N_41448,N_41468);
nand U41524 (N_41524,N_41269,N_41401);
nor U41525 (N_41525,N_41383,N_41431);
nand U41526 (N_41526,N_41420,N_41367);
and U41527 (N_41527,N_41382,N_41350);
xor U41528 (N_41528,N_41303,N_41266);
and U41529 (N_41529,N_41392,N_41298);
and U41530 (N_41530,N_41352,N_41408);
or U41531 (N_41531,N_41313,N_41474);
nor U41532 (N_41532,N_41378,N_41429);
nor U41533 (N_41533,N_41379,N_41339);
nand U41534 (N_41534,N_41490,N_41250);
nor U41535 (N_41535,N_41327,N_41369);
nor U41536 (N_41536,N_41305,N_41477);
xnor U41537 (N_41537,N_41415,N_41364);
xor U41538 (N_41538,N_41341,N_41462);
nor U41539 (N_41539,N_41277,N_41395);
xor U41540 (N_41540,N_41437,N_41322);
xor U41541 (N_41541,N_41342,N_41309);
and U41542 (N_41542,N_41329,N_41438);
nor U41543 (N_41543,N_41432,N_41347);
or U41544 (N_41544,N_41372,N_41485);
xnor U41545 (N_41545,N_41445,N_41486);
and U41546 (N_41546,N_41441,N_41451);
nor U41547 (N_41547,N_41481,N_41256);
xnor U41548 (N_41548,N_41335,N_41348);
and U41549 (N_41549,N_41345,N_41285);
xnor U41550 (N_41550,N_41425,N_41386);
and U41551 (N_41551,N_41362,N_41430);
xor U41552 (N_41552,N_41272,N_41482);
or U41553 (N_41553,N_41267,N_41260);
nor U41554 (N_41554,N_41273,N_41308);
xnor U41555 (N_41555,N_41332,N_41428);
xnor U41556 (N_41556,N_41257,N_41333);
nor U41557 (N_41557,N_41385,N_41371);
or U41558 (N_41558,N_41299,N_41410);
nor U41559 (N_41559,N_41473,N_41316);
nand U41560 (N_41560,N_41280,N_41283);
nor U41561 (N_41561,N_41376,N_41315);
nand U41562 (N_41562,N_41403,N_41471);
xnor U41563 (N_41563,N_41390,N_41317);
xnor U41564 (N_41564,N_41497,N_41291);
nand U41565 (N_41565,N_41358,N_41381);
xor U41566 (N_41566,N_41326,N_41355);
and U41567 (N_41567,N_41466,N_41427);
and U41568 (N_41568,N_41290,N_41498);
nand U41569 (N_41569,N_41433,N_41278);
xnor U41570 (N_41570,N_41251,N_41359);
xor U41571 (N_41571,N_41455,N_41375);
or U41572 (N_41572,N_41495,N_41496);
or U41573 (N_41573,N_41271,N_41447);
and U41574 (N_41574,N_41349,N_41446);
xnor U41575 (N_41575,N_41399,N_41397);
or U41576 (N_41576,N_41293,N_41494);
and U41577 (N_41577,N_41368,N_41353);
nor U41578 (N_41578,N_41417,N_41318);
or U41579 (N_41579,N_41363,N_41454);
nand U41580 (N_41580,N_41423,N_41488);
and U41581 (N_41581,N_41480,N_41470);
and U41582 (N_41582,N_41419,N_41444);
xor U41583 (N_41583,N_41336,N_41478);
nor U41584 (N_41584,N_41344,N_41294);
nor U41585 (N_41585,N_41391,N_41284);
nand U41586 (N_41586,N_41389,N_41301);
xor U41587 (N_41587,N_41463,N_41499);
and U41588 (N_41588,N_41281,N_41354);
xnor U41589 (N_41589,N_41356,N_41422);
or U41590 (N_41590,N_41325,N_41407);
nor U41591 (N_41591,N_41411,N_41314);
xor U41592 (N_41592,N_41340,N_41270);
nand U41593 (N_41593,N_41412,N_41337);
or U41594 (N_41594,N_41459,N_41450);
and U41595 (N_41595,N_41377,N_41443);
nand U41596 (N_41596,N_41338,N_41259);
xor U41597 (N_41597,N_41258,N_41365);
nor U41598 (N_41598,N_41319,N_41274);
nor U41599 (N_41599,N_41402,N_41464);
and U41600 (N_41600,N_41452,N_41357);
and U41601 (N_41601,N_41492,N_41304);
and U41602 (N_41602,N_41312,N_41439);
or U41603 (N_41603,N_41320,N_41300);
xnor U41604 (N_41604,N_41276,N_41275);
xnor U41605 (N_41605,N_41343,N_41440);
or U41606 (N_41606,N_41346,N_41311);
nand U41607 (N_41607,N_41310,N_41418);
or U41608 (N_41608,N_41479,N_41328);
xnor U41609 (N_41609,N_41374,N_41400);
nor U41610 (N_41610,N_41475,N_41295);
and U41611 (N_41611,N_41413,N_41292);
xnor U41612 (N_41612,N_41442,N_41426);
and U41613 (N_41613,N_41465,N_41360);
xor U41614 (N_41614,N_41387,N_41321);
or U41615 (N_41615,N_41380,N_41324);
nand U41616 (N_41616,N_41491,N_41483);
and U41617 (N_41617,N_41361,N_41384);
nor U41618 (N_41618,N_41302,N_41487);
nor U41619 (N_41619,N_41456,N_41351);
xnor U41620 (N_41620,N_41396,N_41373);
or U41621 (N_41621,N_41282,N_41404);
and U41622 (N_41622,N_41476,N_41394);
or U41623 (N_41623,N_41268,N_41416);
nor U41624 (N_41624,N_41330,N_41424);
nand U41625 (N_41625,N_41473,N_41451);
nor U41626 (N_41626,N_41318,N_41387);
nand U41627 (N_41627,N_41493,N_41425);
or U41628 (N_41628,N_41294,N_41310);
nand U41629 (N_41629,N_41342,N_41266);
and U41630 (N_41630,N_41319,N_41374);
or U41631 (N_41631,N_41359,N_41325);
xor U41632 (N_41632,N_41309,N_41325);
or U41633 (N_41633,N_41346,N_41328);
and U41634 (N_41634,N_41482,N_41432);
or U41635 (N_41635,N_41427,N_41473);
nor U41636 (N_41636,N_41280,N_41309);
xnor U41637 (N_41637,N_41250,N_41284);
and U41638 (N_41638,N_41459,N_41268);
nor U41639 (N_41639,N_41269,N_41375);
xnor U41640 (N_41640,N_41318,N_41295);
and U41641 (N_41641,N_41341,N_41474);
or U41642 (N_41642,N_41452,N_41403);
or U41643 (N_41643,N_41337,N_41400);
nor U41644 (N_41644,N_41343,N_41480);
and U41645 (N_41645,N_41396,N_41363);
nor U41646 (N_41646,N_41368,N_41494);
or U41647 (N_41647,N_41393,N_41278);
nor U41648 (N_41648,N_41288,N_41364);
nand U41649 (N_41649,N_41276,N_41476);
nor U41650 (N_41650,N_41316,N_41366);
and U41651 (N_41651,N_41474,N_41446);
and U41652 (N_41652,N_41345,N_41290);
xor U41653 (N_41653,N_41356,N_41469);
and U41654 (N_41654,N_41458,N_41331);
xnor U41655 (N_41655,N_41288,N_41435);
xnor U41656 (N_41656,N_41366,N_41385);
nor U41657 (N_41657,N_41346,N_41441);
and U41658 (N_41658,N_41492,N_41369);
xor U41659 (N_41659,N_41262,N_41432);
or U41660 (N_41660,N_41379,N_41385);
nor U41661 (N_41661,N_41375,N_41383);
xnor U41662 (N_41662,N_41297,N_41447);
nor U41663 (N_41663,N_41369,N_41478);
nor U41664 (N_41664,N_41472,N_41355);
and U41665 (N_41665,N_41486,N_41257);
nor U41666 (N_41666,N_41269,N_41424);
xor U41667 (N_41667,N_41298,N_41350);
and U41668 (N_41668,N_41362,N_41261);
nor U41669 (N_41669,N_41317,N_41448);
xor U41670 (N_41670,N_41423,N_41481);
nand U41671 (N_41671,N_41419,N_41265);
nand U41672 (N_41672,N_41423,N_41306);
xor U41673 (N_41673,N_41392,N_41397);
nor U41674 (N_41674,N_41429,N_41369);
and U41675 (N_41675,N_41377,N_41382);
xnor U41676 (N_41676,N_41370,N_41298);
and U41677 (N_41677,N_41487,N_41376);
nand U41678 (N_41678,N_41424,N_41412);
nand U41679 (N_41679,N_41295,N_41250);
or U41680 (N_41680,N_41325,N_41320);
nor U41681 (N_41681,N_41441,N_41315);
or U41682 (N_41682,N_41478,N_41364);
nand U41683 (N_41683,N_41309,N_41431);
and U41684 (N_41684,N_41379,N_41466);
or U41685 (N_41685,N_41482,N_41385);
or U41686 (N_41686,N_41285,N_41447);
nand U41687 (N_41687,N_41435,N_41457);
nand U41688 (N_41688,N_41329,N_41284);
and U41689 (N_41689,N_41434,N_41330);
and U41690 (N_41690,N_41301,N_41455);
or U41691 (N_41691,N_41365,N_41452);
and U41692 (N_41692,N_41481,N_41482);
nand U41693 (N_41693,N_41346,N_41286);
and U41694 (N_41694,N_41391,N_41305);
or U41695 (N_41695,N_41415,N_41428);
and U41696 (N_41696,N_41425,N_41483);
xor U41697 (N_41697,N_41311,N_41402);
nand U41698 (N_41698,N_41403,N_41386);
nand U41699 (N_41699,N_41489,N_41443);
or U41700 (N_41700,N_41355,N_41409);
or U41701 (N_41701,N_41489,N_41384);
or U41702 (N_41702,N_41334,N_41347);
and U41703 (N_41703,N_41380,N_41322);
xor U41704 (N_41704,N_41434,N_41265);
xnor U41705 (N_41705,N_41329,N_41465);
and U41706 (N_41706,N_41296,N_41367);
nand U41707 (N_41707,N_41317,N_41392);
and U41708 (N_41708,N_41382,N_41353);
or U41709 (N_41709,N_41466,N_41392);
nand U41710 (N_41710,N_41320,N_41337);
nor U41711 (N_41711,N_41452,N_41280);
and U41712 (N_41712,N_41399,N_41382);
or U41713 (N_41713,N_41431,N_41484);
or U41714 (N_41714,N_41384,N_41473);
or U41715 (N_41715,N_41258,N_41395);
or U41716 (N_41716,N_41370,N_41408);
and U41717 (N_41717,N_41386,N_41463);
and U41718 (N_41718,N_41442,N_41384);
nand U41719 (N_41719,N_41302,N_41382);
or U41720 (N_41720,N_41401,N_41288);
xnor U41721 (N_41721,N_41423,N_41448);
nand U41722 (N_41722,N_41313,N_41386);
or U41723 (N_41723,N_41261,N_41302);
nand U41724 (N_41724,N_41450,N_41447);
nand U41725 (N_41725,N_41252,N_41406);
nor U41726 (N_41726,N_41315,N_41344);
or U41727 (N_41727,N_41474,N_41489);
and U41728 (N_41728,N_41405,N_41302);
and U41729 (N_41729,N_41352,N_41436);
nor U41730 (N_41730,N_41345,N_41398);
nor U41731 (N_41731,N_41303,N_41250);
nor U41732 (N_41732,N_41293,N_41410);
nand U41733 (N_41733,N_41432,N_41333);
nor U41734 (N_41734,N_41441,N_41401);
nand U41735 (N_41735,N_41349,N_41408);
xor U41736 (N_41736,N_41406,N_41273);
xnor U41737 (N_41737,N_41294,N_41335);
nor U41738 (N_41738,N_41279,N_41391);
nor U41739 (N_41739,N_41415,N_41251);
and U41740 (N_41740,N_41490,N_41260);
or U41741 (N_41741,N_41436,N_41419);
nor U41742 (N_41742,N_41458,N_41340);
or U41743 (N_41743,N_41386,N_41269);
nor U41744 (N_41744,N_41250,N_41475);
xor U41745 (N_41745,N_41283,N_41415);
nand U41746 (N_41746,N_41337,N_41472);
or U41747 (N_41747,N_41485,N_41262);
nand U41748 (N_41748,N_41485,N_41379);
nor U41749 (N_41749,N_41403,N_41314);
and U41750 (N_41750,N_41740,N_41570);
or U41751 (N_41751,N_41621,N_41505);
xor U41752 (N_41752,N_41622,N_41628);
nand U41753 (N_41753,N_41540,N_41514);
or U41754 (N_41754,N_41536,N_41610);
nor U41755 (N_41755,N_41549,N_41634);
xor U41756 (N_41756,N_41685,N_41704);
nor U41757 (N_41757,N_41544,N_41512);
and U41758 (N_41758,N_41601,N_41609);
or U41759 (N_41759,N_41555,N_41525);
or U41760 (N_41760,N_41551,N_41572);
nand U41761 (N_41761,N_41697,N_41503);
nor U41762 (N_41762,N_41730,N_41595);
nor U41763 (N_41763,N_41640,N_41613);
or U41764 (N_41764,N_41558,N_41743);
or U41765 (N_41765,N_41705,N_41600);
nor U41766 (N_41766,N_41591,N_41585);
nor U41767 (N_41767,N_41552,N_41581);
nor U41768 (N_41768,N_41589,N_41666);
and U41769 (N_41769,N_41664,N_41650);
or U41770 (N_41770,N_41542,N_41627);
nor U41771 (N_41771,N_41508,N_41599);
or U41772 (N_41772,N_41626,N_41729);
xor U41773 (N_41773,N_41559,N_41716);
or U41774 (N_41774,N_41654,N_41594);
and U41775 (N_41775,N_41598,N_41550);
nor U41776 (N_41776,N_41534,N_41547);
nand U41777 (N_41777,N_41562,N_41571);
and U41778 (N_41778,N_41695,N_41513);
and U41779 (N_41779,N_41645,N_41701);
and U41780 (N_41780,N_41588,N_41702);
nor U41781 (N_41781,N_41619,N_41501);
or U41782 (N_41782,N_41708,N_41672);
or U41783 (N_41783,N_41691,N_41633);
xor U41784 (N_41784,N_41733,N_41578);
or U41785 (N_41785,N_41561,N_41735);
or U41786 (N_41786,N_41517,N_41587);
nor U41787 (N_41787,N_41727,N_41745);
and U41788 (N_41788,N_41620,N_41658);
nor U41789 (N_41789,N_41584,N_41742);
nor U41790 (N_41790,N_41644,N_41686);
xor U41791 (N_41791,N_41519,N_41712);
nor U41792 (N_41792,N_41659,N_41535);
nand U41793 (N_41793,N_41582,N_41662);
or U41794 (N_41794,N_41511,N_41749);
or U41795 (N_41795,N_41681,N_41603);
and U41796 (N_41796,N_41728,N_41569);
nor U41797 (N_41797,N_41541,N_41665);
nand U41798 (N_41798,N_41618,N_41698);
nand U41799 (N_41799,N_41631,N_41526);
or U41800 (N_41800,N_41635,N_41671);
nor U41801 (N_41801,N_41639,N_41532);
or U41802 (N_41802,N_41538,N_41683);
or U41803 (N_41803,N_41597,N_41656);
nand U41804 (N_41804,N_41652,N_41586);
xor U41805 (N_41805,N_41611,N_41545);
and U41806 (N_41806,N_41593,N_41673);
nor U41807 (N_41807,N_41524,N_41653);
nor U41808 (N_41808,N_41573,N_41516);
nor U41809 (N_41809,N_41567,N_41509);
xnor U41810 (N_41810,N_41703,N_41692);
or U41811 (N_41811,N_41537,N_41579);
and U41812 (N_41812,N_41630,N_41606);
xnor U41813 (N_41813,N_41518,N_41688);
xnor U41814 (N_41814,N_41713,N_41527);
nor U41815 (N_41815,N_41604,N_41614);
and U41816 (N_41816,N_41707,N_41546);
nand U41817 (N_41817,N_41515,N_41523);
nand U41818 (N_41818,N_41566,N_41649);
xor U41819 (N_41819,N_41677,N_41734);
xnor U41820 (N_41820,N_41646,N_41608);
nand U41821 (N_41821,N_41694,N_41719);
xnor U41822 (N_41822,N_41605,N_41655);
or U41823 (N_41823,N_41636,N_41577);
and U41824 (N_41824,N_41616,N_41739);
or U41825 (N_41825,N_41641,N_41724);
nor U41826 (N_41826,N_41736,N_41741);
nor U41827 (N_41827,N_41720,N_41731);
and U41828 (N_41828,N_41667,N_41732);
xnor U41829 (N_41829,N_41642,N_41590);
xnor U41830 (N_41830,N_41661,N_41583);
xor U41831 (N_41831,N_41564,N_41710);
nand U41832 (N_41832,N_41674,N_41696);
or U41833 (N_41833,N_41592,N_41629);
or U41834 (N_41834,N_41738,N_41543);
and U41835 (N_41835,N_41510,N_41623);
or U41836 (N_41836,N_41596,N_41651);
or U41837 (N_41837,N_41663,N_41647);
and U41838 (N_41838,N_41657,N_41612);
xor U41839 (N_41839,N_41682,N_41747);
nor U41840 (N_41840,N_41721,N_41560);
nand U41841 (N_41841,N_41529,N_41563);
and U41842 (N_41842,N_41748,N_41557);
and U41843 (N_41843,N_41744,N_41675);
nand U41844 (N_41844,N_41531,N_41722);
nor U41845 (N_41845,N_41726,N_41548);
or U41846 (N_41846,N_41507,N_41676);
and U41847 (N_41847,N_41680,N_41615);
or U41848 (N_41848,N_41607,N_41714);
xor U41849 (N_41849,N_41679,N_41746);
nand U41850 (N_41850,N_41556,N_41693);
nor U41851 (N_41851,N_41553,N_41678);
or U41852 (N_41852,N_41687,N_41624);
xnor U41853 (N_41853,N_41709,N_41725);
nor U41854 (N_41854,N_41643,N_41554);
nand U41855 (N_41855,N_41568,N_41520);
or U41856 (N_41856,N_41699,N_41638);
nor U41857 (N_41857,N_41602,N_41580);
xnor U41858 (N_41858,N_41670,N_41723);
or U41859 (N_41859,N_41689,N_41528);
and U41860 (N_41860,N_41668,N_41533);
or U41861 (N_41861,N_41530,N_41706);
and U41862 (N_41862,N_41711,N_41522);
nor U41863 (N_41863,N_41637,N_41700);
nor U41864 (N_41864,N_41576,N_41715);
or U41865 (N_41865,N_41617,N_41521);
nand U41866 (N_41866,N_41575,N_41718);
nor U41867 (N_41867,N_41500,N_41717);
xor U41868 (N_41868,N_41502,N_41632);
nand U41869 (N_41869,N_41574,N_41669);
xor U41870 (N_41870,N_41690,N_41504);
xor U41871 (N_41871,N_41506,N_41648);
or U41872 (N_41872,N_41539,N_41684);
nand U41873 (N_41873,N_41625,N_41660);
nor U41874 (N_41874,N_41737,N_41565);
nand U41875 (N_41875,N_41636,N_41558);
or U41876 (N_41876,N_41699,N_41665);
xor U41877 (N_41877,N_41688,N_41576);
and U41878 (N_41878,N_41720,N_41549);
xor U41879 (N_41879,N_41684,N_41745);
nand U41880 (N_41880,N_41552,N_41688);
or U41881 (N_41881,N_41583,N_41636);
nor U41882 (N_41882,N_41508,N_41563);
xor U41883 (N_41883,N_41731,N_41741);
xnor U41884 (N_41884,N_41552,N_41662);
or U41885 (N_41885,N_41674,N_41516);
nand U41886 (N_41886,N_41714,N_41731);
nor U41887 (N_41887,N_41581,N_41538);
nand U41888 (N_41888,N_41637,N_41740);
nor U41889 (N_41889,N_41523,N_41714);
or U41890 (N_41890,N_41503,N_41556);
xnor U41891 (N_41891,N_41607,N_41649);
nor U41892 (N_41892,N_41518,N_41737);
nand U41893 (N_41893,N_41724,N_41640);
or U41894 (N_41894,N_41571,N_41709);
nor U41895 (N_41895,N_41604,N_41646);
or U41896 (N_41896,N_41578,N_41589);
or U41897 (N_41897,N_41709,N_41527);
and U41898 (N_41898,N_41636,N_41665);
nand U41899 (N_41899,N_41547,N_41572);
nand U41900 (N_41900,N_41559,N_41617);
xnor U41901 (N_41901,N_41665,N_41504);
or U41902 (N_41902,N_41679,N_41516);
and U41903 (N_41903,N_41633,N_41596);
xnor U41904 (N_41904,N_41522,N_41641);
nand U41905 (N_41905,N_41655,N_41597);
nand U41906 (N_41906,N_41694,N_41538);
nor U41907 (N_41907,N_41696,N_41594);
nor U41908 (N_41908,N_41556,N_41739);
or U41909 (N_41909,N_41580,N_41536);
xnor U41910 (N_41910,N_41578,N_41679);
nor U41911 (N_41911,N_41600,N_41740);
nand U41912 (N_41912,N_41581,N_41709);
nor U41913 (N_41913,N_41712,N_41550);
nand U41914 (N_41914,N_41519,N_41513);
xnor U41915 (N_41915,N_41511,N_41660);
and U41916 (N_41916,N_41658,N_41735);
or U41917 (N_41917,N_41639,N_41583);
nor U41918 (N_41918,N_41665,N_41728);
nor U41919 (N_41919,N_41743,N_41500);
xnor U41920 (N_41920,N_41603,N_41599);
xor U41921 (N_41921,N_41581,N_41667);
xnor U41922 (N_41922,N_41530,N_41623);
xnor U41923 (N_41923,N_41603,N_41675);
nand U41924 (N_41924,N_41645,N_41519);
xor U41925 (N_41925,N_41702,N_41638);
or U41926 (N_41926,N_41731,N_41685);
or U41927 (N_41927,N_41645,N_41508);
nor U41928 (N_41928,N_41566,N_41597);
nand U41929 (N_41929,N_41673,N_41736);
or U41930 (N_41930,N_41711,N_41649);
or U41931 (N_41931,N_41628,N_41616);
and U41932 (N_41932,N_41748,N_41649);
xor U41933 (N_41933,N_41657,N_41660);
or U41934 (N_41934,N_41641,N_41572);
xor U41935 (N_41935,N_41533,N_41590);
nand U41936 (N_41936,N_41539,N_41552);
or U41937 (N_41937,N_41515,N_41698);
nor U41938 (N_41938,N_41515,N_41595);
and U41939 (N_41939,N_41700,N_41641);
and U41940 (N_41940,N_41679,N_41720);
xor U41941 (N_41941,N_41652,N_41651);
nand U41942 (N_41942,N_41659,N_41584);
and U41943 (N_41943,N_41672,N_41640);
and U41944 (N_41944,N_41707,N_41639);
xor U41945 (N_41945,N_41718,N_41697);
nor U41946 (N_41946,N_41652,N_41710);
and U41947 (N_41947,N_41620,N_41593);
xnor U41948 (N_41948,N_41517,N_41615);
xor U41949 (N_41949,N_41564,N_41539);
or U41950 (N_41950,N_41513,N_41601);
nand U41951 (N_41951,N_41642,N_41588);
and U41952 (N_41952,N_41659,N_41631);
nand U41953 (N_41953,N_41595,N_41736);
xnor U41954 (N_41954,N_41609,N_41579);
xnor U41955 (N_41955,N_41542,N_41714);
and U41956 (N_41956,N_41620,N_41712);
or U41957 (N_41957,N_41630,N_41642);
nand U41958 (N_41958,N_41749,N_41580);
and U41959 (N_41959,N_41527,N_41562);
xor U41960 (N_41960,N_41510,N_41604);
nor U41961 (N_41961,N_41519,N_41621);
and U41962 (N_41962,N_41734,N_41661);
and U41963 (N_41963,N_41561,N_41733);
or U41964 (N_41964,N_41688,N_41633);
xor U41965 (N_41965,N_41699,N_41550);
and U41966 (N_41966,N_41561,N_41508);
nand U41967 (N_41967,N_41657,N_41564);
and U41968 (N_41968,N_41610,N_41505);
nor U41969 (N_41969,N_41688,N_41506);
and U41970 (N_41970,N_41559,N_41726);
or U41971 (N_41971,N_41623,N_41692);
or U41972 (N_41972,N_41658,N_41644);
or U41973 (N_41973,N_41585,N_41561);
nand U41974 (N_41974,N_41680,N_41683);
and U41975 (N_41975,N_41606,N_41587);
nor U41976 (N_41976,N_41635,N_41696);
and U41977 (N_41977,N_41706,N_41592);
nand U41978 (N_41978,N_41735,N_41562);
or U41979 (N_41979,N_41539,N_41713);
or U41980 (N_41980,N_41745,N_41685);
nor U41981 (N_41981,N_41544,N_41638);
or U41982 (N_41982,N_41644,N_41695);
nand U41983 (N_41983,N_41514,N_41717);
or U41984 (N_41984,N_41642,N_41545);
xnor U41985 (N_41985,N_41717,N_41517);
or U41986 (N_41986,N_41637,N_41718);
or U41987 (N_41987,N_41524,N_41626);
and U41988 (N_41988,N_41595,N_41596);
or U41989 (N_41989,N_41531,N_41671);
nand U41990 (N_41990,N_41599,N_41694);
or U41991 (N_41991,N_41622,N_41570);
and U41992 (N_41992,N_41591,N_41558);
xor U41993 (N_41993,N_41504,N_41545);
nor U41994 (N_41994,N_41699,N_41506);
xnor U41995 (N_41995,N_41589,N_41587);
xor U41996 (N_41996,N_41673,N_41741);
or U41997 (N_41997,N_41690,N_41637);
nand U41998 (N_41998,N_41591,N_41677);
and U41999 (N_41999,N_41717,N_41582);
or U42000 (N_42000,N_41959,N_41794);
xnor U42001 (N_42001,N_41962,N_41758);
and U42002 (N_42002,N_41900,N_41789);
or U42003 (N_42003,N_41927,N_41826);
xnor U42004 (N_42004,N_41818,N_41958);
nor U42005 (N_42005,N_41919,N_41876);
nand U42006 (N_42006,N_41854,N_41879);
nand U42007 (N_42007,N_41866,N_41842);
or U42008 (N_42008,N_41947,N_41841);
nand U42009 (N_42009,N_41825,N_41976);
nand U42010 (N_42010,N_41917,N_41892);
nor U42011 (N_42011,N_41851,N_41961);
nand U42012 (N_42012,N_41817,N_41756);
and U42013 (N_42013,N_41885,N_41881);
nand U42014 (N_42014,N_41869,N_41935);
nand U42015 (N_42015,N_41787,N_41994);
nand U42016 (N_42016,N_41882,N_41824);
and U42017 (N_42017,N_41875,N_41932);
nor U42018 (N_42018,N_41894,N_41844);
xor U42019 (N_42019,N_41920,N_41915);
xor U42020 (N_42020,N_41948,N_41993);
nor U42021 (N_42021,N_41938,N_41857);
xor U42022 (N_42022,N_41849,N_41823);
xnor U42023 (N_42023,N_41904,N_41923);
nand U42024 (N_42024,N_41767,N_41858);
nand U42025 (N_42025,N_41949,N_41788);
nor U42026 (N_42026,N_41783,N_41835);
nor U42027 (N_42027,N_41831,N_41821);
xor U42028 (N_42028,N_41969,N_41804);
or U42029 (N_42029,N_41896,N_41760);
xnor U42030 (N_42030,N_41886,N_41906);
and U42031 (N_42031,N_41769,N_41921);
and U42032 (N_42032,N_41999,N_41863);
nand U42033 (N_42033,N_41889,N_41888);
or U42034 (N_42034,N_41860,N_41991);
nand U42035 (N_42035,N_41805,N_41763);
nor U42036 (N_42036,N_41862,N_41980);
xnor U42037 (N_42037,N_41782,N_41751);
nand U42038 (N_42038,N_41931,N_41806);
and U42039 (N_42039,N_41853,N_41903);
nor U42040 (N_42040,N_41852,N_41759);
and U42041 (N_42041,N_41953,N_41971);
xor U42042 (N_42042,N_41868,N_41890);
nor U42043 (N_42043,N_41790,N_41791);
and U42044 (N_42044,N_41848,N_41928);
xnor U42045 (N_42045,N_41929,N_41954);
nand U42046 (N_42046,N_41984,N_41941);
or U42047 (N_42047,N_41872,N_41752);
and U42048 (N_42048,N_41865,N_41795);
xor U42049 (N_42049,N_41846,N_41796);
and U42050 (N_42050,N_41902,N_41968);
nand U42051 (N_42051,N_41779,N_41770);
nand U42052 (N_42052,N_41891,N_41799);
nor U42053 (N_42053,N_41813,N_41785);
nor U42054 (N_42054,N_41987,N_41803);
or U42055 (N_42055,N_41768,N_41861);
nor U42056 (N_42056,N_41772,N_41916);
nor U42057 (N_42057,N_41833,N_41974);
nor U42058 (N_42058,N_41814,N_41811);
xnor U42059 (N_42059,N_41998,N_41897);
or U42060 (N_42060,N_41992,N_41899);
and U42061 (N_42061,N_41955,N_41859);
xor U42062 (N_42062,N_41855,N_41940);
or U42063 (N_42063,N_41777,N_41942);
nor U42064 (N_42064,N_41981,N_41781);
and U42065 (N_42065,N_41771,N_41778);
or U42066 (N_42066,N_41986,N_41775);
or U42067 (N_42067,N_41887,N_41750);
and U42068 (N_42068,N_41832,N_41944);
and U42069 (N_42069,N_41830,N_41840);
xor U42070 (N_42070,N_41800,N_41989);
and U42071 (N_42071,N_41901,N_41815);
nand U42072 (N_42072,N_41878,N_41913);
and U42073 (N_42073,N_41850,N_41809);
nor U42074 (N_42074,N_41965,N_41978);
nand U42075 (N_42075,N_41952,N_41801);
nor U42076 (N_42076,N_41925,N_41943);
nor U42077 (N_42077,N_41951,N_41977);
nand U42078 (N_42078,N_41979,N_41945);
or U42079 (N_42079,N_41997,N_41983);
nor U42080 (N_42080,N_41930,N_41793);
and U42081 (N_42081,N_41936,N_41757);
or U42082 (N_42082,N_41911,N_41797);
or U42083 (N_42083,N_41922,N_41985);
or U42084 (N_42084,N_41776,N_41773);
nor U42085 (N_42085,N_41963,N_41988);
nand U42086 (N_42086,N_41867,N_41960);
and U42087 (N_42087,N_41926,N_41990);
nand U42088 (N_42088,N_41845,N_41812);
nand U42089 (N_42089,N_41895,N_41972);
and U42090 (N_42090,N_41820,N_41838);
nor U42091 (N_42091,N_41827,N_41964);
nand U42092 (N_42092,N_41754,N_41786);
nor U42093 (N_42093,N_41834,N_41847);
or U42094 (N_42094,N_41950,N_41764);
xnor U42095 (N_42095,N_41880,N_41856);
nand U42096 (N_42096,N_41905,N_41908);
and U42097 (N_42097,N_41924,N_41909);
or U42098 (N_42098,N_41877,N_41873);
xor U42099 (N_42099,N_41808,N_41761);
and U42100 (N_42100,N_41956,N_41807);
xor U42101 (N_42101,N_41762,N_41883);
nor U42102 (N_42102,N_41934,N_41870);
nand U42103 (N_42103,N_41802,N_41798);
nor U42104 (N_42104,N_41816,N_41996);
nor U42105 (N_42105,N_41837,N_41982);
xor U42106 (N_42106,N_41874,N_41939);
xnor U42107 (N_42107,N_41884,N_41864);
nand U42108 (N_42108,N_41907,N_41753);
nand U42109 (N_42109,N_41918,N_41765);
nand U42110 (N_42110,N_41946,N_41914);
nand U42111 (N_42111,N_41822,N_41893);
xor U42112 (N_42112,N_41819,N_41784);
nor U42113 (N_42113,N_41937,N_41973);
nor U42114 (N_42114,N_41810,N_41755);
or U42115 (N_42115,N_41843,N_41766);
xnor U42116 (N_42116,N_41792,N_41828);
xnor U42117 (N_42117,N_41910,N_41970);
or U42118 (N_42118,N_41898,N_41871);
nor U42119 (N_42119,N_41829,N_41966);
nor U42120 (N_42120,N_41975,N_41836);
nand U42121 (N_42121,N_41995,N_41957);
xnor U42122 (N_42122,N_41933,N_41774);
nor U42123 (N_42123,N_41912,N_41780);
xor U42124 (N_42124,N_41967,N_41839);
and U42125 (N_42125,N_41931,N_41866);
xnor U42126 (N_42126,N_41967,N_41836);
xor U42127 (N_42127,N_41760,N_41774);
and U42128 (N_42128,N_41995,N_41795);
nand U42129 (N_42129,N_41891,N_41992);
and U42130 (N_42130,N_41793,N_41812);
nand U42131 (N_42131,N_41914,N_41919);
or U42132 (N_42132,N_41869,N_41918);
nor U42133 (N_42133,N_41868,N_41757);
xnor U42134 (N_42134,N_41949,N_41786);
nor U42135 (N_42135,N_41871,N_41955);
or U42136 (N_42136,N_41790,N_41921);
nand U42137 (N_42137,N_41914,N_41950);
and U42138 (N_42138,N_41783,N_41912);
xor U42139 (N_42139,N_41885,N_41938);
xor U42140 (N_42140,N_41753,N_41786);
nand U42141 (N_42141,N_41826,N_41936);
nand U42142 (N_42142,N_41907,N_41992);
or U42143 (N_42143,N_41798,N_41784);
nor U42144 (N_42144,N_41792,N_41848);
nand U42145 (N_42145,N_41902,N_41927);
and U42146 (N_42146,N_41787,N_41944);
nand U42147 (N_42147,N_41837,N_41848);
nand U42148 (N_42148,N_41965,N_41791);
or U42149 (N_42149,N_41900,N_41888);
nor U42150 (N_42150,N_41879,N_41762);
or U42151 (N_42151,N_41880,N_41797);
nand U42152 (N_42152,N_41981,N_41911);
nand U42153 (N_42153,N_41909,N_41939);
or U42154 (N_42154,N_41957,N_41903);
and U42155 (N_42155,N_41780,N_41927);
nand U42156 (N_42156,N_41965,N_41900);
nor U42157 (N_42157,N_41771,N_41833);
or U42158 (N_42158,N_41826,N_41858);
and U42159 (N_42159,N_41926,N_41841);
nor U42160 (N_42160,N_41802,N_41930);
nand U42161 (N_42161,N_41956,N_41918);
or U42162 (N_42162,N_41842,N_41755);
or U42163 (N_42163,N_41896,N_41846);
nor U42164 (N_42164,N_41980,N_41968);
nor U42165 (N_42165,N_41805,N_41784);
nor U42166 (N_42166,N_41943,N_41964);
xor U42167 (N_42167,N_41816,N_41845);
xor U42168 (N_42168,N_41806,N_41774);
nor U42169 (N_42169,N_41949,N_41987);
xnor U42170 (N_42170,N_41828,N_41905);
and U42171 (N_42171,N_41787,N_41770);
nand U42172 (N_42172,N_41814,N_41812);
nor U42173 (N_42173,N_41941,N_41889);
xnor U42174 (N_42174,N_41821,N_41973);
and U42175 (N_42175,N_41918,N_41954);
nand U42176 (N_42176,N_41834,N_41966);
nand U42177 (N_42177,N_41888,N_41883);
and U42178 (N_42178,N_41943,N_41965);
and U42179 (N_42179,N_41841,N_41980);
and U42180 (N_42180,N_41814,N_41877);
nand U42181 (N_42181,N_41838,N_41794);
nand U42182 (N_42182,N_41797,N_41931);
nor U42183 (N_42183,N_41889,N_41911);
or U42184 (N_42184,N_41954,N_41943);
or U42185 (N_42185,N_41914,N_41849);
xnor U42186 (N_42186,N_41783,N_41905);
nand U42187 (N_42187,N_41762,N_41888);
nor U42188 (N_42188,N_41989,N_41946);
nor U42189 (N_42189,N_41983,N_41942);
nand U42190 (N_42190,N_41908,N_41866);
or U42191 (N_42191,N_41761,N_41955);
nor U42192 (N_42192,N_41924,N_41964);
or U42193 (N_42193,N_41871,N_41945);
nor U42194 (N_42194,N_41861,N_41906);
xnor U42195 (N_42195,N_41768,N_41931);
xor U42196 (N_42196,N_41966,N_41766);
and U42197 (N_42197,N_41828,N_41942);
nand U42198 (N_42198,N_41913,N_41970);
or U42199 (N_42199,N_41993,N_41995);
nand U42200 (N_42200,N_41981,N_41786);
xnor U42201 (N_42201,N_41907,N_41979);
nand U42202 (N_42202,N_41943,N_41942);
xor U42203 (N_42203,N_41863,N_41990);
nand U42204 (N_42204,N_41958,N_41942);
or U42205 (N_42205,N_41799,N_41807);
nand U42206 (N_42206,N_41781,N_41917);
nand U42207 (N_42207,N_41883,N_41828);
nor U42208 (N_42208,N_41978,N_41751);
nor U42209 (N_42209,N_41847,N_41849);
and U42210 (N_42210,N_41988,N_41910);
nor U42211 (N_42211,N_41911,N_41986);
xnor U42212 (N_42212,N_41771,N_41884);
nor U42213 (N_42213,N_41781,N_41886);
and U42214 (N_42214,N_41978,N_41953);
and U42215 (N_42215,N_41760,N_41998);
nor U42216 (N_42216,N_41827,N_41975);
nor U42217 (N_42217,N_41904,N_41772);
or U42218 (N_42218,N_41949,N_41836);
nor U42219 (N_42219,N_41881,N_41768);
nor U42220 (N_42220,N_41924,N_41991);
nand U42221 (N_42221,N_41771,N_41913);
and U42222 (N_42222,N_41778,N_41956);
and U42223 (N_42223,N_41780,N_41751);
nor U42224 (N_42224,N_41769,N_41823);
nor U42225 (N_42225,N_41815,N_41937);
or U42226 (N_42226,N_41886,N_41896);
and U42227 (N_42227,N_41795,N_41875);
nand U42228 (N_42228,N_41915,N_41858);
xor U42229 (N_42229,N_41999,N_41873);
nand U42230 (N_42230,N_41976,N_41944);
nand U42231 (N_42231,N_41826,N_41836);
xor U42232 (N_42232,N_41936,N_41884);
nand U42233 (N_42233,N_41782,N_41903);
nor U42234 (N_42234,N_41777,N_41773);
xor U42235 (N_42235,N_41835,N_41880);
nor U42236 (N_42236,N_41774,N_41910);
nand U42237 (N_42237,N_41824,N_41860);
nor U42238 (N_42238,N_41953,N_41923);
or U42239 (N_42239,N_41804,N_41955);
nor U42240 (N_42240,N_41899,N_41834);
xnor U42241 (N_42241,N_41947,N_41815);
nor U42242 (N_42242,N_41890,N_41913);
nand U42243 (N_42243,N_41997,N_41944);
nor U42244 (N_42244,N_41897,N_41896);
nand U42245 (N_42245,N_41967,N_41850);
or U42246 (N_42246,N_41855,N_41951);
nor U42247 (N_42247,N_41909,N_41789);
and U42248 (N_42248,N_41903,N_41940);
nor U42249 (N_42249,N_41779,N_41946);
nor U42250 (N_42250,N_42104,N_42137);
xnor U42251 (N_42251,N_42192,N_42131);
nor U42252 (N_42252,N_42233,N_42012);
or U42253 (N_42253,N_42117,N_42109);
or U42254 (N_42254,N_42173,N_42010);
xor U42255 (N_42255,N_42157,N_42247);
or U42256 (N_42256,N_42048,N_42070);
xor U42257 (N_42257,N_42001,N_42249);
and U42258 (N_42258,N_42000,N_42176);
or U42259 (N_42259,N_42055,N_42092);
or U42260 (N_42260,N_42130,N_42095);
or U42261 (N_42261,N_42189,N_42182);
and U42262 (N_42262,N_42146,N_42038);
nor U42263 (N_42263,N_42178,N_42172);
nor U42264 (N_42264,N_42188,N_42080);
xnor U42265 (N_42265,N_42236,N_42023);
or U42266 (N_42266,N_42138,N_42198);
nor U42267 (N_42267,N_42083,N_42149);
xor U42268 (N_42268,N_42110,N_42101);
nand U42269 (N_42269,N_42145,N_42240);
nand U42270 (N_42270,N_42125,N_42147);
xor U42271 (N_42271,N_42047,N_42114);
and U42272 (N_42272,N_42091,N_42165);
and U42273 (N_42273,N_42150,N_42015);
nor U42274 (N_42274,N_42021,N_42170);
and U42275 (N_42275,N_42196,N_42013);
and U42276 (N_42276,N_42132,N_42036);
and U42277 (N_42277,N_42209,N_42090);
and U42278 (N_42278,N_42206,N_42052);
nor U42279 (N_42279,N_42089,N_42153);
xnor U42280 (N_42280,N_42190,N_42232);
xor U42281 (N_42281,N_42243,N_42102);
nor U42282 (N_42282,N_42239,N_42241);
or U42283 (N_42283,N_42027,N_42123);
and U42284 (N_42284,N_42111,N_42121);
xor U42285 (N_42285,N_42042,N_42174);
xor U42286 (N_42286,N_42098,N_42113);
and U42287 (N_42287,N_42032,N_42056);
nor U42288 (N_42288,N_42040,N_42016);
nor U42289 (N_42289,N_42009,N_42100);
nor U42290 (N_42290,N_42006,N_42143);
xor U42291 (N_42291,N_42112,N_42028);
or U42292 (N_42292,N_42144,N_42118);
nand U42293 (N_42293,N_42064,N_42007);
or U42294 (N_42294,N_42093,N_42246);
and U42295 (N_42295,N_42078,N_42214);
and U42296 (N_42296,N_42163,N_42034);
nand U42297 (N_42297,N_42162,N_42195);
nor U42298 (N_42298,N_42051,N_42177);
or U42299 (N_42299,N_42031,N_42216);
nor U42300 (N_42300,N_42181,N_42059);
nand U42301 (N_42301,N_42066,N_42008);
nor U42302 (N_42302,N_42079,N_42072);
nand U42303 (N_42303,N_42230,N_42183);
nor U42304 (N_42304,N_42201,N_42075);
or U42305 (N_42305,N_42152,N_42053);
nor U42306 (N_42306,N_42186,N_42218);
nand U42307 (N_42307,N_42030,N_42211);
xor U42308 (N_42308,N_42199,N_42002);
nor U42309 (N_42309,N_42122,N_42203);
nor U42310 (N_42310,N_42107,N_42175);
or U42311 (N_42311,N_42073,N_42019);
nand U42312 (N_42312,N_42069,N_42158);
nand U42313 (N_42313,N_42097,N_42081);
and U42314 (N_42314,N_42180,N_42035);
and U42315 (N_42315,N_42142,N_42215);
or U42316 (N_42316,N_42024,N_42018);
or U42317 (N_42317,N_42129,N_42060);
xnor U42318 (N_42318,N_42088,N_42187);
nor U42319 (N_42319,N_42154,N_42205);
nand U42320 (N_42320,N_42228,N_42161);
nor U42321 (N_42321,N_42245,N_42200);
or U42322 (N_42322,N_42184,N_42194);
nor U42323 (N_42323,N_42108,N_42061);
and U42324 (N_42324,N_42005,N_42223);
or U42325 (N_42325,N_42140,N_42054);
nand U42326 (N_42326,N_42025,N_42076);
and U42327 (N_42327,N_42045,N_42179);
xor U42328 (N_42328,N_42248,N_42139);
xnor U42329 (N_42329,N_42026,N_42065);
nand U42330 (N_42330,N_42231,N_42050);
or U42331 (N_42331,N_42220,N_42085);
nor U42332 (N_42332,N_42128,N_42222);
or U42333 (N_42333,N_42166,N_42197);
xor U42334 (N_42334,N_42116,N_42043);
xor U42335 (N_42335,N_42103,N_42224);
xor U42336 (N_42336,N_42227,N_42039);
and U42337 (N_42337,N_42004,N_42105);
or U42338 (N_42338,N_42234,N_42167);
or U42339 (N_42339,N_42124,N_42164);
xor U42340 (N_42340,N_42014,N_42082);
nor U42341 (N_42341,N_42225,N_42074);
xnor U42342 (N_42342,N_42096,N_42003);
nor U42343 (N_42343,N_42126,N_42219);
nand U42344 (N_42344,N_42046,N_42135);
nor U42345 (N_42345,N_42221,N_42115);
nand U42346 (N_42346,N_42204,N_42160);
or U42347 (N_42347,N_42141,N_42071);
xnor U42348 (N_42348,N_42087,N_42086);
or U42349 (N_42349,N_42029,N_42169);
nand U42350 (N_42350,N_42207,N_42148);
nand U42351 (N_42351,N_42244,N_42242);
nand U42352 (N_42352,N_42067,N_42120);
or U42353 (N_42353,N_42058,N_42063);
nand U42354 (N_42354,N_42068,N_42099);
or U42355 (N_42355,N_42133,N_42057);
or U42356 (N_42356,N_42193,N_42134);
xor U42357 (N_42357,N_42062,N_42022);
xnor U42358 (N_42358,N_42235,N_42077);
and U42359 (N_42359,N_42084,N_42155);
xor U42360 (N_42360,N_42119,N_42168);
nor U42361 (N_42361,N_42044,N_42212);
or U42362 (N_42362,N_42017,N_42185);
xnor U42363 (N_42363,N_42208,N_42171);
or U42364 (N_42364,N_42226,N_42229);
nor U42365 (N_42365,N_42217,N_42151);
nand U42366 (N_42366,N_42106,N_42213);
and U42367 (N_42367,N_42037,N_42127);
xnor U42368 (N_42368,N_42238,N_42033);
xor U42369 (N_42369,N_42191,N_42136);
xor U42370 (N_42370,N_42237,N_42020);
or U42371 (N_42371,N_42210,N_42156);
xor U42372 (N_42372,N_42159,N_42094);
nor U42373 (N_42373,N_42202,N_42049);
nand U42374 (N_42374,N_42041,N_42011);
or U42375 (N_42375,N_42014,N_42130);
nand U42376 (N_42376,N_42190,N_42165);
nor U42377 (N_42377,N_42010,N_42017);
and U42378 (N_42378,N_42031,N_42022);
or U42379 (N_42379,N_42216,N_42141);
and U42380 (N_42380,N_42231,N_42191);
nand U42381 (N_42381,N_42157,N_42246);
nor U42382 (N_42382,N_42170,N_42140);
or U42383 (N_42383,N_42079,N_42026);
nand U42384 (N_42384,N_42239,N_42164);
and U42385 (N_42385,N_42154,N_42098);
nand U42386 (N_42386,N_42046,N_42108);
nor U42387 (N_42387,N_42003,N_42239);
or U42388 (N_42388,N_42183,N_42243);
or U42389 (N_42389,N_42246,N_42175);
nand U42390 (N_42390,N_42199,N_42092);
or U42391 (N_42391,N_42137,N_42129);
xnor U42392 (N_42392,N_42171,N_42006);
or U42393 (N_42393,N_42138,N_42220);
nand U42394 (N_42394,N_42178,N_42174);
xor U42395 (N_42395,N_42157,N_42090);
and U42396 (N_42396,N_42097,N_42134);
nor U42397 (N_42397,N_42153,N_42141);
and U42398 (N_42398,N_42057,N_42223);
or U42399 (N_42399,N_42180,N_42061);
xnor U42400 (N_42400,N_42010,N_42009);
and U42401 (N_42401,N_42213,N_42053);
and U42402 (N_42402,N_42227,N_42049);
or U42403 (N_42403,N_42127,N_42170);
xor U42404 (N_42404,N_42247,N_42236);
nand U42405 (N_42405,N_42211,N_42134);
nor U42406 (N_42406,N_42001,N_42152);
or U42407 (N_42407,N_42190,N_42036);
nor U42408 (N_42408,N_42186,N_42013);
or U42409 (N_42409,N_42119,N_42200);
nand U42410 (N_42410,N_42095,N_42238);
and U42411 (N_42411,N_42134,N_42064);
nor U42412 (N_42412,N_42046,N_42019);
nor U42413 (N_42413,N_42016,N_42221);
nand U42414 (N_42414,N_42031,N_42130);
or U42415 (N_42415,N_42164,N_42237);
nand U42416 (N_42416,N_42031,N_42190);
or U42417 (N_42417,N_42048,N_42137);
nor U42418 (N_42418,N_42145,N_42190);
nor U42419 (N_42419,N_42082,N_42025);
and U42420 (N_42420,N_42022,N_42118);
and U42421 (N_42421,N_42011,N_42181);
or U42422 (N_42422,N_42108,N_42000);
or U42423 (N_42423,N_42035,N_42008);
nor U42424 (N_42424,N_42065,N_42195);
xnor U42425 (N_42425,N_42056,N_42064);
nor U42426 (N_42426,N_42203,N_42049);
or U42427 (N_42427,N_42134,N_42181);
and U42428 (N_42428,N_42119,N_42203);
nor U42429 (N_42429,N_42241,N_42213);
or U42430 (N_42430,N_42144,N_42001);
and U42431 (N_42431,N_42237,N_42104);
or U42432 (N_42432,N_42089,N_42102);
and U42433 (N_42433,N_42105,N_42134);
nor U42434 (N_42434,N_42196,N_42230);
xnor U42435 (N_42435,N_42218,N_42054);
nand U42436 (N_42436,N_42013,N_42045);
xor U42437 (N_42437,N_42013,N_42095);
nand U42438 (N_42438,N_42012,N_42167);
nor U42439 (N_42439,N_42057,N_42216);
nor U42440 (N_42440,N_42116,N_42137);
and U42441 (N_42441,N_42033,N_42194);
nand U42442 (N_42442,N_42018,N_42168);
and U42443 (N_42443,N_42125,N_42118);
or U42444 (N_42444,N_42080,N_42067);
xnor U42445 (N_42445,N_42184,N_42155);
or U42446 (N_42446,N_42164,N_42153);
and U42447 (N_42447,N_42203,N_42012);
nand U42448 (N_42448,N_42047,N_42208);
nand U42449 (N_42449,N_42124,N_42157);
xnor U42450 (N_42450,N_42150,N_42033);
and U42451 (N_42451,N_42055,N_42181);
xnor U42452 (N_42452,N_42224,N_42136);
or U42453 (N_42453,N_42038,N_42167);
or U42454 (N_42454,N_42121,N_42202);
xnor U42455 (N_42455,N_42062,N_42025);
or U42456 (N_42456,N_42223,N_42097);
nand U42457 (N_42457,N_42161,N_42169);
nand U42458 (N_42458,N_42045,N_42088);
and U42459 (N_42459,N_42033,N_42154);
or U42460 (N_42460,N_42088,N_42111);
and U42461 (N_42461,N_42202,N_42158);
or U42462 (N_42462,N_42167,N_42240);
nand U42463 (N_42463,N_42037,N_42192);
xor U42464 (N_42464,N_42101,N_42104);
or U42465 (N_42465,N_42077,N_42083);
nand U42466 (N_42466,N_42070,N_42201);
nor U42467 (N_42467,N_42024,N_42236);
nand U42468 (N_42468,N_42021,N_42125);
or U42469 (N_42469,N_42165,N_42009);
nand U42470 (N_42470,N_42130,N_42100);
nand U42471 (N_42471,N_42055,N_42036);
and U42472 (N_42472,N_42062,N_42202);
or U42473 (N_42473,N_42121,N_42215);
nand U42474 (N_42474,N_42201,N_42243);
xor U42475 (N_42475,N_42199,N_42081);
xor U42476 (N_42476,N_42180,N_42131);
and U42477 (N_42477,N_42022,N_42154);
xor U42478 (N_42478,N_42095,N_42232);
nand U42479 (N_42479,N_42088,N_42101);
nor U42480 (N_42480,N_42190,N_42080);
xnor U42481 (N_42481,N_42222,N_42011);
nand U42482 (N_42482,N_42071,N_42145);
nor U42483 (N_42483,N_42242,N_42192);
and U42484 (N_42484,N_42231,N_42103);
and U42485 (N_42485,N_42010,N_42238);
and U42486 (N_42486,N_42222,N_42196);
or U42487 (N_42487,N_42238,N_42047);
nand U42488 (N_42488,N_42247,N_42186);
xor U42489 (N_42489,N_42019,N_42206);
and U42490 (N_42490,N_42236,N_42123);
nand U42491 (N_42491,N_42131,N_42183);
and U42492 (N_42492,N_42196,N_42070);
nor U42493 (N_42493,N_42080,N_42059);
or U42494 (N_42494,N_42057,N_42235);
or U42495 (N_42495,N_42035,N_42227);
nor U42496 (N_42496,N_42242,N_42059);
nor U42497 (N_42497,N_42064,N_42244);
or U42498 (N_42498,N_42132,N_42183);
or U42499 (N_42499,N_42084,N_42219);
and U42500 (N_42500,N_42351,N_42321);
xnor U42501 (N_42501,N_42473,N_42482);
nand U42502 (N_42502,N_42336,N_42279);
and U42503 (N_42503,N_42440,N_42460);
nor U42504 (N_42504,N_42376,N_42464);
and U42505 (N_42505,N_42450,N_42338);
nor U42506 (N_42506,N_42382,N_42381);
xnor U42507 (N_42507,N_42467,N_42419);
and U42508 (N_42508,N_42379,N_42433);
and U42509 (N_42509,N_42404,N_42295);
and U42510 (N_42510,N_42385,N_42454);
nor U42511 (N_42511,N_42451,N_42253);
nor U42512 (N_42512,N_42493,N_42488);
nand U42513 (N_42513,N_42395,N_42353);
or U42514 (N_42514,N_42416,N_42424);
nand U42515 (N_42515,N_42388,N_42480);
nor U42516 (N_42516,N_42402,N_42337);
xnor U42517 (N_42517,N_42282,N_42400);
xnor U42518 (N_42518,N_42462,N_42259);
xor U42519 (N_42519,N_42341,N_42409);
and U42520 (N_42520,N_42278,N_42357);
xnor U42521 (N_42521,N_42479,N_42463);
nand U42522 (N_42522,N_42334,N_42387);
or U42523 (N_42523,N_42293,N_42324);
nand U42524 (N_42524,N_42481,N_42367);
or U42525 (N_42525,N_42318,N_42486);
xnor U42526 (N_42526,N_42350,N_42390);
and U42527 (N_42527,N_42291,N_42355);
nor U42528 (N_42528,N_42363,N_42372);
nand U42529 (N_42529,N_42301,N_42459);
xnor U42530 (N_42530,N_42446,N_42343);
and U42531 (N_42531,N_42252,N_42359);
nand U42532 (N_42532,N_42270,N_42365);
or U42533 (N_42533,N_42417,N_42292);
nand U42534 (N_42534,N_42375,N_42275);
and U42535 (N_42535,N_42431,N_42313);
xor U42536 (N_42536,N_42352,N_42250);
and U42537 (N_42537,N_42380,N_42333);
and U42538 (N_42538,N_42474,N_42491);
nor U42539 (N_42539,N_42384,N_42420);
xor U42540 (N_42540,N_42429,N_42284);
xor U42541 (N_42541,N_42323,N_42255);
or U42542 (N_42542,N_42347,N_42316);
nand U42543 (N_42543,N_42345,N_42406);
nand U42544 (N_42544,N_42281,N_42271);
nor U42545 (N_42545,N_42344,N_42436);
nand U42546 (N_42546,N_42490,N_42418);
and U42547 (N_42547,N_42399,N_42427);
nor U42548 (N_42548,N_42428,N_42314);
nand U42549 (N_42549,N_42302,N_42311);
xnor U42550 (N_42550,N_42330,N_42398);
or U42551 (N_42551,N_42494,N_42361);
or U42552 (N_42552,N_42413,N_42499);
nand U42553 (N_42553,N_42465,N_42453);
and U42554 (N_42554,N_42447,N_42438);
nand U42555 (N_42555,N_42435,N_42458);
nor U42556 (N_42556,N_42315,N_42368);
and U42557 (N_42557,N_42394,N_42408);
nand U42558 (N_42558,N_42466,N_42448);
nor U42559 (N_42559,N_42423,N_42461);
xor U42560 (N_42560,N_42303,N_42439);
and U42561 (N_42561,N_42331,N_42274);
nand U42562 (N_42562,N_42405,N_42339);
nand U42563 (N_42563,N_42266,N_42412);
or U42564 (N_42564,N_42285,N_42349);
nor U42565 (N_42565,N_42434,N_42469);
and U42566 (N_42566,N_42265,N_42442);
or U42567 (N_42567,N_42422,N_42426);
and U42568 (N_42568,N_42342,N_42470);
or U42569 (N_42569,N_42306,N_42410);
nor U42570 (N_42570,N_42283,N_42298);
nand U42571 (N_42571,N_42319,N_42362);
nand U42572 (N_42572,N_42370,N_42391);
nor U42573 (N_42573,N_42476,N_42322);
and U42574 (N_42574,N_42325,N_42262);
xor U42575 (N_42575,N_42441,N_42307);
xor U42576 (N_42576,N_42421,N_42386);
and U42577 (N_42577,N_42263,N_42437);
nand U42578 (N_42578,N_42378,N_42373);
and U42579 (N_42579,N_42309,N_42492);
or U42580 (N_42580,N_42444,N_42320);
xor U42581 (N_42581,N_42300,N_42468);
and U42582 (N_42582,N_42354,N_42280);
nand U42583 (N_42583,N_42276,N_42327);
or U42584 (N_42584,N_42260,N_42475);
and U42585 (N_42585,N_42407,N_42432);
xnor U42586 (N_42586,N_42335,N_42403);
and U42587 (N_42587,N_42272,N_42267);
and U42588 (N_42588,N_42346,N_42471);
nand U42589 (N_42589,N_42393,N_42425);
xnor U42590 (N_42590,N_42414,N_42358);
xnor U42591 (N_42591,N_42477,N_42340);
nor U42592 (N_42592,N_42366,N_42452);
or U42593 (N_42593,N_42401,N_42288);
xnor U42594 (N_42594,N_42328,N_42397);
or U42595 (N_42595,N_42277,N_42483);
nor U42596 (N_42596,N_42286,N_42411);
nand U42597 (N_42597,N_42369,N_42305);
xnor U42598 (N_42598,N_42257,N_42496);
nor U42599 (N_42599,N_42383,N_42299);
or U42600 (N_42600,N_42392,N_42485);
xor U42601 (N_42601,N_42415,N_42478);
or U42602 (N_42602,N_42294,N_42374);
nor U42603 (N_42603,N_42348,N_42254);
and U42604 (N_42604,N_42489,N_42256);
nor U42605 (N_42605,N_42290,N_42455);
and U42606 (N_42606,N_42430,N_42389);
xor U42607 (N_42607,N_42326,N_42360);
nand U42608 (N_42608,N_42457,N_42487);
and U42609 (N_42609,N_42445,N_42449);
and U42610 (N_42610,N_42317,N_42304);
or U42611 (N_42611,N_42443,N_42377);
nand U42612 (N_42612,N_42296,N_42289);
nand U42613 (N_42613,N_42264,N_42310);
and U42614 (N_42614,N_42268,N_42329);
nand U42615 (N_42615,N_42371,N_42484);
and U42616 (N_42616,N_42297,N_42495);
nand U42617 (N_42617,N_42308,N_42269);
and U42618 (N_42618,N_42396,N_42456);
and U42619 (N_42619,N_42261,N_42258);
nor U42620 (N_42620,N_42497,N_42312);
and U42621 (N_42621,N_42356,N_42498);
xor U42622 (N_42622,N_42332,N_42273);
and U42623 (N_42623,N_42287,N_42472);
and U42624 (N_42624,N_42364,N_42251);
nor U42625 (N_42625,N_42477,N_42411);
nand U42626 (N_42626,N_42403,N_42323);
nor U42627 (N_42627,N_42425,N_42335);
or U42628 (N_42628,N_42409,N_42384);
xnor U42629 (N_42629,N_42323,N_42299);
and U42630 (N_42630,N_42272,N_42386);
xnor U42631 (N_42631,N_42326,N_42423);
nand U42632 (N_42632,N_42347,N_42439);
and U42633 (N_42633,N_42323,N_42473);
nand U42634 (N_42634,N_42393,N_42490);
nand U42635 (N_42635,N_42389,N_42384);
xnor U42636 (N_42636,N_42333,N_42389);
xor U42637 (N_42637,N_42409,N_42282);
nand U42638 (N_42638,N_42412,N_42270);
and U42639 (N_42639,N_42423,N_42394);
nand U42640 (N_42640,N_42373,N_42292);
xor U42641 (N_42641,N_42332,N_42368);
nand U42642 (N_42642,N_42381,N_42363);
and U42643 (N_42643,N_42294,N_42295);
nor U42644 (N_42644,N_42392,N_42352);
nor U42645 (N_42645,N_42425,N_42466);
and U42646 (N_42646,N_42266,N_42440);
or U42647 (N_42647,N_42276,N_42434);
or U42648 (N_42648,N_42371,N_42281);
nand U42649 (N_42649,N_42281,N_42380);
nor U42650 (N_42650,N_42305,N_42378);
and U42651 (N_42651,N_42356,N_42406);
or U42652 (N_42652,N_42258,N_42323);
xnor U42653 (N_42653,N_42496,N_42316);
nand U42654 (N_42654,N_42325,N_42481);
xnor U42655 (N_42655,N_42401,N_42476);
xnor U42656 (N_42656,N_42340,N_42343);
and U42657 (N_42657,N_42258,N_42442);
and U42658 (N_42658,N_42477,N_42373);
nor U42659 (N_42659,N_42299,N_42496);
xor U42660 (N_42660,N_42299,N_42462);
xor U42661 (N_42661,N_42287,N_42403);
or U42662 (N_42662,N_42382,N_42383);
or U42663 (N_42663,N_42359,N_42258);
nand U42664 (N_42664,N_42398,N_42290);
nand U42665 (N_42665,N_42402,N_42320);
nor U42666 (N_42666,N_42372,N_42336);
and U42667 (N_42667,N_42421,N_42491);
nor U42668 (N_42668,N_42298,N_42251);
nand U42669 (N_42669,N_42373,N_42429);
or U42670 (N_42670,N_42289,N_42414);
nor U42671 (N_42671,N_42352,N_42400);
xnor U42672 (N_42672,N_42262,N_42335);
nor U42673 (N_42673,N_42424,N_42275);
xor U42674 (N_42674,N_42340,N_42409);
and U42675 (N_42675,N_42448,N_42429);
nand U42676 (N_42676,N_42297,N_42368);
nor U42677 (N_42677,N_42386,N_42405);
or U42678 (N_42678,N_42353,N_42329);
nand U42679 (N_42679,N_42464,N_42373);
nor U42680 (N_42680,N_42280,N_42310);
nand U42681 (N_42681,N_42288,N_42461);
nand U42682 (N_42682,N_42428,N_42312);
nand U42683 (N_42683,N_42327,N_42485);
nor U42684 (N_42684,N_42352,N_42402);
nor U42685 (N_42685,N_42354,N_42281);
nor U42686 (N_42686,N_42490,N_42430);
or U42687 (N_42687,N_42482,N_42348);
or U42688 (N_42688,N_42453,N_42276);
nor U42689 (N_42689,N_42426,N_42340);
xor U42690 (N_42690,N_42390,N_42492);
xor U42691 (N_42691,N_42317,N_42258);
xor U42692 (N_42692,N_42390,N_42414);
or U42693 (N_42693,N_42480,N_42380);
xnor U42694 (N_42694,N_42331,N_42462);
xor U42695 (N_42695,N_42476,N_42425);
nand U42696 (N_42696,N_42315,N_42316);
nand U42697 (N_42697,N_42388,N_42401);
and U42698 (N_42698,N_42494,N_42269);
nand U42699 (N_42699,N_42339,N_42427);
or U42700 (N_42700,N_42278,N_42499);
xnor U42701 (N_42701,N_42493,N_42278);
nand U42702 (N_42702,N_42326,N_42414);
nor U42703 (N_42703,N_42435,N_42300);
nor U42704 (N_42704,N_42377,N_42300);
nand U42705 (N_42705,N_42467,N_42415);
or U42706 (N_42706,N_42318,N_42360);
nor U42707 (N_42707,N_42464,N_42317);
and U42708 (N_42708,N_42339,N_42489);
nand U42709 (N_42709,N_42396,N_42364);
nand U42710 (N_42710,N_42256,N_42354);
xor U42711 (N_42711,N_42411,N_42489);
and U42712 (N_42712,N_42294,N_42363);
nor U42713 (N_42713,N_42430,N_42493);
and U42714 (N_42714,N_42255,N_42369);
xnor U42715 (N_42715,N_42460,N_42401);
and U42716 (N_42716,N_42276,N_42414);
nand U42717 (N_42717,N_42255,N_42311);
nor U42718 (N_42718,N_42257,N_42295);
nor U42719 (N_42719,N_42306,N_42415);
nor U42720 (N_42720,N_42411,N_42383);
and U42721 (N_42721,N_42370,N_42396);
and U42722 (N_42722,N_42474,N_42445);
xnor U42723 (N_42723,N_42259,N_42349);
or U42724 (N_42724,N_42311,N_42338);
or U42725 (N_42725,N_42258,N_42426);
nor U42726 (N_42726,N_42417,N_42426);
or U42727 (N_42727,N_42442,N_42346);
nor U42728 (N_42728,N_42482,N_42408);
or U42729 (N_42729,N_42272,N_42490);
nor U42730 (N_42730,N_42478,N_42389);
nor U42731 (N_42731,N_42288,N_42255);
nand U42732 (N_42732,N_42263,N_42418);
and U42733 (N_42733,N_42438,N_42303);
or U42734 (N_42734,N_42252,N_42364);
and U42735 (N_42735,N_42349,N_42488);
and U42736 (N_42736,N_42403,N_42464);
and U42737 (N_42737,N_42444,N_42425);
or U42738 (N_42738,N_42339,N_42369);
nor U42739 (N_42739,N_42343,N_42336);
and U42740 (N_42740,N_42259,N_42406);
nor U42741 (N_42741,N_42298,N_42368);
nor U42742 (N_42742,N_42305,N_42260);
or U42743 (N_42743,N_42292,N_42265);
nor U42744 (N_42744,N_42299,N_42436);
and U42745 (N_42745,N_42321,N_42375);
xor U42746 (N_42746,N_42407,N_42476);
or U42747 (N_42747,N_42473,N_42406);
or U42748 (N_42748,N_42435,N_42277);
nand U42749 (N_42749,N_42375,N_42421);
xor U42750 (N_42750,N_42701,N_42514);
nor U42751 (N_42751,N_42713,N_42641);
xor U42752 (N_42752,N_42503,N_42560);
and U42753 (N_42753,N_42502,N_42591);
xor U42754 (N_42754,N_42516,N_42603);
nor U42755 (N_42755,N_42544,N_42570);
nor U42756 (N_42756,N_42558,N_42522);
and U42757 (N_42757,N_42517,N_42608);
nor U42758 (N_42758,N_42737,N_42590);
nand U42759 (N_42759,N_42524,N_42585);
and U42760 (N_42760,N_42647,N_42552);
nand U42761 (N_42761,N_42577,N_42664);
nor U42762 (N_42762,N_42661,N_42575);
xor U42763 (N_42763,N_42696,N_42732);
and U42764 (N_42764,N_42653,N_42512);
or U42765 (N_42765,N_42644,N_42735);
and U42766 (N_42766,N_42550,N_42574);
xnor U42767 (N_42767,N_42614,N_42506);
nor U42768 (N_42768,N_42563,N_42588);
or U42769 (N_42769,N_42626,N_42569);
or U42770 (N_42770,N_42722,N_42674);
and U42771 (N_42771,N_42625,N_42702);
nand U42772 (N_42772,N_42690,N_42704);
nor U42773 (N_42773,N_42685,N_42715);
or U42774 (N_42774,N_42509,N_42531);
nand U42775 (N_42775,N_42636,N_42745);
xnor U42776 (N_42776,N_42637,N_42673);
and U42777 (N_42777,N_42605,N_42688);
or U42778 (N_42778,N_42505,N_42707);
nand U42779 (N_42779,N_42589,N_42501);
nand U42780 (N_42780,N_42659,N_42683);
and U42781 (N_42781,N_42727,N_42621);
nor U42782 (N_42782,N_42518,N_42719);
or U42783 (N_42783,N_42557,N_42597);
or U42784 (N_42784,N_42733,N_42657);
and U42785 (N_42785,N_42547,N_42734);
or U42786 (N_42786,N_42576,N_42689);
and U42787 (N_42787,N_42533,N_42616);
xnor U42788 (N_42788,N_42643,N_42510);
and U42789 (N_42789,N_42692,N_42721);
or U42790 (N_42790,N_42526,N_42666);
nand U42791 (N_42791,N_42611,N_42743);
nand U42792 (N_42792,N_42622,N_42530);
nor U42793 (N_42793,N_42571,N_42619);
xnor U42794 (N_42794,N_42695,N_42698);
nand U42795 (N_42795,N_42573,N_42718);
nor U42796 (N_42796,N_42723,N_42596);
or U42797 (N_42797,N_42618,N_42545);
or U42798 (N_42798,N_42536,N_42598);
and U42799 (N_42799,N_42527,N_42740);
and U42800 (N_42800,N_42582,N_42671);
nor U42801 (N_42801,N_42546,N_42513);
and U42802 (N_42802,N_42584,N_42543);
or U42803 (N_42803,N_42746,N_42586);
nand U42804 (N_42804,N_42594,N_42520);
xor U42805 (N_42805,N_42508,N_42551);
or U42806 (N_42806,N_42649,N_42652);
nor U42807 (N_42807,N_42675,N_42720);
xnor U42808 (N_42808,N_42613,N_42628);
or U42809 (N_42809,N_42606,N_42642);
nor U42810 (N_42810,N_42748,N_42658);
nor U42811 (N_42811,N_42535,N_42581);
or U42812 (N_42812,N_42635,N_42583);
and U42813 (N_42813,N_42630,N_42744);
and U42814 (N_42814,N_42694,N_42724);
or U42815 (N_42815,N_42747,N_42580);
nor U42816 (N_42816,N_42554,N_42556);
xnor U42817 (N_42817,N_42665,N_42699);
or U42818 (N_42818,N_42629,N_42539);
or U42819 (N_42819,N_42525,N_42572);
or U42820 (N_42820,N_42578,N_42729);
or U42821 (N_42821,N_42549,N_42709);
or U42822 (N_42822,N_42739,N_42595);
xor U42823 (N_42823,N_42521,N_42602);
nor U42824 (N_42824,N_42725,N_42663);
or U42825 (N_42825,N_42679,N_42726);
xnor U42826 (N_42826,N_42529,N_42645);
xnor U42827 (N_42827,N_42631,N_42667);
and U42828 (N_42828,N_42601,N_42532);
or U42829 (N_42829,N_42691,N_42607);
nand U42830 (N_42830,N_42538,N_42681);
and U42831 (N_42831,N_42592,N_42623);
nand U42832 (N_42832,N_42676,N_42500);
and U42833 (N_42833,N_42749,N_42624);
or U42834 (N_42834,N_42656,N_42680);
xnor U42835 (N_42835,N_42738,N_42528);
xor U42836 (N_42836,N_42710,N_42627);
nor U42837 (N_42837,N_42615,N_42711);
nor U42838 (N_42838,N_42600,N_42730);
and U42839 (N_42839,N_42742,N_42678);
xnor U42840 (N_42840,N_42566,N_42634);
xor U42841 (N_42841,N_42617,N_42548);
or U42842 (N_42842,N_42677,N_42620);
xnor U42843 (N_42843,N_42537,N_42670);
or U42844 (N_42844,N_42610,N_42555);
and U42845 (N_42845,N_42651,N_42541);
nand U42846 (N_42846,N_42672,N_42736);
nand U42847 (N_42847,N_42639,N_42579);
nand U42848 (N_42848,N_42731,N_42638);
xor U42849 (N_42849,N_42504,N_42587);
xnor U42850 (N_42850,N_42741,N_42682);
xor U42851 (N_42851,N_42712,N_42612);
and U42852 (N_42852,N_42662,N_42559);
xor U42853 (N_42853,N_42604,N_42561);
or U42854 (N_42854,N_42717,N_42609);
or U42855 (N_42855,N_42593,N_42697);
or U42856 (N_42856,N_42599,N_42519);
xnor U42857 (N_42857,N_42716,N_42633);
nor U42858 (N_42858,N_42523,N_42669);
nand U42859 (N_42859,N_42540,N_42553);
and U42860 (N_42860,N_42660,N_42650);
and U42861 (N_42861,N_42686,N_42567);
xnor U42862 (N_42862,N_42646,N_42714);
and U42863 (N_42863,N_42511,N_42703);
nor U42864 (N_42864,N_42705,N_42515);
nor U42865 (N_42865,N_42562,N_42534);
xor U42866 (N_42866,N_42706,N_42708);
and U42867 (N_42867,N_42564,N_42542);
xnor U42868 (N_42868,N_42687,N_42640);
nand U42869 (N_42869,N_42684,N_42632);
or U42870 (N_42870,N_42700,N_42648);
xnor U42871 (N_42871,N_42693,N_42565);
nor U42872 (N_42872,N_42568,N_42668);
xor U42873 (N_42873,N_42728,N_42507);
nor U42874 (N_42874,N_42654,N_42655);
or U42875 (N_42875,N_42509,N_42576);
xor U42876 (N_42876,N_42530,N_42735);
nor U42877 (N_42877,N_42748,N_42504);
nand U42878 (N_42878,N_42714,N_42718);
xor U42879 (N_42879,N_42589,N_42701);
nand U42880 (N_42880,N_42516,N_42504);
or U42881 (N_42881,N_42611,N_42738);
and U42882 (N_42882,N_42561,N_42537);
and U42883 (N_42883,N_42587,N_42749);
nand U42884 (N_42884,N_42654,N_42650);
and U42885 (N_42885,N_42660,N_42673);
nor U42886 (N_42886,N_42733,N_42532);
nand U42887 (N_42887,N_42677,N_42517);
and U42888 (N_42888,N_42683,N_42707);
or U42889 (N_42889,N_42603,N_42748);
xor U42890 (N_42890,N_42692,N_42560);
and U42891 (N_42891,N_42726,N_42522);
xnor U42892 (N_42892,N_42744,N_42670);
and U42893 (N_42893,N_42696,N_42620);
xor U42894 (N_42894,N_42744,N_42501);
or U42895 (N_42895,N_42632,N_42609);
or U42896 (N_42896,N_42630,N_42626);
xor U42897 (N_42897,N_42518,N_42511);
and U42898 (N_42898,N_42629,N_42646);
xor U42899 (N_42899,N_42742,N_42581);
nor U42900 (N_42900,N_42733,N_42542);
or U42901 (N_42901,N_42745,N_42513);
and U42902 (N_42902,N_42507,N_42611);
nor U42903 (N_42903,N_42684,N_42642);
nand U42904 (N_42904,N_42674,N_42719);
xnor U42905 (N_42905,N_42747,N_42707);
xnor U42906 (N_42906,N_42574,N_42538);
nor U42907 (N_42907,N_42675,N_42672);
or U42908 (N_42908,N_42725,N_42579);
or U42909 (N_42909,N_42522,N_42641);
xor U42910 (N_42910,N_42749,N_42737);
xnor U42911 (N_42911,N_42618,N_42632);
or U42912 (N_42912,N_42539,N_42638);
nand U42913 (N_42913,N_42647,N_42571);
and U42914 (N_42914,N_42731,N_42600);
nand U42915 (N_42915,N_42609,N_42743);
nor U42916 (N_42916,N_42682,N_42534);
nand U42917 (N_42917,N_42612,N_42553);
xor U42918 (N_42918,N_42605,N_42580);
and U42919 (N_42919,N_42628,N_42563);
xor U42920 (N_42920,N_42579,N_42678);
and U42921 (N_42921,N_42586,N_42564);
xor U42922 (N_42922,N_42555,N_42613);
nor U42923 (N_42923,N_42678,N_42574);
nand U42924 (N_42924,N_42590,N_42523);
nor U42925 (N_42925,N_42729,N_42561);
nor U42926 (N_42926,N_42642,N_42670);
and U42927 (N_42927,N_42701,N_42711);
nor U42928 (N_42928,N_42640,N_42544);
or U42929 (N_42929,N_42708,N_42699);
or U42930 (N_42930,N_42686,N_42651);
or U42931 (N_42931,N_42747,N_42671);
nand U42932 (N_42932,N_42543,N_42572);
nand U42933 (N_42933,N_42612,N_42688);
nand U42934 (N_42934,N_42653,N_42537);
or U42935 (N_42935,N_42673,N_42511);
or U42936 (N_42936,N_42587,N_42598);
xnor U42937 (N_42937,N_42748,N_42595);
xnor U42938 (N_42938,N_42632,N_42692);
xnor U42939 (N_42939,N_42555,N_42622);
nor U42940 (N_42940,N_42698,N_42747);
and U42941 (N_42941,N_42637,N_42743);
xor U42942 (N_42942,N_42535,N_42748);
and U42943 (N_42943,N_42626,N_42656);
nor U42944 (N_42944,N_42513,N_42654);
xor U42945 (N_42945,N_42671,N_42564);
nand U42946 (N_42946,N_42631,N_42553);
and U42947 (N_42947,N_42723,N_42555);
nor U42948 (N_42948,N_42529,N_42567);
xor U42949 (N_42949,N_42681,N_42610);
or U42950 (N_42950,N_42602,N_42594);
nor U42951 (N_42951,N_42711,N_42515);
nand U42952 (N_42952,N_42523,N_42602);
and U42953 (N_42953,N_42659,N_42551);
nor U42954 (N_42954,N_42665,N_42634);
nand U42955 (N_42955,N_42606,N_42662);
nor U42956 (N_42956,N_42674,N_42630);
nand U42957 (N_42957,N_42605,N_42626);
nand U42958 (N_42958,N_42568,N_42660);
nand U42959 (N_42959,N_42748,N_42557);
xor U42960 (N_42960,N_42661,N_42745);
nand U42961 (N_42961,N_42541,N_42598);
nor U42962 (N_42962,N_42651,N_42502);
xnor U42963 (N_42963,N_42656,N_42577);
or U42964 (N_42964,N_42747,N_42591);
or U42965 (N_42965,N_42719,N_42503);
xnor U42966 (N_42966,N_42620,N_42690);
nand U42967 (N_42967,N_42670,N_42724);
xnor U42968 (N_42968,N_42573,N_42690);
nand U42969 (N_42969,N_42660,N_42599);
nor U42970 (N_42970,N_42599,N_42535);
and U42971 (N_42971,N_42670,N_42575);
xnor U42972 (N_42972,N_42623,N_42685);
xnor U42973 (N_42973,N_42736,N_42518);
nor U42974 (N_42974,N_42720,N_42627);
or U42975 (N_42975,N_42521,N_42543);
or U42976 (N_42976,N_42714,N_42734);
nand U42977 (N_42977,N_42659,N_42670);
and U42978 (N_42978,N_42700,N_42602);
and U42979 (N_42979,N_42564,N_42568);
or U42980 (N_42980,N_42724,N_42579);
nand U42981 (N_42981,N_42644,N_42673);
nor U42982 (N_42982,N_42517,N_42560);
nor U42983 (N_42983,N_42620,N_42603);
or U42984 (N_42984,N_42561,N_42670);
xnor U42985 (N_42985,N_42555,N_42712);
nor U42986 (N_42986,N_42714,N_42521);
or U42987 (N_42987,N_42666,N_42712);
xor U42988 (N_42988,N_42645,N_42741);
xnor U42989 (N_42989,N_42688,N_42717);
nand U42990 (N_42990,N_42654,N_42638);
xor U42991 (N_42991,N_42678,N_42697);
nand U42992 (N_42992,N_42682,N_42607);
nand U42993 (N_42993,N_42626,N_42551);
xnor U42994 (N_42994,N_42577,N_42517);
nand U42995 (N_42995,N_42571,N_42741);
or U42996 (N_42996,N_42696,N_42659);
nand U42997 (N_42997,N_42715,N_42679);
nand U42998 (N_42998,N_42535,N_42608);
nand U42999 (N_42999,N_42647,N_42664);
or U43000 (N_43000,N_42899,N_42843);
nand U43001 (N_43001,N_42814,N_42900);
nor U43002 (N_43002,N_42894,N_42992);
nor U43003 (N_43003,N_42880,N_42958);
or U43004 (N_43004,N_42953,N_42928);
nor U43005 (N_43005,N_42768,N_42811);
xnor U43006 (N_43006,N_42831,N_42872);
nand U43007 (N_43007,N_42927,N_42876);
or U43008 (N_43008,N_42881,N_42991);
nand U43009 (N_43009,N_42865,N_42918);
xor U43010 (N_43010,N_42751,N_42766);
xor U43011 (N_43011,N_42827,N_42837);
and U43012 (N_43012,N_42911,N_42804);
or U43013 (N_43013,N_42866,N_42920);
or U43014 (N_43014,N_42842,N_42966);
and U43015 (N_43015,N_42902,N_42965);
xnor U43016 (N_43016,N_42791,N_42940);
xnor U43017 (N_43017,N_42760,N_42964);
nand U43018 (N_43018,N_42956,N_42971);
xnor U43019 (N_43019,N_42807,N_42771);
nor U43020 (N_43020,N_42821,N_42785);
nand U43021 (N_43021,N_42945,N_42805);
xnor U43022 (N_43022,N_42912,N_42835);
or U43023 (N_43023,N_42803,N_42986);
nand U43024 (N_43024,N_42792,N_42759);
xnor U43025 (N_43025,N_42840,N_42937);
xor U43026 (N_43026,N_42952,N_42853);
nand U43027 (N_43027,N_42884,N_42955);
nor U43028 (N_43028,N_42801,N_42823);
nand U43029 (N_43029,N_42961,N_42769);
and U43030 (N_43030,N_42967,N_42977);
or U43031 (N_43031,N_42856,N_42779);
nor U43032 (N_43032,N_42995,N_42849);
xor U43033 (N_43033,N_42820,N_42931);
nand U43034 (N_43034,N_42948,N_42915);
and U43035 (N_43035,N_42926,N_42762);
or U43036 (N_43036,N_42999,N_42758);
or U43037 (N_43037,N_42822,N_42765);
xor U43038 (N_43038,N_42951,N_42947);
nand U43039 (N_43039,N_42802,N_42776);
nor U43040 (N_43040,N_42763,N_42979);
and U43041 (N_43041,N_42854,N_42809);
nor U43042 (N_43042,N_42824,N_42886);
nand U43043 (N_43043,N_42957,N_42816);
and U43044 (N_43044,N_42910,N_42845);
xor U43045 (N_43045,N_42929,N_42863);
xnor U43046 (N_43046,N_42753,N_42756);
nand U43047 (N_43047,N_42897,N_42846);
nor U43048 (N_43048,N_42901,N_42815);
xor U43049 (N_43049,N_42913,N_42808);
nor U43050 (N_43050,N_42941,N_42784);
and U43051 (N_43051,N_42806,N_42834);
or U43052 (N_43052,N_42851,N_42850);
and U43053 (N_43053,N_42954,N_42982);
nand U43054 (N_43054,N_42778,N_42869);
nand U43055 (N_43055,N_42825,N_42892);
nor U43056 (N_43056,N_42975,N_42819);
or U43057 (N_43057,N_42754,N_42794);
nand U43058 (N_43058,N_42859,N_42860);
xor U43059 (N_43059,N_42833,N_42962);
nand U43060 (N_43060,N_42848,N_42922);
nor U43061 (N_43061,N_42980,N_42755);
or U43062 (N_43062,N_42923,N_42875);
nand U43063 (N_43063,N_42960,N_42887);
or U43064 (N_43064,N_42963,N_42988);
nand U43065 (N_43065,N_42838,N_42878);
and U43066 (N_43066,N_42773,N_42861);
nor U43067 (N_43067,N_42883,N_42987);
nor U43068 (N_43068,N_42857,N_42930);
or U43069 (N_43069,N_42786,N_42997);
nand U43070 (N_43070,N_42906,N_42844);
or U43071 (N_43071,N_42890,N_42864);
nand U43072 (N_43072,N_42932,N_42788);
nor U43073 (N_43073,N_42767,N_42793);
xnor U43074 (N_43074,N_42873,N_42796);
xor U43075 (N_43075,N_42985,N_42798);
xor U43076 (N_43076,N_42830,N_42852);
and U43077 (N_43077,N_42959,N_42855);
xnor U43078 (N_43078,N_42950,N_42973);
or U43079 (N_43079,N_42917,N_42981);
nor U43080 (N_43080,N_42781,N_42871);
and U43081 (N_43081,N_42891,N_42797);
xor U43082 (N_43082,N_42974,N_42836);
or U43083 (N_43083,N_42944,N_42907);
or U43084 (N_43084,N_42895,N_42942);
nand U43085 (N_43085,N_42908,N_42904);
nand U43086 (N_43086,N_42764,N_42782);
xor U43087 (N_43087,N_42998,N_42970);
nand U43088 (N_43088,N_42777,N_42978);
xor U43089 (N_43089,N_42996,N_42934);
or U43090 (N_43090,N_42972,N_42896);
nand U43091 (N_43091,N_42832,N_42888);
nor U43092 (N_43092,N_42874,N_42924);
nand U43093 (N_43093,N_42817,N_42916);
nor U43094 (N_43094,N_42772,N_42770);
or U43095 (N_43095,N_42969,N_42829);
nand U43096 (N_43096,N_42885,N_42909);
and U43097 (N_43097,N_42990,N_42790);
and U43098 (N_43098,N_42752,N_42994);
and U43099 (N_43099,N_42905,N_42847);
or U43100 (N_43100,N_42946,N_42870);
nand U43101 (N_43101,N_42812,N_42877);
nor U43102 (N_43102,N_42789,N_42841);
and U43103 (N_43103,N_42810,N_42939);
or U43104 (N_43104,N_42935,N_42799);
xor U43105 (N_43105,N_42780,N_42976);
nor U43106 (N_43106,N_42949,N_42989);
or U43107 (N_43107,N_42867,N_42858);
or U43108 (N_43108,N_42893,N_42783);
nand U43109 (N_43109,N_42984,N_42795);
nor U43110 (N_43110,N_42813,N_42757);
or U43111 (N_43111,N_42775,N_42921);
nor U43112 (N_43112,N_42774,N_42839);
or U43113 (N_43113,N_42943,N_42914);
or U43114 (N_43114,N_42828,N_42879);
nor U43115 (N_43115,N_42968,N_42933);
nand U43116 (N_43116,N_42938,N_42868);
xor U43117 (N_43117,N_42983,N_42925);
or U43118 (N_43118,N_42818,N_42936);
or U43119 (N_43119,N_42919,N_42787);
xnor U43120 (N_43120,N_42898,N_42761);
and U43121 (N_43121,N_42826,N_42750);
and U43122 (N_43122,N_42800,N_42862);
and U43123 (N_43123,N_42882,N_42889);
or U43124 (N_43124,N_42993,N_42903);
and U43125 (N_43125,N_42876,N_42908);
and U43126 (N_43126,N_42867,N_42776);
nor U43127 (N_43127,N_42770,N_42857);
nand U43128 (N_43128,N_42859,N_42962);
and U43129 (N_43129,N_42834,N_42868);
xnor U43130 (N_43130,N_42801,N_42866);
nand U43131 (N_43131,N_42997,N_42896);
and U43132 (N_43132,N_42909,N_42870);
nand U43133 (N_43133,N_42780,N_42817);
nand U43134 (N_43134,N_42765,N_42887);
nand U43135 (N_43135,N_42759,N_42884);
nand U43136 (N_43136,N_42855,N_42991);
or U43137 (N_43137,N_42948,N_42776);
and U43138 (N_43138,N_42937,N_42923);
and U43139 (N_43139,N_42925,N_42778);
nor U43140 (N_43140,N_42826,N_42827);
xnor U43141 (N_43141,N_42797,N_42806);
xor U43142 (N_43142,N_42996,N_42842);
nand U43143 (N_43143,N_42883,N_42810);
nand U43144 (N_43144,N_42901,N_42810);
or U43145 (N_43145,N_42965,N_42886);
xnor U43146 (N_43146,N_42989,N_42872);
nor U43147 (N_43147,N_42781,N_42792);
nand U43148 (N_43148,N_42794,N_42830);
or U43149 (N_43149,N_42956,N_42830);
nor U43150 (N_43150,N_42839,N_42853);
or U43151 (N_43151,N_42857,N_42895);
nor U43152 (N_43152,N_42766,N_42902);
or U43153 (N_43153,N_42894,N_42961);
or U43154 (N_43154,N_42772,N_42895);
nor U43155 (N_43155,N_42866,N_42881);
and U43156 (N_43156,N_42903,N_42858);
or U43157 (N_43157,N_42829,N_42965);
or U43158 (N_43158,N_42916,N_42983);
and U43159 (N_43159,N_42953,N_42811);
or U43160 (N_43160,N_42812,N_42827);
and U43161 (N_43161,N_42896,N_42862);
or U43162 (N_43162,N_42801,N_42965);
or U43163 (N_43163,N_42884,N_42792);
or U43164 (N_43164,N_42885,N_42784);
or U43165 (N_43165,N_42923,N_42883);
nand U43166 (N_43166,N_42843,N_42975);
nor U43167 (N_43167,N_42847,N_42788);
nand U43168 (N_43168,N_42846,N_42805);
nor U43169 (N_43169,N_42869,N_42792);
xnor U43170 (N_43170,N_42888,N_42843);
nand U43171 (N_43171,N_42946,N_42770);
or U43172 (N_43172,N_42755,N_42995);
and U43173 (N_43173,N_42873,N_42967);
or U43174 (N_43174,N_42942,N_42809);
nor U43175 (N_43175,N_42752,N_42778);
nand U43176 (N_43176,N_42784,N_42923);
or U43177 (N_43177,N_42935,N_42878);
xnor U43178 (N_43178,N_42925,N_42901);
nor U43179 (N_43179,N_42979,N_42928);
nor U43180 (N_43180,N_42758,N_42799);
nand U43181 (N_43181,N_42762,N_42930);
xor U43182 (N_43182,N_42947,N_42975);
nor U43183 (N_43183,N_42772,N_42858);
nor U43184 (N_43184,N_42966,N_42869);
or U43185 (N_43185,N_42863,N_42835);
xor U43186 (N_43186,N_42941,N_42832);
or U43187 (N_43187,N_42991,N_42776);
nor U43188 (N_43188,N_42847,N_42926);
and U43189 (N_43189,N_42838,N_42764);
and U43190 (N_43190,N_42833,N_42873);
nand U43191 (N_43191,N_42999,N_42865);
and U43192 (N_43192,N_42963,N_42967);
and U43193 (N_43193,N_42798,N_42871);
nor U43194 (N_43194,N_42814,N_42854);
and U43195 (N_43195,N_42841,N_42979);
nand U43196 (N_43196,N_42984,N_42779);
and U43197 (N_43197,N_42870,N_42778);
xor U43198 (N_43198,N_42985,N_42864);
nor U43199 (N_43199,N_42981,N_42787);
nor U43200 (N_43200,N_42907,N_42792);
nor U43201 (N_43201,N_42809,N_42805);
nor U43202 (N_43202,N_42952,N_42808);
xor U43203 (N_43203,N_42977,N_42811);
xnor U43204 (N_43204,N_42755,N_42865);
and U43205 (N_43205,N_42915,N_42868);
nor U43206 (N_43206,N_42860,N_42910);
and U43207 (N_43207,N_42807,N_42803);
nand U43208 (N_43208,N_42981,N_42848);
or U43209 (N_43209,N_42906,N_42814);
nor U43210 (N_43210,N_42751,N_42926);
nor U43211 (N_43211,N_42935,N_42970);
nand U43212 (N_43212,N_42793,N_42896);
and U43213 (N_43213,N_42774,N_42818);
or U43214 (N_43214,N_42937,N_42949);
or U43215 (N_43215,N_42843,N_42976);
xnor U43216 (N_43216,N_42970,N_42828);
nand U43217 (N_43217,N_42853,N_42814);
xnor U43218 (N_43218,N_42928,N_42826);
xnor U43219 (N_43219,N_42962,N_42977);
xor U43220 (N_43220,N_42883,N_42831);
nor U43221 (N_43221,N_42993,N_42909);
nand U43222 (N_43222,N_42879,N_42799);
xnor U43223 (N_43223,N_42814,N_42760);
or U43224 (N_43224,N_42839,N_42967);
nand U43225 (N_43225,N_42986,N_42855);
nor U43226 (N_43226,N_42973,N_42891);
or U43227 (N_43227,N_42915,N_42831);
and U43228 (N_43228,N_42941,N_42773);
and U43229 (N_43229,N_42950,N_42787);
nor U43230 (N_43230,N_42798,N_42815);
nand U43231 (N_43231,N_42867,N_42894);
or U43232 (N_43232,N_42836,N_42866);
xnor U43233 (N_43233,N_42765,N_42894);
and U43234 (N_43234,N_42928,N_42984);
nand U43235 (N_43235,N_42756,N_42881);
and U43236 (N_43236,N_42842,N_42979);
xor U43237 (N_43237,N_42993,N_42834);
nor U43238 (N_43238,N_42917,N_42860);
nand U43239 (N_43239,N_42982,N_42757);
and U43240 (N_43240,N_42819,N_42801);
nand U43241 (N_43241,N_42865,N_42953);
or U43242 (N_43242,N_42905,N_42873);
or U43243 (N_43243,N_42943,N_42754);
xnor U43244 (N_43244,N_42764,N_42929);
or U43245 (N_43245,N_42997,N_42875);
xor U43246 (N_43246,N_42805,N_42888);
nor U43247 (N_43247,N_42917,N_42950);
and U43248 (N_43248,N_42849,N_42953);
xor U43249 (N_43249,N_42986,N_42976);
or U43250 (N_43250,N_43077,N_43194);
xor U43251 (N_43251,N_43097,N_43196);
xnor U43252 (N_43252,N_43092,N_43009);
or U43253 (N_43253,N_43018,N_43047);
or U43254 (N_43254,N_43023,N_43191);
nor U43255 (N_43255,N_43022,N_43099);
and U43256 (N_43256,N_43073,N_43039);
nand U43257 (N_43257,N_43007,N_43207);
nand U43258 (N_43258,N_43235,N_43110);
or U43259 (N_43259,N_43079,N_43029);
or U43260 (N_43260,N_43016,N_43143);
nand U43261 (N_43261,N_43100,N_43000);
xor U43262 (N_43262,N_43236,N_43122);
and U43263 (N_43263,N_43134,N_43213);
xor U43264 (N_43264,N_43121,N_43008);
xnor U43265 (N_43265,N_43206,N_43045);
nand U43266 (N_43266,N_43104,N_43169);
and U43267 (N_43267,N_43057,N_43050);
nand U43268 (N_43268,N_43135,N_43070);
nand U43269 (N_43269,N_43200,N_43202);
xnor U43270 (N_43270,N_43247,N_43037);
and U43271 (N_43271,N_43178,N_43132);
or U43272 (N_43272,N_43028,N_43127);
or U43273 (N_43273,N_43154,N_43003);
xnor U43274 (N_43274,N_43067,N_43102);
nor U43275 (N_43275,N_43190,N_43231);
xor U43276 (N_43276,N_43226,N_43056);
nand U43277 (N_43277,N_43150,N_43209);
nand U43278 (N_43278,N_43185,N_43128);
or U43279 (N_43279,N_43164,N_43064);
and U43280 (N_43280,N_43216,N_43068);
nand U43281 (N_43281,N_43225,N_43017);
or U43282 (N_43282,N_43245,N_43032);
and U43283 (N_43283,N_43218,N_43085);
and U43284 (N_43284,N_43118,N_43108);
nor U43285 (N_43285,N_43031,N_43229);
nand U43286 (N_43286,N_43220,N_43152);
or U43287 (N_43287,N_43239,N_43222);
nor U43288 (N_43288,N_43091,N_43112);
nor U43289 (N_43289,N_43042,N_43088);
nor U43290 (N_43290,N_43082,N_43111);
xor U43291 (N_43291,N_43205,N_43026);
nor U43292 (N_43292,N_43162,N_43227);
or U43293 (N_43293,N_43136,N_43014);
or U43294 (N_43294,N_43217,N_43172);
nor U43295 (N_43295,N_43188,N_43040);
xor U43296 (N_43296,N_43138,N_43025);
and U43297 (N_43297,N_43163,N_43147);
nor U43298 (N_43298,N_43033,N_43167);
or U43299 (N_43299,N_43180,N_43005);
or U43300 (N_43300,N_43192,N_43051);
nand U43301 (N_43301,N_43140,N_43210);
xor U43302 (N_43302,N_43001,N_43203);
xor U43303 (N_43303,N_43230,N_43090);
or U43304 (N_43304,N_43081,N_43105);
nand U43305 (N_43305,N_43193,N_43151);
nand U43306 (N_43306,N_43069,N_43024);
nor U43307 (N_43307,N_43123,N_43012);
or U43308 (N_43308,N_43228,N_43170);
nor U43309 (N_43309,N_43071,N_43242);
nand U43310 (N_43310,N_43197,N_43240);
and U43311 (N_43311,N_43093,N_43086);
xnor U43312 (N_43312,N_43211,N_43157);
xor U43313 (N_43313,N_43165,N_43249);
nand U43314 (N_43314,N_43019,N_43160);
nand U43315 (N_43315,N_43078,N_43149);
or U43316 (N_43316,N_43243,N_43189);
or U43317 (N_43317,N_43076,N_43098);
nand U43318 (N_43318,N_43199,N_43089);
nor U43319 (N_43319,N_43113,N_43015);
nor U43320 (N_43320,N_43043,N_43155);
xnor U43321 (N_43321,N_43248,N_43208);
nand U43322 (N_43322,N_43021,N_43195);
nor U43323 (N_43323,N_43141,N_43171);
xnor U43324 (N_43324,N_43133,N_43158);
nand U43325 (N_43325,N_43137,N_43139);
nor U43326 (N_43326,N_43062,N_43052);
xor U43327 (N_43327,N_43101,N_43186);
nand U43328 (N_43328,N_43166,N_43130);
nand U43329 (N_43329,N_43221,N_43212);
nand U43330 (N_43330,N_43030,N_43087);
nor U43331 (N_43331,N_43116,N_43041);
and U43332 (N_43332,N_43115,N_43187);
nor U43333 (N_43333,N_43125,N_43006);
and U43334 (N_43334,N_43074,N_43198);
nor U43335 (N_43335,N_43013,N_43219);
or U43336 (N_43336,N_43061,N_43044);
xnor U43337 (N_43337,N_43053,N_43144);
nor U43338 (N_43338,N_43106,N_43124);
nand U43339 (N_43339,N_43060,N_43103);
nand U43340 (N_43340,N_43145,N_43177);
nand U43341 (N_43341,N_43224,N_43027);
or U43342 (N_43342,N_43084,N_43004);
nand U43343 (N_43343,N_43204,N_43038);
and U43344 (N_43344,N_43072,N_43054);
nor U43345 (N_43345,N_43049,N_43010);
nor U43346 (N_43346,N_43036,N_43168);
xor U43347 (N_43347,N_43035,N_43159);
or U43348 (N_43348,N_43119,N_43034);
nor U43349 (N_43349,N_43181,N_43094);
nand U43350 (N_43350,N_43153,N_43129);
and U43351 (N_43351,N_43179,N_43232);
and U43352 (N_43352,N_43002,N_43215);
xnor U43353 (N_43353,N_43246,N_43184);
xnor U43354 (N_43354,N_43182,N_43146);
or U43355 (N_43355,N_43059,N_43065);
xor U43356 (N_43356,N_43048,N_43055);
and U43357 (N_43357,N_43096,N_43075);
nand U43358 (N_43358,N_43080,N_43083);
xor U43359 (N_43359,N_43063,N_43120);
nor U43360 (N_43360,N_43095,N_43201);
xnor U43361 (N_43361,N_43233,N_43142);
and U43362 (N_43362,N_43173,N_43131);
or U43363 (N_43363,N_43237,N_43244);
xor U43364 (N_43364,N_43176,N_43241);
nand U43365 (N_43365,N_43156,N_43114);
or U43366 (N_43366,N_43020,N_43175);
nand U43367 (N_43367,N_43011,N_43234);
and U43368 (N_43368,N_43126,N_43107);
nor U43369 (N_43369,N_43148,N_43066);
or U43370 (N_43370,N_43109,N_43117);
xor U43371 (N_43371,N_43174,N_43161);
or U43372 (N_43372,N_43223,N_43058);
and U43373 (N_43373,N_43214,N_43238);
nor U43374 (N_43374,N_43183,N_43046);
or U43375 (N_43375,N_43173,N_43110);
or U43376 (N_43376,N_43126,N_43247);
nand U43377 (N_43377,N_43054,N_43139);
nand U43378 (N_43378,N_43097,N_43030);
or U43379 (N_43379,N_43168,N_43165);
nor U43380 (N_43380,N_43177,N_43234);
or U43381 (N_43381,N_43001,N_43085);
nor U43382 (N_43382,N_43221,N_43227);
nor U43383 (N_43383,N_43209,N_43219);
or U43384 (N_43384,N_43034,N_43132);
or U43385 (N_43385,N_43039,N_43108);
nand U43386 (N_43386,N_43126,N_43013);
and U43387 (N_43387,N_43169,N_43033);
nor U43388 (N_43388,N_43004,N_43130);
and U43389 (N_43389,N_43195,N_43169);
xnor U43390 (N_43390,N_43002,N_43114);
xnor U43391 (N_43391,N_43207,N_43101);
and U43392 (N_43392,N_43216,N_43187);
or U43393 (N_43393,N_43063,N_43180);
nor U43394 (N_43394,N_43183,N_43211);
or U43395 (N_43395,N_43191,N_43211);
nor U43396 (N_43396,N_43071,N_43227);
or U43397 (N_43397,N_43057,N_43239);
xor U43398 (N_43398,N_43091,N_43021);
xor U43399 (N_43399,N_43157,N_43215);
xor U43400 (N_43400,N_43019,N_43117);
and U43401 (N_43401,N_43212,N_43033);
or U43402 (N_43402,N_43095,N_43247);
nor U43403 (N_43403,N_43015,N_43143);
nand U43404 (N_43404,N_43225,N_43115);
or U43405 (N_43405,N_43201,N_43118);
nand U43406 (N_43406,N_43223,N_43206);
nor U43407 (N_43407,N_43116,N_43192);
nand U43408 (N_43408,N_43022,N_43089);
xnor U43409 (N_43409,N_43200,N_43214);
nor U43410 (N_43410,N_43245,N_43005);
and U43411 (N_43411,N_43206,N_43180);
xnor U43412 (N_43412,N_43114,N_43216);
nor U43413 (N_43413,N_43047,N_43128);
or U43414 (N_43414,N_43129,N_43010);
or U43415 (N_43415,N_43155,N_43137);
nor U43416 (N_43416,N_43183,N_43004);
xor U43417 (N_43417,N_43207,N_43099);
and U43418 (N_43418,N_43149,N_43033);
or U43419 (N_43419,N_43189,N_43187);
and U43420 (N_43420,N_43127,N_43163);
xor U43421 (N_43421,N_43081,N_43055);
xor U43422 (N_43422,N_43015,N_43058);
nor U43423 (N_43423,N_43197,N_43208);
xnor U43424 (N_43424,N_43009,N_43061);
nand U43425 (N_43425,N_43233,N_43104);
xor U43426 (N_43426,N_43020,N_43192);
nor U43427 (N_43427,N_43211,N_43001);
xor U43428 (N_43428,N_43135,N_43168);
and U43429 (N_43429,N_43179,N_43022);
or U43430 (N_43430,N_43103,N_43210);
nor U43431 (N_43431,N_43045,N_43066);
xnor U43432 (N_43432,N_43104,N_43058);
nand U43433 (N_43433,N_43146,N_43225);
nor U43434 (N_43434,N_43204,N_43033);
or U43435 (N_43435,N_43124,N_43125);
or U43436 (N_43436,N_43213,N_43095);
xnor U43437 (N_43437,N_43102,N_43104);
xnor U43438 (N_43438,N_43174,N_43180);
nor U43439 (N_43439,N_43043,N_43190);
nor U43440 (N_43440,N_43166,N_43086);
or U43441 (N_43441,N_43113,N_43190);
nand U43442 (N_43442,N_43098,N_43050);
and U43443 (N_43443,N_43158,N_43217);
and U43444 (N_43444,N_43237,N_43222);
nor U43445 (N_43445,N_43031,N_43096);
nand U43446 (N_43446,N_43123,N_43105);
and U43447 (N_43447,N_43196,N_43035);
nand U43448 (N_43448,N_43128,N_43203);
xnor U43449 (N_43449,N_43230,N_43049);
or U43450 (N_43450,N_43026,N_43050);
xor U43451 (N_43451,N_43096,N_43062);
nand U43452 (N_43452,N_43105,N_43210);
and U43453 (N_43453,N_43118,N_43085);
and U43454 (N_43454,N_43055,N_43122);
nor U43455 (N_43455,N_43127,N_43043);
nor U43456 (N_43456,N_43066,N_43237);
nor U43457 (N_43457,N_43234,N_43030);
and U43458 (N_43458,N_43202,N_43215);
nand U43459 (N_43459,N_43115,N_43218);
or U43460 (N_43460,N_43091,N_43144);
nand U43461 (N_43461,N_43152,N_43136);
nand U43462 (N_43462,N_43132,N_43138);
xnor U43463 (N_43463,N_43244,N_43133);
and U43464 (N_43464,N_43233,N_43156);
or U43465 (N_43465,N_43226,N_43141);
nor U43466 (N_43466,N_43059,N_43159);
nand U43467 (N_43467,N_43236,N_43108);
nor U43468 (N_43468,N_43054,N_43129);
and U43469 (N_43469,N_43057,N_43074);
xnor U43470 (N_43470,N_43240,N_43090);
and U43471 (N_43471,N_43055,N_43217);
nand U43472 (N_43472,N_43129,N_43182);
xor U43473 (N_43473,N_43014,N_43201);
or U43474 (N_43474,N_43080,N_43010);
xnor U43475 (N_43475,N_43047,N_43161);
nand U43476 (N_43476,N_43244,N_43165);
and U43477 (N_43477,N_43103,N_43003);
or U43478 (N_43478,N_43186,N_43191);
nor U43479 (N_43479,N_43186,N_43066);
xnor U43480 (N_43480,N_43132,N_43187);
nor U43481 (N_43481,N_43166,N_43033);
nand U43482 (N_43482,N_43117,N_43113);
and U43483 (N_43483,N_43211,N_43153);
xnor U43484 (N_43484,N_43114,N_43226);
xor U43485 (N_43485,N_43130,N_43005);
or U43486 (N_43486,N_43188,N_43072);
or U43487 (N_43487,N_43232,N_43071);
xnor U43488 (N_43488,N_43081,N_43086);
nor U43489 (N_43489,N_43002,N_43225);
and U43490 (N_43490,N_43064,N_43092);
xor U43491 (N_43491,N_43005,N_43020);
or U43492 (N_43492,N_43019,N_43116);
and U43493 (N_43493,N_43221,N_43202);
xnor U43494 (N_43494,N_43168,N_43180);
and U43495 (N_43495,N_43213,N_43031);
xnor U43496 (N_43496,N_43191,N_43081);
nand U43497 (N_43497,N_43202,N_43166);
xor U43498 (N_43498,N_43164,N_43166);
nor U43499 (N_43499,N_43084,N_43056);
xnor U43500 (N_43500,N_43430,N_43429);
xnor U43501 (N_43501,N_43297,N_43257);
nor U43502 (N_43502,N_43404,N_43280);
nand U43503 (N_43503,N_43323,N_43364);
xor U43504 (N_43504,N_43326,N_43313);
and U43505 (N_43505,N_43450,N_43361);
xnor U43506 (N_43506,N_43425,N_43387);
or U43507 (N_43507,N_43262,N_43273);
nor U43508 (N_43508,N_43264,N_43274);
nor U43509 (N_43509,N_43296,N_43325);
nor U43510 (N_43510,N_43479,N_43362);
nand U43511 (N_43511,N_43435,N_43254);
and U43512 (N_43512,N_43339,N_43345);
nand U43513 (N_43513,N_43336,N_43371);
nand U43514 (N_43514,N_43347,N_43454);
or U43515 (N_43515,N_43488,N_43443);
xor U43516 (N_43516,N_43487,N_43286);
nor U43517 (N_43517,N_43298,N_43401);
xor U43518 (N_43518,N_43394,N_43341);
nor U43519 (N_43519,N_43373,N_43418);
nor U43520 (N_43520,N_43363,N_43400);
or U43521 (N_43521,N_43481,N_43492);
xor U43522 (N_43522,N_43285,N_43259);
and U43523 (N_43523,N_43374,N_43300);
and U43524 (N_43524,N_43303,N_43448);
xor U43525 (N_43525,N_43301,N_43388);
nor U43526 (N_43526,N_43456,N_43485);
or U43527 (N_43527,N_43310,N_43459);
or U43528 (N_43528,N_43306,N_43496);
and U43529 (N_43529,N_43270,N_43294);
nand U43530 (N_43530,N_43390,N_43399);
xnor U43531 (N_43531,N_43383,N_43366);
or U43532 (N_43532,N_43252,N_43447);
nor U43533 (N_43533,N_43403,N_43410);
xnor U43534 (N_43534,N_43276,N_43378);
xor U43535 (N_43535,N_43382,N_43379);
and U43536 (N_43536,N_43369,N_43269);
and U43537 (N_43537,N_43266,N_43398);
and U43538 (N_43538,N_43486,N_43337);
or U43539 (N_43539,N_43291,N_43320);
nand U43540 (N_43540,N_43489,N_43389);
or U43541 (N_43541,N_43474,N_43302);
or U43542 (N_43542,N_43287,N_43455);
nand U43543 (N_43543,N_43427,N_43331);
xor U43544 (N_43544,N_43472,N_43497);
xnor U43545 (N_43545,N_43463,N_43289);
and U43546 (N_43546,N_43426,N_43278);
xnor U43547 (N_43547,N_43412,N_43392);
nand U43548 (N_43548,N_43368,N_43370);
nor U43549 (N_43549,N_43295,N_43438);
and U43550 (N_43550,N_43355,N_43255);
nor U43551 (N_43551,N_43338,N_43475);
or U43552 (N_43552,N_43309,N_43340);
nand U43553 (N_43553,N_43346,N_43367);
or U43554 (N_43554,N_43490,N_43308);
or U43555 (N_43555,N_43316,N_43359);
xnor U43556 (N_43556,N_43372,N_43250);
and U43557 (N_43557,N_43439,N_43495);
or U43558 (N_43558,N_43491,N_43258);
xnor U43559 (N_43559,N_43482,N_43436);
xnor U43560 (N_43560,N_43396,N_43350);
and U43561 (N_43561,N_43432,N_43253);
nand U43562 (N_43562,N_43263,N_43360);
nand U43563 (N_43563,N_43466,N_43413);
and U43564 (N_43564,N_43480,N_43380);
xor U43565 (N_43565,N_43422,N_43424);
xnor U43566 (N_43566,N_43330,N_43256);
nand U43567 (N_43567,N_43282,N_43344);
nor U43568 (N_43568,N_43445,N_43444);
nor U43569 (N_43569,N_43470,N_43415);
xnor U43570 (N_43570,N_43292,N_43493);
nand U43571 (N_43571,N_43469,N_43460);
nand U43572 (N_43572,N_43411,N_43277);
or U43573 (N_43573,N_43483,N_43329);
or U43574 (N_43574,N_43408,N_43377);
nand U43575 (N_43575,N_43420,N_43304);
nand U43576 (N_43576,N_43423,N_43381);
or U43577 (N_43577,N_43334,N_43314);
nor U43578 (N_43578,N_43484,N_43284);
xor U43579 (N_43579,N_43461,N_43275);
nand U43580 (N_43580,N_43321,N_43307);
nand U43581 (N_43581,N_43452,N_43349);
nor U43582 (N_43582,N_43288,N_43499);
or U43583 (N_43583,N_43332,N_43356);
and U43584 (N_43584,N_43305,N_43437);
and U43585 (N_43585,N_43342,N_43406);
and U43586 (N_43586,N_43402,N_43417);
and U43587 (N_43587,N_43440,N_43414);
and U43588 (N_43588,N_43281,N_43421);
nor U43589 (N_43589,N_43376,N_43317);
or U43590 (N_43590,N_43434,N_43467);
nand U43591 (N_43591,N_43409,N_43328);
nand U43592 (N_43592,N_43449,N_43272);
nor U43593 (N_43593,N_43462,N_43384);
xor U43594 (N_43594,N_43283,N_43293);
nor U43595 (N_43595,N_43494,N_43419);
xor U43596 (N_43596,N_43318,N_43375);
and U43597 (N_43597,N_43457,N_43268);
or U43598 (N_43598,N_43476,N_43385);
and U43599 (N_43599,N_43267,N_43279);
xor U43600 (N_43600,N_43351,N_43290);
nor U43601 (N_43601,N_43431,N_43324);
nor U43602 (N_43602,N_43498,N_43464);
nor U43603 (N_43603,N_43433,N_43442);
nor U43604 (N_43604,N_43251,N_43343);
or U43605 (N_43605,N_43319,N_43333);
nor U43606 (N_43606,N_43458,N_43478);
nand U43607 (N_43607,N_43477,N_43465);
xor U43608 (N_43608,N_43451,N_43416);
nand U43609 (N_43609,N_43358,N_43327);
and U43610 (N_43610,N_43299,N_43261);
nand U43611 (N_43611,N_43428,N_43395);
or U43612 (N_43612,N_43386,N_43271);
xnor U43613 (N_43613,N_43311,N_43353);
and U43614 (N_43614,N_43393,N_43354);
xnor U43615 (N_43615,N_43397,N_43365);
nor U43616 (N_43616,N_43391,N_43260);
nor U43617 (N_43617,N_43335,N_43441);
nor U43618 (N_43618,N_43315,N_43265);
nand U43619 (N_43619,N_43312,N_43357);
nand U43620 (N_43620,N_43407,N_43473);
nand U43621 (N_43621,N_43352,N_43468);
xor U43622 (N_43622,N_43348,N_43453);
nor U43623 (N_43623,N_43405,N_43471);
xor U43624 (N_43624,N_43446,N_43322);
or U43625 (N_43625,N_43450,N_43475);
nor U43626 (N_43626,N_43284,N_43397);
and U43627 (N_43627,N_43468,N_43415);
nand U43628 (N_43628,N_43426,N_43285);
nor U43629 (N_43629,N_43416,N_43299);
and U43630 (N_43630,N_43416,N_43469);
nor U43631 (N_43631,N_43455,N_43341);
xor U43632 (N_43632,N_43479,N_43296);
and U43633 (N_43633,N_43344,N_43414);
xor U43634 (N_43634,N_43420,N_43400);
nand U43635 (N_43635,N_43343,N_43319);
nand U43636 (N_43636,N_43387,N_43354);
nand U43637 (N_43637,N_43467,N_43398);
or U43638 (N_43638,N_43458,N_43477);
or U43639 (N_43639,N_43346,N_43330);
nand U43640 (N_43640,N_43462,N_43467);
and U43641 (N_43641,N_43350,N_43433);
and U43642 (N_43642,N_43312,N_43446);
nor U43643 (N_43643,N_43374,N_43309);
or U43644 (N_43644,N_43320,N_43350);
nor U43645 (N_43645,N_43380,N_43389);
and U43646 (N_43646,N_43366,N_43448);
nand U43647 (N_43647,N_43462,N_43470);
nand U43648 (N_43648,N_43421,N_43398);
nand U43649 (N_43649,N_43422,N_43357);
xnor U43650 (N_43650,N_43304,N_43410);
nand U43651 (N_43651,N_43388,N_43355);
and U43652 (N_43652,N_43493,N_43460);
and U43653 (N_43653,N_43322,N_43342);
and U43654 (N_43654,N_43372,N_43396);
nand U43655 (N_43655,N_43496,N_43454);
nor U43656 (N_43656,N_43340,N_43473);
or U43657 (N_43657,N_43491,N_43260);
nand U43658 (N_43658,N_43443,N_43397);
nor U43659 (N_43659,N_43401,N_43256);
xor U43660 (N_43660,N_43440,N_43497);
xor U43661 (N_43661,N_43430,N_43258);
nor U43662 (N_43662,N_43286,N_43377);
nand U43663 (N_43663,N_43257,N_43365);
xnor U43664 (N_43664,N_43485,N_43449);
xor U43665 (N_43665,N_43345,N_43253);
nor U43666 (N_43666,N_43283,N_43435);
nor U43667 (N_43667,N_43473,N_43288);
xnor U43668 (N_43668,N_43359,N_43498);
or U43669 (N_43669,N_43270,N_43494);
and U43670 (N_43670,N_43334,N_43493);
nand U43671 (N_43671,N_43480,N_43344);
and U43672 (N_43672,N_43378,N_43410);
xnor U43673 (N_43673,N_43260,N_43363);
and U43674 (N_43674,N_43372,N_43296);
or U43675 (N_43675,N_43341,N_43283);
xor U43676 (N_43676,N_43481,N_43280);
and U43677 (N_43677,N_43477,N_43474);
nand U43678 (N_43678,N_43379,N_43448);
xor U43679 (N_43679,N_43250,N_43374);
xnor U43680 (N_43680,N_43265,N_43409);
or U43681 (N_43681,N_43471,N_43439);
nand U43682 (N_43682,N_43266,N_43324);
nor U43683 (N_43683,N_43391,N_43291);
xor U43684 (N_43684,N_43352,N_43336);
nor U43685 (N_43685,N_43439,N_43300);
nand U43686 (N_43686,N_43252,N_43437);
and U43687 (N_43687,N_43442,N_43376);
xnor U43688 (N_43688,N_43278,N_43286);
and U43689 (N_43689,N_43464,N_43454);
nor U43690 (N_43690,N_43366,N_43375);
nor U43691 (N_43691,N_43270,N_43362);
nor U43692 (N_43692,N_43262,N_43376);
nand U43693 (N_43693,N_43267,N_43403);
nand U43694 (N_43694,N_43439,N_43467);
or U43695 (N_43695,N_43276,N_43327);
nand U43696 (N_43696,N_43383,N_43352);
nand U43697 (N_43697,N_43488,N_43284);
and U43698 (N_43698,N_43286,N_43420);
nand U43699 (N_43699,N_43379,N_43397);
and U43700 (N_43700,N_43366,N_43374);
xor U43701 (N_43701,N_43271,N_43260);
or U43702 (N_43702,N_43253,N_43419);
nand U43703 (N_43703,N_43400,N_43307);
or U43704 (N_43704,N_43456,N_43438);
and U43705 (N_43705,N_43445,N_43377);
nand U43706 (N_43706,N_43252,N_43361);
nor U43707 (N_43707,N_43409,N_43295);
nor U43708 (N_43708,N_43366,N_43263);
nand U43709 (N_43709,N_43344,N_43359);
or U43710 (N_43710,N_43386,N_43412);
nor U43711 (N_43711,N_43312,N_43362);
nand U43712 (N_43712,N_43387,N_43410);
and U43713 (N_43713,N_43388,N_43308);
and U43714 (N_43714,N_43462,N_43352);
xor U43715 (N_43715,N_43281,N_43418);
nor U43716 (N_43716,N_43456,N_43385);
nor U43717 (N_43717,N_43253,N_43258);
or U43718 (N_43718,N_43485,N_43371);
or U43719 (N_43719,N_43335,N_43454);
or U43720 (N_43720,N_43435,N_43300);
and U43721 (N_43721,N_43397,N_43277);
nor U43722 (N_43722,N_43382,N_43401);
xor U43723 (N_43723,N_43491,N_43410);
nand U43724 (N_43724,N_43476,N_43253);
xor U43725 (N_43725,N_43427,N_43311);
or U43726 (N_43726,N_43289,N_43499);
nor U43727 (N_43727,N_43350,N_43445);
xnor U43728 (N_43728,N_43352,N_43452);
xor U43729 (N_43729,N_43451,N_43288);
nor U43730 (N_43730,N_43332,N_43252);
xnor U43731 (N_43731,N_43323,N_43265);
and U43732 (N_43732,N_43481,N_43269);
nand U43733 (N_43733,N_43423,N_43352);
and U43734 (N_43734,N_43364,N_43337);
or U43735 (N_43735,N_43383,N_43411);
xnor U43736 (N_43736,N_43453,N_43381);
nand U43737 (N_43737,N_43254,N_43278);
xnor U43738 (N_43738,N_43344,N_43494);
and U43739 (N_43739,N_43397,N_43399);
nand U43740 (N_43740,N_43409,N_43393);
nand U43741 (N_43741,N_43279,N_43290);
nand U43742 (N_43742,N_43481,N_43419);
nand U43743 (N_43743,N_43252,N_43434);
nand U43744 (N_43744,N_43370,N_43469);
or U43745 (N_43745,N_43328,N_43250);
or U43746 (N_43746,N_43431,N_43291);
nand U43747 (N_43747,N_43256,N_43369);
nor U43748 (N_43748,N_43354,N_43279);
xor U43749 (N_43749,N_43449,N_43331);
or U43750 (N_43750,N_43749,N_43677);
or U43751 (N_43751,N_43687,N_43563);
nand U43752 (N_43752,N_43531,N_43686);
nor U43753 (N_43753,N_43701,N_43676);
nand U43754 (N_43754,N_43655,N_43746);
and U43755 (N_43755,N_43748,N_43736);
and U43756 (N_43756,N_43707,N_43501);
nand U43757 (N_43757,N_43550,N_43688);
or U43758 (N_43758,N_43595,N_43647);
xnor U43759 (N_43759,N_43747,N_43740);
nand U43760 (N_43760,N_43510,N_43540);
and U43761 (N_43761,N_43502,N_43616);
nor U43762 (N_43762,N_43671,N_43633);
xnor U43763 (N_43763,N_43567,N_43523);
xor U43764 (N_43764,N_43560,N_43737);
nor U43765 (N_43765,N_43685,N_43675);
xor U43766 (N_43766,N_43614,N_43646);
nand U43767 (N_43767,N_43511,N_43704);
xor U43768 (N_43768,N_43537,N_43706);
xnor U43769 (N_43769,N_43732,N_43515);
nor U43770 (N_43770,N_43582,N_43738);
and U43771 (N_43771,N_43645,N_43679);
nor U43772 (N_43772,N_43503,N_43564);
nor U43773 (N_43773,N_43624,N_43702);
xor U43774 (N_43774,N_43589,N_43545);
nand U43775 (N_43775,N_43650,N_43699);
nand U43776 (N_43776,N_43553,N_43673);
xnor U43777 (N_43777,N_43509,N_43657);
nor U43778 (N_43778,N_43678,N_43535);
nand U43779 (N_43779,N_43727,N_43713);
nor U43780 (N_43780,N_43720,N_43573);
or U43781 (N_43781,N_43725,N_43506);
xnor U43782 (N_43782,N_43643,N_43716);
nor U43783 (N_43783,N_43741,N_43734);
nand U43784 (N_43784,N_43682,N_43692);
and U43785 (N_43785,N_43583,N_43665);
or U43786 (N_43786,N_43521,N_43565);
or U43787 (N_43787,N_43551,N_43705);
or U43788 (N_43788,N_43592,N_43630);
xnor U43789 (N_43789,N_43568,N_43575);
or U43790 (N_43790,N_43680,N_43556);
nand U43791 (N_43791,N_43541,N_43543);
nand U43792 (N_43792,N_43638,N_43651);
xnor U43793 (N_43793,N_43632,N_43598);
nor U43794 (N_43794,N_43518,N_43526);
nor U43795 (N_43795,N_43662,N_43661);
and U43796 (N_43796,N_43695,N_43513);
and U43797 (N_43797,N_43697,N_43533);
xnor U43798 (N_43798,N_43609,N_43528);
nor U43799 (N_43799,N_43664,N_43618);
xor U43800 (N_43800,N_43619,N_43538);
and U43801 (N_43801,N_43574,N_43718);
nor U43802 (N_43802,N_43532,N_43605);
nand U43803 (N_43803,N_43731,N_43539);
or U43804 (N_43804,N_43585,N_43683);
nand U43805 (N_43805,N_43708,N_43656);
and U43806 (N_43806,N_43508,N_43729);
xnor U43807 (N_43807,N_43591,N_43622);
or U43808 (N_43808,N_43612,N_43627);
or U43809 (N_43809,N_43636,N_43519);
or U43810 (N_43810,N_43691,N_43660);
nand U43811 (N_43811,N_43654,N_43681);
nor U43812 (N_43812,N_43640,N_43613);
nor U43813 (N_43813,N_43607,N_43653);
and U43814 (N_43814,N_43674,N_43733);
and U43815 (N_43815,N_43649,N_43709);
nor U43816 (N_43816,N_43621,N_43599);
nor U43817 (N_43817,N_43626,N_43536);
xnor U43818 (N_43818,N_43608,N_43711);
and U43819 (N_43819,N_43712,N_43668);
or U43820 (N_43820,N_43667,N_43505);
xnor U43821 (N_43821,N_43500,N_43586);
nor U43822 (N_43822,N_43610,N_43672);
xor U43823 (N_43823,N_43641,N_43617);
and U43824 (N_43824,N_43517,N_43611);
or U43825 (N_43825,N_43724,N_43639);
xnor U43826 (N_43826,N_43512,N_43594);
or U43827 (N_43827,N_43570,N_43557);
nor U43828 (N_43828,N_43558,N_43615);
nor U43829 (N_43829,N_43603,N_43700);
or U43830 (N_43830,N_43745,N_43717);
and U43831 (N_43831,N_43684,N_43588);
and U43832 (N_43832,N_43690,N_43659);
and U43833 (N_43833,N_43530,N_43590);
xnor U43834 (N_43834,N_43620,N_43730);
and U43835 (N_43835,N_43559,N_43549);
xor U43836 (N_43836,N_43669,N_43721);
xnor U43837 (N_43837,N_43652,N_43555);
nor U43838 (N_43838,N_43584,N_43743);
xnor U43839 (N_43839,N_43561,N_43593);
and U43840 (N_43840,N_43623,N_43648);
or U43841 (N_43841,N_43693,N_43628);
or U43842 (N_43842,N_43597,N_43542);
nor U43843 (N_43843,N_43714,N_43689);
and U43844 (N_43844,N_43602,N_43739);
nor U43845 (N_43845,N_43587,N_43663);
or U43846 (N_43846,N_43723,N_43744);
nand U43847 (N_43847,N_43520,N_43572);
or U43848 (N_43848,N_43534,N_43722);
or U43849 (N_43849,N_43554,N_43562);
and U43850 (N_43850,N_43634,N_43596);
xnor U43851 (N_43851,N_43703,N_43698);
and U43852 (N_43852,N_43576,N_43529);
or U43853 (N_43853,N_43569,N_43525);
nor U43854 (N_43854,N_43524,N_43742);
nand U43855 (N_43855,N_43637,N_43600);
xor U43856 (N_43856,N_43566,N_43544);
xor U43857 (N_43857,N_43670,N_43735);
nand U43858 (N_43858,N_43516,N_43546);
xor U43859 (N_43859,N_43552,N_43547);
nor U43860 (N_43860,N_43631,N_43696);
nand U43861 (N_43861,N_43625,N_43577);
and U43862 (N_43862,N_43710,N_43715);
and U43863 (N_43863,N_43635,N_43606);
and U43864 (N_43864,N_43629,N_43522);
nor U43865 (N_43865,N_43726,N_43642);
and U43866 (N_43866,N_43548,N_43719);
nor U43867 (N_43867,N_43644,N_43571);
or U43868 (N_43868,N_43580,N_43666);
and U43869 (N_43869,N_43658,N_43581);
nand U43870 (N_43870,N_43514,N_43507);
and U43871 (N_43871,N_43527,N_43601);
xnor U43872 (N_43872,N_43728,N_43604);
xor U43873 (N_43873,N_43694,N_43578);
or U43874 (N_43874,N_43504,N_43579);
and U43875 (N_43875,N_43566,N_43545);
or U43876 (N_43876,N_43573,N_43703);
xnor U43877 (N_43877,N_43588,N_43740);
nor U43878 (N_43878,N_43566,N_43647);
and U43879 (N_43879,N_43526,N_43522);
nor U43880 (N_43880,N_43681,N_43533);
or U43881 (N_43881,N_43561,N_43580);
nand U43882 (N_43882,N_43724,N_43741);
or U43883 (N_43883,N_43653,N_43660);
nand U43884 (N_43884,N_43518,N_43582);
nand U43885 (N_43885,N_43738,N_43658);
or U43886 (N_43886,N_43585,N_43564);
xor U43887 (N_43887,N_43708,N_43691);
and U43888 (N_43888,N_43656,N_43633);
nand U43889 (N_43889,N_43709,N_43712);
or U43890 (N_43890,N_43689,N_43710);
nand U43891 (N_43891,N_43621,N_43553);
nand U43892 (N_43892,N_43616,N_43527);
or U43893 (N_43893,N_43541,N_43732);
or U43894 (N_43894,N_43590,N_43529);
and U43895 (N_43895,N_43558,N_43568);
and U43896 (N_43896,N_43685,N_43519);
and U43897 (N_43897,N_43745,N_43670);
and U43898 (N_43898,N_43588,N_43598);
xnor U43899 (N_43899,N_43523,N_43652);
or U43900 (N_43900,N_43711,N_43672);
or U43901 (N_43901,N_43699,N_43676);
xnor U43902 (N_43902,N_43718,N_43573);
xnor U43903 (N_43903,N_43583,N_43549);
xnor U43904 (N_43904,N_43679,N_43642);
nand U43905 (N_43905,N_43714,N_43695);
or U43906 (N_43906,N_43656,N_43711);
or U43907 (N_43907,N_43741,N_43591);
xor U43908 (N_43908,N_43572,N_43573);
nor U43909 (N_43909,N_43628,N_43614);
or U43910 (N_43910,N_43582,N_43698);
xnor U43911 (N_43911,N_43505,N_43592);
nand U43912 (N_43912,N_43564,N_43612);
or U43913 (N_43913,N_43556,N_43701);
or U43914 (N_43914,N_43521,N_43502);
nor U43915 (N_43915,N_43683,N_43635);
xor U43916 (N_43916,N_43722,N_43674);
nor U43917 (N_43917,N_43593,N_43512);
nand U43918 (N_43918,N_43593,N_43716);
xnor U43919 (N_43919,N_43530,N_43531);
nand U43920 (N_43920,N_43547,N_43576);
nor U43921 (N_43921,N_43640,N_43549);
nand U43922 (N_43922,N_43685,N_43607);
and U43923 (N_43923,N_43581,N_43673);
and U43924 (N_43924,N_43672,N_43746);
or U43925 (N_43925,N_43620,N_43749);
and U43926 (N_43926,N_43585,N_43551);
or U43927 (N_43927,N_43600,N_43690);
and U43928 (N_43928,N_43700,N_43720);
nand U43929 (N_43929,N_43743,N_43580);
xor U43930 (N_43930,N_43557,N_43523);
nor U43931 (N_43931,N_43720,N_43632);
nand U43932 (N_43932,N_43554,N_43687);
xor U43933 (N_43933,N_43599,N_43601);
nand U43934 (N_43934,N_43591,N_43563);
nor U43935 (N_43935,N_43654,N_43526);
nor U43936 (N_43936,N_43581,N_43516);
nand U43937 (N_43937,N_43616,N_43514);
nor U43938 (N_43938,N_43537,N_43652);
nor U43939 (N_43939,N_43603,N_43618);
nor U43940 (N_43940,N_43697,N_43581);
nand U43941 (N_43941,N_43580,N_43706);
nand U43942 (N_43942,N_43615,N_43508);
xor U43943 (N_43943,N_43592,N_43518);
nor U43944 (N_43944,N_43646,N_43684);
nor U43945 (N_43945,N_43578,N_43707);
nand U43946 (N_43946,N_43613,N_43541);
nor U43947 (N_43947,N_43678,N_43534);
and U43948 (N_43948,N_43735,N_43702);
or U43949 (N_43949,N_43617,N_43572);
xnor U43950 (N_43950,N_43594,N_43614);
and U43951 (N_43951,N_43617,N_43727);
and U43952 (N_43952,N_43685,N_43603);
and U43953 (N_43953,N_43556,N_43521);
nor U43954 (N_43954,N_43723,N_43616);
nor U43955 (N_43955,N_43728,N_43747);
nand U43956 (N_43956,N_43711,N_43559);
or U43957 (N_43957,N_43654,N_43562);
and U43958 (N_43958,N_43651,N_43694);
or U43959 (N_43959,N_43583,N_43708);
nor U43960 (N_43960,N_43664,N_43656);
or U43961 (N_43961,N_43610,N_43740);
nand U43962 (N_43962,N_43554,N_43691);
nand U43963 (N_43963,N_43557,N_43535);
or U43964 (N_43964,N_43713,N_43654);
and U43965 (N_43965,N_43520,N_43731);
or U43966 (N_43966,N_43643,N_43634);
nand U43967 (N_43967,N_43589,N_43629);
nor U43968 (N_43968,N_43547,N_43732);
and U43969 (N_43969,N_43731,N_43556);
nand U43970 (N_43970,N_43621,N_43604);
nand U43971 (N_43971,N_43719,N_43543);
or U43972 (N_43972,N_43718,N_43598);
nor U43973 (N_43973,N_43568,N_43733);
or U43974 (N_43974,N_43668,N_43572);
nor U43975 (N_43975,N_43535,N_43524);
and U43976 (N_43976,N_43580,N_43719);
nand U43977 (N_43977,N_43715,N_43570);
nand U43978 (N_43978,N_43555,N_43654);
or U43979 (N_43979,N_43510,N_43668);
or U43980 (N_43980,N_43711,N_43678);
xnor U43981 (N_43981,N_43550,N_43723);
nand U43982 (N_43982,N_43535,N_43680);
xor U43983 (N_43983,N_43653,N_43519);
nor U43984 (N_43984,N_43743,N_43683);
nand U43985 (N_43985,N_43668,N_43589);
or U43986 (N_43986,N_43507,N_43631);
and U43987 (N_43987,N_43611,N_43597);
nand U43988 (N_43988,N_43663,N_43705);
xor U43989 (N_43989,N_43590,N_43516);
or U43990 (N_43990,N_43666,N_43712);
xnor U43991 (N_43991,N_43602,N_43616);
or U43992 (N_43992,N_43746,N_43708);
or U43993 (N_43993,N_43667,N_43701);
nor U43994 (N_43994,N_43663,N_43678);
nor U43995 (N_43995,N_43546,N_43606);
nand U43996 (N_43996,N_43507,N_43549);
nor U43997 (N_43997,N_43706,N_43725);
nand U43998 (N_43998,N_43696,N_43541);
nand U43999 (N_43999,N_43684,N_43602);
and U44000 (N_44000,N_43986,N_43899);
nor U44001 (N_44001,N_43954,N_43833);
nor U44002 (N_44002,N_43995,N_43911);
nand U44003 (N_44003,N_43783,N_43982);
and U44004 (N_44004,N_43901,N_43857);
nor U44005 (N_44005,N_43933,N_43798);
xnor U44006 (N_44006,N_43981,N_43809);
or U44007 (N_44007,N_43839,N_43902);
nor U44008 (N_44008,N_43816,N_43904);
xor U44009 (N_44009,N_43814,N_43941);
and U44010 (N_44010,N_43846,N_43907);
or U44011 (N_44011,N_43956,N_43806);
nand U44012 (N_44012,N_43860,N_43823);
and U44013 (N_44013,N_43934,N_43966);
and U44014 (N_44014,N_43920,N_43790);
xnor U44015 (N_44015,N_43879,N_43896);
and U44016 (N_44016,N_43759,N_43926);
nor U44017 (N_44017,N_43804,N_43851);
or U44018 (N_44018,N_43886,N_43938);
and U44019 (N_44019,N_43940,N_43842);
nand U44020 (N_44020,N_43887,N_43789);
and U44021 (N_44021,N_43773,N_43988);
or U44022 (N_44022,N_43867,N_43930);
xor U44023 (N_44023,N_43797,N_43916);
xnor U44024 (N_44024,N_43993,N_43983);
and U44025 (N_44025,N_43870,N_43776);
xor U44026 (N_44026,N_43868,N_43750);
and U44027 (N_44027,N_43862,N_43760);
and U44028 (N_44028,N_43889,N_43869);
or U44029 (N_44029,N_43977,N_43985);
nor U44030 (N_44030,N_43800,N_43754);
and U44031 (N_44031,N_43819,N_43894);
xor U44032 (N_44032,N_43968,N_43762);
xnor U44033 (N_44033,N_43781,N_43818);
or U44034 (N_44034,N_43787,N_43826);
xnor U44035 (N_44035,N_43890,N_43927);
xnor U44036 (N_44036,N_43923,N_43918);
or U44037 (N_44037,N_43791,N_43767);
and U44038 (N_44038,N_43793,N_43950);
and U44039 (N_44039,N_43794,N_43799);
nand U44040 (N_44040,N_43848,N_43900);
and U44041 (N_44041,N_43908,N_43830);
nand U44042 (N_44042,N_43953,N_43929);
xnor U44043 (N_44043,N_43965,N_43771);
nand U44044 (N_44044,N_43855,N_43847);
or U44045 (N_44045,N_43875,N_43775);
nand U44046 (N_44046,N_43925,N_43831);
nand U44047 (N_44047,N_43774,N_43921);
or U44048 (N_44048,N_43764,N_43976);
xor U44049 (N_44049,N_43897,N_43996);
nor U44050 (N_44050,N_43777,N_43992);
nor U44051 (N_44051,N_43970,N_43785);
nand U44052 (N_44052,N_43989,N_43786);
nor U44053 (N_44053,N_43905,N_43963);
xnor U44054 (N_44054,N_43919,N_43866);
nand U44055 (N_44055,N_43884,N_43872);
nand U44056 (N_44056,N_43946,N_43888);
nor U44057 (N_44057,N_43885,N_43917);
nor U44058 (N_44058,N_43844,N_43880);
nor U44059 (N_44059,N_43910,N_43780);
nor U44060 (N_44060,N_43947,N_43998);
nor U44061 (N_44061,N_43757,N_43945);
or U44062 (N_44062,N_43779,N_43778);
or U44063 (N_44063,N_43952,N_43997);
and U44064 (N_44064,N_43937,N_43763);
and U44065 (N_44065,N_43987,N_43815);
and U44066 (N_44066,N_43980,N_43784);
and U44067 (N_44067,N_43770,N_43840);
or U44068 (N_44068,N_43849,N_43974);
or U44069 (N_44069,N_43758,N_43854);
and U44070 (N_44070,N_43939,N_43756);
xor U44071 (N_44071,N_43853,N_43805);
or U44072 (N_44072,N_43994,N_43751);
nor U44073 (N_44073,N_43979,N_43765);
nand U44074 (N_44074,N_43936,N_43972);
nor U44075 (N_44075,N_43755,N_43942);
and U44076 (N_44076,N_43808,N_43864);
or U44077 (N_44077,N_43909,N_43825);
nand U44078 (N_44078,N_43883,N_43820);
nand U44079 (N_44079,N_43878,N_43795);
nand U44080 (N_44080,N_43827,N_43935);
xor U44081 (N_44081,N_43828,N_43821);
and U44082 (N_44082,N_43829,N_43877);
xnor U44083 (N_44083,N_43892,N_43811);
nor U44084 (N_44084,N_43859,N_43876);
xnor U44085 (N_44085,N_43766,N_43969);
nand U44086 (N_44086,N_43792,N_43990);
nand U44087 (N_44087,N_43971,N_43769);
or U44088 (N_44088,N_43943,N_43874);
xnor U44089 (N_44089,N_43817,N_43824);
nand U44090 (N_44090,N_43991,N_43881);
nand U44091 (N_44091,N_43856,N_43801);
or U44092 (N_44092,N_43863,N_43796);
nand U44093 (N_44093,N_43893,N_43958);
or U44094 (N_44094,N_43955,N_43895);
or U44095 (N_44095,N_43865,N_43836);
and U44096 (N_44096,N_43964,N_43999);
nor U44097 (N_44097,N_43837,N_43852);
nand U44098 (N_44098,N_43961,N_43835);
nand U44099 (N_44099,N_43975,N_43822);
xnor U44100 (N_44100,N_43838,N_43948);
and U44101 (N_44101,N_43861,N_43951);
nand U44102 (N_44102,N_43841,N_43761);
xnor U44103 (N_44103,N_43871,N_43915);
nand U44104 (N_44104,N_43850,N_43891);
or U44105 (N_44105,N_43807,N_43922);
or U44106 (N_44106,N_43752,N_43932);
nor U44107 (N_44107,N_43810,N_43782);
and U44108 (N_44108,N_43882,N_43772);
xor U44109 (N_44109,N_43967,N_43928);
nor U44110 (N_44110,N_43802,N_43858);
xnor U44111 (N_44111,N_43924,N_43978);
or U44112 (N_44112,N_43949,N_43768);
nor U44113 (N_44113,N_43813,N_43962);
nand U44114 (N_44114,N_43913,N_43812);
and U44115 (N_44115,N_43788,N_43959);
xnor U44116 (N_44116,N_43873,N_43931);
and U44117 (N_44117,N_43914,N_43906);
xor U44118 (N_44118,N_43832,N_43753);
or U44119 (N_44119,N_43845,N_43973);
nand U44120 (N_44120,N_43912,N_43957);
nand U44121 (N_44121,N_43984,N_43903);
nand U44122 (N_44122,N_43960,N_43834);
and U44123 (N_44123,N_43944,N_43803);
or U44124 (N_44124,N_43843,N_43898);
xor U44125 (N_44125,N_43941,N_43912);
nor U44126 (N_44126,N_43763,N_43966);
nor U44127 (N_44127,N_43928,N_43765);
and U44128 (N_44128,N_43938,N_43930);
nand U44129 (N_44129,N_43898,N_43760);
nor U44130 (N_44130,N_43762,N_43909);
nand U44131 (N_44131,N_43954,N_43925);
xnor U44132 (N_44132,N_43787,N_43868);
xnor U44133 (N_44133,N_43875,N_43961);
and U44134 (N_44134,N_43846,N_43916);
or U44135 (N_44135,N_43829,N_43768);
and U44136 (N_44136,N_43823,N_43958);
and U44137 (N_44137,N_43846,N_43926);
xor U44138 (N_44138,N_43977,N_43919);
nor U44139 (N_44139,N_43956,N_43756);
and U44140 (N_44140,N_43792,N_43910);
xnor U44141 (N_44141,N_43884,N_43780);
nor U44142 (N_44142,N_43797,N_43986);
nor U44143 (N_44143,N_43957,N_43826);
nor U44144 (N_44144,N_43893,N_43948);
nor U44145 (N_44145,N_43822,N_43929);
nor U44146 (N_44146,N_43927,N_43790);
nor U44147 (N_44147,N_43759,N_43872);
nand U44148 (N_44148,N_43774,N_43934);
or U44149 (N_44149,N_43916,N_43777);
nor U44150 (N_44150,N_43902,N_43875);
nand U44151 (N_44151,N_43960,N_43963);
nand U44152 (N_44152,N_43871,N_43801);
or U44153 (N_44153,N_43981,N_43888);
and U44154 (N_44154,N_43855,N_43768);
nand U44155 (N_44155,N_43901,N_43756);
xnor U44156 (N_44156,N_43999,N_43898);
nor U44157 (N_44157,N_43849,N_43903);
xnor U44158 (N_44158,N_43887,N_43832);
xor U44159 (N_44159,N_43978,N_43988);
nand U44160 (N_44160,N_43786,N_43902);
nor U44161 (N_44161,N_43941,N_43942);
xor U44162 (N_44162,N_43806,N_43762);
nand U44163 (N_44163,N_43803,N_43907);
or U44164 (N_44164,N_43817,N_43854);
and U44165 (N_44165,N_43950,N_43893);
and U44166 (N_44166,N_43939,N_43883);
nor U44167 (N_44167,N_43829,N_43972);
xnor U44168 (N_44168,N_43845,N_43939);
nor U44169 (N_44169,N_43808,N_43897);
nand U44170 (N_44170,N_43999,N_43809);
or U44171 (N_44171,N_43998,N_43752);
and U44172 (N_44172,N_43758,N_43971);
or U44173 (N_44173,N_43795,N_43982);
or U44174 (N_44174,N_43797,N_43935);
nand U44175 (N_44175,N_43856,N_43758);
xnor U44176 (N_44176,N_43948,N_43989);
nor U44177 (N_44177,N_43995,N_43752);
xor U44178 (N_44178,N_43907,N_43783);
xnor U44179 (N_44179,N_43808,N_43885);
nor U44180 (N_44180,N_43809,N_43787);
nand U44181 (N_44181,N_43838,N_43770);
xnor U44182 (N_44182,N_43962,N_43951);
xnor U44183 (N_44183,N_43925,N_43763);
nor U44184 (N_44184,N_43773,N_43876);
nor U44185 (N_44185,N_43977,N_43980);
nand U44186 (N_44186,N_43892,N_43824);
nand U44187 (N_44187,N_43861,N_43779);
xnor U44188 (N_44188,N_43943,N_43792);
or U44189 (N_44189,N_43779,N_43787);
xor U44190 (N_44190,N_43824,N_43791);
xnor U44191 (N_44191,N_43776,N_43752);
and U44192 (N_44192,N_43945,N_43837);
nand U44193 (N_44193,N_43854,N_43995);
or U44194 (N_44194,N_43838,N_43832);
or U44195 (N_44195,N_43856,N_43867);
nand U44196 (N_44196,N_43758,N_43889);
xor U44197 (N_44197,N_43803,N_43819);
xnor U44198 (N_44198,N_43814,N_43988);
or U44199 (N_44199,N_43968,N_43908);
xnor U44200 (N_44200,N_43967,N_43862);
nor U44201 (N_44201,N_43778,N_43959);
or U44202 (N_44202,N_43879,N_43856);
or U44203 (N_44203,N_43849,N_43941);
nand U44204 (N_44204,N_43942,N_43865);
or U44205 (N_44205,N_43879,N_43801);
xnor U44206 (N_44206,N_43932,N_43910);
nand U44207 (N_44207,N_43770,N_43877);
nor U44208 (N_44208,N_43789,N_43876);
xor U44209 (N_44209,N_43949,N_43924);
and U44210 (N_44210,N_43774,N_43776);
nor U44211 (N_44211,N_43795,N_43871);
xor U44212 (N_44212,N_43776,N_43901);
xor U44213 (N_44213,N_43775,N_43935);
nand U44214 (N_44214,N_43752,N_43898);
and U44215 (N_44215,N_43760,N_43879);
nand U44216 (N_44216,N_43787,N_43967);
nand U44217 (N_44217,N_43819,N_43824);
nand U44218 (N_44218,N_43888,N_43762);
or U44219 (N_44219,N_43841,N_43943);
or U44220 (N_44220,N_43904,N_43762);
xor U44221 (N_44221,N_43961,N_43833);
xor U44222 (N_44222,N_43919,N_43981);
and U44223 (N_44223,N_43951,N_43888);
nand U44224 (N_44224,N_43762,N_43775);
nor U44225 (N_44225,N_43942,N_43883);
nand U44226 (N_44226,N_43995,N_43814);
xor U44227 (N_44227,N_43950,N_43762);
xnor U44228 (N_44228,N_43919,N_43815);
xnor U44229 (N_44229,N_43871,N_43940);
nand U44230 (N_44230,N_43780,N_43957);
or U44231 (N_44231,N_43847,N_43882);
nor U44232 (N_44232,N_43918,N_43987);
xnor U44233 (N_44233,N_43840,N_43796);
and U44234 (N_44234,N_43989,N_43889);
and U44235 (N_44235,N_43956,N_43985);
xor U44236 (N_44236,N_43994,N_43756);
and U44237 (N_44237,N_43848,N_43956);
and U44238 (N_44238,N_43857,N_43890);
or U44239 (N_44239,N_43912,N_43795);
or U44240 (N_44240,N_43855,N_43951);
and U44241 (N_44241,N_43941,N_43760);
and U44242 (N_44242,N_43830,N_43914);
or U44243 (N_44243,N_43880,N_43930);
and U44244 (N_44244,N_43827,N_43960);
nand U44245 (N_44245,N_43809,N_43883);
or U44246 (N_44246,N_43963,N_43946);
or U44247 (N_44247,N_43881,N_43954);
nand U44248 (N_44248,N_43955,N_43892);
or U44249 (N_44249,N_43887,N_43767);
nand U44250 (N_44250,N_44142,N_44084);
xnor U44251 (N_44251,N_44070,N_44191);
or U44252 (N_44252,N_44232,N_44030);
xnor U44253 (N_44253,N_44151,N_44231);
or U44254 (N_44254,N_44208,N_44080);
or U44255 (N_44255,N_44107,N_44088);
or U44256 (N_44256,N_44121,N_44086);
xnor U44257 (N_44257,N_44021,N_44005);
nand U44258 (N_44258,N_44008,N_44205);
or U44259 (N_44259,N_44152,N_44123);
nor U44260 (N_44260,N_44178,N_44219);
nand U44261 (N_44261,N_44059,N_44003);
or U44262 (N_44262,N_44028,N_44158);
nor U44263 (N_44263,N_44105,N_44194);
nand U44264 (N_44264,N_44124,N_44237);
or U44265 (N_44265,N_44001,N_44122);
and U44266 (N_44266,N_44060,N_44136);
and U44267 (N_44267,N_44144,N_44246);
nor U44268 (N_44268,N_44182,N_44147);
and U44269 (N_44269,N_44118,N_44186);
nand U44270 (N_44270,N_44187,N_44026);
xor U44271 (N_44271,N_44154,N_44055);
nand U44272 (N_44272,N_44047,N_44244);
nand U44273 (N_44273,N_44183,N_44110);
nand U44274 (N_44274,N_44168,N_44020);
xor U44275 (N_44275,N_44193,N_44138);
or U44276 (N_44276,N_44033,N_44104);
and U44277 (N_44277,N_44130,N_44050);
or U44278 (N_44278,N_44019,N_44063);
nor U44279 (N_44279,N_44109,N_44103);
xor U44280 (N_44280,N_44073,N_44155);
nor U44281 (N_44281,N_44024,N_44115);
or U44282 (N_44282,N_44077,N_44101);
xor U44283 (N_44283,N_44017,N_44036);
and U44284 (N_44284,N_44198,N_44102);
xnor U44285 (N_44285,N_44164,N_44169);
and U44286 (N_44286,N_44185,N_44057);
and U44287 (N_44287,N_44096,N_44172);
or U44288 (N_44288,N_44058,N_44175);
nor U44289 (N_44289,N_44240,N_44127);
nor U44290 (N_44290,N_44247,N_44202);
or U44291 (N_44291,N_44010,N_44131);
nand U44292 (N_44292,N_44200,N_44249);
and U44293 (N_44293,N_44224,N_44197);
nor U44294 (N_44294,N_44176,N_44243);
xnor U44295 (N_44295,N_44120,N_44006);
xor U44296 (N_44296,N_44134,N_44211);
nor U44297 (N_44297,N_44072,N_44226);
nand U44298 (N_44298,N_44227,N_44233);
nor U44299 (N_44299,N_44217,N_44149);
or U44300 (N_44300,N_44239,N_44180);
or U44301 (N_44301,N_44038,N_44049);
nand U44302 (N_44302,N_44163,N_44009);
nand U44303 (N_44303,N_44091,N_44052);
xnor U44304 (N_44304,N_44094,N_44081);
xnor U44305 (N_44305,N_44014,N_44238);
xnor U44306 (N_44306,N_44076,N_44002);
nand U44307 (N_44307,N_44166,N_44071);
and U44308 (N_44308,N_44113,N_44220);
nand U44309 (N_44309,N_44184,N_44245);
or U44310 (N_44310,N_44218,N_44048);
nand U44311 (N_44311,N_44011,N_44074);
nor U44312 (N_44312,N_44141,N_44095);
and U44313 (N_44313,N_44087,N_44112);
or U44314 (N_44314,N_44248,N_44129);
and U44315 (N_44315,N_44043,N_44213);
or U44316 (N_44316,N_44106,N_44206);
xnor U44317 (N_44317,N_44126,N_44173);
or U44318 (N_44318,N_44207,N_44181);
xor U44319 (N_44319,N_44190,N_44140);
nand U44320 (N_44320,N_44223,N_44034);
or U44321 (N_44321,N_44125,N_44225);
nor U44322 (N_44322,N_44204,N_44159);
nor U44323 (N_44323,N_44097,N_44156);
and U44324 (N_44324,N_44075,N_44189);
xor U44325 (N_44325,N_44023,N_44090);
and U44326 (N_44326,N_44013,N_44143);
xor U44327 (N_44327,N_44114,N_44203);
or U44328 (N_44328,N_44079,N_44004);
xnor U44329 (N_44329,N_44171,N_44177);
xnor U44330 (N_44330,N_44051,N_44045);
and U44331 (N_44331,N_44221,N_44170);
and U44332 (N_44332,N_44067,N_44148);
nand U44333 (N_44333,N_44242,N_44089);
nand U44334 (N_44334,N_44162,N_44235);
nand U44335 (N_44335,N_44082,N_44117);
and U44336 (N_44336,N_44119,N_44041);
or U44337 (N_44337,N_44025,N_44215);
xor U44338 (N_44338,N_44061,N_44133);
or U44339 (N_44339,N_44108,N_44128);
nand U44340 (N_44340,N_44167,N_44032);
or U44341 (N_44341,N_44146,N_44029);
nor U44342 (N_44342,N_44111,N_44214);
or U44343 (N_44343,N_44031,N_44161);
or U44344 (N_44344,N_44092,N_44015);
nand U44345 (N_44345,N_44195,N_44150);
or U44346 (N_44346,N_44230,N_44099);
nor U44347 (N_44347,N_44139,N_44037);
and U44348 (N_44348,N_44210,N_44132);
and U44349 (N_44349,N_44046,N_44012);
and U44350 (N_44350,N_44216,N_44027);
and U44351 (N_44351,N_44201,N_44153);
nor U44352 (N_44352,N_44100,N_44064);
or U44353 (N_44353,N_44229,N_44157);
xor U44354 (N_44354,N_44234,N_44039);
xnor U44355 (N_44355,N_44068,N_44236);
xor U44356 (N_44356,N_44040,N_44228);
nor U44357 (N_44357,N_44212,N_44199);
and U44358 (N_44358,N_44022,N_44083);
nor U44359 (N_44359,N_44056,N_44000);
nor U44360 (N_44360,N_44078,N_44016);
nor U44361 (N_44361,N_44065,N_44179);
xor U44362 (N_44362,N_44137,N_44007);
nor U44363 (N_44363,N_44209,N_44145);
xor U44364 (N_44364,N_44160,N_44222);
and U44365 (N_44365,N_44135,N_44085);
and U44366 (N_44366,N_44174,N_44066);
nand U44367 (N_44367,N_44192,N_44053);
nand U44368 (N_44368,N_44188,N_44044);
or U44369 (N_44369,N_44116,N_44098);
nand U44370 (N_44370,N_44042,N_44018);
xnor U44371 (N_44371,N_44035,N_44241);
xnor U44372 (N_44372,N_44196,N_44093);
or U44373 (N_44373,N_44069,N_44062);
or U44374 (N_44374,N_44165,N_44054);
nor U44375 (N_44375,N_44211,N_44199);
and U44376 (N_44376,N_44060,N_44125);
nor U44377 (N_44377,N_44118,N_44023);
nand U44378 (N_44378,N_44221,N_44015);
xnor U44379 (N_44379,N_44041,N_44220);
and U44380 (N_44380,N_44084,N_44101);
nor U44381 (N_44381,N_44015,N_44189);
nand U44382 (N_44382,N_44015,N_44078);
xor U44383 (N_44383,N_44125,N_44188);
xnor U44384 (N_44384,N_44239,N_44096);
nor U44385 (N_44385,N_44048,N_44008);
and U44386 (N_44386,N_44023,N_44000);
nand U44387 (N_44387,N_44189,N_44193);
nor U44388 (N_44388,N_44231,N_44076);
xnor U44389 (N_44389,N_44096,N_44148);
and U44390 (N_44390,N_44043,N_44024);
or U44391 (N_44391,N_44239,N_44038);
nor U44392 (N_44392,N_44032,N_44165);
nor U44393 (N_44393,N_44188,N_44089);
nor U44394 (N_44394,N_44219,N_44160);
and U44395 (N_44395,N_44220,N_44098);
and U44396 (N_44396,N_44072,N_44095);
nand U44397 (N_44397,N_44133,N_44039);
and U44398 (N_44398,N_44035,N_44087);
and U44399 (N_44399,N_44232,N_44202);
xnor U44400 (N_44400,N_44247,N_44197);
nor U44401 (N_44401,N_44058,N_44163);
nand U44402 (N_44402,N_44229,N_44049);
or U44403 (N_44403,N_44143,N_44117);
or U44404 (N_44404,N_44197,N_44077);
and U44405 (N_44405,N_44104,N_44078);
and U44406 (N_44406,N_44182,N_44010);
nor U44407 (N_44407,N_44212,N_44184);
nor U44408 (N_44408,N_44002,N_44009);
and U44409 (N_44409,N_44246,N_44011);
and U44410 (N_44410,N_44055,N_44151);
nor U44411 (N_44411,N_44238,N_44166);
and U44412 (N_44412,N_44146,N_44229);
nand U44413 (N_44413,N_44238,N_44215);
nor U44414 (N_44414,N_44241,N_44082);
nor U44415 (N_44415,N_44106,N_44246);
xor U44416 (N_44416,N_44129,N_44131);
nand U44417 (N_44417,N_44004,N_44092);
and U44418 (N_44418,N_44085,N_44060);
or U44419 (N_44419,N_44096,N_44228);
nand U44420 (N_44420,N_44176,N_44223);
nor U44421 (N_44421,N_44236,N_44186);
xnor U44422 (N_44422,N_44054,N_44012);
nand U44423 (N_44423,N_44056,N_44240);
xor U44424 (N_44424,N_44117,N_44023);
nor U44425 (N_44425,N_44159,N_44009);
nor U44426 (N_44426,N_44149,N_44102);
xnor U44427 (N_44427,N_44179,N_44170);
nor U44428 (N_44428,N_44031,N_44187);
and U44429 (N_44429,N_44123,N_44058);
or U44430 (N_44430,N_44158,N_44096);
or U44431 (N_44431,N_44026,N_44190);
xnor U44432 (N_44432,N_44010,N_44190);
nand U44433 (N_44433,N_44071,N_44199);
and U44434 (N_44434,N_44220,N_44153);
nor U44435 (N_44435,N_44222,N_44005);
xnor U44436 (N_44436,N_44223,N_44236);
or U44437 (N_44437,N_44110,N_44055);
nor U44438 (N_44438,N_44112,N_44098);
nor U44439 (N_44439,N_44193,N_44074);
nand U44440 (N_44440,N_44228,N_44214);
and U44441 (N_44441,N_44226,N_44061);
nand U44442 (N_44442,N_44221,N_44091);
nor U44443 (N_44443,N_44122,N_44089);
nand U44444 (N_44444,N_44138,N_44249);
nand U44445 (N_44445,N_44175,N_44130);
and U44446 (N_44446,N_44216,N_44145);
and U44447 (N_44447,N_44225,N_44216);
xor U44448 (N_44448,N_44105,N_44191);
and U44449 (N_44449,N_44186,N_44222);
and U44450 (N_44450,N_44099,N_44024);
nor U44451 (N_44451,N_44213,N_44090);
nor U44452 (N_44452,N_44231,N_44171);
and U44453 (N_44453,N_44008,N_44184);
xor U44454 (N_44454,N_44207,N_44059);
nand U44455 (N_44455,N_44077,N_44212);
nand U44456 (N_44456,N_44156,N_44144);
or U44457 (N_44457,N_44134,N_44118);
xor U44458 (N_44458,N_44223,N_44171);
or U44459 (N_44459,N_44053,N_44155);
nor U44460 (N_44460,N_44142,N_44188);
and U44461 (N_44461,N_44223,N_44002);
and U44462 (N_44462,N_44092,N_44002);
nor U44463 (N_44463,N_44147,N_44102);
or U44464 (N_44464,N_44148,N_44179);
or U44465 (N_44465,N_44232,N_44145);
and U44466 (N_44466,N_44049,N_44202);
or U44467 (N_44467,N_44168,N_44225);
xnor U44468 (N_44468,N_44158,N_44092);
nor U44469 (N_44469,N_44073,N_44154);
xnor U44470 (N_44470,N_44007,N_44188);
or U44471 (N_44471,N_44155,N_44088);
nand U44472 (N_44472,N_44068,N_44140);
and U44473 (N_44473,N_44075,N_44051);
or U44474 (N_44474,N_44113,N_44229);
or U44475 (N_44475,N_44211,N_44084);
nor U44476 (N_44476,N_44091,N_44199);
nor U44477 (N_44477,N_44103,N_44016);
xnor U44478 (N_44478,N_44124,N_44216);
nand U44479 (N_44479,N_44231,N_44083);
nor U44480 (N_44480,N_44101,N_44124);
nor U44481 (N_44481,N_44019,N_44203);
xnor U44482 (N_44482,N_44097,N_44178);
and U44483 (N_44483,N_44141,N_44112);
and U44484 (N_44484,N_44126,N_44072);
nand U44485 (N_44485,N_44075,N_44045);
nor U44486 (N_44486,N_44249,N_44079);
or U44487 (N_44487,N_44026,N_44225);
xnor U44488 (N_44488,N_44003,N_44241);
nor U44489 (N_44489,N_44026,N_44070);
and U44490 (N_44490,N_44017,N_44206);
nor U44491 (N_44491,N_44249,N_44033);
or U44492 (N_44492,N_44045,N_44179);
xnor U44493 (N_44493,N_44230,N_44087);
nor U44494 (N_44494,N_44048,N_44239);
or U44495 (N_44495,N_44022,N_44074);
and U44496 (N_44496,N_44080,N_44047);
nor U44497 (N_44497,N_44007,N_44108);
and U44498 (N_44498,N_44226,N_44179);
or U44499 (N_44499,N_44163,N_44215);
nand U44500 (N_44500,N_44484,N_44425);
nand U44501 (N_44501,N_44462,N_44379);
nor U44502 (N_44502,N_44281,N_44333);
or U44503 (N_44503,N_44414,N_44334);
nand U44504 (N_44504,N_44331,N_44358);
nor U44505 (N_44505,N_44311,N_44361);
nor U44506 (N_44506,N_44261,N_44276);
and U44507 (N_44507,N_44493,N_44445);
nor U44508 (N_44508,N_44316,N_44250);
or U44509 (N_44509,N_44303,N_44465);
xor U44510 (N_44510,N_44475,N_44440);
and U44511 (N_44511,N_44420,N_44289);
or U44512 (N_44512,N_44285,N_44340);
nor U44513 (N_44513,N_44328,N_44399);
nand U44514 (N_44514,N_44388,N_44436);
nor U44515 (N_44515,N_44470,N_44277);
nor U44516 (N_44516,N_44404,N_44429);
nand U44517 (N_44517,N_44374,N_44390);
and U44518 (N_44518,N_44343,N_44325);
nand U44519 (N_44519,N_44430,N_44498);
nand U44520 (N_44520,N_44452,N_44409);
nand U44521 (N_44521,N_44258,N_44392);
xor U44522 (N_44522,N_44299,N_44473);
or U44523 (N_44523,N_44380,N_44356);
nor U44524 (N_44524,N_44265,N_44349);
or U44525 (N_44525,N_44268,N_44278);
and U44526 (N_44526,N_44447,N_44370);
xnor U44527 (N_44527,N_44407,N_44290);
xnor U44528 (N_44528,N_44469,N_44309);
nand U44529 (N_44529,N_44284,N_44454);
xnor U44530 (N_44530,N_44317,N_44294);
and U44531 (N_44531,N_44481,N_44310);
nand U44532 (N_44532,N_44305,N_44342);
or U44533 (N_44533,N_44350,N_44275);
or U44534 (N_44534,N_44413,N_44408);
or U44535 (N_44535,N_44482,N_44422);
or U44536 (N_44536,N_44449,N_44394);
or U44537 (N_44537,N_44458,N_44424);
or U44538 (N_44538,N_44416,N_44496);
or U44539 (N_44539,N_44463,N_44260);
or U44540 (N_44540,N_44400,N_44385);
and U44541 (N_44541,N_44396,N_44485);
or U44542 (N_44542,N_44368,N_44423);
and U44543 (N_44543,N_44417,N_44282);
and U44544 (N_44544,N_44467,N_44348);
xor U44545 (N_44545,N_44369,N_44320);
xnor U44546 (N_44546,N_44491,N_44347);
nand U44547 (N_44547,N_44293,N_44412);
xor U44548 (N_44548,N_44315,N_44327);
or U44549 (N_44549,N_44302,N_44494);
xor U44550 (N_44550,N_44376,N_44357);
and U44551 (N_44551,N_44387,N_44252);
xnor U44552 (N_44552,N_44450,N_44433);
or U44553 (N_44553,N_44345,N_44397);
nand U44554 (N_44554,N_44280,N_44464);
nand U44555 (N_44555,N_44487,N_44259);
nor U44556 (N_44556,N_44418,N_44324);
nor U44557 (N_44557,N_44495,N_44439);
nor U44558 (N_44558,N_44337,N_44480);
xor U44559 (N_44559,N_44314,N_44364);
or U44560 (N_44560,N_44295,N_44474);
xnor U44561 (N_44561,N_44405,N_44352);
nand U44562 (N_44562,N_44319,N_44288);
or U44563 (N_44563,N_44403,N_44483);
nor U44564 (N_44564,N_44323,N_44497);
and U44565 (N_44565,N_44300,N_44393);
and U44566 (N_44566,N_44428,N_44306);
nand U44567 (N_44567,N_44269,N_44382);
nor U44568 (N_44568,N_44460,N_44264);
nand U44569 (N_44569,N_44466,N_44459);
and U44570 (N_44570,N_44410,N_44346);
and U44571 (N_44571,N_44344,N_44451);
nand U44572 (N_44572,N_44271,N_44291);
and U44573 (N_44573,N_44292,N_44395);
and U44574 (N_44574,N_44415,N_44312);
xnor U44575 (N_44575,N_44490,N_44386);
nand U44576 (N_44576,N_44377,N_44365);
xor U44577 (N_44577,N_44402,N_44383);
xor U44578 (N_44578,N_44455,N_44338);
or U44579 (N_44579,N_44472,N_44448);
or U44580 (N_44580,N_44354,N_44360);
nor U44581 (N_44581,N_44499,N_44341);
or U44582 (N_44582,N_44479,N_44362);
and U44583 (N_44583,N_44272,N_44468);
or U44584 (N_44584,N_44427,N_44267);
or U44585 (N_44585,N_44263,N_44286);
nand U44586 (N_44586,N_44330,N_44398);
xor U44587 (N_44587,N_44438,N_44322);
or U44588 (N_44588,N_44266,N_44296);
nor U44589 (N_44589,N_44257,N_44318);
nor U44590 (N_44590,N_44287,N_44371);
and U44591 (N_44591,N_44453,N_44339);
or U44592 (N_44592,N_44461,N_44378);
xor U44593 (N_44593,N_44471,N_44298);
nor U44594 (N_44594,N_44435,N_44419);
nor U44595 (N_44595,N_44434,N_44373);
and U44596 (N_44596,N_44442,N_44366);
and U44597 (N_44597,N_44389,N_44477);
or U44598 (N_44598,N_44273,N_44254);
and U44599 (N_44599,N_44251,N_44351);
nand U44600 (N_44600,N_44426,N_44372);
xnor U44601 (N_44601,N_44279,N_44253);
and U44602 (N_44602,N_44329,N_44488);
and U44603 (N_44603,N_44421,N_44441);
or U44604 (N_44604,N_44355,N_44384);
and U44605 (N_44605,N_44432,N_44336);
nand U44606 (N_44606,N_44478,N_44406);
xor U44607 (N_44607,N_44270,N_44456);
nand U44608 (N_44608,N_44411,N_44437);
nand U44609 (N_44609,N_44367,N_44486);
and U44610 (N_44610,N_44332,N_44476);
or U44611 (N_44611,N_44353,N_44381);
nor U44612 (N_44612,N_44492,N_44363);
xor U44613 (N_44613,N_44457,N_44335);
and U44614 (N_44614,N_44255,N_44359);
or U44615 (N_44615,N_44308,N_44375);
or U44616 (N_44616,N_44256,N_44443);
or U44617 (N_44617,N_44307,N_44304);
nor U44618 (N_44618,N_44489,N_44301);
and U44619 (N_44619,N_44326,N_44391);
and U44620 (N_44620,N_44446,N_44401);
xnor U44621 (N_44621,N_44444,N_44262);
nor U44622 (N_44622,N_44321,N_44313);
xnor U44623 (N_44623,N_44274,N_44297);
nor U44624 (N_44624,N_44283,N_44431);
and U44625 (N_44625,N_44305,N_44400);
nand U44626 (N_44626,N_44444,N_44494);
and U44627 (N_44627,N_44314,N_44429);
or U44628 (N_44628,N_44492,N_44387);
nand U44629 (N_44629,N_44363,N_44301);
nand U44630 (N_44630,N_44442,N_44497);
nor U44631 (N_44631,N_44371,N_44286);
and U44632 (N_44632,N_44464,N_44268);
xnor U44633 (N_44633,N_44481,N_44346);
xnor U44634 (N_44634,N_44286,N_44309);
nor U44635 (N_44635,N_44441,N_44261);
or U44636 (N_44636,N_44307,N_44440);
nor U44637 (N_44637,N_44395,N_44420);
or U44638 (N_44638,N_44393,N_44391);
and U44639 (N_44639,N_44486,N_44499);
xnor U44640 (N_44640,N_44471,N_44428);
nand U44641 (N_44641,N_44323,N_44493);
or U44642 (N_44642,N_44462,N_44331);
nand U44643 (N_44643,N_44259,N_44403);
and U44644 (N_44644,N_44377,N_44277);
nor U44645 (N_44645,N_44425,N_44281);
or U44646 (N_44646,N_44399,N_44290);
and U44647 (N_44647,N_44322,N_44295);
nor U44648 (N_44648,N_44403,N_44322);
nand U44649 (N_44649,N_44364,N_44297);
nand U44650 (N_44650,N_44369,N_44387);
xnor U44651 (N_44651,N_44417,N_44291);
nor U44652 (N_44652,N_44268,N_44397);
and U44653 (N_44653,N_44288,N_44434);
nor U44654 (N_44654,N_44361,N_44472);
xor U44655 (N_44655,N_44417,N_44455);
nand U44656 (N_44656,N_44358,N_44333);
nor U44657 (N_44657,N_44386,N_44306);
nand U44658 (N_44658,N_44290,N_44355);
and U44659 (N_44659,N_44468,N_44287);
xor U44660 (N_44660,N_44394,N_44396);
or U44661 (N_44661,N_44377,N_44372);
nor U44662 (N_44662,N_44420,N_44399);
nand U44663 (N_44663,N_44435,N_44325);
nor U44664 (N_44664,N_44335,N_44371);
nor U44665 (N_44665,N_44265,N_44491);
and U44666 (N_44666,N_44259,N_44453);
nand U44667 (N_44667,N_44460,N_44408);
nand U44668 (N_44668,N_44266,N_44270);
nor U44669 (N_44669,N_44252,N_44371);
nor U44670 (N_44670,N_44312,N_44276);
nor U44671 (N_44671,N_44304,N_44335);
nor U44672 (N_44672,N_44334,N_44261);
nor U44673 (N_44673,N_44379,N_44388);
xor U44674 (N_44674,N_44419,N_44409);
or U44675 (N_44675,N_44277,N_44473);
nand U44676 (N_44676,N_44299,N_44262);
nor U44677 (N_44677,N_44420,N_44400);
or U44678 (N_44678,N_44455,N_44451);
xnor U44679 (N_44679,N_44455,N_44390);
or U44680 (N_44680,N_44399,N_44427);
or U44681 (N_44681,N_44283,N_44322);
nor U44682 (N_44682,N_44255,N_44365);
and U44683 (N_44683,N_44351,N_44355);
and U44684 (N_44684,N_44465,N_44496);
nor U44685 (N_44685,N_44426,N_44289);
nor U44686 (N_44686,N_44382,N_44280);
or U44687 (N_44687,N_44281,N_44254);
nand U44688 (N_44688,N_44253,N_44339);
and U44689 (N_44689,N_44404,N_44342);
nand U44690 (N_44690,N_44336,N_44446);
nand U44691 (N_44691,N_44459,N_44395);
and U44692 (N_44692,N_44275,N_44448);
xor U44693 (N_44693,N_44499,N_44254);
xnor U44694 (N_44694,N_44397,N_44371);
xor U44695 (N_44695,N_44291,N_44355);
nor U44696 (N_44696,N_44464,N_44322);
nor U44697 (N_44697,N_44392,N_44278);
or U44698 (N_44698,N_44251,N_44382);
xor U44699 (N_44699,N_44262,N_44456);
xnor U44700 (N_44700,N_44427,N_44375);
and U44701 (N_44701,N_44414,N_44457);
nor U44702 (N_44702,N_44398,N_44347);
nor U44703 (N_44703,N_44352,N_44354);
nor U44704 (N_44704,N_44339,N_44319);
and U44705 (N_44705,N_44419,N_44319);
nor U44706 (N_44706,N_44373,N_44499);
nand U44707 (N_44707,N_44299,N_44455);
or U44708 (N_44708,N_44437,N_44308);
or U44709 (N_44709,N_44270,N_44497);
nand U44710 (N_44710,N_44284,N_44311);
nand U44711 (N_44711,N_44253,N_44294);
or U44712 (N_44712,N_44291,N_44437);
and U44713 (N_44713,N_44441,N_44340);
xnor U44714 (N_44714,N_44428,N_44312);
or U44715 (N_44715,N_44257,N_44288);
xnor U44716 (N_44716,N_44271,N_44484);
or U44717 (N_44717,N_44289,N_44257);
nand U44718 (N_44718,N_44284,N_44361);
or U44719 (N_44719,N_44405,N_44467);
or U44720 (N_44720,N_44496,N_44302);
nand U44721 (N_44721,N_44427,N_44264);
nand U44722 (N_44722,N_44469,N_44496);
xnor U44723 (N_44723,N_44469,N_44335);
or U44724 (N_44724,N_44320,N_44366);
nand U44725 (N_44725,N_44317,N_44256);
and U44726 (N_44726,N_44402,N_44393);
or U44727 (N_44727,N_44386,N_44414);
and U44728 (N_44728,N_44408,N_44326);
nand U44729 (N_44729,N_44338,N_44488);
or U44730 (N_44730,N_44392,N_44340);
nand U44731 (N_44731,N_44291,N_44380);
nand U44732 (N_44732,N_44411,N_44276);
xor U44733 (N_44733,N_44282,N_44339);
and U44734 (N_44734,N_44456,N_44470);
xor U44735 (N_44735,N_44409,N_44287);
nand U44736 (N_44736,N_44265,N_44395);
or U44737 (N_44737,N_44480,N_44404);
nand U44738 (N_44738,N_44321,N_44364);
or U44739 (N_44739,N_44396,N_44295);
nand U44740 (N_44740,N_44266,N_44418);
and U44741 (N_44741,N_44470,N_44311);
or U44742 (N_44742,N_44469,N_44467);
xor U44743 (N_44743,N_44281,N_44494);
and U44744 (N_44744,N_44369,N_44433);
nor U44745 (N_44745,N_44309,N_44421);
xnor U44746 (N_44746,N_44285,N_44450);
or U44747 (N_44747,N_44434,N_44337);
nor U44748 (N_44748,N_44421,N_44468);
or U44749 (N_44749,N_44384,N_44306);
and U44750 (N_44750,N_44701,N_44646);
nand U44751 (N_44751,N_44685,N_44592);
xnor U44752 (N_44752,N_44571,N_44519);
or U44753 (N_44753,N_44738,N_44748);
and U44754 (N_44754,N_44542,N_44591);
and U44755 (N_44755,N_44640,N_44724);
or U44756 (N_44756,N_44555,N_44512);
nor U44757 (N_44757,N_44507,N_44660);
and U44758 (N_44758,N_44593,N_44671);
nand U44759 (N_44759,N_44536,N_44699);
and U44760 (N_44760,N_44517,N_44672);
xnor U44761 (N_44761,N_44734,N_44632);
or U44762 (N_44762,N_44626,N_44749);
nor U44763 (N_44763,N_44580,N_44655);
and U44764 (N_44764,N_44730,N_44703);
and U44765 (N_44765,N_44621,N_44563);
nor U44766 (N_44766,N_44638,N_44719);
nand U44767 (N_44767,N_44584,N_44746);
nor U44768 (N_44768,N_44642,N_44612);
xor U44769 (N_44769,N_44511,N_44652);
xnor U44770 (N_44770,N_44616,N_44560);
nand U44771 (N_44771,N_44645,N_44704);
nand U44772 (N_44772,N_44595,N_44610);
xor U44773 (N_44773,N_44714,N_44518);
nand U44774 (N_44774,N_44688,N_44682);
nand U44775 (N_44775,N_44596,N_44581);
xnor U44776 (N_44776,N_44594,N_44538);
nand U44777 (N_44777,N_44663,N_44631);
or U44778 (N_44778,N_44679,N_44712);
and U44779 (N_44779,N_44609,N_44624);
or U44780 (N_44780,N_44721,N_44656);
xor U44781 (N_44781,N_44524,N_44617);
nand U44782 (N_44782,N_44668,N_44564);
or U44783 (N_44783,N_44619,N_44601);
nand U44784 (N_44784,N_44557,N_44526);
or U44785 (N_44785,N_44549,N_44692);
xor U44786 (N_44786,N_44653,N_44691);
xnor U44787 (N_44787,N_44503,N_44556);
xnor U44788 (N_44788,N_44669,N_44508);
or U44789 (N_44789,N_44603,N_44681);
and U44790 (N_44790,N_44504,N_44711);
or U44791 (N_44791,N_44558,N_44583);
xnor U44792 (N_44792,N_44540,N_44622);
xnor U44793 (N_44793,N_44598,N_44728);
nand U44794 (N_44794,N_44729,N_44713);
and U44795 (N_44795,N_44725,N_44678);
or U44796 (N_44796,N_44618,N_44522);
nor U44797 (N_44797,N_44569,N_44567);
nand U44798 (N_44798,N_44548,N_44505);
xnor U44799 (N_44799,N_44731,N_44525);
and U44800 (N_44800,N_44551,N_44579);
xnor U44801 (N_44801,N_44572,N_44531);
xor U44802 (N_44802,N_44723,N_44606);
or U44803 (N_44803,N_44546,N_44726);
nor U44804 (N_44804,N_44576,N_44514);
and U44805 (N_44805,N_44667,N_44697);
nand U44806 (N_44806,N_44544,N_44620);
and U44807 (N_44807,N_44597,N_44587);
nor U44808 (N_44808,N_44732,N_44720);
nand U44809 (N_44809,N_44537,N_44707);
or U44810 (N_44810,N_44659,N_44665);
nand U44811 (N_44811,N_44541,N_44589);
nor U44812 (N_44812,N_44575,N_44550);
nor U44813 (N_44813,N_44737,N_44637);
nand U44814 (N_44814,N_44509,N_44705);
xnor U44815 (N_44815,N_44578,N_44528);
xnor U44816 (N_44816,N_44510,N_44561);
xor U44817 (N_44817,N_44670,N_44742);
xnor U44818 (N_44818,N_44658,N_44698);
nor U44819 (N_44819,N_44585,N_44650);
xnor U44820 (N_44820,N_44516,N_44676);
xnor U44821 (N_44821,N_44706,N_44747);
nand U44822 (N_44822,N_44529,N_44717);
nor U44823 (N_44823,N_44552,N_44568);
nand U44824 (N_44824,N_44613,N_44559);
or U44825 (N_44825,N_44684,N_44661);
or U44826 (N_44826,N_44666,N_44677);
nor U44827 (N_44827,N_44735,N_44530);
nand U44828 (N_44828,N_44633,N_44741);
nand U44829 (N_44829,N_44693,N_44696);
nand U44830 (N_44830,N_44644,N_44574);
or U44831 (N_44831,N_44573,N_44590);
nand U44832 (N_44832,N_44521,N_44527);
or U44833 (N_44833,N_44715,N_44623);
xnor U44834 (N_44834,N_44545,N_44700);
or U44835 (N_44835,N_44532,N_44722);
xor U44836 (N_44836,N_44702,N_44648);
xnor U44837 (N_44837,N_44727,N_44586);
and U44838 (N_44838,N_44582,N_44506);
xor U44839 (N_44839,N_44602,N_44639);
nor U44840 (N_44840,N_44554,N_44533);
or U44841 (N_44841,N_44520,N_44740);
or U44842 (N_44842,N_44739,N_44570);
nor U44843 (N_44843,N_44662,N_44736);
xor U44844 (N_44844,N_44625,N_44636);
and U44845 (N_44845,N_44635,N_44654);
and U44846 (N_44846,N_44577,N_44680);
and U44847 (N_44847,N_44502,N_44718);
or U44848 (N_44848,N_44744,N_44694);
nand U44849 (N_44849,N_44641,N_44553);
nor U44850 (N_44850,N_44643,N_44716);
nor U44851 (N_44851,N_44709,N_44614);
and U44852 (N_44852,N_44600,N_44611);
xor U44853 (N_44853,N_44630,N_44615);
nand U44854 (N_44854,N_44733,N_44687);
and U44855 (N_44855,N_44689,N_44566);
nor U44856 (N_44856,N_44690,N_44607);
xor U44857 (N_44857,N_44515,N_44673);
or U44858 (N_44858,N_44664,N_44599);
and U44859 (N_44859,N_44695,N_44604);
and U44860 (N_44860,N_44686,N_44629);
nor U44861 (N_44861,N_44743,N_44535);
xnor U44862 (N_44862,N_44608,N_44647);
nor U44863 (N_44863,N_44539,N_44628);
xor U44864 (N_44864,N_44565,N_44634);
or U44865 (N_44865,N_44675,N_44500);
or U44866 (N_44866,N_44543,N_44710);
or U44867 (N_44867,N_44523,N_44605);
and U44868 (N_44868,N_44745,N_44513);
xor U44869 (N_44869,N_44501,N_44649);
and U44870 (N_44870,N_44534,N_44708);
nor U44871 (N_44871,N_44683,N_44588);
or U44872 (N_44872,N_44651,N_44562);
xnor U44873 (N_44873,N_44657,N_44627);
nand U44874 (N_44874,N_44674,N_44547);
or U44875 (N_44875,N_44584,N_44535);
or U44876 (N_44876,N_44702,N_44578);
nor U44877 (N_44877,N_44666,N_44502);
or U44878 (N_44878,N_44722,N_44749);
nand U44879 (N_44879,N_44597,N_44500);
nand U44880 (N_44880,N_44503,N_44693);
nand U44881 (N_44881,N_44574,N_44517);
nor U44882 (N_44882,N_44643,N_44717);
nand U44883 (N_44883,N_44535,N_44603);
and U44884 (N_44884,N_44565,N_44584);
nor U44885 (N_44885,N_44525,N_44611);
nand U44886 (N_44886,N_44670,N_44710);
xor U44887 (N_44887,N_44725,N_44523);
and U44888 (N_44888,N_44656,N_44613);
or U44889 (N_44889,N_44510,N_44612);
or U44890 (N_44890,N_44686,N_44746);
or U44891 (N_44891,N_44501,N_44628);
and U44892 (N_44892,N_44726,N_44652);
and U44893 (N_44893,N_44726,N_44533);
nand U44894 (N_44894,N_44735,N_44557);
nor U44895 (N_44895,N_44631,N_44636);
nor U44896 (N_44896,N_44723,N_44681);
nand U44897 (N_44897,N_44599,N_44504);
and U44898 (N_44898,N_44549,N_44710);
or U44899 (N_44899,N_44534,N_44581);
nor U44900 (N_44900,N_44629,N_44660);
nor U44901 (N_44901,N_44642,N_44600);
and U44902 (N_44902,N_44643,N_44592);
nor U44903 (N_44903,N_44541,N_44548);
nor U44904 (N_44904,N_44739,N_44585);
nor U44905 (N_44905,N_44585,N_44699);
nand U44906 (N_44906,N_44523,N_44531);
xnor U44907 (N_44907,N_44547,N_44585);
nor U44908 (N_44908,N_44548,N_44746);
and U44909 (N_44909,N_44552,N_44581);
and U44910 (N_44910,N_44514,N_44566);
xnor U44911 (N_44911,N_44643,N_44603);
nor U44912 (N_44912,N_44622,N_44523);
nor U44913 (N_44913,N_44739,N_44696);
nor U44914 (N_44914,N_44723,N_44658);
nand U44915 (N_44915,N_44681,N_44544);
xor U44916 (N_44916,N_44709,N_44617);
nor U44917 (N_44917,N_44713,N_44570);
or U44918 (N_44918,N_44683,N_44600);
or U44919 (N_44919,N_44681,N_44618);
xnor U44920 (N_44920,N_44610,N_44716);
and U44921 (N_44921,N_44607,N_44527);
nand U44922 (N_44922,N_44672,N_44509);
xor U44923 (N_44923,N_44526,N_44548);
nor U44924 (N_44924,N_44689,N_44651);
and U44925 (N_44925,N_44569,N_44745);
nor U44926 (N_44926,N_44718,N_44692);
nor U44927 (N_44927,N_44697,N_44689);
nand U44928 (N_44928,N_44531,N_44654);
nor U44929 (N_44929,N_44531,N_44559);
nand U44930 (N_44930,N_44568,N_44569);
nor U44931 (N_44931,N_44610,N_44526);
and U44932 (N_44932,N_44553,N_44585);
nor U44933 (N_44933,N_44627,N_44656);
or U44934 (N_44934,N_44612,N_44657);
nor U44935 (N_44935,N_44623,N_44661);
xor U44936 (N_44936,N_44633,N_44746);
xnor U44937 (N_44937,N_44608,N_44514);
nand U44938 (N_44938,N_44687,N_44661);
nand U44939 (N_44939,N_44578,N_44632);
or U44940 (N_44940,N_44731,N_44624);
xor U44941 (N_44941,N_44601,N_44640);
nand U44942 (N_44942,N_44512,N_44677);
xor U44943 (N_44943,N_44671,N_44525);
nor U44944 (N_44944,N_44662,N_44583);
xnor U44945 (N_44945,N_44586,N_44741);
xnor U44946 (N_44946,N_44654,N_44515);
or U44947 (N_44947,N_44524,N_44512);
or U44948 (N_44948,N_44502,N_44589);
nor U44949 (N_44949,N_44530,N_44544);
and U44950 (N_44950,N_44741,N_44611);
or U44951 (N_44951,N_44607,N_44686);
nand U44952 (N_44952,N_44641,N_44707);
nor U44953 (N_44953,N_44545,N_44693);
xnor U44954 (N_44954,N_44709,N_44653);
and U44955 (N_44955,N_44527,N_44508);
nand U44956 (N_44956,N_44629,N_44626);
or U44957 (N_44957,N_44703,N_44512);
nor U44958 (N_44958,N_44557,N_44577);
xnor U44959 (N_44959,N_44650,N_44734);
xor U44960 (N_44960,N_44661,N_44504);
and U44961 (N_44961,N_44608,N_44713);
xor U44962 (N_44962,N_44590,N_44686);
and U44963 (N_44963,N_44704,N_44711);
xnor U44964 (N_44964,N_44647,N_44626);
or U44965 (N_44965,N_44570,N_44562);
or U44966 (N_44966,N_44702,N_44714);
or U44967 (N_44967,N_44552,N_44637);
nor U44968 (N_44968,N_44707,N_44704);
or U44969 (N_44969,N_44582,N_44727);
nor U44970 (N_44970,N_44746,N_44551);
nand U44971 (N_44971,N_44609,N_44602);
nand U44972 (N_44972,N_44624,N_44735);
or U44973 (N_44973,N_44719,N_44735);
nand U44974 (N_44974,N_44620,N_44703);
nor U44975 (N_44975,N_44616,N_44711);
nand U44976 (N_44976,N_44623,N_44677);
and U44977 (N_44977,N_44661,N_44539);
xnor U44978 (N_44978,N_44656,N_44538);
or U44979 (N_44979,N_44654,N_44571);
or U44980 (N_44980,N_44695,N_44522);
xnor U44981 (N_44981,N_44658,N_44716);
and U44982 (N_44982,N_44639,N_44731);
or U44983 (N_44983,N_44746,N_44511);
nor U44984 (N_44984,N_44719,N_44509);
and U44985 (N_44985,N_44624,N_44585);
and U44986 (N_44986,N_44561,N_44589);
nand U44987 (N_44987,N_44604,N_44617);
and U44988 (N_44988,N_44528,N_44584);
or U44989 (N_44989,N_44747,N_44578);
and U44990 (N_44990,N_44653,N_44730);
or U44991 (N_44991,N_44537,N_44620);
nand U44992 (N_44992,N_44738,N_44709);
or U44993 (N_44993,N_44517,N_44714);
nor U44994 (N_44994,N_44628,N_44609);
nand U44995 (N_44995,N_44654,N_44519);
xor U44996 (N_44996,N_44567,N_44593);
xnor U44997 (N_44997,N_44621,N_44538);
nor U44998 (N_44998,N_44604,N_44576);
nor U44999 (N_44999,N_44627,N_44618);
or U45000 (N_45000,N_44993,N_44787);
or U45001 (N_45001,N_44894,N_44974);
and U45002 (N_45002,N_44750,N_44819);
and U45003 (N_45003,N_44906,N_44922);
nor U45004 (N_45004,N_44963,N_44961);
nand U45005 (N_45005,N_44820,N_44921);
or U45006 (N_45006,N_44982,N_44970);
nand U45007 (N_45007,N_44941,N_44966);
or U45008 (N_45008,N_44756,N_44859);
xor U45009 (N_45009,N_44927,N_44850);
xnor U45010 (N_45010,N_44962,N_44769);
nor U45011 (N_45011,N_44886,N_44931);
and U45012 (N_45012,N_44971,N_44786);
or U45013 (N_45013,N_44910,N_44918);
nor U45014 (N_45014,N_44881,N_44945);
nand U45015 (N_45015,N_44915,N_44823);
xor U45016 (N_45016,N_44866,N_44847);
and U45017 (N_45017,N_44867,N_44813);
and U45018 (N_45018,N_44784,N_44979);
nor U45019 (N_45019,N_44842,N_44994);
nor U45020 (N_45020,N_44815,N_44925);
xor U45021 (N_45021,N_44800,N_44919);
or U45022 (N_45022,N_44855,N_44949);
and U45023 (N_45023,N_44934,N_44980);
or U45024 (N_45024,N_44990,N_44870);
and U45025 (N_45025,N_44903,N_44871);
and U45026 (N_45026,N_44896,N_44969);
xor U45027 (N_45027,N_44935,N_44795);
nand U45028 (N_45028,N_44785,N_44812);
or U45029 (N_45029,N_44835,N_44798);
or U45030 (N_45030,N_44774,N_44838);
xnor U45031 (N_45031,N_44834,N_44808);
and U45032 (N_45032,N_44865,N_44811);
nand U45033 (N_45033,N_44860,N_44929);
xnor U45034 (N_45034,N_44981,N_44873);
xnor U45035 (N_45035,N_44987,N_44995);
and U45036 (N_45036,N_44939,N_44964);
nand U45037 (N_45037,N_44898,N_44879);
xnor U45038 (N_45038,N_44827,N_44766);
or U45039 (N_45039,N_44923,N_44992);
nor U45040 (N_45040,N_44846,N_44985);
xor U45041 (N_45041,N_44833,N_44796);
or U45042 (N_45042,N_44897,N_44950);
and U45043 (N_45043,N_44912,N_44967);
xor U45044 (N_45044,N_44991,N_44791);
xnor U45045 (N_45045,N_44762,N_44928);
or U45046 (N_45046,N_44810,N_44902);
nor U45047 (N_45047,N_44862,N_44826);
nand U45048 (N_45048,N_44951,N_44771);
xnor U45049 (N_45049,N_44884,N_44764);
or U45050 (N_45050,N_44889,N_44983);
and U45051 (N_45051,N_44904,N_44809);
nand U45052 (N_45052,N_44946,N_44777);
nand U45053 (N_45053,N_44996,N_44978);
and U45054 (N_45054,N_44937,N_44909);
xor U45055 (N_45055,N_44948,N_44947);
nand U45056 (N_45056,N_44876,N_44936);
or U45057 (N_45057,N_44832,N_44958);
or U45058 (N_45058,N_44754,N_44916);
and U45059 (N_45059,N_44861,N_44752);
nand U45060 (N_45060,N_44952,N_44874);
and U45061 (N_45061,N_44887,N_44761);
or U45062 (N_45062,N_44793,N_44763);
or U45063 (N_45063,N_44779,N_44968);
xor U45064 (N_45064,N_44799,N_44882);
nor U45065 (N_45065,N_44942,N_44943);
nand U45066 (N_45066,N_44989,N_44765);
xor U45067 (N_45067,N_44758,N_44857);
nor U45068 (N_45068,N_44755,N_44869);
and U45069 (N_45069,N_44828,N_44851);
or U45070 (N_45070,N_44797,N_44933);
nor U45071 (N_45071,N_44822,N_44908);
and U45072 (N_45072,N_44893,N_44875);
xor U45073 (N_45073,N_44776,N_44790);
or U45074 (N_45074,N_44900,N_44863);
nor U45075 (N_45075,N_44794,N_44883);
xor U45076 (N_45076,N_44973,N_44830);
nor U45077 (N_45077,N_44829,N_44997);
or U45078 (N_45078,N_44770,N_44792);
nand U45079 (N_45079,N_44778,N_44926);
xor U45080 (N_45080,N_44956,N_44914);
or U45081 (N_45081,N_44804,N_44984);
nor U45082 (N_45082,N_44825,N_44901);
xor U45083 (N_45083,N_44852,N_44783);
and U45084 (N_45084,N_44781,N_44824);
and U45085 (N_45085,N_44868,N_44924);
nor U45086 (N_45086,N_44753,N_44789);
nand U45087 (N_45087,N_44805,N_44880);
or U45088 (N_45088,N_44757,N_44960);
nand U45089 (N_45089,N_44888,N_44999);
or U45090 (N_45090,N_44972,N_44891);
and U45091 (N_45091,N_44854,N_44818);
xnor U45092 (N_45092,N_44843,N_44751);
or U45093 (N_45093,N_44885,N_44816);
nor U45094 (N_45094,N_44932,N_44917);
nand U45095 (N_45095,N_44911,N_44775);
and U45096 (N_45096,N_44767,N_44976);
nor U45097 (N_45097,N_44807,N_44849);
xnor U45098 (N_45098,N_44841,N_44877);
nand U45099 (N_45099,N_44821,N_44760);
nor U45100 (N_45100,N_44892,N_44878);
or U45101 (N_45101,N_44959,N_44858);
nand U45102 (N_45102,N_44848,N_44977);
nand U45103 (N_45103,N_44930,N_44954);
or U45104 (N_45104,N_44856,N_44899);
nand U45105 (N_45105,N_44965,N_44988);
nor U45106 (N_45106,N_44782,N_44953);
and U45107 (N_45107,N_44759,N_44839);
xnor U45108 (N_45108,N_44840,N_44905);
xnor U45109 (N_45109,N_44890,N_44940);
nand U45110 (N_45110,N_44895,N_44975);
nand U45111 (N_45111,N_44802,N_44772);
nor U45112 (N_45112,N_44831,N_44872);
nor U45113 (N_45113,N_44864,N_44907);
or U45114 (N_45114,N_44773,N_44844);
and U45115 (N_45115,N_44944,N_44806);
and U45116 (N_45116,N_44998,N_44853);
nor U45117 (N_45117,N_44837,N_44788);
nor U45118 (N_45118,N_44801,N_44780);
and U45119 (N_45119,N_44836,N_44817);
and U45120 (N_45120,N_44814,N_44845);
nor U45121 (N_45121,N_44768,N_44920);
and U45122 (N_45122,N_44957,N_44803);
nor U45123 (N_45123,N_44955,N_44986);
nor U45124 (N_45124,N_44938,N_44913);
and U45125 (N_45125,N_44921,N_44806);
and U45126 (N_45126,N_44885,N_44979);
xor U45127 (N_45127,N_44793,N_44923);
xor U45128 (N_45128,N_44982,N_44851);
or U45129 (N_45129,N_44953,N_44779);
nand U45130 (N_45130,N_44939,N_44990);
and U45131 (N_45131,N_44828,N_44775);
nand U45132 (N_45132,N_44906,N_44844);
nor U45133 (N_45133,N_44758,N_44812);
nand U45134 (N_45134,N_44994,N_44929);
nor U45135 (N_45135,N_44770,N_44973);
and U45136 (N_45136,N_44869,N_44834);
xnor U45137 (N_45137,N_44903,N_44825);
nand U45138 (N_45138,N_44893,N_44851);
xnor U45139 (N_45139,N_44878,N_44983);
xor U45140 (N_45140,N_44973,N_44988);
or U45141 (N_45141,N_44874,N_44819);
nand U45142 (N_45142,N_44804,N_44759);
nor U45143 (N_45143,N_44981,N_44837);
xor U45144 (N_45144,N_44807,N_44914);
or U45145 (N_45145,N_44911,N_44882);
nand U45146 (N_45146,N_44796,N_44805);
and U45147 (N_45147,N_44880,N_44973);
and U45148 (N_45148,N_44891,N_44845);
nor U45149 (N_45149,N_44947,N_44792);
nand U45150 (N_45150,N_44919,N_44976);
or U45151 (N_45151,N_44859,N_44976);
xor U45152 (N_45152,N_44822,N_44931);
and U45153 (N_45153,N_44758,N_44839);
or U45154 (N_45154,N_44850,N_44815);
and U45155 (N_45155,N_44814,N_44960);
xnor U45156 (N_45156,N_44999,N_44833);
nor U45157 (N_45157,N_44908,N_44844);
nor U45158 (N_45158,N_44777,N_44889);
nand U45159 (N_45159,N_44921,N_44940);
or U45160 (N_45160,N_44941,N_44917);
or U45161 (N_45161,N_44798,N_44834);
and U45162 (N_45162,N_44763,N_44852);
or U45163 (N_45163,N_44836,N_44807);
and U45164 (N_45164,N_44965,N_44959);
or U45165 (N_45165,N_44755,N_44800);
and U45166 (N_45166,N_44786,N_44965);
nor U45167 (N_45167,N_44840,N_44861);
xnor U45168 (N_45168,N_44987,N_44759);
nor U45169 (N_45169,N_44871,N_44877);
or U45170 (N_45170,N_44930,N_44919);
and U45171 (N_45171,N_44968,N_44823);
and U45172 (N_45172,N_44944,N_44819);
and U45173 (N_45173,N_44795,N_44751);
xor U45174 (N_45174,N_44949,N_44756);
nand U45175 (N_45175,N_44774,N_44993);
or U45176 (N_45176,N_44790,N_44936);
nor U45177 (N_45177,N_44839,N_44763);
and U45178 (N_45178,N_44966,N_44968);
nor U45179 (N_45179,N_44815,N_44847);
or U45180 (N_45180,N_44751,N_44917);
or U45181 (N_45181,N_44858,N_44851);
nor U45182 (N_45182,N_44851,N_44939);
xnor U45183 (N_45183,N_44861,N_44806);
nor U45184 (N_45184,N_44763,N_44965);
xnor U45185 (N_45185,N_44928,N_44861);
or U45186 (N_45186,N_44791,N_44910);
or U45187 (N_45187,N_44916,N_44771);
or U45188 (N_45188,N_44916,N_44776);
or U45189 (N_45189,N_44966,N_44774);
nand U45190 (N_45190,N_44913,N_44996);
nand U45191 (N_45191,N_44936,N_44982);
and U45192 (N_45192,N_44824,N_44886);
or U45193 (N_45193,N_44989,N_44849);
nand U45194 (N_45194,N_44794,N_44983);
nor U45195 (N_45195,N_44783,N_44752);
xor U45196 (N_45196,N_44908,N_44935);
nand U45197 (N_45197,N_44783,N_44802);
xnor U45198 (N_45198,N_44760,N_44980);
or U45199 (N_45199,N_44812,N_44968);
xnor U45200 (N_45200,N_44779,N_44821);
xor U45201 (N_45201,N_44899,N_44773);
nor U45202 (N_45202,N_44993,N_44942);
or U45203 (N_45203,N_44779,N_44800);
nor U45204 (N_45204,N_44911,N_44800);
and U45205 (N_45205,N_44955,N_44794);
nand U45206 (N_45206,N_44919,N_44979);
xnor U45207 (N_45207,N_44751,N_44873);
xnor U45208 (N_45208,N_44942,N_44779);
or U45209 (N_45209,N_44959,N_44904);
and U45210 (N_45210,N_44764,N_44971);
or U45211 (N_45211,N_44872,N_44884);
nor U45212 (N_45212,N_44961,N_44813);
or U45213 (N_45213,N_44852,N_44924);
and U45214 (N_45214,N_44910,N_44835);
nand U45215 (N_45215,N_44926,N_44984);
or U45216 (N_45216,N_44848,N_44770);
nor U45217 (N_45217,N_44839,N_44987);
nand U45218 (N_45218,N_44791,N_44889);
nand U45219 (N_45219,N_44822,N_44800);
and U45220 (N_45220,N_44793,N_44831);
nand U45221 (N_45221,N_44797,N_44981);
xor U45222 (N_45222,N_44785,N_44981);
nand U45223 (N_45223,N_44808,N_44894);
nand U45224 (N_45224,N_44859,N_44778);
xor U45225 (N_45225,N_44905,N_44781);
and U45226 (N_45226,N_44890,N_44986);
and U45227 (N_45227,N_44836,N_44929);
nand U45228 (N_45228,N_44989,N_44973);
and U45229 (N_45229,N_44943,N_44816);
or U45230 (N_45230,N_44954,N_44990);
nand U45231 (N_45231,N_44937,N_44981);
nor U45232 (N_45232,N_44904,N_44956);
xor U45233 (N_45233,N_44927,N_44942);
nand U45234 (N_45234,N_44854,N_44855);
nor U45235 (N_45235,N_44989,N_44928);
xnor U45236 (N_45236,N_44796,N_44873);
xnor U45237 (N_45237,N_44923,N_44948);
or U45238 (N_45238,N_44905,N_44948);
nor U45239 (N_45239,N_44841,N_44918);
xor U45240 (N_45240,N_44866,N_44973);
nor U45241 (N_45241,N_44914,N_44993);
and U45242 (N_45242,N_44844,N_44910);
or U45243 (N_45243,N_44792,N_44954);
or U45244 (N_45244,N_44758,N_44790);
or U45245 (N_45245,N_44952,N_44944);
or U45246 (N_45246,N_44989,N_44830);
nor U45247 (N_45247,N_44905,N_44862);
and U45248 (N_45248,N_44790,N_44810);
nand U45249 (N_45249,N_44925,N_44873);
and U45250 (N_45250,N_45185,N_45163);
and U45251 (N_45251,N_45096,N_45094);
xnor U45252 (N_45252,N_45130,N_45069);
nor U45253 (N_45253,N_45207,N_45061);
and U45254 (N_45254,N_45161,N_45222);
nor U45255 (N_45255,N_45195,N_45008);
nand U45256 (N_45256,N_45074,N_45224);
nand U45257 (N_45257,N_45243,N_45054);
or U45258 (N_45258,N_45228,N_45165);
or U45259 (N_45259,N_45070,N_45233);
xnor U45260 (N_45260,N_45183,N_45219);
nand U45261 (N_45261,N_45138,N_45077);
xor U45262 (N_45262,N_45026,N_45153);
or U45263 (N_45263,N_45013,N_45100);
and U45264 (N_45264,N_45103,N_45089);
xnor U45265 (N_45265,N_45047,N_45134);
or U45266 (N_45266,N_45015,N_45181);
nor U45267 (N_45267,N_45162,N_45245);
and U45268 (N_45268,N_45006,N_45106);
or U45269 (N_45269,N_45009,N_45129);
xnor U45270 (N_45270,N_45202,N_45188);
or U45271 (N_45271,N_45087,N_45107);
xor U45272 (N_45272,N_45082,N_45039);
nor U45273 (N_45273,N_45223,N_45151);
nand U45274 (N_45274,N_45035,N_45218);
nor U45275 (N_45275,N_45216,N_45097);
xor U45276 (N_45276,N_45120,N_45166);
or U45277 (N_45277,N_45236,N_45158);
nor U45278 (N_45278,N_45196,N_45119);
and U45279 (N_45279,N_45164,N_45080);
or U45280 (N_45280,N_45184,N_45027);
or U45281 (N_45281,N_45237,N_45157);
nor U45282 (N_45282,N_45076,N_45174);
nand U45283 (N_45283,N_45190,N_45105);
nand U45284 (N_45284,N_45179,N_45021);
nand U45285 (N_45285,N_45104,N_45175);
xnor U45286 (N_45286,N_45121,N_45145);
nor U45287 (N_45287,N_45052,N_45149);
xnor U45288 (N_45288,N_45246,N_45221);
and U45289 (N_45289,N_45191,N_45017);
nor U45290 (N_45290,N_45143,N_45172);
nand U45291 (N_45291,N_45095,N_45232);
or U45292 (N_45292,N_45060,N_45108);
and U45293 (N_45293,N_45203,N_45059);
and U45294 (N_45294,N_45063,N_45126);
and U45295 (N_45295,N_45117,N_45018);
or U45296 (N_45296,N_45197,N_45062);
and U45297 (N_45297,N_45014,N_45199);
nor U45298 (N_45298,N_45186,N_45240);
or U45299 (N_45299,N_45213,N_45180);
or U45300 (N_45300,N_45124,N_45125);
nor U45301 (N_45301,N_45109,N_45046);
nand U45302 (N_45302,N_45156,N_45112);
and U45303 (N_45303,N_45075,N_45168);
nand U45304 (N_45304,N_45230,N_45020);
xnor U45305 (N_45305,N_45242,N_45036);
or U45306 (N_45306,N_45248,N_45030);
or U45307 (N_45307,N_45012,N_45226);
nor U45308 (N_45308,N_45155,N_45116);
and U45309 (N_45309,N_45031,N_45048);
and U45310 (N_45310,N_45065,N_45206);
or U45311 (N_45311,N_45132,N_45110);
nand U45312 (N_45312,N_45086,N_45201);
xor U45313 (N_45313,N_45167,N_45139);
nor U45314 (N_45314,N_45081,N_45205);
or U45315 (N_45315,N_45229,N_45016);
nor U45316 (N_45316,N_45022,N_45041);
xor U45317 (N_45317,N_45066,N_45144);
and U45318 (N_45318,N_45135,N_45093);
xor U45319 (N_45319,N_45211,N_45142);
xor U45320 (N_45320,N_45148,N_45025);
nor U45321 (N_45321,N_45118,N_45208);
nor U45322 (N_45322,N_45084,N_45101);
or U45323 (N_45323,N_45071,N_45212);
or U45324 (N_45324,N_45011,N_45053);
nor U45325 (N_45325,N_45136,N_45038);
nor U45326 (N_45326,N_45227,N_45235);
or U45327 (N_45327,N_45122,N_45133);
nand U45328 (N_45328,N_45241,N_45007);
nand U45329 (N_45329,N_45244,N_45249);
or U45330 (N_45330,N_45040,N_45029);
and U45331 (N_45331,N_45072,N_45160);
and U45332 (N_45332,N_45010,N_45215);
nand U45333 (N_45333,N_45150,N_45004);
nand U45334 (N_45334,N_45170,N_45019);
nand U45335 (N_45335,N_45234,N_45127);
nor U45336 (N_45336,N_45099,N_45090);
nand U45337 (N_45337,N_45003,N_45137);
xor U45338 (N_45338,N_45067,N_45173);
or U45339 (N_45339,N_45091,N_45068);
xor U45340 (N_45340,N_45050,N_45079);
xnor U45341 (N_45341,N_45177,N_45123);
and U45342 (N_45342,N_45171,N_45043);
xor U45343 (N_45343,N_45111,N_45005);
or U45344 (N_45344,N_45102,N_45152);
and U45345 (N_45345,N_45037,N_45131);
xor U45346 (N_45346,N_45033,N_45115);
nor U45347 (N_45347,N_45178,N_45189);
nand U45348 (N_45348,N_45045,N_45169);
nor U45349 (N_45349,N_45210,N_45042);
nor U45350 (N_45350,N_45092,N_45024);
xor U45351 (N_45351,N_45217,N_45114);
nor U45352 (N_45352,N_45049,N_45140);
nor U45353 (N_45353,N_45113,N_45088);
nand U45354 (N_45354,N_45051,N_45128);
xnor U45355 (N_45355,N_45055,N_45239);
or U45356 (N_45356,N_45238,N_45057);
and U45357 (N_45357,N_45247,N_45000);
nor U45358 (N_45358,N_45073,N_45085);
xnor U45359 (N_45359,N_45044,N_45141);
nor U45360 (N_45360,N_45056,N_45220);
or U45361 (N_45361,N_45058,N_45198);
xnor U45362 (N_45362,N_45146,N_45001);
xnor U45363 (N_45363,N_45002,N_45064);
xor U45364 (N_45364,N_45231,N_45209);
nor U45365 (N_45365,N_45176,N_45204);
and U45366 (N_45366,N_45225,N_45214);
or U45367 (N_45367,N_45023,N_45034);
nand U45368 (N_45368,N_45194,N_45078);
and U45369 (N_45369,N_45193,N_45032);
or U45370 (N_45370,N_45098,N_45028);
nor U45371 (N_45371,N_45159,N_45154);
xnor U45372 (N_45372,N_45083,N_45147);
and U45373 (N_45373,N_45187,N_45192);
or U45374 (N_45374,N_45200,N_45182);
nor U45375 (N_45375,N_45174,N_45145);
nor U45376 (N_45376,N_45195,N_45246);
or U45377 (N_45377,N_45232,N_45053);
and U45378 (N_45378,N_45089,N_45054);
nor U45379 (N_45379,N_45050,N_45081);
nor U45380 (N_45380,N_45083,N_45171);
nor U45381 (N_45381,N_45057,N_45054);
nand U45382 (N_45382,N_45204,N_45117);
xor U45383 (N_45383,N_45090,N_45124);
or U45384 (N_45384,N_45025,N_45119);
xnor U45385 (N_45385,N_45111,N_45075);
or U45386 (N_45386,N_45165,N_45212);
nor U45387 (N_45387,N_45133,N_45065);
nand U45388 (N_45388,N_45175,N_45173);
xnor U45389 (N_45389,N_45213,N_45129);
xor U45390 (N_45390,N_45099,N_45164);
or U45391 (N_45391,N_45041,N_45130);
xor U45392 (N_45392,N_45081,N_45001);
and U45393 (N_45393,N_45234,N_45077);
or U45394 (N_45394,N_45189,N_45195);
xor U45395 (N_45395,N_45205,N_45242);
xor U45396 (N_45396,N_45010,N_45039);
nand U45397 (N_45397,N_45112,N_45015);
or U45398 (N_45398,N_45208,N_45247);
nand U45399 (N_45399,N_45100,N_45167);
and U45400 (N_45400,N_45106,N_45029);
nor U45401 (N_45401,N_45159,N_45209);
or U45402 (N_45402,N_45038,N_45087);
xnor U45403 (N_45403,N_45231,N_45140);
nor U45404 (N_45404,N_45009,N_45025);
and U45405 (N_45405,N_45089,N_45050);
nor U45406 (N_45406,N_45062,N_45192);
or U45407 (N_45407,N_45158,N_45170);
or U45408 (N_45408,N_45199,N_45148);
or U45409 (N_45409,N_45048,N_45201);
nand U45410 (N_45410,N_45149,N_45093);
xnor U45411 (N_45411,N_45183,N_45158);
or U45412 (N_45412,N_45201,N_45078);
xor U45413 (N_45413,N_45046,N_45055);
nor U45414 (N_45414,N_45040,N_45128);
and U45415 (N_45415,N_45040,N_45196);
or U45416 (N_45416,N_45094,N_45196);
nor U45417 (N_45417,N_45093,N_45216);
or U45418 (N_45418,N_45148,N_45173);
or U45419 (N_45419,N_45009,N_45161);
nand U45420 (N_45420,N_45142,N_45039);
and U45421 (N_45421,N_45043,N_45066);
nor U45422 (N_45422,N_45157,N_45136);
nor U45423 (N_45423,N_45221,N_45210);
or U45424 (N_45424,N_45096,N_45231);
and U45425 (N_45425,N_45157,N_45188);
nand U45426 (N_45426,N_45151,N_45091);
or U45427 (N_45427,N_45223,N_45147);
nand U45428 (N_45428,N_45094,N_45229);
xnor U45429 (N_45429,N_45200,N_45093);
and U45430 (N_45430,N_45231,N_45123);
nor U45431 (N_45431,N_45194,N_45053);
nor U45432 (N_45432,N_45111,N_45207);
or U45433 (N_45433,N_45079,N_45046);
or U45434 (N_45434,N_45226,N_45247);
nand U45435 (N_45435,N_45031,N_45005);
and U45436 (N_45436,N_45037,N_45003);
and U45437 (N_45437,N_45044,N_45084);
nand U45438 (N_45438,N_45166,N_45140);
or U45439 (N_45439,N_45011,N_45217);
and U45440 (N_45440,N_45005,N_45147);
and U45441 (N_45441,N_45101,N_45077);
nor U45442 (N_45442,N_45152,N_45233);
nand U45443 (N_45443,N_45171,N_45112);
nand U45444 (N_45444,N_45067,N_45118);
and U45445 (N_45445,N_45054,N_45099);
nand U45446 (N_45446,N_45033,N_45095);
nor U45447 (N_45447,N_45145,N_45114);
nor U45448 (N_45448,N_45013,N_45092);
or U45449 (N_45449,N_45024,N_45217);
nor U45450 (N_45450,N_45065,N_45244);
and U45451 (N_45451,N_45158,N_45134);
xor U45452 (N_45452,N_45159,N_45149);
nand U45453 (N_45453,N_45110,N_45165);
xnor U45454 (N_45454,N_45241,N_45202);
and U45455 (N_45455,N_45030,N_45120);
nor U45456 (N_45456,N_45114,N_45074);
nor U45457 (N_45457,N_45126,N_45244);
or U45458 (N_45458,N_45074,N_45120);
and U45459 (N_45459,N_45070,N_45017);
and U45460 (N_45460,N_45154,N_45230);
xnor U45461 (N_45461,N_45226,N_45239);
or U45462 (N_45462,N_45208,N_45219);
or U45463 (N_45463,N_45176,N_45163);
nor U45464 (N_45464,N_45194,N_45237);
nand U45465 (N_45465,N_45128,N_45017);
nand U45466 (N_45466,N_45099,N_45041);
nand U45467 (N_45467,N_45117,N_45145);
and U45468 (N_45468,N_45026,N_45147);
or U45469 (N_45469,N_45152,N_45243);
xor U45470 (N_45470,N_45020,N_45121);
nand U45471 (N_45471,N_45098,N_45220);
nand U45472 (N_45472,N_45233,N_45213);
or U45473 (N_45473,N_45045,N_45092);
and U45474 (N_45474,N_45158,N_45076);
xnor U45475 (N_45475,N_45169,N_45219);
xor U45476 (N_45476,N_45051,N_45138);
xor U45477 (N_45477,N_45046,N_45133);
nor U45478 (N_45478,N_45206,N_45058);
nand U45479 (N_45479,N_45225,N_45236);
xnor U45480 (N_45480,N_45006,N_45027);
or U45481 (N_45481,N_45143,N_45097);
xnor U45482 (N_45482,N_45170,N_45223);
nor U45483 (N_45483,N_45015,N_45177);
xor U45484 (N_45484,N_45062,N_45185);
nand U45485 (N_45485,N_45143,N_45053);
xnor U45486 (N_45486,N_45081,N_45036);
and U45487 (N_45487,N_45094,N_45186);
and U45488 (N_45488,N_45214,N_45243);
nand U45489 (N_45489,N_45077,N_45033);
nor U45490 (N_45490,N_45185,N_45183);
and U45491 (N_45491,N_45105,N_45195);
nand U45492 (N_45492,N_45178,N_45237);
and U45493 (N_45493,N_45160,N_45137);
nor U45494 (N_45494,N_45063,N_45080);
xor U45495 (N_45495,N_45211,N_45180);
or U45496 (N_45496,N_45110,N_45238);
and U45497 (N_45497,N_45217,N_45106);
and U45498 (N_45498,N_45132,N_45002);
and U45499 (N_45499,N_45226,N_45122);
nand U45500 (N_45500,N_45293,N_45417);
and U45501 (N_45501,N_45474,N_45262);
nor U45502 (N_45502,N_45275,N_45376);
nand U45503 (N_45503,N_45327,N_45296);
nor U45504 (N_45504,N_45315,N_45395);
or U45505 (N_45505,N_45496,N_45314);
or U45506 (N_45506,N_45398,N_45432);
nor U45507 (N_45507,N_45351,N_45326);
nand U45508 (N_45508,N_45362,N_45464);
or U45509 (N_45509,N_45333,N_45435);
and U45510 (N_45510,N_45388,N_45423);
and U45511 (N_45511,N_45345,N_45468);
nand U45512 (N_45512,N_45456,N_45465);
and U45513 (N_45513,N_45355,N_45338);
or U45514 (N_45514,N_45318,N_45305);
nor U45515 (N_45515,N_45389,N_45348);
or U45516 (N_45516,N_45476,N_45286);
nand U45517 (N_45517,N_45467,N_45431);
nor U45518 (N_45518,N_45434,N_45304);
or U45519 (N_45519,N_45416,N_45442);
and U45520 (N_45520,N_45352,N_45258);
xor U45521 (N_45521,N_45270,N_45320);
nand U45522 (N_45522,N_45340,N_45344);
nand U45523 (N_45523,N_45329,N_45382);
nand U45524 (N_45524,N_45331,N_45366);
nand U45525 (N_45525,N_45273,N_45453);
nand U45526 (N_45526,N_45306,N_45353);
nor U45527 (N_45527,N_45260,N_45299);
and U45528 (N_45528,N_45438,N_45291);
nor U45529 (N_45529,N_45290,N_45497);
and U45530 (N_45530,N_45365,N_45325);
and U45531 (N_45531,N_45261,N_45254);
xnor U45532 (N_45532,N_45408,N_45415);
or U45533 (N_45533,N_45498,N_45283);
xnor U45534 (N_45534,N_45302,N_45419);
nor U45535 (N_45535,N_45390,N_45268);
xor U45536 (N_45536,N_45354,N_45328);
or U45537 (N_45537,N_45255,N_45343);
nor U45538 (N_45538,N_45281,N_45256);
xnor U45539 (N_45539,N_45396,N_45317);
xnor U45540 (N_45540,N_45363,N_45387);
and U45541 (N_45541,N_45466,N_45452);
and U45542 (N_45542,N_45335,N_45319);
nor U45543 (N_45543,N_45364,N_45459);
or U45544 (N_45544,N_45428,N_45359);
and U45545 (N_45545,N_45263,N_45265);
and U45546 (N_45546,N_45490,N_45371);
nand U45547 (N_45547,N_45393,N_45368);
nor U45548 (N_45548,N_45369,N_45404);
and U45549 (N_45549,N_45410,N_45485);
nand U45550 (N_45550,N_45479,N_45370);
nor U45551 (N_45551,N_45483,N_45321);
and U45552 (N_45552,N_45384,N_45400);
and U45553 (N_45553,N_45413,N_45334);
nand U45554 (N_45554,N_45269,N_45499);
and U45555 (N_45555,N_45449,N_45406);
nand U45556 (N_45556,N_45385,N_45494);
or U45557 (N_45557,N_45424,N_45392);
nor U45558 (N_45558,N_45285,N_45295);
or U45559 (N_45559,N_45477,N_45422);
xnor U45560 (N_45560,N_45332,N_45342);
xor U45561 (N_45561,N_45303,N_45357);
xnor U45562 (N_45562,N_45257,N_45475);
or U45563 (N_45563,N_45267,N_45349);
or U45564 (N_45564,N_45309,N_45284);
nand U45565 (N_45565,N_45460,N_45391);
or U45566 (N_45566,N_45488,N_45436);
nor U45567 (N_45567,N_45324,N_45307);
nand U45568 (N_45568,N_45397,N_45380);
nand U45569 (N_45569,N_45405,N_45493);
nand U45570 (N_45570,N_45446,N_45308);
nand U45571 (N_45571,N_45420,N_45276);
nand U45572 (N_45572,N_45495,N_45469);
nor U45573 (N_45573,N_45311,N_45280);
or U45574 (N_45574,N_45418,N_45367);
xor U45575 (N_45575,N_45358,N_45292);
xor U45576 (N_45576,N_45409,N_45489);
xor U45577 (N_45577,N_45282,N_45486);
nand U45578 (N_45578,N_45289,N_45350);
nor U45579 (N_45579,N_45300,N_45401);
nor U45580 (N_45580,N_45274,N_45378);
nand U45581 (N_45581,N_45288,N_45430);
nor U45582 (N_45582,N_45484,N_45414);
xor U45583 (N_45583,N_45341,N_45373);
nor U45584 (N_45584,N_45441,N_45473);
and U45585 (N_45585,N_45425,N_45330);
nor U45586 (N_45586,N_45279,N_45381);
nand U45587 (N_45587,N_45454,N_45323);
nand U45588 (N_45588,N_45437,N_45451);
nand U45589 (N_45589,N_45375,N_45412);
and U45590 (N_45590,N_45471,N_45462);
and U45591 (N_45591,N_45360,N_45266);
nand U45592 (N_45592,N_45251,N_45339);
nor U45593 (N_45593,N_45347,N_45356);
or U45594 (N_45594,N_45287,N_45337);
or U45595 (N_45595,N_45379,N_45407);
and U45596 (N_45596,N_45259,N_45411);
or U45597 (N_45597,N_45377,N_45481);
and U45598 (N_45598,N_45250,N_45458);
nand U45599 (N_45599,N_45336,N_45253);
xnor U45600 (N_45600,N_45346,N_45448);
and U45601 (N_45601,N_45252,N_45482);
nand U45602 (N_45602,N_45470,N_45264);
or U45603 (N_45603,N_45383,N_45278);
nor U45604 (N_45604,N_45301,N_45297);
and U45605 (N_45605,N_45272,N_45310);
nor U45606 (N_45606,N_45421,N_45426);
or U45607 (N_45607,N_45487,N_45316);
nand U45608 (N_45608,N_45294,N_45374);
nor U45609 (N_45609,N_45386,N_45361);
and U45610 (N_45610,N_45492,N_45457);
xnor U45611 (N_45611,N_45402,N_45440);
xnor U45612 (N_45612,N_45399,N_45443);
or U45613 (N_45613,N_45394,N_45429);
nor U45614 (N_45614,N_45298,N_45444);
xnor U45615 (N_45615,N_45271,N_45427);
and U45616 (N_45616,N_45455,N_45372);
nor U45617 (N_45617,N_45491,N_45478);
nand U45618 (N_45618,N_45439,N_45403);
nor U45619 (N_45619,N_45450,N_45277);
nand U45620 (N_45620,N_45313,N_45445);
and U45621 (N_45621,N_45480,N_45322);
and U45622 (N_45622,N_45312,N_45447);
nor U45623 (N_45623,N_45463,N_45472);
nand U45624 (N_45624,N_45461,N_45433);
xnor U45625 (N_45625,N_45421,N_45364);
xnor U45626 (N_45626,N_45404,N_45343);
nand U45627 (N_45627,N_45254,N_45390);
nor U45628 (N_45628,N_45310,N_45259);
xor U45629 (N_45629,N_45256,N_45343);
or U45630 (N_45630,N_45313,N_45355);
nor U45631 (N_45631,N_45460,N_45373);
and U45632 (N_45632,N_45298,N_45466);
nor U45633 (N_45633,N_45379,N_45451);
and U45634 (N_45634,N_45312,N_45432);
and U45635 (N_45635,N_45407,N_45341);
nand U45636 (N_45636,N_45477,N_45448);
nor U45637 (N_45637,N_45409,N_45293);
nand U45638 (N_45638,N_45405,N_45435);
nand U45639 (N_45639,N_45395,N_45254);
nand U45640 (N_45640,N_45422,N_45299);
and U45641 (N_45641,N_45477,N_45494);
xor U45642 (N_45642,N_45432,N_45399);
xor U45643 (N_45643,N_45344,N_45398);
xor U45644 (N_45644,N_45320,N_45278);
and U45645 (N_45645,N_45355,N_45443);
or U45646 (N_45646,N_45445,N_45387);
nor U45647 (N_45647,N_45462,N_45390);
nand U45648 (N_45648,N_45367,N_45436);
xor U45649 (N_45649,N_45295,N_45369);
nand U45650 (N_45650,N_45460,N_45432);
nand U45651 (N_45651,N_45300,N_45374);
xnor U45652 (N_45652,N_45281,N_45363);
or U45653 (N_45653,N_45489,N_45386);
or U45654 (N_45654,N_45386,N_45434);
or U45655 (N_45655,N_45466,N_45250);
nand U45656 (N_45656,N_45408,N_45488);
xor U45657 (N_45657,N_45437,N_45266);
nor U45658 (N_45658,N_45407,N_45336);
or U45659 (N_45659,N_45460,N_45429);
or U45660 (N_45660,N_45318,N_45339);
nor U45661 (N_45661,N_45257,N_45325);
xnor U45662 (N_45662,N_45408,N_45395);
or U45663 (N_45663,N_45296,N_45415);
and U45664 (N_45664,N_45306,N_45252);
xnor U45665 (N_45665,N_45449,N_45429);
and U45666 (N_45666,N_45452,N_45426);
nor U45667 (N_45667,N_45434,N_45270);
or U45668 (N_45668,N_45253,N_45294);
nor U45669 (N_45669,N_45310,N_45422);
and U45670 (N_45670,N_45330,N_45362);
nand U45671 (N_45671,N_45416,N_45253);
xor U45672 (N_45672,N_45303,N_45347);
or U45673 (N_45673,N_45279,N_45278);
and U45674 (N_45674,N_45332,N_45372);
nand U45675 (N_45675,N_45435,N_45288);
nand U45676 (N_45676,N_45312,N_45413);
and U45677 (N_45677,N_45412,N_45409);
or U45678 (N_45678,N_45465,N_45414);
nand U45679 (N_45679,N_45416,N_45472);
xnor U45680 (N_45680,N_45377,N_45469);
and U45681 (N_45681,N_45313,N_45485);
and U45682 (N_45682,N_45316,N_45299);
or U45683 (N_45683,N_45315,N_45479);
or U45684 (N_45684,N_45448,N_45301);
or U45685 (N_45685,N_45277,N_45494);
or U45686 (N_45686,N_45275,N_45439);
and U45687 (N_45687,N_45371,N_45327);
nand U45688 (N_45688,N_45312,N_45290);
and U45689 (N_45689,N_45438,N_45344);
and U45690 (N_45690,N_45384,N_45392);
or U45691 (N_45691,N_45250,N_45362);
and U45692 (N_45692,N_45461,N_45298);
or U45693 (N_45693,N_45436,N_45256);
or U45694 (N_45694,N_45416,N_45478);
or U45695 (N_45695,N_45276,N_45291);
and U45696 (N_45696,N_45311,N_45454);
and U45697 (N_45697,N_45465,N_45326);
nand U45698 (N_45698,N_45383,N_45456);
nand U45699 (N_45699,N_45275,N_45284);
or U45700 (N_45700,N_45344,N_45475);
nor U45701 (N_45701,N_45333,N_45482);
nor U45702 (N_45702,N_45445,N_45330);
and U45703 (N_45703,N_45376,N_45411);
nand U45704 (N_45704,N_45491,N_45352);
nor U45705 (N_45705,N_45277,N_45267);
or U45706 (N_45706,N_45296,N_45471);
xor U45707 (N_45707,N_45438,N_45385);
nand U45708 (N_45708,N_45361,N_45394);
and U45709 (N_45709,N_45294,N_45495);
nor U45710 (N_45710,N_45277,N_45337);
and U45711 (N_45711,N_45482,N_45495);
nand U45712 (N_45712,N_45278,N_45426);
xor U45713 (N_45713,N_45344,N_45325);
nor U45714 (N_45714,N_45393,N_45457);
nand U45715 (N_45715,N_45258,N_45428);
xor U45716 (N_45716,N_45366,N_45360);
and U45717 (N_45717,N_45378,N_45263);
or U45718 (N_45718,N_45312,N_45488);
xor U45719 (N_45719,N_45458,N_45374);
xor U45720 (N_45720,N_45295,N_45286);
nand U45721 (N_45721,N_45416,N_45251);
nand U45722 (N_45722,N_45436,N_45457);
nand U45723 (N_45723,N_45382,N_45287);
nor U45724 (N_45724,N_45310,N_45389);
or U45725 (N_45725,N_45343,N_45401);
or U45726 (N_45726,N_45337,N_45372);
nand U45727 (N_45727,N_45428,N_45391);
xor U45728 (N_45728,N_45479,N_45311);
or U45729 (N_45729,N_45416,N_45267);
xor U45730 (N_45730,N_45393,N_45263);
and U45731 (N_45731,N_45489,N_45260);
and U45732 (N_45732,N_45464,N_45492);
nor U45733 (N_45733,N_45368,N_45461);
nand U45734 (N_45734,N_45473,N_45360);
nor U45735 (N_45735,N_45384,N_45406);
or U45736 (N_45736,N_45432,N_45423);
xor U45737 (N_45737,N_45281,N_45327);
nor U45738 (N_45738,N_45456,N_45426);
xor U45739 (N_45739,N_45459,N_45481);
xor U45740 (N_45740,N_45484,N_45496);
nand U45741 (N_45741,N_45295,N_45263);
or U45742 (N_45742,N_45401,N_45375);
nor U45743 (N_45743,N_45387,N_45318);
or U45744 (N_45744,N_45278,N_45413);
nor U45745 (N_45745,N_45499,N_45382);
and U45746 (N_45746,N_45261,N_45268);
or U45747 (N_45747,N_45339,N_45498);
and U45748 (N_45748,N_45418,N_45283);
xor U45749 (N_45749,N_45297,N_45283);
nor U45750 (N_45750,N_45734,N_45743);
nand U45751 (N_45751,N_45503,N_45737);
nand U45752 (N_45752,N_45541,N_45604);
xnor U45753 (N_45753,N_45622,N_45581);
and U45754 (N_45754,N_45525,N_45689);
and U45755 (N_45755,N_45579,N_45521);
and U45756 (N_45756,N_45654,N_45542);
and U45757 (N_45757,N_45509,N_45739);
and U45758 (N_45758,N_45562,N_45742);
or U45759 (N_45759,N_45502,N_45520);
nor U45760 (N_45760,N_45728,N_45678);
xor U45761 (N_45761,N_45527,N_45740);
xor U45762 (N_45762,N_45582,N_45557);
or U45763 (N_45763,N_45567,N_45636);
and U45764 (N_45764,N_45675,N_45645);
nand U45765 (N_45765,N_45669,N_45656);
nor U45766 (N_45766,N_45580,N_45644);
or U45767 (N_45767,N_45611,N_45613);
xor U45768 (N_45768,N_45570,N_45540);
xnor U45769 (N_45769,N_45606,N_45731);
nand U45770 (N_45770,N_45518,N_45549);
nor U45771 (N_45771,N_45507,N_45707);
nor U45772 (N_45772,N_45664,N_45730);
xor U45773 (N_45773,N_45617,N_45620);
xnor U45774 (N_45774,N_45663,N_45607);
nand U45775 (N_45775,N_45724,N_45523);
nor U45776 (N_45776,N_45706,N_45646);
nand U45777 (N_45777,N_45539,N_45717);
and U45778 (N_45778,N_45558,N_45632);
nand U45779 (N_45779,N_45688,N_45577);
xnor U45780 (N_45780,N_45538,N_45587);
or U45781 (N_45781,N_45714,N_45741);
nor U45782 (N_45782,N_45735,N_45528);
and U45783 (N_45783,N_45594,N_45681);
and U45784 (N_45784,N_45744,N_45680);
nor U45785 (N_45785,N_45510,N_45533);
xor U45786 (N_45786,N_45660,N_45517);
xor U45787 (N_45787,N_45610,N_45713);
and U45788 (N_45788,N_45627,N_45552);
xnor U45789 (N_45789,N_45554,N_45522);
and U45790 (N_45790,N_45519,N_45595);
nor U45791 (N_45791,N_45710,N_45624);
nor U45792 (N_45792,N_45516,N_45605);
xnor U45793 (N_45793,N_45532,N_45619);
xnor U45794 (N_45794,N_45727,N_45609);
or U45795 (N_45795,N_45667,N_45618);
nand U45796 (N_45796,N_45708,N_45561);
and U45797 (N_45797,N_45563,N_45653);
or U45798 (N_45798,N_45531,N_45512);
nor U45799 (N_45799,N_45679,N_45640);
or U45800 (N_45800,N_45631,N_45535);
nor U45801 (N_45801,N_45709,N_45593);
nand U45802 (N_45802,N_45665,N_45677);
xnor U45803 (N_45803,N_45591,N_45712);
or U45804 (N_45804,N_45504,N_45629);
or U45805 (N_45805,N_45699,N_45560);
or U45806 (N_45806,N_45749,N_45583);
nor U45807 (N_45807,N_45530,N_45571);
xnor U45808 (N_45808,N_45686,N_45578);
or U45809 (N_45809,N_45576,N_45553);
nor U45810 (N_45810,N_45683,N_45573);
xnor U45811 (N_45811,N_45723,N_45687);
nand U45812 (N_45812,N_45658,N_45747);
xnor U45813 (N_45813,N_45693,N_45715);
nor U45814 (N_45814,N_45536,N_45720);
xnor U45815 (N_45815,N_45659,N_45625);
and U45816 (N_45816,N_45662,N_45628);
nand U45817 (N_45817,N_45657,N_45614);
nor U45818 (N_45818,N_45633,N_45575);
nor U45819 (N_45819,N_45643,N_45716);
nor U45820 (N_45820,N_45655,N_45572);
nand U45821 (N_45821,N_45615,N_45568);
or U45822 (N_45822,N_45506,N_45634);
and U45823 (N_45823,N_45700,N_45513);
xnor U45824 (N_45824,N_45601,N_45548);
and U45825 (N_45825,N_45602,N_45703);
xor U45826 (N_45826,N_45569,N_45738);
or U45827 (N_45827,N_45585,N_45649);
xnor U45828 (N_45828,N_45729,N_45726);
and U45829 (N_45829,N_45598,N_45526);
and U45830 (N_45830,N_45725,N_45719);
nor U45831 (N_45831,N_45524,N_45685);
nand U45832 (N_45832,N_45668,N_45586);
xor U45833 (N_45833,N_45696,N_45691);
nand U45834 (N_45834,N_45596,N_45543);
and U45835 (N_45835,N_45621,N_45545);
and U45836 (N_45836,N_45555,N_45671);
and U45837 (N_45837,N_45590,N_45698);
and U45838 (N_45838,N_45746,N_45588);
nor U45839 (N_45839,N_45534,N_45565);
nor U45840 (N_45840,N_45546,N_45733);
and U45841 (N_45841,N_45559,N_45589);
or U45842 (N_45842,N_45641,N_45711);
nor U45843 (N_45843,N_45603,N_45702);
or U45844 (N_45844,N_45648,N_45718);
nand U45845 (N_45845,N_45666,N_45623);
nand U45846 (N_45846,N_45682,N_45550);
xnor U45847 (N_45847,N_45574,N_45630);
and U45848 (N_45848,N_45508,N_45564);
and U45849 (N_45849,N_45612,N_45600);
or U45850 (N_45850,N_45650,N_45676);
nor U45851 (N_45851,N_45566,N_45704);
nand U45852 (N_45852,N_45511,N_45695);
and U45853 (N_45853,N_45690,N_45616);
xor U45854 (N_45854,N_45529,N_45501);
xor U45855 (N_45855,N_45652,N_45748);
xnor U45856 (N_45856,N_45647,N_45692);
xnor U45857 (N_45857,N_45551,N_45544);
and U45858 (N_45858,N_45697,N_45642);
xor U45859 (N_45859,N_45637,N_45672);
and U45860 (N_45860,N_45661,N_45673);
or U45861 (N_45861,N_45736,N_45694);
xor U45862 (N_45862,N_45639,N_45592);
nand U45863 (N_45863,N_45626,N_45670);
and U45864 (N_45864,N_45597,N_45721);
nor U45865 (N_45865,N_45745,N_45515);
or U45866 (N_45866,N_45635,N_45705);
nor U45867 (N_45867,N_45608,N_45732);
or U45868 (N_45868,N_45638,N_45651);
xor U45869 (N_45869,N_45537,N_45505);
or U45870 (N_45870,N_45584,N_45547);
and U45871 (N_45871,N_45722,N_45514);
nor U45872 (N_45872,N_45674,N_45701);
xnor U45873 (N_45873,N_45500,N_45684);
nor U45874 (N_45874,N_45556,N_45599);
or U45875 (N_45875,N_45527,N_45573);
xor U45876 (N_45876,N_45616,N_45618);
nand U45877 (N_45877,N_45510,N_45541);
nor U45878 (N_45878,N_45622,N_45668);
nor U45879 (N_45879,N_45566,N_45740);
nor U45880 (N_45880,N_45724,N_45604);
nand U45881 (N_45881,N_45688,N_45642);
and U45882 (N_45882,N_45521,N_45669);
and U45883 (N_45883,N_45547,N_45564);
nor U45884 (N_45884,N_45552,N_45575);
and U45885 (N_45885,N_45618,N_45549);
and U45886 (N_45886,N_45588,N_45661);
nand U45887 (N_45887,N_45543,N_45572);
xor U45888 (N_45888,N_45682,N_45740);
or U45889 (N_45889,N_45709,N_45574);
nand U45890 (N_45890,N_45724,N_45649);
nor U45891 (N_45891,N_45696,N_45684);
nand U45892 (N_45892,N_45679,N_45505);
xnor U45893 (N_45893,N_45546,N_45596);
nor U45894 (N_45894,N_45512,N_45582);
nand U45895 (N_45895,N_45637,N_45576);
and U45896 (N_45896,N_45645,N_45627);
xor U45897 (N_45897,N_45662,N_45597);
nor U45898 (N_45898,N_45658,N_45633);
nor U45899 (N_45899,N_45590,N_45663);
nand U45900 (N_45900,N_45715,N_45585);
xor U45901 (N_45901,N_45579,N_45659);
xor U45902 (N_45902,N_45602,N_45636);
or U45903 (N_45903,N_45571,N_45503);
nand U45904 (N_45904,N_45622,N_45713);
nor U45905 (N_45905,N_45615,N_45714);
nand U45906 (N_45906,N_45519,N_45622);
nand U45907 (N_45907,N_45724,N_45733);
and U45908 (N_45908,N_45670,N_45706);
and U45909 (N_45909,N_45548,N_45564);
nor U45910 (N_45910,N_45593,N_45641);
xnor U45911 (N_45911,N_45604,N_45649);
nor U45912 (N_45912,N_45651,N_45542);
and U45913 (N_45913,N_45515,N_45675);
nor U45914 (N_45914,N_45626,N_45571);
or U45915 (N_45915,N_45732,N_45738);
xnor U45916 (N_45916,N_45573,N_45649);
xor U45917 (N_45917,N_45606,N_45675);
xor U45918 (N_45918,N_45623,N_45545);
or U45919 (N_45919,N_45500,N_45562);
nor U45920 (N_45920,N_45590,N_45602);
nor U45921 (N_45921,N_45525,N_45715);
nor U45922 (N_45922,N_45701,N_45506);
nor U45923 (N_45923,N_45507,N_45521);
nand U45924 (N_45924,N_45697,N_45566);
nand U45925 (N_45925,N_45540,N_45664);
nor U45926 (N_45926,N_45614,N_45671);
and U45927 (N_45927,N_45707,N_45701);
and U45928 (N_45928,N_45553,N_45568);
nor U45929 (N_45929,N_45713,N_45501);
xnor U45930 (N_45930,N_45539,N_45696);
xor U45931 (N_45931,N_45744,N_45547);
and U45932 (N_45932,N_45501,N_45723);
xor U45933 (N_45933,N_45586,N_45583);
xnor U45934 (N_45934,N_45524,N_45577);
xnor U45935 (N_45935,N_45514,N_45518);
nor U45936 (N_45936,N_45546,N_45567);
nor U45937 (N_45937,N_45637,N_45504);
nor U45938 (N_45938,N_45694,N_45524);
nand U45939 (N_45939,N_45739,N_45721);
xnor U45940 (N_45940,N_45745,N_45691);
nand U45941 (N_45941,N_45651,N_45686);
nor U45942 (N_45942,N_45644,N_45561);
and U45943 (N_45943,N_45529,N_45650);
nor U45944 (N_45944,N_45518,N_45728);
nor U45945 (N_45945,N_45523,N_45687);
nand U45946 (N_45946,N_45604,N_45616);
or U45947 (N_45947,N_45652,N_45656);
or U45948 (N_45948,N_45654,N_45668);
xnor U45949 (N_45949,N_45604,N_45560);
nand U45950 (N_45950,N_45625,N_45737);
xor U45951 (N_45951,N_45509,N_45639);
nor U45952 (N_45952,N_45675,N_45548);
or U45953 (N_45953,N_45620,N_45598);
and U45954 (N_45954,N_45666,N_45523);
or U45955 (N_45955,N_45631,N_45683);
nor U45956 (N_45956,N_45525,N_45660);
nor U45957 (N_45957,N_45740,N_45652);
and U45958 (N_45958,N_45554,N_45679);
nand U45959 (N_45959,N_45622,N_45601);
or U45960 (N_45960,N_45593,N_45746);
nor U45961 (N_45961,N_45615,N_45500);
nand U45962 (N_45962,N_45674,N_45602);
nand U45963 (N_45963,N_45560,N_45621);
xnor U45964 (N_45964,N_45569,N_45546);
xnor U45965 (N_45965,N_45649,N_45653);
nor U45966 (N_45966,N_45648,N_45716);
and U45967 (N_45967,N_45651,N_45698);
and U45968 (N_45968,N_45748,N_45626);
and U45969 (N_45969,N_45576,N_45525);
xnor U45970 (N_45970,N_45619,N_45609);
nor U45971 (N_45971,N_45613,N_45607);
and U45972 (N_45972,N_45627,N_45573);
xnor U45973 (N_45973,N_45568,N_45592);
nand U45974 (N_45974,N_45697,N_45689);
nand U45975 (N_45975,N_45701,N_45659);
or U45976 (N_45976,N_45503,N_45626);
xor U45977 (N_45977,N_45508,N_45636);
or U45978 (N_45978,N_45506,N_45682);
and U45979 (N_45979,N_45533,N_45736);
and U45980 (N_45980,N_45573,N_45609);
xor U45981 (N_45981,N_45713,N_45611);
nor U45982 (N_45982,N_45670,N_45585);
xor U45983 (N_45983,N_45624,N_45598);
xor U45984 (N_45984,N_45590,N_45737);
nor U45985 (N_45985,N_45667,N_45513);
and U45986 (N_45986,N_45668,N_45537);
and U45987 (N_45987,N_45721,N_45664);
nor U45988 (N_45988,N_45539,N_45650);
nor U45989 (N_45989,N_45528,N_45553);
nand U45990 (N_45990,N_45584,N_45665);
nor U45991 (N_45991,N_45574,N_45530);
and U45992 (N_45992,N_45672,N_45686);
and U45993 (N_45993,N_45704,N_45615);
nand U45994 (N_45994,N_45556,N_45711);
nor U45995 (N_45995,N_45613,N_45530);
xor U45996 (N_45996,N_45621,N_45610);
and U45997 (N_45997,N_45559,N_45549);
xnor U45998 (N_45998,N_45544,N_45721);
nand U45999 (N_45999,N_45700,N_45604);
and U46000 (N_46000,N_45804,N_45834);
or U46001 (N_46001,N_45977,N_45825);
nand U46002 (N_46002,N_45894,N_45895);
xor U46003 (N_46003,N_45753,N_45822);
or U46004 (N_46004,N_45925,N_45868);
and U46005 (N_46005,N_45930,N_45833);
nand U46006 (N_46006,N_45964,N_45828);
xor U46007 (N_46007,N_45867,N_45896);
nand U46008 (N_46008,N_45952,N_45765);
xnor U46009 (N_46009,N_45794,N_45941);
or U46010 (N_46010,N_45821,N_45806);
xor U46011 (N_46011,N_45876,N_45835);
nand U46012 (N_46012,N_45937,N_45967);
and U46013 (N_46013,N_45798,N_45864);
nand U46014 (N_46014,N_45796,N_45877);
xnor U46015 (N_46015,N_45926,N_45899);
or U46016 (N_46016,N_45792,N_45968);
nor U46017 (N_46017,N_45751,N_45989);
nand U46018 (N_46018,N_45903,N_45971);
nand U46019 (N_46019,N_45756,N_45959);
nor U46020 (N_46020,N_45900,N_45776);
xor U46021 (N_46021,N_45901,N_45815);
xor U46022 (N_46022,N_45832,N_45783);
nor U46023 (N_46023,N_45869,N_45788);
nor U46024 (N_46024,N_45784,N_45885);
xnor U46025 (N_46025,N_45942,N_45778);
or U46026 (N_46026,N_45816,N_45947);
or U46027 (N_46027,N_45787,N_45759);
or U46028 (N_46028,N_45781,N_45923);
xor U46029 (N_46029,N_45767,N_45860);
nor U46030 (N_46030,N_45924,N_45880);
xnor U46031 (N_46031,N_45865,N_45764);
xor U46032 (N_46032,N_45789,N_45760);
and U46033 (N_46033,N_45909,N_45824);
and U46034 (N_46034,N_45809,N_45881);
xnor U46035 (N_46035,N_45842,N_45954);
nand U46036 (N_46036,N_45987,N_45906);
xor U46037 (N_46037,N_45803,N_45916);
nand U46038 (N_46038,N_45827,N_45761);
and U46039 (N_46039,N_45862,N_45848);
and U46040 (N_46040,N_45779,N_45855);
nor U46041 (N_46041,N_45859,N_45893);
nor U46042 (N_46042,N_45863,N_45852);
nand U46043 (N_46043,N_45960,N_45939);
nand U46044 (N_46044,N_45938,N_45853);
or U46045 (N_46045,N_45995,N_45912);
xnor U46046 (N_46046,N_45870,N_45873);
nor U46047 (N_46047,N_45973,N_45883);
nor U46048 (N_46048,N_45858,N_45999);
nor U46049 (N_46049,N_45770,N_45935);
nand U46050 (N_46050,N_45996,N_45969);
nor U46051 (N_46051,N_45990,N_45850);
nand U46052 (N_46052,N_45892,N_45799);
or U46053 (N_46053,N_45948,N_45826);
and U46054 (N_46054,N_45975,N_45933);
or U46055 (N_46055,N_45802,N_45946);
nand U46056 (N_46056,N_45819,N_45890);
and U46057 (N_46057,N_45800,N_45914);
and U46058 (N_46058,N_45985,N_45981);
and U46059 (N_46059,N_45974,N_45979);
and U46060 (N_46060,N_45843,N_45762);
nor U46061 (N_46061,N_45978,N_45904);
xor U46062 (N_46062,N_45884,N_45919);
nand U46063 (N_46063,N_45920,N_45889);
xor U46064 (N_46064,N_45943,N_45829);
nand U46065 (N_46065,N_45810,N_45774);
xnor U46066 (N_46066,N_45839,N_45982);
nor U46067 (N_46067,N_45849,N_45993);
nor U46068 (N_46068,N_45811,N_45992);
and U46069 (N_46069,N_45929,N_45963);
nand U46070 (N_46070,N_45763,N_45908);
nand U46071 (N_46071,N_45813,N_45980);
nor U46072 (N_46072,N_45936,N_45998);
nand U46073 (N_46073,N_45991,N_45951);
xor U46074 (N_46074,N_45861,N_45988);
xnor U46075 (N_46075,N_45797,N_45915);
or U46076 (N_46076,N_45931,N_45805);
nor U46077 (N_46077,N_45782,N_45891);
nor U46078 (N_46078,N_45949,N_45888);
nand U46079 (N_46079,N_45965,N_45785);
nor U46080 (N_46080,N_45857,N_45777);
nand U46081 (N_46081,N_45754,N_45780);
or U46082 (N_46082,N_45773,N_45972);
nand U46083 (N_46083,N_45958,N_45910);
and U46084 (N_46084,N_45817,N_45932);
or U46085 (N_46085,N_45962,N_45872);
nand U46086 (N_46086,N_45838,N_45956);
nor U46087 (N_46087,N_45966,N_45944);
nor U46088 (N_46088,N_45911,N_45878);
xnor U46089 (N_46089,N_45812,N_45752);
nor U46090 (N_46090,N_45841,N_45961);
nand U46091 (N_46091,N_45757,N_45793);
nand U46092 (N_46092,N_45927,N_45918);
xor U46093 (N_46093,N_45984,N_45955);
or U46094 (N_46094,N_45879,N_45934);
nand U46095 (N_46095,N_45854,N_45928);
nand U46096 (N_46096,N_45970,N_45772);
nor U46097 (N_46097,N_45922,N_45840);
or U46098 (N_46098,N_45953,N_45801);
and U46099 (N_46099,N_45818,N_45830);
xnor U46100 (N_46100,N_45847,N_45866);
and U46101 (N_46101,N_45775,N_45814);
or U46102 (N_46102,N_45831,N_45758);
nor U46103 (N_46103,N_45875,N_45886);
nor U46104 (N_46104,N_45940,N_45887);
and U46105 (N_46105,N_45986,N_45976);
nor U46106 (N_46106,N_45913,N_45820);
xnor U46107 (N_46107,N_45856,N_45844);
or U46108 (N_46108,N_45882,N_45917);
nand U46109 (N_46109,N_45950,N_45769);
or U46110 (N_46110,N_45795,N_45790);
or U46111 (N_46111,N_45823,N_45791);
and U46112 (N_46112,N_45845,N_45994);
nand U46113 (N_46113,N_45957,N_45897);
nor U46114 (N_46114,N_45807,N_45786);
and U46115 (N_46115,N_45837,N_45768);
xnor U46116 (N_46116,N_45771,N_45874);
nor U46117 (N_46117,N_45983,N_45945);
and U46118 (N_46118,N_45871,N_45898);
and U46119 (N_46119,N_45766,N_45907);
and U46120 (N_46120,N_45750,N_45836);
nand U46121 (N_46121,N_45921,N_45846);
and U46122 (N_46122,N_45755,N_45997);
nor U46123 (N_46123,N_45808,N_45851);
nand U46124 (N_46124,N_45902,N_45905);
xor U46125 (N_46125,N_45785,N_45908);
or U46126 (N_46126,N_45957,N_45981);
or U46127 (N_46127,N_45796,N_45931);
xor U46128 (N_46128,N_45769,N_45801);
xnor U46129 (N_46129,N_45854,N_45925);
or U46130 (N_46130,N_45902,N_45827);
and U46131 (N_46131,N_45873,N_45794);
xor U46132 (N_46132,N_45856,N_45954);
nand U46133 (N_46133,N_45999,N_45838);
or U46134 (N_46134,N_45913,N_45908);
xor U46135 (N_46135,N_45983,N_45981);
or U46136 (N_46136,N_45938,N_45922);
xor U46137 (N_46137,N_45970,N_45912);
xor U46138 (N_46138,N_45781,N_45852);
and U46139 (N_46139,N_45875,N_45775);
xnor U46140 (N_46140,N_45770,N_45820);
xnor U46141 (N_46141,N_45882,N_45831);
nand U46142 (N_46142,N_45863,N_45937);
or U46143 (N_46143,N_45947,N_45982);
or U46144 (N_46144,N_45817,N_45803);
xor U46145 (N_46145,N_45922,N_45974);
nand U46146 (N_46146,N_45795,N_45887);
nor U46147 (N_46147,N_45942,N_45926);
xor U46148 (N_46148,N_45778,N_45775);
or U46149 (N_46149,N_45950,N_45909);
nand U46150 (N_46150,N_45750,N_45944);
nand U46151 (N_46151,N_45770,N_45842);
xnor U46152 (N_46152,N_45846,N_45964);
nor U46153 (N_46153,N_45834,N_45774);
nor U46154 (N_46154,N_45936,N_45860);
xnor U46155 (N_46155,N_45980,N_45856);
nand U46156 (N_46156,N_45863,N_45952);
or U46157 (N_46157,N_45809,N_45885);
or U46158 (N_46158,N_45877,N_45957);
nand U46159 (N_46159,N_45794,N_45833);
or U46160 (N_46160,N_45935,N_45954);
nor U46161 (N_46161,N_45983,N_45881);
nand U46162 (N_46162,N_45890,N_45823);
xnor U46163 (N_46163,N_45850,N_45937);
nor U46164 (N_46164,N_45753,N_45896);
nand U46165 (N_46165,N_45916,N_45784);
and U46166 (N_46166,N_45757,N_45807);
nand U46167 (N_46167,N_45788,N_45918);
nor U46168 (N_46168,N_45880,N_45872);
nor U46169 (N_46169,N_45943,N_45803);
nand U46170 (N_46170,N_45788,N_45916);
xor U46171 (N_46171,N_45857,N_45760);
and U46172 (N_46172,N_45763,N_45835);
nand U46173 (N_46173,N_45794,N_45955);
nand U46174 (N_46174,N_45881,N_45916);
and U46175 (N_46175,N_45885,N_45983);
and U46176 (N_46176,N_45822,N_45806);
xor U46177 (N_46177,N_45915,N_45972);
nor U46178 (N_46178,N_45942,N_45996);
nor U46179 (N_46179,N_45870,N_45900);
xor U46180 (N_46180,N_45881,N_45753);
nand U46181 (N_46181,N_45966,N_45908);
xor U46182 (N_46182,N_45997,N_45993);
and U46183 (N_46183,N_45945,N_45771);
and U46184 (N_46184,N_45792,N_45795);
or U46185 (N_46185,N_45766,N_45832);
nand U46186 (N_46186,N_45833,N_45877);
nand U46187 (N_46187,N_45994,N_45835);
nor U46188 (N_46188,N_45980,N_45759);
nor U46189 (N_46189,N_45898,N_45757);
xor U46190 (N_46190,N_45793,N_45907);
nand U46191 (N_46191,N_45788,N_45832);
nand U46192 (N_46192,N_45968,N_45830);
xor U46193 (N_46193,N_45985,N_45997);
nand U46194 (N_46194,N_45806,N_45945);
or U46195 (N_46195,N_45802,N_45865);
xnor U46196 (N_46196,N_45887,N_45898);
nand U46197 (N_46197,N_45820,N_45843);
and U46198 (N_46198,N_45860,N_45886);
nand U46199 (N_46199,N_45820,N_45955);
nor U46200 (N_46200,N_45750,N_45837);
nor U46201 (N_46201,N_45839,N_45983);
nor U46202 (N_46202,N_45976,N_45867);
nand U46203 (N_46203,N_45969,N_45795);
xnor U46204 (N_46204,N_45816,N_45977);
xnor U46205 (N_46205,N_45951,N_45986);
nor U46206 (N_46206,N_45803,N_45918);
xor U46207 (N_46207,N_45993,N_45796);
nor U46208 (N_46208,N_45955,N_45896);
xnor U46209 (N_46209,N_45774,N_45929);
nand U46210 (N_46210,N_45810,N_45777);
nor U46211 (N_46211,N_45886,N_45870);
xor U46212 (N_46212,N_45992,N_45937);
nand U46213 (N_46213,N_45787,N_45778);
and U46214 (N_46214,N_45984,N_45839);
nand U46215 (N_46215,N_45951,N_45948);
and U46216 (N_46216,N_45972,N_45774);
nor U46217 (N_46217,N_45918,N_45755);
nor U46218 (N_46218,N_45898,N_45817);
xor U46219 (N_46219,N_45932,N_45950);
xor U46220 (N_46220,N_45837,N_45972);
or U46221 (N_46221,N_45949,N_45889);
nor U46222 (N_46222,N_45778,N_45854);
nand U46223 (N_46223,N_45980,N_45831);
nand U46224 (N_46224,N_45750,N_45762);
nand U46225 (N_46225,N_45753,N_45961);
nor U46226 (N_46226,N_45794,N_45877);
xor U46227 (N_46227,N_45978,N_45757);
or U46228 (N_46228,N_45755,N_45900);
nand U46229 (N_46229,N_45961,N_45890);
xnor U46230 (N_46230,N_45958,N_45951);
nand U46231 (N_46231,N_45792,N_45810);
nand U46232 (N_46232,N_45954,N_45804);
xnor U46233 (N_46233,N_45921,N_45808);
nor U46234 (N_46234,N_45885,N_45822);
xor U46235 (N_46235,N_45756,N_45795);
and U46236 (N_46236,N_45910,N_45995);
xor U46237 (N_46237,N_45800,N_45963);
nand U46238 (N_46238,N_45837,N_45952);
xnor U46239 (N_46239,N_45966,N_45876);
xnor U46240 (N_46240,N_45964,N_45930);
nor U46241 (N_46241,N_45797,N_45759);
and U46242 (N_46242,N_45786,N_45815);
nand U46243 (N_46243,N_45927,N_45764);
and U46244 (N_46244,N_45773,N_45778);
nor U46245 (N_46245,N_45919,N_45866);
xor U46246 (N_46246,N_45944,N_45862);
and U46247 (N_46247,N_45891,N_45804);
and U46248 (N_46248,N_45973,N_45979);
xnor U46249 (N_46249,N_45818,N_45986);
xor U46250 (N_46250,N_46125,N_46003);
nand U46251 (N_46251,N_46058,N_46099);
and U46252 (N_46252,N_46047,N_46034);
and U46253 (N_46253,N_46091,N_46109);
and U46254 (N_46254,N_46180,N_46079);
nand U46255 (N_46255,N_46096,N_46204);
or U46256 (N_46256,N_46106,N_46012);
nand U46257 (N_46257,N_46187,N_46158);
xnor U46258 (N_46258,N_46219,N_46145);
and U46259 (N_46259,N_46082,N_46006);
nand U46260 (N_46260,N_46013,N_46238);
xnor U46261 (N_46261,N_46067,N_46179);
or U46262 (N_46262,N_46051,N_46198);
or U46263 (N_46263,N_46146,N_46170);
or U46264 (N_46264,N_46149,N_46025);
or U46265 (N_46265,N_46244,N_46026);
nor U46266 (N_46266,N_46153,N_46188);
nor U46267 (N_46267,N_46197,N_46032);
and U46268 (N_46268,N_46165,N_46137);
or U46269 (N_46269,N_46039,N_46027);
and U46270 (N_46270,N_46246,N_46084);
nor U46271 (N_46271,N_46065,N_46053);
xor U46272 (N_46272,N_46175,N_46222);
xnor U46273 (N_46273,N_46019,N_46060);
or U46274 (N_46274,N_46057,N_46075);
xor U46275 (N_46275,N_46016,N_46064);
nor U46276 (N_46276,N_46154,N_46235);
xor U46277 (N_46277,N_46209,N_46201);
or U46278 (N_46278,N_46152,N_46218);
nand U46279 (N_46279,N_46052,N_46108);
and U46280 (N_46280,N_46178,N_46011);
or U46281 (N_46281,N_46144,N_46159);
nor U46282 (N_46282,N_46226,N_46206);
and U46283 (N_46283,N_46123,N_46169);
or U46284 (N_46284,N_46164,N_46014);
or U46285 (N_46285,N_46220,N_46161);
nand U46286 (N_46286,N_46128,N_46105);
or U46287 (N_46287,N_46098,N_46166);
xnor U46288 (N_46288,N_46202,N_46157);
nor U46289 (N_46289,N_46054,N_46031);
xor U46290 (N_46290,N_46184,N_46074);
xnor U46291 (N_46291,N_46231,N_46239);
nor U46292 (N_46292,N_46055,N_46121);
xnor U46293 (N_46293,N_46083,N_46010);
xnor U46294 (N_46294,N_46037,N_46035);
nor U46295 (N_46295,N_46212,N_46076);
xor U46296 (N_46296,N_46115,N_46237);
nand U46297 (N_46297,N_46195,N_46189);
and U46298 (N_46298,N_46173,N_46190);
or U46299 (N_46299,N_46101,N_46140);
nand U46300 (N_46300,N_46062,N_46208);
xor U46301 (N_46301,N_46038,N_46048);
nor U46302 (N_46302,N_46131,N_46107);
or U46303 (N_46303,N_46040,N_46232);
xnor U46304 (N_46304,N_46160,N_46205);
nor U46305 (N_46305,N_46071,N_46225);
nor U46306 (N_46306,N_46207,N_46147);
nor U46307 (N_46307,N_46245,N_46095);
xor U46308 (N_46308,N_46033,N_46183);
nand U46309 (N_46309,N_46059,N_46122);
nand U46310 (N_46310,N_46030,N_46217);
and U46311 (N_46311,N_46024,N_46249);
nor U46312 (N_46312,N_46193,N_46148);
nor U46313 (N_46313,N_46174,N_46117);
nand U46314 (N_46314,N_46092,N_46139);
nor U46315 (N_46315,N_46070,N_46168);
nand U46316 (N_46316,N_46241,N_46029);
xor U46317 (N_46317,N_46068,N_46133);
and U46318 (N_46318,N_46097,N_46242);
nor U46319 (N_46319,N_46126,N_46236);
xnor U46320 (N_46320,N_46104,N_46088);
or U46321 (N_46321,N_46136,N_46112);
nor U46322 (N_46322,N_46182,N_46233);
nand U46323 (N_46323,N_46247,N_46211);
and U46324 (N_46324,N_46000,N_46078);
nor U46325 (N_46325,N_46045,N_46020);
nor U46326 (N_46326,N_46110,N_46192);
or U46327 (N_46327,N_46111,N_46094);
or U46328 (N_46328,N_46087,N_46171);
and U46329 (N_46329,N_46234,N_46142);
and U46330 (N_46330,N_46005,N_46213);
xnor U46331 (N_46331,N_46073,N_46118);
nand U46332 (N_46332,N_46085,N_46243);
nor U46333 (N_46333,N_46196,N_46056);
or U46334 (N_46334,N_46018,N_46028);
or U46335 (N_46335,N_46090,N_46176);
nor U46336 (N_46336,N_46066,N_46200);
nor U46337 (N_46337,N_46061,N_46041);
and U46338 (N_46338,N_46130,N_46021);
and U46339 (N_46339,N_46214,N_46156);
or U46340 (N_46340,N_46002,N_46086);
nand U46341 (N_46341,N_46199,N_46080);
or U46342 (N_46342,N_46017,N_46143);
nor U46343 (N_46343,N_46210,N_46001);
nor U46344 (N_46344,N_46223,N_46151);
and U46345 (N_46345,N_46129,N_46043);
or U46346 (N_46346,N_46177,N_46022);
nand U46347 (N_46347,N_46203,N_46186);
or U46348 (N_46348,N_46069,N_46063);
nand U46349 (N_46349,N_46008,N_46102);
or U46350 (N_46350,N_46221,N_46194);
nor U46351 (N_46351,N_46113,N_46089);
or U46352 (N_46352,N_46120,N_46050);
xor U46353 (N_46353,N_46150,N_46103);
and U46354 (N_46354,N_46004,N_46228);
and U46355 (N_46355,N_46191,N_46135);
and U46356 (N_46356,N_46042,N_46124);
xnor U46357 (N_46357,N_46185,N_46007);
xor U46358 (N_46358,N_46155,N_46023);
and U46359 (N_46359,N_46119,N_46081);
nor U46360 (N_46360,N_46163,N_46132);
or U46361 (N_46361,N_46162,N_46172);
or U46362 (N_46362,N_46036,N_46114);
or U46363 (N_46363,N_46072,N_46044);
xor U46364 (N_46364,N_46230,N_46093);
nand U46365 (N_46365,N_46100,N_46240);
xnor U46366 (N_46366,N_46248,N_46224);
and U46367 (N_46367,N_46134,N_46167);
nor U46368 (N_46368,N_46216,N_46181);
nor U46369 (N_46369,N_46077,N_46127);
nor U46370 (N_46370,N_46049,N_46015);
nand U46371 (N_46371,N_46138,N_46116);
nand U46372 (N_46372,N_46229,N_46009);
nor U46373 (N_46373,N_46141,N_46227);
nand U46374 (N_46374,N_46215,N_46046);
and U46375 (N_46375,N_46027,N_46191);
or U46376 (N_46376,N_46137,N_46147);
and U46377 (N_46377,N_46238,N_46234);
nand U46378 (N_46378,N_46115,N_46114);
xnor U46379 (N_46379,N_46087,N_46034);
nor U46380 (N_46380,N_46170,N_46072);
and U46381 (N_46381,N_46086,N_46022);
or U46382 (N_46382,N_46166,N_46144);
nand U46383 (N_46383,N_46232,N_46141);
nand U46384 (N_46384,N_46216,N_46127);
nor U46385 (N_46385,N_46175,N_46124);
or U46386 (N_46386,N_46188,N_46109);
nand U46387 (N_46387,N_46046,N_46023);
or U46388 (N_46388,N_46126,N_46203);
nand U46389 (N_46389,N_46157,N_46190);
xnor U46390 (N_46390,N_46158,N_46116);
xnor U46391 (N_46391,N_46100,N_46027);
xnor U46392 (N_46392,N_46203,N_46223);
nor U46393 (N_46393,N_46221,N_46170);
and U46394 (N_46394,N_46079,N_46231);
or U46395 (N_46395,N_46086,N_46013);
or U46396 (N_46396,N_46210,N_46083);
xor U46397 (N_46397,N_46122,N_46140);
and U46398 (N_46398,N_46131,N_46111);
xor U46399 (N_46399,N_46091,N_46064);
nor U46400 (N_46400,N_46151,N_46139);
xnor U46401 (N_46401,N_46222,N_46019);
xnor U46402 (N_46402,N_46035,N_46136);
xor U46403 (N_46403,N_46215,N_46006);
nand U46404 (N_46404,N_46006,N_46172);
or U46405 (N_46405,N_46140,N_46010);
xor U46406 (N_46406,N_46159,N_46083);
xnor U46407 (N_46407,N_46077,N_46006);
xnor U46408 (N_46408,N_46046,N_46161);
or U46409 (N_46409,N_46231,N_46156);
nand U46410 (N_46410,N_46232,N_46004);
xnor U46411 (N_46411,N_46059,N_46222);
and U46412 (N_46412,N_46248,N_46097);
xor U46413 (N_46413,N_46099,N_46163);
and U46414 (N_46414,N_46073,N_46180);
nor U46415 (N_46415,N_46236,N_46160);
nor U46416 (N_46416,N_46035,N_46176);
nor U46417 (N_46417,N_46002,N_46037);
and U46418 (N_46418,N_46085,N_46151);
xnor U46419 (N_46419,N_46043,N_46164);
nand U46420 (N_46420,N_46152,N_46157);
or U46421 (N_46421,N_46040,N_46090);
and U46422 (N_46422,N_46189,N_46114);
and U46423 (N_46423,N_46215,N_46093);
or U46424 (N_46424,N_46108,N_46147);
nor U46425 (N_46425,N_46197,N_46071);
nor U46426 (N_46426,N_46123,N_46104);
or U46427 (N_46427,N_46096,N_46070);
or U46428 (N_46428,N_46189,N_46109);
nor U46429 (N_46429,N_46060,N_46204);
or U46430 (N_46430,N_46164,N_46190);
xor U46431 (N_46431,N_46181,N_46211);
and U46432 (N_46432,N_46094,N_46055);
and U46433 (N_46433,N_46234,N_46020);
nor U46434 (N_46434,N_46195,N_46109);
xor U46435 (N_46435,N_46177,N_46067);
and U46436 (N_46436,N_46000,N_46141);
nand U46437 (N_46437,N_46140,N_46192);
nor U46438 (N_46438,N_46080,N_46017);
xnor U46439 (N_46439,N_46083,N_46061);
nand U46440 (N_46440,N_46190,N_46147);
and U46441 (N_46441,N_46076,N_46203);
nor U46442 (N_46442,N_46171,N_46240);
and U46443 (N_46443,N_46019,N_46164);
and U46444 (N_46444,N_46135,N_46072);
nor U46445 (N_46445,N_46031,N_46070);
nand U46446 (N_46446,N_46132,N_46155);
nor U46447 (N_46447,N_46175,N_46024);
nand U46448 (N_46448,N_46120,N_46055);
and U46449 (N_46449,N_46225,N_46186);
nor U46450 (N_46450,N_46065,N_46074);
and U46451 (N_46451,N_46184,N_46124);
nand U46452 (N_46452,N_46146,N_46208);
and U46453 (N_46453,N_46217,N_46155);
nand U46454 (N_46454,N_46167,N_46157);
or U46455 (N_46455,N_46065,N_46222);
and U46456 (N_46456,N_46198,N_46144);
xor U46457 (N_46457,N_46192,N_46241);
or U46458 (N_46458,N_46013,N_46100);
xnor U46459 (N_46459,N_46228,N_46173);
xor U46460 (N_46460,N_46237,N_46137);
and U46461 (N_46461,N_46137,N_46140);
xnor U46462 (N_46462,N_46024,N_46206);
and U46463 (N_46463,N_46090,N_46196);
nand U46464 (N_46464,N_46076,N_46030);
nand U46465 (N_46465,N_46142,N_46097);
or U46466 (N_46466,N_46142,N_46197);
and U46467 (N_46467,N_46104,N_46057);
nor U46468 (N_46468,N_46115,N_46131);
or U46469 (N_46469,N_46202,N_46197);
nand U46470 (N_46470,N_46008,N_46177);
and U46471 (N_46471,N_46095,N_46203);
and U46472 (N_46472,N_46024,N_46073);
or U46473 (N_46473,N_46160,N_46116);
xnor U46474 (N_46474,N_46128,N_46196);
nand U46475 (N_46475,N_46155,N_46048);
and U46476 (N_46476,N_46064,N_46018);
or U46477 (N_46477,N_46000,N_46179);
or U46478 (N_46478,N_46185,N_46122);
nand U46479 (N_46479,N_46059,N_46153);
xor U46480 (N_46480,N_46038,N_46094);
nand U46481 (N_46481,N_46014,N_46032);
nand U46482 (N_46482,N_46108,N_46059);
xor U46483 (N_46483,N_46225,N_46027);
nand U46484 (N_46484,N_46078,N_46082);
xor U46485 (N_46485,N_46232,N_46056);
xor U46486 (N_46486,N_46021,N_46209);
and U46487 (N_46487,N_46209,N_46230);
nor U46488 (N_46488,N_46024,N_46052);
xnor U46489 (N_46489,N_46077,N_46064);
nand U46490 (N_46490,N_46199,N_46235);
or U46491 (N_46491,N_46218,N_46249);
and U46492 (N_46492,N_46219,N_46185);
nor U46493 (N_46493,N_46157,N_46045);
nor U46494 (N_46494,N_46150,N_46102);
xnor U46495 (N_46495,N_46160,N_46083);
nor U46496 (N_46496,N_46058,N_46121);
and U46497 (N_46497,N_46156,N_46094);
xor U46498 (N_46498,N_46163,N_46184);
and U46499 (N_46499,N_46055,N_46177);
nand U46500 (N_46500,N_46382,N_46435);
nand U46501 (N_46501,N_46263,N_46306);
nor U46502 (N_46502,N_46292,N_46334);
or U46503 (N_46503,N_46408,N_46467);
xnor U46504 (N_46504,N_46270,N_46446);
and U46505 (N_46505,N_46320,N_46426);
and U46506 (N_46506,N_46287,N_46478);
nor U46507 (N_46507,N_46498,N_46286);
nand U46508 (N_46508,N_46305,N_46416);
xor U46509 (N_46509,N_46399,N_46445);
xnor U46510 (N_46510,N_46473,N_46359);
or U46511 (N_46511,N_46256,N_46415);
xnor U46512 (N_46512,N_46474,N_46462);
xnor U46513 (N_46513,N_46282,N_46295);
and U46514 (N_46514,N_46331,N_46255);
and U46515 (N_46515,N_46332,N_46311);
nor U46516 (N_46516,N_46251,N_46326);
nor U46517 (N_46517,N_46465,N_46372);
nor U46518 (N_46518,N_46375,N_46436);
xnor U46519 (N_46519,N_46314,N_46280);
nand U46520 (N_46520,N_46466,N_46487);
and U46521 (N_46521,N_46387,N_46452);
and U46522 (N_46522,N_46335,N_46421);
nor U46523 (N_46523,N_46479,N_46464);
or U46524 (N_46524,N_46425,N_46343);
or U46525 (N_46525,N_46342,N_46357);
nand U46526 (N_46526,N_46302,N_46406);
or U46527 (N_46527,N_46353,N_46482);
or U46528 (N_46528,N_46497,N_46404);
nor U46529 (N_46529,N_46461,N_46451);
or U46530 (N_46530,N_46312,N_46304);
xor U46531 (N_46531,N_46259,N_46475);
nand U46532 (N_46532,N_46308,N_46257);
nand U46533 (N_46533,N_46325,N_46460);
nor U46534 (N_46534,N_46279,N_46266);
xor U46535 (N_46535,N_46362,N_46373);
and U46536 (N_46536,N_46333,N_46419);
or U46537 (N_46537,N_46293,N_46267);
and U46538 (N_46538,N_46337,N_46485);
xnor U46539 (N_46539,N_46448,N_46420);
and U46540 (N_46540,N_46299,N_46455);
nor U46541 (N_46541,N_46265,N_46427);
nand U46542 (N_46542,N_46431,N_46341);
nand U46543 (N_46543,N_46361,N_46392);
nor U46544 (N_46544,N_46469,N_46271);
nand U46545 (N_46545,N_46397,N_46386);
nor U46546 (N_46546,N_46401,N_46405);
or U46547 (N_46547,N_46403,N_46338);
or U46548 (N_46548,N_46402,N_46481);
nor U46549 (N_46549,N_46422,N_46388);
and U46550 (N_46550,N_46294,N_46400);
or U46551 (N_46551,N_46443,N_46396);
nand U46552 (N_46552,N_46423,N_46364);
nand U46553 (N_46553,N_46490,N_46300);
and U46554 (N_46554,N_46317,N_46477);
nor U46555 (N_46555,N_46269,N_46289);
or U46556 (N_46556,N_46472,N_46275);
and U46557 (N_46557,N_46354,N_46432);
xor U46558 (N_46558,N_46358,N_46458);
or U46559 (N_46559,N_46492,N_46494);
or U46560 (N_46560,N_46339,N_46297);
and U46561 (N_46561,N_46319,N_46355);
xnor U46562 (N_46562,N_46336,N_46395);
xor U46563 (N_46563,N_46322,N_46369);
and U46564 (N_46564,N_46367,N_46380);
nand U46565 (N_46565,N_46301,N_46457);
nand U46566 (N_46566,N_46250,N_46488);
and U46567 (N_46567,N_46454,N_46347);
and U46568 (N_46568,N_46389,N_46328);
and U46569 (N_46569,N_46428,N_46360);
xnor U46570 (N_46570,N_46385,N_46323);
or U46571 (N_46571,N_46418,N_46459);
or U46572 (N_46572,N_46258,N_46316);
xor U46573 (N_46573,N_46313,N_46484);
xnor U46574 (N_46574,N_46398,N_46495);
nand U46575 (N_46575,N_46350,N_46268);
nor U46576 (N_46576,N_46278,N_46381);
or U46577 (N_46577,N_46288,N_46315);
or U46578 (N_46578,N_46424,N_46284);
xor U46579 (N_46579,N_46499,N_46496);
xnor U46580 (N_46580,N_46410,N_46480);
xnor U46581 (N_46581,N_46453,N_46470);
xor U46582 (N_46582,N_46281,N_46413);
and U46583 (N_46583,N_46414,N_46383);
xnor U46584 (N_46584,N_46371,N_46430);
or U46585 (N_46585,N_46352,N_46447);
or U46586 (N_46586,N_46272,N_46391);
nand U46587 (N_46587,N_46262,N_46351);
nand U46588 (N_46588,N_46348,N_46449);
or U46589 (N_46589,N_46476,N_46264);
nand U46590 (N_46590,N_46254,N_46285);
xor U46591 (N_46591,N_46491,N_46273);
and U46592 (N_46592,N_46298,N_46307);
and U46593 (N_46593,N_46433,N_46349);
xnor U46594 (N_46594,N_46411,N_46370);
and U46595 (N_46595,N_46393,N_46468);
nor U46596 (N_46596,N_46471,N_46440);
or U46597 (N_46597,N_46296,N_46377);
nor U46598 (N_46598,N_46442,N_46276);
and U46599 (N_46599,N_46363,N_46378);
nand U46600 (N_46600,N_46309,N_46439);
nor U46601 (N_46601,N_46329,N_46346);
and U46602 (N_46602,N_46409,N_46429);
or U46603 (N_46603,N_46321,N_46366);
or U46604 (N_46604,N_46253,N_46327);
and U46605 (N_46605,N_46390,N_46394);
and U46606 (N_46606,N_46345,N_46260);
nor U46607 (N_46607,N_46291,N_46456);
xnor U46608 (N_46608,N_46252,N_46310);
and U46609 (N_46609,N_46261,N_46463);
xnor U46610 (N_46610,N_46486,N_46303);
and U46611 (N_46611,N_46444,N_46379);
and U46612 (N_46612,N_46344,N_46434);
xor U46613 (N_46613,N_46438,N_46365);
xor U46614 (N_46614,N_46483,N_46324);
nand U46615 (N_46615,N_46318,N_46384);
xnor U46616 (N_46616,N_46356,N_46417);
nor U46617 (N_46617,N_46412,N_46450);
and U46618 (N_46618,N_46283,N_46290);
and U46619 (N_46619,N_46441,N_46407);
xnor U46620 (N_46620,N_46274,N_46493);
and U46621 (N_46621,N_46340,N_46489);
nand U46622 (N_46622,N_46437,N_46368);
nor U46623 (N_46623,N_46374,N_46376);
or U46624 (N_46624,N_46330,N_46277);
and U46625 (N_46625,N_46464,N_46295);
xnor U46626 (N_46626,N_46325,N_46499);
xnor U46627 (N_46627,N_46315,N_46465);
xnor U46628 (N_46628,N_46446,N_46378);
nor U46629 (N_46629,N_46304,N_46306);
or U46630 (N_46630,N_46307,N_46284);
and U46631 (N_46631,N_46313,N_46443);
or U46632 (N_46632,N_46309,N_46483);
or U46633 (N_46633,N_46324,N_46465);
nand U46634 (N_46634,N_46372,N_46421);
and U46635 (N_46635,N_46380,N_46432);
nand U46636 (N_46636,N_46293,N_46478);
or U46637 (N_46637,N_46427,N_46354);
nor U46638 (N_46638,N_46381,N_46372);
nor U46639 (N_46639,N_46319,N_46452);
nand U46640 (N_46640,N_46437,N_46289);
nand U46641 (N_46641,N_46290,N_46435);
xnor U46642 (N_46642,N_46436,N_46316);
nand U46643 (N_46643,N_46498,N_46434);
nand U46644 (N_46644,N_46442,N_46297);
nand U46645 (N_46645,N_46450,N_46435);
and U46646 (N_46646,N_46484,N_46418);
nand U46647 (N_46647,N_46427,N_46426);
or U46648 (N_46648,N_46459,N_46431);
nor U46649 (N_46649,N_46440,N_46261);
xor U46650 (N_46650,N_46337,N_46260);
nand U46651 (N_46651,N_46492,N_46366);
nand U46652 (N_46652,N_46263,N_46454);
xor U46653 (N_46653,N_46269,N_46287);
nand U46654 (N_46654,N_46361,N_46412);
nor U46655 (N_46655,N_46347,N_46461);
xor U46656 (N_46656,N_46341,N_46260);
or U46657 (N_46657,N_46390,N_46359);
nor U46658 (N_46658,N_46459,N_46466);
or U46659 (N_46659,N_46290,N_46370);
and U46660 (N_46660,N_46445,N_46382);
and U46661 (N_46661,N_46416,N_46379);
or U46662 (N_46662,N_46272,N_46466);
xnor U46663 (N_46663,N_46293,N_46445);
nor U46664 (N_46664,N_46300,N_46458);
or U46665 (N_46665,N_46357,N_46462);
nor U46666 (N_46666,N_46484,N_46417);
nor U46667 (N_46667,N_46347,N_46308);
or U46668 (N_46668,N_46452,N_46475);
xnor U46669 (N_46669,N_46430,N_46414);
xnor U46670 (N_46670,N_46431,N_46416);
and U46671 (N_46671,N_46497,N_46336);
nand U46672 (N_46672,N_46328,N_46345);
xnor U46673 (N_46673,N_46443,N_46476);
nand U46674 (N_46674,N_46270,N_46476);
xnor U46675 (N_46675,N_46386,N_46285);
or U46676 (N_46676,N_46449,N_46440);
nor U46677 (N_46677,N_46406,N_46359);
or U46678 (N_46678,N_46392,N_46358);
xor U46679 (N_46679,N_46362,N_46273);
and U46680 (N_46680,N_46441,N_46348);
nand U46681 (N_46681,N_46290,N_46295);
or U46682 (N_46682,N_46412,N_46370);
and U46683 (N_46683,N_46350,N_46434);
nor U46684 (N_46684,N_46285,N_46321);
nand U46685 (N_46685,N_46363,N_46272);
or U46686 (N_46686,N_46492,N_46441);
nor U46687 (N_46687,N_46427,N_46322);
xor U46688 (N_46688,N_46258,N_46385);
xnor U46689 (N_46689,N_46335,N_46255);
xnor U46690 (N_46690,N_46260,N_46373);
and U46691 (N_46691,N_46281,N_46416);
or U46692 (N_46692,N_46265,N_46440);
or U46693 (N_46693,N_46316,N_46290);
or U46694 (N_46694,N_46275,N_46446);
or U46695 (N_46695,N_46275,N_46257);
nand U46696 (N_46696,N_46493,N_46319);
xor U46697 (N_46697,N_46289,N_46305);
and U46698 (N_46698,N_46469,N_46454);
nor U46699 (N_46699,N_46416,N_46327);
nand U46700 (N_46700,N_46392,N_46300);
nor U46701 (N_46701,N_46337,N_46358);
or U46702 (N_46702,N_46415,N_46476);
xnor U46703 (N_46703,N_46322,N_46324);
or U46704 (N_46704,N_46356,N_46354);
or U46705 (N_46705,N_46362,N_46305);
or U46706 (N_46706,N_46441,N_46364);
and U46707 (N_46707,N_46439,N_46430);
xor U46708 (N_46708,N_46436,N_46408);
and U46709 (N_46709,N_46488,N_46256);
nand U46710 (N_46710,N_46429,N_46384);
or U46711 (N_46711,N_46461,N_46445);
xor U46712 (N_46712,N_46332,N_46416);
nor U46713 (N_46713,N_46491,N_46391);
or U46714 (N_46714,N_46316,N_46477);
nand U46715 (N_46715,N_46259,N_46379);
nor U46716 (N_46716,N_46391,N_46409);
and U46717 (N_46717,N_46392,N_46471);
and U46718 (N_46718,N_46495,N_46263);
and U46719 (N_46719,N_46384,N_46462);
nor U46720 (N_46720,N_46294,N_46367);
nor U46721 (N_46721,N_46421,N_46389);
or U46722 (N_46722,N_46461,N_46428);
or U46723 (N_46723,N_46395,N_46425);
or U46724 (N_46724,N_46371,N_46455);
and U46725 (N_46725,N_46368,N_46254);
xor U46726 (N_46726,N_46291,N_46447);
nand U46727 (N_46727,N_46267,N_46271);
xnor U46728 (N_46728,N_46462,N_46377);
or U46729 (N_46729,N_46275,N_46377);
and U46730 (N_46730,N_46269,N_46355);
or U46731 (N_46731,N_46258,N_46419);
xnor U46732 (N_46732,N_46283,N_46480);
xor U46733 (N_46733,N_46343,N_46486);
and U46734 (N_46734,N_46451,N_46370);
nor U46735 (N_46735,N_46493,N_46466);
nor U46736 (N_46736,N_46437,N_46369);
xnor U46737 (N_46737,N_46392,N_46298);
xor U46738 (N_46738,N_46484,N_46360);
nor U46739 (N_46739,N_46279,N_46335);
or U46740 (N_46740,N_46306,N_46255);
nor U46741 (N_46741,N_46295,N_46473);
or U46742 (N_46742,N_46393,N_46482);
nand U46743 (N_46743,N_46489,N_46498);
xnor U46744 (N_46744,N_46467,N_46363);
nor U46745 (N_46745,N_46316,N_46472);
or U46746 (N_46746,N_46362,N_46459);
nor U46747 (N_46747,N_46433,N_46364);
or U46748 (N_46748,N_46432,N_46388);
nand U46749 (N_46749,N_46258,N_46453);
xor U46750 (N_46750,N_46517,N_46688);
or U46751 (N_46751,N_46630,N_46588);
and U46752 (N_46752,N_46509,N_46691);
xor U46753 (N_46753,N_46711,N_46582);
xor U46754 (N_46754,N_46535,N_46689);
and U46755 (N_46755,N_46645,N_46680);
nand U46756 (N_46756,N_46728,N_46508);
and U46757 (N_46757,N_46725,N_46609);
and U46758 (N_46758,N_46667,N_46592);
or U46759 (N_46759,N_46548,N_46614);
nor U46760 (N_46760,N_46610,N_46607);
xor U46761 (N_46761,N_46671,N_46542);
xnor U46762 (N_46762,N_46662,N_46655);
or U46763 (N_46763,N_46749,N_46574);
nor U46764 (N_46764,N_46576,N_46572);
nand U46765 (N_46765,N_46549,N_46726);
xnor U46766 (N_46766,N_46723,N_46637);
nand U46767 (N_46767,N_46577,N_46503);
and U46768 (N_46768,N_46650,N_46589);
and U46769 (N_46769,N_46740,N_46743);
xnor U46770 (N_46770,N_46521,N_46516);
nand U46771 (N_46771,N_46598,N_46616);
nand U46772 (N_46772,N_46674,N_46647);
nor U46773 (N_46773,N_46565,N_46586);
nand U46774 (N_46774,N_46611,N_46651);
or U46775 (N_46775,N_46530,N_46604);
nand U46776 (N_46776,N_46600,N_46608);
or U46777 (N_46777,N_46682,N_46605);
xnor U46778 (N_46778,N_46700,N_46533);
nand U46779 (N_46779,N_46656,N_46677);
nor U46780 (N_46780,N_46665,N_46709);
or U46781 (N_46781,N_46559,N_46522);
nand U46782 (N_46782,N_46715,N_46705);
or U46783 (N_46783,N_46507,N_46718);
nand U46784 (N_46784,N_46623,N_46684);
xor U46785 (N_46785,N_46524,N_46694);
or U46786 (N_46786,N_46707,N_46699);
nand U46787 (N_46787,N_46644,N_46638);
xnor U46788 (N_46788,N_46527,N_46532);
or U46789 (N_46789,N_46547,N_46511);
or U46790 (N_46790,N_46729,N_46666);
or U46791 (N_46791,N_46717,N_46681);
and U46792 (N_46792,N_46561,N_46693);
and U46793 (N_46793,N_46580,N_46599);
xnor U46794 (N_46794,N_46748,N_46668);
and U46795 (N_46795,N_46612,N_46613);
or U46796 (N_46796,N_46735,N_46575);
and U46797 (N_46797,N_46556,N_46624);
nand U46798 (N_46798,N_46730,N_46736);
nand U46799 (N_46799,N_46738,N_46500);
or U46800 (N_46800,N_46529,N_46675);
nor U46801 (N_46801,N_46539,N_46625);
and U46802 (N_46802,N_46722,N_46706);
or U46803 (N_46803,N_46573,N_46652);
xor U46804 (N_46804,N_46659,N_46552);
nor U46805 (N_46805,N_46628,N_46578);
or U46806 (N_46806,N_46678,N_46557);
nor U46807 (N_46807,N_46657,N_46708);
or U46808 (N_46808,N_46569,N_46518);
xnor U46809 (N_46809,N_46734,N_46620);
and U46810 (N_46810,N_46741,N_46502);
xor U46811 (N_46811,N_46713,N_46515);
and U46812 (N_46812,N_46660,N_46550);
nand U46813 (N_46813,N_46727,N_46663);
and U46814 (N_46814,N_46519,N_46544);
nor U46815 (N_46815,N_46510,N_46721);
and U46816 (N_46816,N_46563,N_46568);
nand U46817 (N_46817,N_46546,N_46595);
xnor U46818 (N_46818,N_46746,N_46564);
nor U46819 (N_46819,N_46602,N_46692);
nor U46820 (N_46820,N_46744,N_46618);
nor U46821 (N_46821,N_46731,N_46698);
nor U46822 (N_46822,N_46562,N_46596);
or U46823 (N_46823,N_46583,N_46683);
and U46824 (N_46824,N_46570,N_46501);
or U46825 (N_46825,N_46732,N_46640);
nor U46826 (N_46826,N_46551,N_46635);
or U46827 (N_46827,N_46634,N_46737);
nand U46828 (N_46828,N_46629,N_46615);
xor U46829 (N_46829,N_46538,N_46622);
nand U46830 (N_46830,N_46672,N_46512);
xnor U46831 (N_46831,N_46742,N_46702);
or U46832 (N_46832,N_46653,N_46545);
xor U46833 (N_46833,N_46639,N_46733);
nor U46834 (N_46834,N_46701,N_46579);
xor U46835 (N_46835,N_46581,N_46641);
nor U46836 (N_46836,N_46513,N_46673);
nand U46837 (N_46837,N_46591,N_46670);
xnor U46838 (N_46838,N_46584,N_46719);
and U46839 (N_46839,N_46686,N_46543);
xor U46840 (N_46840,N_46528,N_46523);
and U46841 (N_46841,N_46745,N_46601);
and U46842 (N_46842,N_46654,N_46714);
xor U46843 (N_46843,N_46606,N_46695);
or U46844 (N_46844,N_46593,N_46724);
nor U46845 (N_46845,N_46633,N_46587);
and U46846 (N_46846,N_46649,N_46590);
and U46847 (N_46847,N_46558,N_46676);
xor U46848 (N_46848,N_46526,N_46631);
nand U46849 (N_46849,N_46747,N_46627);
and U46850 (N_46850,N_46617,N_46636);
nand U46851 (N_46851,N_46531,N_46553);
or U46852 (N_46852,N_46504,N_46703);
xor U46853 (N_46853,N_46585,N_46594);
nor U46854 (N_46854,N_46554,N_46739);
xor U46855 (N_46855,N_46669,N_46537);
xor U46856 (N_46856,N_46603,N_46525);
and U46857 (N_46857,N_46712,N_46710);
nand U46858 (N_46858,N_46555,N_46534);
and U46859 (N_46859,N_46505,N_46520);
nor U46860 (N_46860,N_46541,N_46696);
xor U46861 (N_46861,N_46716,N_46679);
nand U46862 (N_46862,N_46632,N_46697);
xor U46863 (N_46863,N_46720,N_46540);
nor U46864 (N_46864,N_46661,N_46536);
nor U46865 (N_46865,N_46626,N_46643);
xnor U46866 (N_46866,N_46664,N_46704);
or U46867 (N_46867,N_46690,N_46567);
nand U46868 (N_46868,N_46658,N_46648);
and U46869 (N_46869,N_46646,N_46619);
xor U46870 (N_46870,N_46687,N_46560);
nand U46871 (N_46871,N_46571,N_46685);
xor U46872 (N_46872,N_46514,N_46621);
and U46873 (N_46873,N_46566,N_46506);
nor U46874 (N_46874,N_46642,N_46597);
and U46875 (N_46875,N_46713,N_46629);
nor U46876 (N_46876,N_46706,N_46549);
nor U46877 (N_46877,N_46589,N_46694);
nand U46878 (N_46878,N_46699,N_46727);
and U46879 (N_46879,N_46524,N_46736);
or U46880 (N_46880,N_46632,N_46600);
nor U46881 (N_46881,N_46663,N_46650);
or U46882 (N_46882,N_46574,N_46652);
nand U46883 (N_46883,N_46555,N_46732);
or U46884 (N_46884,N_46628,N_46654);
nand U46885 (N_46885,N_46553,N_46608);
and U46886 (N_46886,N_46630,N_46695);
nor U46887 (N_46887,N_46563,N_46547);
nor U46888 (N_46888,N_46685,N_46728);
or U46889 (N_46889,N_46702,N_46501);
nand U46890 (N_46890,N_46685,N_46500);
or U46891 (N_46891,N_46583,N_46634);
and U46892 (N_46892,N_46654,N_46691);
and U46893 (N_46893,N_46714,N_46628);
nor U46894 (N_46894,N_46644,N_46562);
nor U46895 (N_46895,N_46520,N_46581);
nor U46896 (N_46896,N_46722,N_46553);
nor U46897 (N_46897,N_46559,N_46675);
xor U46898 (N_46898,N_46587,N_46500);
and U46899 (N_46899,N_46536,N_46694);
xnor U46900 (N_46900,N_46545,N_46673);
xor U46901 (N_46901,N_46510,N_46730);
and U46902 (N_46902,N_46661,N_46649);
and U46903 (N_46903,N_46731,N_46558);
nor U46904 (N_46904,N_46589,N_46676);
nand U46905 (N_46905,N_46578,N_46709);
xnor U46906 (N_46906,N_46749,N_46729);
and U46907 (N_46907,N_46627,N_46665);
or U46908 (N_46908,N_46645,N_46525);
nor U46909 (N_46909,N_46576,N_46558);
and U46910 (N_46910,N_46664,N_46624);
and U46911 (N_46911,N_46589,N_46641);
or U46912 (N_46912,N_46625,N_46502);
nor U46913 (N_46913,N_46687,N_46627);
and U46914 (N_46914,N_46536,N_46599);
nor U46915 (N_46915,N_46700,N_46536);
or U46916 (N_46916,N_46501,N_46689);
xor U46917 (N_46917,N_46665,N_46706);
and U46918 (N_46918,N_46545,N_46626);
or U46919 (N_46919,N_46612,N_46537);
xnor U46920 (N_46920,N_46668,N_46640);
nor U46921 (N_46921,N_46702,N_46591);
or U46922 (N_46922,N_46617,N_46644);
xor U46923 (N_46923,N_46585,N_46693);
or U46924 (N_46924,N_46514,N_46664);
xor U46925 (N_46925,N_46608,N_46748);
or U46926 (N_46926,N_46656,N_46653);
and U46927 (N_46927,N_46548,N_46592);
nor U46928 (N_46928,N_46735,N_46729);
and U46929 (N_46929,N_46632,N_46574);
nor U46930 (N_46930,N_46665,N_46537);
nor U46931 (N_46931,N_46536,N_46545);
or U46932 (N_46932,N_46608,N_46508);
xnor U46933 (N_46933,N_46729,N_46554);
nor U46934 (N_46934,N_46726,N_46525);
nand U46935 (N_46935,N_46693,N_46628);
xnor U46936 (N_46936,N_46644,N_46553);
and U46937 (N_46937,N_46556,N_46676);
or U46938 (N_46938,N_46668,N_46593);
xor U46939 (N_46939,N_46592,N_46587);
nand U46940 (N_46940,N_46590,N_46589);
and U46941 (N_46941,N_46640,N_46538);
xnor U46942 (N_46942,N_46692,N_46635);
xor U46943 (N_46943,N_46698,N_46679);
nand U46944 (N_46944,N_46593,N_46744);
nor U46945 (N_46945,N_46518,N_46523);
nand U46946 (N_46946,N_46547,N_46569);
xnor U46947 (N_46947,N_46516,N_46631);
nor U46948 (N_46948,N_46635,N_46633);
xnor U46949 (N_46949,N_46533,N_46616);
and U46950 (N_46950,N_46610,N_46735);
or U46951 (N_46951,N_46703,N_46645);
or U46952 (N_46952,N_46632,N_46740);
and U46953 (N_46953,N_46588,N_46565);
nand U46954 (N_46954,N_46666,N_46697);
nand U46955 (N_46955,N_46606,N_46568);
nor U46956 (N_46956,N_46614,N_46615);
nand U46957 (N_46957,N_46737,N_46530);
xnor U46958 (N_46958,N_46664,N_46694);
nor U46959 (N_46959,N_46659,N_46686);
and U46960 (N_46960,N_46573,N_46638);
and U46961 (N_46961,N_46623,N_46598);
nor U46962 (N_46962,N_46518,N_46629);
nand U46963 (N_46963,N_46704,N_46722);
nand U46964 (N_46964,N_46667,N_46504);
and U46965 (N_46965,N_46551,N_46704);
nor U46966 (N_46966,N_46664,N_46553);
nor U46967 (N_46967,N_46664,N_46536);
and U46968 (N_46968,N_46694,N_46648);
and U46969 (N_46969,N_46651,N_46647);
xnor U46970 (N_46970,N_46648,N_46721);
and U46971 (N_46971,N_46699,N_46504);
and U46972 (N_46972,N_46639,N_46633);
nor U46973 (N_46973,N_46575,N_46557);
or U46974 (N_46974,N_46717,N_46662);
xor U46975 (N_46975,N_46599,N_46629);
and U46976 (N_46976,N_46516,N_46716);
or U46977 (N_46977,N_46644,N_46524);
nor U46978 (N_46978,N_46524,N_46506);
or U46979 (N_46979,N_46513,N_46548);
or U46980 (N_46980,N_46674,N_46585);
or U46981 (N_46981,N_46555,N_46682);
and U46982 (N_46982,N_46718,N_46559);
nor U46983 (N_46983,N_46684,N_46570);
xnor U46984 (N_46984,N_46543,N_46740);
and U46985 (N_46985,N_46735,N_46587);
nor U46986 (N_46986,N_46676,N_46641);
and U46987 (N_46987,N_46602,N_46678);
nor U46988 (N_46988,N_46676,N_46578);
and U46989 (N_46989,N_46516,N_46663);
nand U46990 (N_46990,N_46643,N_46512);
nor U46991 (N_46991,N_46670,N_46523);
or U46992 (N_46992,N_46558,N_46556);
nor U46993 (N_46993,N_46543,N_46553);
and U46994 (N_46994,N_46681,N_46738);
and U46995 (N_46995,N_46726,N_46550);
and U46996 (N_46996,N_46593,N_46529);
and U46997 (N_46997,N_46731,N_46712);
or U46998 (N_46998,N_46744,N_46740);
xnor U46999 (N_46999,N_46617,N_46578);
nand U47000 (N_47000,N_46808,N_46904);
xnor U47001 (N_47001,N_46906,N_46836);
xor U47002 (N_47002,N_46866,N_46797);
and U47003 (N_47003,N_46873,N_46984);
nand U47004 (N_47004,N_46787,N_46840);
or U47005 (N_47005,N_46767,N_46853);
nor U47006 (N_47006,N_46788,N_46886);
nand U47007 (N_47007,N_46934,N_46884);
nand U47008 (N_47008,N_46789,N_46942);
and U47009 (N_47009,N_46938,N_46895);
or U47010 (N_47010,N_46946,N_46928);
and U47011 (N_47011,N_46969,N_46781);
and U47012 (N_47012,N_46852,N_46911);
and U47013 (N_47013,N_46769,N_46972);
and U47014 (N_47014,N_46939,N_46958);
and U47015 (N_47015,N_46815,N_46790);
nand U47016 (N_47016,N_46779,N_46844);
nor U47017 (N_47017,N_46849,N_46755);
nor U47018 (N_47018,N_46773,N_46801);
xor U47019 (N_47019,N_46960,N_46994);
nor U47020 (N_47020,N_46912,N_46835);
nand U47021 (N_47021,N_46992,N_46964);
xor U47022 (N_47022,N_46855,N_46764);
nor U47023 (N_47023,N_46876,N_46830);
nor U47024 (N_47024,N_46783,N_46763);
nand U47025 (N_47025,N_46976,N_46894);
xnor U47026 (N_47026,N_46899,N_46981);
or U47027 (N_47027,N_46777,N_46967);
xor U47028 (N_47028,N_46890,N_46766);
xnor U47029 (N_47029,N_46988,N_46796);
and U47030 (N_47030,N_46882,N_46881);
nor U47031 (N_47031,N_46819,N_46756);
nor U47032 (N_47032,N_46907,N_46936);
and U47033 (N_47033,N_46803,N_46880);
nand U47034 (N_47034,N_46759,N_46956);
and U47035 (N_47035,N_46903,N_46999);
nand U47036 (N_47036,N_46768,N_46839);
and U47037 (N_47037,N_46891,N_46914);
nand U47038 (N_47038,N_46961,N_46924);
xor U47039 (N_47039,N_46950,N_46814);
nor U47040 (N_47040,N_46918,N_46838);
and U47041 (N_47041,N_46887,N_46971);
nor U47042 (N_47042,N_46774,N_46793);
or U47043 (N_47043,N_46919,N_46871);
xor U47044 (N_47044,N_46868,N_46810);
xnor U47045 (N_47045,N_46879,N_46893);
or U47046 (N_47046,N_46856,N_46975);
and U47047 (N_47047,N_46905,N_46834);
nor U47048 (N_47048,N_46874,N_46983);
nor U47049 (N_47049,N_46927,N_46772);
xnor U47050 (N_47050,N_46888,N_46820);
nand U47051 (N_47051,N_46806,N_46933);
nor U47052 (N_47052,N_46923,N_46799);
nor U47053 (N_47053,N_46862,N_46900);
nand U47054 (N_47054,N_46829,N_46802);
or U47055 (N_47055,N_46869,N_46765);
nor U47056 (N_47056,N_46987,N_46861);
or U47057 (N_47057,N_46997,N_46889);
nor U47058 (N_47058,N_46800,N_46860);
nor U47059 (N_47059,N_46968,N_46935);
nor U47060 (N_47060,N_46877,N_46816);
xor U47061 (N_47061,N_46883,N_46798);
nor U47062 (N_47062,N_46771,N_46753);
nor U47063 (N_47063,N_46822,N_46915);
or U47064 (N_47064,N_46761,N_46752);
xor U47065 (N_47065,N_46782,N_46930);
nand U47066 (N_47066,N_46813,N_46841);
xnor U47067 (N_47067,N_46965,N_46991);
and U47068 (N_47068,N_46979,N_46897);
and U47069 (N_47069,N_46908,N_46986);
and U47070 (N_47070,N_46750,N_46995);
nor U47071 (N_47071,N_46842,N_46843);
or U47072 (N_47072,N_46931,N_46922);
xor U47073 (N_47073,N_46867,N_46809);
nor U47074 (N_47074,N_46825,N_46932);
and U47075 (N_47075,N_46885,N_46947);
nand U47076 (N_47076,N_46859,N_46864);
nor U47077 (N_47077,N_46821,N_46985);
nor U47078 (N_47078,N_46832,N_46952);
nand U47079 (N_47079,N_46827,N_46959);
nor U47080 (N_47080,N_46762,N_46875);
and U47081 (N_47081,N_46949,N_46954);
nand U47082 (N_47082,N_46963,N_46953);
xnor U47083 (N_47083,N_46845,N_46902);
nor U47084 (N_47084,N_46955,N_46831);
and U47085 (N_47085,N_46898,N_46848);
or U47086 (N_47086,N_46920,N_46758);
nor U47087 (N_47087,N_46966,N_46978);
xor U47088 (N_47088,N_46780,N_46754);
nor U47089 (N_47089,N_46917,N_46757);
nor U47090 (N_47090,N_46805,N_46962);
xnor U47091 (N_47091,N_46824,N_46977);
nand U47092 (N_47092,N_46850,N_46998);
and U47093 (N_47093,N_46812,N_46770);
nand U47094 (N_47094,N_46878,N_46785);
nor U47095 (N_47095,N_46943,N_46921);
and U47096 (N_47096,N_46828,N_46851);
nor U47097 (N_47097,N_46926,N_46760);
and U47098 (N_47098,N_46854,N_46823);
or U47099 (N_47099,N_46892,N_46993);
nor U47100 (N_47100,N_46872,N_46973);
nor U47101 (N_47101,N_46982,N_46996);
and U47102 (N_47102,N_46945,N_46807);
xor U47103 (N_47103,N_46865,N_46896);
or U47104 (N_47104,N_46846,N_46944);
or U47105 (N_47105,N_46786,N_46910);
xor U47106 (N_47106,N_46795,N_46990);
xor U47107 (N_47107,N_46775,N_46901);
nor U47108 (N_47108,N_46974,N_46870);
and U47109 (N_47109,N_46794,N_46941);
nand U47110 (N_47110,N_46948,N_46909);
and U47111 (N_47111,N_46925,N_46863);
xor U47112 (N_47112,N_46811,N_46792);
or U47113 (N_47113,N_46940,N_46776);
nor U47114 (N_47114,N_46847,N_46957);
or U47115 (N_47115,N_46916,N_46778);
nor U47116 (N_47116,N_46784,N_46817);
nand U47117 (N_47117,N_46826,N_46857);
nand U47118 (N_47118,N_46818,N_46751);
xnor U47119 (N_47119,N_46989,N_46804);
xor U47120 (N_47120,N_46833,N_46970);
or U47121 (N_47121,N_46980,N_46858);
nor U47122 (N_47122,N_46929,N_46937);
xor U47123 (N_47123,N_46837,N_46913);
and U47124 (N_47124,N_46951,N_46791);
and U47125 (N_47125,N_46909,N_46883);
xor U47126 (N_47126,N_46879,N_46932);
nor U47127 (N_47127,N_46930,N_46911);
nor U47128 (N_47128,N_46751,N_46778);
xnor U47129 (N_47129,N_46850,N_46895);
nand U47130 (N_47130,N_46856,N_46783);
xor U47131 (N_47131,N_46993,N_46891);
xor U47132 (N_47132,N_46887,N_46805);
nor U47133 (N_47133,N_46825,N_46757);
nor U47134 (N_47134,N_46865,N_46770);
or U47135 (N_47135,N_46911,N_46915);
nand U47136 (N_47136,N_46846,N_46985);
and U47137 (N_47137,N_46927,N_46903);
nor U47138 (N_47138,N_46906,N_46838);
and U47139 (N_47139,N_46884,N_46917);
or U47140 (N_47140,N_46915,N_46997);
and U47141 (N_47141,N_46768,N_46844);
and U47142 (N_47142,N_46930,N_46992);
nand U47143 (N_47143,N_46991,N_46997);
or U47144 (N_47144,N_46897,N_46888);
nor U47145 (N_47145,N_46763,N_46776);
nand U47146 (N_47146,N_46786,N_46847);
xnor U47147 (N_47147,N_46956,N_46903);
nor U47148 (N_47148,N_46887,N_46788);
or U47149 (N_47149,N_46753,N_46896);
or U47150 (N_47150,N_46983,N_46796);
xor U47151 (N_47151,N_46901,N_46779);
nand U47152 (N_47152,N_46926,N_46750);
nor U47153 (N_47153,N_46994,N_46912);
nor U47154 (N_47154,N_46922,N_46863);
or U47155 (N_47155,N_46825,N_46872);
nor U47156 (N_47156,N_46958,N_46854);
nand U47157 (N_47157,N_46981,N_46883);
xor U47158 (N_47158,N_46772,N_46750);
nor U47159 (N_47159,N_46861,N_46755);
or U47160 (N_47160,N_46798,N_46759);
or U47161 (N_47161,N_46892,N_46817);
nor U47162 (N_47162,N_46849,N_46793);
or U47163 (N_47163,N_46885,N_46931);
xor U47164 (N_47164,N_46768,N_46927);
nand U47165 (N_47165,N_46786,N_46826);
nand U47166 (N_47166,N_46968,N_46872);
and U47167 (N_47167,N_46943,N_46919);
and U47168 (N_47168,N_46789,N_46983);
nand U47169 (N_47169,N_46868,N_46871);
xor U47170 (N_47170,N_46862,N_46907);
nor U47171 (N_47171,N_46917,N_46985);
nand U47172 (N_47172,N_46770,N_46831);
and U47173 (N_47173,N_46854,N_46774);
nand U47174 (N_47174,N_46956,N_46845);
nand U47175 (N_47175,N_46857,N_46759);
xor U47176 (N_47176,N_46830,N_46950);
nand U47177 (N_47177,N_46821,N_46928);
nor U47178 (N_47178,N_46892,N_46838);
and U47179 (N_47179,N_46851,N_46823);
or U47180 (N_47180,N_46853,N_46793);
or U47181 (N_47181,N_46903,N_46905);
and U47182 (N_47182,N_46973,N_46843);
nor U47183 (N_47183,N_46842,N_46763);
nor U47184 (N_47184,N_46823,N_46927);
xnor U47185 (N_47185,N_46755,N_46854);
nand U47186 (N_47186,N_46916,N_46907);
xnor U47187 (N_47187,N_46976,N_46750);
or U47188 (N_47188,N_46776,N_46804);
or U47189 (N_47189,N_46773,N_46784);
and U47190 (N_47190,N_46883,N_46829);
nand U47191 (N_47191,N_46764,N_46848);
and U47192 (N_47192,N_46751,N_46864);
xnor U47193 (N_47193,N_46930,N_46817);
or U47194 (N_47194,N_46974,N_46781);
nor U47195 (N_47195,N_46872,N_46786);
and U47196 (N_47196,N_46895,N_46913);
or U47197 (N_47197,N_46766,N_46897);
nand U47198 (N_47198,N_46762,N_46969);
nor U47199 (N_47199,N_46854,N_46842);
or U47200 (N_47200,N_46946,N_46999);
nand U47201 (N_47201,N_46941,N_46788);
or U47202 (N_47202,N_46820,N_46917);
or U47203 (N_47203,N_46906,N_46776);
and U47204 (N_47204,N_46885,N_46942);
and U47205 (N_47205,N_46972,N_46750);
nor U47206 (N_47206,N_46928,N_46769);
and U47207 (N_47207,N_46764,N_46951);
or U47208 (N_47208,N_46871,N_46941);
nor U47209 (N_47209,N_46898,N_46816);
or U47210 (N_47210,N_46894,N_46978);
nand U47211 (N_47211,N_46902,N_46831);
and U47212 (N_47212,N_46876,N_46755);
nand U47213 (N_47213,N_46767,N_46894);
nor U47214 (N_47214,N_46843,N_46817);
xnor U47215 (N_47215,N_46796,N_46967);
xor U47216 (N_47216,N_46792,N_46820);
or U47217 (N_47217,N_46791,N_46977);
nor U47218 (N_47218,N_46878,N_46834);
or U47219 (N_47219,N_46989,N_46763);
and U47220 (N_47220,N_46797,N_46895);
xor U47221 (N_47221,N_46786,N_46956);
xnor U47222 (N_47222,N_46913,N_46899);
and U47223 (N_47223,N_46750,N_46817);
and U47224 (N_47224,N_46789,N_46868);
nor U47225 (N_47225,N_46850,N_46797);
nor U47226 (N_47226,N_46775,N_46935);
xor U47227 (N_47227,N_46771,N_46964);
and U47228 (N_47228,N_46828,N_46964);
and U47229 (N_47229,N_46935,N_46846);
and U47230 (N_47230,N_46927,N_46787);
or U47231 (N_47231,N_46925,N_46754);
and U47232 (N_47232,N_46947,N_46898);
or U47233 (N_47233,N_46941,N_46845);
xor U47234 (N_47234,N_46921,N_46797);
and U47235 (N_47235,N_46986,N_46822);
nor U47236 (N_47236,N_46807,N_46888);
nor U47237 (N_47237,N_46947,N_46924);
xnor U47238 (N_47238,N_46974,N_46778);
or U47239 (N_47239,N_46991,N_46787);
nor U47240 (N_47240,N_46886,N_46854);
nor U47241 (N_47241,N_46931,N_46987);
nor U47242 (N_47242,N_46999,N_46937);
xnor U47243 (N_47243,N_46964,N_46757);
or U47244 (N_47244,N_46802,N_46925);
and U47245 (N_47245,N_46912,N_46917);
or U47246 (N_47246,N_46862,N_46798);
nor U47247 (N_47247,N_46954,N_46907);
or U47248 (N_47248,N_46768,N_46918);
xor U47249 (N_47249,N_46759,N_46750);
nand U47250 (N_47250,N_47062,N_47133);
or U47251 (N_47251,N_47045,N_47110);
nor U47252 (N_47252,N_47094,N_47016);
nor U47253 (N_47253,N_47019,N_47187);
nand U47254 (N_47254,N_47178,N_47018);
nand U47255 (N_47255,N_47236,N_47223);
xnor U47256 (N_47256,N_47122,N_47215);
and U47257 (N_47257,N_47202,N_47097);
and U47258 (N_47258,N_47238,N_47130);
xnor U47259 (N_47259,N_47210,N_47084);
and U47260 (N_47260,N_47175,N_47224);
or U47261 (N_47261,N_47172,N_47184);
xor U47262 (N_47262,N_47243,N_47056);
xnor U47263 (N_47263,N_47031,N_47129);
or U47264 (N_47264,N_47154,N_47029);
or U47265 (N_47265,N_47198,N_47149);
xor U47266 (N_47266,N_47103,N_47231);
nand U47267 (N_47267,N_47022,N_47136);
nor U47268 (N_47268,N_47240,N_47244);
and U47269 (N_47269,N_47118,N_47144);
or U47270 (N_47270,N_47035,N_47214);
nand U47271 (N_47271,N_47179,N_47105);
nor U47272 (N_47272,N_47192,N_47235);
and U47273 (N_47273,N_47128,N_47170);
xor U47274 (N_47274,N_47140,N_47125);
nand U47275 (N_47275,N_47003,N_47005);
or U47276 (N_47276,N_47071,N_47162);
nand U47277 (N_47277,N_47226,N_47209);
xor U47278 (N_47278,N_47158,N_47222);
nor U47279 (N_47279,N_47163,N_47063);
nor U47280 (N_47280,N_47119,N_47091);
and U47281 (N_47281,N_47025,N_47239);
xnor U47282 (N_47282,N_47007,N_47190);
and U47283 (N_47283,N_47048,N_47002);
xor U47284 (N_47284,N_47193,N_47123);
nand U47285 (N_47285,N_47164,N_47242);
xor U47286 (N_47286,N_47078,N_47169);
nor U47287 (N_47287,N_47058,N_47180);
nand U47288 (N_47288,N_47150,N_47141);
xnor U47289 (N_47289,N_47027,N_47167);
and U47290 (N_47290,N_47168,N_47127);
nand U47291 (N_47291,N_47032,N_47199);
or U47292 (N_47292,N_47006,N_47088);
nor U47293 (N_47293,N_47039,N_47173);
or U47294 (N_47294,N_47153,N_47038);
xnor U47295 (N_47295,N_47247,N_47213);
xor U47296 (N_47296,N_47092,N_47227);
nor U47297 (N_47297,N_47060,N_47200);
or U47298 (N_47298,N_47036,N_47049);
or U47299 (N_47299,N_47233,N_47040);
or U47300 (N_47300,N_47157,N_47143);
nand U47301 (N_47301,N_47159,N_47237);
nor U47302 (N_47302,N_47126,N_47249);
nand U47303 (N_47303,N_47161,N_47241);
nor U47304 (N_47304,N_47174,N_47013);
xor U47305 (N_47305,N_47204,N_47120);
nand U47306 (N_47306,N_47042,N_47203);
or U47307 (N_47307,N_47081,N_47074);
xnor U47308 (N_47308,N_47121,N_47052);
xor U47309 (N_47309,N_47219,N_47070);
and U47310 (N_47310,N_47107,N_47211);
and U47311 (N_47311,N_47023,N_47218);
and U47312 (N_47312,N_47037,N_47082);
nor U47313 (N_47313,N_47083,N_47185);
xor U47314 (N_47314,N_47044,N_47051);
nor U47315 (N_47315,N_47024,N_47139);
and U47316 (N_47316,N_47101,N_47191);
xor U47317 (N_47317,N_47232,N_47225);
nor U47318 (N_47318,N_47059,N_47248);
xor U47319 (N_47319,N_47017,N_47011);
or U47320 (N_47320,N_47152,N_47196);
xnor U47321 (N_47321,N_47033,N_47061);
or U47322 (N_47322,N_47020,N_47069);
xnor U47323 (N_47323,N_47183,N_47113);
xor U47324 (N_47324,N_47166,N_47212);
nand U47325 (N_47325,N_47068,N_47115);
xor U47326 (N_47326,N_47089,N_47221);
nor U47327 (N_47327,N_47197,N_47230);
xor U47328 (N_47328,N_47234,N_47100);
nand U47329 (N_47329,N_47015,N_47057);
and U47330 (N_47330,N_47028,N_47104);
and U47331 (N_47331,N_47156,N_47102);
nor U47332 (N_47332,N_47181,N_47217);
xor U47333 (N_47333,N_47086,N_47142);
or U47334 (N_47334,N_47077,N_47008);
nor U47335 (N_47335,N_47080,N_47228);
and U47336 (N_47336,N_47114,N_47116);
and U47337 (N_47337,N_47155,N_47009);
nor U47338 (N_47338,N_47041,N_47064);
or U47339 (N_47339,N_47216,N_47021);
xor U47340 (N_47340,N_47053,N_47112);
and U47341 (N_47341,N_47055,N_47186);
nand U47342 (N_47342,N_47066,N_47004);
xor U47343 (N_47343,N_47054,N_47134);
nor U47344 (N_47344,N_47188,N_47067);
or U47345 (N_47345,N_47076,N_47165);
xor U47346 (N_47346,N_47206,N_47117);
or U47347 (N_47347,N_47151,N_47138);
or U47348 (N_47348,N_47245,N_47000);
xor U47349 (N_47349,N_47099,N_47090);
and U47350 (N_47350,N_47109,N_47135);
xor U47351 (N_47351,N_47131,N_47085);
nand U47352 (N_47352,N_47010,N_47098);
and U47353 (N_47353,N_47207,N_47137);
nand U47354 (N_47354,N_47047,N_47079);
nand U47355 (N_47355,N_47096,N_47201);
nor U47356 (N_47356,N_47205,N_47189);
xor U47357 (N_47357,N_47124,N_47012);
nor U47358 (N_47358,N_47026,N_47148);
nand U47359 (N_47359,N_47208,N_47065);
xnor U47360 (N_47360,N_47229,N_47014);
or U47361 (N_47361,N_47132,N_47046);
or U47362 (N_47362,N_47075,N_47246);
xor U47363 (N_47363,N_47043,N_47220);
xor U47364 (N_47364,N_47194,N_47050);
and U47365 (N_47365,N_47176,N_47034);
xnor U47366 (N_47366,N_47072,N_47171);
nor U47367 (N_47367,N_47087,N_47177);
nand U47368 (N_47368,N_47108,N_47030);
or U47369 (N_47369,N_47001,N_47147);
nor U47370 (N_47370,N_47195,N_47146);
nor U47371 (N_47371,N_47111,N_47182);
xor U47372 (N_47372,N_47073,N_47145);
and U47373 (N_47373,N_47095,N_47106);
nor U47374 (N_47374,N_47093,N_47160);
nand U47375 (N_47375,N_47007,N_47206);
and U47376 (N_47376,N_47163,N_47049);
nor U47377 (N_47377,N_47070,N_47017);
or U47378 (N_47378,N_47172,N_47249);
nand U47379 (N_47379,N_47051,N_47020);
or U47380 (N_47380,N_47155,N_47052);
and U47381 (N_47381,N_47036,N_47193);
xor U47382 (N_47382,N_47026,N_47229);
nand U47383 (N_47383,N_47199,N_47117);
nor U47384 (N_47384,N_47180,N_47035);
or U47385 (N_47385,N_47146,N_47214);
nand U47386 (N_47386,N_47007,N_47015);
or U47387 (N_47387,N_47226,N_47218);
or U47388 (N_47388,N_47070,N_47064);
and U47389 (N_47389,N_47217,N_47147);
xnor U47390 (N_47390,N_47156,N_47023);
or U47391 (N_47391,N_47029,N_47226);
nor U47392 (N_47392,N_47009,N_47032);
nand U47393 (N_47393,N_47172,N_47171);
or U47394 (N_47394,N_47095,N_47013);
or U47395 (N_47395,N_47182,N_47056);
and U47396 (N_47396,N_47119,N_47243);
or U47397 (N_47397,N_47123,N_47142);
xnor U47398 (N_47398,N_47034,N_47198);
and U47399 (N_47399,N_47029,N_47033);
nor U47400 (N_47400,N_47026,N_47199);
and U47401 (N_47401,N_47083,N_47008);
and U47402 (N_47402,N_47008,N_47040);
nor U47403 (N_47403,N_47176,N_47233);
nand U47404 (N_47404,N_47179,N_47099);
nand U47405 (N_47405,N_47008,N_47150);
nor U47406 (N_47406,N_47027,N_47096);
xor U47407 (N_47407,N_47233,N_47204);
xor U47408 (N_47408,N_47216,N_47220);
xor U47409 (N_47409,N_47094,N_47216);
and U47410 (N_47410,N_47061,N_47010);
xor U47411 (N_47411,N_47056,N_47145);
and U47412 (N_47412,N_47033,N_47114);
xor U47413 (N_47413,N_47124,N_47091);
xnor U47414 (N_47414,N_47157,N_47079);
nor U47415 (N_47415,N_47235,N_47110);
xor U47416 (N_47416,N_47010,N_47148);
or U47417 (N_47417,N_47167,N_47040);
or U47418 (N_47418,N_47063,N_47195);
or U47419 (N_47419,N_47199,N_47140);
or U47420 (N_47420,N_47029,N_47139);
xnor U47421 (N_47421,N_47011,N_47205);
xor U47422 (N_47422,N_47203,N_47082);
xor U47423 (N_47423,N_47243,N_47246);
nor U47424 (N_47424,N_47020,N_47104);
or U47425 (N_47425,N_47202,N_47092);
nor U47426 (N_47426,N_47096,N_47220);
xor U47427 (N_47427,N_47002,N_47164);
and U47428 (N_47428,N_47071,N_47056);
and U47429 (N_47429,N_47076,N_47154);
xnor U47430 (N_47430,N_47143,N_47093);
and U47431 (N_47431,N_47197,N_47027);
or U47432 (N_47432,N_47172,N_47130);
or U47433 (N_47433,N_47110,N_47176);
or U47434 (N_47434,N_47138,N_47237);
nand U47435 (N_47435,N_47055,N_47067);
nor U47436 (N_47436,N_47014,N_47022);
and U47437 (N_47437,N_47200,N_47174);
nor U47438 (N_47438,N_47005,N_47222);
nand U47439 (N_47439,N_47119,N_47191);
and U47440 (N_47440,N_47123,N_47186);
and U47441 (N_47441,N_47133,N_47201);
nand U47442 (N_47442,N_47248,N_47247);
or U47443 (N_47443,N_47092,N_47204);
nor U47444 (N_47444,N_47030,N_47176);
and U47445 (N_47445,N_47075,N_47048);
nor U47446 (N_47446,N_47096,N_47121);
nor U47447 (N_47447,N_47147,N_47178);
nor U47448 (N_47448,N_47126,N_47071);
nand U47449 (N_47449,N_47037,N_47031);
and U47450 (N_47450,N_47021,N_47024);
and U47451 (N_47451,N_47151,N_47131);
and U47452 (N_47452,N_47128,N_47101);
nor U47453 (N_47453,N_47015,N_47142);
and U47454 (N_47454,N_47093,N_47072);
xnor U47455 (N_47455,N_47209,N_47033);
and U47456 (N_47456,N_47058,N_47081);
nor U47457 (N_47457,N_47240,N_47028);
xor U47458 (N_47458,N_47117,N_47140);
and U47459 (N_47459,N_47129,N_47177);
nand U47460 (N_47460,N_47152,N_47173);
nand U47461 (N_47461,N_47157,N_47023);
and U47462 (N_47462,N_47126,N_47198);
nand U47463 (N_47463,N_47170,N_47027);
nor U47464 (N_47464,N_47134,N_47058);
and U47465 (N_47465,N_47184,N_47177);
nand U47466 (N_47466,N_47223,N_47129);
and U47467 (N_47467,N_47093,N_47071);
nor U47468 (N_47468,N_47035,N_47161);
nor U47469 (N_47469,N_47130,N_47030);
nand U47470 (N_47470,N_47121,N_47141);
or U47471 (N_47471,N_47227,N_47028);
nand U47472 (N_47472,N_47120,N_47112);
nor U47473 (N_47473,N_47147,N_47247);
nor U47474 (N_47474,N_47226,N_47175);
or U47475 (N_47475,N_47093,N_47077);
nand U47476 (N_47476,N_47109,N_47190);
and U47477 (N_47477,N_47135,N_47244);
xnor U47478 (N_47478,N_47046,N_47216);
and U47479 (N_47479,N_47117,N_47097);
nand U47480 (N_47480,N_47233,N_47207);
xor U47481 (N_47481,N_47080,N_47196);
xnor U47482 (N_47482,N_47048,N_47247);
xor U47483 (N_47483,N_47062,N_47091);
or U47484 (N_47484,N_47091,N_47166);
xnor U47485 (N_47485,N_47213,N_47188);
or U47486 (N_47486,N_47151,N_47136);
or U47487 (N_47487,N_47023,N_47247);
or U47488 (N_47488,N_47223,N_47010);
nand U47489 (N_47489,N_47182,N_47046);
and U47490 (N_47490,N_47026,N_47203);
and U47491 (N_47491,N_47095,N_47244);
or U47492 (N_47492,N_47141,N_47057);
xor U47493 (N_47493,N_47059,N_47062);
and U47494 (N_47494,N_47215,N_47052);
nand U47495 (N_47495,N_47243,N_47030);
or U47496 (N_47496,N_47060,N_47244);
nor U47497 (N_47497,N_47105,N_47085);
or U47498 (N_47498,N_47018,N_47033);
xnor U47499 (N_47499,N_47066,N_47184);
xor U47500 (N_47500,N_47339,N_47484);
or U47501 (N_47501,N_47331,N_47417);
xor U47502 (N_47502,N_47372,N_47318);
xor U47503 (N_47503,N_47340,N_47303);
xnor U47504 (N_47504,N_47492,N_47352);
xor U47505 (N_47505,N_47366,N_47351);
xnor U47506 (N_47506,N_47408,N_47281);
or U47507 (N_47507,N_47479,N_47411);
and U47508 (N_47508,N_47427,N_47301);
nand U47509 (N_47509,N_47498,N_47461);
nand U47510 (N_47510,N_47403,N_47380);
nand U47511 (N_47511,N_47368,N_47347);
nand U47512 (N_47512,N_47310,N_47418);
nand U47513 (N_47513,N_47273,N_47291);
xnor U47514 (N_47514,N_47322,N_47425);
nor U47515 (N_47515,N_47353,N_47258);
xor U47516 (N_47516,N_47299,N_47376);
nand U47517 (N_47517,N_47332,N_47496);
nand U47518 (N_47518,N_47442,N_47259);
or U47519 (N_47519,N_47410,N_47487);
xnor U47520 (N_47520,N_47374,N_47428);
nand U47521 (N_47521,N_47334,N_47486);
or U47522 (N_47522,N_47489,N_47356);
nor U47523 (N_47523,N_47337,N_47493);
nor U47524 (N_47524,N_47253,N_47469);
nand U47525 (N_47525,N_47296,N_47468);
xnor U47526 (N_47526,N_47305,N_47270);
and U47527 (N_47527,N_47289,N_47494);
nor U47528 (N_47528,N_47354,N_47321);
nand U47529 (N_47529,N_47422,N_47429);
xor U47530 (N_47530,N_47464,N_47458);
and U47531 (N_47531,N_47459,N_47473);
nor U47532 (N_47532,N_47395,N_47488);
nand U47533 (N_47533,N_47432,N_47371);
xor U47534 (N_47534,N_47381,N_47476);
nand U47535 (N_47535,N_47424,N_47283);
nand U47536 (N_47536,N_47392,N_47415);
and U47537 (N_47537,N_47406,N_47483);
or U47538 (N_47538,N_47387,N_47390);
or U47539 (N_47539,N_47314,N_47388);
xnor U47540 (N_47540,N_47478,N_47325);
nand U47541 (N_47541,N_47295,N_47447);
or U47542 (N_47542,N_47414,N_47364);
nor U47543 (N_47543,N_47306,N_47319);
nor U47544 (N_47544,N_47435,N_47470);
xor U47545 (N_47545,N_47309,N_47378);
xor U47546 (N_47546,N_47383,N_47480);
or U47547 (N_47547,N_47307,N_47402);
or U47548 (N_47548,N_47272,N_47426);
or U47549 (N_47549,N_47385,N_47439);
xor U47550 (N_47550,N_47349,N_47431);
or U47551 (N_47551,N_47419,N_47274);
or U47552 (N_47552,N_47278,N_47257);
or U47553 (N_47553,N_47477,N_47275);
nor U47554 (N_47554,N_47297,N_47269);
nor U47555 (N_47555,N_47328,N_47450);
or U47556 (N_47556,N_47474,N_47370);
nor U47557 (N_47557,N_47443,N_47324);
nor U47558 (N_47558,N_47287,N_47454);
or U47559 (N_47559,N_47290,N_47421);
nor U47560 (N_47560,N_47379,N_47333);
xnor U47561 (N_47561,N_47311,N_47382);
nor U47562 (N_47562,N_47449,N_47455);
nor U47563 (N_47563,N_47327,N_47282);
and U47564 (N_47564,N_47361,N_47495);
xnor U47565 (N_47565,N_47285,N_47377);
or U47566 (N_47566,N_47262,N_47267);
and U47567 (N_47567,N_47467,N_47440);
xor U47568 (N_47568,N_47389,N_47256);
and U47569 (N_47569,N_47280,N_47396);
or U47570 (N_47570,N_47346,N_47350);
xor U47571 (N_47571,N_47336,N_47357);
and U47572 (N_47572,N_47264,N_47263);
and U47573 (N_47573,N_47335,N_47416);
and U47574 (N_47574,N_47386,N_47326);
nand U47575 (N_47575,N_47355,N_47399);
and U47576 (N_47576,N_47279,N_47441);
nand U47577 (N_47577,N_47423,N_47323);
nand U47578 (N_47578,N_47348,N_47313);
nand U47579 (N_47579,N_47452,N_47394);
nand U47580 (N_47580,N_47445,N_47293);
xor U47581 (N_47581,N_47453,N_47292);
xor U47582 (N_47582,N_47300,N_47400);
nor U47583 (N_47583,N_47471,N_47315);
xnor U47584 (N_47584,N_47252,N_47276);
and U47585 (N_47585,N_47491,N_47457);
and U47586 (N_47586,N_47434,N_47451);
and U47587 (N_47587,N_47284,N_47437);
xnor U47588 (N_47588,N_47298,N_47251);
nor U47589 (N_47589,N_47344,N_47260);
nor U47590 (N_47590,N_47456,N_47444);
and U47591 (N_47591,N_47345,N_47413);
nand U47592 (N_47592,N_47482,N_47472);
or U47593 (N_47593,N_47343,N_47294);
or U47594 (N_47594,N_47430,N_47288);
nand U47595 (N_47595,N_47365,N_47433);
and U47596 (N_47596,N_47277,N_47286);
nor U47597 (N_47597,N_47254,N_47490);
xor U47598 (N_47598,N_47317,N_47271);
and U47599 (N_47599,N_47404,N_47463);
xnor U47600 (N_47600,N_47407,N_47250);
nor U47601 (N_47601,N_47363,N_47360);
and U47602 (N_47602,N_47312,N_47420);
nand U47603 (N_47603,N_47261,N_47405);
xor U47604 (N_47604,N_47369,N_47397);
and U47605 (N_47605,N_47412,N_47268);
or U47606 (N_47606,N_47398,N_47448);
nor U47607 (N_47607,N_47409,N_47255);
and U47608 (N_47608,N_47265,N_47329);
nor U47609 (N_47609,N_47266,N_47475);
nand U47610 (N_47610,N_47367,N_47391);
nor U47611 (N_47611,N_47438,N_47316);
nor U47612 (N_47612,N_47338,N_47320);
and U47613 (N_47613,N_47330,N_47465);
nor U47614 (N_47614,N_47393,N_47446);
and U47615 (N_47615,N_47373,N_47460);
and U47616 (N_47616,N_47308,N_47485);
xor U47617 (N_47617,N_47384,N_47304);
nand U47618 (N_47618,N_47359,N_47302);
xnor U47619 (N_47619,N_47436,N_47466);
and U47620 (N_47620,N_47481,N_47497);
nand U47621 (N_47621,N_47401,N_47375);
nor U47622 (N_47622,N_47341,N_47358);
xor U47623 (N_47623,N_47362,N_47499);
nor U47624 (N_47624,N_47342,N_47462);
nand U47625 (N_47625,N_47287,N_47373);
nor U47626 (N_47626,N_47308,N_47263);
or U47627 (N_47627,N_47493,N_47333);
nor U47628 (N_47628,N_47419,N_47307);
and U47629 (N_47629,N_47285,N_47309);
or U47630 (N_47630,N_47416,N_47341);
and U47631 (N_47631,N_47435,N_47358);
nand U47632 (N_47632,N_47383,N_47380);
xor U47633 (N_47633,N_47337,N_47378);
and U47634 (N_47634,N_47372,N_47252);
nor U47635 (N_47635,N_47261,N_47437);
nor U47636 (N_47636,N_47397,N_47291);
xor U47637 (N_47637,N_47377,N_47436);
nor U47638 (N_47638,N_47488,N_47491);
and U47639 (N_47639,N_47388,N_47373);
or U47640 (N_47640,N_47327,N_47489);
or U47641 (N_47641,N_47402,N_47469);
or U47642 (N_47642,N_47374,N_47438);
and U47643 (N_47643,N_47476,N_47280);
nand U47644 (N_47644,N_47492,N_47293);
and U47645 (N_47645,N_47348,N_47470);
or U47646 (N_47646,N_47374,N_47460);
nand U47647 (N_47647,N_47465,N_47430);
and U47648 (N_47648,N_47375,N_47315);
nand U47649 (N_47649,N_47275,N_47426);
or U47650 (N_47650,N_47308,N_47408);
and U47651 (N_47651,N_47307,N_47386);
or U47652 (N_47652,N_47366,N_47299);
and U47653 (N_47653,N_47327,N_47404);
and U47654 (N_47654,N_47424,N_47455);
xnor U47655 (N_47655,N_47355,N_47273);
xnor U47656 (N_47656,N_47402,N_47428);
xnor U47657 (N_47657,N_47446,N_47397);
or U47658 (N_47658,N_47339,N_47420);
xnor U47659 (N_47659,N_47353,N_47461);
xnor U47660 (N_47660,N_47429,N_47447);
nand U47661 (N_47661,N_47333,N_47337);
nand U47662 (N_47662,N_47318,N_47362);
xor U47663 (N_47663,N_47351,N_47432);
or U47664 (N_47664,N_47462,N_47274);
or U47665 (N_47665,N_47310,N_47316);
nor U47666 (N_47666,N_47298,N_47467);
nand U47667 (N_47667,N_47491,N_47270);
nand U47668 (N_47668,N_47310,N_47385);
nor U47669 (N_47669,N_47394,N_47442);
or U47670 (N_47670,N_47385,N_47466);
xor U47671 (N_47671,N_47286,N_47379);
xnor U47672 (N_47672,N_47322,N_47441);
or U47673 (N_47673,N_47374,N_47262);
xor U47674 (N_47674,N_47389,N_47385);
nand U47675 (N_47675,N_47497,N_47305);
xnor U47676 (N_47676,N_47289,N_47444);
xnor U47677 (N_47677,N_47320,N_47495);
xor U47678 (N_47678,N_47318,N_47343);
xor U47679 (N_47679,N_47446,N_47466);
xor U47680 (N_47680,N_47422,N_47439);
nand U47681 (N_47681,N_47275,N_47483);
or U47682 (N_47682,N_47473,N_47338);
or U47683 (N_47683,N_47313,N_47497);
xor U47684 (N_47684,N_47272,N_47293);
xor U47685 (N_47685,N_47287,N_47345);
nand U47686 (N_47686,N_47401,N_47423);
xnor U47687 (N_47687,N_47489,N_47286);
xnor U47688 (N_47688,N_47341,N_47493);
nand U47689 (N_47689,N_47266,N_47385);
xnor U47690 (N_47690,N_47355,N_47334);
nand U47691 (N_47691,N_47494,N_47446);
nand U47692 (N_47692,N_47273,N_47404);
or U47693 (N_47693,N_47469,N_47302);
xnor U47694 (N_47694,N_47368,N_47461);
xnor U47695 (N_47695,N_47341,N_47472);
and U47696 (N_47696,N_47471,N_47311);
nor U47697 (N_47697,N_47396,N_47408);
and U47698 (N_47698,N_47312,N_47278);
or U47699 (N_47699,N_47419,N_47262);
nand U47700 (N_47700,N_47365,N_47385);
xor U47701 (N_47701,N_47446,N_47416);
xor U47702 (N_47702,N_47322,N_47287);
nor U47703 (N_47703,N_47421,N_47494);
nor U47704 (N_47704,N_47462,N_47357);
and U47705 (N_47705,N_47363,N_47435);
or U47706 (N_47706,N_47492,N_47446);
and U47707 (N_47707,N_47310,N_47488);
and U47708 (N_47708,N_47326,N_47282);
nand U47709 (N_47709,N_47362,N_47363);
xnor U47710 (N_47710,N_47404,N_47335);
nor U47711 (N_47711,N_47265,N_47403);
nor U47712 (N_47712,N_47302,N_47464);
nor U47713 (N_47713,N_47304,N_47294);
nor U47714 (N_47714,N_47489,N_47460);
or U47715 (N_47715,N_47324,N_47400);
nor U47716 (N_47716,N_47405,N_47391);
and U47717 (N_47717,N_47265,N_47372);
or U47718 (N_47718,N_47343,N_47359);
nor U47719 (N_47719,N_47267,N_47388);
xnor U47720 (N_47720,N_47434,N_47347);
nand U47721 (N_47721,N_47354,N_47323);
and U47722 (N_47722,N_47396,N_47343);
nor U47723 (N_47723,N_47349,N_47267);
and U47724 (N_47724,N_47268,N_47354);
and U47725 (N_47725,N_47448,N_47283);
xnor U47726 (N_47726,N_47455,N_47473);
or U47727 (N_47727,N_47363,N_47351);
and U47728 (N_47728,N_47265,N_47292);
and U47729 (N_47729,N_47441,N_47346);
and U47730 (N_47730,N_47354,N_47376);
xnor U47731 (N_47731,N_47472,N_47266);
nor U47732 (N_47732,N_47370,N_47490);
xnor U47733 (N_47733,N_47399,N_47482);
xor U47734 (N_47734,N_47346,N_47481);
xnor U47735 (N_47735,N_47283,N_47479);
and U47736 (N_47736,N_47437,N_47448);
or U47737 (N_47737,N_47318,N_47371);
or U47738 (N_47738,N_47464,N_47354);
and U47739 (N_47739,N_47493,N_47410);
nand U47740 (N_47740,N_47425,N_47456);
nor U47741 (N_47741,N_47432,N_47408);
nand U47742 (N_47742,N_47341,N_47300);
and U47743 (N_47743,N_47319,N_47385);
nand U47744 (N_47744,N_47260,N_47488);
nor U47745 (N_47745,N_47387,N_47345);
or U47746 (N_47746,N_47484,N_47480);
nor U47747 (N_47747,N_47481,N_47452);
and U47748 (N_47748,N_47492,N_47353);
xor U47749 (N_47749,N_47390,N_47437);
or U47750 (N_47750,N_47741,N_47591);
or U47751 (N_47751,N_47736,N_47651);
xor U47752 (N_47752,N_47742,N_47590);
nand U47753 (N_47753,N_47508,N_47705);
nand U47754 (N_47754,N_47602,N_47538);
nand U47755 (N_47755,N_47624,N_47711);
xnor U47756 (N_47756,N_47690,N_47504);
nand U47757 (N_47757,N_47635,N_47612);
and U47758 (N_47758,N_47517,N_47731);
nand U47759 (N_47759,N_47580,N_47687);
xnor U47760 (N_47760,N_47672,N_47565);
and U47761 (N_47761,N_47621,N_47664);
and U47762 (N_47762,N_47693,N_47737);
and U47763 (N_47763,N_47540,N_47558);
xnor U47764 (N_47764,N_47725,N_47668);
and U47765 (N_47765,N_47557,N_47746);
and U47766 (N_47766,N_47572,N_47665);
or U47767 (N_47767,N_47537,N_47600);
nand U47768 (N_47768,N_47535,N_47511);
or U47769 (N_47769,N_47619,N_47550);
or U47770 (N_47770,N_47653,N_47729);
or U47771 (N_47771,N_47556,N_47663);
and U47772 (N_47772,N_47534,N_47533);
nor U47773 (N_47773,N_47524,N_47539);
xnor U47774 (N_47774,N_47718,N_47607);
or U47775 (N_47775,N_47543,N_47532);
xnor U47776 (N_47776,N_47544,N_47738);
xor U47777 (N_47777,N_47520,N_47571);
and U47778 (N_47778,N_47573,N_47684);
or U47779 (N_47779,N_47515,N_47643);
nor U47780 (N_47780,N_47654,N_47542);
nor U47781 (N_47781,N_47709,N_47659);
xor U47782 (N_47782,N_47734,N_47747);
xnor U47783 (N_47783,N_47730,N_47715);
and U47784 (N_47784,N_47692,N_47623);
xor U47785 (N_47785,N_47714,N_47502);
xnor U47786 (N_47786,N_47723,N_47599);
xnor U47787 (N_47787,N_47509,N_47642);
or U47788 (N_47788,N_47507,N_47522);
xor U47789 (N_47789,N_47740,N_47547);
xnor U47790 (N_47790,N_47561,N_47581);
nand U47791 (N_47791,N_47649,N_47536);
and U47792 (N_47792,N_47720,N_47677);
and U47793 (N_47793,N_47697,N_47620);
or U47794 (N_47794,N_47548,N_47722);
nand U47795 (N_47795,N_47541,N_47598);
nand U47796 (N_47796,N_47671,N_47529);
xor U47797 (N_47797,N_47613,N_47562);
nand U47798 (N_47798,N_47606,N_47662);
or U47799 (N_47799,N_47566,N_47647);
xnor U47800 (N_47800,N_47685,N_47749);
xor U47801 (N_47801,N_47527,N_47658);
nor U47802 (N_47802,N_47552,N_47691);
xor U47803 (N_47803,N_47576,N_47513);
nand U47804 (N_47804,N_47616,N_47655);
or U47805 (N_47805,N_47501,N_47589);
nand U47806 (N_47806,N_47681,N_47628);
and U47807 (N_47807,N_47564,N_47622);
or U47808 (N_47808,N_47614,N_47500);
and U47809 (N_47809,N_47531,N_47596);
nand U47810 (N_47810,N_47644,N_47526);
nand U47811 (N_47811,N_47512,N_47514);
xnor U47812 (N_47812,N_47701,N_47673);
nand U47813 (N_47813,N_47587,N_47609);
and U47814 (N_47814,N_47639,N_47716);
or U47815 (N_47815,N_47595,N_47739);
and U47816 (N_47816,N_47678,N_47582);
nand U47817 (N_47817,N_47634,N_47676);
and U47818 (N_47818,N_47674,N_47604);
nor U47819 (N_47819,N_47555,N_47516);
nor U47820 (N_47820,N_47545,N_47510);
nor U47821 (N_47821,N_47625,N_47585);
xor U47822 (N_47822,N_47666,N_47583);
xnor U47823 (N_47823,N_47559,N_47577);
nor U47824 (N_47824,N_47611,N_47630);
and U47825 (N_47825,N_47632,N_47633);
or U47826 (N_47826,N_47724,N_47546);
nand U47827 (N_47827,N_47728,N_47615);
xnor U47828 (N_47828,N_47563,N_47650);
or U47829 (N_47829,N_47560,N_47682);
and U47830 (N_47830,N_47618,N_47626);
and U47831 (N_47831,N_47637,N_47610);
nand U47832 (N_47832,N_47719,N_47699);
and U47833 (N_47833,N_47567,N_47695);
nor U47834 (N_47834,N_47503,N_47594);
nand U47835 (N_47835,N_47703,N_47554);
nor U47836 (N_47836,N_47521,N_47704);
and U47837 (N_47837,N_47530,N_47603);
xnor U47838 (N_47838,N_47549,N_47707);
nor U47839 (N_47839,N_47656,N_47574);
nand U47840 (N_47840,N_47641,N_47601);
and U47841 (N_47841,N_47505,N_47575);
or U47842 (N_47842,N_47597,N_47584);
nand U47843 (N_47843,N_47688,N_47579);
and U47844 (N_47844,N_47721,N_47629);
nand U47845 (N_47845,N_47669,N_47702);
nand U47846 (N_47846,N_47679,N_47518);
xor U47847 (N_47847,N_47553,N_47745);
xor U47848 (N_47848,N_47694,N_47708);
or U47849 (N_47849,N_47660,N_47743);
or U47850 (N_47850,N_47578,N_47608);
or U47851 (N_47851,N_47569,N_47657);
or U47852 (N_47852,N_47588,N_47732);
nand U47853 (N_47853,N_47706,N_47661);
nor U47854 (N_47854,N_47645,N_47648);
xnor U47855 (N_47855,N_47675,N_47592);
xor U47856 (N_47856,N_47605,N_47710);
and U47857 (N_47857,N_47640,N_47726);
nand U47858 (N_47858,N_47689,N_47744);
and U47859 (N_47859,N_47586,N_47733);
nor U47860 (N_47860,N_47652,N_47717);
or U47861 (N_47861,N_47627,N_47523);
and U47862 (N_47862,N_47712,N_47735);
or U47863 (N_47863,N_47667,N_47700);
xor U47864 (N_47864,N_47568,N_47551);
and U47865 (N_47865,N_47696,N_47646);
or U47866 (N_47866,N_47698,N_47680);
nor U47867 (N_47867,N_47519,N_47636);
nor U47868 (N_47868,N_47683,N_47713);
or U47869 (N_47869,N_47593,N_47528);
nand U47870 (N_47870,N_47617,N_47570);
or U47871 (N_47871,N_47670,N_47638);
or U47872 (N_47872,N_47686,N_47727);
nand U47873 (N_47873,N_47525,N_47748);
and U47874 (N_47874,N_47631,N_47506);
nand U47875 (N_47875,N_47574,N_47676);
and U47876 (N_47876,N_47577,N_47663);
or U47877 (N_47877,N_47584,N_47511);
and U47878 (N_47878,N_47503,N_47732);
nor U47879 (N_47879,N_47731,N_47567);
xor U47880 (N_47880,N_47537,N_47673);
or U47881 (N_47881,N_47691,N_47613);
xor U47882 (N_47882,N_47604,N_47544);
nor U47883 (N_47883,N_47696,N_47629);
and U47884 (N_47884,N_47531,N_47527);
xnor U47885 (N_47885,N_47629,N_47539);
nor U47886 (N_47886,N_47628,N_47549);
xnor U47887 (N_47887,N_47709,N_47592);
nor U47888 (N_47888,N_47560,N_47646);
xnor U47889 (N_47889,N_47677,N_47718);
xnor U47890 (N_47890,N_47744,N_47559);
xnor U47891 (N_47891,N_47664,N_47673);
nor U47892 (N_47892,N_47512,N_47571);
xnor U47893 (N_47893,N_47580,N_47503);
and U47894 (N_47894,N_47653,N_47616);
nor U47895 (N_47895,N_47713,N_47592);
xor U47896 (N_47896,N_47635,N_47718);
xnor U47897 (N_47897,N_47683,N_47574);
nand U47898 (N_47898,N_47690,N_47511);
and U47899 (N_47899,N_47613,N_47749);
xor U47900 (N_47900,N_47516,N_47605);
nand U47901 (N_47901,N_47600,N_47741);
nor U47902 (N_47902,N_47544,N_47679);
nor U47903 (N_47903,N_47641,N_47552);
nor U47904 (N_47904,N_47629,N_47533);
nor U47905 (N_47905,N_47691,N_47681);
nand U47906 (N_47906,N_47691,N_47745);
nand U47907 (N_47907,N_47735,N_47502);
or U47908 (N_47908,N_47680,N_47722);
and U47909 (N_47909,N_47650,N_47715);
nor U47910 (N_47910,N_47663,N_47694);
nand U47911 (N_47911,N_47516,N_47574);
or U47912 (N_47912,N_47546,N_47573);
and U47913 (N_47913,N_47611,N_47661);
or U47914 (N_47914,N_47540,N_47531);
nand U47915 (N_47915,N_47685,N_47681);
and U47916 (N_47916,N_47528,N_47725);
nand U47917 (N_47917,N_47500,N_47581);
xnor U47918 (N_47918,N_47580,N_47624);
xor U47919 (N_47919,N_47683,N_47567);
or U47920 (N_47920,N_47518,N_47537);
xor U47921 (N_47921,N_47693,N_47530);
and U47922 (N_47922,N_47600,N_47706);
or U47923 (N_47923,N_47708,N_47599);
nor U47924 (N_47924,N_47629,N_47516);
xor U47925 (N_47925,N_47683,N_47661);
nor U47926 (N_47926,N_47670,N_47706);
and U47927 (N_47927,N_47742,N_47666);
nand U47928 (N_47928,N_47620,N_47664);
or U47929 (N_47929,N_47584,N_47665);
xnor U47930 (N_47930,N_47703,N_47672);
and U47931 (N_47931,N_47666,N_47641);
xnor U47932 (N_47932,N_47500,N_47573);
and U47933 (N_47933,N_47615,N_47627);
and U47934 (N_47934,N_47546,N_47643);
and U47935 (N_47935,N_47524,N_47549);
and U47936 (N_47936,N_47665,N_47628);
and U47937 (N_47937,N_47565,N_47720);
nor U47938 (N_47938,N_47631,N_47720);
nor U47939 (N_47939,N_47732,N_47724);
or U47940 (N_47940,N_47721,N_47682);
nand U47941 (N_47941,N_47676,N_47504);
nor U47942 (N_47942,N_47611,N_47539);
or U47943 (N_47943,N_47559,N_47560);
or U47944 (N_47944,N_47711,N_47546);
nand U47945 (N_47945,N_47682,N_47638);
nor U47946 (N_47946,N_47569,N_47702);
and U47947 (N_47947,N_47551,N_47575);
or U47948 (N_47948,N_47578,N_47637);
nand U47949 (N_47949,N_47711,N_47562);
nor U47950 (N_47950,N_47678,N_47565);
nand U47951 (N_47951,N_47544,N_47734);
xor U47952 (N_47952,N_47682,N_47632);
or U47953 (N_47953,N_47667,N_47589);
or U47954 (N_47954,N_47663,N_47603);
or U47955 (N_47955,N_47688,N_47561);
xnor U47956 (N_47956,N_47671,N_47659);
and U47957 (N_47957,N_47511,N_47671);
nand U47958 (N_47958,N_47676,N_47633);
xor U47959 (N_47959,N_47565,N_47515);
and U47960 (N_47960,N_47583,N_47635);
xnor U47961 (N_47961,N_47546,N_47702);
xor U47962 (N_47962,N_47748,N_47733);
nor U47963 (N_47963,N_47656,N_47512);
nor U47964 (N_47964,N_47671,N_47698);
xnor U47965 (N_47965,N_47749,N_47508);
nand U47966 (N_47966,N_47673,N_47629);
nand U47967 (N_47967,N_47658,N_47657);
xnor U47968 (N_47968,N_47605,N_47629);
or U47969 (N_47969,N_47624,N_47646);
and U47970 (N_47970,N_47724,N_47744);
and U47971 (N_47971,N_47709,N_47677);
xnor U47972 (N_47972,N_47704,N_47523);
or U47973 (N_47973,N_47525,N_47606);
nand U47974 (N_47974,N_47664,N_47731);
xnor U47975 (N_47975,N_47744,N_47656);
xor U47976 (N_47976,N_47638,N_47738);
nand U47977 (N_47977,N_47642,N_47709);
and U47978 (N_47978,N_47520,N_47705);
nor U47979 (N_47979,N_47588,N_47595);
and U47980 (N_47980,N_47524,N_47553);
nor U47981 (N_47981,N_47679,N_47604);
or U47982 (N_47982,N_47686,N_47517);
nand U47983 (N_47983,N_47629,N_47506);
xnor U47984 (N_47984,N_47585,N_47610);
nor U47985 (N_47985,N_47596,N_47675);
xnor U47986 (N_47986,N_47573,N_47530);
xnor U47987 (N_47987,N_47649,N_47702);
xnor U47988 (N_47988,N_47517,N_47658);
nand U47989 (N_47989,N_47534,N_47731);
or U47990 (N_47990,N_47611,N_47584);
nand U47991 (N_47991,N_47732,N_47614);
and U47992 (N_47992,N_47599,N_47639);
or U47993 (N_47993,N_47503,N_47621);
and U47994 (N_47994,N_47696,N_47517);
nor U47995 (N_47995,N_47572,N_47534);
and U47996 (N_47996,N_47719,N_47691);
nand U47997 (N_47997,N_47581,N_47592);
or U47998 (N_47998,N_47709,N_47648);
nand U47999 (N_47999,N_47718,N_47739);
xor U48000 (N_48000,N_47908,N_47790);
nor U48001 (N_48001,N_47989,N_47956);
and U48002 (N_48002,N_47944,N_47837);
nand U48003 (N_48003,N_47853,N_47888);
nor U48004 (N_48004,N_47983,N_47965);
or U48005 (N_48005,N_47771,N_47777);
nor U48006 (N_48006,N_47914,N_47834);
and U48007 (N_48007,N_47843,N_47906);
or U48008 (N_48008,N_47907,N_47946);
xor U48009 (N_48009,N_47864,N_47788);
and U48010 (N_48010,N_47930,N_47887);
nand U48011 (N_48011,N_47880,N_47991);
and U48012 (N_48012,N_47918,N_47851);
nand U48013 (N_48013,N_47941,N_47860);
nor U48014 (N_48014,N_47943,N_47804);
nand U48015 (N_48015,N_47940,N_47855);
nor U48016 (N_48016,N_47839,N_47937);
or U48017 (N_48017,N_47847,N_47993);
nand U48018 (N_48018,N_47976,N_47877);
nand U48019 (N_48019,N_47767,N_47927);
or U48020 (N_48020,N_47850,N_47751);
and U48021 (N_48021,N_47878,N_47848);
xnor U48022 (N_48022,N_47960,N_47897);
nand U48023 (N_48023,N_47821,N_47998);
nor U48024 (N_48024,N_47879,N_47799);
xnor U48025 (N_48025,N_47832,N_47859);
or U48026 (N_48026,N_47763,N_47892);
nand U48027 (N_48027,N_47792,N_47980);
nor U48028 (N_48028,N_47978,N_47840);
xnor U48029 (N_48029,N_47948,N_47866);
nor U48030 (N_48030,N_47870,N_47903);
and U48031 (N_48031,N_47768,N_47916);
nand U48032 (N_48032,N_47939,N_47802);
nand U48033 (N_48033,N_47961,N_47753);
and U48034 (N_48034,N_47896,N_47997);
and U48035 (N_48035,N_47833,N_47827);
and U48036 (N_48036,N_47762,N_47935);
or U48037 (N_48037,N_47809,N_47836);
or U48038 (N_48038,N_47829,N_47760);
nor U48039 (N_48039,N_47926,N_47779);
nand U48040 (N_48040,N_47787,N_47830);
and U48041 (N_48041,N_47780,N_47953);
and U48042 (N_48042,N_47871,N_47808);
xor U48043 (N_48043,N_47820,N_47924);
nand U48044 (N_48044,N_47894,N_47919);
and U48045 (N_48045,N_47922,N_47968);
and U48046 (N_48046,N_47890,N_47963);
nand U48047 (N_48047,N_47936,N_47959);
nand U48048 (N_48048,N_47984,N_47752);
xor U48049 (N_48049,N_47945,N_47795);
nor U48050 (N_48050,N_47899,N_47862);
nor U48051 (N_48051,N_47964,N_47754);
and U48052 (N_48052,N_47947,N_47774);
or U48053 (N_48053,N_47800,N_47981);
or U48054 (N_48054,N_47805,N_47987);
xnor U48055 (N_48055,N_47759,N_47882);
xor U48056 (N_48056,N_47967,N_47816);
xnor U48057 (N_48057,N_47949,N_47868);
nor U48058 (N_48058,N_47917,N_47942);
nand U48059 (N_48059,N_47958,N_47758);
xnor U48060 (N_48060,N_47846,N_47814);
nand U48061 (N_48061,N_47867,N_47962);
nor U48062 (N_48062,N_47818,N_47841);
nor U48063 (N_48063,N_47791,N_47977);
nor U48064 (N_48064,N_47782,N_47769);
xor U48065 (N_48065,N_47986,N_47785);
xor U48066 (N_48066,N_47902,N_47770);
nand U48067 (N_48067,N_47921,N_47889);
xnor U48068 (N_48068,N_47773,N_47822);
nand U48069 (N_48069,N_47844,N_47985);
or U48070 (N_48070,N_47973,N_47898);
xnor U48071 (N_48071,N_47934,N_47845);
xnor U48072 (N_48072,N_47856,N_47825);
nor U48073 (N_48073,N_47778,N_47975);
and U48074 (N_48074,N_47781,N_47798);
or U48075 (N_48075,N_47951,N_47789);
xnor U48076 (N_48076,N_47863,N_47994);
nor U48077 (N_48077,N_47910,N_47835);
xnor U48078 (N_48078,N_47786,N_47776);
nand U48079 (N_48079,N_47920,N_47842);
xnor U48080 (N_48080,N_47900,N_47905);
or U48081 (N_48081,N_47904,N_47955);
or U48082 (N_48082,N_47952,N_47988);
xnor U48083 (N_48083,N_47857,N_47971);
nor U48084 (N_48084,N_47876,N_47815);
nand U48085 (N_48085,N_47849,N_47972);
nor U48086 (N_48086,N_47757,N_47838);
nor U48087 (N_48087,N_47923,N_47932);
nand U48088 (N_48088,N_47756,N_47806);
nor U48089 (N_48089,N_47858,N_47893);
and U48090 (N_48090,N_47891,N_47982);
and U48091 (N_48091,N_47761,N_47999);
and U48092 (N_48092,N_47796,N_47823);
and U48093 (N_48093,N_47938,N_47974);
xnor U48094 (N_48094,N_47831,N_47797);
nand U48095 (N_48095,N_47807,N_47915);
or U48096 (N_48096,N_47824,N_47764);
nor U48097 (N_48097,N_47928,N_47957);
nor U48098 (N_48098,N_47813,N_47954);
nor U48099 (N_48099,N_47755,N_47881);
nor U48100 (N_48100,N_47784,N_47925);
or U48101 (N_48101,N_47828,N_47826);
or U48102 (N_48102,N_47995,N_47811);
and U48103 (N_48103,N_47884,N_47979);
nor U48104 (N_48104,N_47909,N_47819);
nor U48105 (N_48105,N_47990,N_47801);
or U48106 (N_48106,N_47873,N_47794);
xnor U48107 (N_48107,N_47883,N_47901);
nor U48108 (N_48108,N_47886,N_47861);
nor U48109 (N_48109,N_47874,N_47854);
xnor U48110 (N_48110,N_47812,N_47913);
and U48111 (N_48111,N_47852,N_47803);
xor U48112 (N_48112,N_47929,N_47969);
nand U48113 (N_48113,N_47992,N_47885);
nor U48114 (N_48114,N_47865,N_47931);
xnor U48115 (N_48115,N_47912,N_47772);
nand U48116 (N_48116,N_47872,N_47775);
or U48117 (N_48117,N_47875,N_47765);
nand U48118 (N_48118,N_47810,N_47783);
xnor U48119 (N_48119,N_47950,N_47869);
nor U48120 (N_48120,N_47895,N_47933);
xor U48121 (N_48121,N_47750,N_47970);
and U48122 (N_48122,N_47996,N_47766);
and U48123 (N_48123,N_47793,N_47911);
nand U48124 (N_48124,N_47966,N_47817);
and U48125 (N_48125,N_47860,N_47867);
nor U48126 (N_48126,N_47767,N_47901);
nand U48127 (N_48127,N_47763,N_47817);
nor U48128 (N_48128,N_47958,N_47839);
or U48129 (N_48129,N_47927,N_47769);
nor U48130 (N_48130,N_47817,N_47825);
and U48131 (N_48131,N_47836,N_47966);
nand U48132 (N_48132,N_47801,N_47767);
nor U48133 (N_48133,N_47808,N_47909);
nand U48134 (N_48134,N_47905,N_47782);
xnor U48135 (N_48135,N_47842,N_47960);
or U48136 (N_48136,N_47961,N_47842);
xnor U48137 (N_48137,N_47981,N_47945);
xor U48138 (N_48138,N_47753,N_47920);
nand U48139 (N_48139,N_47785,N_47893);
nand U48140 (N_48140,N_47822,N_47957);
nor U48141 (N_48141,N_47992,N_47905);
nor U48142 (N_48142,N_47992,N_47787);
xnor U48143 (N_48143,N_47957,N_47867);
and U48144 (N_48144,N_47774,N_47822);
nor U48145 (N_48145,N_47884,N_47974);
nand U48146 (N_48146,N_47812,N_47800);
nand U48147 (N_48147,N_47839,N_47860);
nor U48148 (N_48148,N_47774,N_47815);
xor U48149 (N_48149,N_47817,N_47904);
nand U48150 (N_48150,N_47810,N_47983);
or U48151 (N_48151,N_47797,N_47931);
nor U48152 (N_48152,N_47753,N_47785);
nor U48153 (N_48153,N_47912,N_47843);
nand U48154 (N_48154,N_47852,N_47856);
or U48155 (N_48155,N_47874,N_47863);
nor U48156 (N_48156,N_47970,N_47949);
nor U48157 (N_48157,N_47953,N_47765);
xor U48158 (N_48158,N_47793,N_47888);
nand U48159 (N_48159,N_47958,N_47862);
and U48160 (N_48160,N_47844,N_47787);
xnor U48161 (N_48161,N_47912,N_47914);
or U48162 (N_48162,N_47869,N_47865);
nand U48163 (N_48163,N_47952,N_47876);
xor U48164 (N_48164,N_47844,N_47947);
xnor U48165 (N_48165,N_47869,N_47888);
and U48166 (N_48166,N_47847,N_47912);
or U48167 (N_48167,N_47764,N_47813);
nand U48168 (N_48168,N_47767,N_47761);
and U48169 (N_48169,N_47785,N_47916);
nand U48170 (N_48170,N_47818,N_47803);
nor U48171 (N_48171,N_47816,N_47784);
and U48172 (N_48172,N_47871,N_47877);
xnor U48173 (N_48173,N_47850,N_47777);
and U48174 (N_48174,N_47862,N_47755);
nor U48175 (N_48175,N_47787,N_47952);
xnor U48176 (N_48176,N_47972,N_47753);
nand U48177 (N_48177,N_47931,N_47930);
nor U48178 (N_48178,N_47954,N_47843);
nor U48179 (N_48179,N_47949,N_47858);
xor U48180 (N_48180,N_47894,N_47769);
or U48181 (N_48181,N_47882,N_47932);
or U48182 (N_48182,N_47948,N_47933);
and U48183 (N_48183,N_47981,N_47793);
xnor U48184 (N_48184,N_47841,N_47858);
nand U48185 (N_48185,N_47777,N_47781);
xor U48186 (N_48186,N_47891,N_47871);
and U48187 (N_48187,N_47847,N_47842);
nand U48188 (N_48188,N_47778,N_47990);
nor U48189 (N_48189,N_47753,N_47923);
nor U48190 (N_48190,N_47786,N_47935);
nor U48191 (N_48191,N_47869,N_47976);
and U48192 (N_48192,N_47949,N_47835);
xor U48193 (N_48193,N_47978,N_47887);
xnor U48194 (N_48194,N_47958,N_47876);
xnor U48195 (N_48195,N_47814,N_47904);
or U48196 (N_48196,N_47777,N_47763);
nand U48197 (N_48197,N_47890,N_47764);
or U48198 (N_48198,N_47917,N_47957);
xnor U48199 (N_48199,N_47812,N_47921);
nor U48200 (N_48200,N_47837,N_47777);
and U48201 (N_48201,N_47822,N_47996);
xor U48202 (N_48202,N_47833,N_47878);
or U48203 (N_48203,N_47770,N_47909);
nor U48204 (N_48204,N_47759,N_47972);
nand U48205 (N_48205,N_47792,N_47942);
xor U48206 (N_48206,N_47833,N_47984);
nand U48207 (N_48207,N_47764,N_47918);
or U48208 (N_48208,N_47811,N_47822);
nor U48209 (N_48209,N_47986,N_47847);
and U48210 (N_48210,N_47882,N_47877);
xor U48211 (N_48211,N_47999,N_47863);
or U48212 (N_48212,N_47900,N_47887);
or U48213 (N_48213,N_47850,N_47809);
nor U48214 (N_48214,N_47768,N_47978);
and U48215 (N_48215,N_47781,N_47766);
xor U48216 (N_48216,N_47755,N_47768);
nand U48217 (N_48217,N_47807,N_47792);
xor U48218 (N_48218,N_47990,N_47810);
xnor U48219 (N_48219,N_47903,N_47937);
xor U48220 (N_48220,N_47889,N_47909);
nand U48221 (N_48221,N_47787,N_47980);
and U48222 (N_48222,N_47951,N_47764);
nand U48223 (N_48223,N_47767,N_47759);
or U48224 (N_48224,N_47963,N_47812);
nand U48225 (N_48225,N_47766,N_47956);
and U48226 (N_48226,N_47960,N_47878);
xor U48227 (N_48227,N_47760,N_47947);
xnor U48228 (N_48228,N_47863,N_47820);
and U48229 (N_48229,N_47901,N_47831);
nor U48230 (N_48230,N_47980,N_47941);
or U48231 (N_48231,N_47897,N_47752);
nand U48232 (N_48232,N_47852,N_47939);
nand U48233 (N_48233,N_47761,N_47910);
or U48234 (N_48234,N_47820,N_47903);
and U48235 (N_48235,N_47929,N_47856);
nand U48236 (N_48236,N_47765,N_47913);
and U48237 (N_48237,N_47779,N_47953);
or U48238 (N_48238,N_47781,N_47883);
and U48239 (N_48239,N_47832,N_47879);
or U48240 (N_48240,N_47850,N_47831);
xnor U48241 (N_48241,N_47846,N_47943);
xor U48242 (N_48242,N_47869,N_47785);
and U48243 (N_48243,N_47830,N_47898);
or U48244 (N_48244,N_47807,N_47779);
and U48245 (N_48245,N_47776,N_47872);
or U48246 (N_48246,N_47879,N_47780);
nand U48247 (N_48247,N_47967,N_47944);
nor U48248 (N_48248,N_47932,N_47884);
xor U48249 (N_48249,N_47943,N_47934);
nor U48250 (N_48250,N_48233,N_48121);
or U48251 (N_48251,N_48157,N_48087);
nand U48252 (N_48252,N_48000,N_48062);
or U48253 (N_48253,N_48145,N_48249);
or U48254 (N_48254,N_48015,N_48107);
or U48255 (N_48255,N_48147,N_48020);
xnor U48256 (N_48256,N_48216,N_48092);
or U48257 (N_48257,N_48063,N_48106);
nand U48258 (N_48258,N_48054,N_48070);
nor U48259 (N_48259,N_48030,N_48114);
xnor U48260 (N_48260,N_48071,N_48003);
nor U48261 (N_48261,N_48048,N_48109);
nor U48262 (N_48262,N_48153,N_48139);
or U48263 (N_48263,N_48187,N_48001);
nor U48264 (N_48264,N_48060,N_48064);
xor U48265 (N_48265,N_48206,N_48156);
nor U48266 (N_48266,N_48201,N_48133);
and U48267 (N_48267,N_48155,N_48078);
xnor U48268 (N_48268,N_48152,N_48095);
nand U48269 (N_48269,N_48053,N_48120);
and U48270 (N_48270,N_48150,N_48035);
nand U48271 (N_48271,N_48202,N_48119);
nor U48272 (N_48272,N_48058,N_48191);
or U48273 (N_48273,N_48105,N_48076);
nand U48274 (N_48274,N_48227,N_48246);
nand U48275 (N_48275,N_48019,N_48237);
xnor U48276 (N_48276,N_48032,N_48113);
or U48277 (N_48277,N_48200,N_48068);
or U48278 (N_48278,N_48196,N_48218);
nand U48279 (N_48279,N_48190,N_48103);
nor U48280 (N_48280,N_48044,N_48193);
and U48281 (N_48281,N_48189,N_48008);
nor U48282 (N_48282,N_48141,N_48043);
nand U48283 (N_48283,N_48110,N_48125);
or U48284 (N_48284,N_48031,N_48245);
nor U48285 (N_48285,N_48129,N_48226);
and U48286 (N_48286,N_48069,N_48134);
nand U48287 (N_48287,N_48209,N_48230);
or U48288 (N_48288,N_48163,N_48009);
or U48289 (N_48289,N_48046,N_48184);
nand U48290 (N_48290,N_48059,N_48143);
and U48291 (N_48291,N_48126,N_48234);
nor U48292 (N_48292,N_48111,N_48248);
nand U48293 (N_48293,N_48115,N_48166);
and U48294 (N_48294,N_48239,N_48128);
xnor U48295 (N_48295,N_48224,N_48136);
xnor U48296 (N_48296,N_48075,N_48005);
or U48297 (N_48297,N_48135,N_48217);
nor U48298 (N_48298,N_48082,N_48192);
xor U48299 (N_48299,N_48247,N_48148);
xor U48300 (N_48300,N_48029,N_48026);
or U48301 (N_48301,N_48175,N_48199);
and U48302 (N_48302,N_48102,N_48090);
xor U48303 (N_48303,N_48021,N_48203);
nand U48304 (N_48304,N_48149,N_48047);
or U48305 (N_48305,N_48146,N_48131);
xnor U48306 (N_48306,N_48231,N_48073);
or U48307 (N_48307,N_48004,N_48018);
nor U48308 (N_48308,N_48013,N_48137);
xor U48309 (N_48309,N_48142,N_48056);
or U48310 (N_48310,N_48243,N_48236);
xor U48311 (N_48311,N_48160,N_48240);
and U48312 (N_48312,N_48208,N_48241);
nor U48313 (N_48313,N_48101,N_48117);
nand U48314 (N_48314,N_48214,N_48138);
nand U48315 (N_48315,N_48232,N_48244);
xor U48316 (N_48316,N_48161,N_48023);
nand U48317 (N_48317,N_48219,N_48084);
xnor U48318 (N_48318,N_48154,N_48010);
nand U48319 (N_48319,N_48067,N_48172);
xnor U48320 (N_48320,N_48195,N_48089);
and U48321 (N_48321,N_48198,N_48006);
or U48322 (N_48322,N_48098,N_48097);
and U48323 (N_48323,N_48124,N_48204);
nor U48324 (N_48324,N_48027,N_48215);
nand U48325 (N_48325,N_48212,N_48140);
xor U48326 (N_48326,N_48151,N_48176);
and U48327 (N_48327,N_48037,N_48011);
xnor U48328 (N_48328,N_48038,N_48222);
or U48329 (N_48329,N_48179,N_48229);
xnor U48330 (N_48330,N_48221,N_48159);
or U48331 (N_48331,N_48235,N_48167);
and U48332 (N_48332,N_48158,N_48211);
and U48333 (N_48333,N_48042,N_48186);
nor U48334 (N_48334,N_48210,N_48130);
xnor U48335 (N_48335,N_48091,N_48132);
or U48336 (N_48336,N_48127,N_48116);
or U48337 (N_48337,N_48197,N_48170);
nand U48338 (N_48338,N_48036,N_48242);
nor U48339 (N_48339,N_48178,N_48207);
and U48340 (N_48340,N_48177,N_48066);
and U48341 (N_48341,N_48182,N_48213);
nor U48342 (N_48342,N_48165,N_48088);
or U48343 (N_48343,N_48220,N_48086);
nand U48344 (N_48344,N_48238,N_48017);
and U48345 (N_48345,N_48122,N_48083);
and U48346 (N_48346,N_48079,N_48024);
or U48347 (N_48347,N_48016,N_48168);
and U48348 (N_48348,N_48169,N_48012);
nor U48349 (N_48349,N_48057,N_48225);
nor U48350 (N_48350,N_48223,N_48055);
nand U48351 (N_48351,N_48144,N_48180);
nand U48352 (N_48352,N_48096,N_48002);
or U48353 (N_48353,N_48014,N_48034);
or U48354 (N_48354,N_48052,N_48123);
and U48355 (N_48355,N_48185,N_48173);
or U48356 (N_48356,N_48028,N_48162);
or U48357 (N_48357,N_48074,N_48045);
nor U48358 (N_48358,N_48072,N_48093);
nand U48359 (N_48359,N_48171,N_48183);
or U48360 (N_48360,N_48061,N_48051);
xor U48361 (N_48361,N_48099,N_48100);
nor U48362 (N_48362,N_48025,N_48118);
nor U48363 (N_48363,N_48039,N_48041);
xnor U48364 (N_48364,N_48194,N_48188);
nand U48365 (N_48365,N_48108,N_48104);
or U48366 (N_48366,N_48049,N_48080);
nand U48367 (N_48367,N_48040,N_48085);
nand U48368 (N_48368,N_48065,N_48077);
nor U48369 (N_48369,N_48164,N_48112);
nor U48370 (N_48370,N_48181,N_48094);
and U48371 (N_48371,N_48033,N_48050);
or U48372 (N_48372,N_48081,N_48174);
and U48373 (N_48373,N_48205,N_48007);
xnor U48374 (N_48374,N_48022,N_48228);
nor U48375 (N_48375,N_48228,N_48068);
or U48376 (N_48376,N_48150,N_48072);
and U48377 (N_48377,N_48151,N_48011);
nand U48378 (N_48378,N_48209,N_48046);
and U48379 (N_48379,N_48011,N_48104);
nand U48380 (N_48380,N_48157,N_48015);
or U48381 (N_48381,N_48044,N_48245);
nand U48382 (N_48382,N_48231,N_48168);
or U48383 (N_48383,N_48181,N_48027);
xor U48384 (N_48384,N_48155,N_48142);
nand U48385 (N_48385,N_48190,N_48199);
and U48386 (N_48386,N_48039,N_48106);
and U48387 (N_48387,N_48006,N_48138);
and U48388 (N_48388,N_48170,N_48248);
and U48389 (N_48389,N_48086,N_48221);
xnor U48390 (N_48390,N_48142,N_48080);
or U48391 (N_48391,N_48082,N_48077);
and U48392 (N_48392,N_48097,N_48026);
or U48393 (N_48393,N_48155,N_48231);
and U48394 (N_48394,N_48140,N_48218);
xnor U48395 (N_48395,N_48176,N_48239);
xor U48396 (N_48396,N_48223,N_48016);
nand U48397 (N_48397,N_48226,N_48075);
nand U48398 (N_48398,N_48029,N_48084);
or U48399 (N_48399,N_48043,N_48223);
xnor U48400 (N_48400,N_48205,N_48123);
or U48401 (N_48401,N_48229,N_48237);
or U48402 (N_48402,N_48149,N_48142);
or U48403 (N_48403,N_48235,N_48084);
nand U48404 (N_48404,N_48045,N_48232);
nor U48405 (N_48405,N_48078,N_48240);
nor U48406 (N_48406,N_48058,N_48203);
xor U48407 (N_48407,N_48012,N_48077);
nor U48408 (N_48408,N_48071,N_48051);
xnor U48409 (N_48409,N_48238,N_48083);
and U48410 (N_48410,N_48063,N_48143);
xnor U48411 (N_48411,N_48095,N_48216);
and U48412 (N_48412,N_48166,N_48199);
and U48413 (N_48413,N_48067,N_48188);
nand U48414 (N_48414,N_48214,N_48074);
or U48415 (N_48415,N_48139,N_48092);
nor U48416 (N_48416,N_48069,N_48164);
or U48417 (N_48417,N_48186,N_48177);
xor U48418 (N_48418,N_48005,N_48229);
and U48419 (N_48419,N_48240,N_48227);
nor U48420 (N_48420,N_48128,N_48133);
nand U48421 (N_48421,N_48016,N_48054);
or U48422 (N_48422,N_48173,N_48029);
or U48423 (N_48423,N_48182,N_48052);
nand U48424 (N_48424,N_48046,N_48062);
or U48425 (N_48425,N_48087,N_48038);
nor U48426 (N_48426,N_48114,N_48084);
nor U48427 (N_48427,N_48058,N_48086);
nand U48428 (N_48428,N_48095,N_48243);
nand U48429 (N_48429,N_48186,N_48099);
nor U48430 (N_48430,N_48037,N_48082);
and U48431 (N_48431,N_48014,N_48002);
nand U48432 (N_48432,N_48092,N_48025);
nand U48433 (N_48433,N_48114,N_48018);
and U48434 (N_48434,N_48028,N_48080);
nand U48435 (N_48435,N_48103,N_48123);
and U48436 (N_48436,N_48070,N_48127);
xnor U48437 (N_48437,N_48009,N_48206);
nand U48438 (N_48438,N_48074,N_48034);
or U48439 (N_48439,N_48218,N_48207);
or U48440 (N_48440,N_48237,N_48214);
nand U48441 (N_48441,N_48224,N_48078);
and U48442 (N_48442,N_48155,N_48114);
nor U48443 (N_48443,N_48138,N_48199);
and U48444 (N_48444,N_48081,N_48090);
or U48445 (N_48445,N_48095,N_48082);
and U48446 (N_48446,N_48087,N_48166);
and U48447 (N_48447,N_48038,N_48246);
or U48448 (N_48448,N_48129,N_48060);
or U48449 (N_48449,N_48129,N_48039);
nand U48450 (N_48450,N_48207,N_48094);
nand U48451 (N_48451,N_48132,N_48155);
or U48452 (N_48452,N_48230,N_48164);
or U48453 (N_48453,N_48222,N_48121);
nor U48454 (N_48454,N_48073,N_48099);
nor U48455 (N_48455,N_48014,N_48244);
and U48456 (N_48456,N_48103,N_48176);
or U48457 (N_48457,N_48190,N_48032);
nor U48458 (N_48458,N_48069,N_48191);
xor U48459 (N_48459,N_48184,N_48185);
and U48460 (N_48460,N_48016,N_48125);
nor U48461 (N_48461,N_48127,N_48247);
or U48462 (N_48462,N_48088,N_48134);
nor U48463 (N_48463,N_48077,N_48042);
nor U48464 (N_48464,N_48066,N_48181);
nor U48465 (N_48465,N_48108,N_48089);
nand U48466 (N_48466,N_48000,N_48126);
or U48467 (N_48467,N_48110,N_48192);
and U48468 (N_48468,N_48115,N_48207);
nor U48469 (N_48469,N_48244,N_48007);
xnor U48470 (N_48470,N_48066,N_48137);
and U48471 (N_48471,N_48160,N_48068);
and U48472 (N_48472,N_48124,N_48133);
nand U48473 (N_48473,N_48142,N_48032);
nand U48474 (N_48474,N_48180,N_48115);
nor U48475 (N_48475,N_48069,N_48004);
nand U48476 (N_48476,N_48018,N_48232);
nand U48477 (N_48477,N_48043,N_48233);
nor U48478 (N_48478,N_48215,N_48247);
or U48479 (N_48479,N_48200,N_48067);
xor U48480 (N_48480,N_48219,N_48176);
nand U48481 (N_48481,N_48130,N_48058);
and U48482 (N_48482,N_48029,N_48088);
xor U48483 (N_48483,N_48018,N_48227);
xor U48484 (N_48484,N_48091,N_48076);
nor U48485 (N_48485,N_48147,N_48213);
nand U48486 (N_48486,N_48218,N_48212);
and U48487 (N_48487,N_48175,N_48141);
nand U48488 (N_48488,N_48109,N_48238);
or U48489 (N_48489,N_48176,N_48216);
or U48490 (N_48490,N_48178,N_48019);
and U48491 (N_48491,N_48057,N_48054);
or U48492 (N_48492,N_48227,N_48237);
nor U48493 (N_48493,N_48105,N_48238);
xor U48494 (N_48494,N_48139,N_48112);
nor U48495 (N_48495,N_48105,N_48191);
xnor U48496 (N_48496,N_48174,N_48054);
and U48497 (N_48497,N_48033,N_48119);
nor U48498 (N_48498,N_48116,N_48089);
or U48499 (N_48499,N_48052,N_48176);
and U48500 (N_48500,N_48495,N_48447);
xnor U48501 (N_48501,N_48271,N_48469);
nor U48502 (N_48502,N_48409,N_48301);
nor U48503 (N_48503,N_48470,N_48287);
nand U48504 (N_48504,N_48496,N_48385);
xnor U48505 (N_48505,N_48492,N_48386);
and U48506 (N_48506,N_48452,N_48480);
nor U48507 (N_48507,N_48479,N_48449);
nand U48508 (N_48508,N_48493,N_48277);
nor U48509 (N_48509,N_48347,N_48485);
xnor U48510 (N_48510,N_48466,N_48405);
nand U48511 (N_48511,N_48323,N_48491);
or U48512 (N_48512,N_48355,N_48286);
or U48513 (N_48513,N_48454,N_48423);
nand U48514 (N_48514,N_48362,N_48354);
and U48515 (N_48515,N_48293,N_48372);
xor U48516 (N_48516,N_48300,N_48445);
xor U48517 (N_48517,N_48285,N_48461);
and U48518 (N_48518,N_48269,N_48291);
xor U48519 (N_48519,N_48371,N_48426);
and U48520 (N_48520,N_48476,N_48446);
nor U48521 (N_48521,N_48280,N_48383);
nand U48522 (N_48522,N_48278,N_48375);
or U48523 (N_48523,N_48391,N_48365);
and U48524 (N_48524,N_48296,N_48295);
nand U48525 (N_48525,N_48350,N_48417);
and U48526 (N_48526,N_48361,N_48394);
xor U48527 (N_48527,N_48482,N_48341);
xor U48528 (N_48528,N_48335,N_48315);
and U48529 (N_48529,N_48471,N_48458);
nor U48530 (N_48530,N_48332,N_48265);
xnor U48531 (N_48531,N_48404,N_48419);
nand U48532 (N_48532,N_48322,N_48377);
or U48533 (N_48533,N_48264,N_48415);
and U48534 (N_48534,N_48463,N_48348);
and U48535 (N_48535,N_48465,N_48418);
nor U48536 (N_48536,N_48364,N_48321);
or U48537 (N_48537,N_48282,N_48252);
xor U48538 (N_48538,N_48421,N_48268);
or U48539 (N_48539,N_48381,N_48483);
nand U48540 (N_48540,N_48329,N_48333);
nand U48541 (N_48541,N_48408,N_48369);
nor U48542 (N_48542,N_48360,N_48378);
xnor U48543 (N_48543,N_48498,N_48254);
xnor U48544 (N_48544,N_48260,N_48494);
nand U48545 (N_48545,N_48473,N_48308);
and U48546 (N_48546,N_48303,N_48297);
nor U48547 (N_48547,N_48464,N_48393);
xnor U48548 (N_48548,N_48433,N_48319);
xor U48549 (N_48549,N_48317,N_48487);
nand U48550 (N_48550,N_48429,N_48441);
or U48551 (N_48551,N_48331,N_48478);
nand U48552 (N_48552,N_48437,N_48425);
xnor U48553 (N_48553,N_48486,N_48435);
xnor U48554 (N_48554,N_48316,N_48422);
nor U48555 (N_48555,N_48451,N_48339);
and U48556 (N_48556,N_48304,N_48373);
nor U48557 (N_48557,N_48274,N_48424);
or U48558 (N_48558,N_48399,N_48336);
xor U48559 (N_48559,N_48258,N_48266);
nor U48560 (N_48560,N_48413,N_48284);
nor U48561 (N_48561,N_48376,N_48453);
nor U48562 (N_48562,N_48481,N_48416);
and U48563 (N_48563,N_48477,N_48324);
and U48564 (N_48564,N_48434,N_48427);
and U48565 (N_48565,N_48387,N_48338);
or U48566 (N_48566,N_48411,N_48379);
xnor U48567 (N_48567,N_48459,N_48292);
xnor U48568 (N_48568,N_48294,N_48251);
and U48569 (N_48569,N_48281,N_48356);
xnor U48570 (N_48570,N_48389,N_48275);
or U48571 (N_48571,N_48259,N_48272);
and U48572 (N_48572,N_48309,N_48267);
or U48573 (N_48573,N_48306,N_48402);
or U48574 (N_48574,N_48397,N_48443);
nand U48575 (N_48575,N_48276,N_48310);
and U48576 (N_48576,N_48450,N_48438);
nand U48577 (N_48577,N_48368,N_48359);
or U48578 (N_48578,N_48357,N_48302);
xnor U48579 (N_48579,N_48442,N_48327);
or U48580 (N_48580,N_48484,N_48499);
or U48581 (N_48581,N_48337,N_48314);
and U48582 (N_48582,N_48346,N_48468);
xor U48583 (N_48583,N_48407,N_48288);
and U48584 (N_48584,N_48255,N_48395);
nand U48585 (N_48585,N_48340,N_48444);
xor U48586 (N_48586,N_48401,N_48334);
nor U48587 (N_48587,N_48250,N_48392);
or U48588 (N_48588,N_48488,N_48351);
xnor U48589 (N_48589,N_48455,N_48342);
nor U48590 (N_48590,N_48330,N_48358);
and U48591 (N_48591,N_48253,N_48256);
nor U48592 (N_48592,N_48343,N_48380);
nor U48593 (N_48593,N_48313,N_48403);
xor U48594 (N_48594,N_48431,N_48257);
nor U48595 (N_48595,N_48345,N_48439);
xnor U48596 (N_48596,N_48352,N_48382);
xor U48597 (N_48597,N_48318,N_48305);
nand U48598 (N_48598,N_48279,N_48262);
nand U48599 (N_48599,N_48270,N_48326);
nor U48600 (N_48600,N_48430,N_48436);
and U48601 (N_48601,N_48363,N_48497);
and U48602 (N_48602,N_48344,N_48420);
nor U48603 (N_48603,N_48474,N_48261);
nand U48604 (N_48604,N_48320,N_48388);
and U48605 (N_48605,N_48398,N_48367);
or U48606 (N_48606,N_48366,N_48307);
nand U48607 (N_48607,N_48428,N_48462);
xnor U48608 (N_48608,N_48312,N_48414);
nand U48609 (N_48609,N_48298,N_48406);
nor U48610 (N_48610,N_48456,N_48472);
and U48611 (N_48611,N_48325,N_48289);
or U48612 (N_48612,N_48432,N_48283);
and U48613 (N_48613,N_48396,N_48370);
nor U48614 (N_48614,N_48467,N_48353);
nand U48615 (N_48615,N_48412,N_48489);
nor U48616 (N_48616,N_48311,N_48349);
nand U48617 (N_48617,N_48440,N_48384);
nand U48618 (N_48618,N_48400,N_48263);
and U48619 (N_48619,N_48460,N_48290);
xor U48620 (N_48620,N_48328,N_48457);
xnor U48621 (N_48621,N_48475,N_48299);
nand U48622 (N_48622,N_48490,N_48448);
nand U48623 (N_48623,N_48390,N_48410);
nor U48624 (N_48624,N_48273,N_48374);
or U48625 (N_48625,N_48442,N_48331);
nor U48626 (N_48626,N_48338,N_48473);
or U48627 (N_48627,N_48273,N_48278);
or U48628 (N_48628,N_48307,N_48411);
nor U48629 (N_48629,N_48401,N_48393);
and U48630 (N_48630,N_48448,N_48355);
or U48631 (N_48631,N_48374,N_48354);
nand U48632 (N_48632,N_48278,N_48390);
nand U48633 (N_48633,N_48330,N_48272);
xor U48634 (N_48634,N_48347,N_48417);
nor U48635 (N_48635,N_48488,N_48493);
nand U48636 (N_48636,N_48390,N_48292);
nor U48637 (N_48637,N_48448,N_48478);
or U48638 (N_48638,N_48295,N_48341);
xor U48639 (N_48639,N_48464,N_48467);
nand U48640 (N_48640,N_48401,N_48394);
nand U48641 (N_48641,N_48294,N_48354);
and U48642 (N_48642,N_48291,N_48398);
nand U48643 (N_48643,N_48315,N_48324);
nand U48644 (N_48644,N_48316,N_48314);
nand U48645 (N_48645,N_48396,N_48373);
or U48646 (N_48646,N_48388,N_48483);
or U48647 (N_48647,N_48376,N_48358);
xnor U48648 (N_48648,N_48390,N_48378);
nor U48649 (N_48649,N_48257,N_48344);
or U48650 (N_48650,N_48452,N_48438);
xnor U48651 (N_48651,N_48286,N_48459);
nand U48652 (N_48652,N_48438,N_48433);
nand U48653 (N_48653,N_48415,N_48407);
nand U48654 (N_48654,N_48379,N_48326);
xor U48655 (N_48655,N_48491,N_48273);
nand U48656 (N_48656,N_48456,N_48317);
xor U48657 (N_48657,N_48388,N_48499);
nor U48658 (N_48658,N_48331,N_48423);
nor U48659 (N_48659,N_48381,N_48440);
and U48660 (N_48660,N_48475,N_48294);
nand U48661 (N_48661,N_48276,N_48271);
nand U48662 (N_48662,N_48464,N_48435);
xor U48663 (N_48663,N_48380,N_48376);
nand U48664 (N_48664,N_48385,N_48314);
or U48665 (N_48665,N_48472,N_48438);
nand U48666 (N_48666,N_48444,N_48416);
xor U48667 (N_48667,N_48367,N_48315);
nand U48668 (N_48668,N_48307,N_48315);
and U48669 (N_48669,N_48370,N_48474);
xor U48670 (N_48670,N_48474,N_48469);
nand U48671 (N_48671,N_48410,N_48251);
nand U48672 (N_48672,N_48298,N_48311);
xor U48673 (N_48673,N_48348,N_48289);
xnor U48674 (N_48674,N_48441,N_48381);
and U48675 (N_48675,N_48282,N_48298);
xnor U48676 (N_48676,N_48334,N_48350);
nand U48677 (N_48677,N_48284,N_48388);
nand U48678 (N_48678,N_48365,N_48312);
nor U48679 (N_48679,N_48368,N_48295);
or U48680 (N_48680,N_48374,N_48400);
xnor U48681 (N_48681,N_48477,N_48326);
xor U48682 (N_48682,N_48493,N_48337);
xnor U48683 (N_48683,N_48268,N_48283);
nor U48684 (N_48684,N_48473,N_48270);
nor U48685 (N_48685,N_48405,N_48337);
nand U48686 (N_48686,N_48378,N_48464);
or U48687 (N_48687,N_48264,N_48280);
and U48688 (N_48688,N_48325,N_48451);
nand U48689 (N_48689,N_48296,N_48477);
nor U48690 (N_48690,N_48321,N_48378);
or U48691 (N_48691,N_48379,N_48446);
nor U48692 (N_48692,N_48364,N_48425);
nor U48693 (N_48693,N_48491,N_48383);
nor U48694 (N_48694,N_48351,N_48446);
and U48695 (N_48695,N_48412,N_48432);
or U48696 (N_48696,N_48432,N_48281);
nand U48697 (N_48697,N_48427,N_48357);
nand U48698 (N_48698,N_48366,N_48351);
xor U48699 (N_48699,N_48333,N_48417);
nand U48700 (N_48700,N_48408,N_48284);
nor U48701 (N_48701,N_48439,N_48275);
xnor U48702 (N_48702,N_48450,N_48337);
nand U48703 (N_48703,N_48319,N_48480);
nor U48704 (N_48704,N_48426,N_48308);
and U48705 (N_48705,N_48340,N_48497);
nand U48706 (N_48706,N_48408,N_48497);
and U48707 (N_48707,N_48340,N_48314);
nand U48708 (N_48708,N_48470,N_48400);
xor U48709 (N_48709,N_48496,N_48266);
xnor U48710 (N_48710,N_48420,N_48288);
nor U48711 (N_48711,N_48315,N_48391);
and U48712 (N_48712,N_48383,N_48388);
nand U48713 (N_48713,N_48431,N_48291);
xor U48714 (N_48714,N_48322,N_48450);
and U48715 (N_48715,N_48393,N_48266);
nand U48716 (N_48716,N_48308,N_48443);
nor U48717 (N_48717,N_48337,N_48308);
nor U48718 (N_48718,N_48347,N_48491);
nand U48719 (N_48719,N_48440,N_48374);
nor U48720 (N_48720,N_48290,N_48251);
and U48721 (N_48721,N_48490,N_48311);
and U48722 (N_48722,N_48369,N_48393);
or U48723 (N_48723,N_48286,N_48323);
xor U48724 (N_48724,N_48431,N_48270);
and U48725 (N_48725,N_48453,N_48366);
or U48726 (N_48726,N_48356,N_48306);
or U48727 (N_48727,N_48269,N_48298);
and U48728 (N_48728,N_48354,N_48479);
xnor U48729 (N_48729,N_48253,N_48420);
nor U48730 (N_48730,N_48395,N_48480);
nand U48731 (N_48731,N_48328,N_48269);
or U48732 (N_48732,N_48469,N_48276);
nand U48733 (N_48733,N_48443,N_48342);
nand U48734 (N_48734,N_48480,N_48424);
and U48735 (N_48735,N_48390,N_48301);
nor U48736 (N_48736,N_48277,N_48268);
nand U48737 (N_48737,N_48344,N_48452);
and U48738 (N_48738,N_48255,N_48354);
nor U48739 (N_48739,N_48416,N_48486);
nor U48740 (N_48740,N_48385,N_48293);
nor U48741 (N_48741,N_48270,N_48259);
and U48742 (N_48742,N_48413,N_48458);
xnor U48743 (N_48743,N_48279,N_48454);
or U48744 (N_48744,N_48439,N_48481);
nand U48745 (N_48745,N_48360,N_48450);
or U48746 (N_48746,N_48379,N_48294);
or U48747 (N_48747,N_48494,N_48382);
or U48748 (N_48748,N_48265,N_48303);
nor U48749 (N_48749,N_48331,N_48407);
xnor U48750 (N_48750,N_48661,N_48720);
or U48751 (N_48751,N_48572,N_48636);
nor U48752 (N_48752,N_48587,N_48585);
nor U48753 (N_48753,N_48677,N_48660);
nand U48754 (N_48754,N_48546,N_48675);
and U48755 (N_48755,N_48698,N_48715);
nand U48756 (N_48756,N_48673,N_48598);
xnor U48757 (N_48757,N_48566,N_48601);
nand U48758 (N_48758,N_48516,N_48716);
xnor U48759 (N_48759,N_48522,N_48699);
or U48760 (N_48760,N_48679,N_48500);
and U48761 (N_48761,N_48504,N_48681);
nor U48762 (N_48762,N_48569,N_48696);
xnor U48763 (N_48763,N_48735,N_48605);
xor U48764 (N_48764,N_48653,N_48651);
or U48765 (N_48765,N_48537,N_48656);
or U48766 (N_48766,N_48742,N_48567);
xnor U48767 (N_48767,N_48731,N_48544);
or U48768 (N_48768,N_48640,N_48525);
nor U48769 (N_48769,N_48671,N_48648);
xnor U48770 (N_48770,N_48719,N_48524);
or U48771 (N_48771,N_48508,N_48513);
xor U48772 (N_48772,N_48509,N_48562);
nor U48773 (N_48773,N_48554,N_48702);
and U48774 (N_48774,N_48556,N_48520);
nor U48775 (N_48775,N_48692,N_48652);
nand U48776 (N_48776,N_48521,N_48723);
or U48777 (N_48777,N_48550,N_48725);
nand U48778 (N_48778,N_48705,N_48530);
or U48779 (N_48779,N_48614,N_48644);
nand U48780 (N_48780,N_48539,N_48597);
and U48781 (N_48781,N_48718,N_48734);
nand U48782 (N_48782,N_48529,N_48600);
xor U48783 (N_48783,N_48729,N_48627);
nor U48784 (N_48784,N_48740,N_48704);
and U48785 (N_48785,N_48526,N_48616);
nor U48786 (N_48786,N_48727,N_48642);
and U48787 (N_48787,N_48712,N_48606);
nand U48788 (N_48788,N_48535,N_48564);
and U48789 (N_48789,N_48639,N_48737);
xor U48790 (N_48790,N_48503,N_48749);
nand U48791 (N_48791,N_48728,N_48580);
xnor U48792 (N_48792,N_48528,N_48717);
xnor U48793 (N_48793,N_48560,N_48632);
xnor U48794 (N_48794,N_48573,N_48512);
xnor U48795 (N_48795,N_48577,N_48711);
xor U48796 (N_48796,N_48523,N_48726);
and U48797 (N_48797,N_48634,N_48730);
nor U48798 (N_48798,N_48738,N_48510);
or U48799 (N_48799,N_48533,N_48647);
nand U48800 (N_48800,N_48575,N_48625);
xor U48801 (N_48801,N_48739,N_48633);
and U48802 (N_48802,N_48558,N_48654);
or U48803 (N_48803,N_48590,N_48688);
nor U48804 (N_48804,N_48584,N_48743);
xnor U48805 (N_48805,N_48689,N_48682);
or U48806 (N_48806,N_48511,N_48736);
xnor U48807 (N_48807,N_48568,N_48687);
or U48808 (N_48808,N_48674,N_48592);
and U48809 (N_48809,N_48635,N_48507);
nor U48810 (N_48810,N_48609,N_48545);
or U48811 (N_48811,N_48534,N_48662);
and U48812 (N_48812,N_48666,N_48540);
or U48813 (N_48813,N_48667,N_48626);
nand U48814 (N_48814,N_48561,N_48747);
or U48815 (N_48815,N_48680,N_48571);
or U48816 (N_48816,N_48518,N_48678);
nand U48817 (N_48817,N_48536,N_48663);
and U48818 (N_48818,N_48672,N_48691);
nand U48819 (N_48819,N_48706,N_48620);
xor U48820 (N_48820,N_48732,N_48563);
nor U48821 (N_48821,N_48700,N_48552);
and U48822 (N_48822,N_48659,N_48686);
nand U48823 (N_48823,N_48543,N_48501);
xnor U48824 (N_48824,N_48593,N_48555);
xnor U48825 (N_48825,N_48655,N_48502);
nor U48826 (N_48826,N_48576,N_48570);
and U48827 (N_48827,N_48586,N_48701);
or U48828 (N_48828,N_48542,N_48608);
nor U48829 (N_48829,N_48559,N_48641);
and U48830 (N_48830,N_48714,N_48548);
and U48831 (N_48831,N_48591,N_48713);
or U48832 (N_48832,N_48746,N_48710);
xor U48833 (N_48833,N_48623,N_48578);
xnor U48834 (N_48834,N_48553,N_48541);
or U48835 (N_48835,N_48721,N_48517);
or U48836 (N_48836,N_48693,N_48612);
or U48837 (N_48837,N_48709,N_48733);
xor U48838 (N_48838,N_48684,N_48643);
or U48839 (N_48839,N_48551,N_48602);
nand U48840 (N_48840,N_48610,N_48624);
or U48841 (N_48841,N_48588,N_48613);
and U48842 (N_48842,N_48603,N_48589);
nand U48843 (N_48843,N_48621,N_48596);
nand U48844 (N_48844,N_48748,N_48676);
and U48845 (N_48845,N_48690,N_48724);
nand U48846 (N_48846,N_48611,N_48669);
xor U48847 (N_48847,N_48581,N_48683);
nor U48848 (N_48848,N_48565,N_48607);
xnor U48849 (N_48849,N_48583,N_48594);
and U48850 (N_48850,N_48628,N_48574);
nor U48851 (N_48851,N_48722,N_48599);
xor U48852 (N_48852,N_48506,N_48638);
nand U48853 (N_48853,N_48519,N_48645);
nand U48854 (N_48854,N_48579,N_48741);
and U48855 (N_48855,N_48618,N_48707);
nand U48856 (N_48856,N_48619,N_48665);
and U48857 (N_48857,N_48622,N_48527);
xnor U48858 (N_48858,N_48646,N_48617);
and U48859 (N_48859,N_48657,N_48538);
nand U48860 (N_48860,N_48557,N_48532);
nor U48861 (N_48861,N_48547,N_48595);
nor U48862 (N_48862,N_48631,N_48514);
and U48863 (N_48863,N_48531,N_48668);
xor U48864 (N_48864,N_48694,N_48685);
nor U48865 (N_48865,N_48615,N_48650);
and U48866 (N_48866,N_48664,N_48637);
or U48867 (N_48867,N_48649,N_48582);
or U48868 (N_48868,N_48670,N_48549);
and U48869 (N_48869,N_48658,N_48695);
or U48870 (N_48870,N_48697,N_48515);
or U48871 (N_48871,N_48629,N_48744);
xnor U48872 (N_48872,N_48604,N_48708);
xnor U48873 (N_48873,N_48505,N_48630);
and U48874 (N_48874,N_48703,N_48745);
nor U48875 (N_48875,N_48737,N_48550);
nand U48876 (N_48876,N_48664,N_48591);
and U48877 (N_48877,N_48696,N_48737);
xnor U48878 (N_48878,N_48504,N_48552);
xor U48879 (N_48879,N_48603,N_48566);
nand U48880 (N_48880,N_48656,N_48528);
nor U48881 (N_48881,N_48521,N_48702);
or U48882 (N_48882,N_48748,N_48550);
xor U48883 (N_48883,N_48670,N_48693);
and U48884 (N_48884,N_48586,N_48698);
nor U48885 (N_48885,N_48634,N_48655);
or U48886 (N_48886,N_48710,N_48533);
nand U48887 (N_48887,N_48687,N_48661);
nand U48888 (N_48888,N_48603,N_48561);
xor U48889 (N_48889,N_48701,N_48567);
nor U48890 (N_48890,N_48588,N_48570);
nor U48891 (N_48891,N_48536,N_48608);
xnor U48892 (N_48892,N_48588,N_48629);
nand U48893 (N_48893,N_48683,N_48675);
or U48894 (N_48894,N_48513,N_48544);
nor U48895 (N_48895,N_48631,N_48567);
xor U48896 (N_48896,N_48598,N_48695);
nand U48897 (N_48897,N_48703,N_48692);
and U48898 (N_48898,N_48545,N_48523);
nor U48899 (N_48899,N_48625,N_48697);
nand U48900 (N_48900,N_48680,N_48580);
nor U48901 (N_48901,N_48597,N_48512);
and U48902 (N_48902,N_48685,N_48524);
or U48903 (N_48903,N_48575,N_48573);
nand U48904 (N_48904,N_48526,N_48513);
nor U48905 (N_48905,N_48697,N_48672);
or U48906 (N_48906,N_48518,N_48572);
nand U48907 (N_48907,N_48639,N_48571);
or U48908 (N_48908,N_48659,N_48540);
and U48909 (N_48909,N_48527,N_48597);
xor U48910 (N_48910,N_48722,N_48698);
nor U48911 (N_48911,N_48678,N_48703);
nand U48912 (N_48912,N_48597,N_48566);
xnor U48913 (N_48913,N_48651,N_48674);
and U48914 (N_48914,N_48583,N_48655);
or U48915 (N_48915,N_48642,N_48725);
and U48916 (N_48916,N_48736,N_48651);
and U48917 (N_48917,N_48734,N_48516);
xor U48918 (N_48918,N_48627,N_48655);
and U48919 (N_48919,N_48597,N_48728);
nor U48920 (N_48920,N_48715,N_48508);
xnor U48921 (N_48921,N_48524,N_48748);
and U48922 (N_48922,N_48583,N_48656);
or U48923 (N_48923,N_48628,N_48693);
xnor U48924 (N_48924,N_48630,N_48679);
nor U48925 (N_48925,N_48638,N_48690);
nor U48926 (N_48926,N_48634,N_48710);
or U48927 (N_48927,N_48648,N_48726);
nor U48928 (N_48928,N_48595,N_48585);
or U48929 (N_48929,N_48637,N_48583);
nand U48930 (N_48930,N_48632,N_48686);
xor U48931 (N_48931,N_48565,N_48654);
nor U48932 (N_48932,N_48509,N_48572);
xor U48933 (N_48933,N_48697,N_48506);
or U48934 (N_48934,N_48685,N_48562);
nand U48935 (N_48935,N_48522,N_48732);
nor U48936 (N_48936,N_48525,N_48678);
xor U48937 (N_48937,N_48595,N_48542);
and U48938 (N_48938,N_48748,N_48572);
nand U48939 (N_48939,N_48558,N_48633);
nand U48940 (N_48940,N_48631,N_48646);
and U48941 (N_48941,N_48633,N_48718);
nand U48942 (N_48942,N_48665,N_48679);
and U48943 (N_48943,N_48553,N_48565);
nor U48944 (N_48944,N_48669,N_48698);
xnor U48945 (N_48945,N_48611,N_48589);
or U48946 (N_48946,N_48698,N_48530);
xnor U48947 (N_48947,N_48527,N_48730);
or U48948 (N_48948,N_48690,N_48665);
nor U48949 (N_48949,N_48722,N_48637);
xor U48950 (N_48950,N_48699,N_48505);
nand U48951 (N_48951,N_48520,N_48591);
nand U48952 (N_48952,N_48745,N_48657);
and U48953 (N_48953,N_48571,N_48739);
and U48954 (N_48954,N_48726,N_48642);
and U48955 (N_48955,N_48584,N_48516);
nor U48956 (N_48956,N_48528,N_48585);
or U48957 (N_48957,N_48688,N_48747);
nand U48958 (N_48958,N_48644,N_48553);
nand U48959 (N_48959,N_48628,N_48527);
or U48960 (N_48960,N_48619,N_48579);
nand U48961 (N_48961,N_48632,N_48615);
nand U48962 (N_48962,N_48569,N_48668);
nand U48963 (N_48963,N_48600,N_48591);
xor U48964 (N_48964,N_48609,N_48721);
or U48965 (N_48965,N_48520,N_48604);
xor U48966 (N_48966,N_48705,N_48689);
and U48967 (N_48967,N_48644,N_48679);
and U48968 (N_48968,N_48601,N_48669);
and U48969 (N_48969,N_48528,N_48653);
nand U48970 (N_48970,N_48718,N_48507);
nor U48971 (N_48971,N_48578,N_48747);
nor U48972 (N_48972,N_48510,N_48555);
nor U48973 (N_48973,N_48675,N_48509);
or U48974 (N_48974,N_48634,N_48583);
nand U48975 (N_48975,N_48683,N_48527);
nor U48976 (N_48976,N_48631,N_48536);
xnor U48977 (N_48977,N_48659,N_48647);
or U48978 (N_48978,N_48620,N_48736);
xnor U48979 (N_48979,N_48683,N_48587);
nor U48980 (N_48980,N_48643,N_48744);
and U48981 (N_48981,N_48649,N_48688);
or U48982 (N_48982,N_48719,N_48645);
and U48983 (N_48983,N_48642,N_48525);
and U48984 (N_48984,N_48679,N_48631);
or U48985 (N_48985,N_48623,N_48513);
nor U48986 (N_48986,N_48671,N_48557);
nor U48987 (N_48987,N_48550,N_48590);
nor U48988 (N_48988,N_48502,N_48536);
xnor U48989 (N_48989,N_48655,N_48578);
and U48990 (N_48990,N_48711,N_48540);
xnor U48991 (N_48991,N_48579,N_48661);
xnor U48992 (N_48992,N_48701,N_48684);
or U48993 (N_48993,N_48677,N_48612);
or U48994 (N_48994,N_48717,N_48643);
nand U48995 (N_48995,N_48604,N_48681);
nand U48996 (N_48996,N_48602,N_48614);
xor U48997 (N_48997,N_48597,N_48625);
nor U48998 (N_48998,N_48705,N_48745);
and U48999 (N_48999,N_48565,N_48712);
or U49000 (N_49000,N_48928,N_48857);
and U49001 (N_49001,N_48886,N_48752);
or U49002 (N_49002,N_48927,N_48971);
or U49003 (N_49003,N_48934,N_48755);
xnor U49004 (N_49004,N_48860,N_48826);
xnor U49005 (N_49005,N_48906,N_48781);
xor U49006 (N_49006,N_48929,N_48938);
and U49007 (N_49007,N_48972,N_48979);
nand U49008 (N_49008,N_48894,N_48890);
nand U49009 (N_49009,N_48837,N_48870);
and U49010 (N_49010,N_48863,N_48872);
or U49011 (N_49011,N_48947,N_48763);
or U49012 (N_49012,N_48829,N_48782);
nor U49013 (N_49013,N_48767,N_48759);
nand U49014 (N_49014,N_48962,N_48952);
or U49015 (N_49015,N_48789,N_48823);
nand U49016 (N_49016,N_48840,N_48815);
or U49017 (N_49017,N_48836,N_48808);
or U49018 (N_49018,N_48843,N_48998);
nand U49019 (N_49019,N_48999,N_48940);
xor U49020 (N_49020,N_48909,N_48758);
or U49021 (N_49021,N_48879,N_48768);
or U49022 (N_49022,N_48831,N_48992);
or U49023 (N_49023,N_48757,N_48834);
and U49024 (N_49024,N_48780,N_48858);
xnor U49025 (N_49025,N_48930,N_48916);
or U49026 (N_49026,N_48824,N_48984);
or U49027 (N_49027,N_48931,N_48803);
and U49028 (N_49028,N_48905,N_48822);
nor U49029 (N_49029,N_48765,N_48963);
nor U49030 (N_49030,N_48910,N_48898);
nand U49031 (N_49031,N_48787,N_48964);
and U49032 (N_49032,N_48871,N_48881);
nor U49033 (N_49033,N_48908,N_48957);
nand U49034 (N_49034,N_48853,N_48764);
nor U49035 (N_49035,N_48891,N_48946);
or U49036 (N_49036,N_48897,N_48776);
nor U49037 (N_49037,N_48887,N_48778);
or U49038 (N_49038,N_48986,N_48842);
xor U49039 (N_49039,N_48920,N_48989);
nand U49040 (N_49040,N_48949,N_48895);
and U49041 (N_49041,N_48786,N_48750);
and U49042 (N_49042,N_48922,N_48903);
xnor U49043 (N_49043,N_48771,N_48791);
xnor U49044 (N_49044,N_48914,N_48973);
and U49045 (N_49045,N_48939,N_48802);
xnor U49046 (N_49046,N_48885,N_48797);
nor U49047 (N_49047,N_48987,N_48864);
nor U49048 (N_49048,N_48976,N_48777);
nor U49049 (N_49049,N_48799,N_48805);
or U49050 (N_49050,N_48809,N_48875);
and U49051 (N_49051,N_48865,N_48884);
or U49052 (N_49052,N_48841,N_48762);
and U49053 (N_49053,N_48975,N_48814);
nand U49054 (N_49054,N_48811,N_48882);
and U49055 (N_49055,N_48852,N_48985);
or U49056 (N_49056,N_48937,N_48883);
or U49057 (N_49057,N_48775,N_48925);
nor U49058 (N_49058,N_48790,N_48854);
nand U49059 (N_49059,N_48825,N_48868);
nor U49060 (N_49060,N_48779,N_48848);
nand U49061 (N_49061,N_48954,N_48965);
xnor U49062 (N_49062,N_48935,N_48761);
and U49063 (N_49063,N_48953,N_48770);
and U49064 (N_49064,N_48867,N_48774);
or U49065 (N_49065,N_48974,N_48798);
xor U49066 (N_49066,N_48899,N_48990);
xor U49067 (N_49067,N_48893,N_48996);
nor U49068 (N_49068,N_48810,N_48982);
or U49069 (N_49069,N_48926,N_48941);
xor U49070 (N_49070,N_48933,N_48812);
nand U49071 (N_49071,N_48855,N_48901);
nor U49072 (N_49072,N_48816,N_48783);
xor U49073 (N_49073,N_48889,N_48993);
nand U49074 (N_49074,N_48878,N_48981);
and U49075 (N_49075,N_48994,N_48847);
or U49076 (N_49076,N_48845,N_48955);
or U49077 (N_49077,N_48958,N_48880);
xor U49078 (N_49078,N_48818,N_48801);
nor U49079 (N_49079,N_48850,N_48991);
and U49080 (N_49080,N_48980,N_48856);
and U49081 (N_49081,N_48793,N_48785);
and U49082 (N_49082,N_48912,N_48983);
nor U49083 (N_49083,N_48917,N_48821);
or U49084 (N_49084,N_48806,N_48833);
or U49085 (N_49085,N_48900,N_48943);
or U49086 (N_49086,N_48760,N_48877);
xor U49087 (N_49087,N_48817,N_48966);
or U49088 (N_49088,N_48876,N_48919);
or U49089 (N_49089,N_48936,N_48918);
nand U49090 (N_49090,N_48923,N_48904);
nor U49091 (N_49091,N_48988,N_48862);
xor U49092 (N_49092,N_48896,N_48804);
and U49093 (N_49093,N_48874,N_48948);
nand U49094 (N_49094,N_48861,N_48977);
nor U49095 (N_49095,N_48828,N_48942);
nand U49096 (N_49096,N_48800,N_48788);
xnor U49097 (N_49097,N_48820,N_48915);
or U49098 (N_49098,N_48960,N_48911);
xor U49099 (N_49099,N_48769,N_48772);
nor U49100 (N_49100,N_48969,N_48753);
nand U49101 (N_49101,N_48838,N_48944);
or U49102 (N_49102,N_48807,N_48907);
and U49103 (N_49103,N_48978,N_48839);
xnor U49104 (N_49104,N_48796,N_48792);
xnor U49105 (N_49105,N_48961,N_48921);
nor U49106 (N_49106,N_48819,N_48995);
or U49107 (N_49107,N_48766,N_48866);
or U49108 (N_49108,N_48773,N_48950);
nor U49109 (N_49109,N_48892,N_48997);
and U49110 (N_49110,N_48924,N_48784);
nor U49111 (N_49111,N_48869,N_48913);
and U49112 (N_49112,N_48967,N_48832);
nor U49113 (N_49113,N_48754,N_48859);
or U49114 (N_49114,N_48888,N_48959);
xnor U49115 (N_49115,N_48830,N_48795);
xor U49116 (N_49116,N_48970,N_48945);
xor U49117 (N_49117,N_48756,N_48794);
xnor U49118 (N_49118,N_48932,N_48827);
or U49119 (N_49119,N_48873,N_48902);
nand U49120 (N_49120,N_48956,N_48968);
and U49121 (N_49121,N_48844,N_48849);
and U49122 (N_49122,N_48951,N_48813);
and U49123 (N_49123,N_48846,N_48751);
xnor U49124 (N_49124,N_48835,N_48851);
and U49125 (N_49125,N_48936,N_48976);
nand U49126 (N_49126,N_48980,N_48830);
nand U49127 (N_49127,N_48780,N_48943);
or U49128 (N_49128,N_48752,N_48895);
xnor U49129 (N_49129,N_48856,N_48872);
xor U49130 (N_49130,N_48982,N_48882);
or U49131 (N_49131,N_48784,N_48897);
xor U49132 (N_49132,N_48795,N_48974);
or U49133 (N_49133,N_48867,N_48831);
and U49134 (N_49134,N_48817,N_48842);
nand U49135 (N_49135,N_48828,N_48989);
or U49136 (N_49136,N_48950,N_48826);
or U49137 (N_49137,N_48881,N_48926);
nand U49138 (N_49138,N_48802,N_48791);
or U49139 (N_49139,N_48783,N_48833);
and U49140 (N_49140,N_48825,N_48897);
nor U49141 (N_49141,N_48972,N_48861);
and U49142 (N_49142,N_48944,N_48771);
and U49143 (N_49143,N_48870,N_48823);
xnor U49144 (N_49144,N_48920,N_48892);
and U49145 (N_49145,N_48807,N_48764);
and U49146 (N_49146,N_48891,N_48911);
nor U49147 (N_49147,N_48856,N_48884);
and U49148 (N_49148,N_48928,N_48994);
xor U49149 (N_49149,N_48822,N_48981);
nand U49150 (N_49150,N_48786,N_48922);
or U49151 (N_49151,N_48982,N_48946);
and U49152 (N_49152,N_48997,N_48775);
nand U49153 (N_49153,N_48966,N_48879);
and U49154 (N_49154,N_48919,N_48852);
xnor U49155 (N_49155,N_48831,N_48894);
and U49156 (N_49156,N_48904,N_48961);
xnor U49157 (N_49157,N_48987,N_48819);
or U49158 (N_49158,N_48841,N_48899);
nor U49159 (N_49159,N_48849,N_48820);
and U49160 (N_49160,N_48838,N_48794);
and U49161 (N_49161,N_48869,N_48895);
nor U49162 (N_49162,N_48898,N_48772);
or U49163 (N_49163,N_48958,N_48995);
and U49164 (N_49164,N_48983,N_48840);
or U49165 (N_49165,N_48752,N_48971);
xnor U49166 (N_49166,N_48901,N_48935);
nor U49167 (N_49167,N_48802,N_48840);
xor U49168 (N_49168,N_48959,N_48981);
nand U49169 (N_49169,N_48824,N_48915);
and U49170 (N_49170,N_48918,N_48839);
or U49171 (N_49171,N_48968,N_48949);
xnor U49172 (N_49172,N_48780,N_48915);
nand U49173 (N_49173,N_48842,N_48865);
or U49174 (N_49174,N_48860,N_48900);
nand U49175 (N_49175,N_48865,N_48927);
nor U49176 (N_49176,N_48817,N_48970);
xor U49177 (N_49177,N_48819,N_48953);
and U49178 (N_49178,N_48847,N_48797);
nor U49179 (N_49179,N_48859,N_48794);
nor U49180 (N_49180,N_48866,N_48858);
or U49181 (N_49181,N_48759,N_48893);
or U49182 (N_49182,N_48820,N_48792);
and U49183 (N_49183,N_48854,N_48814);
nor U49184 (N_49184,N_48752,N_48943);
nor U49185 (N_49185,N_48971,N_48761);
nand U49186 (N_49186,N_48754,N_48840);
xnor U49187 (N_49187,N_48967,N_48905);
nor U49188 (N_49188,N_48859,N_48880);
xnor U49189 (N_49189,N_48994,N_48793);
nand U49190 (N_49190,N_48936,N_48922);
nor U49191 (N_49191,N_48858,N_48905);
nor U49192 (N_49192,N_48922,N_48907);
or U49193 (N_49193,N_48828,N_48817);
xnor U49194 (N_49194,N_48913,N_48910);
nor U49195 (N_49195,N_48972,N_48849);
xor U49196 (N_49196,N_48883,N_48970);
xnor U49197 (N_49197,N_48755,N_48766);
and U49198 (N_49198,N_48947,N_48864);
nand U49199 (N_49199,N_48858,N_48870);
nand U49200 (N_49200,N_48966,N_48999);
and U49201 (N_49201,N_48917,N_48765);
nor U49202 (N_49202,N_48756,N_48830);
nor U49203 (N_49203,N_48865,N_48880);
or U49204 (N_49204,N_48997,N_48808);
nand U49205 (N_49205,N_48910,N_48758);
xnor U49206 (N_49206,N_48827,N_48996);
and U49207 (N_49207,N_48872,N_48914);
xor U49208 (N_49208,N_48812,N_48859);
xnor U49209 (N_49209,N_48930,N_48931);
nand U49210 (N_49210,N_48885,N_48864);
and U49211 (N_49211,N_48998,N_48950);
xor U49212 (N_49212,N_48861,N_48979);
xnor U49213 (N_49213,N_48863,N_48895);
or U49214 (N_49214,N_48979,N_48929);
xor U49215 (N_49215,N_48863,N_48926);
or U49216 (N_49216,N_48904,N_48907);
nor U49217 (N_49217,N_48809,N_48822);
and U49218 (N_49218,N_48842,N_48920);
xor U49219 (N_49219,N_48859,N_48802);
and U49220 (N_49220,N_48940,N_48828);
or U49221 (N_49221,N_48751,N_48920);
xnor U49222 (N_49222,N_48824,N_48772);
and U49223 (N_49223,N_48975,N_48951);
nor U49224 (N_49224,N_48989,N_48802);
and U49225 (N_49225,N_48979,N_48840);
xor U49226 (N_49226,N_48990,N_48755);
and U49227 (N_49227,N_48994,N_48815);
and U49228 (N_49228,N_48825,N_48814);
and U49229 (N_49229,N_48993,N_48917);
xnor U49230 (N_49230,N_48871,N_48862);
nor U49231 (N_49231,N_48885,N_48990);
nor U49232 (N_49232,N_48973,N_48815);
and U49233 (N_49233,N_48787,N_48994);
nor U49234 (N_49234,N_48761,N_48896);
nand U49235 (N_49235,N_48995,N_48977);
nand U49236 (N_49236,N_48989,N_48808);
or U49237 (N_49237,N_48866,N_48897);
or U49238 (N_49238,N_48864,N_48774);
or U49239 (N_49239,N_48791,N_48970);
xnor U49240 (N_49240,N_48778,N_48800);
or U49241 (N_49241,N_48755,N_48909);
xnor U49242 (N_49242,N_48764,N_48878);
xor U49243 (N_49243,N_48858,N_48922);
xor U49244 (N_49244,N_48791,N_48972);
xnor U49245 (N_49245,N_48985,N_48977);
and U49246 (N_49246,N_48804,N_48976);
nand U49247 (N_49247,N_48945,N_48872);
and U49248 (N_49248,N_48937,N_48891);
xor U49249 (N_49249,N_48821,N_48971);
and U49250 (N_49250,N_49149,N_49241);
and U49251 (N_49251,N_49073,N_49161);
xor U49252 (N_49252,N_49202,N_49224);
nand U49253 (N_49253,N_49155,N_49021);
or U49254 (N_49254,N_49162,N_49176);
nor U49255 (N_49255,N_49214,N_49197);
and U49256 (N_49256,N_49005,N_49036);
nand U49257 (N_49257,N_49054,N_49025);
and U49258 (N_49258,N_49203,N_49159);
nand U49259 (N_49259,N_49167,N_49110);
nand U49260 (N_49260,N_49218,N_49194);
or U49261 (N_49261,N_49219,N_49153);
or U49262 (N_49262,N_49081,N_49136);
xnor U49263 (N_49263,N_49015,N_49145);
xnor U49264 (N_49264,N_49041,N_49105);
nand U49265 (N_49265,N_49146,N_49029);
xor U49266 (N_49266,N_49121,N_49221);
or U49267 (N_49267,N_49094,N_49068);
nor U49268 (N_49268,N_49130,N_49141);
or U49269 (N_49269,N_49216,N_49051);
nor U49270 (N_49270,N_49037,N_49151);
or U49271 (N_49271,N_49143,N_49038);
nand U49272 (N_49272,N_49229,N_49101);
xnor U49273 (N_49273,N_49012,N_49052);
and U49274 (N_49274,N_49230,N_49011);
or U49275 (N_49275,N_49180,N_49192);
or U49276 (N_49276,N_49215,N_49089);
and U49277 (N_49277,N_49080,N_49236);
xnor U49278 (N_49278,N_49239,N_49211);
nor U49279 (N_49279,N_49075,N_49008);
or U49280 (N_49280,N_49077,N_49160);
nor U49281 (N_49281,N_49246,N_49033);
and U49282 (N_49282,N_49083,N_49126);
xnor U49283 (N_49283,N_49098,N_49165);
xor U49284 (N_49284,N_49193,N_49064);
xnor U49285 (N_49285,N_49240,N_49173);
xnor U49286 (N_49286,N_49132,N_49002);
xor U49287 (N_49287,N_49185,N_49028);
nand U49288 (N_49288,N_49128,N_49040);
nor U49289 (N_49289,N_49009,N_49096);
nand U49290 (N_49290,N_49204,N_49117);
nand U49291 (N_49291,N_49168,N_49006);
nor U49292 (N_49292,N_49024,N_49044);
nand U49293 (N_49293,N_49122,N_49048);
nor U49294 (N_49294,N_49109,N_49062);
nand U49295 (N_49295,N_49129,N_49187);
and U49296 (N_49296,N_49088,N_49099);
nand U49297 (N_49297,N_49183,N_49093);
nor U49298 (N_49298,N_49107,N_49133);
xnor U49299 (N_49299,N_49195,N_49209);
and U49300 (N_49300,N_49220,N_49116);
nor U49301 (N_49301,N_49043,N_49138);
xnor U49302 (N_49302,N_49164,N_49152);
nor U49303 (N_49303,N_49090,N_49057);
nor U49304 (N_49304,N_49147,N_49247);
nand U49305 (N_49305,N_49014,N_49091);
nand U49306 (N_49306,N_49157,N_49156);
and U49307 (N_49307,N_49233,N_49027);
nor U49308 (N_49308,N_49158,N_49030);
and U49309 (N_49309,N_49188,N_49100);
nand U49310 (N_49310,N_49127,N_49184);
nor U49311 (N_49311,N_49119,N_49046);
nor U49312 (N_49312,N_49182,N_49172);
xor U49313 (N_49313,N_49245,N_49243);
nand U49314 (N_49314,N_49106,N_49154);
nand U49315 (N_49315,N_49238,N_49067);
or U49316 (N_49316,N_49069,N_49023);
nor U49317 (N_49317,N_49082,N_49108);
nor U49318 (N_49318,N_49174,N_49178);
nand U49319 (N_49319,N_49104,N_49010);
and U49320 (N_49320,N_49087,N_49072);
and U49321 (N_49321,N_49169,N_49134);
nand U49322 (N_49322,N_49242,N_49125);
and U49323 (N_49323,N_49166,N_49102);
or U49324 (N_49324,N_49163,N_49066);
or U49325 (N_49325,N_49189,N_49179);
xor U49326 (N_49326,N_49206,N_49001);
nor U49327 (N_49327,N_49115,N_49000);
nor U49328 (N_49328,N_49018,N_49234);
xnor U49329 (N_49329,N_49228,N_49056);
nor U49330 (N_49330,N_49017,N_49170);
or U49331 (N_49331,N_49191,N_49013);
or U49332 (N_49332,N_49060,N_49231);
and U49333 (N_49333,N_49227,N_49111);
nor U49334 (N_49334,N_49225,N_49124);
and U49335 (N_49335,N_49200,N_49113);
or U49336 (N_49336,N_49061,N_49059);
and U49337 (N_49337,N_49237,N_49086);
or U49338 (N_49338,N_49144,N_49055);
nor U49339 (N_49339,N_49045,N_49074);
nand U49340 (N_49340,N_49137,N_49065);
or U49341 (N_49341,N_49198,N_49097);
nand U49342 (N_49342,N_49084,N_49213);
xnor U49343 (N_49343,N_49020,N_49235);
or U49344 (N_49344,N_49142,N_49114);
nor U49345 (N_49345,N_49022,N_49007);
nor U49346 (N_49346,N_49207,N_49208);
or U49347 (N_49347,N_49016,N_49076);
xor U49348 (N_49348,N_49131,N_49171);
nand U49349 (N_49349,N_49201,N_49212);
nor U49350 (N_49350,N_49177,N_49123);
and U49351 (N_49351,N_49150,N_49139);
or U49352 (N_49352,N_49079,N_49249);
nor U49353 (N_49353,N_49026,N_49063);
or U49354 (N_49354,N_49135,N_49047);
and U49355 (N_49355,N_49092,N_49181);
xnor U49356 (N_49356,N_49205,N_49223);
xor U49357 (N_49357,N_49118,N_49032);
xor U49358 (N_49358,N_49071,N_49190);
nand U49359 (N_49359,N_49050,N_49095);
nor U49360 (N_49360,N_49217,N_49034);
xnor U49361 (N_49361,N_49186,N_49120);
and U49362 (N_49362,N_49039,N_49058);
nand U49363 (N_49363,N_49049,N_49003);
or U49364 (N_49364,N_49222,N_49019);
xor U49365 (N_49365,N_49244,N_49140);
or U49366 (N_49366,N_49112,N_49078);
xor U49367 (N_49367,N_49004,N_49031);
or U49368 (N_49368,N_49070,N_49085);
nor U49369 (N_49369,N_49226,N_49248);
xor U49370 (N_49370,N_49196,N_49148);
or U49371 (N_49371,N_49210,N_49053);
and U49372 (N_49372,N_49175,N_49042);
nand U49373 (N_49373,N_49103,N_49035);
and U49374 (N_49374,N_49232,N_49199);
nor U49375 (N_49375,N_49047,N_49234);
or U49376 (N_49376,N_49047,N_49032);
nand U49377 (N_49377,N_49182,N_49031);
or U49378 (N_49378,N_49161,N_49218);
nor U49379 (N_49379,N_49147,N_49074);
or U49380 (N_49380,N_49026,N_49008);
and U49381 (N_49381,N_49113,N_49062);
nand U49382 (N_49382,N_49037,N_49122);
xnor U49383 (N_49383,N_49123,N_49017);
or U49384 (N_49384,N_49170,N_49207);
nor U49385 (N_49385,N_49056,N_49024);
xnor U49386 (N_49386,N_49050,N_49180);
and U49387 (N_49387,N_49078,N_49023);
xor U49388 (N_49388,N_49072,N_49150);
nor U49389 (N_49389,N_49143,N_49041);
xor U49390 (N_49390,N_49114,N_49230);
or U49391 (N_49391,N_49153,N_49084);
xnor U49392 (N_49392,N_49007,N_49174);
nor U49393 (N_49393,N_49224,N_49122);
nand U49394 (N_49394,N_49160,N_49091);
and U49395 (N_49395,N_49186,N_49119);
and U49396 (N_49396,N_49059,N_49239);
nand U49397 (N_49397,N_49118,N_49165);
nand U49398 (N_49398,N_49230,N_49142);
nor U49399 (N_49399,N_49025,N_49037);
nand U49400 (N_49400,N_49193,N_49049);
nor U49401 (N_49401,N_49110,N_49145);
nor U49402 (N_49402,N_49094,N_49239);
nor U49403 (N_49403,N_49140,N_49020);
xnor U49404 (N_49404,N_49162,N_49113);
nor U49405 (N_49405,N_49212,N_49154);
nand U49406 (N_49406,N_49073,N_49220);
or U49407 (N_49407,N_49247,N_49122);
xnor U49408 (N_49408,N_49196,N_49057);
nand U49409 (N_49409,N_49168,N_49183);
nor U49410 (N_49410,N_49099,N_49216);
or U49411 (N_49411,N_49246,N_49232);
nand U49412 (N_49412,N_49105,N_49118);
nand U49413 (N_49413,N_49058,N_49107);
nand U49414 (N_49414,N_49104,N_49078);
xnor U49415 (N_49415,N_49198,N_49178);
or U49416 (N_49416,N_49221,N_49065);
nor U49417 (N_49417,N_49166,N_49028);
xnor U49418 (N_49418,N_49026,N_49176);
and U49419 (N_49419,N_49165,N_49100);
and U49420 (N_49420,N_49148,N_49020);
nor U49421 (N_49421,N_49145,N_49143);
or U49422 (N_49422,N_49107,N_49095);
nor U49423 (N_49423,N_49098,N_49143);
and U49424 (N_49424,N_49217,N_49077);
or U49425 (N_49425,N_49248,N_49034);
xnor U49426 (N_49426,N_49043,N_49147);
and U49427 (N_49427,N_49095,N_49011);
nor U49428 (N_49428,N_49018,N_49080);
xor U49429 (N_49429,N_49156,N_49185);
nand U49430 (N_49430,N_49096,N_49183);
xor U49431 (N_49431,N_49049,N_49097);
nor U49432 (N_49432,N_49065,N_49223);
xnor U49433 (N_49433,N_49034,N_49239);
and U49434 (N_49434,N_49214,N_49211);
nor U49435 (N_49435,N_49025,N_49139);
nand U49436 (N_49436,N_49196,N_49020);
nand U49437 (N_49437,N_49127,N_49000);
xnor U49438 (N_49438,N_49172,N_49101);
or U49439 (N_49439,N_49191,N_49065);
nand U49440 (N_49440,N_49013,N_49220);
xnor U49441 (N_49441,N_49242,N_49249);
and U49442 (N_49442,N_49120,N_49004);
and U49443 (N_49443,N_49137,N_49016);
nor U49444 (N_49444,N_49042,N_49215);
nor U49445 (N_49445,N_49035,N_49241);
and U49446 (N_49446,N_49130,N_49043);
or U49447 (N_49447,N_49141,N_49096);
and U49448 (N_49448,N_49068,N_49243);
or U49449 (N_49449,N_49221,N_49218);
nor U49450 (N_49450,N_49230,N_49021);
and U49451 (N_49451,N_49165,N_49018);
and U49452 (N_49452,N_49067,N_49091);
and U49453 (N_49453,N_49162,N_49007);
nand U49454 (N_49454,N_49239,N_49069);
nand U49455 (N_49455,N_49198,N_49189);
nand U49456 (N_49456,N_49058,N_49054);
nand U49457 (N_49457,N_49148,N_49038);
nand U49458 (N_49458,N_49078,N_49010);
and U49459 (N_49459,N_49210,N_49135);
nand U49460 (N_49460,N_49227,N_49001);
or U49461 (N_49461,N_49000,N_49062);
xor U49462 (N_49462,N_49210,N_49042);
xor U49463 (N_49463,N_49114,N_49200);
and U49464 (N_49464,N_49027,N_49196);
nor U49465 (N_49465,N_49034,N_49189);
xnor U49466 (N_49466,N_49041,N_49243);
nand U49467 (N_49467,N_49193,N_49248);
nand U49468 (N_49468,N_49222,N_49159);
xor U49469 (N_49469,N_49093,N_49031);
or U49470 (N_49470,N_49117,N_49028);
nor U49471 (N_49471,N_49022,N_49020);
or U49472 (N_49472,N_49230,N_49034);
nand U49473 (N_49473,N_49034,N_49174);
xnor U49474 (N_49474,N_49049,N_49103);
nor U49475 (N_49475,N_49209,N_49045);
or U49476 (N_49476,N_49247,N_49107);
nor U49477 (N_49477,N_49082,N_49089);
or U49478 (N_49478,N_49048,N_49206);
xnor U49479 (N_49479,N_49161,N_49183);
nor U49480 (N_49480,N_49058,N_49084);
xnor U49481 (N_49481,N_49041,N_49042);
and U49482 (N_49482,N_49036,N_49015);
nor U49483 (N_49483,N_49132,N_49242);
nand U49484 (N_49484,N_49224,N_49130);
or U49485 (N_49485,N_49180,N_49100);
nor U49486 (N_49486,N_49228,N_49010);
nor U49487 (N_49487,N_49122,N_49194);
or U49488 (N_49488,N_49086,N_49030);
xnor U49489 (N_49489,N_49244,N_49023);
xor U49490 (N_49490,N_49166,N_49123);
nand U49491 (N_49491,N_49167,N_49098);
nand U49492 (N_49492,N_49210,N_49128);
nor U49493 (N_49493,N_49044,N_49199);
nor U49494 (N_49494,N_49208,N_49248);
and U49495 (N_49495,N_49051,N_49160);
and U49496 (N_49496,N_49014,N_49188);
or U49497 (N_49497,N_49244,N_49243);
nand U49498 (N_49498,N_49183,N_49052);
and U49499 (N_49499,N_49096,N_49160);
xnor U49500 (N_49500,N_49393,N_49445);
nand U49501 (N_49501,N_49250,N_49268);
nor U49502 (N_49502,N_49339,N_49490);
xor U49503 (N_49503,N_49378,N_49322);
and U49504 (N_49504,N_49447,N_49377);
and U49505 (N_49505,N_49293,N_49416);
xnor U49506 (N_49506,N_49468,N_49381);
or U49507 (N_49507,N_49434,N_49388);
xnor U49508 (N_49508,N_49282,N_49408);
and U49509 (N_49509,N_49478,N_49382);
or U49510 (N_49510,N_49277,N_49261);
and U49511 (N_49511,N_49439,N_49356);
nor U49512 (N_49512,N_49397,N_49488);
xor U49513 (N_49513,N_49302,N_49265);
nand U49514 (N_49514,N_49287,N_49290);
or U49515 (N_49515,N_49319,N_49442);
or U49516 (N_49516,N_49316,N_49274);
and U49517 (N_49517,N_49384,N_49299);
nor U49518 (N_49518,N_49332,N_49495);
xor U49519 (N_49519,N_49491,N_49361);
and U49520 (N_49520,N_49362,N_49320);
nand U49521 (N_49521,N_49459,N_49324);
nand U49522 (N_49522,N_49453,N_49304);
nor U49523 (N_49523,N_49380,N_49266);
xnor U49524 (N_49524,N_49341,N_49404);
or U49525 (N_49525,N_49485,N_49267);
and U49526 (N_49526,N_49461,N_49275);
and U49527 (N_49527,N_49292,N_49374);
xor U49528 (N_49528,N_49481,N_49326);
and U49529 (N_49529,N_49422,N_49463);
nand U49530 (N_49530,N_49263,N_49494);
nand U49531 (N_49531,N_49376,N_49493);
and U49532 (N_49532,N_49333,N_49387);
or U49533 (N_49533,N_49350,N_49371);
xnor U49534 (N_49534,N_49252,N_49348);
nand U49535 (N_49535,N_49497,N_49251);
or U49536 (N_49536,N_49432,N_49424);
nor U49537 (N_49537,N_49480,N_49271);
and U49538 (N_49538,N_49325,N_49345);
and U49539 (N_49539,N_49396,N_49431);
xnor U49540 (N_49540,N_49285,N_49300);
nor U49541 (N_49541,N_49344,N_49270);
or U49542 (N_49542,N_49430,N_49272);
and U49543 (N_49543,N_49449,N_49357);
or U49544 (N_49544,N_49437,N_49417);
nor U49545 (N_49545,N_49343,N_49262);
or U49546 (N_49546,N_49383,N_49429);
and U49547 (N_49547,N_49421,N_49401);
xor U49548 (N_49548,N_49425,N_49342);
nor U49549 (N_49549,N_49406,N_49457);
nor U49550 (N_49550,N_49465,N_49291);
xnor U49551 (N_49551,N_49334,N_49394);
and U49552 (N_49552,N_49476,N_49379);
xnor U49553 (N_49553,N_49471,N_49375);
or U49554 (N_49554,N_49330,N_49276);
or U49555 (N_49555,N_49418,N_49351);
and U49556 (N_49556,N_49255,N_49411);
xor U49557 (N_49557,N_49415,N_49428);
xor U49558 (N_49558,N_49354,N_49456);
nand U49559 (N_49559,N_49349,N_49328);
xnor U49560 (N_49560,N_49368,N_49352);
and U49561 (N_49561,N_49420,N_49256);
and U49562 (N_49562,N_49366,N_49281);
nor U49563 (N_49563,N_49288,N_49338);
nand U49564 (N_49564,N_49310,N_49419);
or U49565 (N_49565,N_49448,N_49413);
xor U49566 (N_49566,N_49372,N_49259);
nand U49567 (N_49567,N_49483,N_49492);
xnor U49568 (N_49568,N_49487,N_49269);
and U49569 (N_49569,N_49409,N_49392);
nand U49570 (N_49570,N_49400,N_49306);
and U49571 (N_49571,N_49405,N_49280);
nand U49572 (N_49572,N_49359,N_49295);
nand U49573 (N_49573,N_49298,N_49279);
nand U49574 (N_49574,N_49323,N_49466);
nand U49575 (N_49575,N_49443,N_49460);
nand U49576 (N_49576,N_49451,N_49347);
or U49577 (N_49577,N_49373,N_49364);
nor U49578 (N_49578,N_49499,N_49412);
nand U49579 (N_49579,N_49260,N_49454);
nor U49580 (N_49580,N_49410,N_49427);
nand U49581 (N_49581,N_49264,N_49278);
or U49582 (N_49582,N_49455,N_49331);
nand U49583 (N_49583,N_49438,N_49395);
nor U49584 (N_49584,N_49475,N_49303);
xor U49585 (N_49585,N_49309,N_49486);
nor U49586 (N_49586,N_49467,N_49473);
nor U49587 (N_49587,N_49367,N_49399);
and U49588 (N_49588,N_49321,N_49390);
nor U49589 (N_49589,N_49391,N_49369);
nand U49590 (N_49590,N_49301,N_49346);
or U49591 (N_49591,N_49469,N_49283);
or U49592 (N_49592,N_49258,N_49440);
nand U49593 (N_49593,N_49423,N_49297);
nor U49594 (N_49594,N_49294,N_49313);
nand U49595 (N_49595,N_49462,N_49477);
nand U49596 (N_49596,N_49441,N_49435);
and U49597 (N_49597,N_49482,N_49426);
or U49598 (N_49598,N_49446,N_49414);
nand U49599 (N_49599,N_49403,N_49370);
nor U49600 (N_49600,N_49284,N_49472);
or U49601 (N_49601,N_49305,N_49358);
nand U49602 (N_49602,N_49307,N_49327);
nand U49603 (N_49603,N_49398,N_49498);
nor U49604 (N_49604,N_49479,N_49273);
nand U49605 (N_49605,N_49312,N_49452);
and U49606 (N_49606,N_49489,N_49314);
or U49607 (N_49607,N_49311,N_49433);
nor U49608 (N_49608,N_49254,N_49365);
or U49609 (N_49609,N_49253,N_49315);
nand U49610 (N_49610,N_49470,N_49286);
nor U49611 (N_49611,N_49360,N_49337);
nand U49612 (N_49612,N_49308,N_49458);
nand U49613 (N_49613,N_49296,N_49385);
nand U49614 (N_49614,N_49335,N_49353);
or U49615 (N_49615,N_49363,N_49318);
nand U49616 (N_49616,N_49484,N_49329);
nand U49617 (N_49617,N_49474,N_49464);
nor U49618 (N_49618,N_49340,N_49257);
nand U49619 (N_49619,N_49444,N_49402);
nand U49620 (N_49620,N_49496,N_49355);
xnor U49621 (N_49621,N_49436,N_49336);
nand U49622 (N_49622,N_49289,N_49389);
nor U49623 (N_49623,N_49450,N_49386);
and U49624 (N_49624,N_49317,N_49407);
and U49625 (N_49625,N_49255,N_49321);
and U49626 (N_49626,N_49430,N_49412);
or U49627 (N_49627,N_49270,N_49250);
nand U49628 (N_49628,N_49463,N_49397);
and U49629 (N_49629,N_49420,N_49281);
nor U49630 (N_49630,N_49332,N_49437);
xnor U49631 (N_49631,N_49255,N_49275);
nand U49632 (N_49632,N_49364,N_49323);
nor U49633 (N_49633,N_49454,N_49387);
nor U49634 (N_49634,N_49403,N_49354);
nor U49635 (N_49635,N_49424,N_49393);
nor U49636 (N_49636,N_49377,N_49267);
or U49637 (N_49637,N_49272,N_49366);
and U49638 (N_49638,N_49327,N_49462);
or U49639 (N_49639,N_49293,N_49330);
and U49640 (N_49640,N_49415,N_49361);
nor U49641 (N_49641,N_49443,N_49393);
nor U49642 (N_49642,N_49391,N_49362);
and U49643 (N_49643,N_49316,N_49424);
nand U49644 (N_49644,N_49358,N_49310);
or U49645 (N_49645,N_49291,N_49337);
xor U49646 (N_49646,N_49294,N_49271);
xor U49647 (N_49647,N_49357,N_49428);
xnor U49648 (N_49648,N_49498,N_49321);
xor U49649 (N_49649,N_49269,N_49474);
or U49650 (N_49650,N_49274,N_49365);
nor U49651 (N_49651,N_49298,N_49483);
and U49652 (N_49652,N_49281,N_49492);
xor U49653 (N_49653,N_49435,N_49492);
nand U49654 (N_49654,N_49267,N_49265);
nand U49655 (N_49655,N_49455,N_49344);
nor U49656 (N_49656,N_49472,N_49270);
and U49657 (N_49657,N_49423,N_49436);
or U49658 (N_49658,N_49320,N_49317);
nor U49659 (N_49659,N_49445,N_49356);
nand U49660 (N_49660,N_49298,N_49468);
or U49661 (N_49661,N_49355,N_49311);
or U49662 (N_49662,N_49250,N_49259);
and U49663 (N_49663,N_49254,N_49369);
nor U49664 (N_49664,N_49444,N_49491);
xnor U49665 (N_49665,N_49267,N_49398);
nor U49666 (N_49666,N_49298,N_49320);
nor U49667 (N_49667,N_49408,N_49361);
xor U49668 (N_49668,N_49271,N_49252);
nor U49669 (N_49669,N_49368,N_49487);
nand U49670 (N_49670,N_49370,N_49277);
and U49671 (N_49671,N_49284,N_49354);
nor U49672 (N_49672,N_49379,N_49272);
nand U49673 (N_49673,N_49389,N_49380);
xnor U49674 (N_49674,N_49371,N_49459);
and U49675 (N_49675,N_49368,N_49419);
or U49676 (N_49676,N_49363,N_49452);
and U49677 (N_49677,N_49475,N_49300);
or U49678 (N_49678,N_49319,N_49265);
nand U49679 (N_49679,N_49421,N_49268);
nand U49680 (N_49680,N_49361,N_49340);
and U49681 (N_49681,N_49347,N_49441);
and U49682 (N_49682,N_49251,N_49271);
xor U49683 (N_49683,N_49482,N_49257);
or U49684 (N_49684,N_49495,N_49459);
and U49685 (N_49685,N_49479,N_49475);
and U49686 (N_49686,N_49454,N_49372);
or U49687 (N_49687,N_49456,N_49379);
or U49688 (N_49688,N_49380,N_49455);
nand U49689 (N_49689,N_49379,N_49346);
nor U49690 (N_49690,N_49496,N_49257);
nand U49691 (N_49691,N_49462,N_49498);
nand U49692 (N_49692,N_49432,N_49332);
xor U49693 (N_49693,N_49289,N_49474);
and U49694 (N_49694,N_49337,N_49275);
xnor U49695 (N_49695,N_49423,N_49293);
nand U49696 (N_49696,N_49336,N_49489);
and U49697 (N_49697,N_49462,N_49450);
nand U49698 (N_49698,N_49451,N_49391);
nor U49699 (N_49699,N_49416,N_49317);
nor U49700 (N_49700,N_49413,N_49466);
nand U49701 (N_49701,N_49343,N_49341);
xnor U49702 (N_49702,N_49496,N_49415);
nor U49703 (N_49703,N_49453,N_49469);
and U49704 (N_49704,N_49452,N_49488);
xor U49705 (N_49705,N_49406,N_49371);
nor U49706 (N_49706,N_49278,N_49378);
and U49707 (N_49707,N_49356,N_49278);
or U49708 (N_49708,N_49400,N_49388);
and U49709 (N_49709,N_49491,N_49305);
nand U49710 (N_49710,N_49420,N_49374);
or U49711 (N_49711,N_49421,N_49361);
nand U49712 (N_49712,N_49380,N_49268);
nand U49713 (N_49713,N_49490,N_49348);
nor U49714 (N_49714,N_49351,N_49499);
nand U49715 (N_49715,N_49377,N_49383);
nor U49716 (N_49716,N_49457,N_49368);
xnor U49717 (N_49717,N_49413,N_49473);
or U49718 (N_49718,N_49451,N_49487);
or U49719 (N_49719,N_49388,N_49281);
nor U49720 (N_49720,N_49348,N_49376);
nand U49721 (N_49721,N_49420,N_49263);
and U49722 (N_49722,N_49333,N_49414);
xor U49723 (N_49723,N_49479,N_49346);
and U49724 (N_49724,N_49335,N_49313);
xor U49725 (N_49725,N_49253,N_49482);
nor U49726 (N_49726,N_49410,N_49395);
and U49727 (N_49727,N_49316,N_49344);
nor U49728 (N_49728,N_49398,N_49377);
nand U49729 (N_49729,N_49305,N_49326);
and U49730 (N_49730,N_49401,N_49320);
and U49731 (N_49731,N_49477,N_49299);
nand U49732 (N_49732,N_49399,N_49426);
and U49733 (N_49733,N_49482,N_49371);
xor U49734 (N_49734,N_49292,N_49290);
xnor U49735 (N_49735,N_49457,N_49335);
nand U49736 (N_49736,N_49388,N_49407);
nand U49737 (N_49737,N_49303,N_49335);
nand U49738 (N_49738,N_49448,N_49265);
nor U49739 (N_49739,N_49446,N_49447);
or U49740 (N_49740,N_49434,N_49473);
and U49741 (N_49741,N_49281,N_49306);
xor U49742 (N_49742,N_49275,N_49479);
xor U49743 (N_49743,N_49344,N_49378);
or U49744 (N_49744,N_49411,N_49388);
nand U49745 (N_49745,N_49438,N_49284);
nand U49746 (N_49746,N_49497,N_49400);
xnor U49747 (N_49747,N_49419,N_49397);
or U49748 (N_49748,N_49444,N_49323);
or U49749 (N_49749,N_49457,N_49377);
and U49750 (N_49750,N_49510,N_49679);
nand U49751 (N_49751,N_49519,N_49573);
nor U49752 (N_49752,N_49613,N_49735);
xnor U49753 (N_49753,N_49520,N_49647);
and U49754 (N_49754,N_49577,N_49713);
nor U49755 (N_49755,N_49702,N_49681);
xnor U49756 (N_49756,N_49598,N_49745);
or U49757 (N_49757,N_49686,N_49700);
or U49758 (N_49758,N_49646,N_49583);
nor U49759 (N_49759,N_49589,N_49665);
xor U49760 (N_49760,N_49563,N_49631);
or U49761 (N_49761,N_49524,N_49678);
and U49762 (N_49762,N_49594,N_49661);
nor U49763 (N_49763,N_49662,N_49606);
or U49764 (N_49764,N_49648,N_49699);
nand U49765 (N_49765,N_49557,N_49636);
nor U49766 (N_49766,N_49623,N_49556);
or U49767 (N_49767,N_49644,N_49714);
or U49768 (N_49768,N_49552,N_49582);
nand U49769 (N_49769,N_49640,N_49579);
nand U49770 (N_49770,N_49592,N_49624);
and U49771 (N_49771,N_49600,N_49709);
nand U49772 (N_49772,N_49639,N_49554);
xor U49773 (N_49773,N_49534,N_49518);
nor U49774 (N_49774,N_49720,N_49742);
xnor U49775 (N_49775,N_49544,N_49551);
nand U49776 (N_49776,N_49673,N_49634);
xor U49777 (N_49777,N_49687,N_49568);
or U49778 (N_49778,N_49569,N_49642);
nand U49779 (N_49779,N_49537,N_49629);
xnor U49780 (N_49780,N_49588,N_49549);
and U49781 (N_49781,N_49509,N_49690);
xor U49782 (N_49782,N_49680,N_49747);
nand U49783 (N_49783,N_49707,N_49587);
nor U49784 (N_49784,N_49739,N_49616);
nor U49785 (N_49785,N_49658,N_49635);
nor U49786 (N_49786,N_49531,N_49710);
or U49787 (N_49787,N_49570,N_49649);
nor U49788 (N_49788,N_49541,N_49604);
or U49789 (N_49789,N_49746,N_49528);
xor U49790 (N_49790,N_49501,N_49610);
nand U49791 (N_49791,N_49572,N_49558);
xnor U49792 (N_49792,N_49715,N_49664);
nor U49793 (N_49793,N_49643,N_49591);
xor U49794 (N_49794,N_49550,N_49535);
nand U49795 (N_49795,N_49744,N_49522);
xor U49796 (N_49796,N_49502,N_49729);
xor U49797 (N_49797,N_49593,N_49605);
nand U49798 (N_49798,N_49612,N_49539);
nor U49799 (N_49799,N_49683,N_49533);
nor U49800 (N_49800,N_49650,N_49601);
nor U49801 (N_49801,N_49712,N_49689);
and U49802 (N_49802,N_49672,N_49618);
nand U49803 (N_49803,N_49676,N_49565);
or U49804 (N_49804,N_49682,N_49743);
and U49805 (N_49805,N_49703,N_49637);
xor U49806 (N_49806,N_49677,N_49660);
or U49807 (N_49807,N_49721,N_49627);
nor U49808 (N_49808,N_49740,N_49607);
and U49809 (N_49809,N_49749,N_49599);
and U49810 (N_49810,N_49657,N_49695);
or U49811 (N_49811,N_49580,N_49711);
nand U49812 (N_49812,N_49726,N_49581);
or U49813 (N_49813,N_49717,N_49693);
xor U49814 (N_49814,N_49728,N_49555);
nor U49815 (N_49815,N_49609,N_49641);
and U49816 (N_49816,N_49685,N_49737);
nand U49817 (N_49817,N_49614,N_49575);
and U49818 (N_49818,N_49645,N_49576);
and U49819 (N_49819,N_49529,N_49608);
and U49820 (N_49820,N_49619,N_49514);
nand U49821 (N_49821,N_49603,N_49698);
xnor U49822 (N_49822,N_49527,N_49675);
nand U49823 (N_49823,N_49595,N_49546);
xnor U49824 (N_49824,N_49622,N_49615);
nor U49825 (N_49825,N_49548,N_49571);
or U49826 (N_49826,N_49512,N_49670);
xor U49827 (N_49827,N_49688,N_49734);
nor U49828 (N_49828,N_49525,N_49655);
xor U49829 (N_49829,N_49585,N_49566);
and U49830 (N_49830,N_49564,N_49532);
or U49831 (N_49831,N_49697,N_49724);
nand U49832 (N_49832,N_49540,N_49567);
and U49833 (N_49833,N_49547,N_49500);
or U49834 (N_49834,N_49517,N_49505);
nor U49835 (N_49835,N_49611,N_49506);
or U49836 (N_49836,N_49719,N_49668);
or U49837 (N_49837,N_49730,N_49716);
xnor U49838 (N_49838,N_49706,N_49536);
nand U49839 (N_49839,N_49621,N_49671);
nor U49840 (N_49840,N_49651,N_49654);
xnor U49841 (N_49841,N_49633,N_49653);
xor U49842 (N_49842,N_49590,N_49523);
and U49843 (N_49843,N_49723,N_49727);
nand U49844 (N_49844,N_49602,N_49578);
nand U49845 (N_49845,N_49722,N_49748);
nand U49846 (N_49846,N_49725,N_49694);
nand U49847 (N_49847,N_49597,N_49538);
or U49848 (N_49848,N_49507,N_49692);
or U49849 (N_49849,N_49516,N_49669);
nor U49850 (N_49850,N_49625,N_49545);
xor U49851 (N_49851,N_49630,N_49626);
or U49852 (N_49852,N_49560,N_49684);
or U49853 (N_49853,N_49515,N_49543);
and U49854 (N_49854,N_49632,N_49574);
or U49855 (N_49855,N_49708,N_49542);
or U49856 (N_49856,N_49704,N_49513);
nor U49857 (N_49857,N_49503,N_49521);
nand U49858 (N_49858,N_49718,N_49666);
xor U49859 (N_49859,N_49628,N_49667);
nand U49860 (N_49860,N_49674,N_49620);
and U49861 (N_49861,N_49596,N_49530);
nand U49862 (N_49862,N_49511,N_49584);
nor U49863 (N_49863,N_49696,N_49586);
xnor U49864 (N_49864,N_49741,N_49559);
nand U49865 (N_49865,N_49732,N_49738);
or U49866 (N_49866,N_49659,N_49731);
xnor U49867 (N_49867,N_49508,N_49638);
nand U49868 (N_49868,N_49656,N_49526);
nand U49869 (N_49869,N_49652,N_49663);
and U49870 (N_49870,N_49736,N_49691);
or U49871 (N_49871,N_49504,N_49705);
nor U49872 (N_49872,N_49553,N_49733);
nand U49873 (N_49873,N_49617,N_49561);
and U49874 (N_49874,N_49562,N_49701);
nand U49875 (N_49875,N_49744,N_49610);
nor U49876 (N_49876,N_49587,N_49575);
or U49877 (N_49877,N_49630,N_49731);
xnor U49878 (N_49878,N_49585,N_49637);
and U49879 (N_49879,N_49517,N_49749);
nor U49880 (N_49880,N_49709,N_49568);
and U49881 (N_49881,N_49514,N_49732);
nor U49882 (N_49882,N_49536,N_49697);
xor U49883 (N_49883,N_49564,N_49686);
or U49884 (N_49884,N_49696,N_49739);
and U49885 (N_49885,N_49650,N_49608);
and U49886 (N_49886,N_49595,N_49525);
xor U49887 (N_49887,N_49717,N_49631);
nor U49888 (N_49888,N_49546,N_49722);
xor U49889 (N_49889,N_49696,N_49649);
nand U49890 (N_49890,N_49599,N_49576);
or U49891 (N_49891,N_49702,N_49717);
xnor U49892 (N_49892,N_49502,N_49588);
xor U49893 (N_49893,N_49698,N_49702);
nor U49894 (N_49894,N_49505,N_49504);
and U49895 (N_49895,N_49735,N_49576);
and U49896 (N_49896,N_49553,N_49602);
nor U49897 (N_49897,N_49720,N_49619);
xnor U49898 (N_49898,N_49674,N_49549);
nand U49899 (N_49899,N_49620,N_49623);
or U49900 (N_49900,N_49660,N_49748);
nand U49901 (N_49901,N_49703,N_49582);
and U49902 (N_49902,N_49603,N_49607);
xnor U49903 (N_49903,N_49598,N_49608);
nor U49904 (N_49904,N_49630,N_49543);
or U49905 (N_49905,N_49684,N_49588);
nand U49906 (N_49906,N_49720,N_49641);
and U49907 (N_49907,N_49515,N_49674);
nand U49908 (N_49908,N_49678,N_49551);
and U49909 (N_49909,N_49522,N_49743);
nor U49910 (N_49910,N_49653,N_49649);
nand U49911 (N_49911,N_49521,N_49662);
and U49912 (N_49912,N_49722,N_49639);
and U49913 (N_49913,N_49513,N_49727);
nand U49914 (N_49914,N_49538,N_49575);
nand U49915 (N_49915,N_49543,N_49688);
nand U49916 (N_49916,N_49683,N_49560);
nor U49917 (N_49917,N_49523,N_49624);
or U49918 (N_49918,N_49648,N_49589);
xor U49919 (N_49919,N_49509,N_49601);
nor U49920 (N_49920,N_49579,N_49636);
nand U49921 (N_49921,N_49533,N_49679);
nor U49922 (N_49922,N_49720,N_49694);
nor U49923 (N_49923,N_49643,N_49500);
nor U49924 (N_49924,N_49552,N_49654);
or U49925 (N_49925,N_49711,N_49518);
and U49926 (N_49926,N_49697,N_49506);
nor U49927 (N_49927,N_49699,N_49540);
xor U49928 (N_49928,N_49703,N_49607);
xor U49929 (N_49929,N_49730,N_49547);
nand U49930 (N_49930,N_49516,N_49689);
nor U49931 (N_49931,N_49710,N_49704);
xor U49932 (N_49932,N_49560,N_49694);
xnor U49933 (N_49933,N_49593,N_49646);
nand U49934 (N_49934,N_49746,N_49740);
xnor U49935 (N_49935,N_49557,N_49534);
xnor U49936 (N_49936,N_49732,N_49683);
xnor U49937 (N_49937,N_49607,N_49733);
nor U49938 (N_49938,N_49522,N_49591);
xnor U49939 (N_49939,N_49516,N_49657);
xnor U49940 (N_49940,N_49518,N_49744);
or U49941 (N_49941,N_49653,N_49617);
nand U49942 (N_49942,N_49560,N_49522);
nand U49943 (N_49943,N_49573,N_49649);
xnor U49944 (N_49944,N_49681,N_49742);
nand U49945 (N_49945,N_49504,N_49653);
or U49946 (N_49946,N_49659,N_49600);
xnor U49947 (N_49947,N_49558,N_49512);
nor U49948 (N_49948,N_49636,N_49718);
xnor U49949 (N_49949,N_49607,N_49641);
nand U49950 (N_49950,N_49573,N_49535);
and U49951 (N_49951,N_49629,N_49508);
nand U49952 (N_49952,N_49727,N_49739);
and U49953 (N_49953,N_49667,N_49640);
and U49954 (N_49954,N_49722,N_49703);
nand U49955 (N_49955,N_49551,N_49724);
nand U49956 (N_49956,N_49626,N_49533);
and U49957 (N_49957,N_49731,N_49547);
xnor U49958 (N_49958,N_49608,N_49611);
nor U49959 (N_49959,N_49577,N_49599);
or U49960 (N_49960,N_49668,N_49677);
and U49961 (N_49961,N_49570,N_49568);
nand U49962 (N_49962,N_49660,N_49578);
nand U49963 (N_49963,N_49660,N_49542);
nor U49964 (N_49964,N_49655,N_49723);
nor U49965 (N_49965,N_49704,N_49512);
nand U49966 (N_49966,N_49514,N_49607);
and U49967 (N_49967,N_49605,N_49587);
or U49968 (N_49968,N_49596,N_49685);
nor U49969 (N_49969,N_49669,N_49693);
nand U49970 (N_49970,N_49593,N_49610);
nor U49971 (N_49971,N_49517,N_49671);
or U49972 (N_49972,N_49638,N_49523);
and U49973 (N_49973,N_49738,N_49571);
xor U49974 (N_49974,N_49654,N_49683);
xor U49975 (N_49975,N_49718,N_49607);
or U49976 (N_49976,N_49713,N_49585);
or U49977 (N_49977,N_49643,N_49632);
nor U49978 (N_49978,N_49663,N_49744);
and U49979 (N_49979,N_49575,N_49585);
xnor U49980 (N_49980,N_49745,N_49523);
nor U49981 (N_49981,N_49522,N_49601);
or U49982 (N_49982,N_49537,N_49538);
nor U49983 (N_49983,N_49506,N_49630);
xor U49984 (N_49984,N_49746,N_49527);
and U49985 (N_49985,N_49538,N_49694);
xnor U49986 (N_49986,N_49643,N_49710);
or U49987 (N_49987,N_49743,N_49521);
nor U49988 (N_49988,N_49684,N_49580);
xor U49989 (N_49989,N_49559,N_49634);
or U49990 (N_49990,N_49627,N_49584);
and U49991 (N_49991,N_49637,N_49574);
nand U49992 (N_49992,N_49675,N_49707);
nor U49993 (N_49993,N_49640,N_49735);
nor U49994 (N_49994,N_49732,N_49735);
xnor U49995 (N_49995,N_49742,N_49679);
nand U49996 (N_49996,N_49701,N_49700);
nor U49997 (N_49997,N_49556,N_49662);
and U49998 (N_49998,N_49588,N_49626);
or U49999 (N_49999,N_49744,N_49531);
nand UO_0 (O_0,N_49883,N_49798);
and UO_1 (O_1,N_49824,N_49925);
xnor UO_2 (O_2,N_49951,N_49888);
nand UO_3 (O_3,N_49949,N_49952);
nor UO_4 (O_4,N_49803,N_49794);
nor UO_5 (O_5,N_49909,N_49942);
and UO_6 (O_6,N_49876,N_49819);
xnor UO_7 (O_7,N_49854,N_49974);
and UO_8 (O_8,N_49979,N_49999);
xnor UO_9 (O_9,N_49840,N_49835);
nor UO_10 (O_10,N_49828,N_49958);
xnor UO_11 (O_11,N_49905,N_49929);
and UO_12 (O_12,N_49832,N_49962);
nor UO_13 (O_13,N_49870,N_49928);
xnor UO_14 (O_14,N_49812,N_49908);
and UO_15 (O_15,N_49838,N_49814);
nor UO_16 (O_16,N_49923,N_49796);
nand UO_17 (O_17,N_49841,N_49892);
or UO_18 (O_18,N_49920,N_49931);
nand UO_19 (O_19,N_49831,N_49849);
nand UO_20 (O_20,N_49914,N_49775);
xnor UO_21 (O_21,N_49807,N_49826);
or UO_22 (O_22,N_49784,N_49953);
and UO_23 (O_23,N_49975,N_49777);
and UO_24 (O_24,N_49948,N_49983);
or UO_25 (O_25,N_49782,N_49894);
and UO_26 (O_26,N_49968,N_49761);
nor UO_27 (O_27,N_49842,N_49904);
or UO_28 (O_28,N_49755,N_49885);
and UO_29 (O_29,N_49785,N_49790);
xnor UO_30 (O_30,N_49800,N_49766);
nor UO_31 (O_31,N_49871,N_49995);
and UO_32 (O_32,N_49887,N_49765);
and UO_33 (O_33,N_49919,N_49865);
or UO_34 (O_34,N_49780,N_49986);
or UO_35 (O_35,N_49940,N_49984);
or UO_36 (O_36,N_49753,N_49882);
and UO_37 (O_37,N_49801,N_49813);
and UO_38 (O_38,N_49980,N_49938);
and UO_39 (O_39,N_49770,N_49936);
nor UO_40 (O_40,N_49950,N_49767);
or UO_41 (O_41,N_49963,N_49774);
nor UO_42 (O_42,N_49837,N_49781);
and UO_43 (O_43,N_49990,N_49965);
xnor UO_44 (O_44,N_49930,N_49976);
xor UO_45 (O_45,N_49866,N_49771);
nand UO_46 (O_46,N_49997,N_49922);
and UO_47 (O_47,N_49805,N_49939);
xnor UO_48 (O_48,N_49998,N_49763);
or UO_49 (O_49,N_49907,N_49847);
or UO_50 (O_50,N_49806,N_49864);
and UO_51 (O_51,N_49880,N_49903);
nor UO_52 (O_52,N_49839,N_49898);
xnor UO_53 (O_53,N_49912,N_49981);
or UO_54 (O_54,N_49833,N_49857);
nand UO_55 (O_55,N_49863,N_49751);
nand UO_56 (O_56,N_49924,N_49941);
and UO_57 (O_57,N_49886,N_49916);
nor UO_58 (O_58,N_49799,N_49897);
nor UO_59 (O_59,N_49985,N_49786);
nor UO_60 (O_60,N_49959,N_49956);
and UO_61 (O_61,N_49966,N_49937);
xnor UO_62 (O_62,N_49867,N_49788);
and UO_63 (O_63,N_49954,N_49756);
nor UO_64 (O_64,N_49964,N_49816);
xnor UO_65 (O_65,N_49988,N_49850);
xor UO_66 (O_66,N_49900,N_49811);
and UO_67 (O_67,N_49844,N_49822);
and UO_68 (O_68,N_49821,N_49890);
nand UO_69 (O_69,N_49817,N_49853);
xor UO_70 (O_70,N_49802,N_49932);
and UO_71 (O_71,N_49830,N_49776);
or UO_72 (O_72,N_49787,N_49757);
or UO_73 (O_73,N_49935,N_49773);
nand UO_74 (O_74,N_49809,N_49759);
nor UO_75 (O_75,N_49915,N_49779);
or UO_76 (O_76,N_49750,N_49795);
xor UO_77 (O_77,N_49827,N_49768);
nor UO_78 (O_78,N_49982,N_49820);
and UO_79 (O_79,N_49851,N_49893);
nor UO_80 (O_80,N_49921,N_49872);
nor UO_81 (O_81,N_49884,N_49933);
nor UO_82 (O_82,N_49996,N_49945);
nand UO_83 (O_83,N_49993,N_49947);
or UO_84 (O_84,N_49791,N_49879);
nor UO_85 (O_85,N_49911,N_49946);
nand UO_86 (O_86,N_49861,N_49772);
and UO_87 (O_87,N_49778,N_49852);
nand UO_88 (O_88,N_49891,N_49955);
or UO_89 (O_89,N_49874,N_49927);
and UO_90 (O_90,N_49856,N_49971);
nor UO_91 (O_91,N_49868,N_49804);
nor UO_92 (O_92,N_49793,N_49918);
xor UO_93 (O_93,N_49846,N_49797);
or UO_94 (O_94,N_49901,N_49792);
and UO_95 (O_95,N_49869,N_49825);
xor UO_96 (O_96,N_49913,N_49758);
and UO_97 (O_97,N_49783,N_49845);
or UO_98 (O_98,N_49943,N_49906);
and UO_99 (O_99,N_49859,N_49823);
and UO_100 (O_100,N_49789,N_49881);
nor UO_101 (O_101,N_49760,N_49808);
or UO_102 (O_102,N_49815,N_49896);
and UO_103 (O_103,N_49862,N_49977);
xnor UO_104 (O_104,N_49899,N_49991);
nand UO_105 (O_105,N_49994,N_49889);
and UO_106 (O_106,N_49860,N_49843);
nor UO_107 (O_107,N_49877,N_49818);
and UO_108 (O_108,N_49944,N_49858);
or UO_109 (O_109,N_49926,N_49873);
and UO_110 (O_110,N_49810,N_49878);
or UO_111 (O_111,N_49969,N_49992);
xnor UO_112 (O_112,N_49957,N_49934);
xnor UO_113 (O_113,N_49910,N_49989);
and UO_114 (O_114,N_49960,N_49917);
nor UO_115 (O_115,N_49764,N_49978);
and UO_116 (O_116,N_49987,N_49829);
or UO_117 (O_117,N_49973,N_49961);
nor UO_118 (O_118,N_49855,N_49752);
nor UO_119 (O_119,N_49972,N_49895);
and UO_120 (O_120,N_49836,N_49769);
and UO_121 (O_121,N_49967,N_49762);
xnor UO_122 (O_122,N_49875,N_49848);
nor UO_123 (O_123,N_49834,N_49902);
xnor UO_124 (O_124,N_49754,N_49970);
nand UO_125 (O_125,N_49929,N_49851);
nor UO_126 (O_126,N_49753,N_49846);
nor UO_127 (O_127,N_49839,N_49816);
xnor UO_128 (O_128,N_49929,N_49895);
xnor UO_129 (O_129,N_49788,N_49949);
xor UO_130 (O_130,N_49908,N_49955);
nand UO_131 (O_131,N_49860,N_49824);
nor UO_132 (O_132,N_49858,N_49891);
nand UO_133 (O_133,N_49893,N_49848);
or UO_134 (O_134,N_49896,N_49880);
xor UO_135 (O_135,N_49798,N_49931);
xor UO_136 (O_136,N_49865,N_49939);
and UO_137 (O_137,N_49927,N_49931);
xor UO_138 (O_138,N_49993,N_49863);
or UO_139 (O_139,N_49894,N_49855);
nor UO_140 (O_140,N_49794,N_49933);
or UO_141 (O_141,N_49902,N_49994);
xnor UO_142 (O_142,N_49962,N_49871);
nor UO_143 (O_143,N_49886,N_49818);
nand UO_144 (O_144,N_49915,N_49778);
nor UO_145 (O_145,N_49902,N_49871);
xnor UO_146 (O_146,N_49774,N_49927);
or UO_147 (O_147,N_49921,N_49997);
nor UO_148 (O_148,N_49894,N_49798);
or UO_149 (O_149,N_49834,N_49943);
or UO_150 (O_150,N_49823,N_49947);
xor UO_151 (O_151,N_49851,N_49846);
and UO_152 (O_152,N_49989,N_49797);
nor UO_153 (O_153,N_49869,N_49933);
nor UO_154 (O_154,N_49923,N_49847);
nor UO_155 (O_155,N_49921,N_49846);
xnor UO_156 (O_156,N_49790,N_49862);
nor UO_157 (O_157,N_49915,N_49942);
and UO_158 (O_158,N_49775,N_49825);
or UO_159 (O_159,N_49901,N_49838);
xor UO_160 (O_160,N_49831,N_49767);
or UO_161 (O_161,N_49842,N_49827);
xor UO_162 (O_162,N_49826,N_49789);
or UO_163 (O_163,N_49891,N_49983);
and UO_164 (O_164,N_49965,N_49839);
or UO_165 (O_165,N_49807,N_49896);
xnor UO_166 (O_166,N_49854,N_49926);
nand UO_167 (O_167,N_49840,N_49774);
xnor UO_168 (O_168,N_49998,N_49874);
nor UO_169 (O_169,N_49841,N_49908);
and UO_170 (O_170,N_49983,N_49994);
xnor UO_171 (O_171,N_49949,N_49917);
and UO_172 (O_172,N_49788,N_49912);
xor UO_173 (O_173,N_49860,N_49911);
or UO_174 (O_174,N_49959,N_49781);
nand UO_175 (O_175,N_49925,N_49917);
and UO_176 (O_176,N_49829,N_49819);
xor UO_177 (O_177,N_49781,N_49997);
xor UO_178 (O_178,N_49984,N_49800);
xor UO_179 (O_179,N_49777,N_49853);
xor UO_180 (O_180,N_49764,N_49950);
nor UO_181 (O_181,N_49790,N_49756);
and UO_182 (O_182,N_49936,N_49791);
nor UO_183 (O_183,N_49987,N_49755);
nand UO_184 (O_184,N_49765,N_49848);
or UO_185 (O_185,N_49963,N_49911);
nand UO_186 (O_186,N_49797,N_49928);
xnor UO_187 (O_187,N_49908,N_49792);
nand UO_188 (O_188,N_49778,N_49933);
and UO_189 (O_189,N_49841,N_49994);
xor UO_190 (O_190,N_49835,N_49876);
and UO_191 (O_191,N_49948,N_49867);
and UO_192 (O_192,N_49820,N_49952);
nand UO_193 (O_193,N_49824,N_49842);
or UO_194 (O_194,N_49931,N_49870);
nand UO_195 (O_195,N_49867,N_49996);
and UO_196 (O_196,N_49763,N_49914);
nand UO_197 (O_197,N_49879,N_49800);
xnor UO_198 (O_198,N_49941,N_49880);
nor UO_199 (O_199,N_49804,N_49855);
nand UO_200 (O_200,N_49841,N_49857);
nand UO_201 (O_201,N_49896,N_49909);
and UO_202 (O_202,N_49828,N_49756);
nand UO_203 (O_203,N_49931,N_49922);
nor UO_204 (O_204,N_49758,N_49975);
xor UO_205 (O_205,N_49958,N_49887);
xnor UO_206 (O_206,N_49808,N_49862);
xnor UO_207 (O_207,N_49972,N_49876);
xor UO_208 (O_208,N_49795,N_49813);
or UO_209 (O_209,N_49753,N_49783);
and UO_210 (O_210,N_49775,N_49857);
xor UO_211 (O_211,N_49919,N_49838);
nor UO_212 (O_212,N_49902,N_49993);
or UO_213 (O_213,N_49863,N_49985);
nor UO_214 (O_214,N_49954,N_49768);
nor UO_215 (O_215,N_49829,N_49881);
nand UO_216 (O_216,N_49767,N_49830);
and UO_217 (O_217,N_49829,N_49954);
or UO_218 (O_218,N_49798,N_49920);
or UO_219 (O_219,N_49750,N_49808);
or UO_220 (O_220,N_49774,N_49932);
and UO_221 (O_221,N_49853,N_49795);
or UO_222 (O_222,N_49762,N_49924);
xor UO_223 (O_223,N_49882,N_49809);
and UO_224 (O_224,N_49929,N_49825);
or UO_225 (O_225,N_49757,N_49894);
and UO_226 (O_226,N_49980,N_49829);
or UO_227 (O_227,N_49984,N_49929);
xor UO_228 (O_228,N_49954,N_49846);
xnor UO_229 (O_229,N_49801,N_49821);
nand UO_230 (O_230,N_49861,N_49954);
nor UO_231 (O_231,N_49751,N_49947);
xnor UO_232 (O_232,N_49923,N_49772);
nand UO_233 (O_233,N_49799,N_49958);
nand UO_234 (O_234,N_49970,N_49812);
or UO_235 (O_235,N_49907,N_49823);
xor UO_236 (O_236,N_49951,N_49838);
nand UO_237 (O_237,N_49808,N_49833);
nor UO_238 (O_238,N_49879,N_49980);
nand UO_239 (O_239,N_49840,N_49798);
nor UO_240 (O_240,N_49899,N_49809);
or UO_241 (O_241,N_49906,N_49968);
nand UO_242 (O_242,N_49900,N_49966);
xor UO_243 (O_243,N_49772,N_49790);
nor UO_244 (O_244,N_49891,N_49889);
nor UO_245 (O_245,N_49890,N_49871);
xnor UO_246 (O_246,N_49824,N_49903);
nor UO_247 (O_247,N_49935,N_49833);
nor UO_248 (O_248,N_49880,N_49974);
or UO_249 (O_249,N_49938,N_49835);
and UO_250 (O_250,N_49943,N_49764);
nand UO_251 (O_251,N_49764,N_49975);
nor UO_252 (O_252,N_49759,N_49838);
or UO_253 (O_253,N_49869,N_49964);
or UO_254 (O_254,N_49831,N_49966);
nand UO_255 (O_255,N_49929,N_49934);
nand UO_256 (O_256,N_49966,N_49989);
or UO_257 (O_257,N_49917,N_49921);
nor UO_258 (O_258,N_49953,N_49881);
nor UO_259 (O_259,N_49887,N_49895);
and UO_260 (O_260,N_49776,N_49989);
nor UO_261 (O_261,N_49830,N_49804);
or UO_262 (O_262,N_49785,N_49799);
or UO_263 (O_263,N_49895,N_49936);
xor UO_264 (O_264,N_49952,N_49922);
nand UO_265 (O_265,N_49863,N_49949);
nor UO_266 (O_266,N_49973,N_49850);
nand UO_267 (O_267,N_49804,N_49884);
or UO_268 (O_268,N_49770,N_49877);
xnor UO_269 (O_269,N_49769,N_49936);
and UO_270 (O_270,N_49834,N_49999);
nor UO_271 (O_271,N_49903,N_49864);
xnor UO_272 (O_272,N_49868,N_49865);
or UO_273 (O_273,N_49947,N_49832);
nor UO_274 (O_274,N_49795,N_49952);
and UO_275 (O_275,N_49856,N_49961);
nor UO_276 (O_276,N_49781,N_49973);
and UO_277 (O_277,N_49904,N_49891);
and UO_278 (O_278,N_49875,N_49767);
xnor UO_279 (O_279,N_49889,N_49817);
and UO_280 (O_280,N_49993,N_49849);
nor UO_281 (O_281,N_49915,N_49899);
nor UO_282 (O_282,N_49824,N_49865);
nor UO_283 (O_283,N_49761,N_49768);
xnor UO_284 (O_284,N_49902,N_49892);
and UO_285 (O_285,N_49868,N_49952);
xor UO_286 (O_286,N_49937,N_49829);
nor UO_287 (O_287,N_49965,N_49878);
and UO_288 (O_288,N_49756,N_49892);
or UO_289 (O_289,N_49941,N_49951);
and UO_290 (O_290,N_49806,N_49961);
nand UO_291 (O_291,N_49847,N_49924);
and UO_292 (O_292,N_49770,N_49891);
and UO_293 (O_293,N_49878,N_49892);
xor UO_294 (O_294,N_49990,N_49960);
xnor UO_295 (O_295,N_49852,N_49826);
nand UO_296 (O_296,N_49885,N_49818);
nand UO_297 (O_297,N_49953,N_49916);
or UO_298 (O_298,N_49843,N_49963);
xnor UO_299 (O_299,N_49991,N_49795);
and UO_300 (O_300,N_49797,N_49773);
and UO_301 (O_301,N_49912,N_49969);
nand UO_302 (O_302,N_49845,N_49878);
nand UO_303 (O_303,N_49994,N_49995);
nor UO_304 (O_304,N_49831,N_49848);
xor UO_305 (O_305,N_49958,N_49902);
and UO_306 (O_306,N_49954,N_49791);
nand UO_307 (O_307,N_49969,N_49790);
and UO_308 (O_308,N_49969,N_49768);
or UO_309 (O_309,N_49865,N_49917);
and UO_310 (O_310,N_49923,N_49781);
and UO_311 (O_311,N_49967,N_49821);
nor UO_312 (O_312,N_49846,N_49779);
nand UO_313 (O_313,N_49801,N_49872);
or UO_314 (O_314,N_49794,N_49781);
or UO_315 (O_315,N_49800,N_49912);
nor UO_316 (O_316,N_49896,N_49797);
or UO_317 (O_317,N_49851,N_49956);
xnor UO_318 (O_318,N_49822,N_49980);
nor UO_319 (O_319,N_49836,N_49933);
or UO_320 (O_320,N_49921,N_49776);
nand UO_321 (O_321,N_49926,N_49884);
or UO_322 (O_322,N_49813,N_49983);
nand UO_323 (O_323,N_49988,N_49998);
nor UO_324 (O_324,N_49979,N_49821);
nand UO_325 (O_325,N_49881,N_49843);
or UO_326 (O_326,N_49824,N_49868);
nand UO_327 (O_327,N_49990,N_49782);
nor UO_328 (O_328,N_49893,N_49791);
and UO_329 (O_329,N_49870,N_49850);
xor UO_330 (O_330,N_49882,N_49954);
and UO_331 (O_331,N_49759,N_49904);
nor UO_332 (O_332,N_49902,N_49919);
nor UO_333 (O_333,N_49864,N_49844);
or UO_334 (O_334,N_49767,N_49883);
and UO_335 (O_335,N_49966,N_49955);
nor UO_336 (O_336,N_49792,N_49878);
xor UO_337 (O_337,N_49763,N_49979);
nor UO_338 (O_338,N_49871,N_49853);
nor UO_339 (O_339,N_49755,N_49862);
xnor UO_340 (O_340,N_49869,N_49769);
nand UO_341 (O_341,N_49875,N_49827);
or UO_342 (O_342,N_49927,N_49992);
nor UO_343 (O_343,N_49982,N_49775);
or UO_344 (O_344,N_49953,N_49751);
and UO_345 (O_345,N_49816,N_49905);
xnor UO_346 (O_346,N_49939,N_49808);
nor UO_347 (O_347,N_49931,N_49877);
and UO_348 (O_348,N_49756,N_49893);
and UO_349 (O_349,N_49932,N_49870);
nand UO_350 (O_350,N_49849,N_49836);
xnor UO_351 (O_351,N_49972,N_49982);
xnor UO_352 (O_352,N_49827,N_49968);
xor UO_353 (O_353,N_49903,N_49794);
nor UO_354 (O_354,N_49782,N_49974);
or UO_355 (O_355,N_49795,N_49876);
and UO_356 (O_356,N_49840,N_49957);
nand UO_357 (O_357,N_49959,N_49859);
nand UO_358 (O_358,N_49836,N_49995);
nor UO_359 (O_359,N_49862,N_49919);
and UO_360 (O_360,N_49791,N_49889);
or UO_361 (O_361,N_49908,N_49758);
and UO_362 (O_362,N_49777,N_49831);
and UO_363 (O_363,N_49765,N_49897);
and UO_364 (O_364,N_49916,N_49923);
and UO_365 (O_365,N_49856,N_49935);
nor UO_366 (O_366,N_49892,N_49775);
nor UO_367 (O_367,N_49936,N_49833);
xor UO_368 (O_368,N_49867,N_49985);
nand UO_369 (O_369,N_49931,N_49911);
xnor UO_370 (O_370,N_49959,N_49752);
xnor UO_371 (O_371,N_49887,N_49872);
or UO_372 (O_372,N_49977,N_49852);
nor UO_373 (O_373,N_49975,N_49846);
nor UO_374 (O_374,N_49967,N_49774);
xnor UO_375 (O_375,N_49859,N_49836);
and UO_376 (O_376,N_49829,N_49872);
and UO_377 (O_377,N_49887,N_49792);
nand UO_378 (O_378,N_49891,N_49995);
or UO_379 (O_379,N_49888,N_49801);
or UO_380 (O_380,N_49864,N_49967);
nor UO_381 (O_381,N_49876,N_49930);
nor UO_382 (O_382,N_49913,N_49950);
and UO_383 (O_383,N_49981,N_49766);
and UO_384 (O_384,N_49859,N_49820);
and UO_385 (O_385,N_49879,N_49783);
or UO_386 (O_386,N_49953,N_49814);
and UO_387 (O_387,N_49875,N_49999);
nor UO_388 (O_388,N_49837,N_49854);
and UO_389 (O_389,N_49991,N_49872);
or UO_390 (O_390,N_49873,N_49845);
and UO_391 (O_391,N_49912,N_49933);
xor UO_392 (O_392,N_49801,N_49944);
nand UO_393 (O_393,N_49934,N_49866);
or UO_394 (O_394,N_49948,N_49897);
nor UO_395 (O_395,N_49984,N_49815);
xor UO_396 (O_396,N_49954,N_49883);
xor UO_397 (O_397,N_49890,N_49917);
nand UO_398 (O_398,N_49865,N_49851);
nand UO_399 (O_399,N_49934,N_49806);
and UO_400 (O_400,N_49774,N_49896);
or UO_401 (O_401,N_49777,N_49790);
nor UO_402 (O_402,N_49983,N_49938);
xor UO_403 (O_403,N_49775,N_49977);
or UO_404 (O_404,N_49938,N_49843);
xnor UO_405 (O_405,N_49918,N_49907);
xor UO_406 (O_406,N_49755,N_49837);
or UO_407 (O_407,N_49759,N_49788);
or UO_408 (O_408,N_49832,N_49867);
and UO_409 (O_409,N_49931,N_49774);
xor UO_410 (O_410,N_49917,N_49905);
nand UO_411 (O_411,N_49941,N_49884);
nor UO_412 (O_412,N_49817,N_49828);
nor UO_413 (O_413,N_49963,N_49998);
or UO_414 (O_414,N_49890,N_49867);
nand UO_415 (O_415,N_49956,N_49777);
and UO_416 (O_416,N_49948,N_49764);
nand UO_417 (O_417,N_49802,N_49764);
and UO_418 (O_418,N_49898,N_49950);
nor UO_419 (O_419,N_49968,N_49964);
xor UO_420 (O_420,N_49826,N_49984);
and UO_421 (O_421,N_49914,N_49888);
nand UO_422 (O_422,N_49819,N_49943);
or UO_423 (O_423,N_49805,N_49792);
and UO_424 (O_424,N_49786,N_49859);
xnor UO_425 (O_425,N_49873,N_49912);
nand UO_426 (O_426,N_49760,N_49885);
and UO_427 (O_427,N_49967,N_49839);
xnor UO_428 (O_428,N_49831,N_49828);
and UO_429 (O_429,N_49770,N_49982);
nor UO_430 (O_430,N_49878,N_49905);
and UO_431 (O_431,N_49910,N_49825);
or UO_432 (O_432,N_49856,N_49795);
and UO_433 (O_433,N_49890,N_49857);
or UO_434 (O_434,N_49773,N_49751);
or UO_435 (O_435,N_49907,N_49831);
nand UO_436 (O_436,N_49777,N_49875);
or UO_437 (O_437,N_49858,N_49826);
or UO_438 (O_438,N_49857,N_49825);
nor UO_439 (O_439,N_49947,N_49905);
and UO_440 (O_440,N_49981,N_49803);
xnor UO_441 (O_441,N_49795,N_49773);
nand UO_442 (O_442,N_49918,N_49829);
nor UO_443 (O_443,N_49924,N_49818);
and UO_444 (O_444,N_49957,N_49788);
or UO_445 (O_445,N_49866,N_49805);
or UO_446 (O_446,N_49864,N_49949);
or UO_447 (O_447,N_49960,N_49982);
nor UO_448 (O_448,N_49858,N_49762);
xor UO_449 (O_449,N_49855,N_49912);
nor UO_450 (O_450,N_49998,N_49996);
and UO_451 (O_451,N_49866,N_49758);
nor UO_452 (O_452,N_49808,N_49830);
and UO_453 (O_453,N_49945,N_49951);
or UO_454 (O_454,N_49779,N_49866);
nand UO_455 (O_455,N_49944,N_49901);
xnor UO_456 (O_456,N_49944,N_49823);
nor UO_457 (O_457,N_49882,N_49771);
and UO_458 (O_458,N_49952,N_49947);
xor UO_459 (O_459,N_49945,N_49982);
or UO_460 (O_460,N_49829,N_49923);
xor UO_461 (O_461,N_49861,N_49944);
xor UO_462 (O_462,N_49753,N_49992);
nand UO_463 (O_463,N_49895,N_49878);
nand UO_464 (O_464,N_49928,N_49815);
xor UO_465 (O_465,N_49914,N_49960);
and UO_466 (O_466,N_49832,N_49770);
xnor UO_467 (O_467,N_49882,N_49780);
nor UO_468 (O_468,N_49986,N_49759);
xor UO_469 (O_469,N_49965,N_49905);
xor UO_470 (O_470,N_49976,N_49961);
nand UO_471 (O_471,N_49875,N_49785);
nor UO_472 (O_472,N_49772,N_49993);
xor UO_473 (O_473,N_49900,N_49785);
or UO_474 (O_474,N_49843,N_49962);
nand UO_475 (O_475,N_49964,N_49791);
nor UO_476 (O_476,N_49784,N_49853);
and UO_477 (O_477,N_49779,N_49771);
or UO_478 (O_478,N_49871,N_49812);
or UO_479 (O_479,N_49770,N_49975);
nand UO_480 (O_480,N_49771,N_49803);
xnor UO_481 (O_481,N_49981,N_49924);
nor UO_482 (O_482,N_49852,N_49780);
nor UO_483 (O_483,N_49851,N_49866);
nor UO_484 (O_484,N_49836,N_49860);
nand UO_485 (O_485,N_49837,N_49778);
xor UO_486 (O_486,N_49973,N_49809);
nor UO_487 (O_487,N_49822,N_49900);
or UO_488 (O_488,N_49898,N_49933);
nor UO_489 (O_489,N_49751,N_49896);
xor UO_490 (O_490,N_49971,N_49823);
nand UO_491 (O_491,N_49995,N_49972);
and UO_492 (O_492,N_49764,N_49956);
xnor UO_493 (O_493,N_49891,N_49778);
xnor UO_494 (O_494,N_49964,N_49890);
xnor UO_495 (O_495,N_49922,N_49981);
nand UO_496 (O_496,N_49855,N_49901);
nor UO_497 (O_497,N_49862,N_49983);
nand UO_498 (O_498,N_49952,N_49856);
xnor UO_499 (O_499,N_49944,N_49908);
xnor UO_500 (O_500,N_49802,N_49961);
or UO_501 (O_501,N_49750,N_49886);
or UO_502 (O_502,N_49865,N_49781);
xnor UO_503 (O_503,N_49858,N_49979);
or UO_504 (O_504,N_49935,N_49938);
nor UO_505 (O_505,N_49970,N_49806);
xnor UO_506 (O_506,N_49916,N_49825);
or UO_507 (O_507,N_49782,N_49993);
nand UO_508 (O_508,N_49998,N_49840);
nor UO_509 (O_509,N_49789,N_49906);
xor UO_510 (O_510,N_49944,N_49966);
xnor UO_511 (O_511,N_49861,N_49974);
and UO_512 (O_512,N_49880,N_49945);
xnor UO_513 (O_513,N_49916,N_49863);
or UO_514 (O_514,N_49775,N_49894);
nand UO_515 (O_515,N_49899,N_49755);
nor UO_516 (O_516,N_49794,N_49756);
and UO_517 (O_517,N_49935,N_49757);
nand UO_518 (O_518,N_49898,N_49836);
nand UO_519 (O_519,N_49959,N_49814);
and UO_520 (O_520,N_49983,N_49771);
and UO_521 (O_521,N_49757,N_49838);
or UO_522 (O_522,N_49929,N_49915);
or UO_523 (O_523,N_49859,N_49890);
or UO_524 (O_524,N_49991,N_49866);
nand UO_525 (O_525,N_49824,N_49761);
xor UO_526 (O_526,N_49915,N_49874);
nand UO_527 (O_527,N_49870,N_49872);
or UO_528 (O_528,N_49787,N_49762);
nor UO_529 (O_529,N_49830,N_49847);
and UO_530 (O_530,N_49798,N_49906);
or UO_531 (O_531,N_49814,N_49858);
nand UO_532 (O_532,N_49982,N_49936);
nor UO_533 (O_533,N_49850,N_49918);
nor UO_534 (O_534,N_49977,N_49927);
xor UO_535 (O_535,N_49776,N_49848);
xor UO_536 (O_536,N_49751,N_49937);
nor UO_537 (O_537,N_49989,N_49783);
or UO_538 (O_538,N_49858,N_49825);
or UO_539 (O_539,N_49910,N_49796);
and UO_540 (O_540,N_49796,N_49871);
xor UO_541 (O_541,N_49930,N_49839);
or UO_542 (O_542,N_49817,N_49950);
nor UO_543 (O_543,N_49787,N_49986);
and UO_544 (O_544,N_49991,N_49877);
and UO_545 (O_545,N_49959,N_49977);
nor UO_546 (O_546,N_49775,N_49958);
or UO_547 (O_547,N_49933,N_49958);
or UO_548 (O_548,N_49833,N_49918);
nor UO_549 (O_549,N_49815,N_49765);
nor UO_550 (O_550,N_49956,N_49893);
and UO_551 (O_551,N_49979,N_49854);
nand UO_552 (O_552,N_49991,N_49927);
or UO_553 (O_553,N_49850,N_49947);
nand UO_554 (O_554,N_49980,N_49942);
or UO_555 (O_555,N_49801,N_49896);
nor UO_556 (O_556,N_49920,N_49904);
or UO_557 (O_557,N_49941,N_49795);
nand UO_558 (O_558,N_49920,N_49924);
or UO_559 (O_559,N_49799,N_49878);
nand UO_560 (O_560,N_49914,N_49944);
xnor UO_561 (O_561,N_49797,N_49931);
nand UO_562 (O_562,N_49913,N_49815);
xor UO_563 (O_563,N_49752,N_49797);
and UO_564 (O_564,N_49797,N_49997);
nor UO_565 (O_565,N_49848,N_49863);
and UO_566 (O_566,N_49946,N_49773);
nor UO_567 (O_567,N_49958,N_49892);
nand UO_568 (O_568,N_49852,N_49871);
or UO_569 (O_569,N_49769,N_49996);
nor UO_570 (O_570,N_49761,N_49995);
or UO_571 (O_571,N_49788,N_49987);
xnor UO_572 (O_572,N_49919,N_49791);
nor UO_573 (O_573,N_49931,N_49987);
or UO_574 (O_574,N_49792,N_49794);
xor UO_575 (O_575,N_49865,N_49887);
and UO_576 (O_576,N_49924,N_49828);
or UO_577 (O_577,N_49750,N_49927);
and UO_578 (O_578,N_49902,N_49762);
and UO_579 (O_579,N_49967,N_49885);
or UO_580 (O_580,N_49968,N_49922);
and UO_581 (O_581,N_49833,N_49879);
nand UO_582 (O_582,N_49998,N_49809);
nor UO_583 (O_583,N_49837,N_49919);
and UO_584 (O_584,N_49844,N_49887);
xnor UO_585 (O_585,N_49913,N_49920);
xor UO_586 (O_586,N_49808,N_49813);
xnor UO_587 (O_587,N_49769,N_49783);
or UO_588 (O_588,N_49968,N_49903);
xor UO_589 (O_589,N_49786,N_49970);
xnor UO_590 (O_590,N_49813,N_49850);
xor UO_591 (O_591,N_49808,N_49773);
nand UO_592 (O_592,N_49921,N_49935);
and UO_593 (O_593,N_49968,N_49810);
nor UO_594 (O_594,N_49854,N_49943);
xor UO_595 (O_595,N_49950,N_49808);
nor UO_596 (O_596,N_49870,N_49859);
nor UO_597 (O_597,N_49918,N_49933);
or UO_598 (O_598,N_49850,N_49795);
nand UO_599 (O_599,N_49846,N_49885);
nand UO_600 (O_600,N_49792,N_49871);
and UO_601 (O_601,N_49810,N_49821);
nand UO_602 (O_602,N_49966,N_49840);
nor UO_603 (O_603,N_49873,N_49792);
or UO_604 (O_604,N_49929,N_49908);
nand UO_605 (O_605,N_49771,N_49825);
and UO_606 (O_606,N_49998,N_49893);
or UO_607 (O_607,N_49901,N_49942);
or UO_608 (O_608,N_49860,N_49898);
or UO_609 (O_609,N_49812,N_49938);
or UO_610 (O_610,N_49786,N_49895);
or UO_611 (O_611,N_49951,N_49795);
xnor UO_612 (O_612,N_49779,N_49825);
and UO_613 (O_613,N_49909,N_49817);
nor UO_614 (O_614,N_49763,N_49995);
nand UO_615 (O_615,N_49837,N_49935);
nor UO_616 (O_616,N_49946,N_49926);
or UO_617 (O_617,N_49874,N_49917);
nand UO_618 (O_618,N_49929,N_49903);
and UO_619 (O_619,N_49985,N_49961);
xor UO_620 (O_620,N_49993,N_49946);
nor UO_621 (O_621,N_49881,N_49896);
and UO_622 (O_622,N_49771,N_49812);
and UO_623 (O_623,N_49818,N_49768);
or UO_624 (O_624,N_49865,N_49882);
and UO_625 (O_625,N_49752,N_49946);
nand UO_626 (O_626,N_49780,N_49773);
nor UO_627 (O_627,N_49900,N_49864);
nand UO_628 (O_628,N_49821,N_49925);
xnor UO_629 (O_629,N_49819,N_49874);
or UO_630 (O_630,N_49966,N_49876);
nand UO_631 (O_631,N_49953,N_49922);
and UO_632 (O_632,N_49764,N_49944);
nand UO_633 (O_633,N_49869,N_49783);
nand UO_634 (O_634,N_49834,N_49976);
and UO_635 (O_635,N_49797,N_49957);
and UO_636 (O_636,N_49929,N_49774);
and UO_637 (O_637,N_49760,N_49997);
and UO_638 (O_638,N_49927,N_49873);
nand UO_639 (O_639,N_49826,N_49884);
nand UO_640 (O_640,N_49861,N_49904);
xor UO_641 (O_641,N_49797,N_49955);
xnor UO_642 (O_642,N_49851,N_49784);
or UO_643 (O_643,N_49775,N_49954);
xor UO_644 (O_644,N_49905,N_49950);
nor UO_645 (O_645,N_49877,N_49923);
nor UO_646 (O_646,N_49997,N_49972);
or UO_647 (O_647,N_49877,N_49957);
xor UO_648 (O_648,N_49790,N_49878);
nand UO_649 (O_649,N_49868,N_49881);
nor UO_650 (O_650,N_49815,N_49752);
and UO_651 (O_651,N_49887,N_49869);
or UO_652 (O_652,N_49856,N_49972);
or UO_653 (O_653,N_49875,N_49870);
and UO_654 (O_654,N_49831,N_49916);
nand UO_655 (O_655,N_49915,N_49969);
nor UO_656 (O_656,N_49925,N_49931);
nand UO_657 (O_657,N_49957,N_49783);
nand UO_658 (O_658,N_49951,N_49977);
xnor UO_659 (O_659,N_49952,N_49812);
or UO_660 (O_660,N_49918,N_49972);
nor UO_661 (O_661,N_49907,N_49819);
and UO_662 (O_662,N_49902,N_49825);
and UO_663 (O_663,N_49826,N_49758);
nand UO_664 (O_664,N_49781,N_49926);
xnor UO_665 (O_665,N_49926,N_49827);
nor UO_666 (O_666,N_49860,N_49966);
nand UO_667 (O_667,N_49852,N_49754);
and UO_668 (O_668,N_49949,N_49974);
xor UO_669 (O_669,N_49842,N_49775);
nor UO_670 (O_670,N_49915,N_49863);
nand UO_671 (O_671,N_49921,N_49871);
xnor UO_672 (O_672,N_49948,N_49874);
nor UO_673 (O_673,N_49954,N_49993);
nor UO_674 (O_674,N_49961,N_49792);
xnor UO_675 (O_675,N_49825,N_49959);
xor UO_676 (O_676,N_49954,N_49790);
nand UO_677 (O_677,N_49939,N_49976);
xnor UO_678 (O_678,N_49809,N_49876);
and UO_679 (O_679,N_49975,N_49971);
nor UO_680 (O_680,N_49823,N_49841);
and UO_681 (O_681,N_49918,N_49797);
nor UO_682 (O_682,N_49963,N_49955);
and UO_683 (O_683,N_49801,N_49862);
nand UO_684 (O_684,N_49807,N_49837);
and UO_685 (O_685,N_49917,N_49906);
nand UO_686 (O_686,N_49867,N_49765);
and UO_687 (O_687,N_49833,N_49959);
xor UO_688 (O_688,N_49967,N_49827);
nand UO_689 (O_689,N_49796,N_49780);
nand UO_690 (O_690,N_49866,N_49996);
xnor UO_691 (O_691,N_49868,N_49911);
nor UO_692 (O_692,N_49987,N_49756);
or UO_693 (O_693,N_49885,N_49893);
and UO_694 (O_694,N_49932,N_49836);
or UO_695 (O_695,N_49972,N_49911);
nand UO_696 (O_696,N_49810,N_49934);
or UO_697 (O_697,N_49770,N_49909);
or UO_698 (O_698,N_49988,N_49906);
nor UO_699 (O_699,N_49875,N_49993);
or UO_700 (O_700,N_49917,N_49809);
nand UO_701 (O_701,N_49841,N_49931);
nand UO_702 (O_702,N_49986,N_49805);
xor UO_703 (O_703,N_49763,N_49800);
and UO_704 (O_704,N_49819,N_49784);
xnor UO_705 (O_705,N_49988,N_49997);
nor UO_706 (O_706,N_49980,N_49841);
nor UO_707 (O_707,N_49940,N_49810);
and UO_708 (O_708,N_49931,N_49902);
nand UO_709 (O_709,N_49812,N_49824);
or UO_710 (O_710,N_49892,N_49849);
nor UO_711 (O_711,N_49835,N_49948);
and UO_712 (O_712,N_49917,N_49892);
nand UO_713 (O_713,N_49752,N_49817);
xor UO_714 (O_714,N_49765,N_49795);
xor UO_715 (O_715,N_49834,N_49856);
and UO_716 (O_716,N_49761,N_49988);
nor UO_717 (O_717,N_49860,N_49774);
nor UO_718 (O_718,N_49769,N_49961);
nand UO_719 (O_719,N_49824,N_49760);
xor UO_720 (O_720,N_49854,N_49758);
xor UO_721 (O_721,N_49965,N_49941);
and UO_722 (O_722,N_49882,N_49982);
and UO_723 (O_723,N_49953,N_49927);
nand UO_724 (O_724,N_49817,N_49981);
nand UO_725 (O_725,N_49784,N_49877);
xor UO_726 (O_726,N_49788,N_49809);
nand UO_727 (O_727,N_49844,N_49919);
xor UO_728 (O_728,N_49998,N_49775);
and UO_729 (O_729,N_49986,N_49829);
or UO_730 (O_730,N_49806,N_49977);
nand UO_731 (O_731,N_49792,N_49944);
xor UO_732 (O_732,N_49925,N_49945);
nor UO_733 (O_733,N_49845,N_49859);
xnor UO_734 (O_734,N_49835,N_49785);
and UO_735 (O_735,N_49756,N_49957);
nand UO_736 (O_736,N_49879,N_49834);
nand UO_737 (O_737,N_49842,N_49947);
or UO_738 (O_738,N_49914,N_49795);
xor UO_739 (O_739,N_49762,N_49941);
nand UO_740 (O_740,N_49773,N_49757);
nor UO_741 (O_741,N_49752,N_49906);
nand UO_742 (O_742,N_49836,N_49817);
and UO_743 (O_743,N_49811,N_49870);
or UO_744 (O_744,N_49777,N_49870);
nand UO_745 (O_745,N_49828,N_49952);
and UO_746 (O_746,N_49869,N_49849);
nand UO_747 (O_747,N_49950,N_49816);
and UO_748 (O_748,N_49811,N_49909);
or UO_749 (O_749,N_49932,N_49906);
and UO_750 (O_750,N_49940,N_49953);
nand UO_751 (O_751,N_49770,N_49808);
nor UO_752 (O_752,N_49999,N_49957);
and UO_753 (O_753,N_49847,N_49988);
and UO_754 (O_754,N_49987,N_49833);
or UO_755 (O_755,N_49872,N_49808);
or UO_756 (O_756,N_49800,N_49964);
and UO_757 (O_757,N_49796,N_49853);
and UO_758 (O_758,N_49844,N_49831);
nand UO_759 (O_759,N_49932,N_49992);
nor UO_760 (O_760,N_49956,N_49968);
nor UO_761 (O_761,N_49827,N_49982);
and UO_762 (O_762,N_49775,N_49905);
and UO_763 (O_763,N_49841,N_49754);
nand UO_764 (O_764,N_49889,N_49950);
nor UO_765 (O_765,N_49827,N_49774);
and UO_766 (O_766,N_49900,N_49804);
xnor UO_767 (O_767,N_49752,N_49985);
or UO_768 (O_768,N_49975,N_49876);
or UO_769 (O_769,N_49940,N_49751);
and UO_770 (O_770,N_49859,N_49897);
xnor UO_771 (O_771,N_49877,N_49843);
nand UO_772 (O_772,N_49913,N_49966);
and UO_773 (O_773,N_49842,N_49799);
nor UO_774 (O_774,N_49963,N_49870);
nor UO_775 (O_775,N_49818,N_49801);
nor UO_776 (O_776,N_49915,N_49789);
xor UO_777 (O_777,N_49960,N_49771);
or UO_778 (O_778,N_49963,N_49860);
xor UO_779 (O_779,N_49979,N_49750);
and UO_780 (O_780,N_49976,N_49752);
nand UO_781 (O_781,N_49841,N_49807);
xnor UO_782 (O_782,N_49791,N_49984);
and UO_783 (O_783,N_49812,N_49807);
or UO_784 (O_784,N_49980,N_49781);
xnor UO_785 (O_785,N_49919,N_49942);
nor UO_786 (O_786,N_49965,N_49786);
xor UO_787 (O_787,N_49885,N_49827);
nor UO_788 (O_788,N_49963,N_49916);
xnor UO_789 (O_789,N_49754,N_49984);
and UO_790 (O_790,N_49957,N_49890);
nor UO_791 (O_791,N_49872,N_49998);
nor UO_792 (O_792,N_49915,N_49870);
or UO_793 (O_793,N_49837,N_49963);
nor UO_794 (O_794,N_49923,N_49963);
xnor UO_795 (O_795,N_49994,N_49835);
nor UO_796 (O_796,N_49877,N_49904);
and UO_797 (O_797,N_49925,N_49877);
nor UO_798 (O_798,N_49953,N_49890);
xor UO_799 (O_799,N_49812,N_49873);
and UO_800 (O_800,N_49988,N_49775);
or UO_801 (O_801,N_49992,N_49938);
nand UO_802 (O_802,N_49953,N_49998);
nand UO_803 (O_803,N_49902,N_49750);
nand UO_804 (O_804,N_49833,N_49913);
nand UO_805 (O_805,N_49963,N_49982);
and UO_806 (O_806,N_49928,N_49776);
or UO_807 (O_807,N_49995,N_49969);
and UO_808 (O_808,N_49889,N_49859);
nor UO_809 (O_809,N_49813,N_49972);
or UO_810 (O_810,N_49990,N_49848);
xnor UO_811 (O_811,N_49918,N_49788);
nand UO_812 (O_812,N_49866,N_49963);
or UO_813 (O_813,N_49991,N_49756);
xor UO_814 (O_814,N_49933,N_49871);
and UO_815 (O_815,N_49848,N_49935);
nand UO_816 (O_816,N_49755,N_49980);
or UO_817 (O_817,N_49902,N_49987);
and UO_818 (O_818,N_49786,N_49767);
nand UO_819 (O_819,N_49782,N_49888);
and UO_820 (O_820,N_49835,N_49899);
and UO_821 (O_821,N_49974,N_49813);
and UO_822 (O_822,N_49990,N_49930);
or UO_823 (O_823,N_49822,N_49802);
nand UO_824 (O_824,N_49949,N_49854);
or UO_825 (O_825,N_49770,N_49771);
and UO_826 (O_826,N_49775,N_49808);
nor UO_827 (O_827,N_49922,N_49801);
or UO_828 (O_828,N_49861,N_49923);
xnor UO_829 (O_829,N_49850,N_49985);
nand UO_830 (O_830,N_49756,N_49915);
and UO_831 (O_831,N_49865,N_49954);
or UO_832 (O_832,N_49955,N_49869);
or UO_833 (O_833,N_49970,N_49778);
xor UO_834 (O_834,N_49865,N_49950);
or UO_835 (O_835,N_49818,N_49937);
nand UO_836 (O_836,N_49937,N_49803);
or UO_837 (O_837,N_49985,N_49805);
nand UO_838 (O_838,N_49963,N_49954);
nor UO_839 (O_839,N_49781,N_49792);
or UO_840 (O_840,N_49803,N_49965);
xor UO_841 (O_841,N_49790,N_49799);
nor UO_842 (O_842,N_49805,N_49929);
nor UO_843 (O_843,N_49904,N_49999);
nor UO_844 (O_844,N_49923,N_49821);
xor UO_845 (O_845,N_49996,N_49753);
nand UO_846 (O_846,N_49809,N_49997);
nand UO_847 (O_847,N_49796,N_49998);
nand UO_848 (O_848,N_49828,N_49961);
nor UO_849 (O_849,N_49919,N_49864);
and UO_850 (O_850,N_49753,N_49941);
and UO_851 (O_851,N_49909,N_49785);
xnor UO_852 (O_852,N_49916,N_49786);
nor UO_853 (O_853,N_49760,N_49790);
xnor UO_854 (O_854,N_49941,N_49943);
nand UO_855 (O_855,N_49907,N_49902);
or UO_856 (O_856,N_49951,N_49985);
or UO_857 (O_857,N_49931,N_49763);
and UO_858 (O_858,N_49777,N_49794);
nand UO_859 (O_859,N_49928,N_49760);
xnor UO_860 (O_860,N_49923,N_49952);
and UO_861 (O_861,N_49934,N_49827);
and UO_862 (O_862,N_49804,N_49984);
xnor UO_863 (O_863,N_49766,N_49852);
nand UO_864 (O_864,N_49948,N_49829);
and UO_865 (O_865,N_49843,N_49948);
xnor UO_866 (O_866,N_49862,N_49769);
xnor UO_867 (O_867,N_49863,N_49770);
or UO_868 (O_868,N_49867,N_49849);
nand UO_869 (O_869,N_49887,N_49892);
nor UO_870 (O_870,N_49762,N_49833);
nor UO_871 (O_871,N_49866,N_49980);
and UO_872 (O_872,N_49864,N_49789);
nor UO_873 (O_873,N_49794,N_49994);
nor UO_874 (O_874,N_49860,N_49768);
nand UO_875 (O_875,N_49936,N_49956);
nor UO_876 (O_876,N_49994,N_49750);
and UO_877 (O_877,N_49770,N_49819);
nor UO_878 (O_878,N_49972,N_49842);
and UO_879 (O_879,N_49869,N_49908);
and UO_880 (O_880,N_49992,N_49826);
and UO_881 (O_881,N_49894,N_49780);
or UO_882 (O_882,N_49843,N_49857);
and UO_883 (O_883,N_49841,N_49945);
xnor UO_884 (O_884,N_49808,N_49835);
nand UO_885 (O_885,N_49777,N_49909);
xnor UO_886 (O_886,N_49830,N_49873);
xnor UO_887 (O_887,N_49925,N_49816);
nor UO_888 (O_888,N_49887,N_49963);
nand UO_889 (O_889,N_49981,N_49785);
or UO_890 (O_890,N_49893,N_49929);
xnor UO_891 (O_891,N_49909,N_49794);
nand UO_892 (O_892,N_49857,N_49817);
nor UO_893 (O_893,N_49834,N_49862);
and UO_894 (O_894,N_49970,N_49916);
and UO_895 (O_895,N_49787,N_49753);
and UO_896 (O_896,N_49769,N_49993);
nor UO_897 (O_897,N_49867,N_49937);
or UO_898 (O_898,N_49849,N_49750);
and UO_899 (O_899,N_49834,N_49761);
nand UO_900 (O_900,N_49764,N_49798);
nor UO_901 (O_901,N_49903,N_49896);
nor UO_902 (O_902,N_49905,N_49853);
and UO_903 (O_903,N_49995,N_49866);
nor UO_904 (O_904,N_49998,N_49807);
and UO_905 (O_905,N_49882,N_49968);
xor UO_906 (O_906,N_49952,N_49988);
nor UO_907 (O_907,N_49786,N_49991);
xor UO_908 (O_908,N_49754,N_49768);
and UO_909 (O_909,N_49861,N_49901);
and UO_910 (O_910,N_49892,N_49899);
nand UO_911 (O_911,N_49796,N_49912);
or UO_912 (O_912,N_49881,N_49794);
nand UO_913 (O_913,N_49954,N_49943);
or UO_914 (O_914,N_49777,N_49967);
nor UO_915 (O_915,N_49930,N_49928);
and UO_916 (O_916,N_49850,N_49826);
nor UO_917 (O_917,N_49873,N_49770);
xnor UO_918 (O_918,N_49806,N_49818);
xor UO_919 (O_919,N_49766,N_49860);
and UO_920 (O_920,N_49885,N_49932);
and UO_921 (O_921,N_49939,N_49952);
and UO_922 (O_922,N_49985,N_49959);
and UO_923 (O_923,N_49936,N_49909);
and UO_924 (O_924,N_49877,N_49754);
nand UO_925 (O_925,N_49806,N_49881);
nor UO_926 (O_926,N_49910,N_49859);
xnor UO_927 (O_927,N_49801,N_49930);
nor UO_928 (O_928,N_49836,N_49889);
and UO_929 (O_929,N_49780,N_49917);
or UO_930 (O_930,N_49838,N_49900);
or UO_931 (O_931,N_49917,N_49784);
xor UO_932 (O_932,N_49940,N_49898);
or UO_933 (O_933,N_49994,N_49808);
nor UO_934 (O_934,N_49863,N_49816);
xnor UO_935 (O_935,N_49882,N_49814);
nand UO_936 (O_936,N_49916,N_49891);
xor UO_937 (O_937,N_49759,N_49993);
and UO_938 (O_938,N_49893,N_49837);
or UO_939 (O_939,N_49932,N_49829);
nor UO_940 (O_940,N_49812,N_49918);
and UO_941 (O_941,N_49935,N_49813);
and UO_942 (O_942,N_49971,N_49943);
or UO_943 (O_943,N_49769,N_49952);
or UO_944 (O_944,N_49791,N_49993);
or UO_945 (O_945,N_49924,N_49835);
nand UO_946 (O_946,N_49766,N_49764);
xor UO_947 (O_947,N_49880,N_49917);
xor UO_948 (O_948,N_49991,N_49757);
nand UO_949 (O_949,N_49977,N_49855);
nor UO_950 (O_950,N_49967,N_49893);
nand UO_951 (O_951,N_49858,N_49953);
nand UO_952 (O_952,N_49819,N_49976);
or UO_953 (O_953,N_49828,N_49975);
xnor UO_954 (O_954,N_49788,N_49980);
nand UO_955 (O_955,N_49816,N_49811);
nand UO_956 (O_956,N_49919,N_49772);
nor UO_957 (O_957,N_49879,N_49751);
or UO_958 (O_958,N_49876,N_49921);
nor UO_959 (O_959,N_49958,N_49785);
nand UO_960 (O_960,N_49843,N_49995);
nor UO_961 (O_961,N_49932,N_49830);
or UO_962 (O_962,N_49958,N_49848);
nor UO_963 (O_963,N_49881,N_49752);
nand UO_964 (O_964,N_49858,N_49784);
nand UO_965 (O_965,N_49997,N_49805);
or UO_966 (O_966,N_49811,N_49805);
and UO_967 (O_967,N_49855,N_49926);
nor UO_968 (O_968,N_49760,N_49809);
or UO_969 (O_969,N_49843,N_49926);
nand UO_970 (O_970,N_49860,N_49905);
or UO_971 (O_971,N_49987,N_49832);
and UO_972 (O_972,N_49849,N_49945);
xnor UO_973 (O_973,N_49856,N_49927);
or UO_974 (O_974,N_49987,N_49794);
and UO_975 (O_975,N_49805,N_49907);
xor UO_976 (O_976,N_49836,N_49866);
xnor UO_977 (O_977,N_49981,N_49802);
xor UO_978 (O_978,N_49911,N_49903);
nand UO_979 (O_979,N_49838,N_49768);
and UO_980 (O_980,N_49872,N_49953);
nor UO_981 (O_981,N_49751,N_49795);
and UO_982 (O_982,N_49967,N_49911);
or UO_983 (O_983,N_49867,N_49932);
or UO_984 (O_984,N_49770,N_49790);
or UO_985 (O_985,N_49793,N_49847);
or UO_986 (O_986,N_49959,N_49899);
or UO_987 (O_987,N_49984,N_49904);
or UO_988 (O_988,N_49833,N_49843);
nor UO_989 (O_989,N_49786,N_49920);
or UO_990 (O_990,N_49894,N_49983);
and UO_991 (O_991,N_49821,N_49978);
and UO_992 (O_992,N_49960,N_49954);
nand UO_993 (O_993,N_49778,N_49893);
nand UO_994 (O_994,N_49916,N_49930);
or UO_995 (O_995,N_49861,N_49849);
and UO_996 (O_996,N_49842,N_49899);
or UO_997 (O_997,N_49960,N_49830);
or UO_998 (O_998,N_49762,N_49921);
xor UO_999 (O_999,N_49753,N_49986);
and UO_1000 (O_1000,N_49987,N_49908);
nand UO_1001 (O_1001,N_49802,N_49840);
and UO_1002 (O_1002,N_49935,N_49916);
and UO_1003 (O_1003,N_49950,N_49976);
and UO_1004 (O_1004,N_49834,N_49934);
and UO_1005 (O_1005,N_49819,N_49830);
or UO_1006 (O_1006,N_49872,N_49844);
and UO_1007 (O_1007,N_49947,N_49937);
xor UO_1008 (O_1008,N_49886,N_49933);
nand UO_1009 (O_1009,N_49778,N_49849);
xnor UO_1010 (O_1010,N_49944,N_49794);
or UO_1011 (O_1011,N_49979,N_49850);
nor UO_1012 (O_1012,N_49968,N_49913);
nor UO_1013 (O_1013,N_49895,N_49904);
nor UO_1014 (O_1014,N_49979,N_49972);
or UO_1015 (O_1015,N_49958,N_49980);
nand UO_1016 (O_1016,N_49903,N_49937);
or UO_1017 (O_1017,N_49756,N_49997);
or UO_1018 (O_1018,N_49922,N_49888);
xor UO_1019 (O_1019,N_49931,N_49839);
nand UO_1020 (O_1020,N_49986,N_49841);
nand UO_1021 (O_1021,N_49975,N_49813);
nor UO_1022 (O_1022,N_49794,N_49793);
nor UO_1023 (O_1023,N_49755,N_49967);
or UO_1024 (O_1024,N_49830,N_49959);
nor UO_1025 (O_1025,N_49950,N_49902);
nand UO_1026 (O_1026,N_49790,N_49839);
nor UO_1027 (O_1027,N_49948,N_49753);
nor UO_1028 (O_1028,N_49795,N_49763);
nor UO_1029 (O_1029,N_49839,N_49973);
xnor UO_1030 (O_1030,N_49811,N_49822);
xor UO_1031 (O_1031,N_49891,N_49833);
xnor UO_1032 (O_1032,N_49986,N_49869);
and UO_1033 (O_1033,N_49860,N_49999);
xor UO_1034 (O_1034,N_49894,N_49911);
or UO_1035 (O_1035,N_49861,N_49966);
or UO_1036 (O_1036,N_49957,N_49782);
xor UO_1037 (O_1037,N_49773,N_49817);
and UO_1038 (O_1038,N_49814,N_49984);
and UO_1039 (O_1039,N_49970,N_49801);
nand UO_1040 (O_1040,N_49813,N_49995);
nor UO_1041 (O_1041,N_49773,N_49810);
nor UO_1042 (O_1042,N_49829,N_49893);
nor UO_1043 (O_1043,N_49772,N_49836);
xor UO_1044 (O_1044,N_49838,N_49840);
nor UO_1045 (O_1045,N_49974,N_49954);
xor UO_1046 (O_1046,N_49983,N_49775);
nor UO_1047 (O_1047,N_49979,N_49898);
nor UO_1048 (O_1048,N_49915,N_49958);
nor UO_1049 (O_1049,N_49862,N_49836);
nor UO_1050 (O_1050,N_49858,N_49996);
or UO_1051 (O_1051,N_49974,N_49844);
xnor UO_1052 (O_1052,N_49789,N_49978);
nor UO_1053 (O_1053,N_49774,N_49879);
nor UO_1054 (O_1054,N_49855,N_49853);
nor UO_1055 (O_1055,N_49836,N_49907);
nor UO_1056 (O_1056,N_49828,N_49882);
nand UO_1057 (O_1057,N_49953,N_49974);
nand UO_1058 (O_1058,N_49978,N_49823);
xnor UO_1059 (O_1059,N_49822,N_49799);
or UO_1060 (O_1060,N_49806,N_49998);
or UO_1061 (O_1061,N_49891,N_49920);
and UO_1062 (O_1062,N_49968,N_49997);
xor UO_1063 (O_1063,N_49793,N_49824);
or UO_1064 (O_1064,N_49815,N_49810);
xnor UO_1065 (O_1065,N_49806,N_49969);
and UO_1066 (O_1066,N_49754,N_49968);
and UO_1067 (O_1067,N_49773,N_49929);
xnor UO_1068 (O_1068,N_49802,N_49884);
xor UO_1069 (O_1069,N_49787,N_49832);
xnor UO_1070 (O_1070,N_49926,N_49917);
xnor UO_1071 (O_1071,N_49893,N_49945);
nand UO_1072 (O_1072,N_49945,N_49797);
nor UO_1073 (O_1073,N_49888,N_49822);
or UO_1074 (O_1074,N_49856,N_49963);
or UO_1075 (O_1075,N_49832,N_49982);
nand UO_1076 (O_1076,N_49823,N_49994);
or UO_1077 (O_1077,N_49895,N_49794);
and UO_1078 (O_1078,N_49853,N_49774);
nor UO_1079 (O_1079,N_49888,N_49837);
nand UO_1080 (O_1080,N_49933,N_49963);
or UO_1081 (O_1081,N_49937,N_49949);
nor UO_1082 (O_1082,N_49898,N_49798);
and UO_1083 (O_1083,N_49883,N_49852);
nand UO_1084 (O_1084,N_49843,N_49802);
nand UO_1085 (O_1085,N_49982,N_49969);
nand UO_1086 (O_1086,N_49805,N_49840);
or UO_1087 (O_1087,N_49940,N_49813);
and UO_1088 (O_1088,N_49963,N_49798);
xnor UO_1089 (O_1089,N_49918,N_49920);
nand UO_1090 (O_1090,N_49782,N_49780);
and UO_1091 (O_1091,N_49774,N_49943);
nand UO_1092 (O_1092,N_49925,N_49794);
or UO_1093 (O_1093,N_49858,N_49919);
nor UO_1094 (O_1094,N_49860,N_49935);
nand UO_1095 (O_1095,N_49814,N_49991);
or UO_1096 (O_1096,N_49915,N_49775);
nand UO_1097 (O_1097,N_49834,N_49776);
or UO_1098 (O_1098,N_49961,N_49805);
or UO_1099 (O_1099,N_49852,N_49805);
and UO_1100 (O_1100,N_49847,N_49915);
or UO_1101 (O_1101,N_49918,N_49911);
or UO_1102 (O_1102,N_49857,N_49768);
and UO_1103 (O_1103,N_49819,N_49757);
nand UO_1104 (O_1104,N_49884,N_49768);
or UO_1105 (O_1105,N_49925,N_49788);
nor UO_1106 (O_1106,N_49985,N_49823);
xnor UO_1107 (O_1107,N_49815,N_49869);
and UO_1108 (O_1108,N_49874,N_49925);
xor UO_1109 (O_1109,N_49846,N_49973);
nand UO_1110 (O_1110,N_49907,N_49969);
xor UO_1111 (O_1111,N_49999,N_49965);
xor UO_1112 (O_1112,N_49998,N_49958);
and UO_1113 (O_1113,N_49871,N_49801);
xnor UO_1114 (O_1114,N_49930,N_49837);
nor UO_1115 (O_1115,N_49974,N_49931);
nor UO_1116 (O_1116,N_49794,N_49963);
nand UO_1117 (O_1117,N_49961,N_49959);
xor UO_1118 (O_1118,N_49956,N_49833);
or UO_1119 (O_1119,N_49801,N_49940);
or UO_1120 (O_1120,N_49811,N_49941);
xnor UO_1121 (O_1121,N_49939,N_49783);
xor UO_1122 (O_1122,N_49975,N_49850);
and UO_1123 (O_1123,N_49829,N_49920);
or UO_1124 (O_1124,N_49772,N_49976);
or UO_1125 (O_1125,N_49935,N_49786);
nand UO_1126 (O_1126,N_49793,N_49831);
or UO_1127 (O_1127,N_49871,N_49822);
and UO_1128 (O_1128,N_49800,N_49899);
nand UO_1129 (O_1129,N_49783,N_49904);
xnor UO_1130 (O_1130,N_49934,N_49872);
nand UO_1131 (O_1131,N_49828,N_49877);
and UO_1132 (O_1132,N_49951,N_49828);
nor UO_1133 (O_1133,N_49956,N_49826);
xnor UO_1134 (O_1134,N_49861,N_49853);
or UO_1135 (O_1135,N_49925,N_49969);
nor UO_1136 (O_1136,N_49935,N_49787);
and UO_1137 (O_1137,N_49795,N_49917);
nand UO_1138 (O_1138,N_49908,N_49874);
or UO_1139 (O_1139,N_49902,N_49838);
nor UO_1140 (O_1140,N_49776,N_49917);
nand UO_1141 (O_1141,N_49966,N_49809);
or UO_1142 (O_1142,N_49967,N_49805);
and UO_1143 (O_1143,N_49867,N_49805);
and UO_1144 (O_1144,N_49847,N_49853);
nand UO_1145 (O_1145,N_49796,N_49900);
nand UO_1146 (O_1146,N_49760,N_49843);
nor UO_1147 (O_1147,N_49980,N_49922);
nand UO_1148 (O_1148,N_49937,N_49982);
nand UO_1149 (O_1149,N_49893,N_49955);
nand UO_1150 (O_1150,N_49774,N_49918);
or UO_1151 (O_1151,N_49842,N_49846);
or UO_1152 (O_1152,N_49791,N_49831);
and UO_1153 (O_1153,N_49898,N_49830);
nor UO_1154 (O_1154,N_49866,N_49798);
nor UO_1155 (O_1155,N_49809,N_49937);
and UO_1156 (O_1156,N_49790,N_49974);
and UO_1157 (O_1157,N_49993,N_49862);
nand UO_1158 (O_1158,N_49760,N_49962);
or UO_1159 (O_1159,N_49806,N_49880);
or UO_1160 (O_1160,N_49841,N_49871);
xor UO_1161 (O_1161,N_49928,N_49885);
or UO_1162 (O_1162,N_49944,N_49992);
or UO_1163 (O_1163,N_49977,N_49975);
xor UO_1164 (O_1164,N_49988,N_49829);
xnor UO_1165 (O_1165,N_49817,N_49867);
nand UO_1166 (O_1166,N_49963,N_49959);
xnor UO_1167 (O_1167,N_49944,N_49784);
or UO_1168 (O_1168,N_49971,N_49809);
xor UO_1169 (O_1169,N_49939,N_49838);
nand UO_1170 (O_1170,N_49816,N_49806);
nor UO_1171 (O_1171,N_49986,N_49920);
nand UO_1172 (O_1172,N_49778,N_49757);
nor UO_1173 (O_1173,N_49751,N_49884);
and UO_1174 (O_1174,N_49828,N_49779);
or UO_1175 (O_1175,N_49753,N_49855);
or UO_1176 (O_1176,N_49908,N_49899);
and UO_1177 (O_1177,N_49877,N_49802);
and UO_1178 (O_1178,N_49912,N_49797);
nor UO_1179 (O_1179,N_49873,N_49971);
or UO_1180 (O_1180,N_49769,N_49851);
xor UO_1181 (O_1181,N_49823,N_49853);
xnor UO_1182 (O_1182,N_49909,N_49810);
xor UO_1183 (O_1183,N_49974,N_49771);
nand UO_1184 (O_1184,N_49807,N_49959);
nand UO_1185 (O_1185,N_49989,N_49908);
nand UO_1186 (O_1186,N_49894,N_49872);
nor UO_1187 (O_1187,N_49900,N_49801);
xor UO_1188 (O_1188,N_49851,N_49888);
or UO_1189 (O_1189,N_49878,N_49876);
nor UO_1190 (O_1190,N_49859,N_49963);
or UO_1191 (O_1191,N_49838,N_49937);
nor UO_1192 (O_1192,N_49786,N_49891);
xor UO_1193 (O_1193,N_49994,N_49890);
xor UO_1194 (O_1194,N_49975,N_49776);
xnor UO_1195 (O_1195,N_49825,N_49962);
xnor UO_1196 (O_1196,N_49930,N_49895);
or UO_1197 (O_1197,N_49776,N_49907);
nand UO_1198 (O_1198,N_49761,N_49991);
nor UO_1199 (O_1199,N_49992,N_49852);
nor UO_1200 (O_1200,N_49920,N_49756);
nand UO_1201 (O_1201,N_49964,N_49820);
or UO_1202 (O_1202,N_49802,N_49867);
or UO_1203 (O_1203,N_49835,N_49983);
nor UO_1204 (O_1204,N_49918,N_49798);
and UO_1205 (O_1205,N_49925,N_49762);
xnor UO_1206 (O_1206,N_49940,N_49802);
and UO_1207 (O_1207,N_49931,N_49801);
nor UO_1208 (O_1208,N_49792,N_49809);
xnor UO_1209 (O_1209,N_49940,N_49959);
nor UO_1210 (O_1210,N_49822,N_49917);
nor UO_1211 (O_1211,N_49781,N_49831);
and UO_1212 (O_1212,N_49868,N_49934);
nand UO_1213 (O_1213,N_49805,N_49990);
xnor UO_1214 (O_1214,N_49882,N_49927);
nor UO_1215 (O_1215,N_49754,N_49961);
xor UO_1216 (O_1216,N_49832,N_49999);
nor UO_1217 (O_1217,N_49946,N_49999);
xor UO_1218 (O_1218,N_49852,N_49966);
nor UO_1219 (O_1219,N_49830,N_49951);
xor UO_1220 (O_1220,N_49902,N_49884);
xor UO_1221 (O_1221,N_49812,N_49944);
nand UO_1222 (O_1222,N_49903,N_49919);
and UO_1223 (O_1223,N_49861,N_49978);
and UO_1224 (O_1224,N_49931,N_49907);
xor UO_1225 (O_1225,N_49882,N_49883);
and UO_1226 (O_1226,N_49760,N_49926);
nor UO_1227 (O_1227,N_49920,N_49988);
or UO_1228 (O_1228,N_49886,N_49757);
or UO_1229 (O_1229,N_49793,N_49920);
nand UO_1230 (O_1230,N_49842,N_49944);
nor UO_1231 (O_1231,N_49762,N_49755);
nand UO_1232 (O_1232,N_49886,N_49871);
nand UO_1233 (O_1233,N_49997,N_49900);
nand UO_1234 (O_1234,N_49946,N_49854);
and UO_1235 (O_1235,N_49832,N_49845);
xor UO_1236 (O_1236,N_49971,N_49801);
nor UO_1237 (O_1237,N_49932,N_49865);
xor UO_1238 (O_1238,N_49809,N_49850);
nor UO_1239 (O_1239,N_49757,N_49826);
or UO_1240 (O_1240,N_49784,N_49796);
xor UO_1241 (O_1241,N_49887,N_49988);
nand UO_1242 (O_1242,N_49781,N_49910);
and UO_1243 (O_1243,N_49957,N_49854);
xor UO_1244 (O_1244,N_49982,N_49812);
and UO_1245 (O_1245,N_49784,N_49939);
and UO_1246 (O_1246,N_49840,N_49780);
or UO_1247 (O_1247,N_49986,N_49908);
or UO_1248 (O_1248,N_49896,N_49850);
or UO_1249 (O_1249,N_49877,N_49973);
nor UO_1250 (O_1250,N_49988,N_49796);
nand UO_1251 (O_1251,N_49763,N_49924);
or UO_1252 (O_1252,N_49912,N_49872);
nor UO_1253 (O_1253,N_49875,N_49881);
or UO_1254 (O_1254,N_49900,N_49817);
nand UO_1255 (O_1255,N_49999,N_49761);
or UO_1256 (O_1256,N_49891,N_49923);
xor UO_1257 (O_1257,N_49996,N_49982);
nor UO_1258 (O_1258,N_49801,N_49756);
and UO_1259 (O_1259,N_49989,N_49964);
xor UO_1260 (O_1260,N_49825,N_49809);
nor UO_1261 (O_1261,N_49937,N_49925);
nor UO_1262 (O_1262,N_49967,N_49976);
nand UO_1263 (O_1263,N_49977,N_49895);
and UO_1264 (O_1264,N_49836,N_49788);
and UO_1265 (O_1265,N_49846,N_49876);
xor UO_1266 (O_1266,N_49889,N_49964);
xor UO_1267 (O_1267,N_49838,N_49940);
and UO_1268 (O_1268,N_49906,N_49826);
or UO_1269 (O_1269,N_49783,N_49948);
xor UO_1270 (O_1270,N_49979,N_49934);
or UO_1271 (O_1271,N_49763,N_49879);
nand UO_1272 (O_1272,N_49920,N_49990);
or UO_1273 (O_1273,N_49801,N_49868);
nand UO_1274 (O_1274,N_49979,N_49930);
nand UO_1275 (O_1275,N_49917,N_49752);
nor UO_1276 (O_1276,N_49862,N_49998);
and UO_1277 (O_1277,N_49818,N_49971);
nor UO_1278 (O_1278,N_49802,N_49957);
nor UO_1279 (O_1279,N_49795,N_49756);
and UO_1280 (O_1280,N_49835,N_49849);
xnor UO_1281 (O_1281,N_49832,N_49795);
nand UO_1282 (O_1282,N_49927,N_49917);
nor UO_1283 (O_1283,N_49785,N_49847);
xor UO_1284 (O_1284,N_49895,N_49853);
xor UO_1285 (O_1285,N_49960,N_49875);
xor UO_1286 (O_1286,N_49891,N_49876);
xor UO_1287 (O_1287,N_49998,N_49858);
xnor UO_1288 (O_1288,N_49891,N_49816);
or UO_1289 (O_1289,N_49776,N_49926);
nor UO_1290 (O_1290,N_49970,N_49816);
nor UO_1291 (O_1291,N_49977,N_49898);
or UO_1292 (O_1292,N_49783,N_49852);
xor UO_1293 (O_1293,N_49913,N_49941);
and UO_1294 (O_1294,N_49980,N_49952);
xnor UO_1295 (O_1295,N_49968,N_49914);
xor UO_1296 (O_1296,N_49914,N_49893);
xnor UO_1297 (O_1297,N_49944,N_49849);
nor UO_1298 (O_1298,N_49894,N_49874);
or UO_1299 (O_1299,N_49778,N_49859);
nor UO_1300 (O_1300,N_49758,N_49948);
xnor UO_1301 (O_1301,N_49798,N_49893);
xor UO_1302 (O_1302,N_49937,N_49946);
xor UO_1303 (O_1303,N_49851,N_49768);
nor UO_1304 (O_1304,N_49997,N_49865);
nand UO_1305 (O_1305,N_49982,N_49810);
and UO_1306 (O_1306,N_49929,N_49832);
nand UO_1307 (O_1307,N_49782,N_49816);
nor UO_1308 (O_1308,N_49876,N_49926);
xor UO_1309 (O_1309,N_49964,N_49895);
nor UO_1310 (O_1310,N_49758,N_49883);
xnor UO_1311 (O_1311,N_49866,N_49830);
or UO_1312 (O_1312,N_49779,N_49854);
xor UO_1313 (O_1313,N_49831,N_49897);
nor UO_1314 (O_1314,N_49846,N_49774);
nor UO_1315 (O_1315,N_49949,N_49994);
xnor UO_1316 (O_1316,N_49774,N_49759);
nand UO_1317 (O_1317,N_49942,N_49773);
and UO_1318 (O_1318,N_49851,N_49896);
nor UO_1319 (O_1319,N_49812,N_49808);
xor UO_1320 (O_1320,N_49817,N_49837);
nor UO_1321 (O_1321,N_49890,N_49940);
or UO_1322 (O_1322,N_49777,N_49854);
xnor UO_1323 (O_1323,N_49862,N_49925);
xnor UO_1324 (O_1324,N_49971,N_49933);
or UO_1325 (O_1325,N_49878,N_49817);
or UO_1326 (O_1326,N_49800,N_49840);
xor UO_1327 (O_1327,N_49983,N_49827);
nor UO_1328 (O_1328,N_49895,N_49821);
or UO_1329 (O_1329,N_49772,N_49754);
nand UO_1330 (O_1330,N_49826,N_49778);
or UO_1331 (O_1331,N_49950,N_49917);
and UO_1332 (O_1332,N_49762,N_49918);
or UO_1333 (O_1333,N_49986,N_49886);
nor UO_1334 (O_1334,N_49758,N_49769);
xor UO_1335 (O_1335,N_49930,N_49978);
and UO_1336 (O_1336,N_49947,N_49990);
or UO_1337 (O_1337,N_49988,N_49891);
or UO_1338 (O_1338,N_49963,N_49799);
nand UO_1339 (O_1339,N_49828,N_49900);
and UO_1340 (O_1340,N_49782,N_49962);
and UO_1341 (O_1341,N_49767,N_49876);
and UO_1342 (O_1342,N_49920,N_49989);
or UO_1343 (O_1343,N_49868,N_49781);
nand UO_1344 (O_1344,N_49784,N_49884);
nand UO_1345 (O_1345,N_49917,N_49912);
and UO_1346 (O_1346,N_49787,N_49985);
and UO_1347 (O_1347,N_49786,N_49838);
nand UO_1348 (O_1348,N_49876,N_49751);
and UO_1349 (O_1349,N_49860,N_49982);
and UO_1350 (O_1350,N_49909,N_49791);
and UO_1351 (O_1351,N_49787,N_49851);
nor UO_1352 (O_1352,N_49774,N_49819);
nand UO_1353 (O_1353,N_49929,N_49945);
xor UO_1354 (O_1354,N_49860,N_49769);
nand UO_1355 (O_1355,N_49811,N_49980);
nor UO_1356 (O_1356,N_49783,N_49925);
nand UO_1357 (O_1357,N_49850,N_49814);
xor UO_1358 (O_1358,N_49867,N_49824);
nor UO_1359 (O_1359,N_49882,N_49751);
nor UO_1360 (O_1360,N_49790,N_49959);
nor UO_1361 (O_1361,N_49969,N_49860);
nor UO_1362 (O_1362,N_49964,N_49875);
or UO_1363 (O_1363,N_49786,N_49932);
xor UO_1364 (O_1364,N_49847,N_49794);
xor UO_1365 (O_1365,N_49949,N_49969);
nand UO_1366 (O_1366,N_49892,N_49884);
xor UO_1367 (O_1367,N_49930,N_49795);
xnor UO_1368 (O_1368,N_49870,N_49934);
and UO_1369 (O_1369,N_49835,N_49767);
and UO_1370 (O_1370,N_49892,N_49912);
or UO_1371 (O_1371,N_49906,N_49929);
xor UO_1372 (O_1372,N_49840,N_49846);
or UO_1373 (O_1373,N_49944,N_49875);
and UO_1374 (O_1374,N_49951,N_49846);
xor UO_1375 (O_1375,N_49751,N_49798);
or UO_1376 (O_1376,N_49765,N_49879);
nor UO_1377 (O_1377,N_49928,N_49762);
xor UO_1378 (O_1378,N_49839,N_49758);
nand UO_1379 (O_1379,N_49916,N_49756);
xnor UO_1380 (O_1380,N_49890,N_49969);
nor UO_1381 (O_1381,N_49951,N_49753);
or UO_1382 (O_1382,N_49934,N_49901);
and UO_1383 (O_1383,N_49934,N_49997);
xor UO_1384 (O_1384,N_49776,N_49782);
and UO_1385 (O_1385,N_49844,N_49763);
xor UO_1386 (O_1386,N_49792,N_49949);
xnor UO_1387 (O_1387,N_49978,N_49890);
nor UO_1388 (O_1388,N_49897,N_49970);
xor UO_1389 (O_1389,N_49938,N_49780);
xnor UO_1390 (O_1390,N_49887,N_49795);
or UO_1391 (O_1391,N_49813,N_49885);
nor UO_1392 (O_1392,N_49826,N_49882);
nor UO_1393 (O_1393,N_49874,N_49980);
nor UO_1394 (O_1394,N_49920,N_49899);
xnor UO_1395 (O_1395,N_49933,N_49807);
or UO_1396 (O_1396,N_49914,N_49911);
or UO_1397 (O_1397,N_49843,N_49918);
nand UO_1398 (O_1398,N_49808,N_49920);
nor UO_1399 (O_1399,N_49851,N_49991);
nand UO_1400 (O_1400,N_49774,N_49848);
and UO_1401 (O_1401,N_49961,N_49901);
and UO_1402 (O_1402,N_49881,N_49830);
or UO_1403 (O_1403,N_49777,N_49954);
or UO_1404 (O_1404,N_49765,N_49904);
nor UO_1405 (O_1405,N_49849,N_49874);
nor UO_1406 (O_1406,N_49861,N_49970);
or UO_1407 (O_1407,N_49860,N_49779);
nor UO_1408 (O_1408,N_49944,N_49758);
xnor UO_1409 (O_1409,N_49908,N_49800);
nand UO_1410 (O_1410,N_49996,N_49775);
nor UO_1411 (O_1411,N_49781,N_49915);
nand UO_1412 (O_1412,N_49796,N_49999);
nor UO_1413 (O_1413,N_49986,N_49976);
xnor UO_1414 (O_1414,N_49924,N_49863);
xor UO_1415 (O_1415,N_49983,N_49934);
nor UO_1416 (O_1416,N_49755,N_49814);
or UO_1417 (O_1417,N_49821,N_49869);
and UO_1418 (O_1418,N_49901,N_49845);
or UO_1419 (O_1419,N_49974,N_49824);
nor UO_1420 (O_1420,N_49905,N_49948);
nor UO_1421 (O_1421,N_49795,N_49894);
or UO_1422 (O_1422,N_49847,N_49894);
nor UO_1423 (O_1423,N_49832,N_49993);
and UO_1424 (O_1424,N_49786,N_49919);
and UO_1425 (O_1425,N_49872,N_49863);
xor UO_1426 (O_1426,N_49999,N_49763);
and UO_1427 (O_1427,N_49843,N_49977);
and UO_1428 (O_1428,N_49983,N_49944);
nand UO_1429 (O_1429,N_49941,N_49976);
or UO_1430 (O_1430,N_49817,N_49995);
nor UO_1431 (O_1431,N_49995,N_49879);
or UO_1432 (O_1432,N_49928,N_49798);
xnor UO_1433 (O_1433,N_49767,N_49909);
nor UO_1434 (O_1434,N_49806,N_49885);
xor UO_1435 (O_1435,N_49772,N_49855);
nand UO_1436 (O_1436,N_49879,N_49801);
and UO_1437 (O_1437,N_49921,N_49788);
xnor UO_1438 (O_1438,N_49966,N_49975);
nand UO_1439 (O_1439,N_49765,N_49833);
and UO_1440 (O_1440,N_49841,N_49847);
and UO_1441 (O_1441,N_49849,N_49792);
xnor UO_1442 (O_1442,N_49969,N_49851);
and UO_1443 (O_1443,N_49801,N_49787);
nor UO_1444 (O_1444,N_49926,N_49849);
and UO_1445 (O_1445,N_49950,N_49915);
nor UO_1446 (O_1446,N_49753,N_49838);
xnor UO_1447 (O_1447,N_49768,N_49946);
or UO_1448 (O_1448,N_49895,N_49892);
and UO_1449 (O_1449,N_49793,N_49899);
nor UO_1450 (O_1450,N_49815,N_49936);
and UO_1451 (O_1451,N_49787,N_49828);
nor UO_1452 (O_1452,N_49911,N_49904);
nor UO_1453 (O_1453,N_49999,N_49775);
xor UO_1454 (O_1454,N_49765,N_49814);
and UO_1455 (O_1455,N_49821,N_49903);
nand UO_1456 (O_1456,N_49943,N_49820);
nand UO_1457 (O_1457,N_49968,N_49796);
nor UO_1458 (O_1458,N_49941,N_49834);
nand UO_1459 (O_1459,N_49763,N_49887);
or UO_1460 (O_1460,N_49864,N_49848);
nand UO_1461 (O_1461,N_49973,N_49900);
nor UO_1462 (O_1462,N_49915,N_49857);
nand UO_1463 (O_1463,N_49996,N_49916);
nand UO_1464 (O_1464,N_49792,N_49881);
and UO_1465 (O_1465,N_49982,N_49866);
nor UO_1466 (O_1466,N_49850,N_49880);
nand UO_1467 (O_1467,N_49802,N_49984);
nand UO_1468 (O_1468,N_49816,N_49763);
xnor UO_1469 (O_1469,N_49859,N_49766);
nor UO_1470 (O_1470,N_49864,N_49781);
nor UO_1471 (O_1471,N_49895,N_49828);
xor UO_1472 (O_1472,N_49860,N_49771);
nor UO_1473 (O_1473,N_49790,N_49886);
nor UO_1474 (O_1474,N_49778,N_49802);
or UO_1475 (O_1475,N_49940,N_49904);
xor UO_1476 (O_1476,N_49861,N_49784);
nand UO_1477 (O_1477,N_49801,N_49960);
nor UO_1478 (O_1478,N_49925,N_49906);
nor UO_1479 (O_1479,N_49922,N_49891);
xnor UO_1480 (O_1480,N_49804,N_49927);
nor UO_1481 (O_1481,N_49813,N_49868);
nand UO_1482 (O_1482,N_49927,N_49792);
nor UO_1483 (O_1483,N_49884,N_49750);
and UO_1484 (O_1484,N_49766,N_49887);
or UO_1485 (O_1485,N_49945,N_49755);
nor UO_1486 (O_1486,N_49845,N_49957);
nor UO_1487 (O_1487,N_49859,N_49821);
and UO_1488 (O_1488,N_49818,N_49895);
xnor UO_1489 (O_1489,N_49998,N_49875);
nand UO_1490 (O_1490,N_49870,N_49842);
nor UO_1491 (O_1491,N_49876,N_49948);
nand UO_1492 (O_1492,N_49844,N_49812);
nand UO_1493 (O_1493,N_49951,N_49913);
nand UO_1494 (O_1494,N_49896,N_49888);
nand UO_1495 (O_1495,N_49959,N_49933);
nand UO_1496 (O_1496,N_49905,N_49932);
nor UO_1497 (O_1497,N_49900,N_49888);
nor UO_1498 (O_1498,N_49868,N_49799);
nor UO_1499 (O_1499,N_49950,N_49972);
xnor UO_1500 (O_1500,N_49820,N_49791);
or UO_1501 (O_1501,N_49840,N_49996);
and UO_1502 (O_1502,N_49812,N_49837);
nand UO_1503 (O_1503,N_49915,N_49845);
nor UO_1504 (O_1504,N_49956,N_49788);
or UO_1505 (O_1505,N_49965,N_49960);
nor UO_1506 (O_1506,N_49855,N_49825);
xnor UO_1507 (O_1507,N_49943,N_49916);
nand UO_1508 (O_1508,N_49947,N_49846);
xor UO_1509 (O_1509,N_49942,N_49782);
or UO_1510 (O_1510,N_49790,N_49814);
nor UO_1511 (O_1511,N_49973,N_49980);
and UO_1512 (O_1512,N_49857,N_49839);
or UO_1513 (O_1513,N_49850,N_49817);
and UO_1514 (O_1514,N_49830,N_49768);
or UO_1515 (O_1515,N_49894,N_49859);
and UO_1516 (O_1516,N_49991,N_49842);
nor UO_1517 (O_1517,N_49892,N_49764);
nor UO_1518 (O_1518,N_49794,N_49898);
or UO_1519 (O_1519,N_49773,N_49992);
nor UO_1520 (O_1520,N_49874,N_49950);
and UO_1521 (O_1521,N_49991,N_49970);
nor UO_1522 (O_1522,N_49900,N_49974);
nor UO_1523 (O_1523,N_49814,N_49899);
nor UO_1524 (O_1524,N_49954,N_49965);
nor UO_1525 (O_1525,N_49894,N_49910);
nand UO_1526 (O_1526,N_49855,N_49980);
and UO_1527 (O_1527,N_49987,N_49806);
nor UO_1528 (O_1528,N_49801,N_49935);
xnor UO_1529 (O_1529,N_49764,N_49971);
nand UO_1530 (O_1530,N_49881,N_49758);
or UO_1531 (O_1531,N_49900,N_49910);
nor UO_1532 (O_1532,N_49807,N_49981);
xnor UO_1533 (O_1533,N_49963,N_49902);
nor UO_1534 (O_1534,N_49790,N_49973);
and UO_1535 (O_1535,N_49827,N_49776);
nand UO_1536 (O_1536,N_49925,N_49858);
and UO_1537 (O_1537,N_49962,N_49889);
or UO_1538 (O_1538,N_49960,N_49956);
xor UO_1539 (O_1539,N_49797,N_49804);
xor UO_1540 (O_1540,N_49754,N_49794);
xnor UO_1541 (O_1541,N_49920,N_49751);
xor UO_1542 (O_1542,N_49864,N_49990);
or UO_1543 (O_1543,N_49898,N_49808);
nor UO_1544 (O_1544,N_49978,N_49863);
nor UO_1545 (O_1545,N_49795,N_49980);
xnor UO_1546 (O_1546,N_49980,N_49771);
or UO_1547 (O_1547,N_49939,N_49766);
xor UO_1548 (O_1548,N_49750,N_49982);
or UO_1549 (O_1549,N_49859,N_49896);
nor UO_1550 (O_1550,N_49754,N_49835);
and UO_1551 (O_1551,N_49939,N_49768);
xnor UO_1552 (O_1552,N_49840,N_49811);
and UO_1553 (O_1553,N_49786,N_49844);
or UO_1554 (O_1554,N_49867,N_49816);
nor UO_1555 (O_1555,N_49928,N_49969);
xor UO_1556 (O_1556,N_49934,N_49756);
nor UO_1557 (O_1557,N_49933,N_49788);
nor UO_1558 (O_1558,N_49993,N_49815);
and UO_1559 (O_1559,N_49845,N_49791);
nor UO_1560 (O_1560,N_49799,N_49865);
nand UO_1561 (O_1561,N_49922,N_49917);
nor UO_1562 (O_1562,N_49966,N_49921);
or UO_1563 (O_1563,N_49862,N_49916);
xor UO_1564 (O_1564,N_49789,N_49969);
or UO_1565 (O_1565,N_49763,N_49847);
and UO_1566 (O_1566,N_49778,N_49931);
nand UO_1567 (O_1567,N_49935,N_49958);
nor UO_1568 (O_1568,N_49869,N_49863);
or UO_1569 (O_1569,N_49795,N_49821);
or UO_1570 (O_1570,N_49897,N_49807);
or UO_1571 (O_1571,N_49852,N_49926);
and UO_1572 (O_1572,N_49838,N_49925);
or UO_1573 (O_1573,N_49815,N_49770);
xor UO_1574 (O_1574,N_49847,N_49803);
nor UO_1575 (O_1575,N_49861,N_49941);
and UO_1576 (O_1576,N_49853,N_49789);
or UO_1577 (O_1577,N_49796,N_49804);
or UO_1578 (O_1578,N_49992,N_49808);
nand UO_1579 (O_1579,N_49961,N_49810);
or UO_1580 (O_1580,N_49864,N_49818);
and UO_1581 (O_1581,N_49884,N_49776);
nand UO_1582 (O_1582,N_49832,N_49979);
or UO_1583 (O_1583,N_49975,N_49763);
or UO_1584 (O_1584,N_49960,N_49792);
or UO_1585 (O_1585,N_49915,N_49788);
nand UO_1586 (O_1586,N_49923,N_49890);
and UO_1587 (O_1587,N_49917,N_49867);
and UO_1588 (O_1588,N_49939,N_49837);
or UO_1589 (O_1589,N_49791,N_49921);
and UO_1590 (O_1590,N_49886,N_49824);
and UO_1591 (O_1591,N_49979,N_49826);
nor UO_1592 (O_1592,N_49905,N_49895);
and UO_1593 (O_1593,N_49770,N_49791);
and UO_1594 (O_1594,N_49782,N_49772);
nand UO_1595 (O_1595,N_49918,N_49849);
nor UO_1596 (O_1596,N_49853,N_49824);
nor UO_1597 (O_1597,N_49935,N_49788);
xnor UO_1598 (O_1598,N_49847,N_49825);
xnor UO_1599 (O_1599,N_49975,N_49862);
xor UO_1600 (O_1600,N_49838,N_49896);
nand UO_1601 (O_1601,N_49935,N_49864);
and UO_1602 (O_1602,N_49875,N_49991);
or UO_1603 (O_1603,N_49935,N_49791);
nand UO_1604 (O_1604,N_49885,N_49952);
and UO_1605 (O_1605,N_49909,N_49963);
nor UO_1606 (O_1606,N_49860,N_49945);
xnor UO_1607 (O_1607,N_49894,N_49766);
xnor UO_1608 (O_1608,N_49927,N_49811);
xor UO_1609 (O_1609,N_49843,N_49968);
xor UO_1610 (O_1610,N_49970,N_49956);
and UO_1611 (O_1611,N_49956,N_49909);
nor UO_1612 (O_1612,N_49859,N_49916);
nand UO_1613 (O_1613,N_49914,N_49773);
nor UO_1614 (O_1614,N_49962,N_49971);
nor UO_1615 (O_1615,N_49782,N_49895);
xnor UO_1616 (O_1616,N_49758,N_49829);
xor UO_1617 (O_1617,N_49992,N_49887);
or UO_1618 (O_1618,N_49996,N_49906);
or UO_1619 (O_1619,N_49806,N_49804);
or UO_1620 (O_1620,N_49962,N_49982);
xnor UO_1621 (O_1621,N_49885,N_49991);
nand UO_1622 (O_1622,N_49997,N_49782);
nand UO_1623 (O_1623,N_49953,N_49952);
nor UO_1624 (O_1624,N_49959,N_49776);
and UO_1625 (O_1625,N_49753,N_49758);
nor UO_1626 (O_1626,N_49790,N_49872);
nand UO_1627 (O_1627,N_49979,N_49794);
xnor UO_1628 (O_1628,N_49910,N_49804);
and UO_1629 (O_1629,N_49890,N_49879);
and UO_1630 (O_1630,N_49948,N_49978);
nand UO_1631 (O_1631,N_49954,N_49941);
and UO_1632 (O_1632,N_49943,N_49928);
xor UO_1633 (O_1633,N_49805,N_49860);
and UO_1634 (O_1634,N_49894,N_49962);
or UO_1635 (O_1635,N_49856,N_49783);
xor UO_1636 (O_1636,N_49816,N_49807);
and UO_1637 (O_1637,N_49908,N_49824);
xor UO_1638 (O_1638,N_49816,N_49838);
and UO_1639 (O_1639,N_49905,N_49997);
nor UO_1640 (O_1640,N_49908,N_49972);
or UO_1641 (O_1641,N_49848,N_49912);
nor UO_1642 (O_1642,N_49890,N_49824);
nand UO_1643 (O_1643,N_49793,N_49841);
xor UO_1644 (O_1644,N_49752,N_49787);
or UO_1645 (O_1645,N_49953,N_49878);
or UO_1646 (O_1646,N_49924,N_49817);
or UO_1647 (O_1647,N_49860,N_49942);
or UO_1648 (O_1648,N_49915,N_49981);
or UO_1649 (O_1649,N_49974,N_49936);
nand UO_1650 (O_1650,N_49967,N_49995);
nor UO_1651 (O_1651,N_49964,N_49924);
nand UO_1652 (O_1652,N_49779,N_49835);
nor UO_1653 (O_1653,N_49944,N_49771);
nor UO_1654 (O_1654,N_49853,N_49766);
nand UO_1655 (O_1655,N_49803,N_49811);
nand UO_1656 (O_1656,N_49951,N_49752);
nand UO_1657 (O_1657,N_49927,N_49784);
or UO_1658 (O_1658,N_49947,N_49898);
nand UO_1659 (O_1659,N_49760,N_49810);
nand UO_1660 (O_1660,N_49860,N_49964);
xor UO_1661 (O_1661,N_49981,N_49995);
xnor UO_1662 (O_1662,N_49841,N_49837);
or UO_1663 (O_1663,N_49933,N_49920);
nor UO_1664 (O_1664,N_49947,N_49851);
nand UO_1665 (O_1665,N_49846,N_49784);
nand UO_1666 (O_1666,N_49948,N_49859);
xor UO_1667 (O_1667,N_49826,N_49753);
xor UO_1668 (O_1668,N_49876,N_49764);
nor UO_1669 (O_1669,N_49889,N_49892);
and UO_1670 (O_1670,N_49789,N_49765);
and UO_1671 (O_1671,N_49995,N_49776);
or UO_1672 (O_1672,N_49935,N_49953);
nor UO_1673 (O_1673,N_49935,N_49898);
and UO_1674 (O_1674,N_49863,N_49910);
nand UO_1675 (O_1675,N_49982,N_49865);
and UO_1676 (O_1676,N_49759,N_49881);
or UO_1677 (O_1677,N_49929,N_49882);
and UO_1678 (O_1678,N_49775,N_49896);
and UO_1679 (O_1679,N_49863,N_49826);
xnor UO_1680 (O_1680,N_49938,N_49763);
xnor UO_1681 (O_1681,N_49932,N_49968);
nand UO_1682 (O_1682,N_49991,N_49752);
xor UO_1683 (O_1683,N_49965,N_49883);
or UO_1684 (O_1684,N_49900,N_49928);
nor UO_1685 (O_1685,N_49843,N_49823);
nand UO_1686 (O_1686,N_49922,N_49835);
nor UO_1687 (O_1687,N_49875,N_49948);
or UO_1688 (O_1688,N_49844,N_49780);
or UO_1689 (O_1689,N_49781,N_49943);
nor UO_1690 (O_1690,N_49885,N_49931);
nand UO_1691 (O_1691,N_49957,N_49873);
nor UO_1692 (O_1692,N_49759,N_49791);
xor UO_1693 (O_1693,N_49906,N_49975);
nand UO_1694 (O_1694,N_49899,N_49815);
nor UO_1695 (O_1695,N_49780,N_49947);
nor UO_1696 (O_1696,N_49773,N_49828);
and UO_1697 (O_1697,N_49805,N_49862);
nand UO_1698 (O_1698,N_49751,N_49755);
and UO_1699 (O_1699,N_49928,N_49945);
nand UO_1700 (O_1700,N_49926,N_49820);
and UO_1701 (O_1701,N_49760,N_49804);
nor UO_1702 (O_1702,N_49854,N_49966);
and UO_1703 (O_1703,N_49783,N_49800);
or UO_1704 (O_1704,N_49922,N_49754);
and UO_1705 (O_1705,N_49799,N_49968);
nand UO_1706 (O_1706,N_49983,N_49962);
or UO_1707 (O_1707,N_49962,N_49869);
or UO_1708 (O_1708,N_49826,N_49774);
xnor UO_1709 (O_1709,N_49808,N_49895);
and UO_1710 (O_1710,N_49976,N_49963);
xnor UO_1711 (O_1711,N_49786,N_49769);
xnor UO_1712 (O_1712,N_49970,N_49927);
nor UO_1713 (O_1713,N_49826,N_49981);
xnor UO_1714 (O_1714,N_49796,N_49954);
nand UO_1715 (O_1715,N_49838,N_49924);
or UO_1716 (O_1716,N_49772,N_49932);
nor UO_1717 (O_1717,N_49811,N_49806);
or UO_1718 (O_1718,N_49996,N_49860);
and UO_1719 (O_1719,N_49936,N_49903);
nand UO_1720 (O_1720,N_49889,N_49904);
and UO_1721 (O_1721,N_49898,N_49845);
nor UO_1722 (O_1722,N_49952,N_49788);
nand UO_1723 (O_1723,N_49905,N_49941);
nor UO_1724 (O_1724,N_49983,N_49978);
nor UO_1725 (O_1725,N_49835,N_49771);
xor UO_1726 (O_1726,N_49902,N_49833);
or UO_1727 (O_1727,N_49934,N_49998);
or UO_1728 (O_1728,N_49958,N_49811);
xnor UO_1729 (O_1729,N_49900,N_49782);
xor UO_1730 (O_1730,N_49753,N_49969);
xor UO_1731 (O_1731,N_49845,N_49822);
xnor UO_1732 (O_1732,N_49969,N_49951);
nand UO_1733 (O_1733,N_49762,N_49917);
xor UO_1734 (O_1734,N_49895,N_49920);
or UO_1735 (O_1735,N_49894,N_49929);
nor UO_1736 (O_1736,N_49822,N_49853);
or UO_1737 (O_1737,N_49853,N_49885);
and UO_1738 (O_1738,N_49997,N_49778);
or UO_1739 (O_1739,N_49984,N_49973);
or UO_1740 (O_1740,N_49872,N_49849);
xnor UO_1741 (O_1741,N_49844,N_49980);
xnor UO_1742 (O_1742,N_49776,N_49815);
xnor UO_1743 (O_1743,N_49998,N_49891);
nand UO_1744 (O_1744,N_49806,N_49910);
nor UO_1745 (O_1745,N_49791,N_49779);
nand UO_1746 (O_1746,N_49915,N_49910);
or UO_1747 (O_1747,N_49986,N_49973);
nor UO_1748 (O_1748,N_49822,N_49952);
and UO_1749 (O_1749,N_49894,N_49991);
or UO_1750 (O_1750,N_49939,N_49916);
or UO_1751 (O_1751,N_49930,N_49822);
nand UO_1752 (O_1752,N_49936,N_49891);
or UO_1753 (O_1753,N_49809,N_49999);
or UO_1754 (O_1754,N_49927,N_49755);
xor UO_1755 (O_1755,N_49906,N_49911);
xor UO_1756 (O_1756,N_49888,N_49955);
nand UO_1757 (O_1757,N_49916,N_49838);
xnor UO_1758 (O_1758,N_49835,N_49789);
nand UO_1759 (O_1759,N_49833,N_49786);
or UO_1760 (O_1760,N_49878,N_49835);
and UO_1761 (O_1761,N_49800,N_49882);
nand UO_1762 (O_1762,N_49867,N_49755);
xor UO_1763 (O_1763,N_49973,N_49997);
nand UO_1764 (O_1764,N_49963,N_49899);
nor UO_1765 (O_1765,N_49864,N_49913);
xnor UO_1766 (O_1766,N_49927,N_49759);
nand UO_1767 (O_1767,N_49915,N_49773);
and UO_1768 (O_1768,N_49768,N_49840);
nand UO_1769 (O_1769,N_49764,N_49901);
and UO_1770 (O_1770,N_49946,N_49952);
nor UO_1771 (O_1771,N_49931,N_49832);
xnor UO_1772 (O_1772,N_49835,N_49970);
nand UO_1773 (O_1773,N_49981,N_49758);
nor UO_1774 (O_1774,N_49869,N_49950);
and UO_1775 (O_1775,N_49956,N_49812);
and UO_1776 (O_1776,N_49758,N_49856);
and UO_1777 (O_1777,N_49783,N_49950);
and UO_1778 (O_1778,N_49957,N_49865);
nor UO_1779 (O_1779,N_49888,N_49972);
or UO_1780 (O_1780,N_49905,N_49823);
or UO_1781 (O_1781,N_49877,N_49990);
nand UO_1782 (O_1782,N_49919,N_49908);
nor UO_1783 (O_1783,N_49774,N_49955);
or UO_1784 (O_1784,N_49869,N_49803);
nand UO_1785 (O_1785,N_49945,N_49816);
xnor UO_1786 (O_1786,N_49849,N_49887);
or UO_1787 (O_1787,N_49902,N_49882);
or UO_1788 (O_1788,N_49956,N_49895);
nor UO_1789 (O_1789,N_49840,N_49770);
and UO_1790 (O_1790,N_49783,N_49873);
nand UO_1791 (O_1791,N_49791,N_49992);
nand UO_1792 (O_1792,N_49860,N_49830);
nand UO_1793 (O_1793,N_49846,N_49818);
or UO_1794 (O_1794,N_49873,N_49996);
nand UO_1795 (O_1795,N_49923,N_49946);
xnor UO_1796 (O_1796,N_49755,N_49803);
xnor UO_1797 (O_1797,N_49872,N_49753);
nor UO_1798 (O_1798,N_49976,N_49999);
and UO_1799 (O_1799,N_49927,N_49937);
or UO_1800 (O_1800,N_49759,N_49895);
and UO_1801 (O_1801,N_49856,N_49892);
xnor UO_1802 (O_1802,N_49771,N_49849);
nor UO_1803 (O_1803,N_49902,N_49784);
nand UO_1804 (O_1804,N_49935,N_49907);
nand UO_1805 (O_1805,N_49967,N_49887);
nor UO_1806 (O_1806,N_49793,N_49952);
and UO_1807 (O_1807,N_49952,N_49972);
or UO_1808 (O_1808,N_49988,N_49856);
nand UO_1809 (O_1809,N_49852,N_49855);
xnor UO_1810 (O_1810,N_49901,N_49964);
or UO_1811 (O_1811,N_49750,N_49803);
or UO_1812 (O_1812,N_49824,N_49781);
or UO_1813 (O_1813,N_49828,N_49808);
xor UO_1814 (O_1814,N_49820,N_49803);
nor UO_1815 (O_1815,N_49915,N_49917);
and UO_1816 (O_1816,N_49997,N_49823);
xnor UO_1817 (O_1817,N_49986,N_49883);
nand UO_1818 (O_1818,N_49804,N_49773);
and UO_1819 (O_1819,N_49775,N_49968);
nor UO_1820 (O_1820,N_49901,N_49768);
or UO_1821 (O_1821,N_49764,N_49993);
nand UO_1822 (O_1822,N_49835,N_49932);
xnor UO_1823 (O_1823,N_49983,N_49779);
nor UO_1824 (O_1824,N_49816,N_49903);
nand UO_1825 (O_1825,N_49852,N_49817);
xnor UO_1826 (O_1826,N_49817,N_49860);
nand UO_1827 (O_1827,N_49762,N_49851);
and UO_1828 (O_1828,N_49834,N_49750);
nand UO_1829 (O_1829,N_49798,N_49935);
nor UO_1830 (O_1830,N_49791,N_49962);
xor UO_1831 (O_1831,N_49892,N_49893);
nand UO_1832 (O_1832,N_49796,N_49818);
or UO_1833 (O_1833,N_49917,N_49852);
nor UO_1834 (O_1834,N_49943,N_49980);
and UO_1835 (O_1835,N_49808,N_49913);
or UO_1836 (O_1836,N_49806,N_49947);
nand UO_1837 (O_1837,N_49847,N_49842);
and UO_1838 (O_1838,N_49887,N_49914);
and UO_1839 (O_1839,N_49936,N_49811);
nor UO_1840 (O_1840,N_49892,N_49933);
nor UO_1841 (O_1841,N_49839,N_49833);
nand UO_1842 (O_1842,N_49969,N_49827);
or UO_1843 (O_1843,N_49763,N_49756);
nand UO_1844 (O_1844,N_49789,N_49901);
nand UO_1845 (O_1845,N_49805,N_49983);
and UO_1846 (O_1846,N_49782,N_49850);
or UO_1847 (O_1847,N_49757,N_49810);
nor UO_1848 (O_1848,N_49926,N_49879);
nand UO_1849 (O_1849,N_49838,N_49809);
nor UO_1850 (O_1850,N_49782,N_49937);
and UO_1851 (O_1851,N_49857,N_49900);
or UO_1852 (O_1852,N_49977,N_49829);
xor UO_1853 (O_1853,N_49790,N_49898);
and UO_1854 (O_1854,N_49953,N_49768);
nor UO_1855 (O_1855,N_49891,N_49959);
xor UO_1856 (O_1856,N_49800,N_49975);
nor UO_1857 (O_1857,N_49818,N_49936);
nor UO_1858 (O_1858,N_49979,N_49955);
and UO_1859 (O_1859,N_49944,N_49963);
and UO_1860 (O_1860,N_49892,N_49914);
nor UO_1861 (O_1861,N_49787,N_49921);
and UO_1862 (O_1862,N_49794,N_49763);
and UO_1863 (O_1863,N_49782,N_49760);
nand UO_1864 (O_1864,N_49951,N_49841);
nor UO_1865 (O_1865,N_49984,N_49874);
and UO_1866 (O_1866,N_49846,N_49844);
and UO_1867 (O_1867,N_49777,N_49750);
nand UO_1868 (O_1868,N_49782,N_49947);
xor UO_1869 (O_1869,N_49927,N_49795);
nor UO_1870 (O_1870,N_49836,N_49823);
and UO_1871 (O_1871,N_49840,N_49809);
or UO_1872 (O_1872,N_49762,N_49870);
and UO_1873 (O_1873,N_49823,N_49918);
or UO_1874 (O_1874,N_49879,N_49838);
nand UO_1875 (O_1875,N_49824,N_49857);
and UO_1876 (O_1876,N_49775,N_49774);
and UO_1877 (O_1877,N_49983,N_49884);
and UO_1878 (O_1878,N_49821,N_49930);
and UO_1879 (O_1879,N_49908,N_49811);
nand UO_1880 (O_1880,N_49977,N_49963);
nand UO_1881 (O_1881,N_49983,N_49792);
and UO_1882 (O_1882,N_49887,N_49909);
or UO_1883 (O_1883,N_49826,N_49998);
xor UO_1884 (O_1884,N_49897,N_49865);
xor UO_1885 (O_1885,N_49926,N_49982);
and UO_1886 (O_1886,N_49777,N_49835);
or UO_1887 (O_1887,N_49986,N_49887);
or UO_1888 (O_1888,N_49827,N_49916);
nor UO_1889 (O_1889,N_49986,N_49939);
xnor UO_1890 (O_1890,N_49964,N_49872);
and UO_1891 (O_1891,N_49881,N_49763);
xnor UO_1892 (O_1892,N_49880,N_49778);
or UO_1893 (O_1893,N_49830,N_49796);
nor UO_1894 (O_1894,N_49820,N_49908);
or UO_1895 (O_1895,N_49903,N_49886);
nand UO_1896 (O_1896,N_49891,N_49992);
nor UO_1897 (O_1897,N_49775,N_49951);
and UO_1898 (O_1898,N_49878,N_49968);
and UO_1899 (O_1899,N_49825,N_49805);
and UO_1900 (O_1900,N_49898,N_49918);
xnor UO_1901 (O_1901,N_49932,N_49769);
and UO_1902 (O_1902,N_49901,N_49816);
nor UO_1903 (O_1903,N_49894,N_49934);
nand UO_1904 (O_1904,N_49926,N_49974);
and UO_1905 (O_1905,N_49900,N_49862);
xor UO_1906 (O_1906,N_49764,N_49897);
or UO_1907 (O_1907,N_49859,N_49981);
or UO_1908 (O_1908,N_49823,N_49900);
and UO_1909 (O_1909,N_49941,N_49774);
nand UO_1910 (O_1910,N_49978,N_49819);
nor UO_1911 (O_1911,N_49921,N_49875);
xor UO_1912 (O_1912,N_49929,N_49890);
nand UO_1913 (O_1913,N_49937,N_49896);
nor UO_1914 (O_1914,N_49866,N_49964);
and UO_1915 (O_1915,N_49868,N_49977);
and UO_1916 (O_1916,N_49940,N_49793);
xor UO_1917 (O_1917,N_49772,N_49765);
and UO_1918 (O_1918,N_49826,N_49983);
nor UO_1919 (O_1919,N_49962,N_49872);
xor UO_1920 (O_1920,N_49928,N_49912);
or UO_1921 (O_1921,N_49870,N_49751);
or UO_1922 (O_1922,N_49796,N_49981);
and UO_1923 (O_1923,N_49879,N_49889);
nand UO_1924 (O_1924,N_49982,N_49892);
nor UO_1925 (O_1925,N_49808,N_49977);
and UO_1926 (O_1926,N_49902,N_49879);
nor UO_1927 (O_1927,N_49876,N_49899);
nand UO_1928 (O_1928,N_49852,N_49765);
xnor UO_1929 (O_1929,N_49958,N_49891);
and UO_1930 (O_1930,N_49897,N_49939);
nor UO_1931 (O_1931,N_49763,N_49845);
xnor UO_1932 (O_1932,N_49903,N_49771);
nand UO_1933 (O_1933,N_49836,N_49919);
xnor UO_1934 (O_1934,N_49824,N_49861);
xnor UO_1935 (O_1935,N_49938,N_49994);
xor UO_1936 (O_1936,N_49843,N_49864);
xnor UO_1937 (O_1937,N_49863,N_49908);
and UO_1938 (O_1938,N_49913,N_49843);
xor UO_1939 (O_1939,N_49975,N_49965);
and UO_1940 (O_1940,N_49910,N_49884);
nor UO_1941 (O_1941,N_49880,N_49845);
and UO_1942 (O_1942,N_49954,N_49787);
and UO_1943 (O_1943,N_49973,N_49779);
and UO_1944 (O_1944,N_49913,N_49769);
nand UO_1945 (O_1945,N_49897,N_49876);
or UO_1946 (O_1946,N_49910,N_49800);
xor UO_1947 (O_1947,N_49970,N_49863);
xnor UO_1948 (O_1948,N_49852,N_49913);
nor UO_1949 (O_1949,N_49780,N_49949);
nor UO_1950 (O_1950,N_49756,N_49864);
nand UO_1951 (O_1951,N_49828,N_49771);
nor UO_1952 (O_1952,N_49774,N_49977);
and UO_1953 (O_1953,N_49950,N_49900);
nand UO_1954 (O_1954,N_49794,N_49786);
xnor UO_1955 (O_1955,N_49780,N_49959);
xnor UO_1956 (O_1956,N_49979,N_49755);
nand UO_1957 (O_1957,N_49883,N_49774);
or UO_1958 (O_1958,N_49878,N_49948);
nand UO_1959 (O_1959,N_49898,N_49996);
or UO_1960 (O_1960,N_49788,N_49883);
xor UO_1961 (O_1961,N_49780,N_49777);
xnor UO_1962 (O_1962,N_49758,N_49840);
xnor UO_1963 (O_1963,N_49913,N_49872);
xnor UO_1964 (O_1964,N_49861,N_49787);
xnor UO_1965 (O_1965,N_49961,N_49957);
and UO_1966 (O_1966,N_49970,N_49900);
nor UO_1967 (O_1967,N_49776,N_49817);
nand UO_1968 (O_1968,N_49998,N_49882);
xor UO_1969 (O_1969,N_49814,N_49826);
and UO_1970 (O_1970,N_49946,N_49931);
xor UO_1971 (O_1971,N_49900,N_49772);
xor UO_1972 (O_1972,N_49780,N_49874);
xnor UO_1973 (O_1973,N_49996,N_49901);
and UO_1974 (O_1974,N_49946,N_49971);
nor UO_1975 (O_1975,N_49800,N_49806);
nor UO_1976 (O_1976,N_49767,N_49864);
nand UO_1977 (O_1977,N_49920,N_49995);
nand UO_1978 (O_1978,N_49836,N_49852);
and UO_1979 (O_1979,N_49803,N_49833);
and UO_1980 (O_1980,N_49926,N_49954);
or UO_1981 (O_1981,N_49915,N_49801);
and UO_1982 (O_1982,N_49825,N_49899);
xor UO_1983 (O_1983,N_49768,N_49876);
and UO_1984 (O_1984,N_49865,N_49889);
nand UO_1985 (O_1985,N_49772,N_49825);
or UO_1986 (O_1986,N_49971,N_49790);
xor UO_1987 (O_1987,N_49767,N_49921);
xor UO_1988 (O_1988,N_49780,N_49962);
and UO_1989 (O_1989,N_49754,N_49792);
or UO_1990 (O_1990,N_49987,N_49781);
nand UO_1991 (O_1991,N_49770,N_49884);
nand UO_1992 (O_1992,N_49832,N_49856);
nor UO_1993 (O_1993,N_49985,N_49904);
xnor UO_1994 (O_1994,N_49913,N_49801);
xor UO_1995 (O_1995,N_49928,N_49786);
nand UO_1996 (O_1996,N_49984,N_49965);
nand UO_1997 (O_1997,N_49990,N_49966);
nand UO_1998 (O_1998,N_49863,N_49954);
xor UO_1999 (O_1999,N_49792,N_49928);
or UO_2000 (O_2000,N_49933,N_49927);
nand UO_2001 (O_2001,N_49950,N_49983);
or UO_2002 (O_2002,N_49790,N_49831);
nor UO_2003 (O_2003,N_49808,N_49815);
nor UO_2004 (O_2004,N_49871,N_49974);
or UO_2005 (O_2005,N_49872,N_49765);
or UO_2006 (O_2006,N_49765,N_49812);
xor UO_2007 (O_2007,N_49769,N_49879);
xnor UO_2008 (O_2008,N_49821,N_49804);
or UO_2009 (O_2009,N_49938,N_49868);
nor UO_2010 (O_2010,N_49939,N_49978);
nor UO_2011 (O_2011,N_49979,N_49769);
nand UO_2012 (O_2012,N_49871,N_49891);
nand UO_2013 (O_2013,N_49926,N_49966);
xnor UO_2014 (O_2014,N_49957,N_49954);
or UO_2015 (O_2015,N_49957,N_49774);
and UO_2016 (O_2016,N_49888,N_49954);
nand UO_2017 (O_2017,N_49796,N_49811);
nor UO_2018 (O_2018,N_49836,N_49929);
nand UO_2019 (O_2019,N_49995,N_49775);
xnor UO_2020 (O_2020,N_49951,N_49928);
nand UO_2021 (O_2021,N_49988,N_49919);
nand UO_2022 (O_2022,N_49952,N_49950);
and UO_2023 (O_2023,N_49837,N_49917);
nand UO_2024 (O_2024,N_49760,N_49958);
xor UO_2025 (O_2025,N_49777,N_49952);
xnor UO_2026 (O_2026,N_49954,N_49774);
and UO_2027 (O_2027,N_49919,N_49954);
nor UO_2028 (O_2028,N_49844,N_49952);
nor UO_2029 (O_2029,N_49828,N_49986);
and UO_2030 (O_2030,N_49924,N_49914);
and UO_2031 (O_2031,N_49764,N_49859);
nand UO_2032 (O_2032,N_49970,N_49847);
xnor UO_2033 (O_2033,N_49775,N_49877);
or UO_2034 (O_2034,N_49939,N_49801);
or UO_2035 (O_2035,N_49751,N_49914);
nor UO_2036 (O_2036,N_49837,N_49895);
and UO_2037 (O_2037,N_49904,N_49924);
and UO_2038 (O_2038,N_49777,N_49959);
xor UO_2039 (O_2039,N_49962,N_49916);
nand UO_2040 (O_2040,N_49919,N_49850);
xnor UO_2041 (O_2041,N_49934,N_49865);
nor UO_2042 (O_2042,N_49912,N_49877);
and UO_2043 (O_2043,N_49898,N_49782);
and UO_2044 (O_2044,N_49863,N_49849);
or UO_2045 (O_2045,N_49939,N_49951);
and UO_2046 (O_2046,N_49879,N_49917);
nand UO_2047 (O_2047,N_49895,N_49779);
nor UO_2048 (O_2048,N_49779,N_49967);
nand UO_2049 (O_2049,N_49903,N_49908);
nor UO_2050 (O_2050,N_49929,N_49762);
nand UO_2051 (O_2051,N_49890,N_49975);
xnor UO_2052 (O_2052,N_49813,N_49992);
nand UO_2053 (O_2053,N_49850,N_49822);
nand UO_2054 (O_2054,N_49824,N_49804);
or UO_2055 (O_2055,N_49768,N_49793);
nand UO_2056 (O_2056,N_49920,N_49922);
or UO_2057 (O_2057,N_49897,N_49921);
nor UO_2058 (O_2058,N_49786,N_49868);
nand UO_2059 (O_2059,N_49885,N_49958);
nor UO_2060 (O_2060,N_49842,N_49934);
or UO_2061 (O_2061,N_49942,N_49853);
nand UO_2062 (O_2062,N_49847,N_49888);
and UO_2063 (O_2063,N_49854,N_49824);
and UO_2064 (O_2064,N_49936,N_49776);
nand UO_2065 (O_2065,N_49847,N_49846);
xnor UO_2066 (O_2066,N_49853,N_49762);
and UO_2067 (O_2067,N_49790,N_49838);
nand UO_2068 (O_2068,N_49993,N_49968);
or UO_2069 (O_2069,N_49818,N_49916);
or UO_2070 (O_2070,N_49944,N_49928);
or UO_2071 (O_2071,N_49807,N_49780);
nand UO_2072 (O_2072,N_49879,N_49886);
xor UO_2073 (O_2073,N_49984,N_49854);
nand UO_2074 (O_2074,N_49982,N_49874);
or UO_2075 (O_2075,N_49909,N_49946);
or UO_2076 (O_2076,N_49819,N_49787);
or UO_2077 (O_2077,N_49819,N_49772);
nand UO_2078 (O_2078,N_49978,N_49791);
xnor UO_2079 (O_2079,N_49766,N_49799);
and UO_2080 (O_2080,N_49760,N_49780);
xor UO_2081 (O_2081,N_49811,N_49750);
nor UO_2082 (O_2082,N_49969,N_49901);
or UO_2083 (O_2083,N_49917,N_49854);
nand UO_2084 (O_2084,N_49967,N_49826);
nand UO_2085 (O_2085,N_49980,N_49838);
or UO_2086 (O_2086,N_49813,N_49804);
nor UO_2087 (O_2087,N_49927,N_49876);
and UO_2088 (O_2088,N_49757,N_49956);
nand UO_2089 (O_2089,N_49881,N_49773);
nand UO_2090 (O_2090,N_49893,N_49768);
nand UO_2091 (O_2091,N_49832,N_49915);
and UO_2092 (O_2092,N_49892,N_49937);
nand UO_2093 (O_2093,N_49959,N_49845);
or UO_2094 (O_2094,N_49773,N_49904);
nand UO_2095 (O_2095,N_49874,N_49882);
nand UO_2096 (O_2096,N_49882,N_49921);
nor UO_2097 (O_2097,N_49951,N_49874);
nor UO_2098 (O_2098,N_49976,N_49962);
nor UO_2099 (O_2099,N_49988,N_49976);
or UO_2100 (O_2100,N_49966,N_49804);
nor UO_2101 (O_2101,N_49844,N_49759);
or UO_2102 (O_2102,N_49903,N_49847);
or UO_2103 (O_2103,N_49955,N_49751);
nor UO_2104 (O_2104,N_49911,N_49988);
nor UO_2105 (O_2105,N_49884,N_49796);
or UO_2106 (O_2106,N_49885,N_49904);
xor UO_2107 (O_2107,N_49916,N_49864);
nor UO_2108 (O_2108,N_49916,N_49840);
nand UO_2109 (O_2109,N_49876,N_49952);
nand UO_2110 (O_2110,N_49952,N_49865);
nor UO_2111 (O_2111,N_49837,N_49760);
nor UO_2112 (O_2112,N_49860,N_49840);
nand UO_2113 (O_2113,N_49754,N_49914);
nor UO_2114 (O_2114,N_49987,N_49750);
or UO_2115 (O_2115,N_49952,N_49961);
and UO_2116 (O_2116,N_49768,N_49878);
nor UO_2117 (O_2117,N_49829,N_49855);
and UO_2118 (O_2118,N_49876,N_49988);
and UO_2119 (O_2119,N_49895,N_49962);
xor UO_2120 (O_2120,N_49988,N_49975);
and UO_2121 (O_2121,N_49979,N_49956);
nand UO_2122 (O_2122,N_49770,N_49847);
or UO_2123 (O_2123,N_49794,N_49932);
or UO_2124 (O_2124,N_49919,N_49950);
and UO_2125 (O_2125,N_49985,N_49770);
and UO_2126 (O_2126,N_49915,N_49907);
xor UO_2127 (O_2127,N_49774,N_49926);
xor UO_2128 (O_2128,N_49770,N_49948);
nand UO_2129 (O_2129,N_49940,N_49755);
xnor UO_2130 (O_2130,N_49943,N_49777);
nor UO_2131 (O_2131,N_49789,N_49932);
nor UO_2132 (O_2132,N_49847,N_49943);
nor UO_2133 (O_2133,N_49952,N_49963);
or UO_2134 (O_2134,N_49785,N_49883);
or UO_2135 (O_2135,N_49827,N_49845);
or UO_2136 (O_2136,N_49804,N_49911);
nor UO_2137 (O_2137,N_49853,N_49851);
or UO_2138 (O_2138,N_49843,N_49989);
and UO_2139 (O_2139,N_49768,N_49949);
and UO_2140 (O_2140,N_49801,N_49882);
and UO_2141 (O_2141,N_49857,N_49941);
or UO_2142 (O_2142,N_49826,N_49961);
xnor UO_2143 (O_2143,N_49953,N_49840);
or UO_2144 (O_2144,N_49985,N_49761);
xor UO_2145 (O_2145,N_49922,N_49907);
or UO_2146 (O_2146,N_49830,N_49991);
and UO_2147 (O_2147,N_49786,N_49834);
or UO_2148 (O_2148,N_49966,N_49982);
and UO_2149 (O_2149,N_49899,N_49756);
nor UO_2150 (O_2150,N_49897,N_49829);
and UO_2151 (O_2151,N_49945,N_49904);
nor UO_2152 (O_2152,N_49977,N_49882);
nand UO_2153 (O_2153,N_49931,N_49856);
nor UO_2154 (O_2154,N_49829,N_49785);
nand UO_2155 (O_2155,N_49801,N_49948);
or UO_2156 (O_2156,N_49804,N_49836);
and UO_2157 (O_2157,N_49864,N_49888);
or UO_2158 (O_2158,N_49928,N_49756);
nand UO_2159 (O_2159,N_49772,N_49962);
xnor UO_2160 (O_2160,N_49976,N_49876);
nand UO_2161 (O_2161,N_49757,N_49922);
nor UO_2162 (O_2162,N_49937,N_49978);
or UO_2163 (O_2163,N_49985,N_49983);
and UO_2164 (O_2164,N_49767,N_49980);
or UO_2165 (O_2165,N_49983,N_49922);
nor UO_2166 (O_2166,N_49751,N_49994);
and UO_2167 (O_2167,N_49887,N_49953);
or UO_2168 (O_2168,N_49927,N_49764);
or UO_2169 (O_2169,N_49988,N_49915);
or UO_2170 (O_2170,N_49995,N_49945);
or UO_2171 (O_2171,N_49831,N_49970);
nor UO_2172 (O_2172,N_49778,N_49862);
xnor UO_2173 (O_2173,N_49956,N_49915);
nand UO_2174 (O_2174,N_49832,N_49841);
or UO_2175 (O_2175,N_49823,N_49915);
nand UO_2176 (O_2176,N_49758,N_49970);
nor UO_2177 (O_2177,N_49953,N_49862);
xor UO_2178 (O_2178,N_49875,N_49770);
or UO_2179 (O_2179,N_49774,N_49823);
nand UO_2180 (O_2180,N_49810,N_49978);
xor UO_2181 (O_2181,N_49876,N_49824);
xor UO_2182 (O_2182,N_49792,N_49953);
nor UO_2183 (O_2183,N_49831,N_49933);
or UO_2184 (O_2184,N_49971,N_49900);
or UO_2185 (O_2185,N_49889,N_49923);
or UO_2186 (O_2186,N_49879,N_49796);
and UO_2187 (O_2187,N_49775,N_49918);
nand UO_2188 (O_2188,N_49825,N_49755);
xor UO_2189 (O_2189,N_49773,N_49982);
nor UO_2190 (O_2190,N_49785,N_49823);
and UO_2191 (O_2191,N_49982,N_49799);
and UO_2192 (O_2192,N_49869,N_49999);
or UO_2193 (O_2193,N_49889,N_49845);
and UO_2194 (O_2194,N_49915,N_49815);
xor UO_2195 (O_2195,N_49902,N_49766);
nor UO_2196 (O_2196,N_49911,N_49796);
nand UO_2197 (O_2197,N_49767,N_49917);
and UO_2198 (O_2198,N_49877,N_49779);
and UO_2199 (O_2199,N_49909,N_49922);
nor UO_2200 (O_2200,N_49884,N_49900);
or UO_2201 (O_2201,N_49964,N_49931);
nor UO_2202 (O_2202,N_49751,N_49776);
or UO_2203 (O_2203,N_49999,N_49988);
or UO_2204 (O_2204,N_49955,N_49967);
and UO_2205 (O_2205,N_49907,N_49990);
nand UO_2206 (O_2206,N_49939,N_49943);
nor UO_2207 (O_2207,N_49896,N_49786);
nand UO_2208 (O_2208,N_49821,N_49826);
nand UO_2209 (O_2209,N_49875,N_49920);
nand UO_2210 (O_2210,N_49859,N_49994);
nand UO_2211 (O_2211,N_49925,N_49914);
nor UO_2212 (O_2212,N_49758,N_49774);
nand UO_2213 (O_2213,N_49952,N_49767);
or UO_2214 (O_2214,N_49988,N_49898);
or UO_2215 (O_2215,N_49790,N_49913);
or UO_2216 (O_2216,N_49852,N_49970);
or UO_2217 (O_2217,N_49819,N_49929);
or UO_2218 (O_2218,N_49856,N_49876);
nor UO_2219 (O_2219,N_49793,N_49773);
nand UO_2220 (O_2220,N_49990,N_49999);
nand UO_2221 (O_2221,N_49814,N_49979);
nand UO_2222 (O_2222,N_49945,N_49898);
nor UO_2223 (O_2223,N_49955,N_49882);
and UO_2224 (O_2224,N_49781,N_49953);
xnor UO_2225 (O_2225,N_49895,N_49969);
xor UO_2226 (O_2226,N_49867,N_49910);
nor UO_2227 (O_2227,N_49996,N_49968);
and UO_2228 (O_2228,N_49874,N_49811);
or UO_2229 (O_2229,N_49897,N_49888);
xor UO_2230 (O_2230,N_49812,N_49770);
or UO_2231 (O_2231,N_49845,N_49920);
nor UO_2232 (O_2232,N_49842,N_49763);
or UO_2233 (O_2233,N_49915,N_49820);
nand UO_2234 (O_2234,N_49932,N_49767);
xnor UO_2235 (O_2235,N_49851,N_49781);
nor UO_2236 (O_2236,N_49796,N_49908);
xor UO_2237 (O_2237,N_49965,N_49763);
and UO_2238 (O_2238,N_49915,N_49786);
or UO_2239 (O_2239,N_49880,N_49978);
nand UO_2240 (O_2240,N_49924,N_49806);
nor UO_2241 (O_2241,N_49879,N_49975);
or UO_2242 (O_2242,N_49967,N_49982);
nand UO_2243 (O_2243,N_49924,N_49865);
and UO_2244 (O_2244,N_49997,N_49806);
xnor UO_2245 (O_2245,N_49831,N_49865);
nand UO_2246 (O_2246,N_49811,N_49859);
and UO_2247 (O_2247,N_49766,N_49990);
nor UO_2248 (O_2248,N_49850,N_49897);
and UO_2249 (O_2249,N_49931,N_49755);
nand UO_2250 (O_2250,N_49823,N_49767);
xor UO_2251 (O_2251,N_49921,N_49947);
nand UO_2252 (O_2252,N_49859,N_49809);
xor UO_2253 (O_2253,N_49912,N_49834);
or UO_2254 (O_2254,N_49836,N_49894);
and UO_2255 (O_2255,N_49931,N_49847);
and UO_2256 (O_2256,N_49826,N_49752);
xnor UO_2257 (O_2257,N_49974,N_49951);
and UO_2258 (O_2258,N_49871,N_49821);
nand UO_2259 (O_2259,N_49960,N_49945);
xor UO_2260 (O_2260,N_49770,N_49915);
xnor UO_2261 (O_2261,N_49943,N_49859);
or UO_2262 (O_2262,N_49877,N_49928);
xor UO_2263 (O_2263,N_49892,N_49991);
nor UO_2264 (O_2264,N_49986,N_49761);
nand UO_2265 (O_2265,N_49829,N_49789);
or UO_2266 (O_2266,N_49930,N_49790);
nand UO_2267 (O_2267,N_49978,N_49766);
nand UO_2268 (O_2268,N_49783,N_49912);
xor UO_2269 (O_2269,N_49969,N_49980);
or UO_2270 (O_2270,N_49822,N_49767);
nand UO_2271 (O_2271,N_49873,N_49779);
nor UO_2272 (O_2272,N_49861,N_49830);
nand UO_2273 (O_2273,N_49867,N_49973);
or UO_2274 (O_2274,N_49993,N_49992);
or UO_2275 (O_2275,N_49880,N_49755);
nand UO_2276 (O_2276,N_49960,N_49800);
xor UO_2277 (O_2277,N_49884,N_49935);
and UO_2278 (O_2278,N_49869,N_49834);
or UO_2279 (O_2279,N_49992,N_49979);
nand UO_2280 (O_2280,N_49905,N_49771);
nand UO_2281 (O_2281,N_49929,N_49785);
xor UO_2282 (O_2282,N_49961,N_49921);
and UO_2283 (O_2283,N_49785,N_49779);
and UO_2284 (O_2284,N_49984,N_49958);
and UO_2285 (O_2285,N_49944,N_49891);
or UO_2286 (O_2286,N_49976,N_49798);
and UO_2287 (O_2287,N_49907,N_49910);
xnor UO_2288 (O_2288,N_49959,N_49954);
nor UO_2289 (O_2289,N_49766,N_49998);
nor UO_2290 (O_2290,N_49973,N_49882);
and UO_2291 (O_2291,N_49887,N_49905);
xnor UO_2292 (O_2292,N_49884,N_49832);
nor UO_2293 (O_2293,N_49844,N_49854);
and UO_2294 (O_2294,N_49894,N_49778);
nand UO_2295 (O_2295,N_49908,N_49833);
nand UO_2296 (O_2296,N_49875,N_49795);
or UO_2297 (O_2297,N_49838,N_49803);
or UO_2298 (O_2298,N_49947,N_49965);
and UO_2299 (O_2299,N_49871,N_49916);
xnor UO_2300 (O_2300,N_49803,N_49805);
or UO_2301 (O_2301,N_49968,N_49803);
xor UO_2302 (O_2302,N_49965,N_49974);
or UO_2303 (O_2303,N_49943,N_49801);
xnor UO_2304 (O_2304,N_49908,N_49802);
nand UO_2305 (O_2305,N_49834,N_49859);
or UO_2306 (O_2306,N_49852,N_49866);
or UO_2307 (O_2307,N_49863,N_49960);
xnor UO_2308 (O_2308,N_49833,N_49898);
xor UO_2309 (O_2309,N_49971,N_49847);
xor UO_2310 (O_2310,N_49813,N_49842);
nand UO_2311 (O_2311,N_49794,N_49981);
and UO_2312 (O_2312,N_49919,N_49861);
nor UO_2313 (O_2313,N_49996,N_49960);
nand UO_2314 (O_2314,N_49859,N_49925);
nor UO_2315 (O_2315,N_49869,N_49932);
and UO_2316 (O_2316,N_49798,N_49891);
nand UO_2317 (O_2317,N_49832,N_49855);
and UO_2318 (O_2318,N_49811,N_49862);
nand UO_2319 (O_2319,N_49968,N_49942);
and UO_2320 (O_2320,N_49805,N_49980);
xor UO_2321 (O_2321,N_49996,N_49918);
or UO_2322 (O_2322,N_49934,N_49813);
nand UO_2323 (O_2323,N_49801,N_49994);
nor UO_2324 (O_2324,N_49841,N_49998);
nor UO_2325 (O_2325,N_49788,N_49899);
and UO_2326 (O_2326,N_49995,N_49998);
nor UO_2327 (O_2327,N_49900,N_49759);
or UO_2328 (O_2328,N_49966,N_49932);
and UO_2329 (O_2329,N_49754,N_49908);
nand UO_2330 (O_2330,N_49923,N_49875);
nor UO_2331 (O_2331,N_49902,N_49921);
nor UO_2332 (O_2332,N_49823,N_49989);
and UO_2333 (O_2333,N_49879,N_49863);
nand UO_2334 (O_2334,N_49985,N_49892);
or UO_2335 (O_2335,N_49935,N_49881);
and UO_2336 (O_2336,N_49820,N_49936);
xnor UO_2337 (O_2337,N_49959,N_49844);
nand UO_2338 (O_2338,N_49843,N_49953);
or UO_2339 (O_2339,N_49832,N_49942);
xor UO_2340 (O_2340,N_49974,N_49865);
nand UO_2341 (O_2341,N_49901,N_49922);
nand UO_2342 (O_2342,N_49864,N_49835);
nor UO_2343 (O_2343,N_49934,N_49880);
and UO_2344 (O_2344,N_49980,N_49931);
nand UO_2345 (O_2345,N_49864,N_49807);
and UO_2346 (O_2346,N_49962,N_49883);
nor UO_2347 (O_2347,N_49999,N_49845);
nand UO_2348 (O_2348,N_49915,N_49918);
or UO_2349 (O_2349,N_49837,N_49999);
nor UO_2350 (O_2350,N_49997,N_49848);
and UO_2351 (O_2351,N_49976,N_49793);
nand UO_2352 (O_2352,N_49937,N_49788);
and UO_2353 (O_2353,N_49970,N_49933);
nor UO_2354 (O_2354,N_49764,N_49900);
xnor UO_2355 (O_2355,N_49807,N_49988);
nand UO_2356 (O_2356,N_49806,N_49995);
xor UO_2357 (O_2357,N_49779,N_49976);
or UO_2358 (O_2358,N_49772,N_49890);
or UO_2359 (O_2359,N_49793,N_49928);
xnor UO_2360 (O_2360,N_49932,N_49889);
or UO_2361 (O_2361,N_49826,N_49962);
nand UO_2362 (O_2362,N_49772,N_49899);
or UO_2363 (O_2363,N_49972,N_49867);
xor UO_2364 (O_2364,N_49769,N_49881);
or UO_2365 (O_2365,N_49939,N_49793);
or UO_2366 (O_2366,N_49922,N_49830);
and UO_2367 (O_2367,N_49908,N_49909);
and UO_2368 (O_2368,N_49987,N_49988);
or UO_2369 (O_2369,N_49914,N_49937);
and UO_2370 (O_2370,N_49872,N_49822);
nand UO_2371 (O_2371,N_49880,N_49864);
nand UO_2372 (O_2372,N_49947,N_49974);
xor UO_2373 (O_2373,N_49879,N_49816);
xnor UO_2374 (O_2374,N_49907,N_49755);
xnor UO_2375 (O_2375,N_49949,N_49811);
nand UO_2376 (O_2376,N_49878,N_49888);
or UO_2377 (O_2377,N_49785,N_49953);
or UO_2378 (O_2378,N_49877,N_49906);
nor UO_2379 (O_2379,N_49759,N_49824);
nor UO_2380 (O_2380,N_49944,N_49970);
nand UO_2381 (O_2381,N_49826,N_49775);
or UO_2382 (O_2382,N_49893,N_49754);
nor UO_2383 (O_2383,N_49974,N_49983);
xnor UO_2384 (O_2384,N_49817,N_49992);
or UO_2385 (O_2385,N_49976,N_49873);
or UO_2386 (O_2386,N_49937,N_49857);
xnor UO_2387 (O_2387,N_49871,N_49940);
nand UO_2388 (O_2388,N_49754,N_49830);
nand UO_2389 (O_2389,N_49926,N_49752);
nor UO_2390 (O_2390,N_49969,N_49854);
and UO_2391 (O_2391,N_49751,N_49873);
nand UO_2392 (O_2392,N_49754,N_49833);
nor UO_2393 (O_2393,N_49763,N_49891);
or UO_2394 (O_2394,N_49818,N_49965);
nand UO_2395 (O_2395,N_49834,N_49784);
xnor UO_2396 (O_2396,N_49978,N_49836);
and UO_2397 (O_2397,N_49807,N_49770);
or UO_2398 (O_2398,N_49834,N_49830);
or UO_2399 (O_2399,N_49884,N_49801);
xor UO_2400 (O_2400,N_49836,N_49776);
or UO_2401 (O_2401,N_49926,N_49816);
xor UO_2402 (O_2402,N_49846,N_49751);
or UO_2403 (O_2403,N_49793,N_49772);
and UO_2404 (O_2404,N_49940,N_49970);
xor UO_2405 (O_2405,N_49944,N_49765);
nand UO_2406 (O_2406,N_49841,N_49912);
nor UO_2407 (O_2407,N_49809,N_49994);
or UO_2408 (O_2408,N_49846,N_49972);
nand UO_2409 (O_2409,N_49883,N_49867);
xor UO_2410 (O_2410,N_49806,N_49814);
nand UO_2411 (O_2411,N_49776,N_49966);
nor UO_2412 (O_2412,N_49954,N_49987);
or UO_2413 (O_2413,N_49968,N_49951);
or UO_2414 (O_2414,N_49954,N_49782);
nor UO_2415 (O_2415,N_49809,N_49963);
nand UO_2416 (O_2416,N_49827,N_49929);
or UO_2417 (O_2417,N_49869,N_49914);
nand UO_2418 (O_2418,N_49880,N_49753);
or UO_2419 (O_2419,N_49808,N_49788);
and UO_2420 (O_2420,N_49817,N_49766);
nand UO_2421 (O_2421,N_49938,N_49889);
nor UO_2422 (O_2422,N_49833,N_49887);
and UO_2423 (O_2423,N_49960,N_49953);
and UO_2424 (O_2424,N_49915,N_49822);
or UO_2425 (O_2425,N_49819,N_49750);
and UO_2426 (O_2426,N_49909,N_49999);
or UO_2427 (O_2427,N_49890,N_49967);
nor UO_2428 (O_2428,N_49787,N_49816);
or UO_2429 (O_2429,N_49812,N_49859);
xnor UO_2430 (O_2430,N_49850,N_49898);
nor UO_2431 (O_2431,N_49850,N_49901);
and UO_2432 (O_2432,N_49862,N_49807);
or UO_2433 (O_2433,N_49785,N_49820);
and UO_2434 (O_2434,N_49940,N_49764);
or UO_2435 (O_2435,N_49846,N_49995);
nor UO_2436 (O_2436,N_49935,N_49828);
xnor UO_2437 (O_2437,N_49788,N_49948);
nor UO_2438 (O_2438,N_49782,N_49834);
nand UO_2439 (O_2439,N_49849,N_49804);
nor UO_2440 (O_2440,N_49867,N_49868);
nor UO_2441 (O_2441,N_49923,N_49961);
or UO_2442 (O_2442,N_49925,N_49798);
xor UO_2443 (O_2443,N_49995,N_49757);
and UO_2444 (O_2444,N_49857,N_49855);
or UO_2445 (O_2445,N_49825,N_49838);
nor UO_2446 (O_2446,N_49992,N_49839);
nand UO_2447 (O_2447,N_49908,N_49884);
or UO_2448 (O_2448,N_49855,N_49869);
nor UO_2449 (O_2449,N_49942,N_49868);
nor UO_2450 (O_2450,N_49816,N_49899);
or UO_2451 (O_2451,N_49789,N_49825);
and UO_2452 (O_2452,N_49864,N_49791);
or UO_2453 (O_2453,N_49866,N_49936);
nand UO_2454 (O_2454,N_49883,N_49766);
xor UO_2455 (O_2455,N_49880,N_49811);
xor UO_2456 (O_2456,N_49994,N_49858);
xnor UO_2457 (O_2457,N_49841,N_49949);
or UO_2458 (O_2458,N_49751,N_49778);
or UO_2459 (O_2459,N_49918,N_49922);
or UO_2460 (O_2460,N_49949,N_49888);
nor UO_2461 (O_2461,N_49893,N_49786);
and UO_2462 (O_2462,N_49864,N_49824);
nand UO_2463 (O_2463,N_49878,N_49855);
xnor UO_2464 (O_2464,N_49797,N_49883);
and UO_2465 (O_2465,N_49823,N_49935);
or UO_2466 (O_2466,N_49834,N_49835);
and UO_2467 (O_2467,N_49896,N_49987);
and UO_2468 (O_2468,N_49803,N_49843);
or UO_2469 (O_2469,N_49782,N_49914);
nor UO_2470 (O_2470,N_49888,N_49824);
or UO_2471 (O_2471,N_49974,N_49940);
nor UO_2472 (O_2472,N_49863,N_49809);
and UO_2473 (O_2473,N_49970,N_49872);
xor UO_2474 (O_2474,N_49830,N_49907);
xnor UO_2475 (O_2475,N_49821,N_49832);
xor UO_2476 (O_2476,N_49863,N_49836);
or UO_2477 (O_2477,N_49760,N_49918);
xnor UO_2478 (O_2478,N_49970,N_49885);
xnor UO_2479 (O_2479,N_49845,N_49965);
xnor UO_2480 (O_2480,N_49818,N_49909);
nand UO_2481 (O_2481,N_49884,N_49753);
or UO_2482 (O_2482,N_49764,N_49980);
nor UO_2483 (O_2483,N_49774,N_49908);
and UO_2484 (O_2484,N_49882,N_49877);
or UO_2485 (O_2485,N_49832,N_49916);
and UO_2486 (O_2486,N_49842,N_49868);
xor UO_2487 (O_2487,N_49826,N_49929);
xnor UO_2488 (O_2488,N_49877,N_49938);
or UO_2489 (O_2489,N_49846,N_49998);
and UO_2490 (O_2490,N_49827,N_49837);
and UO_2491 (O_2491,N_49848,N_49799);
and UO_2492 (O_2492,N_49994,N_49850);
and UO_2493 (O_2493,N_49913,N_49860);
xor UO_2494 (O_2494,N_49960,N_49967);
nor UO_2495 (O_2495,N_49865,N_49848);
or UO_2496 (O_2496,N_49867,N_49760);
nor UO_2497 (O_2497,N_49897,N_49950);
nand UO_2498 (O_2498,N_49960,N_49821);
nand UO_2499 (O_2499,N_49840,N_49988);
and UO_2500 (O_2500,N_49829,N_49805);
xor UO_2501 (O_2501,N_49820,N_49932);
nand UO_2502 (O_2502,N_49886,N_49907);
nor UO_2503 (O_2503,N_49851,N_49881);
xnor UO_2504 (O_2504,N_49912,N_49818);
or UO_2505 (O_2505,N_49944,N_49989);
nand UO_2506 (O_2506,N_49940,N_49924);
nand UO_2507 (O_2507,N_49790,N_49977);
and UO_2508 (O_2508,N_49812,N_49973);
and UO_2509 (O_2509,N_49864,N_49778);
xor UO_2510 (O_2510,N_49824,N_49817);
nor UO_2511 (O_2511,N_49876,N_49818);
xor UO_2512 (O_2512,N_49819,N_49776);
or UO_2513 (O_2513,N_49863,N_49888);
nor UO_2514 (O_2514,N_49962,N_49937);
nand UO_2515 (O_2515,N_49837,N_49942);
nor UO_2516 (O_2516,N_49963,N_49806);
nor UO_2517 (O_2517,N_49884,N_49847);
and UO_2518 (O_2518,N_49918,N_49757);
and UO_2519 (O_2519,N_49785,N_49833);
and UO_2520 (O_2520,N_49869,N_49823);
and UO_2521 (O_2521,N_49891,N_49985);
xnor UO_2522 (O_2522,N_49804,N_49755);
nand UO_2523 (O_2523,N_49813,N_49884);
or UO_2524 (O_2524,N_49775,N_49751);
and UO_2525 (O_2525,N_49756,N_49861);
nor UO_2526 (O_2526,N_49826,N_49932);
nand UO_2527 (O_2527,N_49843,N_49919);
nand UO_2528 (O_2528,N_49905,N_49757);
and UO_2529 (O_2529,N_49785,N_49850);
nand UO_2530 (O_2530,N_49895,N_49764);
or UO_2531 (O_2531,N_49796,N_49952);
nand UO_2532 (O_2532,N_49803,N_49873);
or UO_2533 (O_2533,N_49908,N_49850);
nor UO_2534 (O_2534,N_49879,N_49759);
nor UO_2535 (O_2535,N_49847,N_49774);
or UO_2536 (O_2536,N_49829,N_49890);
nor UO_2537 (O_2537,N_49773,N_49816);
or UO_2538 (O_2538,N_49839,N_49922);
or UO_2539 (O_2539,N_49807,N_49991);
nand UO_2540 (O_2540,N_49777,N_49844);
nand UO_2541 (O_2541,N_49807,N_49872);
nor UO_2542 (O_2542,N_49860,N_49827);
or UO_2543 (O_2543,N_49970,N_49829);
nor UO_2544 (O_2544,N_49757,N_49940);
or UO_2545 (O_2545,N_49983,N_49965);
and UO_2546 (O_2546,N_49949,N_49989);
and UO_2547 (O_2547,N_49814,N_49864);
and UO_2548 (O_2548,N_49800,N_49935);
xnor UO_2549 (O_2549,N_49914,N_49972);
and UO_2550 (O_2550,N_49807,N_49819);
nor UO_2551 (O_2551,N_49883,N_49914);
or UO_2552 (O_2552,N_49885,N_49949);
or UO_2553 (O_2553,N_49804,N_49894);
nor UO_2554 (O_2554,N_49956,N_49889);
nand UO_2555 (O_2555,N_49779,N_49836);
and UO_2556 (O_2556,N_49998,N_49925);
and UO_2557 (O_2557,N_49824,N_49800);
nor UO_2558 (O_2558,N_49911,N_49826);
nor UO_2559 (O_2559,N_49990,N_49887);
or UO_2560 (O_2560,N_49824,N_49827);
xor UO_2561 (O_2561,N_49864,N_49971);
xnor UO_2562 (O_2562,N_49830,N_49763);
xnor UO_2563 (O_2563,N_49876,N_49892);
xnor UO_2564 (O_2564,N_49800,N_49997);
nor UO_2565 (O_2565,N_49914,N_49921);
nor UO_2566 (O_2566,N_49868,N_49910);
and UO_2567 (O_2567,N_49799,N_49846);
or UO_2568 (O_2568,N_49863,N_49871);
and UO_2569 (O_2569,N_49790,N_49791);
xor UO_2570 (O_2570,N_49866,N_49930);
xor UO_2571 (O_2571,N_49774,N_49962);
xor UO_2572 (O_2572,N_49988,N_49867);
nand UO_2573 (O_2573,N_49850,N_49928);
or UO_2574 (O_2574,N_49860,N_49884);
or UO_2575 (O_2575,N_49963,N_49924);
xor UO_2576 (O_2576,N_49950,N_49780);
and UO_2577 (O_2577,N_49969,N_49785);
xor UO_2578 (O_2578,N_49762,N_49764);
nand UO_2579 (O_2579,N_49885,N_49883);
and UO_2580 (O_2580,N_49940,N_49980);
xor UO_2581 (O_2581,N_49858,N_49819);
nand UO_2582 (O_2582,N_49827,N_49930);
xor UO_2583 (O_2583,N_49997,N_49845);
nor UO_2584 (O_2584,N_49842,N_49981);
nor UO_2585 (O_2585,N_49802,N_49857);
and UO_2586 (O_2586,N_49798,N_49887);
nor UO_2587 (O_2587,N_49887,N_49956);
or UO_2588 (O_2588,N_49941,N_49750);
or UO_2589 (O_2589,N_49845,N_49757);
nor UO_2590 (O_2590,N_49809,N_49845);
nand UO_2591 (O_2591,N_49992,N_49988);
nor UO_2592 (O_2592,N_49805,N_49902);
or UO_2593 (O_2593,N_49788,N_49812);
nor UO_2594 (O_2594,N_49957,N_49824);
xor UO_2595 (O_2595,N_49969,N_49803);
nor UO_2596 (O_2596,N_49886,N_49968);
nor UO_2597 (O_2597,N_49750,N_49952);
xor UO_2598 (O_2598,N_49995,N_49943);
nand UO_2599 (O_2599,N_49825,N_49973);
and UO_2600 (O_2600,N_49899,N_49970);
nor UO_2601 (O_2601,N_49876,N_49815);
xor UO_2602 (O_2602,N_49909,N_49771);
and UO_2603 (O_2603,N_49878,N_49873);
nor UO_2604 (O_2604,N_49988,N_49942);
or UO_2605 (O_2605,N_49793,N_49895);
or UO_2606 (O_2606,N_49860,N_49812);
and UO_2607 (O_2607,N_49955,N_49885);
nand UO_2608 (O_2608,N_49775,N_49827);
or UO_2609 (O_2609,N_49893,N_49814);
nand UO_2610 (O_2610,N_49869,N_49995);
or UO_2611 (O_2611,N_49789,N_49796);
xnor UO_2612 (O_2612,N_49902,N_49877);
nor UO_2613 (O_2613,N_49765,N_49805);
and UO_2614 (O_2614,N_49819,N_49869);
xor UO_2615 (O_2615,N_49942,N_49805);
nor UO_2616 (O_2616,N_49863,N_49990);
and UO_2617 (O_2617,N_49826,N_49989);
and UO_2618 (O_2618,N_49795,N_49797);
nand UO_2619 (O_2619,N_49965,N_49879);
nand UO_2620 (O_2620,N_49969,N_49955);
nor UO_2621 (O_2621,N_49843,N_49807);
xor UO_2622 (O_2622,N_49768,N_49803);
or UO_2623 (O_2623,N_49771,N_49774);
xnor UO_2624 (O_2624,N_49936,N_49849);
xor UO_2625 (O_2625,N_49866,N_49953);
nor UO_2626 (O_2626,N_49925,N_49771);
nor UO_2627 (O_2627,N_49787,N_49840);
nor UO_2628 (O_2628,N_49863,N_49808);
or UO_2629 (O_2629,N_49816,N_49918);
xor UO_2630 (O_2630,N_49860,N_49803);
or UO_2631 (O_2631,N_49851,N_49880);
nand UO_2632 (O_2632,N_49843,N_49865);
nor UO_2633 (O_2633,N_49832,N_49891);
xnor UO_2634 (O_2634,N_49909,N_49873);
and UO_2635 (O_2635,N_49879,N_49792);
nand UO_2636 (O_2636,N_49943,N_49991);
nand UO_2637 (O_2637,N_49910,N_49943);
nand UO_2638 (O_2638,N_49760,N_49988);
xnor UO_2639 (O_2639,N_49982,N_49985);
nand UO_2640 (O_2640,N_49774,N_49919);
xnor UO_2641 (O_2641,N_49896,N_49771);
nor UO_2642 (O_2642,N_49969,N_49926);
nor UO_2643 (O_2643,N_49896,N_49990);
xor UO_2644 (O_2644,N_49783,N_49844);
nand UO_2645 (O_2645,N_49751,N_49891);
nor UO_2646 (O_2646,N_49766,N_49963);
nor UO_2647 (O_2647,N_49957,N_49892);
xor UO_2648 (O_2648,N_49901,N_49932);
xor UO_2649 (O_2649,N_49936,N_49863);
nand UO_2650 (O_2650,N_49771,N_49888);
nor UO_2651 (O_2651,N_49791,N_49804);
xnor UO_2652 (O_2652,N_49859,N_49927);
nor UO_2653 (O_2653,N_49777,N_49925);
nand UO_2654 (O_2654,N_49909,N_49758);
xor UO_2655 (O_2655,N_49754,N_49920);
or UO_2656 (O_2656,N_49847,N_49863);
and UO_2657 (O_2657,N_49874,N_49983);
xor UO_2658 (O_2658,N_49969,N_49814);
and UO_2659 (O_2659,N_49833,N_49798);
and UO_2660 (O_2660,N_49874,N_49881);
nand UO_2661 (O_2661,N_49905,N_49826);
nand UO_2662 (O_2662,N_49763,N_49960);
nor UO_2663 (O_2663,N_49770,N_49792);
nor UO_2664 (O_2664,N_49825,N_49773);
and UO_2665 (O_2665,N_49811,N_49843);
and UO_2666 (O_2666,N_49980,N_49827);
and UO_2667 (O_2667,N_49993,N_49951);
xor UO_2668 (O_2668,N_49849,N_49939);
nor UO_2669 (O_2669,N_49937,N_49766);
nand UO_2670 (O_2670,N_49934,N_49956);
xnor UO_2671 (O_2671,N_49755,N_49896);
and UO_2672 (O_2672,N_49837,N_49846);
nand UO_2673 (O_2673,N_49873,N_49793);
nor UO_2674 (O_2674,N_49914,N_49804);
and UO_2675 (O_2675,N_49906,N_49885);
or UO_2676 (O_2676,N_49919,N_49872);
nor UO_2677 (O_2677,N_49917,N_49814);
xnor UO_2678 (O_2678,N_49924,N_49829);
or UO_2679 (O_2679,N_49758,N_49812);
xnor UO_2680 (O_2680,N_49949,N_49990);
nor UO_2681 (O_2681,N_49885,N_49903);
nand UO_2682 (O_2682,N_49937,N_49958);
xor UO_2683 (O_2683,N_49991,N_49945);
nor UO_2684 (O_2684,N_49760,N_49798);
and UO_2685 (O_2685,N_49978,N_49878);
or UO_2686 (O_2686,N_49808,N_49991);
or UO_2687 (O_2687,N_49820,N_49890);
nand UO_2688 (O_2688,N_49845,N_49930);
or UO_2689 (O_2689,N_49809,N_49820);
nand UO_2690 (O_2690,N_49876,N_49924);
nand UO_2691 (O_2691,N_49955,N_49895);
and UO_2692 (O_2692,N_49943,N_49955);
nor UO_2693 (O_2693,N_49917,N_49856);
nor UO_2694 (O_2694,N_49821,N_49845);
or UO_2695 (O_2695,N_49769,N_49921);
nand UO_2696 (O_2696,N_49882,N_49812);
and UO_2697 (O_2697,N_49900,N_49985);
nand UO_2698 (O_2698,N_49973,N_49920);
and UO_2699 (O_2699,N_49964,N_49812);
and UO_2700 (O_2700,N_49835,N_49782);
nand UO_2701 (O_2701,N_49941,N_49868);
and UO_2702 (O_2702,N_49962,N_49951);
nand UO_2703 (O_2703,N_49883,N_49922);
or UO_2704 (O_2704,N_49931,N_49760);
nand UO_2705 (O_2705,N_49998,N_49781);
xor UO_2706 (O_2706,N_49992,N_49920);
or UO_2707 (O_2707,N_49887,N_49996);
or UO_2708 (O_2708,N_49854,N_49850);
or UO_2709 (O_2709,N_49933,N_49939);
and UO_2710 (O_2710,N_49964,N_49883);
xor UO_2711 (O_2711,N_49959,N_49895);
xnor UO_2712 (O_2712,N_49755,N_49773);
nor UO_2713 (O_2713,N_49992,N_49830);
nand UO_2714 (O_2714,N_49990,N_49925);
nor UO_2715 (O_2715,N_49910,N_49904);
nor UO_2716 (O_2716,N_49810,N_49764);
xnor UO_2717 (O_2717,N_49759,N_49936);
or UO_2718 (O_2718,N_49876,N_49922);
and UO_2719 (O_2719,N_49881,N_49778);
or UO_2720 (O_2720,N_49969,N_49904);
nor UO_2721 (O_2721,N_49765,N_49880);
xor UO_2722 (O_2722,N_49838,N_49815);
nand UO_2723 (O_2723,N_49768,N_49974);
nor UO_2724 (O_2724,N_49795,N_49997);
and UO_2725 (O_2725,N_49877,N_49829);
and UO_2726 (O_2726,N_49774,N_49893);
nand UO_2727 (O_2727,N_49800,N_49895);
nor UO_2728 (O_2728,N_49847,N_49844);
and UO_2729 (O_2729,N_49796,N_49819);
and UO_2730 (O_2730,N_49872,N_49988);
or UO_2731 (O_2731,N_49797,N_49765);
nor UO_2732 (O_2732,N_49815,N_49873);
and UO_2733 (O_2733,N_49807,N_49947);
xor UO_2734 (O_2734,N_49766,N_49952);
nand UO_2735 (O_2735,N_49962,N_49758);
nand UO_2736 (O_2736,N_49847,N_49985);
and UO_2737 (O_2737,N_49985,N_49911);
nor UO_2738 (O_2738,N_49944,N_49995);
nor UO_2739 (O_2739,N_49962,N_49908);
xnor UO_2740 (O_2740,N_49760,N_49896);
nand UO_2741 (O_2741,N_49999,N_49865);
nor UO_2742 (O_2742,N_49889,N_49825);
xnor UO_2743 (O_2743,N_49761,N_49847);
nand UO_2744 (O_2744,N_49788,N_49855);
xnor UO_2745 (O_2745,N_49983,N_49966);
nor UO_2746 (O_2746,N_49886,N_49926);
xnor UO_2747 (O_2747,N_49888,N_49983);
nor UO_2748 (O_2748,N_49946,N_49981);
nor UO_2749 (O_2749,N_49918,N_49869);
xor UO_2750 (O_2750,N_49807,N_49785);
xor UO_2751 (O_2751,N_49994,N_49979);
nand UO_2752 (O_2752,N_49876,N_49769);
xor UO_2753 (O_2753,N_49959,N_49995);
and UO_2754 (O_2754,N_49827,N_49786);
nand UO_2755 (O_2755,N_49967,N_49837);
nor UO_2756 (O_2756,N_49869,N_49915);
or UO_2757 (O_2757,N_49841,N_49985);
nand UO_2758 (O_2758,N_49826,N_49783);
nand UO_2759 (O_2759,N_49864,N_49895);
and UO_2760 (O_2760,N_49965,N_49894);
and UO_2761 (O_2761,N_49844,N_49862);
and UO_2762 (O_2762,N_49884,N_49909);
and UO_2763 (O_2763,N_49828,N_49842);
or UO_2764 (O_2764,N_49876,N_49756);
nand UO_2765 (O_2765,N_49781,N_49914);
or UO_2766 (O_2766,N_49791,N_49905);
nor UO_2767 (O_2767,N_49919,N_49794);
nand UO_2768 (O_2768,N_49999,N_49854);
or UO_2769 (O_2769,N_49904,N_49772);
nor UO_2770 (O_2770,N_49867,N_49798);
nor UO_2771 (O_2771,N_49852,N_49980);
nor UO_2772 (O_2772,N_49837,N_49826);
nand UO_2773 (O_2773,N_49909,N_49848);
nor UO_2774 (O_2774,N_49968,N_49778);
and UO_2775 (O_2775,N_49894,N_49922);
nor UO_2776 (O_2776,N_49821,N_49943);
nor UO_2777 (O_2777,N_49993,N_49916);
and UO_2778 (O_2778,N_49922,N_49940);
nor UO_2779 (O_2779,N_49795,N_49965);
or UO_2780 (O_2780,N_49809,N_49778);
xor UO_2781 (O_2781,N_49848,N_49785);
and UO_2782 (O_2782,N_49767,N_49840);
nand UO_2783 (O_2783,N_49949,N_49803);
xnor UO_2784 (O_2784,N_49967,N_49776);
xnor UO_2785 (O_2785,N_49807,N_49781);
or UO_2786 (O_2786,N_49931,N_49858);
and UO_2787 (O_2787,N_49805,N_49876);
nor UO_2788 (O_2788,N_49948,N_49970);
xnor UO_2789 (O_2789,N_49837,N_49948);
xor UO_2790 (O_2790,N_49856,N_49779);
nand UO_2791 (O_2791,N_49926,N_49791);
or UO_2792 (O_2792,N_49798,N_49950);
nand UO_2793 (O_2793,N_49982,N_49949);
nor UO_2794 (O_2794,N_49871,N_49988);
xor UO_2795 (O_2795,N_49957,N_49871);
xor UO_2796 (O_2796,N_49919,N_49764);
or UO_2797 (O_2797,N_49989,N_49751);
xnor UO_2798 (O_2798,N_49813,N_49978);
xor UO_2799 (O_2799,N_49821,N_49858);
xnor UO_2800 (O_2800,N_49800,N_49980);
and UO_2801 (O_2801,N_49823,N_49827);
xor UO_2802 (O_2802,N_49917,N_49801);
nand UO_2803 (O_2803,N_49848,N_49826);
nand UO_2804 (O_2804,N_49896,N_49943);
xnor UO_2805 (O_2805,N_49954,N_49908);
and UO_2806 (O_2806,N_49867,N_49751);
and UO_2807 (O_2807,N_49948,N_49790);
or UO_2808 (O_2808,N_49914,N_49794);
xor UO_2809 (O_2809,N_49853,N_49899);
nor UO_2810 (O_2810,N_49808,N_49948);
and UO_2811 (O_2811,N_49991,N_49938);
xor UO_2812 (O_2812,N_49787,N_49988);
xor UO_2813 (O_2813,N_49825,N_49813);
or UO_2814 (O_2814,N_49879,N_49968);
nand UO_2815 (O_2815,N_49960,N_49822);
and UO_2816 (O_2816,N_49917,N_49946);
xor UO_2817 (O_2817,N_49907,N_49899);
or UO_2818 (O_2818,N_49919,N_49787);
nor UO_2819 (O_2819,N_49815,N_49946);
and UO_2820 (O_2820,N_49885,N_49960);
nor UO_2821 (O_2821,N_49769,N_49821);
or UO_2822 (O_2822,N_49857,N_49872);
or UO_2823 (O_2823,N_49877,N_49776);
or UO_2824 (O_2824,N_49953,N_49909);
and UO_2825 (O_2825,N_49904,N_49767);
or UO_2826 (O_2826,N_49803,N_49982);
nand UO_2827 (O_2827,N_49920,N_49916);
and UO_2828 (O_2828,N_49900,N_49779);
nand UO_2829 (O_2829,N_49754,N_49909);
xnor UO_2830 (O_2830,N_49828,N_49864);
and UO_2831 (O_2831,N_49763,N_49950);
and UO_2832 (O_2832,N_49967,N_49903);
xor UO_2833 (O_2833,N_49989,N_49837);
or UO_2834 (O_2834,N_49891,N_49879);
xnor UO_2835 (O_2835,N_49883,N_49886);
nor UO_2836 (O_2836,N_49899,N_49885);
nor UO_2837 (O_2837,N_49909,N_49938);
xor UO_2838 (O_2838,N_49939,N_49929);
or UO_2839 (O_2839,N_49851,N_49826);
nor UO_2840 (O_2840,N_49853,N_49898);
xor UO_2841 (O_2841,N_49766,N_49961);
xnor UO_2842 (O_2842,N_49932,N_49875);
nor UO_2843 (O_2843,N_49809,N_49977);
or UO_2844 (O_2844,N_49855,N_49810);
and UO_2845 (O_2845,N_49751,N_49814);
xor UO_2846 (O_2846,N_49833,N_49917);
nor UO_2847 (O_2847,N_49827,N_49893);
and UO_2848 (O_2848,N_49879,N_49827);
nor UO_2849 (O_2849,N_49995,N_49756);
nand UO_2850 (O_2850,N_49922,N_49869);
and UO_2851 (O_2851,N_49868,N_49862);
nand UO_2852 (O_2852,N_49929,N_49923);
and UO_2853 (O_2853,N_49869,N_49885);
nor UO_2854 (O_2854,N_49871,N_49894);
and UO_2855 (O_2855,N_49832,N_49992);
nand UO_2856 (O_2856,N_49917,N_49931);
or UO_2857 (O_2857,N_49957,N_49985);
nor UO_2858 (O_2858,N_49912,N_49886);
nor UO_2859 (O_2859,N_49795,N_49769);
nand UO_2860 (O_2860,N_49816,N_49932);
and UO_2861 (O_2861,N_49992,N_49922);
or UO_2862 (O_2862,N_49920,N_49850);
nor UO_2863 (O_2863,N_49984,N_49959);
and UO_2864 (O_2864,N_49828,N_49834);
or UO_2865 (O_2865,N_49873,N_49948);
nor UO_2866 (O_2866,N_49938,N_49769);
and UO_2867 (O_2867,N_49819,N_49898);
nand UO_2868 (O_2868,N_49917,N_49834);
nand UO_2869 (O_2869,N_49956,N_49984);
nand UO_2870 (O_2870,N_49890,N_49782);
nor UO_2871 (O_2871,N_49926,N_49906);
nand UO_2872 (O_2872,N_49919,N_49770);
or UO_2873 (O_2873,N_49955,N_49759);
and UO_2874 (O_2874,N_49859,N_49842);
nand UO_2875 (O_2875,N_49853,N_49809);
nor UO_2876 (O_2876,N_49752,N_49940);
and UO_2877 (O_2877,N_49850,N_49764);
xnor UO_2878 (O_2878,N_49932,N_49898);
nand UO_2879 (O_2879,N_49960,N_49808);
and UO_2880 (O_2880,N_49853,N_49900);
nor UO_2881 (O_2881,N_49870,N_49877);
xor UO_2882 (O_2882,N_49803,N_49863);
nand UO_2883 (O_2883,N_49848,N_49888);
and UO_2884 (O_2884,N_49931,N_49766);
and UO_2885 (O_2885,N_49875,N_49806);
nor UO_2886 (O_2886,N_49788,N_49795);
and UO_2887 (O_2887,N_49888,N_49948);
and UO_2888 (O_2888,N_49764,N_49915);
nor UO_2889 (O_2889,N_49816,N_49878);
and UO_2890 (O_2890,N_49974,N_49987);
nor UO_2891 (O_2891,N_49943,N_49840);
nand UO_2892 (O_2892,N_49922,N_49781);
nor UO_2893 (O_2893,N_49929,N_49999);
nor UO_2894 (O_2894,N_49797,N_49842);
or UO_2895 (O_2895,N_49820,N_49900);
and UO_2896 (O_2896,N_49775,N_49903);
or UO_2897 (O_2897,N_49959,N_49930);
xnor UO_2898 (O_2898,N_49787,N_49785);
nand UO_2899 (O_2899,N_49869,N_49813);
and UO_2900 (O_2900,N_49911,N_49865);
or UO_2901 (O_2901,N_49896,N_49931);
nand UO_2902 (O_2902,N_49786,N_49775);
xnor UO_2903 (O_2903,N_49890,N_49913);
xnor UO_2904 (O_2904,N_49766,N_49792);
or UO_2905 (O_2905,N_49815,N_49868);
nand UO_2906 (O_2906,N_49798,N_49930);
or UO_2907 (O_2907,N_49756,N_49962);
or UO_2908 (O_2908,N_49842,N_49879);
and UO_2909 (O_2909,N_49820,N_49903);
xor UO_2910 (O_2910,N_49758,N_49789);
or UO_2911 (O_2911,N_49808,N_49878);
or UO_2912 (O_2912,N_49889,N_49882);
or UO_2913 (O_2913,N_49975,N_49899);
nor UO_2914 (O_2914,N_49786,N_49869);
xnor UO_2915 (O_2915,N_49782,N_49783);
and UO_2916 (O_2916,N_49799,N_49947);
or UO_2917 (O_2917,N_49762,N_49998);
and UO_2918 (O_2918,N_49767,N_49930);
and UO_2919 (O_2919,N_49884,N_49824);
and UO_2920 (O_2920,N_49750,N_49759);
and UO_2921 (O_2921,N_49810,N_49949);
xor UO_2922 (O_2922,N_49918,N_49828);
and UO_2923 (O_2923,N_49978,N_49958);
and UO_2924 (O_2924,N_49844,N_49760);
nand UO_2925 (O_2925,N_49995,N_49909);
xor UO_2926 (O_2926,N_49830,N_49824);
or UO_2927 (O_2927,N_49805,N_49822);
and UO_2928 (O_2928,N_49797,N_49788);
or UO_2929 (O_2929,N_49937,N_49776);
xnor UO_2930 (O_2930,N_49951,N_49909);
and UO_2931 (O_2931,N_49877,N_49788);
and UO_2932 (O_2932,N_49965,N_49869);
nand UO_2933 (O_2933,N_49756,N_49878);
nor UO_2934 (O_2934,N_49954,N_49826);
or UO_2935 (O_2935,N_49839,N_49936);
nand UO_2936 (O_2936,N_49868,N_49810);
nand UO_2937 (O_2937,N_49863,N_49783);
nand UO_2938 (O_2938,N_49755,N_49840);
xnor UO_2939 (O_2939,N_49939,N_49765);
xnor UO_2940 (O_2940,N_49852,N_49860);
nand UO_2941 (O_2941,N_49863,N_49758);
or UO_2942 (O_2942,N_49760,N_49921);
nand UO_2943 (O_2943,N_49801,N_49851);
xor UO_2944 (O_2944,N_49785,N_49828);
nor UO_2945 (O_2945,N_49948,N_49767);
and UO_2946 (O_2946,N_49869,N_49804);
xor UO_2947 (O_2947,N_49854,N_49962);
nand UO_2948 (O_2948,N_49968,N_49847);
and UO_2949 (O_2949,N_49891,N_49890);
or UO_2950 (O_2950,N_49810,N_49846);
or UO_2951 (O_2951,N_49904,N_49829);
or UO_2952 (O_2952,N_49795,N_49803);
nand UO_2953 (O_2953,N_49968,N_49860);
nand UO_2954 (O_2954,N_49905,N_49847);
nor UO_2955 (O_2955,N_49758,N_49891);
and UO_2956 (O_2956,N_49839,N_49873);
nand UO_2957 (O_2957,N_49793,N_49979);
nor UO_2958 (O_2958,N_49758,N_49931);
nor UO_2959 (O_2959,N_49970,N_49994);
or UO_2960 (O_2960,N_49896,N_49829);
xor UO_2961 (O_2961,N_49982,N_49847);
xor UO_2962 (O_2962,N_49963,N_49901);
and UO_2963 (O_2963,N_49830,N_49953);
or UO_2964 (O_2964,N_49913,N_49875);
and UO_2965 (O_2965,N_49960,N_49805);
and UO_2966 (O_2966,N_49835,N_49843);
xnor UO_2967 (O_2967,N_49796,N_49943);
xnor UO_2968 (O_2968,N_49884,N_49953);
and UO_2969 (O_2969,N_49976,N_49992);
nand UO_2970 (O_2970,N_49766,N_49816);
and UO_2971 (O_2971,N_49851,N_49786);
xor UO_2972 (O_2972,N_49993,N_49985);
xnor UO_2973 (O_2973,N_49888,N_49967);
and UO_2974 (O_2974,N_49910,N_49773);
or UO_2975 (O_2975,N_49818,N_49859);
and UO_2976 (O_2976,N_49898,N_49944);
nand UO_2977 (O_2977,N_49772,N_49913);
nor UO_2978 (O_2978,N_49787,N_49965);
and UO_2979 (O_2979,N_49932,N_49917);
xnor UO_2980 (O_2980,N_49806,N_49994);
and UO_2981 (O_2981,N_49945,N_49817);
and UO_2982 (O_2982,N_49964,N_49804);
or UO_2983 (O_2983,N_49975,N_49998);
nor UO_2984 (O_2984,N_49948,N_49988);
or UO_2985 (O_2985,N_49799,N_49914);
and UO_2986 (O_2986,N_49955,N_49821);
nand UO_2987 (O_2987,N_49833,N_49873);
nor UO_2988 (O_2988,N_49801,N_49826);
and UO_2989 (O_2989,N_49881,N_49853);
or UO_2990 (O_2990,N_49892,N_49945);
nor UO_2991 (O_2991,N_49837,N_49864);
xnor UO_2992 (O_2992,N_49801,N_49986);
and UO_2993 (O_2993,N_49971,N_49950);
xnor UO_2994 (O_2994,N_49752,N_49790);
and UO_2995 (O_2995,N_49913,N_49961);
or UO_2996 (O_2996,N_49881,N_49831);
and UO_2997 (O_2997,N_49879,N_49909);
or UO_2998 (O_2998,N_49931,N_49765);
nand UO_2999 (O_2999,N_49964,N_49790);
xor UO_3000 (O_3000,N_49894,N_49972);
or UO_3001 (O_3001,N_49826,N_49843);
and UO_3002 (O_3002,N_49777,N_49868);
nor UO_3003 (O_3003,N_49842,N_49825);
nand UO_3004 (O_3004,N_49861,N_49979);
xor UO_3005 (O_3005,N_49777,N_49920);
xnor UO_3006 (O_3006,N_49893,N_49871);
and UO_3007 (O_3007,N_49936,N_49966);
xnor UO_3008 (O_3008,N_49949,N_49984);
and UO_3009 (O_3009,N_49776,N_49934);
or UO_3010 (O_3010,N_49846,N_49953);
nor UO_3011 (O_3011,N_49929,N_49976);
or UO_3012 (O_3012,N_49839,N_49783);
or UO_3013 (O_3013,N_49953,N_49836);
nor UO_3014 (O_3014,N_49916,N_49752);
or UO_3015 (O_3015,N_49869,N_49939);
xnor UO_3016 (O_3016,N_49855,N_49771);
or UO_3017 (O_3017,N_49803,N_49875);
nand UO_3018 (O_3018,N_49982,N_49785);
and UO_3019 (O_3019,N_49944,N_49882);
xnor UO_3020 (O_3020,N_49857,N_49990);
nand UO_3021 (O_3021,N_49892,N_49828);
xnor UO_3022 (O_3022,N_49896,N_49840);
or UO_3023 (O_3023,N_49858,N_49756);
and UO_3024 (O_3024,N_49943,N_49768);
nor UO_3025 (O_3025,N_49804,N_49759);
and UO_3026 (O_3026,N_49911,N_49961);
nor UO_3027 (O_3027,N_49761,N_49998);
nand UO_3028 (O_3028,N_49777,N_49879);
nand UO_3029 (O_3029,N_49785,N_49844);
and UO_3030 (O_3030,N_49795,N_49992);
and UO_3031 (O_3031,N_49776,N_49763);
and UO_3032 (O_3032,N_49875,N_49797);
nand UO_3033 (O_3033,N_49985,N_49943);
nand UO_3034 (O_3034,N_49857,N_49814);
and UO_3035 (O_3035,N_49787,N_49913);
xnor UO_3036 (O_3036,N_49806,N_49957);
nand UO_3037 (O_3037,N_49752,N_49840);
nor UO_3038 (O_3038,N_49854,N_49891);
nor UO_3039 (O_3039,N_49828,N_49906);
or UO_3040 (O_3040,N_49947,N_49954);
nand UO_3041 (O_3041,N_49872,N_49924);
or UO_3042 (O_3042,N_49959,N_49915);
nand UO_3043 (O_3043,N_49816,N_49979);
nand UO_3044 (O_3044,N_49751,N_49753);
xnor UO_3045 (O_3045,N_49915,N_49945);
xnor UO_3046 (O_3046,N_49993,N_49761);
nand UO_3047 (O_3047,N_49950,N_49993);
nand UO_3048 (O_3048,N_49894,N_49943);
xor UO_3049 (O_3049,N_49784,N_49998);
nor UO_3050 (O_3050,N_49847,N_49913);
and UO_3051 (O_3051,N_49958,N_49792);
nor UO_3052 (O_3052,N_49780,N_49908);
xnor UO_3053 (O_3053,N_49776,N_49970);
nand UO_3054 (O_3054,N_49956,N_49978);
and UO_3055 (O_3055,N_49958,N_49929);
xor UO_3056 (O_3056,N_49829,N_49870);
nor UO_3057 (O_3057,N_49938,N_49888);
nand UO_3058 (O_3058,N_49963,N_49821);
nand UO_3059 (O_3059,N_49988,N_49991);
and UO_3060 (O_3060,N_49972,N_49788);
and UO_3061 (O_3061,N_49944,N_49755);
nor UO_3062 (O_3062,N_49886,N_49759);
nor UO_3063 (O_3063,N_49920,N_49849);
or UO_3064 (O_3064,N_49923,N_49969);
nand UO_3065 (O_3065,N_49797,N_49815);
xnor UO_3066 (O_3066,N_49788,N_49789);
xnor UO_3067 (O_3067,N_49752,N_49944);
and UO_3068 (O_3068,N_49800,N_49860);
or UO_3069 (O_3069,N_49796,N_49994);
nor UO_3070 (O_3070,N_49795,N_49935);
and UO_3071 (O_3071,N_49801,N_49947);
and UO_3072 (O_3072,N_49774,N_49830);
nand UO_3073 (O_3073,N_49978,N_49936);
nand UO_3074 (O_3074,N_49972,N_49780);
nor UO_3075 (O_3075,N_49878,N_49786);
and UO_3076 (O_3076,N_49806,N_49786);
and UO_3077 (O_3077,N_49847,N_49797);
xor UO_3078 (O_3078,N_49845,N_49981);
and UO_3079 (O_3079,N_49806,N_49954);
and UO_3080 (O_3080,N_49838,N_49893);
xor UO_3081 (O_3081,N_49773,N_49846);
or UO_3082 (O_3082,N_49863,N_49800);
or UO_3083 (O_3083,N_49919,N_49765);
or UO_3084 (O_3084,N_49800,N_49963);
xnor UO_3085 (O_3085,N_49898,N_49910);
nor UO_3086 (O_3086,N_49759,N_49995);
and UO_3087 (O_3087,N_49810,N_49798);
nor UO_3088 (O_3088,N_49919,N_49928);
xnor UO_3089 (O_3089,N_49941,N_49826);
nor UO_3090 (O_3090,N_49750,N_49971);
and UO_3091 (O_3091,N_49859,N_49995);
xnor UO_3092 (O_3092,N_49948,N_49761);
and UO_3093 (O_3093,N_49963,N_49839);
xor UO_3094 (O_3094,N_49907,N_49760);
and UO_3095 (O_3095,N_49800,N_49812);
nor UO_3096 (O_3096,N_49980,N_49982);
xor UO_3097 (O_3097,N_49973,N_49987);
and UO_3098 (O_3098,N_49795,N_49811);
nand UO_3099 (O_3099,N_49897,N_49930);
and UO_3100 (O_3100,N_49924,N_49993);
or UO_3101 (O_3101,N_49766,N_49888);
nor UO_3102 (O_3102,N_49972,N_49809);
nand UO_3103 (O_3103,N_49806,N_49923);
or UO_3104 (O_3104,N_49991,N_49926);
nand UO_3105 (O_3105,N_49892,N_49903);
and UO_3106 (O_3106,N_49807,N_49857);
and UO_3107 (O_3107,N_49888,N_49781);
and UO_3108 (O_3108,N_49951,N_49844);
and UO_3109 (O_3109,N_49838,N_49974);
and UO_3110 (O_3110,N_49778,N_49817);
or UO_3111 (O_3111,N_49836,N_49914);
and UO_3112 (O_3112,N_49987,N_49838);
and UO_3113 (O_3113,N_49917,N_49908);
or UO_3114 (O_3114,N_49792,N_49750);
nand UO_3115 (O_3115,N_49869,N_49762);
nor UO_3116 (O_3116,N_49914,N_49776);
nor UO_3117 (O_3117,N_49860,N_49936);
and UO_3118 (O_3118,N_49783,N_49858);
and UO_3119 (O_3119,N_49866,N_49884);
and UO_3120 (O_3120,N_49873,N_49918);
and UO_3121 (O_3121,N_49919,N_49818);
nor UO_3122 (O_3122,N_49971,N_49848);
nor UO_3123 (O_3123,N_49755,N_49976);
and UO_3124 (O_3124,N_49911,N_49884);
xor UO_3125 (O_3125,N_49763,N_49770);
xnor UO_3126 (O_3126,N_49769,N_49971);
nor UO_3127 (O_3127,N_49974,N_49996);
xor UO_3128 (O_3128,N_49819,N_49967);
xor UO_3129 (O_3129,N_49872,N_49950);
xnor UO_3130 (O_3130,N_49808,N_49946);
nor UO_3131 (O_3131,N_49811,N_49777);
nor UO_3132 (O_3132,N_49947,N_49903);
and UO_3133 (O_3133,N_49951,N_49886);
nand UO_3134 (O_3134,N_49943,N_49785);
and UO_3135 (O_3135,N_49774,N_49939);
or UO_3136 (O_3136,N_49971,N_49882);
and UO_3137 (O_3137,N_49937,N_49943);
nand UO_3138 (O_3138,N_49920,N_49873);
and UO_3139 (O_3139,N_49818,N_49807);
and UO_3140 (O_3140,N_49857,N_49859);
nor UO_3141 (O_3141,N_49809,N_49762);
and UO_3142 (O_3142,N_49806,N_49855);
nand UO_3143 (O_3143,N_49788,N_49989);
nand UO_3144 (O_3144,N_49841,N_49753);
nor UO_3145 (O_3145,N_49913,N_49949);
nand UO_3146 (O_3146,N_49889,N_49890);
xnor UO_3147 (O_3147,N_49969,N_49917);
or UO_3148 (O_3148,N_49979,N_49946);
xnor UO_3149 (O_3149,N_49920,N_49908);
nand UO_3150 (O_3150,N_49817,N_49979);
xor UO_3151 (O_3151,N_49934,N_49785);
nand UO_3152 (O_3152,N_49810,N_49844);
nor UO_3153 (O_3153,N_49952,N_49884);
nand UO_3154 (O_3154,N_49954,N_49868);
or UO_3155 (O_3155,N_49981,N_49840);
and UO_3156 (O_3156,N_49784,N_49782);
or UO_3157 (O_3157,N_49823,N_49755);
nor UO_3158 (O_3158,N_49785,N_49801);
and UO_3159 (O_3159,N_49874,N_49902);
and UO_3160 (O_3160,N_49901,N_49960);
xor UO_3161 (O_3161,N_49948,N_49845);
or UO_3162 (O_3162,N_49823,N_49796);
and UO_3163 (O_3163,N_49994,N_49820);
nor UO_3164 (O_3164,N_49888,N_49821);
nand UO_3165 (O_3165,N_49804,N_49943);
xnor UO_3166 (O_3166,N_49926,N_49773);
and UO_3167 (O_3167,N_49777,N_49781);
and UO_3168 (O_3168,N_49809,N_49821);
nand UO_3169 (O_3169,N_49892,N_49928);
nor UO_3170 (O_3170,N_49941,N_49816);
or UO_3171 (O_3171,N_49926,N_49882);
nand UO_3172 (O_3172,N_49892,N_49925);
and UO_3173 (O_3173,N_49956,N_49998);
and UO_3174 (O_3174,N_49866,N_49946);
nand UO_3175 (O_3175,N_49826,N_49994);
or UO_3176 (O_3176,N_49863,N_49880);
nor UO_3177 (O_3177,N_49858,N_49934);
nor UO_3178 (O_3178,N_49848,N_49890);
and UO_3179 (O_3179,N_49922,N_49768);
or UO_3180 (O_3180,N_49932,N_49982);
or UO_3181 (O_3181,N_49770,N_49933);
nor UO_3182 (O_3182,N_49790,N_49822);
nand UO_3183 (O_3183,N_49935,N_49799);
or UO_3184 (O_3184,N_49864,N_49931);
xor UO_3185 (O_3185,N_49786,N_49979);
nor UO_3186 (O_3186,N_49852,N_49763);
or UO_3187 (O_3187,N_49866,N_49829);
nor UO_3188 (O_3188,N_49897,N_49782);
or UO_3189 (O_3189,N_49869,N_49752);
xor UO_3190 (O_3190,N_49993,N_49837);
xor UO_3191 (O_3191,N_49857,N_49848);
xnor UO_3192 (O_3192,N_49802,N_49967);
xor UO_3193 (O_3193,N_49772,N_49950);
and UO_3194 (O_3194,N_49991,N_49815);
nand UO_3195 (O_3195,N_49928,N_49910);
nand UO_3196 (O_3196,N_49874,N_49752);
nand UO_3197 (O_3197,N_49833,N_49827);
nor UO_3198 (O_3198,N_49907,N_49917);
or UO_3199 (O_3199,N_49928,N_49819);
nand UO_3200 (O_3200,N_49796,N_49942);
nand UO_3201 (O_3201,N_49820,N_49821);
nor UO_3202 (O_3202,N_49773,N_49896);
and UO_3203 (O_3203,N_49930,N_49777);
and UO_3204 (O_3204,N_49792,N_49987);
or UO_3205 (O_3205,N_49891,N_49896);
xnor UO_3206 (O_3206,N_49969,N_49802);
nand UO_3207 (O_3207,N_49953,N_49979);
and UO_3208 (O_3208,N_49931,N_49806);
nand UO_3209 (O_3209,N_49880,N_49813);
or UO_3210 (O_3210,N_49822,N_49857);
nor UO_3211 (O_3211,N_49777,N_49774);
nand UO_3212 (O_3212,N_49942,N_49953);
xor UO_3213 (O_3213,N_49917,N_49916);
nand UO_3214 (O_3214,N_49880,N_49940);
nand UO_3215 (O_3215,N_49898,N_49890);
nor UO_3216 (O_3216,N_49895,N_49949);
or UO_3217 (O_3217,N_49947,N_49967);
nor UO_3218 (O_3218,N_49893,N_49900);
or UO_3219 (O_3219,N_49966,N_49942);
nor UO_3220 (O_3220,N_49775,N_49792);
or UO_3221 (O_3221,N_49881,N_49782);
and UO_3222 (O_3222,N_49826,N_49829);
nor UO_3223 (O_3223,N_49971,N_49937);
nor UO_3224 (O_3224,N_49924,N_49905);
or UO_3225 (O_3225,N_49843,N_49774);
nor UO_3226 (O_3226,N_49782,N_49758);
and UO_3227 (O_3227,N_49794,N_49952);
nand UO_3228 (O_3228,N_49889,N_49896);
and UO_3229 (O_3229,N_49955,N_49841);
and UO_3230 (O_3230,N_49816,N_49887);
and UO_3231 (O_3231,N_49853,N_49982);
nand UO_3232 (O_3232,N_49834,N_49855);
nor UO_3233 (O_3233,N_49977,N_49916);
and UO_3234 (O_3234,N_49762,N_49798);
and UO_3235 (O_3235,N_49897,N_49814);
and UO_3236 (O_3236,N_49813,N_49779);
nand UO_3237 (O_3237,N_49960,N_49803);
nor UO_3238 (O_3238,N_49817,N_49834);
and UO_3239 (O_3239,N_49881,N_49923);
nand UO_3240 (O_3240,N_49767,N_49872);
xor UO_3241 (O_3241,N_49950,N_49883);
nand UO_3242 (O_3242,N_49954,N_49955);
or UO_3243 (O_3243,N_49784,N_49882);
nand UO_3244 (O_3244,N_49904,N_49954);
nand UO_3245 (O_3245,N_49997,N_49887);
and UO_3246 (O_3246,N_49970,N_49844);
nor UO_3247 (O_3247,N_49897,N_49984);
or UO_3248 (O_3248,N_49809,N_49802);
and UO_3249 (O_3249,N_49925,N_49981);
xor UO_3250 (O_3250,N_49988,N_49866);
and UO_3251 (O_3251,N_49925,N_49996);
xor UO_3252 (O_3252,N_49895,N_49862);
and UO_3253 (O_3253,N_49828,N_49979);
nand UO_3254 (O_3254,N_49775,N_49978);
xor UO_3255 (O_3255,N_49861,N_49793);
or UO_3256 (O_3256,N_49986,N_49956);
nand UO_3257 (O_3257,N_49826,N_49769);
or UO_3258 (O_3258,N_49795,N_49861);
or UO_3259 (O_3259,N_49877,N_49987);
or UO_3260 (O_3260,N_49900,N_49894);
or UO_3261 (O_3261,N_49919,N_49769);
nand UO_3262 (O_3262,N_49955,N_49973);
and UO_3263 (O_3263,N_49845,N_49926);
or UO_3264 (O_3264,N_49951,N_49944);
and UO_3265 (O_3265,N_49769,N_49887);
and UO_3266 (O_3266,N_49839,N_49842);
and UO_3267 (O_3267,N_49896,N_49899);
nor UO_3268 (O_3268,N_49942,N_49986);
nand UO_3269 (O_3269,N_49805,N_49984);
nand UO_3270 (O_3270,N_49936,N_49874);
nand UO_3271 (O_3271,N_49826,N_49846);
or UO_3272 (O_3272,N_49899,N_49827);
nand UO_3273 (O_3273,N_49992,N_49950);
xor UO_3274 (O_3274,N_49829,N_49935);
nand UO_3275 (O_3275,N_49999,N_49948);
and UO_3276 (O_3276,N_49954,N_49779);
or UO_3277 (O_3277,N_49775,N_49879);
or UO_3278 (O_3278,N_49856,N_49998);
or UO_3279 (O_3279,N_49922,N_49999);
or UO_3280 (O_3280,N_49906,N_49883);
nand UO_3281 (O_3281,N_49828,N_49807);
or UO_3282 (O_3282,N_49851,N_49933);
xnor UO_3283 (O_3283,N_49827,N_49962);
nand UO_3284 (O_3284,N_49865,N_49859);
or UO_3285 (O_3285,N_49871,N_49777);
and UO_3286 (O_3286,N_49762,N_49926);
xor UO_3287 (O_3287,N_49956,N_49784);
or UO_3288 (O_3288,N_49976,N_49754);
xor UO_3289 (O_3289,N_49852,N_49925);
and UO_3290 (O_3290,N_49837,N_49862);
xor UO_3291 (O_3291,N_49898,N_49972);
xnor UO_3292 (O_3292,N_49949,N_49980);
nand UO_3293 (O_3293,N_49969,N_49989);
xnor UO_3294 (O_3294,N_49890,N_49766);
xor UO_3295 (O_3295,N_49922,N_49751);
or UO_3296 (O_3296,N_49864,N_49908);
or UO_3297 (O_3297,N_49851,N_49916);
and UO_3298 (O_3298,N_49828,N_49812);
and UO_3299 (O_3299,N_49751,N_49827);
xor UO_3300 (O_3300,N_49977,N_49826);
nor UO_3301 (O_3301,N_49994,N_49952);
nor UO_3302 (O_3302,N_49823,N_49973);
nand UO_3303 (O_3303,N_49843,N_49899);
nand UO_3304 (O_3304,N_49865,N_49760);
or UO_3305 (O_3305,N_49980,N_49914);
xor UO_3306 (O_3306,N_49913,N_49846);
xnor UO_3307 (O_3307,N_49990,N_49878);
and UO_3308 (O_3308,N_49857,N_49902);
xnor UO_3309 (O_3309,N_49908,N_49840);
or UO_3310 (O_3310,N_49892,N_49960);
xor UO_3311 (O_3311,N_49754,N_49943);
nor UO_3312 (O_3312,N_49939,N_49987);
and UO_3313 (O_3313,N_49989,N_49845);
or UO_3314 (O_3314,N_49822,N_49885);
and UO_3315 (O_3315,N_49826,N_49916);
nor UO_3316 (O_3316,N_49909,N_49866);
nand UO_3317 (O_3317,N_49901,N_49783);
and UO_3318 (O_3318,N_49796,N_49974);
xor UO_3319 (O_3319,N_49766,N_49785);
xor UO_3320 (O_3320,N_49943,N_49904);
and UO_3321 (O_3321,N_49933,N_49968);
nand UO_3322 (O_3322,N_49804,N_49811);
nor UO_3323 (O_3323,N_49975,N_49897);
nand UO_3324 (O_3324,N_49888,N_49842);
and UO_3325 (O_3325,N_49938,N_49942);
or UO_3326 (O_3326,N_49851,N_49878);
xor UO_3327 (O_3327,N_49905,N_49966);
nand UO_3328 (O_3328,N_49987,N_49993);
xor UO_3329 (O_3329,N_49980,N_49779);
nor UO_3330 (O_3330,N_49815,N_49886);
nand UO_3331 (O_3331,N_49984,N_49969);
nand UO_3332 (O_3332,N_49933,N_49985);
nor UO_3333 (O_3333,N_49958,N_49888);
nand UO_3334 (O_3334,N_49932,N_49808);
nor UO_3335 (O_3335,N_49939,N_49915);
nor UO_3336 (O_3336,N_49929,N_49838);
or UO_3337 (O_3337,N_49898,N_49878);
and UO_3338 (O_3338,N_49991,N_49813);
or UO_3339 (O_3339,N_49985,N_49757);
and UO_3340 (O_3340,N_49833,N_49978);
and UO_3341 (O_3341,N_49831,N_49772);
and UO_3342 (O_3342,N_49955,N_49996);
nor UO_3343 (O_3343,N_49947,N_49857);
nor UO_3344 (O_3344,N_49905,N_49868);
or UO_3345 (O_3345,N_49844,N_49997);
or UO_3346 (O_3346,N_49758,N_49837);
or UO_3347 (O_3347,N_49805,N_49773);
nand UO_3348 (O_3348,N_49811,N_49993);
xor UO_3349 (O_3349,N_49955,N_49927);
xnor UO_3350 (O_3350,N_49778,N_49828);
and UO_3351 (O_3351,N_49902,N_49835);
nor UO_3352 (O_3352,N_49954,N_49784);
xor UO_3353 (O_3353,N_49908,N_49804);
nor UO_3354 (O_3354,N_49824,N_49988);
nand UO_3355 (O_3355,N_49905,N_49822);
xnor UO_3356 (O_3356,N_49936,N_49961);
nand UO_3357 (O_3357,N_49914,N_49961);
xnor UO_3358 (O_3358,N_49797,N_49821);
or UO_3359 (O_3359,N_49806,N_49765);
xnor UO_3360 (O_3360,N_49842,N_49896);
nand UO_3361 (O_3361,N_49851,N_49789);
nand UO_3362 (O_3362,N_49851,N_49848);
nor UO_3363 (O_3363,N_49775,N_49767);
nor UO_3364 (O_3364,N_49802,N_49803);
nor UO_3365 (O_3365,N_49834,N_49988);
nor UO_3366 (O_3366,N_49889,N_49989);
or UO_3367 (O_3367,N_49792,N_49898);
nor UO_3368 (O_3368,N_49834,N_49909);
xor UO_3369 (O_3369,N_49836,N_49971);
xor UO_3370 (O_3370,N_49971,N_49964);
nand UO_3371 (O_3371,N_49830,N_49962);
or UO_3372 (O_3372,N_49906,N_49859);
or UO_3373 (O_3373,N_49970,N_49950);
and UO_3374 (O_3374,N_49991,N_49773);
and UO_3375 (O_3375,N_49881,N_49918);
or UO_3376 (O_3376,N_49913,N_49841);
xnor UO_3377 (O_3377,N_49813,N_49890);
xnor UO_3378 (O_3378,N_49980,N_49887);
xor UO_3379 (O_3379,N_49798,N_49902);
nand UO_3380 (O_3380,N_49965,N_49781);
xor UO_3381 (O_3381,N_49962,N_49815);
nor UO_3382 (O_3382,N_49842,N_49832);
or UO_3383 (O_3383,N_49870,N_49781);
nand UO_3384 (O_3384,N_49962,N_49819);
and UO_3385 (O_3385,N_49860,N_49787);
and UO_3386 (O_3386,N_49997,N_49837);
nand UO_3387 (O_3387,N_49810,N_49939);
nor UO_3388 (O_3388,N_49991,N_49852);
xnor UO_3389 (O_3389,N_49799,N_49870);
nor UO_3390 (O_3390,N_49776,N_49807);
xnor UO_3391 (O_3391,N_49757,N_49983);
xnor UO_3392 (O_3392,N_49978,N_49986);
nor UO_3393 (O_3393,N_49804,N_49932);
and UO_3394 (O_3394,N_49751,N_49788);
or UO_3395 (O_3395,N_49765,N_49989);
xnor UO_3396 (O_3396,N_49765,N_49844);
or UO_3397 (O_3397,N_49846,N_49820);
and UO_3398 (O_3398,N_49816,N_49852);
nor UO_3399 (O_3399,N_49897,N_49892);
nand UO_3400 (O_3400,N_49807,N_49950);
nor UO_3401 (O_3401,N_49883,N_49958);
xnor UO_3402 (O_3402,N_49757,N_49885);
nand UO_3403 (O_3403,N_49813,N_49764);
nor UO_3404 (O_3404,N_49967,N_49877);
and UO_3405 (O_3405,N_49810,N_49893);
or UO_3406 (O_3406,N_49930,N_49883);
or UO_3407 (O_3407,N_49954,N_49763);
xor UO_3408 (O_3408,N_49886,N_49858);
xor UO_3409 (O_3409,N_49955,N_49950);
xor UO_3410 (O_3410,N_49951,N_49798);
xnor UO_3411 (O_3411,N_49954,N_49783);
or UO_3412 (O_3412,N_49838,N_49999);
or UO_3413 (O_3413,N_49946,N_49802);
and UO_3414 (O_3414,N_49816,N_49995);
or UO_3415 (O_3415,N_49759,N_49906);
or UO_3416 (O_3416,N_49881,N_49844);
or UO_3417 (O_3417,N_49929,N_49786);
xnor UO_3418 (O_3418,N_49898,N_49873);
nor UO_3419 (O_3419,N_49819,N_49921);
and UO_3420 (O_3420,N_49829,N_49788);
and UO_3421 (O_3421,N_49941,N_49961);
nor UO_3422 (O_3422,N_49777,N_49751);
or UO_3423 (O_3423,N_49809,N_49812);
nand UO_3424 (O_3424,N_49998,N_49782);
nor UO_3425 (O_3425,N_49852,N_49982);
or UO_3426 (O_3426,N_49903,N_49758);
xnor UO_3427 (O_3427,N_49962,N_49751);
or UO_3428 (O_3428,N_49872,N_49782);
and UO_3429 (O_3429,N_49917,N_49757);
xor UO_3430 (O_3430,N_49802,N_49873);
and UO_3431 (O_3431,N_49884,N_49888);
nand UO_3432 (O_3432,N_49792,N_49954);
or UO_3433 (O_3433,N_49855,N_49760);
nor UO_3434 (O_3434,N_49919,N_49802);
xnor UO_3435 (O_3435,N_49848,N_49982);
or UO_3436 (O_3436,N_49792,N_49894);
xnor UO_3437 (O_3437,N_49893,N_49932);
nand UO_3438 (O_3438,N_49947,N_49944);
nand UO_3439 (O_3439,N_49941,N_49866);
or UO_3440 (O_3440,N_49996,N_49757);
nand UO_3441 (O_3441,N_49882,N_49915);
nand UO_3442 (O_3442,N_49992,N_49874);
or UO_3443 (O_3443,N_49966,N_49798);
and UO_3444 (O_3444,N_49954,N_49840);
nand UO_3445 (O_3445,N_49972,N_49910);
and UO_3446 (O_3446,N_49886,N_49930);
and UO_3447 (O_3447,N_49954,N_49936);
or UO_3448 (O_3448,N_49885,N_49875);
or UO_3449 (O_3449,N_49832,N_49792);
xor UO_3450 (O_3450,N_49806,N_49918);
and UO_3451 (O_3451,N_49873,N_49828);
xnor UO_3452 (O_3452,N_49820,N_49868);
or UO_3453 (O_3453,N_49884,N_49906);
xnor UO_3454 (O_3454,N_49851,N_49998);
nor UO_3455 (O_3455,N_49922,N_49895);
nand UO_3456 (O_3456,N_49876,N_49989);
nor UO_3457 (O_3457,N_49928,N_49923);
or UO_3458 (O_3458,N_49915,N_49970);
nor UO_3459 (O_3459,N_49761,N_49759);
xnor UO_3460 (O_3460,N_49818,N_49999);
and UO_3461 (O_3461,N_49898,N_49750);
xor UO_3462 (O_3462,N_49946,N_49756);
or UO_3463 (O_3463,N_49798,N_49841);
nor UO_3464 (O_3464,N_49844,N_49856);
and UO_3465 (O_3465,N_49811,N_49850);
nand UO_3466 (O_3466,N_49803,N_49899);
or UO_3467 (O_3467,N_49838,N_49958);
or UO_3468 (O_3468,N_49995,N_49771);
and UO_3469 (O_3469,N_49765,N_49782);
nand UO_3470 (O_3470,N_49988,N_49951);
nand UO_3471 (O_3471,N_49906,N_49781);
nor UO_3472 (O_3472,N_49909,N_49894);
and UO_3473 (O_3473,N_49965,N_49957);
or UO_3474 (O_3474,N_49974,N_49798);
and UO_3475 (O_3475,N_49945,N_49953);
nand UO_3476 (O_3476,N_49850,N_49827);
xor UO_3477 (O_3477,N_49987,N_49799);
or UO_3478 (O_3478,N_49938,N_49953);
or UO_3479 (O_3479,N_49866,N_49906);
xnor UO_3480 (O_3480,N_49906,N_49855);
and UO_3481 (O_3481,N_49902,N_49898);
nor UO_3482 (O_3482,N_49811,N_49830);
or UO_3483 (O_3483,N_49897,N_49893);
nor UO_3484 (O_3484,N_49892,N_49898);
nor UO_3485 (O_3485,N_49790,N_49961);
and UO_3486 (O_3486,N_49830,N_49982);
xor UO_3487 (O_3487,N_49787,N_49768);
nand UO_3488 (O_3488,N_49807,N_49992);
xnor UO_3489 (O_3489,N_49842,N_49802);
and UO_3490 (O_3490,N_49878,N_49999);
or UO_3491 (O_3491,N_49789,N_49963);
and UO_3492 (O_3492,N_49907,N_49942);
xnor UO_3493 (O_3493,N_49938,N_49993);
xnor UO_3494 (O_3494,N_49962,N_49873);
nor UO_3495 (O_3495,N_49907,N_49801);
nor UO_3496 (O_3496,N_49817,N_49960);
nand UO_3497 (O_3497,N_49980,N_49842);
nand UO_3498 (O_3498,N_49822,N_49846);
nand UO_3499 (O_3499,N_49947,N_49996);
and UO_3500 (O_3500,N_49751,N_49862);
nor UO_3501 (O_3501,N_49829,N_49931);
or UO_3502 (O_3502,N_49793,N_49785);
and UO_3503 (O_3503,N_49875,N_49860);
or UO_3504 (O_3504,N_49799,N_49922);
xor UO_3505 (O_3505,N_49837,N_49757);
xor UO_3506 (O_3506,N_49769,N_49960);
and UO_3507 (O_3507,N_49769,N_49763);
xor UO_3508 (O_3508,N_49788,N_49985);
nand UO_3509 (O_3509,N_49909,N_49878);
nand UO_3510 (O_3510,N_49891,N_49838);
nand UO_3511 (O_3511,N_49951,N_49922);
or UO_3512 (O_3512,N_49915,N_49877);
nor UO_3513 (O_3513,N_49770,N_49917);
xnor UO_3514 (O_3514,N_49783,N_49793);
and UO_3515 (O_3515,N_49967,N_49954);
and UO_3516 (O_3516,N_49782,N_49792);
xor UO_3517 (O_3517,N_49899,N_49905);
nand UO_3518 (O_3518,N_49860,N_49899);
nor UO_3519 (O_3519,N_49839,N_49935);
and UO_3520 (O_3520,N_49997,N_49999);
xnor UO_3521 (O_3521,N_49919,N_49812);
nand UO_3522 (O_3522,N_49894,N_49840);
xnor UO_3523 (O_3523,N_49750,N_49868);
nor UO_3524 (O_3524,N_49963,N_49905);
nor UO_3525 (O_3525,N_49978,N_49959);
or UO_3526 (O_3526,N_49894,N_49880);
or UO_3527 (O_3527,N_49895,N_49915);
xnor UO_3528 (O_3528,N_49982,N_49837);
xor UO_3529 (O_3529,N_49968,N_49807);
or UO_3530 (O_3530,N_49811,N_49929);
nor UO_3531 (O_3531,N_49763,N_49978);
and UO_3532 (O_3532,N_49969,N_49769);
nand UO_3533 (O_3533,N_49792,N_49930);
or UO_3534 (O_3534,N_49981,N_49949);
or UO_3535 (O_3535,N_49940,N_49998);
xnor UO_3536 (O_3536,N_49885,N_49973);
and UO_3537 (O_3537,N_49797,N_49960);
xor UO_3538 (O_3538,N_49976,N_49795);
or UO_3539 (O_3539,N_49847,N_49904);
nand UO_3540 (O_3540,N_49848,N_49936);
xor UO_3541 (O_3541,N_49879,N_49982);
or UO_3542 (O_3542,N_49923,N_49832);
nor UO_3543 (O_3543,N_49786,N_49756);
nor UO_3544 (O_3544,N_49885,N_49987);
xnor UO_3545 (O_3545,N_49922,N_49848);
xor UO_3546 (O_3546,N_49830,N_49938);
or UO_3547 (O_3547,N_49949,N_49781);
nand UO_3548 (O_3548,N_49790,N_49803);
or UO_3549 (O_3549,N_49817,N_49997);
nand UO_3550 (O_3550,N_49787,N_49926);
nor UO_3551 (O_3551,N_49937,N_49991);
nand UO_3552 (O_3552,N_49755,N_49939);
and UO_3553 (O_3553,N_49928,N_49942);
nor UO_3554 (O_3554,N_49974,N_49849);
nor UO_3555 (O_3555,N_49983,N_49897);
and UO_3556 (O_3556,N_49897,N_49832);
nor UO_3557 (O_3557,N_49865,N_49821);
or UO_3558 (O_3558,N_49953,N_49903);
nor UO_3559 (O_3559,N_49954,N_49913);
or UO_3560 (O_3560,N_49819,N_49824);
nand UO_3561 (O_3561,N_49812,N_49887);
nand UO_3562 (O_3562,N_49987,N_49822);
nor UO_3563 (O_3563,N_49854,N_49908);
and UO_3564 (O_3564,N_49810,N_49967);
or UO_3565 (O_3565,N_49970,N_49780);
or UO_3566 (O_3566,N_49905,N_49922);
xnor UO_3567 (O_3567,N_49998,N_49982);
xor UO_3568 (O_3568,N_49931,N_49986);
and UO_3569 (O_3569,N_49803,N_49806);
nand UO_3570 (O_3570,N_49870,N_49925);
nand UO_3571 (O_3571,N_49982,N_49954);
or UO_3572 (O_3572,N_49898,N_49799);
or UO_3573 (O_3573,N_49940,N_49913);
xor UO_3574 (O_3574,N_49982,N_49944);
xor UO_3575 (O_3575,N_49898,N_49751);
nand UO_3576 (O_3576,N_49788,N_49968);
nand UO_3577 (O_3577,N_49886,N_49980);
nand UO_3578 (O_3578,N_49850,N_49926);
or UO_3579 (O_3579,N_49794,N_49880);
xor UO_3580 (O_3580,N_49980,N_49763);
or UO_3581 (O_3581,N_49984,N_49918);
nor UO_3582 (O_3582,N_49951,N_49956);
nand UO_3583 (O_3583,N_49865,N_49951);
nor UO_3584 (O_3584,N_49760,N_49949);
xor UO_3585 (O_3585,N_49900,N_49987);
xnor UO_3586 (O_3586,N_49895,N_49911);
nand UO_3587 (O_3587,N_49889,N_49760);
nand UO_3588 (O_3588,N_49983,N_49976);
nand UO_3589 (O_3589,N_49865,N_49973);
nand UO_3590 (O_3590,N_49961,N_49775);
and UO_3591 (O_3591,N_49955,N_49769);
or UO_3592 (O_3592,N_49798,N_49933);
or UO_3593 (O_3593,N_49986,N_49815);
or UO_3594 (O_3594,N_49916,N_49934);
or UO_3595 (O_3595,N_49754,N_49930);
nor UO_3596 (O_3596,N_49917,N_49857);
nand UO_3597 (O_3597,N_49771,N_49816);
or UO_3598 (O_3598,N_49984,N_49911);
and UO_3599 (O_3599,N_49803,N_49892);
or UO_3600 (O_3600,N_49966,N_49792);
or UO_3601 (O_3601,N_49789,N_49850);
or UO_3602 (O_3602,N_49935,N_49889);
nor UO_3603 (O_3603,N_49822,N_49812);
or UO_3604 (O_3604,N_49897,N_49848);
xor UO_3605 (O_3605,N_49866,N_49899);
nor UO_3606 (O_3606,N_49790,N_49899);
nor UO_3607 (O_3607,N_49755,N_49918);
and UO_3608 (O_3608,N_49789,N_49922);
nor UO_3609 (O_3609,N_49908,N_49848);
or UO_3610 (O_3610,N_49935,N_49972);
and UO_3611 (O_3611,N_49831,N_49787);
nand UO_3612 (O_3612,N_49752,N_49872);
or UO_3613 (O_3613,N_49991,N_49827);
or UO_3614 (O_3614,N_49750,N_49814);
or UO_3615 (O_3615,N_49783,N_49767);
nor UO_3616 (O_3616,N_49999,N_49908);
xor UO_3617 (O_3617,N_49876,N_49771);
nor UO_3618 (O_3618,N_49987,N_49994);
nor UO_3619 (O_3619,N_49910,N_49942);
and UO_3620 (O_3620,N_49786,N_49981);
xor UO_3621 (O_3621,N_49884,N_49904);
and UO_3622 (O_3622,N_49942,N_49814);
xnor UO_3623 (O_3623,N_49924,N_49854);
and UO_3624 (O_3624,N_49860,N_49906);
or UO_3625 (O_3625,N_49936,N_49819);
and UO_3626 (O_3626,N_49830,N_49821);
xnor UO_3627 (O_3627,N_49943,N_49970);
or UO_3628 (O_3628,N_49822,N_49780);
and UO_3629 (O_3629,N_49901,N_49760);
xnor UO_3630 (O_3630,N_49782,N_49961);
or UO_3631 (O_3631,N_49802,N_49762);
or UO_3632 (O_3632,N_49807,N_49927);
nand UO_3633 (O_3633,N_49953,N_49874);
and UO_3634 (O_3634,N_49988,N_49936);
or UO_3635 (O_3635,N_49803,N_49764);
xor UO_3636 (O_3636,N_49782,N_49984);
xor UO_3637 (O_3637,N_49950,N_49791);
and UO_3638 (O_3638,N_49789,N_49898);
nor UO_3639 (O_3639,N_49801,N_49981);
nand UO_3640 (O_3640,N_49868,N_49823);
nor UO_3641 (O_3641,N_49876,N_49813);
or UO_3642 (O_3642,N_49768,N_49791);
and UO_3643 (O_3643,N_49898,N_49801);
or UO_3644 (O_3644,N_49903,N_49825);
xnor UO_3645 (O_3645,N_49863,N_49955);
and UO_3646 (O_3646,N_49823,N_49778);
or UO_3647 (O_3647,N_49756,N_49982);
and UO_3648 (O_3648,N_49757,N_49967);
nor UO_3649 (O_3649,N_49857,N_49844);
or UO_3650 (O_3650,N_49999,N_49868);
or UO_3651 (O_3651,N_49842,N_49767);
nor UO_3652 (O_3652,N_49759,N_49811);
and UO_3653 (O_3653,N_49977,N_49813);
nor UO_3654 (O_3654,N_49992,N_49843);
nor UO_3655 (O_3655,N_49799,N_49887);
nand UO_3656 (O_3656,N_49900,N_49769);
nor UO_3657 (O_3657,N_49810,N_49828);
nand UO_3658 (O_3658,N_49789,N_49770);
nor UO_3659 (O_3659,N_49889,N_49844);
and UO_3660 (O_3660,N_49759,N_49764);
or UO_3661 (O_3661,N_49792,N_49934);
xnor UO_3662 (O_3662,N_49900,N_49954);
xor UO_3663 (O_3663,N_49867,N_49873);
and UO_3664 (O_3664,N_49877,N_49949);
nand UO_3665 (O_3665,N_49895,N_49917);
nor UO_3666 (O_3666,N_49957,N_49933);
or UO_3667 (O_3667,N_49994,N_49968);
xnor UO_3668 (O_3668,N_49887,N_49879);
nor UO_3669 (O_3669,N_49987,N_49999);
nand UO_3670 (O_3670,N_49869,N_49858);
nor UO_3671 (O_3671,N_49873,N_49913);
and UO_3672 (O_3672,N_49866,N_49939);
or UO_3673 (O_3673,N_49817,N_49906);
nand UO_3674 (O_3674,N_49841,N_49997);
and UO_3675 (O_3675,N_49835,N_49880);
nand UO_3676 (O_3676,N_49951,N_49998);
and UO_3677 (O_3677,N_49815,N_49898);
nor UO_3678 (O_3678,N_49790,N_49916);
xnor UO_3679 (O_3679,N_49759,N_49971);
or UO_3680 (O_3680,N_49801,N_49800);
nand UO_3681 (O_3681,N_49817,N_49777);
nor UO_3682 (O_3682,N_49928,N_49924);
nand UO_3683 (O_3683,N_49795,N_49884);
or UO_3684 (O_3684,N_49859,N_49983);
and UO_3685 (O_3685,N_49773,N_49811);
nor UO_3686 (O_3686,N_49757,N_49855);
nand UO_3687 (O_3687,N_49919,N_49993);
xnor UO_3688 (O_3688,N_49984,N_49900);
nor UO_3689 (O_3689,N_49912,N_49910);
or UO_3690 (O_3690,N_49868,N_49943);
nand UO_3691 (O_3691,N_49944,N_49785);
and UO_3692 (O_3692,N_49971,N_49930);
nor UO_3693 (O_3693,N_49860,N_49901);
nand UO_3694 (O_3694,N_49885,N_49976);
nor UO_3695 (O_3695,N_49768,N_49759);
xnor UO_3696 (O_3696,N_49801,N_49778);
nand UO_3697 (O_3697,N_49887,N_49758);
xnor UO_3698 (O_3698,N_49981,N_49839);
nand UO_3699 (O_3699,N_49855,N_49817);
nor UO_3700 (O_3700,N_49840,N_49825);
xnor UO_3701 (O_3701,N_49904,N_49899);
xor UO_3702 (O_3702,N_49918,N_49766);
or UO_3703 (O_3703,N_49997,N_49886);
and UO_3704 (O_3704,N_49930,N_49954);
or UO_3705 (O_3705,N_49853,N_49955);
or UO_3706 (O_3706,N_49830,N_49877);
and UO_3707 (O_3707,N_49825,N_49924);
and UO_3708 (O_3708,N_49762,N_49847);
nor UO_3709 (O_3709,N_49844,N_49784);
nand UO_3710 (O_3710,N_49915,N_49829);
nand UO_3711 (O_3711,N_49895,N_49799);
nand UO_3712 (O_3712,N_49802,N_49786);
nand UO_3713 (O_3713,N_49820,N_49775);
nor UO_3714 (O_3714,N_49937,N_49922);
xnor UO_3715 (O_3715,N_49988,N_49981);
and UO_3716 (O_3716,N_49879,N_49959);
and UO_3717 (O_3717,N_49866,N_49950);
xnor UO_3718 (O_3718,N_49777,N_49847);
and UO_3719 (O_3719,N_49854,N_49752);
or UO_3720 (O_3720,N_49803,N_49961);
nand UO_3721 (O_3721,N_49812,N_49789);
or UO_3722 (O_3722,N_49874,N_49827);
xnor UO_3723 (O_3723,N_49769,N_49893);
or UO_3724 (O_3724,N_49867,N_49837);
nand UO_3725 (O_3725,N_49775,N_49875);
nand UO_3726 (O_3726,N_49978,N_49798);
nand UO_3727 (O_3727,N_49995,N_49820);
and UO_3728 (O_3728,N_49829,N_49946);
nand UO_3729 (O_3729,N_49758,N_49849);
nand UO_3730 (O_3730,N_49803,N_49974);
and UO_3731 (O_3731,N_49924,N_49884);
nand UO_3732 (O_3732,N_49936,N_49816);
and UO_3733 (O_3733,N_49984,N_49830);
nand UO_3734 (O_3734,N_49925,N_49754);
nand UO_3735 (O_3735,N_49847,N_49948);
nor UO_3736 (O_3736,N_49900,N_49994);
and UO_3737 (O_3737,N_49768,N_49965);
nand UO_3738 (O_3738,N_49772,N_49959);
or UO_3739 (O_3739,N_49840,N_49963);
nand UO_3740 (O_3740,N_49823,N_49988);
or UO_3741 (O_3741,N_49911,N_49945);
nand UO_3742 (O_3742,N_49870,N_49865);
nand UO_3743 (O_3743,N_49960,N_49900);
nand UO_3744 (O_3744,N_49990,N_49812);
nand UO_3745 (O_3745,N_49956,N_49780);
xnor UO_3746 (O_3746,N_49808,N_49767);
nor UO_3747 (O_3747,N_49801,N_49847);
and UO_3748 (O_3748,N_49918,N_49862);
nor UO_3749 (O_3749,N_49891,N_49937);
and UO_3750 (O_3750,N_49983,N_49778);
or UO_3751 (O_3751,N_49757,N_49913);
xor UO_3752 (O_3752,N_49872,N_49923);
nor UO_3753 (O_3753,N_49896,N_49918);
nand UO_3754 (O_3754,N_49858,N_49813);
xor UO_3755 (O_3755,N_49984,N_49995);
and UO_3756 (O_3756,N_49865,N_49933);
nor UO_3757 (O_3757,N_49973,N_49893);
nor UO_3758 (O_3758,N_49868,N_49827);
and UO_3759 (O_3759,N_49870,N_49831);
and UO_3760 (O_3760,N_49853,N_49966);
xnor UO_3761 (O_3761,N_49867,N_49875);
and UO_3762 (O_3762,N_49857,N_49821);
and UO_3763 (O_3763,N_49758,N_49771);
nand UO_3764 (O_3764,N_49966,N_49915);
xor UO_3765 (O_3765,N_49858,N_49754);
and UO_3766 (O_3766,N_49956,N_49801);
xnor UO_3767 (O_3767,N_49811,N_49800);
or UO_3768 (O_3768,N_49774,N_49813);
nand UO_3769 (O_3769,N_49977,N_49814);
xor UO_3770 (O_3770,N_49963,N_49930);
xor UO_3771 (O_3771,N_49791,N_49801);
nor UO_3772 (O_3772,N_49966,N_49828);
and UO_3773 (O_3773,N_49752,N_49750);
nor UO_3774 (O_3774,N_49776,N_49794);
xnor UO_3775 (O_3775,N_49991,N_49759);
and UO_3776 (O_3776,N_49757,N_49874);
nand UO_3777 (O_3777,N_49989,N_49836);
nor UO_3778 (O_3778,N_49852,N_49792);
or UO_3779 (O_3779,N_49795,N_49871);
and UO_3780 (O_3780,N_49992,N_49857);
and UO_3781 (O_3781,N_49885,N_49817);
xnor UO_3782 (O_3782,N_49868,N_49784);
and UO_3783 (O_3783,N_49839,N_49776);
nand UO_3784 (O_3784,N_49853,N_49916);
xnor UO_3785 (O_3785,N_49875,N_49980);
or UO_3786 (O_3786,N_49854,N_49923);
nand UO_3787 (O_3787,N_49800,N_49809);
xnor UO_3788 (O_3788,N_49966,N_49943);
xnor UO_3789 (O_3789,N_49874,N_49897);
nand UO_3790 (O_3790,N_49957,N_49989);
xor UO_3791 (O_3791,N_49940,N_49874);
xnor UO_3792 (O_3792,N_49937,N_49888);
nand UO_3793 (O_3793,N_49753,N_49896);
nor UO_3794 (O_3794,N_49973,N_49860);
xor UO_3795 (O_3795,N_49776,N_49956);
and UO_3796 (O_3796,N_49956,N_49854);
and UO_3797 (O_3797,N_49985,N_49820);
or UO_3798 (O_3798,N_49925,N_49903);
and UO_3799 (O_3799,N_49764,N_49968);
xor UO_3800 (O_3800,N_49945,N_49895);
nor UO_3801 (O_3801,N_49863,N_49911);
xor UO_3802 (O_3802,N_49958,N_49966);
nand UO_3803 (O_3803,N_49766,N_49775);
xnor UO_3804 (O_3804,N_49927,N_49893);
xnor UO_3805 (O_3805,N_49869,N_49981);
and UO_3806 (O_3806,N_49867,N_49825);
or UO_3807 (O_3807,N_49763,N_49764);
nand UO_3808 (O_3808,N_49935,N_49776);
and UO_3809 (O_3809,N_49974,N_49858);
and UO_3810 (O_3810,N_49880,N_49987);
nand UO_3811 (O_3811,N_49857,N_49811);
nand UO_3812 (O_3812,N_49839,N_49765);
or UO_3813 (O_3813,N_49791,N_49792);
and UO_3814 (O_3814,N_49809,N_49842);
xnor UO_3815 (O_3815,N_49902,N_49850);
or UO_3816 (O_3816,N_49804,N_49885);
nand UO_3817 (O_3817,N_49760,N_49913);
or UO_3818 (O_3818,N_49864,N_49783);
nor UO_3819 (O_3819,N_49812,N_49972);
nor UO_3820 (O_3820,N_49752,N_49891);
or UO_3821 (O_3821,N_49914,N_49933);
nor UO_3822 (O_3822,N_49886,N_49789);
and UO_3823 (O_3823,N_49969,N_49797);
xor UO_3824 (O_3824,N_49881,N_49926);
nand UO_3825 (O_3825,N_49857,N_49940);
xor UO_3826 (O_3826,N_49893,N_49864);
and UO_3827 (O_3827,N_49755,N_49868);
nand UO_3828 (O_3828,N_49781,N_49783);
and UO_3829 (O_3829,N_49870,N_49761);
or UO_3830 (O_3830,N_49836,N_49795);
and UO_3831 (O_3831,N_49944,N_49960);
and UO_3832 (O_3832,N_49809,N_49784);
nor UO_3833 (O_3833,N_49799,N_49867);
and UO_3834 (O_3834,N_49812,N_49757);
nor UO_3835 (O_3835,N_49911,N_49792);
nand UO_3836 (O_3836,N_49810,N_49922);
and UO_3837 (O_3837,N_49846,N_49919);
nand UO_3838 (O_3838,N_49839,N_49856);
nor UO_3839 (O_3839,N_49780,N_49801);
nand UO_3840 (O_3840,N_49949,N_49945);
or UO_3841 (O_3841,N_49954,N_49839);
nand UO_3842 (O_3842,N_49774,N_49789);
nor UO_3843 (O_3843,N_49912,N_49757);
nor UO_3844 (O_3844,N_49801,N_49989);
and UO_3845 (O_3845,N_49783,N_49919);
xnor UO_3846 (O_3846,N_49970,N_49827);
nor UO_3847 (O_3847,N_49845,N_49795);
or UO_3848 (O_3848,N_49838,N_49950);
xnor UO_3849 (O_3849,N_49831,N_49771);
nor UO_3850 (O_3850,N_49785,N_49892);
or UO_3851 (O_3851,N_49751,N_49991);
nand UO_3852 (O_3852,N_49949,N_49869);
xor UO_3853 (O_3853,N_49790,N_49793);
nand UO_3854 (O_3854,N_49853,N_49858);
nand UO_3855 (O_3855,N_49901,N_49801);
xor UO_3856 (O_3856,N_49856,N_49789);
or UO_3857 (O_3857,N_49759,N_49785);
or UO_3858 (O_3858,N_49985,N_49916);
or UO_3859 (O_3859,N_49982,N_49981);
or UO_3860 (O_3860,N_49757,N_49914);
nor UO_3861 (O_3861,N_49793,N_49833);
and UO_3862 (O_3862,N_49997,N_49835);
nor UO_3863 (O_3863,N_49835,N_49821);
and UO_3864 (O_3864,N_49969,N_49956);
xnor UO_3865 (O_3865,N_49897,N_49887);
nand UO_3866 (O_3866,N_49834,N_49848);
nand UO_3867 (O_3867,N_49911,N_49793);
nor UO_3868 (O_3868,N_49804,N_49777);
xor UO_3869 (O_3869,N_49834,N_49888);
or UO_3870 (O_3870,N_49826,N_49974);
and UO_3871 (O_3871,N_49999,N_49751);
nor UO_3872 (O_3872,N_49973,N_49854);
xor UO_3873 (O_3873,N_49960,N_49931);
xor UO_3874 (O_3874,N_49828,N_49811);
or UO_3875 (O_3875,N_49883,N_49984);
nand UO_3876 (O_3876,N_49791,N_49970);
or UO_3877 (O_3877,N_49755,N_49951);
or UO_3878 (O_3878,N_49908,N_49974);
and UO_3879 (O_3879,N_49875,N_49835);
xnor UO_3880 (O_3880,N_49819,N_49789);
nand UO_3881 (O_3881,N_49898,N_49786);
and UO_3882 (O_3882,N_49760,N_49883);
xnor UO_3883 (O_3883,N_49766,N_49972);
or UO_3884 (O_3884,N_49955,N_49902);
nand UO_3885 (O_3885,N_49906,N_49753);
nor UO_3886 (O_3886,N_49804,N_49834);
and UO_3887 (O_3887,N_49994,N_49975);
nor UO_3888 (O_3888,N_49982,N_49974);
xor UO_3889 (O_3889,N_49750,N_49896);
xnor UO_3890 (O_3890,N_49803,N_49757);
or UO_3891 (O_3891,N_49980,N_49903);
nand UO_3892 (O_3892,N_49893,N_49948);
nor UO_3893 (O_3893,N_49921,N_49880);
xor UO_3894 (O_3894,N_49932,N_49790);
nor UO_3895 (O_3895,N_49943,N_49860);
or UO_3896 (O_3896,N_49981,N_49886);
nand UO_3897 (O_3897,N_49960,N_49773);
or UO_3898 (O_3898,N_49806,N_49928);
nand UO_3899 (O_3899,N_49991,N_49890);
or UO_3900 (O_3900,N_49986,N_49854);
xor UO_3901 (O_3901,N_49992,N_49959);
xnor UO_3902 (O_3902,N_49933,N_49873);
nor UO_3903 (O_3903,N_49889,N_49822);
nand UO_3904 (O_3904,N_49876,N_49839);
nand UO_3905 (O_3905,N_49878,N_49976);
nor UO_3906 (O_3906,N_49831,N_49974);
and UO_3907 (O_3907,N_49906,N_49969);
and UO_3908 (O_3908,N_49927,N_49950);
nor UO_3909 (O_3909,N_49880,N_49788);
xor UO_3910 (O_3910,N_49855,N_49856);
and UO_3911 (O_3911,N_49832,N_49965);
or UO_3912 (O_3912,N_49996,N_49850);
xor UO_3913 (O_3913,N_49827,N_49769);
and UO_3914 (O_3914,N_49976,N_49996);
or UO_3915 (O_3915,N_49780,N_49963);
nor UO_3916 (O_3916,N_49766,N_49947);
and UO_3917 (O_3917,N_49770,N_49782);
nand UO_3918 (O_3918,N_49755,N_49955);
nor UO_3919 (O_3919,N_49997,N_49802);
and UO_3920 (O_3920,N_49959,N_49998);
and UO_3921 (O_3921,N_49861,N_49845);
nor UO_3922 (O_3922,N_49869,N_49827);
xor UO_3923 (O_3923,N_49913,N_49804);
and UO_3924 (O_3924,N_49944,N_49988);
and UO_3925 (O_3925,N_49938,N_49958);
nor UO_3926 (O_3926,N_49857,N_49888);
or UO_3927 (O_3927,N_49893,N_49995);
and UO_3928 (O_3928,N_49889,N_49783);
nor UO_3929 (O_3929,N_49978,N_49952);
and UO_3930 (O_3930,N_49780,N_49885);
and UO_3931 (O_3931,N_49933,N_49994);
xnor UO_3932 (O_3932,N_49941,N_49844);
and UO_3933 (O_3933,N_49835,N_49799);
xnor UO_3934 (O_3934,N_49840,N_49857);
or UO_3935 (O_3935,N_49795,N_49802);
nor UO_3936 (O_3936,N_49808,N_49759);
nor UO_3937 (O_3937,N_49780,N_49971);
nand UO_3938 (O_3938,N_49912,N_49953);
xor UO_3939 (O_3939,N_49926,N_49757);
xnor UO_3940 (O_3940,N_49753,N_49973);
nand UO_3941 (O_3941,N_49880,N_49826);
and UO_3942 (O_3942,N_49959,N_49951);
xor UO_3943 (O_3943,N_49798,N_49774);
or UO_3944 (O_3944,N_49753,N_49754);
and UO_3945 (O_3945,N_49919,N_49766);
xor UO_3946 (O_3946,N_49865,N_49841);
xnor UO_3947 (O_3947,N_49837,N_49914);
nor UO_3948 (O_3948,N_49900,N_49979);
and UO_3949 (O_3949,N_49847,N_49947);
xnor UO_3950 (O_3950,N_49918,N_49826);
nand UO_3951 (O_3951,N_49804,N_49794);
nor UO_3952 (O_3952,N_49943,N_49923);
or UO_3953 (O_3953,N_49824,N_49875);
xor UO_3954 (O_3954,N_49920,N_49796);
and UO_3955 (O_3955,N_49995,N_49751);
or UO_3956 (O_3956,N_49874,N_49885);
or UO_3957 (O_3957,N_49949,N_49812);
nand UO_3958 (O_3958,N_49811,N_49790);
nor UO_3959 (O_3959,N_49977,N_49964);
and UO_3960 (O_3960,N_49909,N_49987);
nand UO_3961 (O_3961,N_49788,N_49786);
nor UO_3962 (O_3962,N_49820,N_49823);
and UO_3963 (O_3963,N_49860,N_49854);
xor UO_3964 (O_3964,N_49814,N_49922);
xnor UO_3965 (O_3965,N_49817,N_49958);
or UO_3966 (O_3966,N_49993,N_49937);
nand UO_3967 (O_3967,N_49781,N_49819);
xnor UO_3968 (O_3968,N_49891,N_49989);
nor UO_3969 (O_3969,N_49962,N_49794);
or UO_3970 (O_3970,N_49950,N_49819);
and UO_3971 (O_3971,N_49835,N_49980);
xnor UO_3972 (O_3972,N_49851,N_49807);
nor UO_3973 (O_3973,N_49821,N_49770);
nand UO_3974 (O_3974,N_49911,N_49992);
and UO_3975 (O_3975,N_49927,N_49821);
nand UO_3976 (O_3976,N_49862,N_49816);
and UO_3977 (O_3977,N_49808,N_49756);
or UO_3978 (O_3978,N_49778,N_49833);
nand UO_3979 (O_3979,N_49814,N_49800);
or UO_3980 (O_3980,N_49779,N_49906);
xor UO_3981 (O_3981,N_49815,N_49790);
or UO_3982 (O_3982,N_49862,N_49913);
xor UO_3983 (O_3983,N_49944,N_49985);
nor UO_3984 (O_3984,N_49903,N_49764);
and UO_3985 (O_3985,N_49857,N_49858);
xor UO_3986 (O_3986,N_49781,N_49898);
xor UO_3987 (O_3987,N_49952,N_49770);
xnor UO_3988 (O_3988,N_49933,N_49776);
xnor UO_3989 (O_3989,N_49947,N_49914);
or UO_3990 (O_3990,N_49789,N_49919);
or UO_3991 (O_3991,N_49873,N_49784);
nand UO_3992 (O_3992,N_49787,N_49975);
and UO_3993 (O_3993,N_49967,N_49883);
and UO_3994 (O_3994,N_49848,N_49819);
nand UO_3995 (O_3995,N_49944,N_49990);
xnor UO_3996 (O_3996,N_49910,N_49792);
or UO_3997 (O_3997,N_49761,N_49977);
nand UO_3998 (O_3998,N_49869,N_49811);
and UO_3999 (O_3999,N_49920,N_49981);
xor UO_4000 (O_4000,N_49835,N_49977);
xnor UO_4001 (O_4001,N_49836,N_49762);
nor UO_4002 (O_4002,N_49785,N_49865);
nor UO_4003 (O_4003,N_49980,N_49959);
and UO_4004 (O_4004,N_49998,N_49774);
xor UO_4005 (O_4005,N_49779,N_49857);
xor UO_4006 (O_4006,N_49751,N_49963);
and UO_4007 (O_4007,N_49908,N_49766);
or UO_4008 (O_4008,N_49993,N_49854);
nor UO_4009 (O_4009,N_49959,N_49873);
and UO_4010 (O_4010,N_49975,N_49788);
nand UO_4011 (O_4011,N_49892,N_49881);
xor UO_4012 (O_4012,N_49942,N_49936);
xor UO_4013 (O_4013,N_49752,N_49811);
nor UO_4014 (O_4014,N_49887,N_49950);
nor UO_4015 (O_4015,N_49931,N_49782);
or UO_4016 (O_4016,N_49921,N_49824);
nor UO_4017 (O_4017,N_49956,N_49888);
xor UO_4018 (O_4018,N_49840,N_49941);
nor UO_4019 (O_4019,N_49974,N_49888);
and UO_4020 (O_4020,N_49946,N_49767);
xor UO_4021 (O_4021,N_49918,N_49768);
xor UO_4022 (O_4022,N_49754,N_49785);
xor UO_4023 (O_4023,N_49841,N_49891);
and UO_4024 (O_4024,N_49827,N_49959);
nand UO_4025 (O_4025,N_49834,N_49845);
nor UO_4026 (O_4026,N_49795,N_49948);
xor UO_4027 (O_4027,N_49941,N_49818);
or UO_4028 (O_4028,N_49847,N_49755);
nor UO_4029 (O_4029,N_49961,N_49962);
xor UO_4030 (O_4030,N_49874,N_49775);
and UO_4031 (O_4031,N_49899,N_49966);
nor UO_4032 (O_4032,N_49884,N_49978);
xnor UO_4033 (O_4033,N_49800,N_49951);
nand UO_4034 (O_4034,N_49844,N_49888);
nand UO_4035 (O_4035,N_49987,N_49769);
and UO_4036 (O_4036,N_49816,N_49755);
xnor UO_4037 (O_4037,N_49952,N_49824);
or UO_4038 (O_4038,N_49836,N_49970);
nand UO_4039 (O_4039,N_49938,N_49874);
xor UO_4040 (O_4040,N_49906,N_49772);
nor UO_4041 (O_4041,N_49883,N_49900);
nand UO_4042 (O_4042,N_49832,N_49936);
nor UO_4043 (O_4043,N_49936,N_49812);
nand UO_4044 (O_4044,N_49915,N_49900);
and UO_4045 (O_4045,N_49986,N_49894);
xor UO_4046 (O_4046,N_49897,N_49879);
nor UO_4047 (O_4047,N_49929,N_49796);
and UO_4048 (O_4048,N_49827,N_49966);
and UO_4049 (O_4049,N_49840,N_49970);
nor UO_4050 (O_4050,N_49782,N_49775);
and UO_4051 (O_4051,N_49815,N_49754);
or UO_4052 (O_4052,N_49821,N_49990);
or UO_4053 (O_4053,N_49799,N_49881);
and UO_4054 (O_4054,N_49972,N_49896);
xor UO_4055 (O_4055,N_49864,N_49922);
or UO_4056 (O_4056,N_49835,N_49794);
or UO_4057 (O_4057,N_49866,N_49910);
or UO_4058 (O_4058,N_49997,N_49750);
and UO_4059 (O_4059,N_49901,N_49787);
or UO_4060 (O_4060,N_49770,N_49935);
xnor UO_4061 (O_4061,N_49752,N_49871);
xnor UO_4062 (O_4062,N_49782,N_49761);
nor UO_4063 (O_4063,N_49896,N_49907);
xor UO_4064 (O_4064,N_49756,N_49886);
xnor UO_4065 (O_4065,N_49875,N_49872);
nand UO_4066 (O_4066,N_49955,N_49818);
nand UO_4067 (O_4067,N_49903,N_49894);
and UO_4068 (O_4068,N_49846,N_49980);
nand UO_4069 (O_4069,N_49992,N_49765);
nand UO_4070 (O_4070,N_49801,N_49992);
nor UO_4071 (O_4071,N_49848,N_49914);
xnor UO_4072 (O_4072,N_49986,N_49765);
nor UO_4073 (O_4073,N_49766,N_49830);
nand UO_4074 (O_4074,N_49856,N_49954);
xnor UO_4075 (O_4075,N_49881,N_49885);
nand UO_4076 (O_4076,N_49927,N_49988);
nand UO_4077 (O_4077,N_49846,N_49940);
nand UO_4078 (O_4078,N_49891,N_49827);
xor UO_4079 (O_4079,N_49836,N_49881);
or UO_4080 (O_4080,N_49759,N_49973);
xor UO_4081 (O_4081,N_49937,N_49910);
nor UO_4082 (O_4082,N_49770,N_49839);
and UO_4083 (O_4083,N_49882,N_49860);
nand UO_4084 (O_4084,N_49883,N_49827);
nand UO_4085 (O_4085,N_49763,N_49982);
xnor UO_4086 (O_4086,N_49983,N_49820);
and UO_4087 (O_4087,N_49918,N_49836);
nor UO_4088 (O_4088,N_49812,N_49845);
nor UO_4089 (O_4089,N_49848,N_49855);
xor UO_4090 (O_4090,N_49754,N_49788);
xor UO_4091 (O_4091,N_49852,N_49833);
and UO_4092 (O_4092,N_49966,N_49934);
xnor UO_4093 (O_4093,N_49974,N_49778);
xor UO_4094 (O_4094,N_49990,N_49813);
nor UO_4095 (O_4095,N_49962,N_49789);
xor UO_4096 (O_4096,N_49795,N_49834);
or UO_4097 (O_4097,N_49888,N_49960);
nor UO_4098 (O_4098,N_49870,N_49901);
or UO_4099 (O_4099,N_49840,N_49879);
xor UO_4100 (O_4100,N_49843,N_49753);
nor UO_4101 (O_4101,N_49788,N_49983);
nand UO_4102 (O_4102,N_49971,N_49835);
nor UO_4103 (O_4103,N_49931,N_49843);
nor UO_4104 (O_4104,N_49883,N_49876);
or UO_4105 (O_4105,N_49839,N_49945);
nand UO_4106 (O_4106,N_49774,N_49766);
nor UO_4107 (O_4107,N_49993,N_49911);
and UO_4108 (O_4108,N_49975,N_49953);
xor UO_4109 (O_4109,N_49769,N_49771);
nor UO_4110 (O_4110,N_49998,N_49824);
xor UO_4111 (O_4111,N_49907,N_49986);
nand UO_4112 (O_4112,N_49798,N_49977);
or UO_4113 (O_4113,N_49779,N_49764);
or UO_4114 (O_4114,N_49880,N_49796);
or UO_4115 (O_4115,N_49899,N_49964);
nand UO_4116 (O_4116,N_49839,N_49809);
nor UO_4117 (O_4117,N_49954,N_49918);
xor UO_4118 (O_4118,N_49938,N_49926);
nand UO_4119 (O_4119,N_49825,N_49965);
or UO_4120 (O_4120,N_49980,N_49944);
xor UO_4121 (O_4121,N_49809,N_49814);
xor UO_4122 (O_4122,N_49841,N_49843);
or UO_4123 (O_4123,N_49820,N_49818);
nor UO_4124 (O_4124,N_49879,N_49804);
and UO_4125 (O_4125,N_49976,N_49769);
nand UO_4126 (O_4126,N_49971,N_49961);
nand UO_4127 (O_4127,N_49789,N_49984);
nor UO_4128 (O_4128,N_49878,N_49981);
and UO_4129 (O_4129,N_49845,N_49852);
nand UO_4130 (O_4130,N_49919,N_49979);
or UO_4131 (O_4131,N_49760,N_49930);
xor UO_4132 (O_4132,N_49878,N_49988);
nand UO_4133 (O_4133,N_49760,N_49890);
or UO_4134 (O_4134,N_49901,N_49884);
xor UO_4135 (O_4135,N_49831,N_49786);
and UO_4136 (O_4136,N_49894,N_49764);
and UO_4137 (O_4137,N_49771,N_49963);
nand UO_4138 (O_4138,N_49841,N_49873);
or UO_4139 (O_4139,N_49793,N_49758);
and UO_4140 (O_4140,N_49981,N_49877);
xor UO_4141 (O_4141,N_49938,N_49863);
or UO_4142 (O_4142,N_49994,N_49964);
nand UO_4143 (O_4143,N_49760,N_49998);
nand UO_4144 (O_4144,N_49847,N_49817);
and UO_4145 (O_4145,N_49899,N_49976);
xor UO_4146 (O_4146,N_49750,N_49859);
xnor UO_4147 (O_4147,N_49905,N_49969);
nor UO_4148 (O_4148,N_49945,N_49999);
or UO_4149 (O_4149,N_49760,N_49817);
and UO_4150 (O_4150,N_49809,N_49816);
nor UO_4151 (O_4151,N_49914,N_49789);
and UO_4152 (O_4152,N_49986,N_49997);
and UO_4153 (O_4153,N_49870,N_49784);
and UO_4154 (O_4154,N_49879,N_49967);
and UO_4155 (O_4155,N_49909,N_49893);
xor UO_4156 (O_4156,N_49818,N_49997);
nor UO_4157 (O_4157,N_49811,N_49861);
or UO_4158 (O_4158,N_49916,N_49983);
nand UO_4159 (O_4159,N_49889,N_49804);
nor UO_4160 (O_4160,N_49773,N_49997);
or UO_4161 (O_4161,N_49751,N_49782);
xnor UO_4162 (O_4162,N_49860,N_49893);
nand UO_4163 (O_4163,N_49763,N_49805);
and UO_4164 (O_4164,N_49813,N_49784);
nor UO_4165 (O_4165,N_49885,N_49998);
nor UO_4166 (O_4166,N_49957,N_49921);
or UO_4167 (O_4167,N_49924,N_49774);
nand UO_4168 (O_4168,N_49884,N_49966);
nand UO_4169 (O_4169,N_49987,N_49862);
nand UO_4170 (O_4170,N_49983,N_49990);
xnor UO_4171 (O_4171,N_49812,N_49992);
or UO_4172 (O_4172,N_49887,N_49760);
nand UO_4173 (O_4173,N_49955,N_49941);
nor UO_4174 (O_4174,N_49839,N_49889);
nor UO_4175 (O_4175,N_49794,N_49761);
xor UO_4176 (O_4176,N_49876,N_49956);
nand UO_4177 (O_4177,N_49965,N_49808);
and UO_4178 (O_4178,N_49778,N_49953);
nor UO_4179 (O_4179,N_49795,N_49805);
or UO_4180 (O_4180,N_49937,N_49999);
nand UO_4181 (O_4181,N_49800,N_49875);
nand UO_4182 (O_4182,N_49832,N_49973);
or UO_4183 (O_4183,N_49768,N_49798);
and UO_4184 (O_4184,N_49912,N_49785);
or UO_4185 (O_4185,N_49812,N_49834);
or UO_4186 (O_4186,N_49825,N_49817);
or UO_4187 (O_4187,N_49858,N_49992);
nand UO_4188 (O_4188,N_49811,N_49992);
nand UO_4189 (O_4189,N_49781,N_49952);
nor UO_4190 (O_4190,N_49877,N_49896);
xnor UO_4191 (O_4191,N_49962,N_49969);
nor UO_4192 (O_4192,N_49921,N_49888);
nor UO_4193 (O_4193,N_49955,N_49792);
nor UO_4194 (O_4194,N_49827,N_49944);
nor UO_4195 (O_4195,N_49822,N_49909);
xnor UO_4196 (O_4196,N_49847,N_49979);
or UO_4197 (O_4197,N_49847,N_49779);
or UO_4198 (O_4198,N_49826,N_49767);
and UO_4199 (O_4199,N_49852,N_49903);
or UO_4200 (O_4200,N_49821,N_49848);
and UO_4201 (O_4201,N_49879,N_49771);
or UO_4202 (O_4202,N_49796,N_49971);
xor UO_4203 (O_4203,N_49828,N_49804);
nand UO_4204 (O_4204,N_49991,N_49828);
or UO_4205 (O_4205,N_49974,N_49909);
and UO_4206 (O_4206,N_49887,N_49903);
nand UO_4207 (O_4207,N_49988,N_49877);
and UO_4208 (O_4208,N_49902,N_49913);
and UO_4209 (O_4209,N_49756,N_49966);
xor UO_4210 (O_4210,N_49756,N_49839);
nand UO_4211 (O_4211,N_49777,N_49779);
or UO_4212 (O_4212,N_49778,N_49835);
and UO_4213 (O_4213,N_49874,N_49886);
and UO_4214 (O_4214,N_49849,N_49782);
nor UO_4215 (O_4215,N_49759,N_49981);
or UO_4216 (O_4216,N_49784,N_49937);
nor UO_4217 (O_4217,N_49976,N_49845);
or UO_4218 (O_4218,N_49768,N_49816);
nor UO_4219 (O_4219,N_49989,N_49866);
or UO_4220 (O_4220,N_49769,N_49891);
and UO_4221 (O_4221,N_49926,N_49804);
nand UO_4222 (O_4222,N_49856,N_49979);
nor UO_4223 (O_4223,N_49755,N_49765);
xor UO_4224 (O_4224,N_49771,N_49865);
xnor UO_4225 (O_4225,N_49844,N_49758);
or UO_4226 (O_4226,N_49975,N_49778);
nor UO_4227 (O_4227,N_49969,N_49952);
and UO_4228 (O_4228,N_49921,N_49753);
nand UO_4229 (O_4229,N_49842,N_49848);
xnor UO_4230 (O_4230,N_49808,N_49817);
and UO_4231 (O_4231,N_49945,N_49907);
nor UO_4232 (O_4232,N_49841,N_49948);
xnor UO_4233 (O_4233,N_49823,N_49894);
nand UO_4234 (O_4234,N_49849,N_49795);
nand UO_4235 (O_4235,N_49904,N_49855);
or UO_4236 (O_4236,N_49755,N_49843);
nand UO_4237 (O_4237,N_49889,N_49991);
xor UO_4238 (O_4238,N_49990,N_49768);
xor UO_4239 (O_4239,N_49846,N_49878);
or UO_4240 (O_4240,N_49864,N_49938);
nand UO_4241 (O_4241,N_49769,N_49759);
xor UO_4242 (O_4242,N_49825,N_49759);
or UO_4243 (O_4243,N_49953,N_49821);
nand UO_4244 (O_4244,N_49923,N_49766);
nand UO_4245 (O_4245,N_49931,N_49800);
and UO_4246 (O_4246,N_49939,N_49896);
and UO_4247 (O_4247,N_49927,N_49889);
nand UO_4248 (O_4248,N_49912,N_49908);
and UO_4249 (O_4249,N_49814,N_49756);
xnor UO_4250 (O_4250,N_49897,N_49999);
nand UO_4251 (O_4251,N_49895,N_49869);
and UO_4252 (O_4252,N_49901,N_49818);
or UO_4253 (O_4253,N_49792,N_49799);
xnor UO_4254 (O_4254,N_49895,N_49860);
nor UO_4255 (O_4255,N_49820,N_49882);
nor UO_4256 (O_4256,N_49903,N_49866);
nor UO_4257 (O_4257,N_49975,N_49848);
xor UO_4258 (O_4258,N_49891,N_49977);
nor UO_4259 (O_4259,N_49768,N_49935);
xor UO_4260 (O_4260,N_49874,N_49869);
nand UO_4261 (O_4261,N_49991,N_49770);
xnor UO_4262 (O_4262,N_49782,N_49820);
or UO_4263 (O_4263,N_49880,N_49865);
nor UO_4264 (O_4264,N_49788,N_49861);
and UO_4265 (O_4265,N_49993,N_49980);
nor UO_4266 (O_4266,N_49989,N_49762);
xor UO_4267 (O_4267,N_49813,N_49979);
xnor UO_4268 (O_4268,N_49885,N_49796);
nand UO_4269 (O_4269,N_49820,N_49906);
and UO_4270 (O_4270,N_49965,N_49846);
or UO_4271 (O_4271,N_49816,N_49815);
xor UO_4272 (O_4272,N_49782,N_49837);
or UO_4273 (O_4273,N_49946,N_49874);
nand UO_4274 (O_4274,N_49951,N_49943);
and UO_4275 (O_4275,N_49763,N_49893);
nor UO_4276 (O_4276,N_49817,N_49813);
and UO_4277 (O_4277,N_49869,N_49765);
nand UO_4278 (O_4278,N_49974,N_49807);
or UO_4279 (O_4279,N_49925,N_49760);
or UO_4280 (O_4280,N_49943,N_49972);
nand UO_4281 (O_4281,N_49987,N_49843);
xor UO_4282 (O_4282,N_49888,N_49827);
or UO_4283 (O_4283,N_49823,N_49750);
nand UO_4284 (O_4284,N_49903,N_49799);
nand UO_4285 (O_4285,N_49970,N_49911);
or UO_4286 (O_4286,N_49924,N_49881);
xor UO_4287 (O_4287,N_49765,N_49836);
or UO_4288 (O_4288,N_49822,N_49756);
nor UO_4289 (O_4289,N_49990,N_49832);
nand UO_4290 (O_4290,N_49975,N_49903);
xnor UO_4291 (O_4291,N_49760,N_49942);
xor UO_4292 (O_4292,N_49957,N_49914);
or UO_4293 (O_4293,N_49907,N_49948);
and UO_4294 (O_4294,N_49844,N_49774);
nand UO_4295 (O_4295,N_49853,N_49845);
and UO_4296 (O_4296,N_49874,N_49926);
nor UO_4297 (O_4297,N_49856,N_49877);
xnor UO_4298 (O_4298,N_49950,N_49859);
nand UO_4299 (O_4299,N_49877,N_49948);
nand UO_4300 (O_4300,N_49998,N_49804);
and UO_4301 (O_4301,N_49912,N_49828);
xnor UO_4302 (O_4302,N_49992,N_49904);
or UO_4303 (O_4303,N_49898,N_49992);
nand UO_4304 (O_4304,N_49938,N_49979);
and UO_4305 (O_4305,N_49751,N_49803);
or UO_4306 (O_4306,N_49836,N_49937);
xor UO_4307 (O_4307,N_49948,N_49903);
nor UO_4308 (O_4308,N_49777,N_49962);
or UO_4309 (O_4309,N_49885,N_49750);
and UO_4310 (O_4310,N_49884,N_49848);
xor UO_4311 (O_4311,N_49977,N_49755);
nand UO_4312 (O_4312,N_49901,N_49759);
xnor UO_4313 (O_4313,N_49955,N_49933);
and UO_4314 (O_4314,N_49791,N_49833);
nand UO_4315 (O_4315,N_49873,N_49984);
xnor UO_4316 (O_4316,N_49975,N_49786);
nand UO_4317 (O_4317,N_49816,N_49898);
nand UO_4318 (O_4318,N_49832,N_49878);
xor UO_4319 (O_4319,N_49856,N_49957);
xnor UO_4320 (O_4320,N_49782,N_49819);
or UO_4321 (O_4321,N_49841,N_49974);
or UO_4322 (O_4322,N_49973,N_49919);
nor UO_4323 (O_4323,N_49782,N_49971);
and UO_4324 (O_4324,N_49987,N_49915);
or UO_4325 (O_4325,N_49925,N_49929);
xnor UO_4326 (O_4326,N_49914,N_49946);
nor UO_4327 (O_4327,N_49839,N_49826);
xnor UO_4328 (O_4328,N_49981,N_49917);
and UO_4329 (O_4329,N_49853,N_49929);
nand UO_4330 (O_4330,N_49813,N_49967);
and UO_4331 (O_4331,N_49840,N_49845);
and UO_4332 (O_4332,N_49759,N_49933);
or UO_4333 (O_4333,N_49974,N_49770);
or UO_4334 (O_4334,N_49976,N_49918);
or UO_4335 (O_4335,N_49788,N_49971);
xor UO_4336 (O_4336,N_49842,N_49796);
or UO_4337 (O_4337,N_49885,N_49999);
and UO_4338 (O_4338,N_49839,N_49794);
nor UO_4339 (O_4339,N_49880,N_49942);
nor UO_4340 (O_4340,N_49993,N_49975);
nand UO_4341 (O_4341,N_49750,N_49928);
nor UO_4342 (O_4342,N_49987,N_49963);
or UO_4343 (O_4343,N_49864,N_49966);
nor UO_4344 (O_4344,N_49912,N_49887);
nor UO_4345 (O_4345,N_49786,N_49815);
xnor UO_4346 (O_4346,N_49857,N_49957);
xor UO_4347 (O_4347,N_49987,N_49920);
nor UO_4348 (O_4348,N_49962,N_49938);
nand UO_4349 (O_4349,N_49957,N_49964);
xnor UO_4350 (O_4350,N_49909,N_49982);
nand UO_4351 (O_4351,N_49900,N_49757);
nor UO_4352 (O_4352,N_49894,N_49928);
xor UO_4353 (O_4353,N_49899,N_49787);
nand UO_4354 (O_4354,N_49918,N_49997);
or UO_4355 (O_4355,N_49973,N_49901);
or UO_4356 (O_4356,N_49966,N_49799);
xor UO_4357 (O_4357,N_49833,N_49806);
and UO_4358 (O_4358,N_49969,N_49767);
xnor UO_4359 (O_4359,N_49847,N_49752);
nand UO_4360 (O_4360,N_49977,N_49883);
nand UO_4361 (O_4361,N_49777,N_49981);
and UO_4362 (O_4362,N_49755,N_49968);
nand UO_4363 (O_4363,N_49839,N_49830);
and UO_4364 (O_4364,N_49794,N_49802);
or UO_4365 (O_4365,N_49935,N_49763);
or UO_4366 (O_4366,N_49927,N_49762);
or UO_4367 (O_4367,N_49942,N_49947);
nand UO_4368 (O_4368,N_49934,N_49841);
and UO_4369 (O_4369,N_49993,N_49940);
nor UO_4370 (O_4370,N_49926,N_49988);
and UO_4371 (O_4371,N_49769,N_49959);
xor UO_4372 (O_4372,N_49914,N_49882);
nand UO_4373 (O_4373,N_49768,N_49967);
and UO_4374 (O_4374,N_49780,N_49853);
nand UO_4375 (O_4375,N_49750,N_49930);
xnor UO_4376 (O_4376,N_49903,N_49859);
nand UO_4377 (O_4377,N_49925,N_49867);
or UO_4378 (O_4378,N_49992,N_49983);
nand UO_4379 (O_4379,N_49894,N_49807);
or UO_4380 (O_4380,N_49767,N_49837);
nor UO_4381 (O_4381,N_49926,N_49880);
and UO_4382 (O_4382,N_49913,N_49995);
nor UO_4383 (O_4383,N_49767,N_49829);
nor UO_4384 (O_4384,N_49945,N_49754);
and UO_4385 (O_4385,N_49877,N_49895);
xor UO_4386 (O_4386,N_49818,N_49795);
xor UO_4387 (O_4387,N_49959,N_49997);
and UO_4388 (O_4388,N_49883,N_49819);
nand UO_4389 (O_4389,N_49871,N_49815);
and UO_4390 (O_4390,N_49806,N_49801);
nand UO_4391 (O_4391,N_49847,N_49795);
and UO_4392 (O_4392,N_49843,N_49781);
or UO_4393 (O_4393,N_49904,N_49894);
nand UO_4394 (O_4394,N_49890,N_49776);
nand UO_4395 (O_4395,N_49957,N_49963);
or UO_4396 (O_4396,N_49910,N_49820);
or UO_4397 (O_4397,N_49883,N_49948);
nor UO_4398 (O_4398,N_49815,N_49901);
xnor UO_4399 (O_4399,N_49949,N_49777);
xnor UO_4400 (O_4400,N_49965,N_49956);
nor UO_4401 (O_4401,N_49825,N_49819);
nor UO_4402 (O_4402,N_49865,N_49836);
nor UO_4403 (O_4403,N_49861,N_49977);
xor UO_4404 (O_4404,N_49971,N_49941);
nor UO_4405 (O_4405,N_49867,N_49980);
nand UO_4406 (O_4406,N_49816,N_49904);
and UO_4407 (O_4407,N_49871,N_49818);
or UO_4408 (O_4408,N_49844,N_49920);
nand UO_4409 (O_4409,N_49842,N_49924);
or UO_4410 (O_4410,N_49943,N_49818);
nor UO_4411 (O_4411,N_49961,N_49915);
and UO_4412 (O_4412,N_49811,N_49945);
and UO_4413 (O_4413,N_49762,N_49751);
nor UO_4414 (O_4414,N_49789,N_49975);
nand UO_4415 (O_4415,N_49858,N_49963);
and UO_4416 (O_4416,N_49865,N_49753);
xnor UO_4417 (O_4417,N_49763,N_49990);
and UO_4418 (O_4418,N_49947,N_49854);
nor UO_4419 (O_4419,N_49946,N_49818);
and UO_4420 (O_4420,N_49758,N_49790);
nand UO_4421 (O_4421,N_49957,N_49996);
xnor UO_4422 (O_4422,N_49912,N_49820);
nor UO_4423 (O_4423,N_49964,N_49917);
and UO_4424 (O_4424,N_49829,N_49800);
or UO_4425 (O_4425,N_49940,N_49826);
and UO_4426 (O_4426,N_49936,N_49842);
xnor UO_4427 (O_4427,N_49904,N_49850);
nand UO_4428 (O_4428,N_49916,N_49987);
and UO_4429 (O_4429,N_49983,N_49853);
or UO_4430 (O_4430,N_49944,N_49838);
xor UO_4431 (O_4431,N_49815,N_49971);
or UO_4432 (O_4432,N_49862,N_49958);
nand UO_4433 (O_4433,N_49904,N_49788);
xor UO_4434 (O_4434,N_49856,N_49831);
or UO_4435 (O_4435,N_49885,N_49829);
nor UO_4436 (O_4436,N_49890,N_49956);
nand UO_4437 (O_4437,N_49823,N_49934);
xor UO_4438 (O_4438,N_49853,N_49921);
xnor UO_4439 (O_4439,N_49917,N_49864);
nor UO_4440 (O_4440,N_49807,N_49787);
nor UO_4441 (O_4441,N_49805,N_49869);
xnor UO_4442 (O_4442,N_49891,N_49861);
xor UO_4443 (O_4443,N_49878,N_49837);
nor UO_4444 (O_4444,N_49954,N_49843);
nor UO_4445 (O_4445,N_49922,N_49802);
xnor UO_4446 (O_4446,N_49815,N_49964);
nand UO_4447 (O_4447,N_49818,N_49829);
nor UO_4448 (O_4448,N_49854,N_49905);
nor UO_4449 (O_4449,N_49962,N_49960);
or UO_4450 (O_4450,N_49964,N_49780);
or UO_4451 (O_4451,N_49814,N_49761);
or UO_4452 (O_4452,N_49860,N_49902);
and UO_4453 (O_4453,N_49917,N_49813);
nor UO_4454 (O_4454,N_49811,N_49934);
nand UO_4455 (O_4455,N_49990,N_49937);
xor UO_4456 (O_4456,N_49758,N_49757);
nor UO_4457 (O_4457,N_49822,N_49848);
nor UO_4458 (O_4458,N_49965,N_49885);
or UO_4459 (O_4459,N_49836,N_49844);
nand UO_4460 (O_4460,N_49947,N_49894);
or UO_4461 (O_4461,N_49907,N_49992);
and UO_4462 (O_4462,N_49764,N_49958);
nor UO_4463 (O_4463,N_49792,N_49752);
or UO_4464 (O_4464,N_49993,N_49978);
nor UO_4465 (O_4465,N_49779,N_49774);
nor UO_4466 (O_4466,N_49760,N_49833);
nor UO_4467 (O_4467,N_49845,N_49856);
nand UO_4468 (O_4468,N_49984,N_49877);
or UO_4469 (O_4469,N_49952,N_49944);
and UO_4470 (O_4470,N_49798,N_49939);
and UO_4471 (O_4471,N_49897,N_49929);
and UO_4472 (O_4472,N_49866,N_49937);
nor UO_4473 (O_4473,N_49927,N_49895);
xnor UO_4474 (O_4474,N_49861,N_49914);
nand UO_4475 (O_4475,N_49985,N_49902);
xnor UO_4476 (O_4476,N_49775,N_49829);
nor UO_4477 (O_4477,N_49925,N_49768);
and UO_4478 (O_4478,N_49935,N_49831);
nor UO_4479 (O_4479,N_49846,N_49880);
nand UO_4480 (O_4480,N_49863,N_49857);
nand UO_4481 (O_4481,N_49883,N_49932);
or UO_4482 (O_4482,N_49854,N_49921);
or UO_4483 (O_4483,N_49751,N_49905);
nand UO_4484 (O_4484,N_49825,N_49798);
nand UO_4485 (O_4485,N_49850,N_49913);
nor UO_4486 (O_4486,N_49850,N_49869);
nor UO_4487 (O_4487,N_49956,N_49948);
or UO_4488 (O_4488,N_49951,N_49816);
xnor UO_4489 (O_4489,N_49921,N_49950);
nor UO_4490 (O_4490,N_49882,N_49966);
nand UO_4491 (O_4491,N_49918,N_49931);
or UO_4492 (O_4492,N_49996,N_49892);
xor UO_4493 (O_4493,N_49867,N_49842);
xnor UO_4494 (O_4494,N_49930,N_49852);
xnor UO_4495 (O_4495,N_49765,N_49883);
and UO_4496 (O_4496,N_49785,N_49975);
or UO_4497 (O_4497,N_49786,N_49810);
and UO_4498 (O_4498,N_49989,N_49938);
nand UO_4499 (O_4499,N_49832,N_49966);
nor UO_4500 (O_4500,N_49836,N_49834);
nand UO_4501 (O_4501,N_49786,N_49761);
nor UO_4502 (O_4502,N_49830,N_49758);
nor UO_4503 (O_4503,N_49752,N_49785);
or UO_4504 (O_4504,N_49909,N_49824);
nor UO_4505 (O_4505,N_49830,N_49952);
xnor UO_4506 (O_4506,N_49973,N_49969);
nor UO_4507 (O_4507,N_49902,N_49810);
and UO_4508 (O_4508,N_49893,N_49926);
nor UO_4509 (O_4509,N_49800,N_49930);
or UO_4510 (O_4510,N_49999,N_49822);
nand UO_4511 (O_4511,N_49920,N_49835);
and UO_4512 (O_4512,N_49985,N_49878);
or UO_4513 (O_4513,N_49970,N_49865);
nand UO_4514 (O_4514,N_49760,N_49904);
xor UO_4515 (O_4515,N_49822,N_49926);
or UO_4516 (O_4516,N_49814,N_49842);
nor UO_4517 (O_4517,N_49787,N_49995);
nor UO_4518 (O_4518,N_49790,N_49956);
nand UO_4519 (O_4519,N_49963,N_49873);
xor UO_4520 (O_4520,N_49984,N_49762);
or UO_4521 (O_4521,N_49994,N_49810);
nor UO_4522 (O_4522,N_49759,N_49999);
xnor UO_4523 (O_4523,N_49785,N_49879);
nand UO_4524 (O_4524,N_49813,N_49952);
xnor UO_4525 (O_4525,N_49967,N_49858);
xor UO_4526 (O_4526,N_49775,N_49863);
nor UO_4527 (O_4527,N_49892,N_49848);
and UO_4528 (O_4528,N_49830,N_49930);
and UO_4529 (O_4529,N_49836,N_49882);
nand UO_4530 (O_4530,N_49859,N_49751);
and UO_4531 (O_4531,N_49938,N_49936);
nor UO_4532 (O_4532,N_49838,N_49909);
nor UO_4533 (O_4533,N_49803,N_49930);
or UO_4534 (O_4534,N_49925,N_49767);
nor UO_4535 (O_4535,N_49753,N_49985);
nor UO_4536 (O_4536,N_49929,N_49883);
nand UO_4537 (O_4537,N_49990,N_49800);
nor UO_4538 (O_4538,N_49774,N_49872);
xnor UO_4539 (O_4539,N_49799,N_49902);
nand UO_4540 (O_4540,N_49986,N_49846);
or UO_4541 (O_4541,N_49766,N_49953);
or UO_4542 (O_4542,N_49916,N_49810);
or UO_4543 (O_4543,N_49984,N_49868);
and UO_4544 (O_4544,N_49952,N_49880);
and UO_4545 (O_4545,N_49813,N_49835);
nand UO_4546 (O_4546,N_49864,N_49974);
nand UO_4547 (O_4547,N_49965,N_49939);
and UO_4548 (O_4548,N_49774,N_49835);
xnor UO_4549 (O_4549,N_49761,N_49752);
xor UO_4550 (O_4550,N_49824,N_49792);
xnor UO_4551 (O_4551,N_49834,N_49831);
nor UO_4552 (O_4552,N_49889,N_49840);
xor UO_4553 (O_4553,N_49946,N_49777);
or UO_4554 (O_4554,N_49765,N_49777);
xor UO_4555 (O_4555,N_49804,N_49754);
and UO_4556 (O_4556,N_49930,N_49764);
nor UO_4557 (O_4557,N_49942,N_49965);
xnor UO_4558 (O_4558,N_49878,N_49758);
nor UO_4559 (O_4559,N_49890,N_49860);
and UO_4560 (O_4560,N_49764,N_49977);
xor UO_4561 (O_4561,N_49924,N_49931);
xor UO_4562 (O_4562,N_49876,N_49961);
or UO_4563 (O_4563,N_49995,N_49760);
xor UO_4564 (O_4564,N_49784,N_49856);
or UO_4565 (O_4565,N_49858,N_49789);
nor UO_4566 (O_4566,N_49980,N_49796);
and UO_4567 (O_4567,N_49807,N_49801);
nand UO_4568 (O_4568,N_49757,N_49772);
nand UO_4569 (O_4569,N_49975,N_49856);
or UO_4570 (O_4570,N_49855,N_49925);
xor UO_4571 (O_4571,N_49864,N_49866);
or UO_4572 (O_4572,N_49841,N_49952);
and UO_4573 (O_4573,N_49933,N_49832);
nand UO_4574 (O_4574,N_49758,N_49968);
and UO_4575 (O_4575,N_49925,N_49893);
or UO_4576 (O_4576,N_49865,N_49755);
nor UO_4577 (O_4577,N_49856,N_49918);
nand UO_4578 (O_4578,N_49815,N_49878);
or UO_4579 (O_4579,N_49906,N_49939);
and UO_4580 (O_4580,N_49861,N_49992);
nand UO_4581 (O_4581,N_49798,N_49895);
and UO_4582 (O_4582,N_49967,N_49814);
nand UO_4583 (O_4583,N_49941,N_49822);
xor UO_4584 (O_4584,N_49880,N_49752);
or UO_4585 (O_4585,N_49964,N_49963);
nor UO_4586 (O_4586,N_49842,N_49873);
nor UO_4587 (O_4587,N_49981,N_49852);
or UO_4588 (O_4588,N_49767,N_49809);
and UO_4589 (O_4589,N_49892,N_49946);
xor UO_4590 (O_4590,N_49909,N_49828);
xor UO_4591 (O_4591,N_49937,N_49756);
xnor UO_4592 (O_4592,N_49990,N_49867);
nor UO_4593 (O_4593,N_49819,N_49831);
nand UO_4594 (O_4594,N_49879,N_49927);
or UO_4595 (O_4595,N_49756,N_49986);
or UO_4596 (O_4596,N_49940,N_49925);
xnor UO_4597 (O_4597,N_49954,N_49927);
xor UO_4598 (O_4598,N_49998,N_49999);
xnor UO_4599 (O_4599,N_49963,N_49823);
and UO_4600 (O_4600,N_49849,N_49940);
nand UO_4601 (O_4601,N_49825,N_49793);
or UO_4602 (O_4602,N_49908,N_49831);
or UO_4603 (O_4603,N_49892,N_49860);
nand UO_4604 (O_4604,N_49886,N_49783);
or UO_4605 (O_4605,N_49909,N_49885);
nand UO_4606 (O_4606,N_49977,N_49925);
or UO_4607 (O_4607,N_49950,N_49929);
nor UO_4608 (O_4608,N_49792,N_49769);
or UO_4609 (O_4609,N_49940,N_49833);
xnor UO_4610 (O_4610,N_49774,N_49776);
nor UO_4611 (O_4611,N_49788,N_49833);
xnor UO_4612 (O_4612,N_49853,N_49947);
or UO_4613 (O_4613,N_49875,N_49937);
xnor UO_4614 (O_4614,N_49951,N_49908);
nand UO_4615 (O_4615,N_49947,N_49911);
nor UO_4616 (O_4616,N_49999,N_49896);
nand UO_4617 (O_4617,N_49949,N_49987);
and UO_4618 (O_4618,N_49831,N_49823);
or UO_4619 (O_4619,N_49844,N_49818);
nor UO_4620 (O_4620,N_49853,N_49826);
xnor UO_4621 (O_4621,N_49948,N_49902);
and UO_4622 (O_4622,N_49976,N_49998);
nand UO_4623 (O_4623,N_49812,N_49896);
or UO_4624 (O_4624,N_49805,N_49871);
nor UO_4625 (O_4625,N_49781,N_49890);
xor UO_4626 (O_4626,N_49817,N_49912);
nor UO_4627 (O_4627,N_49858,N_49908);
xnor UO_4628 (O_4628,N_49833,N_49905);
and UO_4629 (O_4629,N_49930,N_49923);
xor UO_4630 (O_4630,N_49971,N_49938);
and UO_4631 (O_4631,N_49916,N_49955);
and UO_4632 (O_4632,N_49779,N_49887);
xnor UO_4633 (O_4633,N_49907,N_49851);
nor UO_4634 (O_4634,N_49780,N_49805);
and UO_4635 (O_4635,N_49947,N_49891);
or UO_4636 (O_4636,N_49815,N_49933);
and UO_4637 (O_4637,N_49962,N_49867);
and UO_4638 (O_4638,N_49798,N_49797);
nor UO_4639 (O_4639,N_49838,N_49996);
nand UO_4640 (O_4640,N_49770,N_49858);
nand UO_4641 (O_4641,N_49917,N_49797);
xor UO_4642 (O_4642,N_49873,N_49795);
nor UO_4643 (O_4643,N_49854,N_49928);
nand UO_4644 (O_4644,N_49814,N_49907);
and UO_4645 (O_4645,N_49930,N_49752);
xor UO_4646 (O_4646,N_49774,N_49801);
xnor UO_4647 (O_4647,N_49880,N_49885);
and UO_4648 (O_4648,N_49881,N_49771);
and UO_4649 (O_4649,N_49878,N_49841);
nor UO_4650 (O_4650,N_49990,N_49814);
xnor UO_4651 (O_4651,N_49783,N_49842);
nand UO_4652 (O_4652,N_49990,N_49934);
nor UO_4653 (O_4653,N_49883,N_49805);
and UO_4654 (O_4654,N_49784,N_49770);
nand UO_4655 (O_4655,N_49935,N_49780);
or UO_4656 (O_4656,N_49758,N_49801);
and UO_4657 (O_4657,N_49900,N_49755);
nor UO_4658 (O_4658,N_49966,N_49976);
xnor UO_4659 (O_4659,N_49763,N_49854);
nand UO_4660 (O_4660,N_49754,N_49948);
or UO_4661 (O_4661,N_49892,N_49994);
or UO_4662 (O_4662,N_49954,N_49949);
nor UO_4663 (O_4663,N_49980,N_49820);
nor UO_4664 (O_4664,N_49783,N_49824);
or UO_4665 (O_4665,N_49839,N_49825);
and UO_4666 (O_4666,N_49792,N_49846);
nor UO_4667 (O_4667,N_49902,N_49859);
nand UO_4668 (O_4668,N_49928,N_49908);
xnor UO_4669 (O_4669,N_49937,N_49926);
or UO_4670 (O_4670,N_49825,N_49900);
or UO_4671 (O_4671,N_49894,N_49933);
xor UO_4672 (O_4672,N_49769,N_49822);
nor UO_4673 (O_4673,N_49881,N_49834);
nand UO_4674 (O_4674,N_49899,N_49910);
nand UO_4675 (O_4675,N_49912,N_49934);
and UO_4676 (O_4676,N_49806,N_49979);
xnor UO_4677 (O_4677,N_49778,N_49987);
nor UO_4678 (O_4678,N_49794,N_49900);
nor UO_4679 (O_4679,N_49782,N_49846);
or UO_4680 (O_4680,N_49832,N_49858);
xnor UO_4681 (O_4681,N_49797,N_49840);
nor UO_4682 (O_4682,N_49980,N_49872);
xnor UO_4683 (O_4683,N_49957,N_49828);
xnor UO_4684 (O_4684,N_49871,N_49788);
nor UO_4685 (O_4685,N_49795,N_49766);
nand UO_4686 (O_4686,N_49861,N_49838);
nor UO_4687 (O_4687,N_49842,N_49816);
and UO_4688 (O_4688,N_49922,N_49889);
xnor UO_4689 (O_4689,N_49968,N_49790);
or UO_4690 (O_4690,N_49857,N_49921);
or UO_4691 (O_4691,N_49919,N_49944);
or UO_4692 (O_4692,N_49862,N_49806);
xnor UO_4693 (O_4693,N_49866,N_49785);
nand UO_4694 (O_4694,N_49969,N_49761);
xor UO_4695 (O_4695,N_49820,N_49916);
nand UO_4696 (O_4696,N_49880,N_49785);
xor UO_4697 (O_4697,N_49945,N_49864);
xor UO_4698 (O_4698,N_49807,N_49876);
or UO_4699 (O_4699,N_49824,N_49918);
and UO_4700 (O_4700,N_49808,N_49766);
or UO_4701 (O_4701,N_49754,N_49903);
or UO_4702 (O_4702,N_49752,N_49921);
xnor UO_4703 (O_4703,N_49768,N_49932);
or UO_4704 (O_4704,N_49970,N_49797);
xor UO_4705 (O_4705,N_49934,N_49794);
or UO_4706 (O_4706,N_49900,N_49866);
xor UO_4707 (O_4707,N_49885,N_49915);
and UO_4708 (O_4708,N_49864,N_49991);
xor UO_4709 (O_4709,N_49979,N_49931);
nand UO_4710 (O_4710,N_49998,N_49993);
xnor UO_4711 (O_4711,N_49924,N_49888);
or UO_4712 (O_4712,N_49856,N_49911);
or UO_4713 (O_4713,N_49972,N_49985);
nor UO_4714 (O_4714,N_49931,N_49959);
xnor UO_4715 (O_4715,N_49868,N_49890);
nor UO_4716 (O_4716,N_49838,N_49763);
nand UO_4717 (O_4717,N_49913,N_49816);
xor UO_4718 (O_4718,N_49786,N_49903);
nor UO_4719 (O_4719,N_49758,N_49859);
and UO_4720 (O_4720,N_49868,N_49787);
xor UO_4721 (O_4721,N_49816,N_49966);
xor UO_4722 (O_4722,N_49983,N_49905);
nor UO_4723 (O_4723,N_49940,N_49847);
or UO_4724 (O_4724,N_49986,N_49839);
xnor UO_4725 (O_4725,N_49801,N_49961);
or UO_4726 (O_4726,N_49794,N_49838);
or UO_4727 (O_4727,N_49850,N_49765);
or UO_4728 (O_4728,N_49984,N_49758);
xnor UO_4729 (O_4729,N_49807,N_49846);
nand UO_4730 (O_4730,N_49894,N_49770);
or UO_4731 (O_4731,N_49857,N_49770);
nand UO_4732 (O_4732,N_49876,N_49755);
nand UO_4733 (O_4733,N_49921,N_49940);
xnor UO_4734 (O_4734,N_49987,N_49884);
nand UO_4735 (O_4735,N_49846,N_49760);
nand UO_4736 (O_4736,N_49936,N_49852);
nand UO_4737 (O_4737,N_49971,N_49840);
xnor UO_4738 (O_4738,N_49931,N_49752);
nand UO_4739 (O_4739,N_49861,N_49835);
xor UO_4740 (O_4740,N_49795,N_49957);
nand UO_4741 (O_4741,N_49856,N_49768);
nor UO_4742 (O_4742,N_49753,N_49939);
or UO_4743 (O_4743,N_49903,N_49999);
or UO_4744 (O_4744,N_49796,N_49783);
nor UO_4745 (O_4745,N_49821,N_49757);
and UO_4746 (O_4746,N_49933,N_49755);
nand UO_4747 (O_4747,N_49916,N_49895);
xor UO_4748 (O_4748,N_49982,N_49786);
and UO_4749 (O_4749,N_49830,N_49874);
nand UO_4750 (O_4750,N_49922,N_49985);
or UO_4751 (O_4751,N_49899,N_49750);
nor UO_4752 (O_4752,N_49959,N_49887);
xor UO_4753 (O_4753,N_49876,N_49984);
xnor UO_4754 (O_4754,N_49805,N_49948);
and UO_4755 (O_4755,N_49980,N_49812);
xor UO_4756 (O_4756,N_49860,N_49786);
nor UO_4757 (O_4757,N_49861,N_49928);
nor UO_4758 (O_4758,N_49848,N_49793);
nand UO_4759 (O_4759,N_49957,N_49761);
nor UO_4760 (O_4760,N_49845,N_49994);
and UO_4761 (O_4761,N_49804,N_49815);
nand UO_4762 (O_4762,N_49773,N_49838);
or UO_4763 (O_4763,N_49974,N_49901);
xor UO_4764 (O_4764,N_49850,N_49845);
nand UO_4765 (O_4765,N_49989,N_49775);
or UO_4766 (O_4766,N_49880,N_49857);
and UO_4767 (O_4767,N_49788,N_49776);
and UO_4768 (O_4768,N_49951,N_49912);
xnor UO_4769 (O_4769,N_49975,N_49830);
or UO_4770 (O_4770,N_49838,N_49898);
and UO_4771 (O_4771,N_49861,N_49937);
xor UO_4772 (O_4772,N_49809,N_49790);
and UO_4773 (O_4773,N_49765,N_49845);
nor UO_4774 (O_4774,N_49798,N_49824);
or UO_4775 (O_4775,N_49860,N_49772);
xor UO_4776 (O_4776,N_49886,N_49819);
nand UO_4777 (O_4777,N_49810,N_49988);
nand UO_4778 (O_4778,N_49925,N_49810);
and UO_4779 (O_4779,N_49835,N_49848);
nor UO_4780 (O_4780,N_49780,N_49909);
nor UO_4781 (O_4781,N_49892,N_49844);
or UO_4782 (O_4782,N_49822,N_49831);
nor UO_4783 (O_4783,N_49971,N_49934);
nor UO_4784 (O_4784,N_49972,N_49825);
or UO_4785 (O_4785,N_49924,N_49956);
xnor UO_4786 (O_4786,N_49962,N_49857);
nor UO_4787 (O_4787,N_49810,N_49774);
nand UO_4788 (O_4788,N_49935,N_49855);
and UO_4789 (O_4789,N_49781,N_49782);
nor UO_4790 (O_4790,N_49906,N_49888);
xor UO_4791 (O_4791,N_49894,N_49879);
or UO_4792 (O_4792,N_49887,N_49791);
or UO_4793 (O_4793,N_49843,N_49922);
nor UO_4794 (O_4794,N_49775,N_49839);
xnor UO_4795 (O_4795,N_49962,N_49762);
and UO_4796 (O_4796,N_49902,N_49927);
and UO_4797 (O_4797,N_49853,N_49785);
xor UO_4798 (O_4798,N_49882,N_49761);
xor UO_4799 (O_4799,N_49882,N_49807);
nand UO_4800 (O_4800,N_49831,N_49835);
nand UO_4801 (O_4801,N_49864,N_49762);
xnor UO_4802 (O_4802,N_49834,N_49971);
or UO_4803 (O_4803,N_49756,N_49903);
or UO_4804 (O_4804,N_49920,N_49917);
and UO_4805 (O_4805,N_49924,N_49855);
nor UO_4806 (O_4806,N_49966,N_49995);
xor UO_4807 (O_4807,N_49892,N_49852);
nand UO_4808 (O_4808,N_49917,N_49970);
xnor UO_4809 (O_4809,N_49969,N_49964);
nand UO_4810 (O_4810,N_49969,N_49835);
nor UO_4811 (O_4811,N_49896,N_49788);
xnor UO_4812 (O_4812,N_49787,N_49844);
and UO_4813 (O_4813,N_49992,N_49912);
nor UO_4814 (O_4814,N_49839,N_49750);
or UO_4815 (O_4815,N_49811,N_49938);
nand UO_4816 (O_4816,N_49759,N_49885);
nand UO_4817 (O_4817,N_49987,N_49831);
nor UO_4818 (O_4818,N_49952,N_49774);
and UO_4819 (O_4819,N_49860,N_49822);
and UO_4820 (O_4820,N_49829,N_49751);
nor UO_4821 (O_4821,N_49819,N_49888);
and UO_4822 (O_4822,N_49995,N_49898);
and UO_4823 (O_4823,N_49995,N_49755);
nor UO_4824 (O_4824,N_49862,N_49793);
xnor UO_4825 (O_4825,N_49870,N_49797);
nor UO_4826 (O_4826,N_49846,N_49757);
or UO_4827 (O_4827,N_49882,N_49815);
and UO_4828 (O_4828,N_49982,N_49938);
or UO_4829 (O_4829,N_49916,N_49879);
nor UO_4830 (O_4830,N_49884,N_49772);
xor UO_4831 (O_4831,N_49910,N_49765);
or UO_4832 (O_4832,N_49819,N_49840);
or UO_4833 (O_4833,N_49914,N_49854);
nand UO_4834 (O_4834,N_49910,N_49924);
xor UO_4835 (O_4835,N_49869,N_49921);
and UO_4836 (O_4836,N_49836,N_49794);
xor UO_4837 (O_4837,N_49832,N_49905);
or UO_4838 (O_4838,N_49952,N_49877);
xnor UO_4839 (O_4839,N_49907,N_49807);
and UO_4840 (O_4840,N_49959,N_49877);
xor UO_4841 (O_4841,N_49767,N_49931);
xor UO_4842 (O_4842,N_49871,N_49797);
nor UO_4843 (O_4843,N_49944,N_49938);
nor UO_4844 (O_4844,N_49779,N_49761);
nand UO_4845 (O_4845,N_49809,N_49982);
and UO_4846 (O_4846,N_49891,N_49787);
nor UO_4847 (O_4847,N_49963,N_49875);
and UO_4848 (O_4848,N_49802,N_49879);
nand UO_4849 (O_4849,N_49921,N_49937);
nor UO_4850 (O_4850,N_49880,N_49751);
and UO_4851 (O_4851,N_49939,N_49785);
xnor UO_4852 (O_4852,N_49845,N_49956);
xor UO_4853 (O_4853,N_49896,N_49863);
nor UO_4854 (O_4854,N_49900,N_49774);
or UO_4855 (O_4855,N_49768,N_49834);
xnor UO_4856 (O_4856,N_49851,N_49898);
xor UO_4857 (O_4857,N_49982,N_49919);
nor UO_4858 (O_4858,N_49967,N_49988);
or UO_4859 (O_4859,N_49838,N_49977);
nor UO_4860 (O_4860,N_49846,N_49852);
or UO_4861 (O_4861,N_49966,N_49813);
nor UO_4862 (O_4862,N_49803,N_49870);
xor UO_4863 (O_4863,N_49799,N_49956);
nand UO_4864 (O_4864,N_49873,N_49760);
nand UO_4865 (O_4865,N_49819,N_49956);
nor UO_4866 (O_4866,N_49830,N_49791);
xor UO_4867 (O_4867,N_49880,N_49906);
and UO_4868 (O_4868,N_49836,N_49822);
and UO_4869 (O_4869,N_49919,N_49963);
nand UO_4870 (O_4870,N_49868,N_49796);
xnor UO_4871 (O_4871,N_49764,N_49966);
or UO_4872 (O_4872,N_49839,N_49808);
or UO_4873 (O_4873,N_49908,N_49925);
nand UO_4874 (O_4874,N_49927,N_49963);
xnor UO_4875 (O_4875,N_49914,N_49851);
nand UO_4876 (O_4876,N_49940,N_49902);
or UO_4877 (O_4877,N_49757,N_49861);
and UO_4878 (O_4878,N_49871,N_49869);
nor UO_4879 (O_4879,N_49958,N_49906);
and UO_4880 (O_4880,N_49833,N_49864);
nand UO_4881 (O_4881,N_49869,N_49968);
xnor UO_4882 (O_4882,N_49967,N_49790);
xor UO_4883 (O_4883,N_49785,N_49979);
nand UO_4884 (O_4884,N_49802,N_49782);
or UO_4885 (O_4885,N_49986,N_49933);
or UO_4886 (O_4886,N_49763,N_49787);
and UO_4887 (O_4887,N_49826,N_49754);
nand UO_4888 (O_4888,N_49976,N_49884);
or UO_4889 (O_4889,N_49932,N_49915);
and UO_4890 (O_4890,N_49875,N_49879);
nor UO_4891 (O_4891,N_49880,N_49943);
and UO_4892 (O_4892,N_49812,N_49752);
xnor UO_4893 (O_4893,N_49762,N_49781);
or UO_4894 (O_4894,N_49886,N_49943);
and UO_4895 (O_4895,N_49966,N_49775);
nand UO_4896 (O_4896,N_49889,N_49770);
and UO_4897 (O_4897,N_49968,N_49853);
nor UO_4898 (O_4898,N_49878,N_49793);
nor UO_4899 (O_4899,N_49874,N_49899);
nor UO_4900 (O_4900,N_49807,N_49987);
xor UO_4901 (O_4901,N_49805,N_49813);
or UO_4902 (O_4902,N_49756,N_49860);
and UO_4903 (O_4903,N_49872,N_49781);
or UO_4904 (O_4904,N_49929,N_49750);
or UO_4905 (O_4905,N_49961,N_49949);
nor UO_4906 (O_4906,N_49969,N_49762);
nand UO_4907 (O_4907,N_49846,N_49802);
xor UO_4908 (O_4908,N_49922,N_49773);
nand UO_4909 (O_4909,N_49933,N_49874);
xor UO_4910 (O_4910,N_49928,N_49977);
or UO_4911 (O_4911,N_49797,N_49813);
or UO_4912 (O_4912,N_49787,N_49904);
or UO_4913 (O_4913,N_49951,N_49810);
nor UO_4914 (O_4914,N_49979,N_49981);
nand UO_4915 (O_4915,N_49924,N_49793);
xnor UO_4916 (O_4916,N_49817,N_49879);
or UO_4917 (O_4917,N_49876,N_49953);
or UO_4918 (O_4918,N_49877,N_49903);
and UO_4919 (O_4919,N_49984,N_49763);
nand UO_4920 (O_4920,N_49891,N_49860);
nand UO_4921 (O_4921,N_49983,N_49815);
nand UO_4922 (O_4922,N_49910,N_49750);
and UO_4923 (O_4923,N_49995,N_49834);
and UO_4924 (O_4924,N_49913,N_49952);
and UO_4925 (O_4925,N_49756,N_49771);
nor UO_4926 (O_4926,N_49937,N_49938);
nand UO_4927 (O_4927,N_49772,N_49818);
nand UO_4928 (O_4928,N_49941,N_49781);
xor UO_4929 (O_4929,N_49981,N_49944);
nand UO_4930 (O_4930,N_49753,N_49954);
and UO_4931 (O_4931,N_49863,N_49790);
nor UO_4932 (O_4932,N_49892,N_49901);
xnor UO_4933 (O_4933,N_49977,N_49955);
and UO_4934 (O_4934,N_49811,N_49833);
nand UO_4935 (O_4935,N_49885,N_49839);
xor UO_4936 (O_4936,N_49811,N_49963);
xor UO_4937 (O_4937,N_49929,N_49804);
nor UO_4938 (O_4938,N_49940,N_49918);
nand UO_4939 (O_4939,N_49991,N_49871);
xnor UO_4940 (O_4940,N_49901,N_49912);
nor UO_4941 (O_4941,N_49869,N_49890);
xnor UO_4942 (O_4942,N_49826,N_49759);
and UO_4943 (O_4943,N_49935,N_49827);
nor UO_4944 (O_4944,N_49790,N_49827);
nand UO_4945 (O_4945,N_49912,N_49978);
and UO_4946 (O_4946,N_49971,N_49909);
nand UO_4947 (O_4947,N_49920,N_49862);
or UO_4948 (O_4948,N_49757,N_49824);
and UO_4949 (O_4949,N_49784,N_49905);
or UO_4950 (O_4950,N_49822,N_49927);
and UO_4951 (O_4951,N_49870,N_49961);
xor UO_4952 (O_4952,N_49799,N_49841);
nor UO_4953 (O_4953,N_49800,N_49946);
nand UO_4954 (O_4954,N_49906,N_49919);
or UO_4955 (O_4955,N_49783,N_49970);
nand UO_4956 (O_4956,N_49858,N_49815);
nand UO_4957 (O_4957,N_49793,N_49786);
nor UO_4958 (O_4958,N_49813,N_49973);
and UO_4959 (O_4959,N_49945,N_49966);
nand UO_4960 (O_4960,N_49867,N_49874);
and UO_4961 (O_4961,N_49972,N_49987);
nor UO_4962 (O_4962,N_49789,N_49897);
nand UO_4963 (O_4963,N_49780,N_49989);
or UO_4964 (O_4964,N_49758,N_49785);
nand UO_4965 (O_4965,N_49990,N_49917);
and UO_4966 (O_4966,N_49994,N_49969);
xnor UO_4967 (O_4967,N_49769,N_49808);
xnor UO_4968 (O_4968,N_49902,N_49794);
nand UO_4969 (O_4969,N_49976,N_49916);
nor UO_4970 (O_4970,N_49833,N_49947);
and UO_4971 (O_4971,N_49917,N_49975);
nor UO_4972 (O_4972,N_49830,N_49769);
nand UO_4973 (O_4973,N_49755,N_49813);
xnor UO_4974 (O_4974,N_49774,N_49803);
nor UO_4975 (O_4975,N_49880,N_49962);
and UO_4976 (O_4976,N_49784,N_49814);
nor UO_4977 (O_4977,N_49828,N_49813);
nand UO_4978 (O_4978,N_49882,N_49904);
and UO_4979 (O_4979,N_49897,N_49890);
nor UO_4980 (O_4980,N_49989,N_49855);
nor UO_4981 (O_4981,N_49810,N_49883);
xor UO_4982 (O_4982,N_49772,N_49854);
or UO_4983 (O_4983,N_49795,N_49858);
nor UO_4984 (O_4984,N_49855,N_49850);
nand UO_4985 (O_4985,N_49921,N_49774);
nand UO_4986 (O_4986,N_49958,N_49814);
and UO_4987 (O_4987,N_49779,N_49795);
xor UO_4988 (O_4988,N_49947,N_49767);
nor UO_4989 (O_4989,N_49804,N_49761);
nand UO_4990 (O_4990,N_49933,N_49900);
and UO_4991 (O_4991,N_49812,N_49820);
and UO_4992 (O_4992,N_49933,N_49877);
or UO_4993 (O_4993,N_49883,N_49983);
nor UO_4994 (O_4994,N_49969,N_49752);
xor UO_4995 (O_4995,N_49983,N_49876);
nor UO_4996 (O_4996,N_49920,N_49959);
xor UO_4997 (O_4997,N_49812,N_49909);
nand UO_4998 (O_4998,N_49895,N_49776);
and UO_4999 (O_4999,N_49755,N_49920);
endmodule