module basic_1000_10000_1500_4_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_684,In_155);
or U1 (N_1,In_305,In_846);
nand U2 (N_2,In_613,In_517);
nor U3 (N_3,In_552,In_304);
and U4 (N_4,In_71,In_405);
nand U5 (N_5,In_972,In_875);
nor U6 (N_6,In_625,In_136);
nand U7 (N_7,In_248,In_599);
xor U8 (N_8,In_825,In_505);
and U9 (N_9,In_96,In_981);
nor U10 (N_10,In_72,In_342);
nor U11 (N_11,In_103,In_420);
nand U12 (N_12,In_432,In_231);
and U13 (N_13,In_462,In_435);
and U14 (N_14,In_757,In_827);
and U15 (N_15,In_196,In_0);
and U16 (N_16,In_53,In_532);
nand U17 (N_17,In_399,In_646);
and U18 (N_18,In_54,In_597);
nand U19 (N_19,In_261,In_851);
or U20 (N_20,In_117,In_689);
or U21 (N_21,In_535,In_915);
or U22 (N_22,In_402,In_42);
nor U23 (N_23,In_102,In_37);
nand U24 (N_24,In_35,In_549);
nand U25 (N_25,In_327,In_956);
nor U26 (N_26,In_13,In_112);
or U27 (N_27,In_667,In_310);
and U28 (N_28,In_282,In_217);
and U29 (N_29,In_735,In_387);
nor U30 (N_30,In_19,In_131);
and U31 (N_31,In_538,In_714);
nor U32 (N_32,In_339,In_108);
and U33 (N_33,In_609,In_640);
nand U34 (N_34,In_760,In_180);
and U35 (N_35,In_897,In_606);
and U36 (N_36,In_911,In_645);
nor U37 (N_37,In_985,In_292);
nor U38 (N_38,In_622,In_750);
nand U39 (N_39,In_464,In_586);
or U40 (N_40,In_783,In_811);
or U41 (N_41,In_543,In_433);
nor U42 (N_42,In_73,In_145);
nand U43 (N_43,In_293,In_78);
nor U44 (N_44,In_234,In_439);
or U45 (N_45,In_480,In_224);
nor U46 (N_46,In_694,In_186);
nand U47 (N_47,In_861,In_977);
and U48 (N_48,In_307,In_813);
and U49 (N_49,In_266,In_545);
nand U50 (N_50,In_283,In_742);
nor U51 (N_51,In_182,In_437);
nor U52 (N_52,In_942,In_643);
nor U53 (N_53,In_928,In_837);
nor U54 (N_54,In_796,In_573);
and U55 (N_55,In_766,In_162);
or U56 (N_56,In_501,In_22);
nor U57 (N_57,In_934,In_470);
nor U58 (N_58,In_756,In_263);
nand U59 (N_59,In_780,In_338);
nand U60 (N_60,In_670,In_719);
nand U61 (N_61,In_577,In_840);
and U62 (N_62,In_101,In_895);
nor U63 (N_63,In_192,In_682);
nor U64 (N_64,In_880,In_82);
nor U65 (N_65,In_690,In_461);
nor U66 (N_66,In_578,In_968);
xnor U67 (N_67,In_489,In_699);
nand U68 (N_68,In_635,In_28);
or U69 (N_69,In_417,In_70);
or U70 (N_70,In_408,In_332);
and U71 (N_71,In_493,In_955);
nand U72 (N_72,In_158,In_236);
xnor U73 (N_73,In_596,In_588);
nor U74 (N_74,In_316,In_375);
and U75 (N_75,In_10,In_716);
or U76 (N_76,In_485,In_127);
nor U77 (N_77,In_152,In_808);
nor U78 (N_78,In_534,In_975);
and U79 (N_79,In_841,In_914);
nand U80 (N_80,In_468,In_215);
and U81 (N_81,In_84,In_451);
or U82 (N_82,In_378,In_59);
or U83 (N_83,In_250,In_376);
or U84 (N_84,In_287,In_881);
nand U85 (N_85,In_513,In_503);
or U86 (N_86,In_963,In_529);
nor U87 (N_87,In_494,In_401);
and U88 (N_88,In_3,In_497);
nand U89 (N_89,In_842,In_495);
xnor U90 (N_90,In_41,In_644);
nand U91 (N_91,In_797,In_321);
nand U92 (N_92,In_326,In_809);
nor U93 (N_93,In_804,In_658);
and U94 (N_94,In_87,In_185);
or U95 (N_95,In_371,In_969);
or U96 (N_96,In_971,In_927);
nor U97 (N_97,In_441,In_739);
nand U98 (N_98,In_33,In_720);
nor U99 (N_99,In_718,In_121);
or U100 (N_100,In_424,In_569);
nand U101 (N_101,In_478,In_729);
and U102 (N_102,In_454,In_329);
nor U103 (N_103,In_567,In_360);
nor U104 (N_104,In_508,In_64);
or U105 (N_105,In_600,In_821);
nand U106 (N_106,In_536,In_228);
nor U107 (N_107,In_492,In_772);
nand U108 (N_108,In_165,In_223);
or U109 (N_109,In_564,In_615);
nor U110 (N_110,In_776,In_657);
and U111 (N_111,In_666,In_982);
nor U112 (N_112,In_257,In_687);
and U113 (N_113,In_479,In_983);
and U114 (N_114,In_651,In_671);
and U115 (N_115,In_738,In_741);
nand U116 (N_116,In_523,In_369);
and U117 (N_117,In_466,In_410);
or U118 (N_118,In_425,In_950);
nand U119 (N_119,In_159,In_562);
nand U120 (N_120,In_949,In_700);
nand U121 (N_121,In_334,In_184);
or U122 (N_122,In_820,In_852);
nor U123 (N_123,In_886,In_873);
nor U124 (N_124,In_979,In_980);
or U125 (N_125,In_672,In_710);
and U126 (N_126,In_740,In_752);
or U127 (N_127,In_572,In_550);
nand U128 (N_128,In_987,In_795);
and U129 (N_129,In_863,In_785);
or U130 (N_130,In_322,In_782);
nor U131 (N_131,In_730,In_372);
and U132 (N_132,In_869,In_436);
and U133 (N_133,In_707,In_362);
and U134 (N_134,In_413,In_918);
or U135 (N_135,In_514,In_260);
or U136 (N_136,In_659,In_724);
nor U137 (N_137,In_252,In_421);
or U138 (N_138,In_1,In_531);
nand U139 (N_139,In_616,In_16);
or U140 (N_140,In_935,In_291);
nor U141 (N_141,In_768,In_770);
nor U142 (N_142,In_188,In_619);
or U143 (N_143,In_359,In_498);
or U144 (N_144,In_389,In_116);
nand U145 (N_145,In_902,In_818);
nor U146 (N_146,In_507,In_591);
nor U147 (N_147,In_636,In_747);
nand U148 (N_148,In_794,In_879);
and U149 (N_149,In_9,In_618);
or U150 (N_150,In_128,In_888);
or U151 (N_151,In_605,In_571);
nand U152 (N_152,In_124,In_105);
and U153 (N_153,In_661,In_132);
xor U154 (N_154,In_452,In_633);
nand U155 (N_155,In_793,In_685);
or U156 (N_156,In_118,In_926);
nand U157 (N_157,In_208,In_426);
or U158 (N_158,In_930,In_801);
or U159 (N_159,In_395,In_213);
and U160 (N_160,In_664,In_522);
nand U161 (N_161,In_153,In_500);
and U162 (N_162,In_107,In_47);
or U163 (N_163,In_922,In_406);
nor U164 (N_164,In_167,In_758);
nor U165 (N_165,In_836,In_692);
nand U166 (N_166,In_126,In_848);
and U167 (N_167,In_348,In_815);
nand U168 (N_168,In_568,In_726);
nor U169 (N_169,In_792,In_330);
or U170 (N_170,In_920,In_674);
nand U171 (N_171,In_995,In_465);
and U172 (N_172,In_237,In_11);
nand U173 (N_173,In_755,In_488);
and U174 (N_174,In_876,In_574);
or U175 (N_175,In_120,In_515);
or U176 (N_176,In_207,In_746);
and U177 (N_177,In_25,In_333);
nor U178 (N_178,In_973,In_702);
or U179 (N_179,In_411,In_253);
nand U180 (N_180,In_916,In_168);
nand U181 (N_181,In_274,In_356);
nor U182 (N_182,In_784,In_473);
nand U183 (N_183,In_303,In_864);
nor U184 (N_184,In_431,In_129);
or U185 (N_185,In_669,In_12);
or U186 (N_186,In_397,In_308);
and U187 (N_187,In_55,In_99);
and U188 (N_188,In_859,In_512);
nor U189 (N_189,In_381,In_113);
and U190 (N_190,In_581,In_403);
and U191 (N_191,In_909,In_510);
or U192 (N_192,In_368,In_100);
and U193 (N_193,In_314,In_798);
nor U194 (N_194,In_824,In_556);
nand U195 (N_195,In_992,In_210);
nand U196 (N_196,In_46,In_176);
and U197 (N_197,In_166,In_88);
nor U198 (N_198,In_891,In_483);
and U199 (N_199,In_731,In_450);
nand U200 (N_200,In_937,In_541);
nor U201 (N_201,In_476,In_986);
or U202 (N_202,In_697,In_265);
nand U203 (N_203,In_874,In_161);
nor U204 (N_204,In_268,In_219);
or U205 (N_205,In_678,In_86);
nand U206 (N_206,In_530,In_151);
nand U207 (N_207,In_90,In_528);
or U208 (N_208,In_504,In_351);
and U209 (N_209,In_839,In_313);
nand U210 (N_210,In_50,In_805);
nand U211 (N_211,In_416,In_892);
and U212 (N_212,In_903,In_831);
or U213 (N_213,In_400,In_249);
nor U214 (N_214,In_233,In_761);
nor U215 (N_215,In_819,In_347);
nand U216 (N_216,In_156,In_775);
nor U217 (N_217,In_172,In_834);
or U218 (N_218,In_952,In_789);
and U219 (N_219,In_448,In_323);
nor U220 (N_220,In_885,In_364);
and U221 (N_221,In_85,In_647);
nor U222 (N_222,In_154,In_23);
and U223 (N_223,In_681,In_21);
nand U224 (N_224,In_900,In_953);
nand U225 (N_225,In_270,In_771);
nor U226 (N_226,In_443,In_810);
and U227 (N_227,In_559,In_883);
nand U228 (N_228,In_79,In_370);
nor U229 (N_229,In_134,In_717);
and U230 (N_230,In_45,In_8);
nor U231 (N_231,In_662,In_743);
nor U232 (N_232,In_26,In_749);
or U233 (N_233,In_214,In_607);
nand U234 (N_234,In_668,In_40);
and U235 (N_235,In_6,In_20);
or U236 (N_236,In_524,In_373);
and U237 (N_237,In_216,In_511);
xor U238 (N_238,In_311,In_936);
nor U239 (N_239,In_943,In_533);
nor U240 (N_240,In_829,In_904);
and U241 (N_241,In_264,In_294);
and U242 (N_242,In_350,In_713);
nand U243 (N_243,In_830,In_601);
nor U244 (N_244,In_227,In_367);
xor U245 (N_245,In_469,In_639);
nand U246 (N_246,In_762,In_390);
nor U247 (N_247,In_773,In_183);
nor U248 (N_248,In_655,In_620);
and U249 (N_249,In_944,In_142);
nor U250 (N_250,In_458,In_247);
and U251 (N_251,In_656,In_898);
or U252 (N_252,In_832,In_141);
nand U253 (N_253,In_769,In_382);
or U254 (N_254,In_737,In_964);
nand U255 (N_255,In_80,In_147);
and U256 (N_256,In_286,In_778);
or U257 (N_257,In_81,In_709);
nand U258 (N_258,In_958,In_175);
and U259 (N_259,In_853,In_477);
and U260 (N_260,In_525,In_868);
nand U261 (N_261,In_967,In_51);
xor U262 (N_262,In_959,In_229);
and U263 (N_263,In_558,In_345);
nor U264 (N_264,In_52,In_608);
and U265 (N_265,In_624,In_4);
or U266 (N_266,In_66,In_537);
and U267 (N_267,In_806,In_276);
nor U268 (N_268,In_945,In_463);
nor U269 (N_269,In_62,In_712);
nor U270 (N_270,In_114,In_634);
or U271 (N_271,In_519,In_910);
and U272 (N_272,In_858,In_164);
or U273 (N_273,In_343,In_324);
nor U274 (N_274,In_843,In_923);
nor U275 (N_275,In_563,In_887);
nand U276 (N_276,In_301,In_48);
or U277 (N_277,In_960,In_56);
and U278 (N_278,In_97,In_77);
nand U279 (N_279,In_384,In_765);
or U280 (N_280,In_92,In_546);
nor U281 (N_281,In_409,In_774);
nor U282 (N_282,In_414,In_976);
nor U283 (N_283,In_866,In_496);
or U284 (N_284,In_457,In_882);
nor U285 (N_285,In_391,In_392);
nand U286 (N_286,In_427,In_627);
or U287 (N_287,In_901,In_111);
or U288 (N_288,In_698,In_27);
nor U289 (N_289,In_732,In_595);
nor U290 (N_290,In_855,In_849);
nor U291 (N_291,In_18,In_246);
nand U292 (N_292,In_238,In_125);
nor U293 (N_293,In_506,In_998);
and U294 (N_294,In_857,In_150);
nor U295 (N_295,In_833,In_239);
nand U296 (N_296,In_455,In_75);
nor U297 (N_297,In_941,In_143);
nor U298 (N_298,In_931,In_68);
nor U299 (N_299,In_225,In_104);
or U300 (N_300,In_315,In_221);
nor U301 (N_301,In_211,In_940);
or U302 (N_302,In_913,In_598);
or U303 (N_303,In_422,In_845);
and U304 (N_304,In_862,In_961);
or U305 (N_305,In_242,In_5);
or U306 (N_306,In_440,In_222);
and U307 (N_307,In_119,In_991);
nand U308 (N_308,In_361,In_996);
nand U309 (N_309,In_244,In_94);
or U310 (N_310,In_814,In_865);
and U311 (N_311,In_575,In_933);
nor U312 (N_312,In_110,In_49);
nor U313 (N_313,In_727,In_412);
nor U314 (N_314,In_553,In_560);
or U315 (N_315,In_585,In_499);
xnor U316 (N_316,In_807,In_653);
and U317 (N_317,In_921,In_281);
nand U318 (N_318,In_331,In_415);
nand U319 (N_319,In_894,In_540);
nor U320 (N_320,In_98,In_146);
or U321 (N_321,In_521,In_896);
and U322 (N_322,In_491,In_123);
and U323 (N_323,In_691,In_61);
and U324 (N_324,In_255,In_95);
nand U325 (N_325,In_803,In_148);
nand U326 (N_326,In_60,In_939);
nor U327 (N_327,In_178,In_14);
nand U328 (N_328,In_790,In_191);
or U329 (N_329,In_63,In_877);
and U330 (N_330,In_200,In_786);
nand U331 (N_331,In_802,In_352);
and U332 (N_332,In_544,In_272);
nand U333 (N_333,In_917,In_978);
nand U334 (N_334,In_15,In_611);
and U335 (N_335,In_31,In_366);
and U336 (N_336,In_576,In_140);
nand U337 (N_337,In_204,In_763);
nor U338 (N_338,In_988,In_144);
nor U339 (N_339,In_999,In_340);
or U340 (N_340,In_854,In_642);
and U341 (N_341,In_44,In_520);
nor U342 (N_342,In_115,In_76);
or U343 (N_343,In_357,In_823);
or U344 (N_344,In_688,In_472);
nor U345 (N_345,In_349,In_650);
nand U346 (N_346,In_663,In_665);
nand U347 (N_347,In_856,In_335);
and U348 (N_348,In_446,In_679);
and U349 (N_349,In_174,In_481);
nor U350 (N_350,In_285,In_309);
nand U351 (N_351,In_482,In_889);
nor U352 (N_352,In_404,In_602);
and U353 (N_353,In_474,In_383);
or U354 (N_354,In_754,In_302);
and U355 (N_355,In_518,In_566);
nand U356 (N_356,In_194,In_871);
and U357 (N_357,In_83,In_201);
nand U358 (N_358,In_948,In_966);
nand U359 (N_359,In_69,In_377);
and U360 (N_360,In_442,In_965);
and U361 (N_361,In_838,In_394);
and U362 (N_362,In_187,In_212);
and U363 (N_363,In_38,In_905);
nand U364 (N_364,In_583,In_318);
nand U365 (N_365,In_723,In_767);
and U366 (N_366,In_954,In_130);
nand U367 (N_367,In_759,In_899);
or U368 (N_368,In_587,In_438);
nor U369 (N_369,In_693,In_705);
nor U370 (N_370,In_295,In_277);
and U371 (N_371,In_908,In_336);
nor U372 (N_372,In_34,In_736);
or U373 (N_373,In_812,In_610);
nor U374 (N_374,In_641,In_133);
and U375 (N_375,In_946,In_365);
or U376 (N_376,In_721,In_555);
nor U377 (N_377,In_346,In_695);
or U378 (N_378,In_704,In_328);
nor U379 (N_379,In_363,In_547);
nor U380 (N_380,In_938,In_460);
nor U381 (N_381,In_502,In_241);
and U382 (N_382,In_893,In_288);
and U383 (N_383,In_195,In_870);
nor U384 (N_384,In_993,In_445);
nand U385 (N_385,In_299,In_170);
or U386 (N_386,In_631,In_379);
nand U387 (N_387,In_486,In_557);
and U388 (N_388,In_269,In_284);
nand U389 (N_389,In_554,In_579);
nand U390 (N_390,In_660,In_683);
nand U391 (N_391,In_181,In_58);
or U392 (N_392,In_256,In_997);
nor U393 (N_393,In_594,In_230);
or U394 (N_394,In_358,In_262);
or U395 (N_395,In_300,In_487);
or U396 (N_396,In_527,In_816);
or U397 (N_397,In_844,In_734);
or U398 (N_398,In_177,In_418);
and U399 (N_399,In_733,In_199);
or U400 (N_400,In_787,In_703);
nor U401 (N_401,In_551,In_509);
or U402 (N_402,In_149,In_711);
nand U403 (N_403,In_490,In_206);
and U404 (N_404,In_706,In_380);
and U405 (N_405,In_565,In_628);
and U406 (N_406,In_254,In_344);
or U407 (N_407,In_925,In_580);
and U408 (N_408,In_205,In_139);
nor U409 (N_409,In_632,In_799);
xnor U410 (N_410,In_725,In_43);
nor U411 (N_411,In_385,In_279);
nor U412 (N_412,In_36,In_516);
or U413 (N_413,In_561,In_275);
and U414 (N_414,In_648,In_273);
nor U415 (N_415,In_271,In_974);
nand U416 (N_416,In_267,In_290);
nor U417 (N_417,In_924,In_817);
nor U418 (N_418,In_722,In_198);
nor U419 (N_419,In_542,In_163);
and U420 (N_420,In_297,In_449);
or U421 (N_421,In_89,In_612);
nor U422 (N_422,In_748,In_957);
nand U423 (N_423,In_919,In_453);
nor U424 (N_424,In_444,In_189);
nor U425 (N_425,In_777,In_428);
or U426 (N_426,In_278,In_24);
or U427 (N_427,In_744,In_745);
nor U428 (N_428,In_289,In_57);
nand U429 (N_429,In_169,In_29);
and U430 (N_430,In_878,In_374);
nor U431 (N_431,In_584,In_475);
and U432 (N_432,In_419,In_109);
nand U433 (N_433,In_429,In_341);
or U434 (N_434,In_614,In_243);
or U435 (N_435,In_280,In_764);
nor U436 (N_436,In_298,In_354);
nand U437 (N_437,In_386,In_912);
and U438 (N_438,In_74,In_686);
and U439 (N_439,In_994,In_800);
or U440 (N_440,In_867,In_355);
nor U441 (N_441,In_788,In_654);
nand U442 (N_442,In_708,In_202);
and U443 (N_443,In_637,In_160);
nor U444 (N_444,In_629,In_638);
nor U445 (N_445,In_226,In_122);
nand U446 (N_446,In_220,In_30);
nand U447 (N_447,In_434,In_791);
and U448 (N_448,In_592,In_106);
nor U449 (N_449,In_135,In_259);
and U450 (N_450,In_623,In_984);
or U451 (N_451,In_312,In_467);
nor U452 (N_452,In_539,In_296);
nand U453 (N_453,In_456,In_396);
and U454 (N_454,In_320,In_582);
nor U455 (N_455,In_822,In_884);
nor U456 (N_456,In_317,In_39);
and U457 (N_457,In_626,In_929);
and U458 (N_458,In_337,In_388);
nor U459 (N_459,In_835,In_590);
or U460 (N_460,In_32,In_675);
and U461 (N_461,In_753,In_676);
or U462 (N_462,In_93,In_728);
nor U463 (N_463,In_593,In_138);
nor U464 (N_464,In_232,In_951);
nand U465 (N_465,In_393,In_677);
and U466 (N_466,In_319,In_906);
or U467 (N_467,In_423,In_484);
nand U468 (N_468,In_91,In_828);
xnor U469 (N_469,In_17,In_589);
nand U470 (N_470,In_447,In_715);
nor U471 (N_471,In_471,In_932);
or U472 (N_472,In_652,In_240);
nand U473 (N_473,In_989,In_137);
or U474 (N_474,In_398,In_850);
nor U475 (N_475,In_65,In_604);
nand U476 (N_476,In_751,In_907);
or U477 (N_477,In_258,In_990);
nor U478 (N_478,In_570,In_325);
nor U479 (N_479,In_67,In_179);
or U480 (N_480,In_617,In_459);
nor U481 (N_481,In_306,In_630);
or U482 (N_482,In_251,In_171);
nor U483 (N_483,In_872,In_701);
nor U484 (N_484,In_218,In_649);
or U485 (N_485,In_353,In_847);
nor U486 (N_486,In_603,In_890);
nand U487 (N_487,In_2,In_947);
nand U488 (N_488,In_962,In_245);
nand U489 (N_489,In_209,In_7);
nand U490 (N_490,In_193,In_970);
and U491 (N_491,In_779,In_430);
or U492 (N_492,In_173,In_526);
or U493 (N_493,In_407,In_673);
and U494 (N_494,In_621,In_781);
nand U495 (N_495,In_826,In_860);
or U496 (N_496,In_548,In_696);
nor U497 (N_497,In_157,In_203);
nor U498 (N_498,In_680,In_190);
nand U499 (N_499,In_235,In_197);
or U500 (N_500,In_920,In_230);
or U501 (N_501,In_112,In_172);
or U502 (N_502,In_152,In_718);
or U503 (N_503,In_139,In_844);
nand U504 (N_504,In_760,In_251);
and U505 (N_505,In_553,In_716);
nor U506 (N_506,In_496,In_3);
nor U507 (N_507,In_271,In_138);
and U508 (N_508,In_495,In_574);
nor U509 (N_509,In_704,In_931);
nor U510 (N_510,In_466,In_419);
nand U511 (N_511,In_394,In_552);
nor U512 (N_512,In_872,In_227);
nor U513 (N_513,In_492,In_580);
nor U514 (N_514,In_565,In_932);
or U515 (N_515,In_217,In_658);
and U516 (N_516,In_656,In_513);
nand U517 (N_517,In_763,In_861);
nand U518 (N_518,In_347,In_390);
and U519 (N_519,In_680,In_831);
and U520 (N_520,In_156,In_753);
and U521 (N_521,In_247,In_262);
nand U522 (N_522,In_870,In_868);
nor U523 (N_523,In_263,In_396);
or U524 (N_524,In_893,In_550);
nor U525 (N_525,In_495,In_751);
nor U526 (N_526,In_638,In_82);
nor U527 (N_527,In_381,In_475);
or U528 (N_528,In_535,In_965);
nor U529 (N_529,In_72,In_999);
or U530 (N_530,In_825,In_746);
nand U531 (N_531,In_805,In_98);
nand U532 (N_532,In_765,In_87);
or U533 (N_533,In_178,In_590);
or U534 (N_534,In_604,In_950);
nor U535 (N_535,In_365,In_827);
nor U536 (N_536,In_313,In_55);
and U537 (N_537,In_763,In_534);
and U538 (N_538,In_37,In_717);
nor U539 (N_539,In_173,In_187);
nand U540 (N_540,In_757,In_947);
and U541 (N_541,In_391,In_354);
or U542 (N_542,In_337,In_888);
or U543 (N_543,In_978,In_381);
nor U544 (N_544,In_524,In_864);
and U545 (N_545,In_918,In_470);
nor U546 (N_546,In_818,In_178);
nor U547 (N_547,In_656,In_179);
nor U548 (N_548,In_700,In_722);
and U549 (N_549,In_616,In_851);
nor U550 (N_550,In_679,In_803);
nand U551 (N_551,In_823,In_279);
and U552 (N_552,In_584,In_954);
or U553 (N_553,In_689,In_299);
nor U554 (N_554,In_603,In_107);
nor U555 (N_555,In_807,In_540);
nand U556 (N_556,In_128,In_155);
and U557 (N_557,In_646,In_120);
nor U558 (N_558,In_900,In_686);
nand U559 (N_559,In_201,In_750);
or U560 (N_560,In_486,In_226);
or U561 (N_561,In_140,In_209);
nand U562 (N_562,In_184,In_569);
and U563 (N_563,In_419,In_385);
and U564 (N_564,In_368,In_475);
nand U565 (N_565,In_496,In_822);
and U566 (N_566,In_306,In_185);
nor U567 (N_567,In_30,In_66);
or U568 (N_568,In_47,In_984);
or U569 (N_569,In_242,In_226);
or U570 (N_570,In_33,In_887);
or U571 (N_571,In_592,In_89);
or U572 (N_572,In_88,In_635);
and U573 (N_573,In_811,In_414);
and U574 (N_574,In_836,In_929);
or U575 (N_575,In_46,In_181);
nand U576 (N_576,In_3,In_22);
and U577 (N_577,In_906,In_357);
or U578 (N_578,In_292,In_872);
and U579 (N_579,In_942,In_403);
or U580 (N_580,In_538,In_444);
xor U581 (N_581,In_956,In_655);
nor U582 (N_582,In_879,In_149);
nand U583 (N_583,In_291,In_919);
and U584 (N_584,In_320,In_74);
or U585 (N_585,In_697,In_94);
and U586 (N_586,In_892,In_262);
or U587 (N_587,In_542,In_99);
or U588 (N_588,In_613,In_381);
or U589 (N_589,In_453,In_377);
nor U590 (N_590,In_857,In_962);
nor U591 (N_591,In_868,In_42);
nand U592 (N_592,In_695,In_826);
or U593 (N_593,In_333,In_232);
nand U594 (N_594,In_84,In_832);
nand U595 (N_595,In_706,In_46);
or U596 (N_596,In_693,In_109);
and U597 (N_597,In_496,In_754);
nor U598 (N_598,In_350,In_139);
and U599 (N_599,In_208,In_214);
and U600 (N_600,In_624,In_354);
nor U601 (N_601,In_202,In_517);
nor U602 (N_602,In_741,In_43);
nor U603 (N_603,In_798,In_112);
nor U604 (N_604,In_156,In_446);
and U605 (N_605,In_664,In_99);
nor U606 (N_606,In_701,In_529);
or U607 (N_607,In_284,In_739);
or U608 (N_608,In_270,In_645);
and U609 (N_609,In_81,In_724);
and U610 (N_610,In_882,In_959);
xnor U611 (N_611,In_669,In_493);
and U612 (N_612,In_959,In_244);
and U613 (N_613,In_959,In_964);
and U614 (N_614,In_470,In_600);
nand U615 (N_615,In_120,In_482);
nor U616 (N_616,In_246,In_840);
or U617 (N_617,In_602,In_946);
nand U618 (N_618,In_72,In_432);
nand U619 (N_619,In_310,In_460);
and U620 (N_620,In_623,In_368);
and U621 (N_621,In_488,In_920);
nand U622 (N_622,In_653,In_414);
nand U623 (N_623,In_148,In_688);
or U624 (N_624,In_127,In_246);
or U625 (N_625,In_722,In_783);
nor U626 (N_626,In_134,In_31);
and U627 (N_627,In_656,In_168);
and U628 (N_628,In_871,In_643);
nand U629 (N_629,In_201,In_525);
and U630 (N_630,In_236,In_547);
or U631 (N_631,In_802,In_460);
nor U632 (N_632,In_845,In_975);
nor U633 (N_633,In_879,In_359);
or U634 (N_634,In_639,In_717);
and U635 (N_635,In_477,In_335);
or U636 (N_636,In_742,In_853);
and U637 (N_637,In_541,In_387);
nor U638 (N_638,In_932,In_26);
nor U639 (N_639,In_166,In_208);
nor U640 (N_640,In_592,In_223);
nor U641 (N_641,In_579,In_442);
nand U642 (N_642,In_678,In_403);
nand U643 (N_643,In_327,In_510);
and U644 (N_644,In_138,In_865);
or U645 (N_645,In_216,In_35);
and U646 (N_646,In_432,In_525);
and U647 (N_647,In_865,In_583);
or U648 (N_648,In_314,In_375);
or U649 (N_649,In_600,In_603);
xor U650 (N_650,In_267,In_559);
nor U651 (N_651,In_153,In_338);
nor U652 (N_652,In_854,In_543);
nor U653 (N_653,In_735,In_711);
nor U654 (N_654,In_820,In_41);
and U655 (N_655,In_556,In_761);
nor U656 (N_656,In_920,In_524);
nor U657 (N_657,In_39,In_935);
and U658 (N_658,In_395,In_134);
and U659 (N_659,In_674,In_566);
nor U660 (N_660,In_304,In_243);
nand U661 (N_661,In_577,In_9);
nand U662 (N_662,In_307,In_38);
and U663 (N_663,In_436,In_924);
nor U664 (N_664,In_25,In_484);
nor U665 (N_665,In_365,In_158);
nor U666 (N_666,In_284,In_700);
and U667 (N_667,In_459,In_904);
nor U668 (N_668,In_851,In_333);
nand U669 (N_669,In_815,In_166);
nor U670 (N_670,In_936,In_379);
nor U671 (N_671,In_494,In_107);
nor U672 (N_672,In_24,In_413);
nand U673 (N_673,In_699,In_336);
and U674 (N_674,In_499,In_688);
nor U675 (N_675,In_809,In_522);
nand U676 (N_676,In_206,In_542);
or U677 (N_677,In_830,In_424);
and U678 (N_678,In_43,In_723);
or U679 (N_679,In_597,In_373);
nand U680 (N_680,In_617,In_487);
or U681 (N_681,In_71,In_386);
nor U682 (N_682,In_85,In_880);
and U683 (N_683,In_972,In_726);
nand U684 (N_684,In_254,In_704);
nor U685 (N_685,In_619,In_856);
or U686 (N_686,In_285,In_925);
and U687 (N_687,In_287,In_188);
and U688 (N_688,In_107,In_652);
nor U689 (N_689,In_748,In_687);
and U690 (N_690,In_766,In_836);
and U691 (N_691,In_408,In_213);
nand U692 (N_692,In_60,In_712);
nand U693 (N_693,In_433,In_798);
xor U694 (N_694,In_73,In_33);
nor U695 (N_695,In_186,In_280);
or U696 (N_696,In_870,In_767);
or U697 (N_697,In_743,In_723);
nand U698 (N_698,In_304,In_241);
and U699 (N_699,In_89,In_562);
and U700 (N_700,In_215,In_221);
nor U701 (N_701,In_326,In_580);
and U702 (N_702,In_591,In_844);
nor U703 (N_703,In_565,In_901);
xnor U704 (N_704,In_701,In_991);
nand U705 (N_705,In_16,In_300);
or U706 (N_706,In_790,In_31);
nor U707 (N_707,In_607,In_436);
and U708 (N_708,In_937,In_365);
or U709 (N_709,In_883,In_64);
nand U710 (N_710,In_581,In_923);
or U711 (N_711,In_368,In_442);
nand U712 (N_712,In_519,In_171);
or U713 (N_713,In_818,In_600);
nand U714 (N_714,In_64,In_882);
or U715 (N_715,In_730,In_139);
and U716 (N_716,In_885,In_625);
or U717 (N_717,In_681,In_801);
nor U718 (N_718,In_954,In_454);
nor U719 (N_719,In_187,In_885);
nand U720 (N_720,In_491,In_360);
and U721 (N_721,In_322,In_158);
and U722 (N_722,In_105,In_457);
or U723 (N_723,In_194,In_809);
and U724 (N_724,In_575,In_825);
nor U725 (N_725,In_25,In_753);
and U726 (N_726,In_994,In_918);
nand U727 (N_727,In_417,In_396);
or U728 (N_728,In_687,In_222);
nand U729 (N_729,In_90,In_573);
or U730 (N_730,In_804,In_404);
nand U731 (N_731,In_305,In_547);
nand U732 (N_732,In_983,In_823);
or U733 (N_733,In_225,In_443);
or U734 (N_734,In_569,In_880);
and U735 (N_735,In_417,In_79);
nor U736 (N_736,In_383,In_8);
or U737 (N_737,In_546,In_789);
nor U738 (N_738,In_129,In_621);
or U739 (N_739,In_511,In_444);
nor U740 (N_740,In_297,In_204);
nand U741 (N_741,In_420,In_243);
nor U742 (N_742,In_41,In_870);
nor U743 (N_743,In_141,In_835);
and U744 (N_744,In_907,In_701);
and U745 (N_745,In_809,In_11);
nand U746 (N_746,In_311,In_874);
nor U747 (N_747,In_3,In_686);
and U748 (N_748,In_579,In_529);
nand U749 (N_749,In_713,In_214);
or U750 (N_750,In_151,In_319);
nand U751 (N_751,In_330,In_661);
nand U752 (N_752,In_896,In_398);
and U753 (N_753,In_691,In_696);
nand U754 (N_754,In_515,In_403);
or U755 (N_755,In_56,In_419);
or U756 (N_756,In_482,In_714);
and U757 (N_757,In_883,In_417);
or U758 (N_758,In_732,In_199);
or U759 (N_759,In_589,In_376);
nand U760 (N_760,In_153,In_620);
or U761 (N_761,In_60,In_448);
or U762 (N_762,In_163,In_624);
and U763 (N_763,In_413,In_158);
and U764 (N_764,In_370,In_592);
nand U765 (N_765,In_866,In_865);
nand U766 (N_766,In_450,In_323);
or U767 (N_767,In_398,In_448);
nand U768 (N_768,In_982,In_425);
nor U769 (N_769,In_954,In_369);
and U770 (N_770,In_973,In_7);
and U771 (N_771,In_780,In_467);
and U772 (N_772,In_338,In_790);
nand U773 (N_773,In_931,In_5);
nand U774 (N_774,In_117,In_281);
and U775 (N_775,In_69,In_556);
and U776 (N_776,In_793,In_357);
nand U777 (N_777,In_185,In_736);
or U778 (N_778,In_363,In_830);
nand U779 (N_779,In_857,In_177);
nor U780 (N_780,In_845,In_138);
or U781 (N_781,In_875,In_691);
nor U782 (N_782,In_275,In_246);
and U783 (N_783,In_329,In_833);
and U784 (N_784,In_532,In_101);
nor U785 (N_785,In_423,In_866);
and U786 (N_786,In_945,In_104);
nor U787 (N_787,In_998,In_661);
or U788 (N_788,In_870,In_375);
and U789 (N_789,In_911,In_348);
nor U790 (N_790,In_725,In_518);
and U791 (N_791,In_124,In_217);
and U792 (N_792,In_379,In_34);
nor U793 (N_793,In_961,In_44);
or U794 (N_794,In_790,In_468);
or U795 (N_795,In_349,In_716);
and U796 (N_796,In_781,In_702);
nand U797 (N_797,In_840,In_644);
and U798 (N_798,In_564,In_705);
and U799 (N_799,In_606,In_283);
nor U800 (N_800,In_949,In_932);
or U801 (N_801,In_355,In_921);
and U802 (N_802,In_862,In_840);
and U803 (N_803,In_197,In_548);
xor U804 (N_804,In_402,In_220);
or U805 (N_805,In_198,In_205);
nand U806 (N_806,In_620,In_832);
or U807 (N_807,In_291,In_485);
nand U808 (N_808,In_959,In_785);
nand U809 (N_809,In_702,In_461);
nor U810 (N_810,In_469,In_981);
and U811 (N_811,In_273,In_899);
and U812 (N_812,In_512,In_793);
and U813 (N_813,In_978,In_132);
nor U814 (N_814,In_373,In_761);
and U815 (N_815,In_307,In_370);
nand U816 (N_816,In_513,In_285);
nor U817 (N_817,In_757,In_733);
nor U818 (N_818,In_843,In_359);
nand U819 (N_819,In_924,In_651);
or U820 (N_820,In_733,In_365);
nand U821 (N_821,In_363,In_9);
or U822 (N_822,In_218,In_604);
nand U823 (N_823,In_48,In_266);
and U824 (N_824,In_796,In_448);
or U825 (N_825,In_149,In_582);
nand U826 (N_826,In_396,In_168);
or U827 (N_827,In_459,In_513);
nand U828 (N_828,In_765,In_899);
nor U829 (N_829,In_781,In_821);
and U830 (N_830,In_329,In_792);
nand U831 (N_831,In_322,In_905);
nand U832 (N_832,In_304,In_687);
nor U833 (N_833,In_756,In_709);
or U834 (N_834,In_668,In_965);
nand U835 (N_835,In_489,In_563);
nand U836 (N_836,In_409,In_753);
or U837 (N_837,In_378,In_372);
nand U838 (N_838,In_646,In_31);
and U839 (N_839,In_582,In_228);
and U840 (N_840,In_558,In_949);
and U841 (N_841,In_263,In_971);
nand U842 (N_842,In_252,In_556);
or U843 (N_843,In_840,In_121);
and U844 (N_844,In_862,In_190);
and U845 (N_845,In_504,In_249);
or U846 (N_846,In_991,In_771);
nor U847 (N_847,In_892,In_567);
or U848 (N_848,In_177,In_927);
or U849 (N_849,In_850,In_702);
and U850 (N_850,In_288,In_198);
or U851 (N_851,In_175,In_826);
and U852 (N_852,In_887,In_324);
or U853 (N_853,In_128,In_118);
or U854 (N_854,In_283,In_879);
or U855 (N_855,In_523,In_181);
or U856 (N_856,In_271,In_217);
and U857 (N_857,In_235,In_374);
nand U858 (N_858,In_995,In_211);
nor U859 (N_859,In_243,In_88);
nor U860 (N_860,In_980,In_673);
nand U861 (N_861,In_626,In_687);
or U862 (N_862,In_576,In_740);
nor U863 (N_863,In_90,In_956);
and U864 (N_864,In_452,In_512);
and U865 (N_865,In_656,In_223);
or U866 (N_866,In_395,In_899);
or U867 (N_867,In_352,In_809);
or U868 (N_868,In_683,In_405);
nor U869 (N_869,In_50,In_74);
or U870 (N_870,In_258,In_291);
nand U871 (N_871,In_972,In_85);
or U872 (N_872,In_777,In_734);
and U873 (N_873,In_676,In_485);
or U874 (N_874,In_921,In_85);
nand U875 (N_875,In_170,In_639);
or U876 (N_876,In_920,In_139);
or U877 (N_877,In_899,In_942);
or U878 (N_878,In_803,In_381);
xor U879 (N_879,In_208,In_742);
nand U880 (N_880,In_356,In_156);
nand U881 (N_881,In_461,In_745);
or U882 (N_882,In_878,In_238);
nand U883 (N_883,In_610,In_666);
nand U884 (N_884,In_42,In_810);
nand U885 (N_885,In_647,In_2);
nor U886 (N_886,In_368,In_160);
and U887 (N_887,In_399,In_850);
nand U888 (N_888,In_595,In_110);
nor U889 (N_889,In_584,In_104);
or U890 (N_890,In_677,In_292);
nor U891 (N_891,In_880,In_20);
and U892 (N_892,In_386,In_703);
nand U893 (N_893,In_804,In_591);
nand U894 (N_894,In_194,In_384);
and U895 (N_895,In_472,In_992);
nand U896 (N_896,In_779,In_151);
nand U897 (N_897,In_351,In_841);
nand U898 (N_898,In_721,In_731);
and U899 (N_899,In_123,In_808);
nor U900 (N_900,In_864,In_439);
or U901 (N_901,In_62,In_275);
nor U902 (N_902,In_209,In_143);
or U903 (N_903,In_277,In_951);
and U904 (N_904,In_782,In_209);
nand U905 (N_905,In_87,In_96);
or U906 (N_906,In_44,In_384);
nor U907 (N_907,In_687,In_616);
xnor U908 (N_908,In_934,In_737);
or U909 (N_909,In_507,In_417);
or U910 (N_910,In_560,In_499);
and U911 (N_911,In_120,In_423);
nor U912 (N_912,In_454,In_749);
nand U913 (N_913,In_237,In_639);
and U914 (N_914,In_73,In_467);
nor U915 (N_915,In_604,In_405);
or U916 (N_916,In_701,In_895);
or U917 (N_917,In_171,In_303);
or U918 (N_918,In_664,In_847);
and U919 (N_919,In_310,In_615);
and U920 (N_920,In_459,In_54);
or U921 (N_921,In_698,In_298);
nor U922 (N_922,In_460,In_724);
or U923 (N_923,In_330,In_120);
and U924 (N_924,In_360,In_49);
or U925 (N_925,In_413,In_998);
and U926 (N_926,In_289,In_240);
or U927 (N_927,In_32,In_549);
nand U928 (N_928,In_828,In_956);
and U929 (N_929,In_447,In_125);
nor U930 (N_930,In_378,In_664);
and U931 (N_931,In_594,In_573);
nor U932 (N_932,In_796,In_210);
and U933 (N_933,In_176,In_113);
nor U934 (N_934,In_173,In_430);
and U935 (N_935,In_892,In_380);
and U936 (N_936,In_524,In_945);
and U937 (N_937,In_939,In_3);
or U938 (N_938,In_347,In_285);
and U939 (N_939,In_195,In_784);
nor U940 (N_940,In_128,In_460);
nor U941 (N_941,In_702,In_222);
nor U942 (N_942,In_288,In_214);
nor U943 (N_943,In_421,In_730);
and U944 (N_944,In_805,In_262);
nor U945 (N_945,In_511,In_946);
nand U946 (N_946,In_173,In_938);
or U947 (N_947,In_585,In_435);
nor U948 (N_948,In_107,In_808);
or U949 (N_949,In_179,In_139);
or U950 (N_950,In_581,In_347);
and U951 (N_951,In_646,In_737);
and U952 (N_952,In_59,In_451);
and U953 (N_953,In_853,In_442);
or U954 (N_954,In_960,In_910);
nor U955 (N_955,In_666,In_343);
or U956 (N_956,In_312,In_739);
and U957 (N_957,In_602,In_221);
nor U958 (N_958,In_903,In_59);
or U959 (N_959,In_831,In_407);
nand U960 (N_960,In_715,In_782);
or U961 (N_961,In_362,In_69);
nand U962 (N_962,In_93,In_432);
nand U963 (N_963,In_339,In_311);
nand U964 (N_964,In_548,In_202);
nor U965 (N_965,In_173,In_212);
or U966 (N_966,In_202,In_296);
or U967 (N_967,In_715,In_63);
or U968 (N_968,In_469,In_495);
nand U969 (N_969,In_264,In_578);
nor U970 (N_970,In_629,In_174);
and U971 (N_971,In_140,In_417);
or U972 (N_972,In_771,In_501);
and U973 (N_973,In_123,In_355);
nand U974 (N_974,In_233,In_228);
or U975 (N_975,In_909,In_810);
or U976 (N_976,In_733,In_586);
nand U977 (N_977,In_867,In_802);
nor U978 (N_978,In_188,In_879);
nor U979 (N_979,In_493,In_492);
and U980 (N_980,In_266,In_619);
nand U981 (N_981,In_703,In_12);
or U982 (N_982,In_764,In_225);
and U983 (N_983,In_899,In_601);
or U984 (N_984,In_427,In_951);
or U985 (N_985,In_284,In_970);
nor U986 (N_986,In_686,In_744);
or U987 (N_987,In_584,In_798);
and U988 (N_988,In_537,In_981);
or U989 (N_989,In_318,In_28);
or U990 (N_990,In_123,In_164);
or U991 (N_991,In_306,In_224);
and U992 (N_992,In_663,In_228);
or U993 (N_993,In_521,In_793);
or U994 (N_994,In_393,In_344);
nor U995 (N_995,In_911,In_420);
and U996 (N_996,In_580,In_237);
and U997 (N_997,In_593,In_880);
and U998 (N_998,In_23,In_345);
xor U999 (N_999,In_531,In_443);
nand U1000 (N_1000,In_574,In_802);
nand U1001 (N_1001,In_187,In_686);
and U1002 (N_1002,In_201,In_351);
and U1003 (N_1003,In_613,In_837);
or U1004 (N_1004,In_632,In_209);
and U1005 (N_1005,In_321,In_27);
and U1006 (N_1006,In_228,In_225);
and U1007 (N_1007,In_999,In_723);
and U1008 (N_1008,In_361,In_360);
nor U1009 (N_1009,In_856,In_627);
and U1010 (N_1010,In_78,In_151);
or U1011 (N_1011,In_283,In_972);
nand U1012 (N_1012,In_196,In_234);
nor U1013 (N_1013,In_151,In_305);
or U1014 (N_1014,In_604,In_110);
or U1015 (N_1015,In_149,In_39);
or U1016 (N_1016,In_91,In_811);
nor U1017 (N_1017,In_840,In_311);
or U1018 (N_1018,In_515,In_673);
or U1019 (N_1019,In_379,In_529);
or U1020 (N_1020,In_282,In_361);
nand U1021 (N_1021,In_820,In_554);
or U1022 (N_1022,In_778,In_801);
and U1023 (N_1023,In_261,In_589);
and U1024 (N_1024,In_939,In_498);
nor U1025 (N_1025,In_997,In_939);
nor U1026 (N_1026,In_196,In_496);
nand U1027 (N_1027,In_491,In_283);
nor U1028 (N_1028,In_615,In_257);
and U1029 (N_1029,In_98,In_743);
nor U1030 (N_1030,In_879,In_860);
or U1031 (N_1031,In_46,In_249);
nor U1032 (N_1032,In_847,In_787);
and U1033 (N_1033,In_448,In_838);
and U1034 (N_1034,In_171,In_596);
or U1035 (N_1035,In_948,In_984);
nor U1036 (N_1036,In_171,In_164);
nand U1037 (N_1037,In_73,In_600);
and U1038 (N_1038,In_196,In_568);
and U1039 (N_1039,In_428,In_359);
or U1040 (N_1040,In_859,In_38);
or U1041 (N_1041,In_316,In_145);
nand U1042 (N_1042,In_301,In_598);
or U1043 (N_1043,In_487,In_939);
and U1044 (N_1044,In_787,In_919);
nand U1045 (N_1045,In_940,In_51);
nand U1046 (N_1046,In_126,In_269);
nor U1047 (N_1047,In_957,In_270);
or U1048 (N_1048,In_510,In_989);
nand U1049 (N_1049,In_412,In_593);
or U1050 (N_1050,In_537,In_18);
nand U1051 (N_1051,In_723,In_757);
nand U1052 (N_1052,In_384,In_881);
or U1053 (N_1053,In_675,In_579);
or U1054 (N_1054,In_207,In_174);
or U1055 (N_1055,In_128,In_135);
nor U1056 (N_1056,In_237,In_88);
nand U1057 (N_1057,In_404,In_336);
nand U1058 (N_1058,In_632,In_601);
nand U1059 (N_1059,In_547,In_933);
and U1060 (N_1060,In_602,In_519);
nor U1061 (N_1061,In_113,In_238);
or U1062 (N_1062,In_764,In_258);
nand U1063 (N_1063,In_800,In_673);
nand U1064 (N_1064,In_540,In_409);
or U1065 (N_1065,In_416,In_267);
nand U1066 (N_1066,In_392,In_867);
nand U1067 (N_1067,In_457,In_428);
nor U1068 (N_1068,In_36,In_174);
nand U1069 (N_1069,In_237,In_915);
and U1070 (N_1070,In_796,In_618);
or U1071 (N_1071,In_530,In_93);
or U1072 (N_1072,In_308,In_702);
or U1073 (N_1073,In_624,In_925);
and U1074 (N_1074,In_643,In_880);
nand U1075 (N_1075,In_694,In_482);
or U1076 (N_1076,In_875,In_439);
and U1077 (N_1077,In_259,In_506);
and U1078 (N_1078,In_335,In_253);
nand U1079 (N_1079,In_700,In_41);
or U1080 (N_1080,In_855,In_544);
and U1081 (N_1081,In_465,In_775);
and U1082 (N_1082,In_895,In_996);
nand U1083 (N_1083,In_57,In_743);
nand U1084 (N_1084,In_3,In_235);
or U1085 (N_1085,In_616,In_236);
nand U1086 (N_1086,In_656,In_733);
nor U1087 (N_1087,In_221,In_746);
or U1088 (N_1088,In_327,In_239);
or U1089 (N_1089,In_162,In_784);
nor U1090 (N_1090,In_102,In_487);
or U1091 (N_1091,In_39,In_547);
and U1092 (N_1092,In_343,In_347);
or U1093 (N_1093,In_669,In_504);
nand U1094 (N_1094,In_635,In_90);
nand U1095 (N_1095,In_768,In_290);
and U1096 (N_1096,In_393,In_748);
or U1097 (N_1097,In_650,In_900);
nand U1098 (N_1098,In_754,In_570);
nor U1099 (N_1099,In_410,In_362);
nand U1100 (N_1100,In_975,In_464);
or U1101 (N_1101,In_734,In_133);
nand U1102 (N_1102,In_352,In_653);
xnor U1103 (N_1103,In_887,In_548);
or U1104 (N_1104,In_142,In_873);
or U1105 (N_1105,In_255,In_698);
nand U1106 (N_1106,In_760,In_410);
nand U1107 (N_1107,In_354,In_989);
or U1108 (N_1108,In_96,In_272);
nand U1109 (N_1109,In_321,In_975);
nand U1110 (N_1110,In_789,In_393);
nand U1111 (N_1111,In_610,In_952);
nand U1112 (N_1112,In_748,In_675);
and U1113 (N_1113,In_227,In_204);
nor U1114 (N_1114,In_6,In_242);
or U1115 (N_1115,In_91,In_658);
nor U1116 (N_1116,In_721,In_720);
and U1117 (N_1117,In_125,In_849);
nand U1118 (N_1118,In_684,In_8);
nor U1119 (N_1119,In_588,In_597);
or U1120 (N_1120,In_751,In_834);
or U1121 (N_1121,In_531,In_802);
or U1122 (N_1122,In_15,In_756);
or U1123 (N_1123,In_892,In_362);
nand U1124 (N_1124,In_450,In_348);
nand U1125 (N_1125,In_252,In_33);
and U1126 (N_1126,In_758,In_343);
nand U1127 (N_1127,In_512,In_238);
nor U1128 (N_1128,In_64,In_703);
or U1129 (N_1129,In_200,In_534);
nor U1130 (N_1130,In_505,In_127);
nand U1131 (N_1131,In_203,In_835);
and U1132 (N_1132,In_871,In_365);
and U1133 (N_1133,In_934,In_809);
or U1134 (N_1134,In_535,In_767);
or U1135 (N_1135,In_203,In_461);
or U1136 (N_1136,In_863,In_656);
and U1137 (N_1137,In_891,In_846);
or U1138 (N_1138,In_589,In_175);
nor U1139 (N_1139,In_688,In_846);
or U1140 (N_1140,In_615,In_601);
nand U1141 (N_1141,In_441,In_157);
or U1142 (N_1142,In_480,In_242);
or U1143 (N_1143,In_677,In_593);
nand U1144 (N_1144,In_392,In_374);
and U1145 (N_1145,In_345,In_579);
nand U1146 (N_1146,In_416,In_759);
nand U1147 (N_1147,In_276,In_268);
nor U1148 (N_1148,In_331,In_891);
nand U1149 (N_1149,In_258,In_304);
nand U1150 (N_1150,In_786,In_592);
and U1151 (N_1151,In_721,In_128);
and U1152 (N_1152,In_310,In_494);
or U1153 (N_1153,In_962,In_576);
and U1154 (N_1154,In_181,In_824);
nor U1155 (N_1155,In_546,In_191);
nor U1156 (N_1156,In_151,In_805);
or U1157 (N_1157,In_501,In_852);
nor U1158 (N_1158,In_669,In_722);
or U1159 (N_1159,In_636,In_296);
or U1160 (N_1160,In_125,In_41);
nand U1161 (N_1161,In_776,In_639);
nor U1162 (N_1162,In_854,In_713);
and U1163 (N_1163,In_507,In_610);
nand U1164 (N_1164,In_605,In_397);
nand U1165 (N_1165,In_453,In_346);
nor U1166 (N_1166,In_584,In_308);
or U1167 (N_1167,In_705,In_90);
or U1168 (N_1168,In_218,In_514);
nand U1169 (N_1169,In_101,In_484);
nand U1170 (N_1170,In_599,In_210);
or U1171 (N_1171,In_652,In_343);
nand U1172 (N_1172,In_138,In_452);
and U1173 (N_1173,In_17,In_6);
and U1174 (N_1174,In_160,In_967);
nor U1175 (N_1175,In_871,In_157);
nor U1176 (N_1176,In_29,In_58);
nor U1177 (N_1177,In_35,In_846);
nor U1178 (N_1178,In_587,In_294);
nand U1179 (N_1179,In_906,In_347);
nor U1180 (N_1180,In_112,In_187);
and U1181 (N_1181,In_810,In_193);
nor U1182 (N_1182,In_104,In_788);
and U1183 (N_1183,In_702,In_52);
nor U1184 (N_1184,In_555,In_686);
and U1185 (N_1185,In_611,In_744);
or U1186 (N_1186,In_103,In_339);
nand U1187 (N_1187,In_460,In_105);
nand U1188 (N_1188,In_327,In_698);
nand U1189 (N_1189,In_206,In_794);
and U1190 (N_1190,In_686,In_50);
nand U1191 (N_1191,In_81,In_55);
nand U1192 (N_1192,In_30,In_827);
or U1193 (N_1193,In_492,In_352);
nor U1194 (N_1194,In_373,In_822);
and U1195 (N_1195,In_337,In_181);
nand U1196 (N_1196,In_383,In_163);
nand U1197 (N_1197,In_134,In_487);
nor U1198 (N_1198,In_360,In_301);
nand U1199 (N_1199,In_500,In_328);
nor U1200 (N_1200,In_282,In_261);
nand U1201 (N_1201,In_828,In_54);
nor U1202 (N_1202,In_591,In_495);
nor U1203 (N_1203,In_893,In_494);
or U1204 (N_1204,In_538,In_515);
nand U1205 (N_1205,In_3,In_781);
nor U1206 (N_1206,In_590,In_792);
and U1207 (N_1207,In_583,In_607);
xor U1208 (N_1208,In_703,In_411);
nor U1209 (N_1209,In_562,In_117);
nand U1210 (N_1210,In_398,In_803);
or U1211 (N_1211,In_122,In_994);
and U1212 (N_1212,In_516,In_751);
and U1213 (N_1213,In_11,In_31);
and U1214 (N_1214,In_822,In_694);
and U1215 (N_1215,In_456,In_866);
nor U1216 (N_1216,In_642,In_992);
nor U1217 (N_1217,In_554,In_301);
nand U1218 (N_1218,In_237,In_514);
or U1219 (N_1219,In_76,In_669);
nand U1220 (N_1220,In_903,In_299);
or U1221 (N_1221,In_420,In_594);
nor U1222 (N_1222,In_288,In_917);
nand U1223 (N_1223,In_80,In_159);
or U1224 (N_1224,In_341,In_108);
nand U1225 (N_1225,In_938,In_494);
and U1226 (N_1226,In_186,In_208);
nand U1227 (N_1227,In_65,In_190);
and U1228 (N_1228,In_537,In_730);
nand U1229 (N_1229,In_557,In_541);
nand U1230 (N_1230,In_637,In_914);
nand U1231 (N_1231,In_275,In_590);
nand U1232 (N_1232,In_347,In_672);
and U1233 (N_1233,In_680,In_328);
nand U1234 (N_1234,In_438,In_966);
nor U1235 (N_1235,In_321,In_351);
nor U1236 (N_1236,In_461,In_479);
nor U1237 (N_1237,In_948,In_857);
or U1238 (N_1238,In_11,In_456);
and U1239 (N_1239,In_748,In_403);
nor U1240 (N_1240,In_422,In_766);
or U1241 (N_1241,In_205,In_16);
and U1242 (N_1242,In_733,In_672);
or U1243 (N_1243,In_324,In_531);
nand U1244 (N_1244,In_391,In_229);
nand U1245 (N_1245,In_942,In_910);
nand U1246 (N_1246,In_199,In_459);
and U1247 (N_1247,In_270,In_329);
nand U1248 (N_1248,In_538,In_16);
and U1249 (N_1249,In_68,In_672);
or U1250 (N_1250,In_479,In_381);
or U1251 (N_1251,In_370,In_466);
nor U1252 (N_1252,In_606,In_457);
nand U1253 (N_1253,In_941,In_462);
nor U1254 (N_1254,In_953,In_78);
nand U1255 (N_1255,In_939,In_688);
nor U1256 (N_1256,In_542,In_534);
or U1257 (N_1257,In_970,In_816);
and U1258 (N_1258,In_822,In_608);
nor U1259 (N_1259,In_643,In_472);
nor U1260 (N_1260,In_836,In_740);
or U1261 (N_1261,In_339,In_922);
nand U1262 (N_1262,In_983,In_703);
nand U1263 (N_1263,In_391,In_284);
nor U1264 (N_1264,In_314,In_132);
nor U1265 (N_1265,In_725,In_848);
and U1266 (N_1266,In_908,In_210);
nor U1267 (N_1267,In_122,In_317);
or U1268 (N_1268,In_545,In_329);
or U1269 (N_1269,In_132,In_464);
nor U1270 (N_1270,In_297,In_80);
nor U1271 (N_1271,In_72,In_834);
nor U1272 (N_1272,In_38,In_735);
or U1273 (N_1273,In_778,In_10);
xor U1274 (N_1274,In_787,In_970);
nand U1275 (N_1275,In_419,In_694);
or U1276 (N_1276,In_732,In_846);
nand U1277 (N_1277,In_499,In_339);
or U1278 (N_1278,In_15,In_784);
and U1279 (N_1279,In_311,In_948);
and U1280 (N_1280,In_105,In_317);
and U1281 (N_1281,In_883,In_880);
nand U1282 (N_1282,In_164,In_15);
nor U1283 (N_1283,In_826,In_152);
and U1284 (N_1284,In_390,In_742);
nand U1285 (N_1285,In_919,In_93);
nor U1286 (N_1286,In_335,In_31);
nand U1287 (N_1287,In_754,In_473);
nor U1288 (N_1288,In_733,In_18);
and U1289 (N_1289,In_99,In_546);
and U1290 (N_1290,In_635,In_770);
and U1291 (N_1291,In_106,In_182);
or U1292 (N_1292,In_919,In_35);
nor U1293 (N_1293,In_927,In_817);
or U1294 (N_1294,In_20,In_770);
nor U1295 (N_1295,In_676,In_559);
nor U1296 (N_1296,In_321,In_103);
or U1297 (N_1297,In_590,In_860);
nand U1298 (N_1298,In_374,In_418);
nand U1299 (N_1299,In_104,In_579);
nand U1300 (N_1300,In_379,In_903);
nand U1301 (N_1301,In_361,In_858);
or U1302 (N_1302,In_132,In_964);
nor U1303 (N_1303,In_14,In_799);
nand U1304 (N_1304,In_169,In_22);
xor U1305 (N_1305,In_2,In_28);
nor U1306 (N_1306,In_617,In_460);
nor U1307 (N_1307,In_749,In_781);
nand U1308 (N_1308,In_204,In_104);
nor U1309 (N_1309,In_234,In_258);
and U1310 (N_1310,In_684,In_848);
and U1311 (N_1311,In_689,In_804);
and U1312 (N_1312,In_409,In_896);
nor U1313 (N_1313,In_84,In_93);
or U1314 (N_1314,In_42,In_679);
and U1315 (N_1315,In_169,In_556);
nor U1316 (N_1316,In_464,In_492);
nand U1317 (N_1317,In_281,In_465);
nor U1318 (N_1318,In_739,In_416);
or U1319 (N_1319,In_90,In_861);
or U1320 (N_1320,In_657,In_882);
nand U1321 (N_1321,In_687,In_469);
nand U1322 (N_1322,In_547,In_434);
and U1323 (N_1323,In_443,In_227);
nand U1324 (N_1324,In_452,In_66);
nand U1325 (N_1325,In_830,In_18);
nor U1326 (N_1326,In_602,In_523);
nor U1327 (N_1327,In_110,In_271);
nand U1328 (N_1328,In_519,In_33);
nand U1329 (N_1329,In_37,In_633);
and U1330 (N_1330,In_22,In_741);
nand U1331 (N_1331,In_742,In_497);
or U1332 (N_1332,In_622,In_239);
nor U1333 (N_1333,In_539,In_419);
or U1334 (N_1334,In_931,In_812);
or U1335 (N_1335,In_396,In_394);
and U1336 (N_1336,In_768,In_512);
nand U1337 (N_1337,In_21,In_143);
nand U1338 (N_1338,In_374,In_380);
nor U1339 (N_1339,In_435,In_5);
and U1340 (N_1340,In_703,In_158);
nor U1341 (N_1341,In_517,In_637);
and U1342 (N_1342,In_325,In_710);
nand U1343 (N_1343,In_724,In_416);
nor U1344 (N_1344,In_471,In_38);
nor U1345 (N_1345,In_173,In_493);
nand U1346 (N_1346,In_233,In_575);
nor U1347 (N_1347,In_747,In_110);
nand U1348 (N_1348,In_396,In_863);
nor U1349 (N_1349,In_754,In_210);
and U1350 (N_1350,In_10,In_825);
and U1351 (N_1351,In_274,In_677);
nor U1352 (N_1352,In_48,In_356);
nor U1353 (N_1353,In_905,In_605);
or U1354 (N_1354,In_205,In_563);
nand U1355 (N_1355,In_668,In_873);
nor U1356 (N_1356,In_568,In_975);
or U1357 (N_1357,In_330,In_782);
nor U1358 (N_1358,In_245,In_504);
and U1359 (N_1359,In_865,In_575);
or U1360 (N_1360,In_281,In_857);
nor U1361 (N_1361,In_189,In_895);
or U1362 (N_1362,In_593,In_683);
or U1363 (N_1363,In_141,In_698);
or U1364 (N_1364,In_730,In_151);
and U1365 (N_1365,In_303,In_393);
and U1366 (N_1366,In_172,In_47);
nand U1367 (N_1367,In_747,In_54);
nor U1368 (N_1368,In_998,In_113);
nor U1369 (N_1369,In_889,In_520);
nor U1370 (N_1370,In_318,In_48);
or U1371 (N_1371,In_91,In_555);
nand U1372 (N_1372,In_150,In_663);
and U1373 (N_1373,In_832,In_484);
nor U1374 (N_1374,In_643,In_92);
and U1375 (N_1375,In_118,In_240);
nor U1376 (N_1376,In_989,In_446);
or U1377 (N_1377,In_453,In_340);
and U1378 (N_1378,In_152,In_503);
and U1379 (N_1379,In_914,In_870);
nand U1380 (N_1380,In_802,In_268);
or U1381 (N_1381,In_253,In_865);
or U1382 (N_1382,In_627,In_934);
nand U1383 (N_1383,In_228,In_939);
nor U1384 (N_1384,In_705,In_794);
or U1385 (N_1385,In_332,In_915);
or U1386 (N_1386,In_6,In_226);
nand U1387 (N_1387,In_968,In_742);
nor U1388 (N_1388,In_359,In_554);
nor U1389 (N_1389,In_123,In_855);
or U1390 (N_1390,In_197,In_352);
or U1391 (N_1391,In_565,In_383);
and U1392 (N_1392,In_343,In_180);
nor U1393 (N_1393,In_480,In_943);
nor U1394 (N_1394,In_482,In_944);
or U1395 (N_1395,In_601,In_613);
and U1396 (N_1396,In_463,In_336);
or U1397 (N_1397,In_570,In_990);
nor U1398 (N_1398,In_576,In_446);
and U1399 (N_1399,In_641,In_727);
nor U1400 (N_1400,In_633,In_848);
nor U1401 (N_1401,In_947,In_562);
and U1402 (N_1402,In_335,In_688);
and U1403 (N_1403,In_823,In_707);
and U1404 (N_1404,In_246,In_103);
or U1405 (N_1405,In_32,In_300);
nand U1406 (N_1406,In_964,In_616);
and U1407 (N_1407,In_308,In_745);
nor U1408 (N_1408,In_177,In_866);
nand U1409 (N_1409,In_368,In_358);
or U1410 (N_1410,In_112,In_227);
nor U1411 (N_1411,In_810,In_615);
nor U1412 (N_1412,In_480,In_356);
or U1413 (N_1413,In_641,In_285);
or U1414 (N_1414,In_452,In_974);
and U1415 (N_1415,In_196,In_520);
nand U1416 (N_1416,In_249,In_88);
or U1417 (N_1417,In_947,In_593);
and U1418 (N_1418,In_788,In_21);
or U1419 (N_1419,In_775,In_206);
nor U1420 (N_1420,In_795,In_508);
or U1421 (N_1421,In_414,In_410);
and U1422 (N_1422,In_505,In_227);
or U1423 (N_1423,In_482,In_416);
and U1424 (N_1424,In_715,In_826);
or U1425 (N_1425,In_797,In_120);
and U1426 (N_1426,In_436,In_451);
nand U1427 (N_1427,In_384,In_214);
nor U1428 (N_1428,In_889,In_69);
nor U1429 (N_1429,In_673,In_848);
or U1430 (N_1430,In_141,In_7);
and U1431 (N_1431,In_289,In_843);
nand U1432 (N_1432,In_448,In_452);
nand U1433 (N_1433,In_221,In_719);
nand U1434 (N_1434,In_374,In_371);
nand U1435 (N_1435,In_761,In_107);
nor U1436 (N_1436,In_715,In_52);
and U1437 (N_1437,In_791,In_366);
or U1438 (N_1438,In_131,In_358);
nand U1439 (N_1439,In_418,In_156);
nand U1440 (N_1440,In_63,In_245);
nand U1441 (N_1441,In_405,In_264);
nor U1442 (N_1442,In_921,In_210);
and U1443 (N_1443,In_215,In_731);
nand U1444 (N_1444,In_792,In_498);
nor U1445 (N_1445,In_314,In_307);
or U1446 (N_1446,In_32,In_235);
or U1447 (N_1447,In_641,In_378);
or U1448 (N_1448,In_65,In_157);
or U1449 (N_1449,In_797,In_832);
nand U1450 (N_1450,In_353,In_734);
or U1451 (N_1451,In_510,In_468);
and U1452 (N_1452,In_487,In_312);
nor U1453 (N_1453,In_854,In_990);
or U1454 (N_1454,In_383,In_446);
nand U1455 (N_1455,In_386,In_797);
or U1456 (N_1456,In_899,In_716);
or U1457 (N_1457,In_722,In_610);
or U1458 (N_1458,In_199,In_321);
nand U1459 (N_1459,In_197,In_980);
or U1460 (N_1460,In_621,In_486);
and U1461 (N_1461,In_771,In_837);
or U1462 (N_1462,In_597,In_917);
or U1463 (N_1463,In_575,In_170);
xnor U1464 (N_1464,In_346,In_301);
and U1465 (N_1465,In_584,In_262);
and U1466 (N_1466,In_191,In_793);
nand U1467 (N_1467,In_209,In_547);
and U1468 (N_1468,In_215,In_125);
or U1469 (N_1469,In_113,In_887);
or U1470 (N_1470,In_242,In_44);
nand U1471 (N_1471,In_857,In_200);
or U1472 (N_1472,In_855,In_636);
nand U1473 (N_1473,In_873,In_136);
nor U1474 (N_1474,In_122,In_106);
nand U1475 (N_1475,In_237,In_868);
nand U1476 (N_1476,In_396,In_959);
and U1477 (N_1477,In_19,In_465);
or U1478 (N_1478,In_601,In_374);
and U1479 (N_1479,In_128,In_945);
and U1480 (N_1480,In_509,In_658);
nor U1481 (N_1481,In_647,In_729);
nand U1482 (N_1482,In_837,In_648);
nor U1483 (N_1483,In_354,In_869);
or U1484 (N_1484,In_200,In_760);
or U1485 (N_1485,In_385,In_142);
or U1486 (N_1486,In_866,In_260);
or U1487 (N_1487,In_973,In_703);
nor U1488 (N_1488,In_10,In_588);
and U1489 (N_1489,In_720,In_799);
or U1490 (N_1490,In_439,In_68);
nor U1491 (N_1491,In_875,In_4);
nand U1492 (N_1492,In_435,In_495);
xor U1493 (N_1493,In_70,In_305);
or U1494 (N_1494,In_817,In_816);
or U1495 (N_1495,In_127,In_533);
or U1496 (N_1496,In_979,In_387);
nor U1497 (N_1497,In_917,In_465);
nand U1498 (N_1498,In_468,In_904);
nand U1499 (N_1499,In_352,In_842);
xnor U1500 (N_1500,In_630,In_698);
nand U1501 (N_1501,In_939,In_728);
and U1502 (N_1502,In_296,In_362);
and U1503 (N_1503,In_239,In_605);
or U1504 (N_1504,In_468,In_185);
nand U1505 (N_1505,In_609,In_55);
nor U1506 (N_1506,In_556,In_458);
nor U1507 (N_1507,In_94,In_505);
or U1508 (N_1508,In_770,In_866);
nor U1509 (N_1509,In_340,In_761);
nor U1510 (N_1510,In_833,In_840);
nand U1511 (N_1511,In_166,In_490);
and U1512 (N_1512,In_541,In_804);
nand U1513 (N_1513,In_898,In_976);
nor U1514 (N_1514,In_35,In_717);
or U1515 (N_1515,In_673,In_389);
nand U1516 (N_1516,In_113,In_792);
or U1517 (N_1517,In_707,In_251);
nand U1518 (N_1518,In_919,In_575);
xnor U1519 (N_1519,In_934,In_813);
and U1520 (N_1520,In_608,In_650);
and U1521 (N_1521,In_741,In_949);
and U1522 (N_1522,In_179,In_456);
nand U1523 (N_1523,In_235,In_709);
and U1524 (N_1524,In_198,In_772);
and U1525 (N_1525,In_360,In_975);
and U1526 (N_1526,In_875,In_83);
nand U1527 (N_1527,In_91,In_477);
nand U1528 (N_1528,In_631,In_949);
nand U1529 (N_1529,In_235,In_267);
or U1530 (N_1530,In_858,In_346);
or U1531 (N_1531,In_690,In_345);
nor U1532 (N_1532,In_515,In_864);
and U1533 (N_1533,In_660,In_867);
and U1534 (N_1534,In_405,In_623);
nand U1535 (N_1535,In_220,In_856);
or U1536 (N_1536,In_17,In_960);
and U1537 (N_1537,In_738,In_216);
nor U1538 (N_1538,In_324,In_991);
and U1539 (N_1539,In_574,In_352);
and U1540 (N_1540,In_728,In_721);
or U1541 (N_1541,In_279,In_487);
or U1542 (N_1542,In_296,In_879);
nand U1543 (N_1543,In_96,In_531);
nor U1544 (N_1544,In_822,In_771);
nor U1545 (N_1545,In_309,In_574);
nor U1546 (N_1546,In_280,In_811);
or U1547 (N_1547,In_717,In_45);
or U1548 (N_1548,In_55,In_283);
nor U1549 (N_1549,In_854,In_186);
and U1550 (N_1550,In_850,In_104);
nand U1551 (N_1551,In_971,In_493);
and U1552 (N_1552,In_266,In_626);
and U1553 (N_1553,In_846,In_896);
nand U1554 (N_1554,In_424,In_313);
or U1555 (N_1555,In_145,In_604);
or U1556 (N_1556,In_163,In_446);
and U1557 (N_1557,In_433,In_200);
or U1558 (N_1558,In_340,In_365);
nor U1559 (N_1559,In_129,In_471);
and U1560 (N_1560,In_924,In_126);
or U1561 (N_1561,In_156,In_543);
and U1562 (N_1562,In_336,In_236);
nor U1563 (N_1563,In_716,In_542);
and U1564 (N_1564,In_800,In_285);
nand U1565 (N_1565,In_583,In_743);
and U1566 (N_1566,In_609,In_765);
nand U1567 (N_1567,In_210,In_968);
nor U1568 (N_1568,In_626,In_961);
and U1569 (N_1569,In_641,In_397);
nand U1570 (N_1570,In_818,In_866);
nor U1571 (N_1571,In_364,In_675);
nor U1572 (N_1572,In_294,In_66);
nor U1573 (N_1573,In_871,In_481);
or U1574 (N_1574,In_456,In_674);
and U1575 (N_1575,In_372,In_703);
nand U1576 (N_1576,In_800,In_614);
nor U1577 (N_1577,In_383,In_60);
nand U1578 (N_1578,In_847,In_574);
or U1579 (N_1579,In_298,In_632);
or U1580 (N_1580,In_161,In_304);
nor U1581 (N_1581,In_42,In_586);
nand U1582 (N_1582,In_34,In_526);
or U1583 (N_1583,In_523,In_299);
or U1584 (N_1584,In_264,In_961);
nand U1585 (N_1585,In_700,In_931);
or U1586 (N_1586,In_741,In_377);
nand U1587 (N_1587,In_513,In_10);
or U1588 (N_1588,In_0,In_540);
and U1589 (N_1589,In_538,In_150);
nand U1590 (N_1590,In_399,In_565);
and U1591 (N_1591,In_45,In_361);
and U1592 (N_1592,In_628,In_238);
or U1593 (N_1593,In_80,In_301);
nor U1594 (N_1594,In_574,In_360);
or U1595 (N_1595,In_215,In_107);
or U1596 (N_1596,In_13,In_672);
nor U1597 (N_1597,In_809,In_327);
nor U1598 (N_1598,In_566,In_953);
and U1599 (N_1599,In_815,In_739);
and U1600 (N_1600,In_255,In_344);
and U1601 (N_1601,In_770,In_120);
nand U1602 (N_1602,In_483,In_618);
or U1603 (N_1603,In_572,In_503);
nand U1604 (N_1604,In_612,In_283);
xnor U1605 (N_1605,In_891,In_148);
or U1606 (N_1606,In_148,In_882);
nor U1607 (N_1607,In_959,In_296);
or U1608 (N_1608,In_656,In_347);
or U1609 (N_1609,In_105,In_841);
nand U1610 (N_1610,In_907,In_734);
nor U1611 (N_1611,In_982,In_623);
nand U1612 (N_1612,In_271,In_648);
nor U1613 (N_1613,In_818,In_439);
or U1614 (N_1614,In_812,In_118);
nor U1615 (N_1615,In_556,In_343);
nand U1616 (N_1616,In_894,In_685);
nand U1617 (N_1617,In_785,In_836);
nand U1618 (N_1618,In_381,In_366);
or U1619 (N_1619,In_188,In_918);
nand U1620 (N_1620,In_9,In_546);
or U1621 (N_1621,In_284,In_946);
nor U1622 (N_1622,In_512,In_27);
nor U1623 (N_1623,In_864,In_288);
or U1624 (N_1624,In_556,In_763);
nand U1625 (N_1625,In_143,In_714);
nor U1626 (N_1626,In_45,In_195);
or U1627 (N_1627,In_49,In_605);
and U1628 (N_1628,In_523,In_184);
nor U1629 (N_1629,In_10,In_405);
nor U1630 (N_1630,In_147,In_815);
or U1631 (N_1631,In_315,In_496);
nand U1632 (N_1632,In_247,In_264);
and U1633 (N_1633,In_273,In_662);
nor U1634 (N_1634,In_155,In_330);
or U1635 (N_1635,In_119,In_757);
or U1636 (N_1636,In_673,In_363);
nor U1637 (N_1637,In_605,In_711);
or U1638 (N_1638,In_19,In_474);
and U1639 (N_1639,In_684,In_800);
or U1640 (N_1640,In_195,In_171);
nor U1641 (N_1641,In_159,In_541);
and U1642 (N_1642,In_655,In_583);
or U1643 (N_1643,In_843,In_826);
or U1644 (N_1644,In_861,In_947);
or U1645 (N_1645,In_863,In_456);
nor U1646 (N_1646,In_36,In_478);
or U1647 (N_1647,In_485,In_176);
nor U1648 (N_1648,In_211,In_869);
nor U1649 (N_1649,In_316,In_0);
nand U1650 (N_1650,In_366,In_579);
nor U1651 (N_1651,In_861,In_957);
nor U1652 (N_1652,In_495,In_227);
and U1653 (N_1653,In_383,In_609);
nor U1654 (N_1654,In_588,In_355);
nor U1655 (N_1655,In_46,In_887);
and U1656 (N_1656,In_649,In_437);
or U1657 (N_1657,In_976,In_887);
nand U1658 (N_1658,In_743,In_847);
and U1659 (N_1659,In_905,In_407);
nor U1660 (N_1660,In_369,In_266);
nor U1661 (N_1661,In_197,In_2);
or U1662 (N_1662,In_895,In_848);
nor U1663 (N_1663,In_286,In_489);
nor U1664 (N_1664,In_710,In_527);
nor U1665 (N_1665,In_519,In_302);
nand U1666 (N_1666,In_457,In_113);
nor U1667 (N_1667,In_719,In_274);
nand U1668 (N_1668,In_802,In_893);
or U1669 (N_1669,In_297,In_487);
nor U1670 (N_1670,In_57,In_969);
or U1671 (N_1671,In_188,In_454);
or U1672 (N_1672,In_115,In_596);
and U1673 (N_1673,In_824,In_881);
nor U1674 (N_1674,In_112,In_50);
and U1675 (N_1675,In_956,In_289);
and U1676 (N_1676,In_772,In_507);
and U1677 (N_1677,In_446,In_944);
nand U1678 (N_1678,In_372,In_518);
nand U1679 (N_1679,In_654,In_348);
or U1680 (N_1680,In_795,In_548);
and U1681 (N_1681,In_161,In_630);
and U1682 (N_1682,In_468,In_226);
or U1683 (N_1683,In_699,In_922);
or U1684 (N_1684,In_291,In_859);
and U1685 (N_1685,In_952,In_473);
nor U1686 (N_1686,In_234,In_416);
or U1687 (N_1687,In_243,In_736);
and U1688 (N_1688,In_188,In_659);
nor U1689 (N_1689,In_866,In_375);
nand U1690 (N_1690,In_293,In_861);
nor U1691 (N_1691,In_892,In_999);
nand U1692 (N_1692,In_76,In_355);
or U1693 (N_1693,In_985,In_126);
and U1694 (N_1694,In_29,In_124);
and U1695 (N_1695,In_131,In_868);
or U1696 (N_1696,In_959,In_586);
and U1697 (N_1697,In_153,In_693);
nor U1698 (N_1698,In_233,In_658);
or U1699 (N_1699,In_612,In_82);
nand U1700 (N_1700,In_799,In_639);
and U1701 (N_1701,In_728,In_464);
or U1702 (N_1702,In_544,In_600);
nor U1703 (N_1703,In_222,In_750);
nor U1704 (N_1704,In_523,In_161);
nor U1705 (N_1705,In_665,In_710);
nor U1706 (N_1706,In_295,In_58);
nor U1707 (N_1707,In_917,In_292);
nor U1708 (N_1708,In_791,In_118);
or U1709 (N_1709,In_454,In_286);
nor U1710 (N_1710,In_666,In_719);
or U1711 (N_1711,In_343,In_105);
nand U1712 (N_1712,In_165,In_836);
or U1713 (N_1713,In_423,In_497);
or U1714 (N_1714,In_293,In_422);
and U1715 (N_1715,In_549,In_922);
nor U1716 (N_1716,In_707,In_534);
and U1717 (N_1717,In_430,In_0);
nor U1718 (N_1718,In_759,In_578);
nand U1719 (N_1719,In_356,In_822);
nor U1720 (N_1720,In_15,In_483);
nor U1721 (N_1721,In_8,In_87);
or U1722 (N_1722,In_655,In_714);
nor U1723 (N_1723,In_920,In_134);
or U1724 (N_1724,In_790,In_12);
nor U1725 (N_1725,In_152,In_735);
or U1726 (N_1726,In_289,In_887);
and U1727 (N_1727,In_383,In_221);
nand U1728 (N_1728,In_404,In_89);
xor U1729 (N_1729,In_184,In_652);
nand U1730 (N_1730,In_593,In_699);
or U1731 (N_1731,In_675,In_431);
or U1732 (N_1732,In_679,In_754);
nor U1733 (N_1733,In_523,In_687);
nand U1734 (N_1734,In_669,In_166);
and U1735 (N_1735,In_134,In_259);
nand U1736 (N_1736,In_994,In_19);
nor U1737 (N_1737,In_94,In_695);
nand U1738 (N_1738,In_837,In_73);
nand U1739 (N_1739,In_283,In_170);
nand U1740 (N_1740,In_405,In_947);
and U1741 (N_1741,In_465,In_10);
nand U1742 (N_1742,In_145,In_255);
nor U1743 (N_1743,In_771,In_865);
nor U1744 (N_1744,In_673,In_610);
or U1745 (N_1745,In_122,In_577);
or U1746 (N_1746,In_280,In_379);
nand U1747 (N_1747,In_290,In_200);
and U1748 (N_1748,In_225,In_456);
or U1749 (N_1749,In_42,In_950);
or U1750 (N_1750,In_749,In_652);
nand U1751 (N_1751,In_896,In_437);
nor U1752 (N_1752,In_866,In_424);
and U1753 (N_1753,In_865,In_148);
nand U1754 (N_1754,In_681,In_139);
nor U1755 (N_1755,In_47,In_450);
and U1756 (N_1756,In_982,In_275);
nor U1757 (N_1757,In_16,In_114);
or U1758 (N_1758,In_740,In_461);
nor U1759 (N_1759,In_982,In_848);
nor U1760 (N_1760,In_559,In_613);
nand U1761 (N_1761,In_42,In_724);
nand U1762 (N_1762,In_247,In_595);
nand U1763 (N_1763,In_371,In_57);
xnor U1764 (N_1764,In_224,In_628);
and U1765 (N_1765,In_764,In_532);
nand U1766 (N_1766,In_826,In_652);
nor U1767 (N_1767,In_683,In_831);
nand U1768 (N_1768,In_921,In_634);
or U1769 (N_1769,In_451,In_396);
and U1770 (N_1770,In_12,In_531);
and U1771 (N_1771,In_209,In_948);
and U1772 (N_1772,In_826,In_464);
nor U1773 (N_1773,In_637,In_202);
nand U1774 (N_1774,In_533,In_3);
and U1775 (N_1775,In_28,In_8);
or U1776 (N_1776,In_867,In_468);
or U1777 (N_1777,In_337,In_33);
and U1778 (N_1778,In_853,In_87);
nand U1779 (N_1779,In_968,In_431);
and U1780 (N_1780,In_96,In_462);
or U1781 (N_1781,In_312,In_0);
or U1782 (N_1782,In_160,In_74);
nor U1783 (N_1783,In_635,In_338);
and U1784 (N_1784,In_861,In_185);
and U1785 (N_1785,In_530,In_444);
or U1786 (N_1786,In_746,In_365);
nand U1787 (N_1787,In_305,In_174);
nor U1788 (N_1788,In_241,In_555);
and U1789 (N_1789,In_71,In_756);
nor U1790 (N_1790,In_334,In_628);
and U1791 (N_1791,In_933,In_761);
nor U1792 (N_1792,In_642,In_413);
or U1793 (N_1793,In_519,In_521);
or U1794 (N_1794,In_715,In_631);
and U1795 (N_1795,In_96,In_149);
or U1796 (N_1796,In_697,In_508);
xor U1797 (N_1797,In_489,In_334);
and U1798 (N_1798,In_37,In_888);
nor U1799 (N_1799,In_243,In_869);
and U1800 (N_1800,In_913,In_660);
or U1801 (N_1801,In_695,In_830);
nand U1802 (N_1802,In_636,In_11);
nor U1803 (N_1803,In_310,In_597);
nand U1804 (N_1804,In_316,In_430);
or U1805 (N_1805,In_782,In_668);
nand U1806 (N_1806,In_420,In_335);
and U1807 (N_1807,In_317,In_921);
and U1808 (N_1808,In_190,In_134);
nand U1809 (N_1809,In_301,In_769);
nand U1810 (N_1810,In_78,In_8);
nor U1811 (N_1811,In_856,In_814);
and U1812 (N_1812,In_660,In_451);
or U1813 (N_1813,In_357,In_255);
nor U1814 (N_1814,In_234,In_536);
and U1815 (N_1815,In_799,In_468);
and U1816 (N_1816,In_144,In_17);
or U1817 (N_1817,In_749,In_106);
and U1818 (N_1818,In_126,In_634);
nand U1819 (N_1819,In_83,In_473);
or U1820 (N_1820,In_746,In_62);
or U1821 (N_1821,In_206,In_528);
nand U1822 (N_1822,In_331,In_819);
and U1823 (N_1823,In_173,In_82);
and U1824 (N_1824,In_36,In_0);
nor U1825 (N_1825,In_418,In_587);
or U1826 (N_1826,In_884,In_674);
nand U1827 (N_1827,In_151,In_688);
and U1828 (N_1828,In_117,In_115);
xor U1829 (N_1829,In_245,In_208);
nand U1830 (N_1830,In_996,In_734);
or U1831 (N_1831,In_141,In_979);
and U1832 (N_1832,In_131,In_476);
and U1833 (N_1833,In_749,In_83);
and U1834 (N_1834,In_916,In_616);
nor U1835 (N_1835,In_995,In_476);
nand U1836 (N_1836,In_853,In_301);
or U1837 (N_1837,In_29,In_292);
or U1838 (N_1838,In_343,In_283);
nand U1839 (N_1839,In_132,In_348);
and U1840 (N_1840,In_421,In_443);
and U1841 (N_1841,In_270,In_219);
or U1842 (N_1842,In_223,In_137);
nand U1843 (N_1843,In_496,In_922);
or U1844 (N_1844,In_165,In_210);
and U1845 (N_1845,In_668,In_364);
or U1846 (N_1846,In_366,In_352);
and U1847 (N_1847,In_801,In_541);
nor U1848 (N_1848,In_180,In_706);
nor U1849 (N_1849,In_515,In_38);
nand U1850 (N_1850,In_344,In_10);
and U1851 (N_1851,In_152,In_751);
and U1852 (N_1852,In_136,In_908);
or U1853 (N_1853,In_230,In_677);
nor U1854 (N_1854,In_387,In_144);
and U1855 (N_1855,In_21,In_623);
nand U1856 (N_1856,In_90,In_291);
nor U1857 (N_1857,In_242,In_386);
nor U1858 (N_1858,In_811,In_501);
or U1859 (N_1859,In_536,In_321);
nor U1860 (N_1860,In_940,In_63);
nor U1861 (N_1861,In_938,In_623);
nor U1862 (N_1862,In_767,In_458);
and U1863 (N_1863,In_902,In_401);
or U1864 (N_1864,In_332,In_243);
and U1865 (N_1865,In_516,In_908);
and U1866 (N_1866,In_524,In_582);
or U1867 (N_1867,In_791,In_62);
nor U1868 (N_1868,In_822,In_458);
nor U1869 (N_1869,In_524,In_760);
nor U1870 (N_1870,In_751,In_928);
or U1871 (N_1871,In_980,In_760);
nand U1872 (N_1872,In_651,In_456);
or U1873 (N_1873,In_413,In_346);
and U1874 (N_1874,In_911,In_996);
or U1875 (N_1875,In_577,In_944);
and U1876 (N_1876,In_529,In_94);
nor U1877 (N_1877,In_422,In_307);
nand U1878 (N_1878,In_620,In_367);
nand U1879 (N_1879,In_581,In_917);
or U1880 (N_1880,In_703,In_29);
nor U1881 (N_1881,In_451,In_641);
and U1882 (N_1882,In_174,In_651);
or U1883 (N_1883,In_776,In_122);
nor U1884 (N_1884,In_669,In_357);
and U1885 (N_1885,In_748,In_292);
and U1886 (N_1886,In_224,In_803);
nand U1887 (N_1887,In_447,In_984);
nand U1888 (N_1888,In_952,In_806);
nor U1889 (N_1889,In_602,In_42);
nand U1890 (N_1890,In_935,In_946);
nand U1891 (N_1891,In_673,In_731);
and U1892 (N_1892,In_347,In_949);
xnor U1893 (N_1893,In_251,In_986);
and U1894 (N_1894,In_640,In_401);
nor U1895 (N_1895,In_499,In_19);
nor U1896 (N_1896,In_435,In_459);
nand U1897 (N_1897,In_671,In_957);
and U1898 (N_1898,In_240,In_920);
and U1899 (N_1899,In_609,In_899);
or U1900 (N_1900,In_425,In_924);
and U1901 (N_1901,In_576,In_454);
and U1902 (N_1902,In_52,In_158);
nor U1903 (N_1903,In_47,In_466);
nand U1904 (N_1904,In_26,In_504);
or U1905 (N_1905,In_590,In_951);
and U1906 (N_1906,In_814,In_815);
and U1907 (N_1907,In_313,In_470);
nand U1908 (N_1908,In_361,In_81);
and U1909 (N_1909,In_562,In_923);
nor U1910 (N_1910,In_92,In_854);
nor U1911 (N_1911,In_424,In_156);
nand U1912 (N_1912,In_850,In_689);
nand U1913 (N_1913,In_855,In_656);
nand U1914 (N_1914,In_932,In_362);
nand U1915 (N_1915,In_815,In_743);
nand U1916 (N_1916,In_598,In_225);
nand U1917 (N_1917,In_419,In_525);
nor U1918 (N_1918,In_678,In_128);
and U1919 (N_1919,In_351,In_349);
nor U1920 (N_1920,In_659,In_173);
or U1921 (N_1921,In_427,In_746);
nand U1922 (N_1922,In_292,In_177);
nor U1923 (N_1923,In_313,In_623);
or U1924 (N_1924,In_643,In_172);
and U1925 (N_1925,In_965,In_28);
and U1926 (N_1926,In_173,In_226);
nor U1927 (N_1927,In_512,In_74);
nand U1928 (N_1928,In_0,In_919);
or U1929 (N_1929,In_553,In_676);
and U1930 (N_1930,In_822,In_528);
and U1931 (N_1931,In_886,In_119);
nor U1932 (N_1932,In_804,In_464);
nand U1933 (N_1933,In_615,In_916);
nand U1934 (N_1934,In_914,In_673);
or U1935 (N_1935,In_599,In_126);
nand U1936 (N_1936,In_831,In_149);
nand U1937 (N_1937,In_403,In_375);
or U1938 (N_1938,In_43,In_848);
nor U1939 (N_1939,In_476,In_732);
or U1940 (N_1940,In_376,In_63);
or U1941 (N_1941,In_542,In_518);
nand U1942 (N_1942,In_586,In_378);
and U1943 (N_1943,In_154,In_123);
nor U1944 (N_1944,In_212,In_669);
and U1945 (N_1945,In_576,In_769);
and U1946 (N_1946,In_252,In_140);
nand U1947 (N_1947,In_205,In_576);
nand U1948 (N_1948,In_821,In_290);
or U1949 (N_1949,In_593,In_842);
and U1950 (N_1950,In_780,In_201);
and U1951 (N_1951,In_401,In_853);
or U1952 (N_1952,In_102,In_277);
nand U1953 (N_1953,In_268,In_770);
nor U1954 (N_1954,In_904,In_326);
nand U1955 (N_1955,In_564,In_173);
nor U1956 (N_1956,In_212,In_779);
or U1957 (N_1957,In_960,In_378);
nor U1958 (N_1958,In_385,In_349);
or U1959 (N_1959,In_878,In_880);
nand U1960 (N_1960,In_270,In_363);
nand U1961 (N_1961,In_153,In_790);
nor U1962 (N_1962,In_80,In_334);
nand U1963 (N_1963,In_913,In_385);
nand U1964 (N_1964,In_360,In_639);
nor U1965 (N_1965,In_980,In_298);
nor U1966 (N_1966,In_697,In_576);
nor U1967 (N_1967,In_220,In_943);
and U1968 (N_1968,In_71,In_125);
nor U1969 (N_1969,In_977,In_244);
nor U1970 (N_1970,In_988,In_18);
or U1971 (N_1971,In_949,In_657);
nand U1972 (N_1972,In_361,In_408);
nor U1973 (N_1973,In_828,In_935);
nand U1974 (N_1974,In_697,In_493);
and U1975 (N_1975,In_349,In_412);
nor U1976 (N_1976,In_953,In_67);
or U1977 (N_1977,In_794,In_134);
and U1978 (N_1978,In_595,In_717);
and U1979 (N_1979,In_17,In_730);
or U1980 (N_1980,In_880,In_6);
and U1981 (N_1981,In_767,In_313);
and U1982 (N_1982,In_345,In_727);
nor U1983 (N_1983,In_773,In_909);
nor U1984 (N_1984,In_182,In_289);
and U1985 (N_1985,In_964,In_567);
or U1986 (N_1986,In_986,In_794);
nor U1987 (N_1987,In_988,In_866);
xnor U1988 (N_1988,In_612,In_426);
and U1989 (N_1989,In_732,In_126);
nand U1990 (N_1990,In_117,In_957);
or U1991 (N_1991,In_673,In_894);
or U1992 (N_1992,In_478,In_914);
nand U1993 (N_1993,In_412,In_856);
and U1994 (N_1994,In_700,In_85);
or U1995 (N_1995,In_950,In_335);
or U1996 (N_1996,In_785,In_397);
nor U1997 (N_1997,In_920,In_797);
nor U1998 (N_1998,In_578,In_811);
or U1999 (N_1999,In_342,In_882);
nand U2000 (N_2000,In_448,In_45);
and U2001 (N_2001,In_758,In_706);
nor U2002 (N_2002,In_954,In_335);
nand U2003 (N_2003,In_478,In_604);
and U2004 (N_2004,In_739,In_347);
nor U2005 (N_2005,In_917,In_647);
nand U2006 (N_2006,In_128,In_820);
nand U2007 (N_2007,In_194,In_334);
nand U2008 (N_2008,In_176,In_351);
nand U2009 (N_2009,In_377,In_860);
nand U2010 (N_2010,In_707,In_302);
nand U2011 (N_2011,In_276,In_458);
nor U2012 (N_2012,In_137,In_509);
nor U2013 (N_2013,In_3,In_119);
nor U2014 (N_2014,In_385,In_957);
or U2015 (N_2015,In_18,In_217);
nor U2016 (N_2016,In_715,In_946);
nor U2017 (N_2017,In_647,In_66);
and U2018 (N_2018,In_666,In_35);
or U2019 (N_2019,In_195,In_468);
or U2020 (N_2020,In_72,In_839);
nor U2021 (N_2021,In_9,In_816);
and U2022 (N_2022,In_360,In_809);
and U2023 (N_2023,In_92,In_718);
or U2024 (N_2024,In_830,In_453);
nor U2025 (N_2025,In_359,In_677);
or U2026 (N_2026,In_445,In_518);
nand U2027 (N_2027,In_354,In_510);
nand U2028 (N_2028,In_419,In_706);
and U2029 (N_2029,In_244,In_481);
or U2030 (N_2030,In_752,In_110);
nand U2031 (N_2031,In_645,In_971);
nor U2032 (N_2032,In_729,In_506);
and U2033 (N_2033,In_16,In_437);
nand U2034 (N_2034,In_749,In_955);
nand U2035 (N_2035,In_52,In_515);
nor U2036 (N_2036,In_157,In_28);
or U2037 (N_2037,In_673,In_104);
nand U2038 (N_2038,In_46,In_442);
or U2039 (N_2039,In_296,In_404);
or U2040 (N_2040,In_163,In_675);
and U2041 (N_2041,In_681,In_815);
nand U2042 (N_2042,In_594,In_416);
nand U2043 (N_2043,In_447,In_41);
nor U2044 (N_2044,In_727,In_286);
and U2045 (N_2045,In_136,In_924);
nand U2046 (N_2046,In_117,In_409);
nor U2047 (N_2047,In_997,In_454);
nor U2048 (N_2048,In_919,In_856);
or U2049 (N_2049,In_857,In_461);
xnor U2050 (N_2050,In_899,In_949);
or U2051 (N_2051,In_7,In_144);
or U2052 (N_2052,In_751,In_269);
and U2053 (N_2053,In_865,In_783);
nor U2054 (N_2054,In_667,In_2);
or U2055 (N_2055,In_710,In_822);
or U2056 (N_2056,In_964,In_66);
and U2057 (N_2057,In_466,In_375);
nor U2058 (N_2058,In_634,In_937);
and U2059 (N_2059,In_897,In_358);
or U2060 (N_2060,In_66,In_368);
nand U2061 (N_2061,In_241,In_419);
nand U2062 (N_2062,In_978,In_814);
nor U2063 (N_2063,In_676,In_703);
nor U2064 (N_2064,In_386,In_983);
or U2065 (N_2065,In_443,In_614);
nor U2066 (N_2066,In_507,In_416);
and U2067 (N_2067,In_337,In_994);
nor U2068 (N_2068,In_617,In_264);
or U2069 (N_2069,In_413,In_923);
or U2070 (N_2070,In_502,In_939);
or U2071 (N_2071,In_798,In_975);
nor U2072 (N_2072,In_576,In_480);
xor U2073 (N_2073,In_896,In_921);
nand U2074 (N_2074,In_98,In_960);
nor U2075 (N_2075,In_302,In_409);
nand U2076 (N_2076,In_756,In_376);
and U2077 (N_2077,In_442,In_504);
nor U2078 (N_2078,In_715,In_3);
nor U2079 (N_2079,In_42,In_598);
nand U2080 (N_2080,In_112,In_205);
and U2081 (N_2081,In_372,In_123);
or U2082 (N_2082,In_138,In_45);
nor U2083 (N_2083,In_555,In_382);
nand U2084 (N_2084,In_197,In_369);
nand U2085 (N_2085,In_868,In_953);
or U2086 (N_2086,In_767,In_510);
nor U2087 (N_2087,In_42,In_74);
nor U2088 (N_2088,In_144,In_619);
nand U2089 (N_2089,In_264,In_666);
nor U2090 (N_2090,In_593,In_222);
or U2091 (N_2091,In_827,In_801);
nand U2092 (N_2092,In_397,In_555);
nand U2093 (N_2093,In_764,In_378);
and U2094 (N_2094,In_568,In_47);
nor U2095 (N_2095,In_650,In_309);
or U2096 (N_2096,In_525,In_775);
nor U2097 (N_2097,In_242,In_299);
nand U2098 (N_2098,In_639,In_81);
xor U2099 (N_2099,In_500,In_800);
and U2100 (N_2100,In_485,In_476);
or U2101 (N_2101,In_967,In_358);
and U2102 (N_2102,In_116,In_27);
and U2103 (N_2103,In_744,In_672);
nor U2104 (N_2104,In_649,In_601);
nor U2105 (N_2105,In_286,In_206);
and U2106 (N_2106,In_376,In_571);
xnor U2107 (N_2107,In_270,In_176);
and U2108 (N_2108,In_994,In_98);
nand U2109 (N_2109,In_434,In_800);
nor U2110 (N_2110,In_269,In_607);
and U2111 (N_2111,In_437,In_409);
nand U2112 (N_2112,In_32,In_83);
and U2113 (N_2113,In_500,In_918);
and U2114 (N_2114,In_675,In_548);
and U2115 (N_2115,In_689,In_819);
and U2116 (N_2116,In_238,In_236);
and U2117 (N_2117,In_832,In_621);
nand U2118 (N_2118,In_153,In_149);
or U2119 (N_2119,In_906,In_699);
nand U2120 (N_2120,In_787,In_578);
nor U2121 (N_2121,In_359,In_834);
nand U2122 (N_2122,In_530,In_90);
or U2123 (N_2123,In_146,In_891);
nor U2124 (N_2124,In_256,In_796);
and U2125 (N_2125,In_629,In_751);
nand U2126 (N_2126,In_563,In_303);
nor U2127 (N_2127,In_863,In_146);
nor U2128 (N_2128,In_304,In_950);
nor U2129 (N_2129,In_469,In_13);
nand U2130 (N_2130,In_907,In_372);
or U2131 (N_2131,In_856,In_392);
and U2132 (N_2132,In_510,In_585);
nor U2133 (N_2133,In_119,In_445);
nor U2134 (N_2134,In_779,In_207);
nand U2135 (N_2135,In_814,In_650);
nand U2136 (N_2136,In_845,In_280);
and U2137 (N_2137,In_888,In_13);
nor U2138 (N_2138,In_160,In_365);
nor U2139 (N_2139,In_202,In_18);
and U2140 (N_2140,In_225,In_605);
nand U2141 (N_2141,In_833,In_48);
and U2142 (N_2142,In_804,In_316);
and U2143 (N_2143,In_580,In_329);
nor U2144 (N_2144,In_842,In_80);
nor U2145 (N_2145,In_179,In_453);
or U2146 (N_2146,In_109,In_68);
or U2147 (N_2147,In_411,In_970);
nor U2148 (N_2148,In_784,In_82);
nand U2149 (N_2149,In_345,In_14);
nor U2150 (N_2150,In_702,In_916);
nand U2151 (N_2151,In_558,In_222);
and U2152 (N_2152,In_941,In_732);
nand U2153 (N_2153,In_550,In_324);
nand U2154 (N_2154,In_785,In_578);
and U2155 (N_2155,In_440,In_811);
and U2156 (N_2156,In_132,In_333);
or U2157 (N_2157,In_902,In_105);
nand U2158 (N_2158,In_58,In_120);
nor U2159 (N_2159,In_700,In_307);
and U2160 (N_2160,In_16,In_417);
and U2161 (N_2161,In_642,In_924);
nand U2162 (N_2162,In_114,In_573);
nor U2163 (N_2163,In_566,In_337);
or U2164 (N_2164,In_277,In_8);
and U2165 (N_2165,In_615,In_218);
nor U2166 (N_2166,In_697,In_43);
or U2167 (N_2167,In_99,In_911);
and U2168 (N_2168,In_199,In_637);
or U2169 (N_2169,In_416,In_116);
and U2170 (N_2170,In_774,In_990);
nand U2171 (N_2171,In_742,In_146);
and U2172 (N_2172,In_306,In_807);
and U2173 (N_2173,In_772,In_368);
or U2174 (N_2174,In_7,In_231);
nor U2175 (N_2175,In_402,In_282);
nor U2176 (N_2176,In_383,In_88);
and U2177 (N_2177,In_38,In_853);
and U2178 (N_2178,In_897,In_376);
nand U2179 (N_2179,In_362,In_439);
and U2180 (N_2180,In_646,In_837);
nand U2181 (N_2181,In_658,In_358);
nand U2182 (N_2182,In_512,In_18);
or U2183 (N_2183,In_489,In_324);
and U2184 (N_2184,In_560,In_972);
nor U2185 (N_2185,In_53,In_144);
or U2186 (N_2186,In_44,In_936);
or U2187 (N_2187,In_779,In_991);
nor U2188 (N_2188,In_476,In_216);
or U2189 (N_2189,In_921,In_240);
nand U2190 (N_2190,In_183,In_199);
xor U2191 (N_2191,In_565,In_592);
nor U2192 (N_2192,In_506,In_647);
nor U2193 (N_2193,In_350,In_652);
nor U2194 (N_2194,In_79,In_94);
and U2195 (N_2195,In_309,In_587);
nand U2196 (N_2196,In_386,In_771);
nand U2197 (N_2197,In_775,In_253);
and U2198 (N_2198,In_851,In_663);
nor U2199 (N_2199,In_709,In_160);
nand U2200 (N_2200,In_26,In_684);
or U2201 (N_2201,In_729,In_524);
or U2202 (N_2202,In_233,In_410);
and U2203 (N_2203,In_587,In_84);
or U2204 (N_2204,In_491,In_893);
nor U2205 (N_2205,In_598,In_296);
and U2206 (N_2206,In_259,In_903);
or U2207 (N_2207,In_277,In_836);
and U2208 (N_2208,In_495,In_449);
and U2209 (N_2209,In_713,In_70);
and U2210 (N_2210,In_589,In_233);
and U2211 (N_2211,In_625,In_499);
and U2212 (N_2212,In_13,In_579);
and U2213 (N_2213,In_448,In_562);
nand U2214 (N_2214,In_395,In_790);
or U2215 (N_2215,In_666,In_842);
and U2216 (N_2216,In_734,In_149);
or U2217 (N_2217,In_288,In_488);
or U2218 (N_2218,In_967,In_248);
or U2219 (N_2219,In_215,In_532);
or U2220 (N_2220,In_61,In_724);
nand U2221 (N_2221,In_172,In_514);
nand U2222 (N_2222,In_284,In_359);
and U2223 (N_2223,In_738,In_158);
or U2224 (N_2224,In_828,In_816);
nand U2225 (N_2225,In_44,In_988);
and U2226 (N_2226,In_503,In_175);
nor U2227 (N_2227,In_627,In_181);
or U2228 (N_2228,In_500,In_491);
and U2229 (N_2229,In_618,In_677);
and U2230 (N_2230,In_458,In_300);
and U2231 (N_2231,In_972,In_977);
nand U2232 (N_2232,In_50,In_692);
nand U2233 (N_2233,In_826,In_254);
nand U2234 (N_2234,In_234,In_73);
and U2235 (N_2235,In_921,In_849);
xnor U2236 (N_2236,In_997,In_386);
nand U2237 (N_2237,In_511,In_2);
or U2238 (N_2238,In_119,In_147);
and U2239 (N_2239,In_888,In_884);
nor U2240 (N_2240,In_321,In_871);
nand U2241 (N_2241,In_776,In_535);
nor U2242 (N_2242,In_336,In_622);
xor U2243 (N_2243,In_581,In_436);
or U2244 (N_2244,In_78,In_308);
nor U2245 (N_2245,In_663,In_38);
and U2246 (N_2246,In_702,In_26);
nor U2247 (N_2247,In_527,In_287);
or U2248 (N_2248,In_460,In_75);
nor U2249 (N_2249,In_620,In_834);
nand U2250 (N_2250,In_149,In_925);
and U2251 (N_2251,In_138,In_486);
nand U2252 (N_2252,In_42,In_599);
nand U2253 (N_2253,In_795,In_886);
or U2254 (N_2254,In_144,In_532);
nand U2255 (N_2255,In_921,In_724);
and U2256 (N_2256,In_663,In_745);
nand U2257 (N_2257,In_498,In_563);
nor U2258 (N_2258,In_361,In_552);
nor U2259 (N_2259,In_898,In_682);
and U2260 (N_2260,In_741,In_932);
and U2261 (N_2261,In_472,In_247);
nor U2262 (N_2262,In_571,In_132);
nand U2263 (N_2263,In_683,In_618);
nand U2264 (N_2264,In_757,In_401);
or U2265 (N_2265,In_546,In_543);
nand U2266 (N_2266,In_370,In_321);
nor U2267 (N_2267,In_482,In_210);
and U2268 (N_2268,In_711,In_675);
or U2269 (N_2269,In_518,In_346);
and U2270 (N_2270,In_716,In_177);
nor U2271 (N_2271,In_953,In_348);
or U2272 (N_2272,In_727,In_832);
nand U2273 (N_2273,In_895,In_714);
nand U2274 (N_2274,In_427,In_20);
and U2275 (N_2275,In_997,In_510);
and U2276 (N_2276,In_900,In_701);
or U2277 (N_2277,In_724,In_555);
or U2278 (N_2278,In_189,In_242);
nor U2279 (N_2279,In_17,In_654);
or U2280 (N_2280,In_418,In_748);
or U2281 (N_2281,In_802,In_886);
or U2282 (N_2282,In_907,In_837);
nand U2283 (N_2283,In_100,In_82);
nor U2284 (N_2284,In_406,In_723);
or U2285 (N_2285,In_713,In_218);
and U2286 (N_2286,In_96,In_830);
and U2287 (N_2287,In_370,In_214);
or U2288 (N_2288,In_66,In_811);
or U2289 (N_2289,In_245,In_486);
nand U2290 (N_2290,In_912,In_311);
and U2291 (N_2291,In_767,In_986);
nor U2292 (N_2292,In_415,In_393);
nand U2293 (N_2293,In_786,In_337);
nand U2294 (N_2294,In_822,In_487);
nand U2295 (N_2295,In_631,In_691);
or U2296 (N_2296,In_685,In_119);
or U2297 (N_2297,In_262,In_219);
nand U2298 (N_2298,In_863,In_199);
nand U2299 (N_2299,In_578,In_151);
nand U2300 (N_2300,In_936,In_229);
nor U2301 (N_2301,In_307,In_698);
and U2302 (N_2302,In_150,In_652);
nor U2303 (N_2303,In_203,In_257);
and U2304 (N_2304,In_754,In_439);
nand U2305 (N_2305,In_533,In_126);
or U2306 (N_2306,In_378,In_561);
or U2307 (N_2307,In_829,In_418);
nor U2308 (N_2308,In_586,In_827);
nand U2309 (N_2309,In_412,In_907);
nand U2310 (N_2310,In_325,In_799);
nor U2311 (N_2311,In_948,In_531);
and U2312 (N_2312,In_282,In_767);
nor U2313 (N_2313,In_52,In_325);
nand U2314 (N_2314,In_654,In_809);
nand U2315 (N_2315,In_245,In_892);
and U2316 (N_2316,In_325,In_11);
and U2317 (N_2317,In_299,In_716);
and U2318 (N_2318,In_121,In_436);
and U2319 (N_2319,In_76,In_372);
or U2320 (N_2320,In_916,In_706);
nand U2321 (N_2321,In_72,In_637);
nand U2322 (N_2322,In_85,In_951);
or U2323 (N_2323,In_975,In_693);
or U2324 (N_2324,In_408,In_743);
nand U2325 (N_2325,In_199,In_567);
or U2326 (N_2326,In_917,In_869);
or U2327 (N_2327,In_268,In_440);
nand U2328 (N_2328,In_451,In_743);
nand U2329 (N_2329,In_272,In_67);
or U2330 (N_2330,In_563,In_648);
nor U2331 (N_2331,In_659,In_240);
nand U2332 (N_2332,In_262,In_104);
and U2333 (N_2333,In_502,In_962);
nor U2334 (N_2334,In_305,In_879);
and U2335 (N_2335,In_633,In_977);
or U2336 (N_2336,In_128,In_10);
and U2337 (N_2337,In_997,In_433);
or U2338 (N_2338,In_451,In_546);
or U2339 (N_2339,In_660,In_136);
nand U2340 (N_2340,In_736,In_745);
and U2341 (N_2341,In_439,In_572);
nand U2342 (N_2342,In_985,In_791);
and U2343 (N_2343,In_40,In_51);
or U2344 (N_2344,In_278,In_147);
and U2345 (N_2345,In_45,In_323);
or U2346 (N_2346,In_205,In_175);
nor U2347 (N_2347,In_636,In_930);
or U2348 (N_2348,In_500,In_548);
nor U2349 (N_2349,In_605,In_420);
and U2350 (N_2350,In_621,In_830);
nor U2351 (N_2351,In_367,In_284);
and U2352 (N_2352,In_503,In_681);
and U2353 (N_2353,In_141,In_96);
nand U2354 (N_2354,In_234,In_140);
nor U2355 (N_2355,In_263,In_132);
and U2356 (N_2356,In_561,In_711);
nor U2357 (N_2357,In_813,In_493);
and U2358 (N_2358,In_19,In_945);
nor U2359 (N_2359,In_9,In_648);
nand U2360 (N_2360,In_715,In_776);
or U2361 (N_2361,In_747,In_12);
nor U2362 (N_2362,In_534,In_987);
nor U2363 (N_2363,In_209,In_943);
nand U2364 (N_2364,In_163,In_762);
nor U2365 (N_2365,In_560,In_42);
or U2366 (N_2366,In_302,In_959);
or U2367 (N_2367,In_841,In_198);
or U2368 (N_2368,In_332,In_91);
nand U2369 (N_2369,In_900,In_658);
nor U2370 (N_2370,In_65,In_696);
or U2371 (N_2371,In_478,In_387);
or U2372 (N_2372,In_756,In_223);
or U2373 (N_2373,In_796,In_94);
nor U2374 (N_2374,In_877,In_987);
nand U2375 (N_2375,In_789,In_374);
and U2376 (N_2376,In_546,In_965);
and U2377 (N_2377,In_651,In_858);
nor U2378 (N_2378,In_958,In_997);
and U2379 (N_2379,In_943,In_813);
and U2380 (N_2380,In_19,In_412);
or U2381 (N_2381,In_49,In_806);
nand U2382 (N_2382,In_32,In_869);
and U2383 (N_2383,In_378,In_893);
nand U2384 (N_2384,In_200,In_771);
and U2385 (N_2385,In_461,In_281);
or U2386 (N_2386,In_501,In_315);
and U2387 (N_2387,In_471,In_721);
and U2388 (N_2388,In_856,In_184);
nand U2389 (N_2389,In_513,In_80);
nand U2390 (N_2390,In_405,In_984);
nor U2391 (N_2391,In_691,In_987);
or U2392 (N_2392,In_485,In_639);
or U2393 (N_2393,In_543,In_798);
or U2394 (N_2394,In_382,In_230);
nor U2395 (N_2395,In_650,In_437);
or U2396 (N_2396,In_150,In_163);
nor U2397 (N_2397,In_801,In_148);
or U2398 (N_2398,In_647,In_309);
and U2399 (N_2399,In_109,In_433);
nor U2400 (N_2400,In_71,In_149);
nor U2401 (N_2401,In_410,In_144);
or U2402 (N_2402,In_277,In_750);
and U2403 (N_2403,In_151,In_177);
nand U2404 (N_2404,In_708,In_324);
nand U2405 (N_2405,In_920,In_467);
nand U2406 (N_2406,In_571,In_193);
nor U2407 (N_2407,In_66,In_894);
or U2408 (N_2408,In_216,In_295);
or U2409 (N_2409,In_588,In_980);
nor U2410 (N_2410,In_938,In_612);
and U2411 (N_2411,In_620,In_524);
nor U2412 (N_2412,In_355,In_152);
or U2413 (N_2413,In_34,In_411);
nand U2414 (N_2414,In_645,In_378);
nor U2415 (N_2415,In_347,In_253);
and U2416 (N_2416,In_100,In_561);
or U2417 (N_2417,In_706,In_872);
xnor U2418 (N_2418,In_694,In_534);
nand U2419 (N_2419,In_574,In_758);
nor U2420 (N_2420,In_373,In_375);
and U2421 (N_2421,In_544,In_92);
nor U2422 (N_2422,In_15,In_755);
nor U2423 (N_2423,In_976,In_506);
and U2424 (N_2424,In_900,In_53);
nand U2425 (N_2425,In_366,In_397);
or U2426 (N_2426,In_608,In_405);
nor U2427 (N_2427,In_285,In_853);
nand U2428 (N_2428,In_700,In_181);
and U2429 (N_2429,In_962,In_418);
and U2430 (N_2430,In_590,In_365);
nand U2431 (N_2431,In_389,In_783);
and U2432 (N_2432,In_339,In_93);
nand U2433 (N_2433,In_810,In_115);
nor U2434 (N_2434,In_528,In_883);
or U2435 (N_2435,In_142,In_231);
xor U2436 (N_2436,In_436,In_606);
nor U2437 (N_2437,In_233,In_836);
nand U2438 (N_2438,In_552,In_255);
and U2439 (N_2439,In_587,In_211);
nand U2440 (N_2440,In_146,In_464);
nor U2441 (N_2441,In_345,In_714);
and U2442 (N_2442,In_628,In_735);
nand U2443 (N_2443,In_793,In_250);
nor U2444 (N_2444,In_762,In_552);
nand U2445 (N_2445,In_544,In_526);
nand U2446 (N_2446,In_328,In_519);
or U2447 (N_2447,In_840,In_908);
or U2448 (N_2448,In_672,In_14);
or U2449 (N_2449,In_300,In_74);
or U2450 (N_2450,In_170,In_747);
or U2451 (N_2451,In_934,In_669);
or U2452 (N_2452,In_793,In_361);
nor U2453 (N_2453,In_159,In_825);
nor U2454 (N_2454,In_933,In_503);
nand U2455 (N_2455,In_773,In_28);
or U2456 (N_2456,In_935,In_365);
nor U2457 (N_2457,In_474,In_955);
and U2458 (N_2458,In_582,In_765);
and U2459 (N_2459,In_397,In_169);
and U2460 (N_2460,In_733,In_196);
nand U2461 (N_2461,In_27,In_759);
or U2462 (N_2462,In_668,In_828);
nand U2463 (N_2463,In_596,In_508);
or U2464 (N_2464,In_169,In_334);
nand U2465 (N_2465,In_860,In_49);
nor U2466 (N_2466,In_835,In_81);
and U2467 (N_2467,In_235,In_38);
nor U2468 (N_2468,In_307,In_882);
nor U2469 (N_2469,In_62,In_22);
nand U2470 (N_2470,In_407,In_435);
nand U2471 (N_2471,In_571,In_507);
nand U2472 (N_2472,In_864,In_914);
and U2473 (N_2473,In_487,In_627);
nor U2474 (N_2474,In_349,In_586);
or U2475 (N_2475,In_80,In_525);
and U2476 (N_2476,In_737,In_323);
and U2477 (N_2477,In_385,In_370);
nor U2478 (N_2478,In_317,In_404);
nand U2479 (N_2479,In_561,In_987);
nor U2480 (N_2480,In_524,In_27);
nand U2481 (N_2481,In_613,In_9);
xnor U2482 (N_2482,In_696,In_402);
and U2483 (N_2483,In_91,In_768);
or U2484 (N_2484,In_59,In_930);
nand U2485 (N_2485,In_76,In_389);
and U2486 (N_2486,In_943,In_919);
nand U2487 (N_2487,In_147,In_209);
and U2488 (N_2488,In_390,In_481);
and U2489 (N_2489,In_581,In_602);
or U2490 (N_2490,In_130,In_944);
nor U2491 (N_2491,In_158,In_396);
nand U2492 (N_2492,In_413,In_32);
or U2493 (N_2493,In_122,In_895);
nand U2494 (N_2494,In_434,In_872);
nor U2495 (N_2495,In_482,In_212);
nand U2496 (N_2496,In_994,In_679);
nand U2497 (N_2497,In_765,In_677);
or U2498 (N_2498,In_700,In_33);
or U2499 (N_2499,In_229,In_544);
nor U2500 (N_2500,N_1470,N_880);
nor U2501 (N_2501,N_596,N_683);
nor U2502 (N_2502,N_1221,N_1859);
and U2503 (N_2503,N_2115,N_1002);
or U2504 (N_2504,N_415,N_360);
nor U2505 (N_2505,N_1566,N_2339);
or U2506 (N_2506,N_806,N_615);
nor U2507 (N_2507,N_1630,N_1706);
and U2508 (N_2508,N_1633,N_592);
and U2509 (N_2509,N_1372,N_514);
nor U2510 (N_2510,N_656,N_794);
nor U2511 (N_2511,N_1635,N_2237);
nor U2512 (N_2512,N_1933,N_758);
nor U2513 (N_2513,N_1342,N_1245);
nand U2514 (N_2514,N_525,N_2247);
nor U2515 (N_2515,N_1853,N_1409);
or U2516 (N_2516,N_1850,N_1541);
or U2517 (N_2517,N_561,N_608);
nand U2518 (N_2518,N_432,N_2417);
nor U2519 (N_2519,N_1425,N_646);
nand U2520 (N_2520,N_696,N_1291);
or U2521 (N_2521,N_1448,N_2252);
or U2522 (N_2522,N_776,N_1754);
nand U2523 (N_2523,N_850,N_1513);
or U2524 (N_2524,N_1436,N_649);
and U2525 (N_2525,N_326,N_1044);
nand U2526 (N_2526,N_2206,N_1921);
and U2527 (N_2527,N_1177,N_2432);
and U2528 (N_2528,N_1136,N_1900);
nand U2529 (N_2529,N_963,N_129);
nand U2530 (N_2530,N_1627,N_2126);
nand U2531 (N_2531,N_1621,N_185);
nand U2532 (N_2532,N_2134,N_2324);
and U2533 (N_2533,N_2446,N_1942);
nor U2534 (N_2534,N_1651,N_1550);
or U2535 (N_2535,N_372,N_1258);
or U2536 (N_2536,N_1060,N_32);
nor U2537 (N_2537,N_637,N_1306);
or U2538 (N_2538,N_429,N_290);
or U2539 (N_2539,N_737,N_945);
and U2540 (N_2540,N_1107,N_1368);
nand U2541 (N_2541,N_523,N_2371);
and U2542 (N_2542,N_417,N_252);
or U2543 (N_2543,N_1223,N_687);
or U2544 (N_2544,N_566,N_1288);
or U2545 (N_2545,N_887,N_2447);
or U2546 (N_2546,N_414,N_1776);
and U2547 (N_2547,N_1601,N_1901);
nor U2548 (N_2548,N_468,N_984);
nand U2549 (N_2549,N_807,N_1847);
nor U2550 (N_2550,N_507,N_1611);
or U2551 (N_2551,N_308,N_2210);
nor U2552 (N_2552,N_1255,N_426);
nor U2553 (N_2553,N_1990,N_2458);
nor U2554 (N_2554,N_855,N_1769);
nand U2555 (N_2555,N_184,N_146);
nand U2556 (N_2556,N_2168,N_1637);
and U2557 (N_2557,N_761,N_2166);
nand U2558 (N_2558,N_1095,N_438);
or U2559 (N_2559,N_2039,N_1344);
or U2560 (N_2560,N_1434,N_2125);
nor U2561 (N_2561,N_933,N_893);
xnor U2562 (N_2562,N_2144,N_227);
nor U2563 (N_2563,N_682,N_1093);
and U2564 (N_2564,N_2470,N_1388);
and U2565 (N_2565,N_851,N_2288);
or U2566 (N_2566,N_1832,N_1457);
and U2567 (N_2567,N_352,N_151);
and U2568 (N_2568,N_285,N_1313);
and U2569 (N_2569,N_1432,N_2120);
nor U2570 (N_2570,N_2194,N_1569);
or U2571 (N_2571,N_64,N_1035);
or U2572 (N_2572,N_2037,N_1539);
xor U2573 (N_2573,N_1906,N_1682);
nand U2574 (N_2574,N_375,N_313);
nor U2575 (N_2575,N_1262,N_344);
and U2576 (N_2576,N_228,N_2157);
nand U2577 (N_2577,N_469,N_1839);
nor U2578 (N_2578,N_1840,N_1760);
and U2579 (N_2579,N_1773,N_2379);
or U2580 (N_2580,N_1261,N_1994);
nand U2581 (N_2581,N_2251,N_1064);
nand U2582 (N_2582,N_741,N_467);
nand U2583 (N_2583,N_323,N_1155);
nand U2584 (N_2584,N_1399,N_1522);
nand U2585 (N_2585,N_2423,N_139);
nand U2586 (N_2586,N_991,N_2087);
or U2587 (N_2587,N_1753,N_2047);
nor U2588 (N_2588,N_1157,N_54);
nand U2589 (N_2589,N_401,N_2232);
and U2590 (N_2590,N_908,N_330);
or U2591 (N_2591,N_1881,N_424);
nor U2592 (N_2592,N_2071,N_1338);
nand U2593 (N_2593,N_1631,N_2114);
and U2594 (N_2594,N_2171,N_69);
and U2595 (N_2595,N_985,N_1251);
nor U2596 (N_2596,N_1384,N_1855);
and U2597 (N_2597,N_643,N_833);
and U2598 (N_2598,N_695,N_2351);
and U2599 (N_2599,N_2367,N_2113);
and U2600 (N_2600,N_1340,N_800);
and U2601 (N_2601,N_1632,N_1273);
xor U2602 (N_2602,N_818,N_445);
or U2603 (N_2603,N_759,N_1620);
and U2604 (N_2604,N_2053,N_2401);
nand U2605 (N_2605,N_977,N_1200);
or U2606 (N_2606,N_292,N_1961);
nor U2607 (N_2607,N_123,N_499);
nand U2608 (N_2608,N_2298,N_2045);
nand U2609 (N_2609,N_1722,N_2142);
or U2610 (N_2610,N_715,N_2170);
nand U2611 (N_2611,N_810,N_728);
nand U2612 (N_2612,N_2372,N_1312);
or U2613 (N_2613,N_1912,N_1424);
or U2614 (N_2614,N_2208,N_2133);
nand U2615 (N_2615,N_941,N_754);
nor U2616 (N_2616,N_358,N_200);
nand U2617 (N_2617,N_1700,N_2286);
and U2618 (N_2618,N_1130,N_922);
or U2619 (N_2619,N_2487,N_1973);
nand U2620 (N_2620,N_2436,N_2414);
nor U2621 (N_2621,N_2050,N_1995);
nand U2622 (N_2622,N_1898,N_942);
nand U2623 (N_2623,N_760,N_116);
nor U2624 (N_2624,N_1547,N_973);
and U2625 (N_2625,N_1718,N_1579);
or U2626 (N_2626,N_341,N_780);
nand U2627 (N_2627,N_466,N_2409);
nor U2628 (N_2628,N_1201,N_1336);
nor U2629 (N_2629,N_168,N_273);
nor U2630 (N_2630,N_678,N_988);
or U2631 (N_2631,N_1693,N_726);
or U2632 (N_2632,N_164,N_2433);
xor U2633 (N_2633,N_1816,N_1887);
nor U2634 (N_2634,N_1226,N_2069);
nor U2635 (N_2635,N_2457,N_791);
nand U2636 (N_2636,N_774,N_1979);
and U2637 (N_2637,N_1624,N_1841);
and U2638 (N_2638,N_2364,N_1894);
or U2639 (N_2639,N_1787,N_822);
nand U2640 (N_2640,N_2308,N_1305);
nand U2641 (N_2641,N_700,N_1061);
nor U2642 (N_2642,N_2280,N_316);
or U2643 (N_2643,N_1899,N_713);
nor U2644 (N_2644,N_1439,N_1561);
or U2645 (N_2645,N_419,N_881);
nand U2646 (N_2646,N_2389,N_271);
and U2647 (N_2647,N_1355,N_2257);
nor U2648 (N_2648,N_1999,N_1199);
nor U2649 (N_2649,N_1751,N_2192);
or U2650 (N_2650,N_957,N_845);
nand U2651 (N_2651,N_958,N_298);
and U2652 (N_2652,N_2240,N_2112);
nand U2653 (N_2653,N_2305,N_2346);
or U2654 (N_2654,N_1167,N_2195);
nor U2655 (N_2655,N_1966,N_1366);
nand U2656 (N_2656,N_2107,N_543);
nand U2657 (N_2657,N_2416,N_910);
nand U2658 (N_2658,N_2201,N_755);
or U2659 (N_2659,N_1389,N_42);
nor U2660 (N_2660,N_1408,N_1230);
and U2661 (N_2661,N_2466,N_2493);
nor U2662 (N_2662,N_581,N_837);
and U2663 (N_2663,N_98,N_2062);
or U2664 (N_2664,N_510,N_877);
or U2665 (N_2665,N_1799,N_256);
nor U2666 (N_2666,N_422,N_1863);
nand U2667 (N_2667,N_2478,N_2336);
and U2668 (N_2668,N_1535,N_1676);
and U2669 (N_2669,N_627,N_2083);
or U2670 (N_2670,N_1852,N_1510);
or U2671 (N_2671,N_1247,N_296);
or U2672 (N_2672,N_1458,N_137);
or U2673 (N_2673,N_2182,N_399);
and U2674 (N_2674,N_707,N_11);
and U2675 (N_2675,N_2400,N_1952);
nor U2676 (N_2676,N_165,N_593);
and U2677 (N_2677,N_1810,N_2078);
or U2678 (N_2678,N_2174,N_1928);
and U2679 (N_2679,N_1178,N_2321);
and U2680 (N_2680,N_1211,N_504);
or U2681 (N_2681,N_1750,N_412);
nor U2682 (N_2682,N_1166,N_1087);
nand U2683 (N_2683,N_584,N_288);
nor U2684 (N_2684,N_757,N_2186);
nand U2685 (N_2685,N_1075,N_1654);
and U2686 (N_2686,N_269,N_2329);
or U2687 (N_2687,N_744,N_1652);
and U2688 (N_2688,N_2405,N_2393);
nor U2689 (N_2689,N_1484,N_975);
or U2690 (N_2690,N_1345,N_1517);
or U2691 (N_2691,N_530,N_478);
or U2692 (N_2692,N_586,N_1820);
and U2693 (N_2693,N_2334,N_2007);
or U2694 (N_2694,N_2220,N_1565);
and U2695 (N_2695,N_178,N_2026);
or U2696 (N_2696,N_127,N_953);
or U2697 (N_2697,N_1934,N_1016);
or U2698 (N_2698,N_1743,N_1828);
and U2699 (N_2699,N_1604,N_740);
or U2700 (N_2700,N_1804,N_2193);
nand U2701 (N_2701,N_1055,N_2070);
nor U2702 (N_2702,N_1057,N_639);
nand U2703 (N_2703,N_1024,N_2185);
nand U2704 (N_2704,N_311,N_2154);
or U2705 (N_2705,N_2332,N_2046);
nor U2706 (N_2706,N_206,N_12);
or U2707 (N_2707,N_1260,N_1465);
or U2708 (N_2708,N_2385,N_1418);
and U2709 (N_2709,N_411,N_2230);
nand U2710 (N_2710,N_1814,N_8);
nand U2711 (N_2711,N_669,N_2061);
nor U2712 (N_2712,N_2451,N_1834);
nand U2713 (N_2713,N_1378,N_1354);
nand U2714 (N_2714,N_915,N_657);
nor U2715 (N_2715,N_551,N_84);
and U2716 (N_2716,N_1556,N_1655);
or U2717 (N_2717,N_2277,N_274);
nand U2718 (N_2718,N_240,N_152);
or U2719 (N_2719,N_2213,N_970);
or U2720 (N_2720,N_1501,N_578);
and U2721 (N_2721,N_2052,N_663);
nor U2722 (N_2722,N_31,N_948);
nand U2723 (N_2723,N_1189,N_932);
nand U2724 (N_2724,N_1032,N_2236);
or U2725 (N_2725,N_2076,N_94);
or U2726 (N_2726,N_1334,N_1460);
and U2727 (N_2727,N_1642,N_378);
nor U2728 (N_2728,N_1842,N_2179);
nor U2729 (N_2729,N_1381,N_66);
nor U2730 (N_2730,N_1739,N_1913);
nand U2731 (N_2731,N_1697,N_36);
nor U2732 (N_2732,N_2489,N_2307);
nor U2733 (N_2733,N_1857,N_1412);
nor U2734 (N_2734,N_1735,N_1516);
nand U2735 (N_2735,N_1416,N_1640);
or U2736 (N_2736,N_1709,N_2108);
nor U2737 (N_2737,N_795,N_2456);
nand U2738 (N_2738,N_2381,N_1451);
xor U2739 (N_2739,N_380,N_1647);
nor U2740 (N_2740,N_2119,N_2323);
and U2741 (N_2741,N_2234,N_1151);
or U2742 (N_2742,N_475,N_331);
nand U2743 (N_2743,N_2435,N_729);
nor U2744 (N_2744,N_706,N_2420);
nor U2745 (N_2745,N_1085,N_1259);
and U2746 (N_2746,N_710,N_1858);
and U2747 (N_2747,N_453,N_2003);
nor U2748 (N_2748,N_1573,N_2290);
nand U2749 (N_2749,N_470,N_1008);
or U2750 (N_2750,N_1673,N_490);
or U2751 (N_2751,N_2072,N_1475);
and U2752 (N_2752,N_1675,N_620);
nand U2753 (N_2753,N_1925,N_1321);
or U2754 (N_2754,N_1158,N_1626);
and U2755 (N_2755,N_310,N_2049);
and U2756 (N_2756,N_340,N_752);
and U2757 (N_2757,N_193,N_978);
nor U2758 (N_2758,N_383,N_1184);
nor U2759 (N_2759,N_1781,N_2105);
or U2760 (N_2760,N_1586,N_121);
or U2761 (N_2761,N_2127,N_690);
or U2762 (N_2762,N_1919,N_542);
nand U2763 (N_2763,N_1920,N_1872);
or U2764 (N_2764,N_2143,N_1555);
nand U2765 (N_2765,N_2136,N_2441);
and U2766 (N_2766,N_2101,N_1891);
nand U2767 (N_2767,N_1109,N_763);
nor U2768 (N_2768,N_1698,N_1144);
or U2769 (N_2769,N_633,N_1888);
and U2770 (N_2770,N_398,N_2445);
nor U2771 (N_2771,N_559,N_2139);
and U2772 (N_2772,N_346,N_109);
and U2773 (N_2773,N_314,N_265);
nor U2774 (N_2774,N_161,N_1171);
nor U2775 (N_2775,N_1512,N_2454);
nor U2776 (N_2776,N_1037,N_1011);
and U2777 (N_2777,N_1974,N_659);
or U2778 (N_2778,N_405,N_2248);
or U2779 (N_2779,N_2394,N_205);
nand U2780 (N_2780,N_348,N_1975);
nand U2781 (N_2781,N_911,N_2282);
and U2782 (N_2782,N_1352,N_2468);
nand U2783 (N_2783,N_1600,N_1134);
or U2784 (N_2784,N_2088,N_374);
nand U2785 (N_2785,N_1643,N_2057);
nor U2786 (N_2786,N_270,N_1712);
nand U2787 (N_2787,N_799,N_2162);
nor U2788 (N_2788,N_935,N_1431);
xnor U2789 (N_2789,N_1217,N_1433);
nor U2790 (N_2790,N_1756,N_521);
nand U2791 (N_2791,N_2431,N_1492);
nand U2792 (N_2792,N_212,N_483);
xnor U2793 (N_2793,N_2268,N_1065);
nand U2794 (N_2794,N_1279,N_1013);
and U2795 (N_2795,N_250,N_1227);
nor U2796 (N_2796,N_2304,N_1455);
nor U2797 (N_2797,N_128,N_106);
and U2798 (N_2798,N_2359,N_1935);
nand U2799 (N_2799,N_838,N_1534);
nor U2800 (N_2800,N_105,N_730);
and U2801 (N_2801,N_2411,N_76);
or U2802 (N_2802,N_937,N_81);
nand U2803 (N_2803,N_1968,N_2130);
or U2804 (N_2804,N_1194,N_1792);
and U2805 (N_2805,N_1536,N_1530);
nor U2806 (N_2806,N_177,N_766);
or U2807 (N_2807,N_709,N_1932);
nand U2808 (N_2808,N_955,N_1580);
nand U2809 (N_2809,N_1719,N_2422);
or U2810 (N_2810,N_1128,N_1613);
nor U2811 (N_2811,N_772,N_225);
and U2812 (N_2812,N_428,N_1304);
nor U2813 (N_2813,N_243,N_1821);
nand U2814 (N_2814,N_1477,N_1489);
nor U2815 (N_2815,N_267,N_2345);
nand U2816 (N_2816,N_1328,N_2205);
nand U2817 (N_2817,N_808,N_80);
nand U2818 (N_2818,N_907,N_986);
or U2819 (N_2819,N_1940,N_2328);
or U2820 (N_2820,N_1165,N_110);
nand U2821 (N_2821,N_2019,N_1490);
nand U2822 (N_2822,N_904,N_1319);
nand U2823 (N_2823,N_2073,N_319);
or U2824 (N_2824,N_1361,N_1656);
and U2825 (N_2825,N_1951,N_291);
nor U2826 (N_2826,N_384,N_18);
or U2827 (N_2827,N_1474,N_2102);
nor U2828 (N_2828,N_1190,N_2137);
nor U2829 (N_2829,N_1950,N_2342);
and U2830 (N_2830,N_1007,N_1082);
nand U2831 (N_2831,N_1339,N_498);
nand U2832 (N_2832,N_482,N_644);
or U2833 (N_2833,N_1081,N_173);
or U2834 (N_2834,N_1377,N_1915);
and U2835 (N_2835,N_2473,N_343);
or U2836 (N_2836,N_2044,N_1337);
nor U2837 (N_2837,N_2480,N_617);
nand U2838 (N_2838,N_527,N_1977);
nand U2839 (N_2839,N_430,N_2249);
and U2840 (N_2840,N_373,N_1263);
nand U2841 (N_2841,N_1498,N_1195);
nand U2842 (N_2842,N_1004,N_2094);
or U2843 (N_2843,N_2153,N_59);
or U2844 (N_2844,N_847,N_815);
nand U2845 (N_2845,N_437,N_183);
nand U2846 (N_2846,N_1317,N_816);
xnor U2847 (N_2847,N_2318,N_88);
or U2848 (N_2848,N_732,N_1998);
and U2849 (N_2849,N_1202,N_436);
or U2850 (N_2850,N_1599,N_1419);
xor U2851 (N_2851,N_480,N_2055);
or U2852 (N_2852,N_361,N_1404);
or U2853 (N_2853,N_2375,N_2481);
or U2854 (N_2854,N_149,N_2449);
nand U2855 (N_2855,N_117,N_255);
and U2856 (N_2856,N_145,N_2207);
and U2857 (N_2857,N_1,N_2419);
or U2858 (N_2858,N_1967,N_1825);
nor U2859 (N_2859,N_156,N_2299);
nor U2860 (N_2860,N_2337,N_875);
nand U2861 (N_2861,N_964,N_1143);
nor U2862 (N_2862,N_1567,N_1428);
and U2863 (N_2863,N_2164,N_2273);
and U2864 (N_2864,N_2149,N_2098);
nand U2865 (N_2865,N_1575,N_829);
or U2866 (N_2866,N_2455,N_1023);
and U2867 (N_2867,N_443,N_92);
or U2868 (N_2868,N_1022,N_503);
nor U2869 (N_2869,N_1716,N_863);
nand U2870 (N_2870,N_2148,N_2175);
and U2871 (N_2871,N_871,N_1156);
or U2872 (N_2872,N_278,N_1710);
or U2873 (N_2873,N_70,N_1333);
nor U2874 (N_2874,N_990,N_387);
nand U2875 (N_2875,N_2437,N_2250);
nand U2876 (N_2876,N_1971,N_1614);
nand U2877 (N_2877,N_1976,N_2218);
nor U2878 (N_2878,N_2460,N_281);
and U2879 (N_2879,N_1954,N_823);
nand U2880 (N_2880,N_1382,N_1964);
and U2881 (N_2881,N_1066,N_1910);
nand U2882 (N_2882,N_1854,N_824);
nand U2883 (N_2883,N_2110,N_2368);
or U2884 (N_2884,N_148,N_679);
nand U2885 (N_2885,N_572,N_366);
nand U2886 (N_2886,N_1272,N_2089);
or U2887 (N_2887,N_517,N_1192);
or U2888 (N_2888,N_1789,N_724);
and U2889 (N_2889,N_464,N_747);
nor U2890 (N_2890,N_175,N_300);
and U2891 (N_2891,N_2264,N_2227);
or U2892 (N_2892,N_51,N_781);
nor U2893 (N_2893,N_841,N_355);
and U2894 (N_2894,N_2172,N_951);
nor U2895 (N_2895,N_996,N_321);
nand U2896 (N_2896,N_1407,N_886);
or U2897 (N_2897,N_1268,N_956);
or U2898 (N_2898,N_1274,N_1672);
or U2899 (N_2899,N_364,N_1746);
nand U2900 (N_2900,N_368,N_144);
or U2901 (N_2901,N_681,N_2129);
nand U2902 (N_2902,N_1692,N_925);
and U2903 (N_2903,N_632,N_1824);
nand U2904 (N_2904,N_1286,N_618);
and U2905 (N_2905,N_869,N_28);
and U2906 (N_2906,N_122,N_789);
or U2907 (N_2907,N_556,N_1509);
or U2908 (N_2908,N_512,N_2353);
or U2909 (N_2909,N_1362,N_86);
or U2910 (N_2910,N_749,N_2322);
and U2911 (N_2911,N_1807,N_260);
nor U2912 (N_2912,N_1256,N_1838);
nor U2913 (N_2913,N_2283,N_585);
nand U2914 (N_2914,N_397,N_1752);
nor U2915 (N_2915,N_1882,N_1936);
nor U2916 (N_2916,N_1105,N_753);
nand U2917 (N_2917,N_2074,N_1401);
nand U2918 (N_2918,N_1027,N_55);
or U2919 (N_2919,N_718,N_1603);
nand U2920 (N_2920,N_2256,N_1727);
nand U2921 (N_2921,N_236,N_1861);
or U2922 (N_2922,N_2067,N_2279);
or U2923 (N_2923,N_1941,N_554);
nand U2924 (N_2924,N_242,N_897);
and U2925 (N_2925,N_1294,N_1644);
nor U2926 (N_2926,N_22,N_1320);
and U2927 (N_2927,N_967,N_1802);
nand U2928 (N_2928,N_2147,N_961);
xor U2929 (N_2929,N_135,N_809);
nand U2930 (N_2930,N_976,N_2386);
or U2931 (N_2931,N_1815,N_111);
nor U2932 (N_2932,N_712,N_1996);
and U2933 (N_2933,N_2326,N_2199);
and U2934 (N_2934,N_1042,N_1454);
or U2935 (N_2935,N_882,N_141);
and U2936 (N_2936,N_702,N_1257);
nor U2937 (N_2937,N_1949,N_1552);
and U2938 (N_2938,N_15,N_392);
nor U2939 (N_2939,N_1285,N_811);
nor U2940 (N_2940,N_2335,N_251);
nor U2941 (N_2941,N_1759,N_1531);
nor U2942 (N_2942,N_1187,N_153);
nand U2943 (N_2943,N_1302,N_287);
or U2944 (N_2944,N_409,N_529);
or U2945 (N_2945,N_2428,N_2358);
nor U2946 (N_2946,N_1559,N_1124);
or U2947 (N_2947,N_376,N_134);
and U2948 (N_2948,N_1323,N_1736);
and U2949 (N_2949,N_458,N_934);
and U2950 (N_2950,N_1266,N_686);
nand U2951 (N_2951,N_2010,N_1026);
nand U2952 (N_2952,N_2284,N_474);
and U2953 (N_2953,N_2032,N_2302);
and U2954 (N_2954,N_21,N_697);
nor U2955 (N_2955,N_1080,N_1058);
or U2956 (N_2956,N_677,N_2035);
nand U2957 (N_2957,N_187,N_812);
or U2958 (N_2958,N_1835,N_1937);
nor U2959 (N_2959,N_2095,N_565);
or U2960 (N_2960,N_1734,N_1186);
nand U2961 (N_2961,N_1957,N_1958);
or U2962 (N_2962,N_1768,N_1708);
nor U2963 (N_2963,N_295,N_2278);
or U2964 (N_2964,N_68,N_692);
and U2965 (N_2965,N_2382,N_16);
nor U2966 (N_2966,N_1593,N_1707);
or U2967 (N_2967,N_1390,N_614);
or U2968 (N_2968,N_580,N_96);
and U2969 (N_2969,N_112,N_701);
or U2970 (N_2970,N_853,N_2293);
nand U2971 (N_2971,N_1182,N_2140);
nand U2972 (N_2972,N_719,N_1083);
nor U2973 (N_2973,N_2012,N_2287);
or U2974 (N_2974,N_406,N_67);
nor U2975 (N_2975,N_1036,N_485);
or U2976 (N_2976,N_539,N_1907);
nor U2977 (N_2977,N_1529,N_805);
or U2978 (N_2978,N_320,N_1984);
nand U2979 (N_2979,N_418,N_777);
nand U2980 (N_2980,N_1293,N_1717);
nor U2981 (N_2981,N_35,N_2016);
nor U2982 (N_2982,N_38,N_2384);
nand U2983 (N_2983,N_1846,N_492);
and U2984 (N_2984,N_447,N_782);
nor U2985 (N_2985,N_1574,N_1544);
nand U2986 (N_2986,N_13,N_545);
nand U2987 (N_2987,N_377,N_506);
xor U2988 (N_2988,N_20,N_2306);
nand U2989 (N_2989,N_1356,N_1125);
nand U2990 (N_2990,N_1959,N_1496);
nor U2991 (N_2991,N_1373,N_1346);
nor U2992 (N_2992,N_17,N_1406);
and U2993 (N_2993,N_1745,N_58);
and U2994 (N_2994,N_2292,N_2097);
and U2995 (N_2995,N_515,N_1594);
and U2996 (N_2996,N_1123,N_393);
and U2997 (N_2997,N_1299,N_1507);
nor U2998 (N_2998,N_2459,N_655);
and U2999 (N_2999,N_540,N_921);
or U3000 (N_3000,N_1092,N_524);
nand U3001 (N_3001,N_247,N_1325);
or U3002 (N_3002,N_722,N_1122);
and U3003 (N_3003,N_1622,N_1473);
or U3004 (N_3004,N_1733,N_1141);
and U3005 (N_3005,N_1231,N_2155);
and U3006 (N_3006,N_1153,N_1056);
or U3007 (N_3007,N_2009,N_1191);
nand U3008 (N_3008,N_1548,N_1918);
and U3009 (N_3009,N_47,N_1343);
or U3010 (N_3010,N_2316,N_979);
or U3011 (N_3011,N_797,N_983);
and U3012 (N_3012,N_2091,N_528);
nor U3013 (N_3013,N_1062,N_1193);
and U3014 (N_3014,N_2398,N_1364);
nand U3015 (N_3015,N_335,N_2015);
nor U3016 (N_3016,N_629,N_2141);
and U3017 (N_3017,N_1472,N_557);
nor U3018 (N_3018,N_263,N_302);
and U3019 (N_3019,N_159,N_2439);
nand U3020 (N_3020,N_1238,N_1324);
nor U3021 (N_3021,N_1909,N_929);
nor U3022 (N_3022,N_1445,N_1000);
nor U3023 (N_3023,N_234,N_1363);
nand U3024 (N_3024,N_1243,N_1437);
and U3025 (N_3025,N_1376,N_303);
nand U3026 (N_3026,N_1878,N_2497);
nand U3027 (N_3027,N_1545,N_667);
nor U3028 (N_3028,N_773,N_1916);
nor U3029 (N_3029,N_1091,N_820);
or U3030 (N_3030,N_2357,N_1006);
nor U3031 (N_3031,N_1890,N_1265);
nor U3032 (N_3032,N_1283,N_79);
nor U3033 (N_3033,N_1782,N_119);
and U3034 (N_3034,N_658,N_2158);
nand U3035 (N_3035,N_1711,N_1904);
nand U3036 (N_3036,N_938,N_2320);
nor U3037 (N_3037,N_2221,N_56);
nor U3038 (N_3038,N_1298,N_2294);
nor U3039 (N_3039,N_1870,N_1102);
and U3040 (N_3040,N_583,N_1054);
and U3041 (N_3041,N_714,N_2151);
or U3042 (N_3042,N_2370,N_564);
nor U3043 (N_3043,N_75,N_1468);
nor U3044 (N_3044,N_531,N_261);
or U3045 (N_3045,N_708,N_981);
and U3046 (N_3046,N_878,N_1084);
nand U3047 (N_3047,N_1664,N_2259);
and U3048 (N_3048,N_1738,N_218);
and U3049 (N_3049,N_1737,N_1301);
nor U3050 (N_3050,N_2356,N_1677);
or U3051 (N_3051,N_885,N_2027);
nor U3052 (N_3052,N_2059,N_1755);
nand U3053 (N_3053,N_1980,N_1089);
nor U3054 (N_3054,N_1139,N_1237);
and U3055 (N_3055,N_1253,N_2116);
and U3056 (N_3056,N_1370,N_2024);
and U3057 (N_3057,N_1371,N_1715);
nor U3058 (N_3058,N_913,N_1459);
and U3059 (N_3059,N_2412,N_2387);
or U3060 (N_3060,N_591,N_231);
or U3061 (N_3061,N_1583,N_1653);
nand U3062 (N_3062,N_1827,N_989);
nor U3063 (N_3063,N_1220,N_635);
or U3064 (N_3064,N_1557,N_10);
nand U3065 (N_3065,N_662,N_1188);
nor U3066 (N_3066,N_1449,N_1943);
nor U3067 (N_3067,N_420,N_2029);
and U3068 (N_3068,N_385,N_1309);
nor U3069 (N_3069,N_860,N_2163);
nand U3070 (N_3070,N_155,N_2404);
and U3071 (N_3071,N_739,N_790);
nand U3072 (N_3072,N_237,N_693);
and U3073 (N_3073,N_338,N_721);
nand U3074 (N_3074,N_2092,N_534);
nand U3075 (N_3075,N_1300,N_125);
or U3076 (N_3076,N_1772,N_1246);
or U3077 (N_3077,N_1350,N_731);
nor U3078 (N_3078,N_1533,N_1369);
or U3079 (N_3079,N_2080,N_421);
or U3080 (N_3080,N_1040,N_1052);
nand U3081 (N_3081,N_381,N_920);
nand U3082 (N_3082,N_2225,N_2377);
and U3083 (N_3083,N_751,N_456);
and U3084 (N_3084,N_204,N_391);
or U3085 (N_3085,N_1387,N_74);
nor U3086 (N_3086,N_917,N_2060);
or U3087 (N_3087,N_1775,N_1025);
nand U3088 (N_3088,N_2469,N_214);
nor U3089 (N_3089,N_7,N_2281);
or U3090 (N_3090,N_1795,N_1248);
or U3091 (N_3091,N_1161,N_2025);
or U3092 (N_3092,N_1380,N_1646);
nor U3093 (N_3093,N_997,N_2109);
and U3094 (N_3094,N_560,N_1689);
nand U3095 (N_3095,N_971,N_1028);
or U3096 (N_3096,N_410,N_1741);
and U3097 (N_3097,N_1017,N_2418);
or U3098 (N_3098,N_1744,N_2106);
nand U3099 (N_3099,N_1314,N_2467);
nor U3100 (N_3100,N_579,N_2442);
nand U3101 (N_3101,N_334,N_1069);
and U3102 (N_3102,N_1868,N_2319);
and U3103 (N_3103,N_587,N_258);
nor U3104 (N_3104,N_1502,N_1822);
nor U3105 (N_3105,N_661,N_1796);
nor U3106 (N_3106,N_500,N_1596);
nor U3107 (N_3107,N_1790,N_217);
nand U3108 (N_3108,N_213,N_85);
and U3109 (N_3109,N_1045,N_1794);
nor U3110 (N_3110,N_336,N_2471);
nor U3111 (N_3111,N_2312,N_2224);
nor U3112 (N_3112,N_1528,N_440);
nand U3113 (N_3113,N_1578,N_1880);
nand U3114 (N_3114,N_750,N_93);
nand U3115 (N_3115,N_625,N_1405);
or U3116 (N_3116,N_1665,N_268);
xnor U3117 (N_3117,N_1121,N_1059);
nor U3118 (N_3118,N_793,N_2380);
nor U3119 (N_3119,N_526,N_345);
and U3120 (N_3120,N_457,N_407);
or U3121 (N_3121,N_402,N_416);
or U3122 (N_3122,N_1871,N_2464);
nor U3123 (N_3123,N_1546,N_1926);
xnor U3124 (N_3124,N_648,N_1831);
nand U3125 (N_3125,N_450,N_2313);
nand U3126 (N_3126,N_1104,N_1033);
nor U3127 (N_3127,N_645,N_1931);
or U3128 (N_3128,N_2369,N_143);
and U3129 (N_3129,N_1577,N_1290);
nand U3130 (N_3130,N_1411,N_1721);
and U3131 (N_3131,N_1292,N_317);
and U3132 (N_3132,N_1978,N_454);
nand U3133 (N_3133,N_1420,N_1953);
nor U3134 (N_3134,N_1303,N_2267);
nor U3135 (N_3135,N_2219,N_1020);
or U3136 (N_3136,N_849,N_779);
and U3137 (N_3137,N_1829,N_2450);
nand U3138 (N_3138,N_209,N_1591);
and U3139 (N_3139,N_1427,N_2014);
or U3140 (N_3140,N_198,N_1705);
nand U3141 (N_3141,N_2474,N_1435);
or U3142 (N_3142,N_2241,N_1280);
nand U3143 (N_3143,N_65,N_181);
and U3144 (N_3144,N_489,N_2397);
or U3145 (N_3145,N_1679,N_2344);
and U3146 (N_3146,N_1295,N_1275);
and U3147 (N_3147,N_1763,N_1562);
nor U3148 (N_3148,N_1009,N_1176);
or U3149 (N_3149,N_2486,N_2479);
nor U3150 (N_3150,N_166,N_1170);
nand U3151 (N_3151,N_704,N_974);
nor U3152 (N_3152,N_2269,N_286);
or U3153 (N_3153,N_1780,N_960);
nand U3154 (N_3154,N_1267,N_832);
and U3155 (N_3155,N_817,N_1851);
nor U3156 (N_3156,N_1917,N_1740);
or U3157 (N_3157,N_202,N_0);
nor U3158 (N_3158,N_1695,N_864);
nor U3159 (N_3159,N_1638,N_2233);
and U3160 (N_3160,N_670,N_1173);
and U3161 (N_3161,N_481,N_2254);
or U3162 (N_3162,N_299,N_2407);
nand U3163 (N_3163,N_1276,N_1330);
and U3164 (N_3164,N_115,N_1658);
and U3165 (N_3165,N_778,N_257);
nand U3166 (N_3166,N_1726,N_1168);
nor U3167 (N_3167,N_668,N_1786);
nor U3168 (N_3168,N_1844,N_1197);
nand U3169 (N_3169,N_768,N_1674);
and U3170 (N_3170,N_611,N_1284);
or U3171 (N_3171,N_322,N_2427);
or U3172 (N_3172,N_1228,N_1965);
nor U3173 (N_3173,N_612,N_189);
nor U3174 (N_3174,N_353,N_705);
or U3175 (N_3175,N_2002,N_488);
or U3176 (N_3176,N_2034,N_1848);
nand U3177 (N_3177,N_473,N_223);
nor U3178 (N_3178,N_196,N_1239);
nand U3179 (N_3179,N_1823,N_546);
or U3180 (N_3180,N_2383,N_1902);
and U3181 (N_3181,N_2231,N_2348);
and U3182 (N_3182,N_840,N_673);
nand U3183 (N_3183,N_1359,N_276);
nor U3184 (N_3184,N_2476,N_462);
and U3185 (N_3185,N_1494,N_2352);
nor U3186 (N_3186,N_497,N_1793);
and U3187 (N_3187,N_444,N_1930);
nand U3188 (N_3188,N_2462,N_2217);
nand U3189 (N_3189,N_1270,N_26);
nand U3190 (N_3190,N_902,N_289);
nor U3191 (N_3191,N_1108,N_866);
nor U3192 (N_3192,N_1703,N_472);
or U3193 (N_3193,N_699,N_1504);
nand U3194 (N_3194,N_2465,N_771);
and U3195 (N_3195,N_2295,N_157);
nor U3196 (N_3196,N_1254,N_1609);
nor U3197 (N_3197,N_2311,N_1518);
nand U3198 (N_3198,N_1924,N_1415);
or U3199 (N_3199,N_1410,N_44);
and U3200 (N_3200,N_1985,N_224);
nor U3201 (N_3201,N_2424,N_2178);
nand U3202 (N_3202,N_2363,N_275);
or U3203 (N_3203,N_1969,N_2330);
and U3204 (N_3204,N_2238,N_2085);
nor U3205 (N_3205,N_1956,N_1118);
nor U3206 (N_3206,N_362,N_1154);
nor U3207 (N_3207,N_1629,N_2160);
nand U3208 (N_3208,N_1777,N_2146);
and U3209 (N_3209,N_2243,N_918);
or U3210 (N_3210,N_1224,N_896);
or U3211 (N_3211,N_1113,N_1450);
nand U3212 (N_3212,N_404,N_1204);
and U3213 (N_3213,N_315,N_1766);
or U3214 (N_3214,N_1101,N_104);
nor U3215 (N_3215,N_52,N_2017);
or U3216 (N_3216,N_626,N_91);
or U3217 (N_3217,N_203,N_1225);
nand U3218 (N_3218,N_1172,N_1469);
nand U3219 (N_3219,N_854,N_954);
nor U3220 (N_3220,N_1648,N_2421);
xor U3221 (N_3221,N_952,N_827);
nor U3222 (N_3222,N_1694,N_1132);
nor U3223 (N_3223,N_1873,N_282);
nor U3224 (N_3224,N_2434,N_2122);
or U3225 (N_3225,N_1791,N_1568);
nand U3226 (N_3226,N_1866,N_558);
nor U3227 (N_3227,N_1955,N_238);
or U3228 (N_3228,N_1463,N_1326);
and U3229 (N_3229,N_2461,N_2096);
nand U3230 (N_3230,N_37,N_516);
nand U3231 (N_3231,N_2075,N_927);
nand U3232 (N_3232,N_118,N_1068);
or U3233 (N_3233,N_1869,N_1576);
and U3234 (N_3234,N_494,N_982);
nand U3235 (N_3235,N_1413,N_1402);
nor U3236 (N_3236,N_2338,N_995);
and U3237 (N_3237,N_870,N_154);
and U3238 (N_3238,N_2190,N_1482);
or U3239 (N_3239,N_171,N_1488);
and U3240 (N_3240,N_1686,N_1625);
xor U3241 (N_3241,N_182,N_1519);
nand U3242 (N_3242,N_2123,N_723);
or U3243 (N_3243,N_548,N_2472);
or U3244 (N_3244,N_2373,N_642);
nand U3245 (N_3245,N_87,N_1426);
nand U3246 (N_3246,N_199,N_1031);
nand U3247 (N_3247,N_40,N_60);
nand U3248 (N_3248,N_1150,N_2042);
nor U3249 (N_3249,N_89,N_1003);
xor U3250 (N_3250,N_2100,N_821);
or U3251 (N_3251,N_1830,N_1970);
or U3252 (N_3252,N_550,N_6);
or U3253 (N_3253,N_533,N_1923);
nand U3254 (N_3254,N_2399,N_190);
nor U3255 (N_3255,N_727,N_1047);
and U3256 (N_3256,N_801,N_1142);
or U3257 (N_3257,N_965,N_597);
or U3258 (N_3258,N_337,N_1809);
nor U3259 (N_3259,N_1515,N_131);
nor U3260 (N_3260,N_1329,N_210);
nor U3261 (N_3261,N_390,N_460);
nor U3262 (N_3262,N_1503,N_449);
nand U3263 (N_3263,N_1927,N_1762);
and U3264 (N_3264,N_966,N_107);
and U3265 (N_3265,N_1229,N_895);
nor U3266 (N_3266,N_1208,N_1467);
nor U3267 (N_3267,N_2413,N_1690);
nand U3268 (N_3268,N_2200,N_1099);
nor U3269 (N_3269,N_1634,N_891);
nor U3270 (N_3270,N_1982,N_1374);
and U3271 (N_3271,N_858,N_905);
nand U3272 (N_3272,N_1714,N_221);
nand U3273 (N_3273,N_898,N_738);
and U3274 (N_3274,N_1571,N_2030);
nand U3275 (N_3275,N_1607,N_2360);
or U3276 (N_3276,N_1233,N_174);
and U3277 (N_3277,N_1801,N_582);
or U3278 (N_3278,N_1615,N_312);
nand U3279 (N_3279,N_1070,N_1322);
nor U3280 (N_3280,N_588,N_1471);
or U3281 (N_3281,N_520,N_1071);
nor U3282 (N_3282,N_2485,N_1386);
and U3283 (N_3283,N_1685,N_2054);
nor U3284 (N_3284,N_1817,N_487);
nand U3285 (N_3285,N_775,N_1063);
or U3286 (N_3286,N_2040,N_280);
or U3287 (N_3287,N_328,N_555);
nor U3288 (N_3288,N_1946,N_180);
and U3289 (N_3289,N_1667,N_2124);
or U3290 (N_3290,N_2477,N_1179);
or U3291 (N_3291,N_1526,N_628);
nor U3292 (N_3292,N_1862,N_1696);
and U3293 (N_3293,N_2212,N_433);
or U3294 (N_3294,N_1244,N_2366);
nor U3295 (N_3295,N_798,N_1988);
or U3296 (N_3296,N_2229,N_2303);
nor U3297 (N_3297,N_451,N_1440);
nand U3298 (N_3298,N_1897,N_1441);
nor U3299 (N_3299,N_1106,N_930);
or U3300 (N_3300,N_607,N_1523);
or U3301 (N_3301,N_1989,N_1281);
or U3302 (N_3302,N_170,N_1205);
and U3303 (N_3303,N_103,N_2093);
nor U3304 (N_3304,N_1181,N_562);
nand U3305 (N_3305,N_2262,N_1865);
nor U3306 (N_3306,N_354,N_1360);
nand U3307 (N_3307,N_73,N_1678);
nand U3308 (N_3308,N_1497,N_2081);
nor U3309 (N_3309,N_868,N_1836);
nand U3310 (N_3310,N_980,N_1423);
and U3311 (N_3311,N_2365,N_717);
nand U3312 (N_3312,N_100,N_688);
or U3313 (N_3313,N_912,N_2272);
nand U3314 (N_3314,N_1948,N_1287);
and U3315 (N_3315,N_819,N_1249);
nor U3316 (N_3316,N_1147,N_1308);
and U3317 (N_3317,N_142,N_599);
and U3318 (N_3318,N_9,N_423);
or U3319 (N_3319,N_1582,N_2415);
and U3320 (N_3320,N_826,N_1845);
nor U3321 (N_3321,N_901,N_873);
nand U3322 (N_3322,N_2043,N_1421);
nand U3323 (N_3323,N_2177,N_1723);
or U3324 (N_3324,N_1560,N_575);
or U3325 (N_3325,N_1551,N_1819);
nand U3326 (N_3326,N_992,N_2145);
and U3327 (N_3327,N_698,N_2265);
nor U3328 (N_3328,N_1145,N_571);
and U3329 (N_3329,N_2118,N_126);
or U3330 (N_3330,N_1086,N_613);
nand U3331 (N_3331,N_532,N_1466);
or U3332 (N_3332,N_1005,N_1701);
or U3333 (N_3333,N_843,N_2079);
nand U3334 (N_3334,N_1043,N_1542);
nor U3335 (N_3335,N_2228,N_666);
nand U3336 (N_3336,N_1905,N_689);
and U3337 (N_3337,N_2488,N_2403);
nand U3338 (N_3338,N_604,N_1641);
nand U3339 (N_3339,N_1014,N_1096);
and U3340 (N_3340,N_1947,N_1987);
or U3341 (N_3341,N_1860,N_1724);
nor U3342 (N_3342,N_1895,N_1683);
or U3343 (N_3343,N_463,N_2204);
nand U3344 (N_3344,N_1602,N_147);
nand U3345 (N_3345,N_883,N_99);
and U3346 (N_3346,N_660,N_1945);
or U3347 (N_3347,N_2008,N_636);
nand U3348 (N_3348,N_2340,N_272);
xor U3349 (N_3349,N_2202,N_501);
or U3350 (N_3350,N_2271,N_2209);
nor U3351 (N_3351,N_1012,N_786);
or U3352 (N_3352,N_264,N_2444);
nand U3353 (N_3353,N_1438,N_1619);
nor U3354 (N_3354,N_1843,N_568);
nand U3355 (N_3355,N_1180,N_53);
nand U3356 (N_3356,N_304,N_77);
or U3357 (N_3357,N_2408,N_1148);
or U3358 (N_3358,N_947,N_802);
nand U3359 (N_3359,N_651,N_859);
and U3360 (N_3360,N_2188,N_1779);
nor U3361 (N_3361,N_2331,N_598);
and U3362 (N_3362,N_324,N_2138);
or U3363 (N_3363,N_349,N_1725);
nor U3364 (N_3364,N_1608,N_2020);
nand U3365 (N_3365,N_90,N_2440);
nand U3366 (N_3366,N_857,N_972);
nor U3367 (N_3367,N_1077,N_347);
nand U3368 (N_3368,N_1478,N_1806);
and U3369 (N_3369,N_2310,N_1662);
and U3370 (N_3370,N_2289,N_62);
nand U3371 (N_3371,N_114,N_553);
nand U3372 (N_3372,N_602,N_476);
and U3373 (N_3373,N_1296,N_1264);
nor U3374 (N_3374,N_1617,N_294);
nand U3375 (N_3375,N_852,N_486);
nor U3376 (N_3376,N_765,N_1307);
or U3377 (N_3377,N_1616,N_2425);
nor U3378 (N_3378,N_1383,N_1447);
nor U3379 (N_3379,N_735,N_1481);
nor U3380 (N_3380,N_538,N_439);
and U3381 (N_3381,N_685,N_1729);
xnor U3382 (N_3382,N_19,N_1289);
or U3383 (N_3383,N_2022,N_1476);
nor U3384 (N_3384,N_2392,N_1039);
or U3385 (N_3385,N_2309,N_999);
and U3386 (N_3386,N_1277,N_519);
nand U3387 (N_3387,N_998,N_279);
nand U3388 (N_3388,N_1271,N_1929);
nor U3389 (N_3389,N_284,N_245);
or U3390 (N_3390,N_1203,N_1922);
nor U3391 (N_3391,N_914,N_434);
nor U3392 (N_3392,N_946,N_2491);
or U3393 (N_3393,N_191,N_743);
or U3394 (N_3394,N_219,N_150);
nor U3395 (N_3395,N_442,N_216);
nor U3396 (N_3396,N_2077,N_890);
or U3397 (N_3397,N_2245,N_2317);
nor U3398 (N_3398,N_671,N_746);
nand U3399 (N_3399,N_2296,N_46);
nor U3400 (N_3400,N_830,N_484);
and U3401 (N_3401,N_783,N_505);
nand U3402 (N_3402,N_188,N_1767);
or U3403 (N_3403,N_1282,N_814);
and U3404 (N_3404,N_459,N_49);
and U3405 (N_3405,N_2082,N_2065);
nand U3406 (N_3406,N_2189,N_944);
and U3407 (N_3407,N_725,N_1680);
nand U3408 (N_3408,N_1650,N_389);
and U3409 (N_3409,N_672,N_876);
and U3410 (N_3410,N_940,N_1397);
nor U3411 (N_3411,N_653,N_2376);
or U3412 (N_3412,N_1403,N_124);
and U3413 (N_3413,N_163,N_455);
and U3414 (N_3414,N_1385,N_899);
and U3415 (N_3415,N_1162,N_2135);
nand U3416 (N_3416,N_408,N_2242);
and U3417 (N_3417,N_513,N_1537);
nand U3418 (N_3418,N_936,N_552);
and U3419 (N_3419,N_195,N_828);
or U3420 (N_3420,N_1668,N_1525);
nand U3421 (N_3421,N_865,N_1797);
and U3422 (N_3422,N_441,N_1097);
nand U3423 (N_3423,N_664,N_1444);
nor U3424 (N_3424,N_448,N_351);
nand U3425 (N_3425,N_1030,N_1367);
and U3426 (N_3426,N_1649,N_1341);
or U3427 (N_3427,N_2,N_518);
or U3428 (N_3428,N_1088,N_1453);
and U3429 (N_3429,N_2343,N_2378);
or U3430 (N_3430,N_2258,N_1213);
and U3431 (N_3431,N_939,N_1349);
nand U3432 (N_3432,N_1311,N_241);
and U3433 (N_3433,N_2214,N_1076);
and U3434 (N_3434,N_570,N_425);
nand U3435 (N_3435,N_1749,N_1327);
and U3436 (N_3436,N_1198,N_1100);
and U3437 (N_3437,N_836,N_471);
and U3438 (N_3438,N_1669,N_1131);
or U3439 (N_3439,N_803,N_71);
and U3440 (N_3440,N_511,N_770);
nand U3441 (N_3441,N_327,N_1398);
nor U3442 (N_3442,N_1137,N_888);
or U3443 (N_3443,N_1117,N_1078);
nor U3444 (N_3444,N_253,N_1278);
or U3445 (N_3445,N_2314,N_2395);
or U3446 (N_3446,N_2361,N_1116);
nand U3447 (N_3447,N_2058,N_1462);
nor U3448 (N_3448,N_1543,N_197);
or U3449 (N_3449,N_194,N_2152);
or U3450 (N_3450,N_1684,N_2064);
or U3451 (N_3451,N_461,N_674);
xnor U3452 (N_3452,N_2132,N_1219);
nand U3453 (N_3453,N_874,N_1598);
nor U3454 (N_3454,N_2391,N_2499);
or U3455 (N_3455,N_1618,N_762);
and U3456 (N_3456,N_595,N_835);
nor U3457 (N_3457,N_2297,N_1394);
or U3458 (N_3458,N_733,N_2492);
or U3459 (N_3459,N_1704,N_609);
and U3460 (N_3460,N_619,N_691);
nand U3461 (N_3461,N_839,N_589);
and U3462 (N_3462,N_382,N_2463);
xnor U3463 (N_3463,N_1222,N_1732);
and U3464 (N_3464,N_1588,N_1549);
nor U3465 (N_3465,N_2084,N_1169);
nor U3466 (N_3466,N_2184,N_1422);
nand U3467 (N_3467,N_889,N_78);
nor U3468 (N_3468,N_61,N_959);
nor U3469 (N_3469,N_928,N_1884);
nor U3470 (N_3470,N_1883,N_120);
and U3471 (N_3471,N_842,N_2169);
or U3472 (N_3472,N_684,N_1939);
nor U3473 (N_3473,N_2041,N_493);
nor U3474 (N_3474,N_1639,N_1315);
or U3475 (N_3475,N_1540,N_924);
nor U3476 (N_3476,N_1713,N_1893);
or U3477 (N_3477,N_2496,N_1183);
and U3478 (N_3478,N_650,N_1681);
and U3479 (N_3479,N_1110,N_1720);
or U3480 (N_3480,N_2156,N_616);
and U3481 (N_3481,N_283,N_1316);
nor U3482 (N_3482,N_2448,N_1558);
nand U3483 (N_3483,N_2275,N_665);
nor U3484 (N_3484,N_1053,N_63);
nand U3485 (N_3485,N_45,N_1414);
nand U3486 (N_3486,N_215,N_1612);
nand U3487 (N_3487,N_1495,N_1538);
nand U3488 (N_3488,N_1357,N_1670);
nor U3489 (N_3489,N_306,N_1446);
nor U3490 (N_3490,N_1396,N_634);
nand U3491 (N_3491,N_136,N_1748);
nor U3492 (N_3492,N_1112,N_1889);
nor U3493 (N_3493,N_1353,N_1564);
or U3494 (N_3494,N_25,N_796);
or U3495 (N_3495,N_1826,N_1521);
and U3496 (N_3496,N_1236,N_1218);
nand U3497 (N_3497,N_509,N_1146);
or U3498 (N_3498,N_1164,N_813);
or U3499 (N_3499,N_2197,N_1331);
nor U3500 (N_3500,N_357,N_1347);
and U3501 (N_3501,N_547,N_325);
or U3502 (N_3502,N_1879,N_307);
or U3503 (N_3503,N_2117,N_113);
or U3504 (N_3504,N_491,N_1803);
or U3505 (N_3505,N_2426,N_1699);
nand U3506 (N_3506,N_2000,N_1375);
and U3507 (N_3507,N_1997,N_943);
nand U3508 (N_3508,N_2033,N_2203);
and U3509 (N_3509,N_305,N_1479);
nand U3510 (N_3510,N_1442,N_477);
and U3511 (N_3511,N_101,N_606);
nor U3512 (N_3512,N_1520,N_631);
or U3513 (N_3513,N_2266,N_356);
and U3514 (N_3514,N_39,N_2090);
and U3515 (N_3515,N_2390,N_446);
nand U3516 (N_3516,N_884,N_1532);
nand U3517 (N_3517,N_1250,N_711);
nand U3518 (N_3518,N_369,N_2036);
nor U3519 (N_3519,N_1757,N_1597);
nor U3520 (N_3520,N_610,N_720);
and U3521 (N_3521,N_573,N_2216);
and U3522 (N_3522,N_2253,N_1553);
or U3523 (N_3523,N_2347,N_1914);
or U3524 (N_3524,N_844,N_716);
or U3525 (N_3525,N_1944,N_179);
nand U3526 (N_3526,N_861,N_329);
nand U3527 (N_3527,N_208,N_97);
nor U3528 (N_3528,N_1046,N_30);
and U3529 (N_3529,N_2276,N_576);
nor U3530 (N_3530,N_1963,N_160);
nor U3531 (N_3531,N_1351,N_544);
nand U3532 (N_3532,N_867,N_1960);
nor U3533 (N_3533,N_2495,N_792);
nor U3534 (N_3534,N_1661,N_2051);
nor U3535 (N_3535,N_1010,N_1778);
and U3536 (N_3536,N_736,N_2111);
nand U3537 (N_3537,N_600,N_2438);
and U3538 (N_3538,N_1358,N_318);
or U3539 (N_3539,N_2270,N_1365);
nand U3540 (N_3540,N_2056,N_537);
xnor U3541 (N_3541,N_623,N_2235);
and U3542 (N_3542,N_2196,N_2349);
xnor U3543 (N_3543,N_1133,N_1657);
and U3544 (N_3544,N_1570,N_1595);
and U3545 (N_3545,N_1041,N_1671);
and U3546 (N_3546,N_2301,N_2410);
or U3547 (N_3547,N_207,N_968);
or U3548 (N_3548,N_2121,N_1742);
nor U3549 (N_3549,N_363,N_386);
nand U3550 (N_3550,N_1864,N_2244);
nor U3551 (N_3551,N_239,N_259);
nand U3552 (N_3552,N_1645,N_522);
nor U3553 (N_3553,N_1210,N_1393);
nand U3554 (N_3554,N_2167,N_787);
nor U3555 (N_3555,N_622,N_2429);
nand U3556 (N_3556,N_734,N_413);
nand U3557 (N_3557,N_1581,N_567);
nor U3558 (N_3558,N_452,N_2150);
nand U3559 (N_3559,N_1636,N_1252);
or U3560 (N_3560,N_1232,N_2099);
nand U3561 (N_3561,N_1115,N_2226);
and U3562 (N_3562,N_1051,N_742);
or U3563 (N_3563,N_2086,N_479);
and U3564 (N_3564,N_748,N_630);
and U3565 (N_3565,N_2374,N_745);
nor U3566 (N_3566,N_784,N_2004);
nor U3567 (N_3567,N_230,N_1892);
or U3568 (N_3568,N_2173,N_5);
nor U3569 (N_3569,N_703,N_1429);
or U3570 (N_3570,N_1215,N_1206);
nor U3571 (N_3571,N_785,N_1348);
nor U3572 (N_3572,N_2038,N_1771);
nor U3573 (N_3573,N_394,N_654);
nor U3574 (N_3574,N_1310,N_138);
or U3575 (N_3575,N_1185,N_41);
nor U3576 (N_3576,N_1764,N_2274);
nor U3577 (N_3577,N_2104,N_919);
and U3578 (N_3578,N_1983,N_132);
and U3579 (N_3579,N_1805,N_1505);
nand U3580 (N_3580,N_133,N_50);
nor U3581 (N_3581,N_1297,N_1379);
nor U3582 (N_3582,N_1140,N_2255);
and U3583 (N_3583,N_266,N_2362);
or U3584 (N_3584,N_1886,N_694);
nor U3585 (N_3585,N_201,N_848);
nand U3586 (N_3586,N_652,N_2181);
and U3587 (N_3587,N_1554,N_246);
and U3588 (N_3588,N_371,N_1938);
and U3589 (N_3589,N_1728,N_1784);
or U3590 (N_3590,N_2406,N_350);
nand U3591 (N_3591,N_403,N_1152);
or U3592 (N_3592,N_1127,N_367);
nor U3593 (N_3593,N_1758,N_1072);
and U3594 (N_3594,N_1687,N_431);
nor U3595 (N_3595,N_2341,N_395);
and U3596 (N_3596,N_2263,N_879);
or U3597 (N_3597,N_1212,N_756);
or U3598 (N_3598,N_1335,N_903);
nand U3599 (N_3599,N_365,N_388);
xor U3600 (N_3600,N_2498,N_2018);
or U3601 (N_3601,N_1018,N_1666);
and U3602 (N_3602,N_162,N_2031);
nand U3603 (N_3603,N_254,N_1876);
nor U3604 (N_3604,N_1443,N_1103);
nand U3605 (N_3605,N_894,N_1770);
and U3606 (N_3606,N_14,N_1034);
nand U3607 (N_3607,N_1464,N_400);
nand U3608 (N_3608,N_2103,N_1589);
nor U3609 (N_3609,N_2396,N_1765);
nor U3610 (N_3610,N_2159,N_102);
and U3611 (N_3611,N_2239,N_680);
nand U3612 (N_3612,N_764,N_1663);
and U3613 (N_3613,N_1605,N_2333);
or U3614 (N_3614,N_675,N_2354);
nor U3615 (N_3615,N_594,N_495);
and U3616 (N_3616,N_1073,N_950);
nor U3617 (N_3617,N_1079,N_2028);
or U3618 (N_3618,N_1175,N_1048);
nand U3619 (N_3619,N_1500,N_1659);
xnor U3620 (N_3620,N_1111,N_2131);
nor U3621 (N_3621,N_1456,N_846);
nor U3622 (N_3622,N_2300,N_508);
or U3623 (N_3623,N_1837,N_1610);
nor U3624 (N_3624,N_1029,N_1508);
nor U3625 (N_3625,N_590,N_43);
or U3626 (N_3626,N_892,N_1856);
or U3627 (N_3627,N_220,N_1972);
nor U3628 (N_3628,N_57,N_1098);
and U3629 (N_3629,N_1491,N_1992);
nand U3630 (N_3630,N_211,N_235);
nand U3631 (N_3631,N_605,N_2261);
nor U3632 (N_3632,N_27,N_1235);
and U3633 (N_3633,N_1480,N_834);
nor U3634 (N_3634,N_2066,N_1430);
nand U3635 (N_3635,N_379,N_541);
nand U3636 (N_3636,N_2388,N_169);
nand U3637 (N_3637,N_872,N_1993);
or U3638 (N_3638,N_621,N_569);
nand U3639 (N_3639,N_1242,N_1590);
nand U3640 (N_3640,N_186,N_825);
nand U3641 (N_3641,N_1015,N_2260);
or U3642 (N_3642,N_1135,N_2475);
and U3643 (N_3643,N_1234,N_788);
nand U3644 (N_3644,N_1867,N_563);
and U3645 (N_3645,N_856,N_1021);
or U3646 (N_3646,N_2430,N_1962);
or U3647 (N_3647,N_158,N_1818);
nor U3648 (N_3648,N_248,N_2327);
nand U3649 (N_3649,N_2211,N_435);
and U3650 (N_3650,N_1019,N_2246);
nor U3651 (N_3651,N_370,N_1660);
and U3652 (N_3652,N_2453,N_1214);
nand U3653 (N_3653,N_603,N_95);
and U3654 (N_3654,N_1493,N_1149);
nand U3655 (N_3655,N_1395,N_862);
nand U3656 (N_3656,N_1730,N_34);
nand U3657 (N_3657,N_2482,N_1981);
nor U3658 (N_3658,N_226,N_1731);
and U3659 (N_3659,N_647,N_769);
or U3660 (N_3660,N_577,N_1461);
nand U3661 (N_3661,N_1318,N_2176);
and U3662 (N_3662,N_2023,N_2006);
or U3663 (N_3663,N_1159,N_1511);
nand U3664 (N_3664,N_962,N_1991);
nand U3665 (N_3665,N_931,N_1120);
nand U3666 (N_3666,N_2215,N_624);
and U3667 (N_3667,N_1788,N_2001);
nand U3668 (N_3668,N_1592,N_1485);
or U3669 (N_3669,N_1527,N_1783);
or U3670 (N_3670,N_229,N_676);
nor U3671 (N_3671,N_2443,N_2021);
xnor U3672 (N_3672,N_33,N_1487);
nand U3673 (N_3673,N_1563,N_1067);
and U3674 (N_3674,N_2291,N_277);
or U3675 (N_3675,N_1216,N_1049);
and U3676 (N_3676,N_359,N_2350);
nand U3677 (N_3677,N_1038,N_2285);
nand U3678 (N_3678,N_2191,N_249);
nand U3679 (N_3679,N_1877,N_167);
nor U3680 (N_3680,N_1903,N_1196);
nand U3681 (N_3681,N_1119,N_1785);
nand U3682 (N_3682,N_2128,N_1240);
or U3683 (N_3683,N_1691,N_1908);
or U3684 (N_3684,N_1747,N_1514);
and U3685 (N_3685,N_3,N_1090);
nor U3686 (N_3686,N_535,N_172);
and U3687 (N_3687,N_1209,N_48);
or U3688 (N_3688,N_4,N_2048);
nor U3689 (N_3689,N_342,N_2484);
nor U3690 (N_3690,N_140,N_1875);
or U3691 (N_3691,N_1761,N_1074);
nor U3692 (N_3692,N_549,N_638);
or U3693 (N_3693,N_72,N_1911);
nand U3694 (N_3694,N_2165,N_987);
nand U3695 (N_3695,N_222,N_1688);
and U3696 (N_3696,N_24,N_83);
nor U3697 (N_3697,N_994,N_301);
and U3698 (N_3698,N_2198,N_640);
or U3699 (N_3699,N_2315,N_262);
or U3700 (N_3700,N_1483,N_108);
nor U3701 (N_3701,N_297,N_2068);
nand U3702 (N_3702,N_1813,N_1174);
nor U3703 (N_3703,N_23,N_2490);
and U3704 (N_3704,N_2005,N_332);
and U3705 (N_3705,N_1001,N_916);
or U3706 (N_3706,N_192,N_1524);
nor U3707 (N_3707,N_574,N_1896);
and U3708 (N_3708,N_2222,N_233);
and U3709 (N_3709,N_1417,N_1874);
nor U3710 (N_3710,N_2452,N_1138);
or U3711 (N_3711,N_1833,N_969);
nand U3712 (N_3712,N_339,N_2355);
and U3713 (N_3713,N_1094,N_1986);
xor U3714 (N_3714,N_923,N_1774);
or U3715 (N_3715,N_1798,N_1572);
nor U3716 (N_3716,N_831,N_2161);
or U3717 (N_3717,N_29,N_1849);
and U3718 (N_3718,N_1114,N_1452);
and U3719 (N_3719,N_641,N_767);
nand U3720 (N_3720,N_1623,N_1499);
and U3721 (N_3721,N_1129,N_1050);
and U3722 (N_3722,N_82,N_1391);
or U3723 (N_3723,N_1811,N_1269);
nand U3724 (N_3724,N_1400,N_2180);
nand U3725 (N_3725,N_1606,N_1800);
and U3726 (N_3726,N_1506,N_130);
nor U3727 (N_3727,N_2011,N_2063);
or U3728 (N_3728,N_2402,N_2325);
and U3729 (N_3729,N_1812,N_906);
and U3730 (N_3730,N_1392,N_1808);
or U3731 (N_3731,N_293,N_2013);
nor U3732 (N_3732,N_309,N_1702);
nand U3733 (N_3733,N_601,N_900);
xnor U3734 (N_3734,N_1241,N_1207);
and U3735 (N_3735,N_232,N_909);
nor U3736 (N_3736,N_2483,N_1486);
nor U3737 (N_3737,N_1628,N_1885);
nor U3738 (N_3738,N_1585,N_1126);
nor U3739 (N_3739,N_244,N_1587);
nor U3740 (N_3740,N_2187,N_2183);
and U3741 (N_3741,N_926,N_804);
or U3742 (N_3742,N_427,N_465);
and U3743 (N_3743,N_1163,N_1584);
or U3744 (N_3744,N_333,N_396);
nand U3745 (N_3745,N_993,N_176);
and U3746 (N_3746,N_949,N_496);
nand U3747 (N_3747,N_2223,N_1160);
nand U3748 (N_3748,N_536,N_502);
nor U3749 (N_3749,N_1332,N_2494);
and U3750 (N_3750,N_1662,N_1555);
nor U3751 (N_3751,N_2482,N_581);
or U3752 (N_3752,N_2007,N_1660);
nand U3753 (N_3753,N_1532,N_1643);
and U3754 (N_3754,N_42,N_1905);
nor U3755 (N_3755,N_2262,N_1031);
and U3756 (N_3756,N_731,N_1789);
nor U3757 (N_3757,N_308,N_1021);
and U3758 (N_3758,N_645,N_1528);
nand U3759 (N_3759,N_983,N_1034);
nand U3760 (N_3760,N_405,N_2494);
xnor U3761 (N_3761,N_1856,N_1441);
and U3762 (N_3762,N_1430,N_1447);
or U3763 (N_3763,N_1634,N_441);
and U3764 (N_3764,N_451,N_351);
or U3765 (N_3765,N_509,N_1964);
nand U3766 (N_3766,N_282,N_708);
or U3767 (N_3767,N_1661,N_1048);
and U3768 (N_3768,N_2486,N_693);
or U3769 (N_3769,N_244,N_2237);
nor U3770 (N_3770,N_1034,N_2430);
nor U3771 (N_3771,N_1863,N_2319);
or U3772 (N_3772,N_2450,N_597);
nand U3773 (N_3773,N_659,N_1390);
or U3774 (N_3774,N_2307,N_2407);
and U3775 (N_3775,N_157,N_1284);
or U3776 (N_3776,N_980,N_2443);
or U3777 (N_3777,N_1433,N_2281);
or U3778 (N_3778,N_1434,N_1810);
and U3779 (N_3779,N_456,N_716);
and U3780 (N_3780,N_1312,N_613);
nor U3781 (N_3781,N_17,N_910);
nor U3782 (N_3782,N_1255,N_1094);
nand U3783 (N_3783,N_828,N_2185);
and U3784 (N_3784,N_480,N_1040);
or U3785 (N_3785,N_1998,N_534);
or U3786 (N_3786,N_1745,N_1866);
nor U3787 (N_3787,N_80,N_1249);
nand U3788 (N_3788,N_186,N_62);
nand U3789 (N_3789,N_1266,N_1552);
nand U3790 (N_3790,N_2310,N_2476);
nor U3791 (N_3791,N_2170,N_2279);
and U3792 (N_3792,N_59,N_792);
nand U3793 (N_3793,N_1426,N_479);
nor U3794 (N_3794,N_687,N_2126);
and U3795 (N_3795,N_770,N_2236);
nand U3796 (N_3796,N_2011,N_244);
nor U3797 (N_3797,N_596,N_1361);
nand U3798 (N_3798,N_216,N_2224);
nor U3799 (N_3799,N_763,N_2162);
nand U3800 (N_3800,N_2480,N_682);
or U3801 (N_3801,N_1882,N_2208);
or U3802 (N_3802,N_1405,N_979);
and U3803 (N_3803,N_640,N_1315);
or U3804 (N_3804,N_2278,N_317);
or U3805 (N_3805,N_316,N_1816);
nand U3806 (N_3806,N_571,N_613);
nand U3807 (N_3807,N_2124,N_2102);
and U3808 (N_3808,N_1285,N_2111);
nand U3809 (N_3809,N_1895,N_1110);
nand U3810 (N_3810,N_875,N_1028);
and U3811 (N_3811,N_1887,N_1700);
nor U3812 (N_3812,N_282,N_743);
and U3813 (N_3813,N_5,N_2294);
and U3814 (N_3814,N_1951,N_1498);
nor U3815 (N_3815,N_1568,N_466);
or U3816 (N_3816,N_1263,N_2105);
or U3817 (N_3817,N_840,N_883);
and U3818 (N_3818,N_1674,N_1091);
or U3819 (N_3819,N_1752,N_398);
and U3820 (N_3820,N_2250,N_147);
and U3821 (N_3821,N_2207,N_1530);
or U3822 (N_3822,N_2173,N_1122);
or U3823 (N_3823,N_1436,N_255);
or U3824 (N_3824,N_1475,N_1298);
nand U3825 (N_3825,N_354,N_1173);
nor U3826 (N_3826,N_1671,N_1297);
or U3827 (N_3827,N_2037,N_615);
nand U3828 (N_3828,N_2362,N_1147);
and U3829 (N_3829,N_1449,N_833);
nor U3830 (N_3830,N_1498,N_1419);
nand U3831 (N_3831,N_1691,N_2123);
nand U3832 (N_3832,N_1828,N_1273);
nor U3833 (N_3833,N_195,N_575);
nor U3834 (N_3834,N_493,N_918);
or U3835 (N_3835,N_1746,N_327);
and U3836 (N_3836,N_1365,N_1327);
or U3837 (N_3837,N_2153,N_869);
nand U3838 (N_3838,N_1391,N_367);
nor U3839 (N_3839,N_779,N_1437);
or U3840 (N_3840,N_1688,N_174);
nor U3841 (N_3841,N_1971,N_2021);
or U3842 (N_3842,N_1222,N_649);
or U3843 (N_3843,N_2012,N_2359);
and U3844 (N_3844,N_912,N_1712);
nand U3845 (N_3845,N_768,N_1923);
or U3846 (N_3846,N_419,N_1077);
nand U3847 (N_3847,N_515,N_95);
nand U3848 (N_3848,N_1263,N_1064);
or U3849 (N_3849,N_2268,N_21);
nor U3850 (N_3850,N_135,N_221);
and U3851 (N_3851,N_2321,N_1446);
and U3852 (N_3852,N_1116,N_600);
nor U3853 (N_3853,N_484,N_1755);
xnor U3854 (N_3854,N_2196,N_209);
nand U3855 (N_3855,N_1417,N_1960);
nor U3856 (N_3856,N_1933,N_700);
nor U3857 (N_3857,N_542,N_2435);
nor U3858 (N_3858,N_2459,N_1067);
nand U3859 (N_3859,N_1050,N_461);
and U3860 (N_3860,N_2449,N_795);
and U3861 (N_3861,N_91,N_120);
nand U3862 (N_3862,N_952,N_1526);
or U3863 (N_3863,N_2259,N_2215);
nor U3864 (N_3864,N_1799,N_297);
nor U3865 (N_3865,N_1973,N_2472);
or U3866 (N_3866,N_688,N_162);
or U3867 (N_3867,N_2208,N_1687);
or U3868 (N_3868,N_2494,N_289);
or U3869 (N_3869,N_1521,N_1360);
and U3870 (N_3870,N_224,N_1558);
nor U3871 (N_3871,N_693,N_2336);
nor U3872 (N_3872,N_1413,N_1663);
or U3873 (N_3873,N_675,N_416);
nand U3874 (N_3874,N_420,N_1568);
xor U3875 (N_3875,N_693,N_62);
and U3876 (N_3876,N_1009,N_253);
nand U3877 (N_3877,N_1258,N_992);
nand U3878 (N_3878,N_2328,N_2148);
nor U3879 (N_3879,N_1294,N_1678);
and U3880 (N_3880,N_888,N_850);
or U3881 (N_3881,N_2397,N_1821);
and U3882 (N_3882,N_2343,N_1056);
nand U3883 (N_3883,N_1105,N_1801);
or U3884 (N_3884,N_2063,N_506);
or U3885 (N_3885,N_347,N_1504);
nand U3886 (N_3886,N_522,N_1672);
or U3887 (N_3887,N_2125,N_451);
and U3888 (N_3888,N_1490,N_669);
nand U3889 (N_3889,N_584,N_2456);
and U3890 (N_3890,N_754,N_222);
nand U3891 (N_3891,N_2165,N_15);
or U3892 (N_3892,N_337,N_1783);
and U3893 (N_3893,N_1509,N_183);
nand U3894 (N_3894,N_1360,N_715);
nor U3895 (N_3895,N_1483,N_2354);
nor U3896 (N_3896,N_714,N_2461);
nand U3897 (N_3897,N_261,N_1789);
or U3898 (N_3898,N_1957,N_1273);
nor U3899 (N_3899,N_865,N_1847);
or U3900 (N_3900,N_589,N_1339);
nand U3901 (N_3901,N_347,N_459);
and U3902 (N_3902,N_64,N_1658);
and U3903 (N_3903,N_932,N_1763);
nor U3904 (N_3904,N_653,N_1104);
nand U3905 (N_3905,N_344,N_1733);
and U3906 (N_3906,N_137,N_1832);
nor U3907 (N_3907,N_2295,N_1860);
nor U3908 (N_3908,N_1482,N_226);
nor U3909 (N_3909,N_1599,N_2168);
xnor U3910 (N_3910,N_2016,N_1180);
nor U3911 (N_3911,N_1295,N_1301);
nand U3912 (N_3912,N_624,N_360);
and U3913 (N_3913,N_1847,N_801);
and U3914 (N_3914,N_1706,N_1862);
nor U3915 (N_3915,N_1197,N_1940);
nor U3916 (N_3916,N_1890,N_892);
nor U3917 (N_3917,N_1622,N_2437);
nand U3918 (N_3918,N_2450,N_2165);
nor U3919 (N_3919,N_1387,N_1095);
nor U3920 (N_3920,N_906,N_1633);
nand U3921 (N_3921,N_453,N_2113);
nor U3922 (N_3922,N_223,N_2385);
nor U3923 (N_3923,N_2137,N_1102);
and U3924 (N_3924,N_1183,N_1536);
nand U3925 (N_3925,N_1466,N_1827);
and U3926 (N_3926,N_2015,N_1923);
nor U3927 (N_3927,N_395,N_2053);
or U3928 (N_3928,N_732,N_2218);
nand U3929 (N_3929,N_897,N_415);
and U3930 (N_3930,N_1583,N_1472);
and U3931 (N_3931,N_646,N_1887);
or U3932 (N_3932,N_544,N_2240);
and U3933 (N_3933,N_1974,N_2178);
and U3934 (N_3934,N_1163,N_1075);
or U3935 (N_3935,N_1759,N_1692);
and U3936 (N_3936,N_1704,N_2367);
nand U3937 (N_3937,N_1880,N_469);
or U3938 (N_3938,N_480,N_751);
nor U3939 (N_3939,N_1400,N_1798);
nand U3940 (N_3940,N_1701,N_100);
or U3941 (N_3941,N_1559,N_341);
or U3942 (N_3942,N_1870,N_1460);
nand U3943 (N_3943,N_2166,N_771);
nor U3944 (N_3944,N_771,N_1778);
or U3945 (N_3945,N_1864,N_1638);
and U3946 (N_3946,N_1178,N_2344);
and U3947 (N_3947,N_2399,N_1587);
nand U3948 (N_3948,N_1626,N_1430);
or U3949 (N_3949,N_375,N_58);
nand U3950 (N_3950,N_2217,N_1592);
and U3951 (N_3951,N_2342,N_353);
nor U3952 (N_3952,N_1491,N_1726);
nor U3953 (N_3953,N_788,N_2058);
or U3954 (N_3954,N_895,N_1407);
or U3955 (N_3955,N_252,N_18);
nand U3956 (N_3956,N_991,N_304);
nor U3957 (N_3957,N_223,N_1456);
or U3958 (N_3958,N_1065,N_991);
nor U3959 (N_3959,N_926,N_649);
nor U3960 (N_3960,N_1279,N_2234);
nor U3961 (N_3961,N_2163,N_2215);
nand U3962 (N_3962,N_1555,N_2405);
or U3963 (N_3963,N_1004,N_315);
nor U3964 (N_3964,N_924,N_2146);
and U3965 (N_3965,N_2051,N_1574);
nor U3966 (N_3966,N_1050,N_1713);
nor U3967 (N_3967,N_258,N_113);
nand U3968 (N_3968,N_1123,N_1853);
nand U3969 (N_3969,N_1980,N_649);
nor U3970 (N_3970,N_416,N_2174);
or U3971 (N_3971,N_1791,N_1952);
and U3972 (N_3972,N_1117,N_1792);
nor U3973 (N_3973,N_899,N_481);
nand U3974 (N_3974,N_2011,N_1917);
and U3975 (N_3975,N_1324,N_17);
nand U3976 (N_3976,N_142,N_2069);
or U3977 (N_3977,N_1731,N_277);
or U3978 (N_3978,N_306,N_108);
and U3979 (N_3979,N_1601,N_730);
nor U3980 (N_3980,N_1499,N_2287);
nand U3981 (N_3981,N_471,N_2390);
and U3982 (N_3982,N_214,N_2244);
or U3983 (N_3983,N_1074,N_445);
nor U3984 (N_3984,N_207,N_363);
nand U3985 (N_3985,N_2003,N_1753);
or U3986 (N_3986,N_1094,N_1950);
nand U3987 (N_3987,N_2290,N_57);
and U3988 (N_3988,N_306,N_1660);
nor U3989 (N_3989,N_2235,N_1555);
nand U3990 (N_3990,N_22,N_2045);
or U3991 (N_3991,N_1527,N_2316);
and U3992 (N_3992,N_637,N_2410);
xor U3993 (N_3993,N_1151,N_826);
and U3994 (N_3994,N_1740,N_360);
or U3995 (N_3995,N_967,N_65);
nand U3996 (N_3996,N_276,N_1854);
or U3997 (N_3997,N_1405,N_1549);
nor U3998 (N_3998,N_2302,N_348);
and U3999 (N_3999,N_746,N_1764);
nor U4000 (N_4000,N_603,N_2032);
and U4001 (N_4001,N_1075,N_2409);
or U4002 (N_4002,N_90,N_1032);
or U4003 (N_4003,N_2251,N_1453);
nor U4004 (N_4004,N_1736,N_2041);
nor U4005 (N_4005,N_358,N_2236);
and U4006 (N_4006,N_1012,N_805);
nand U4007 (N_4007,N_343,N_1842);
nor U4008 (N_4008,N_793,N_934);
nor U4009 (N_4009,N_45,N_2444);
and U4010 (N_4010,N_61,N_2219);
and U4011 (N_4011,N_10,N_1513);
nand U4012 (N_4012,N_1561,N_1550);
nand U4013 (N_4013,N_819,N_848);
nor U4014 (N_4014,N_2189,N_2390);
nor U4015 (N_4015,N_1560,N_2312);
nand U4016 (N_4016,N_891,N_1242);
and U4017 (N_4017,N_1600,N_2157);
and U4018 (N_4018,N_194,N_2239);
and U4019 (N_4019,N_2043,N_2169);
or U4020 (N_4020,N_961,N_787);
nor U4021 (N_4021,N_1491,N_2078);
nor U4022 (N_4022,N_902,N_1191);
or U4023 (N_4023,N_692,N_1889);
nor U4024 (N_4024,N_69,N_1349);
nor U4025 (N_4025,N_2407,N_2260);
nand U4026 (N_4026,N_1060,N_1418);
nor U4027 (N_4027,N_825,N_1521);
nand U4028 (N_4028,N_2405,N_575);
or U4029 (N_4029,N_1762,N_1288);
or U4030 (N_4030,N_945,N_1305);
and U4031 (N_4031,N_1867,N_944);
nand U4032 (N_4032,N_1570,N_1516);
and U4033 (N_4033,N_1888,N_260);
nor U4034 (N_4034,N_756,N_1517);
or U4035 (N_4035,N_2116,N_2287);
or U4036 (N_4036,N_332,N_834);
and U4037 (N_4037,N_2499,N_1246);
nand U4038 (N_4038,N_1504,N_2441);
or U4039 (N_4039,N_1257,N_1);
nand U4040 (N_4040,N_1007,N_2000);
nor U4041 (N_4041,N_1571,N_1848);
nand U4042 (N_4042,N_1955,N_215);
or U4043 (N_4043,N_189,N_498);
nor U4044 (N_4044,N_430,N_203);
or U4045 (N_4045,N_2241,N_1171);
and U4046 (N_4046,N_707,N_1138);
or U4047 (N_4047,N_2387,N_2231);
and U4048 (N_4048,N_1026,N_1816);
nor U4049 (N_4049,N_1821,N_285);
and U4050 (N_4050,N_1701,N_1613);
nand U4051 (N_4051,N_1598,N_1094);
or U4052 (N_4052,N_2125,N_1190);
xor U4053 (N_4053,N_847,N_792);
or U4054 (N_4054,N_2343,N_1002);
nor U4055 (N_4055,N_1039,N_1072);
nand U4056 (N_4056,N_462,N_707);
and U4057 (N_4057,N_217,N_727);
nand U4058 (N_4058,N_396,N_1814);
nor U4059 (N_4059,N_2234,N_1970);
or U4060 (N_4060,N_415,N_553);
nor U4061 (N_4061,N_977,N_758);
nand U4062 (N_4062,N_716,N_2496);
nor U4063 (N_4063,N_688,N_2342);
nor U4064 (N_4064,N_2172,N_1299);
nand U4065 (N_4065,N_2319,N_1621);
and U4066 (N_4066,N_2027,N_950);
nor U4067 (N_4067,N_2086,N_360);
or U4068 (N_4068,N_2116,N_1257);
nor U4069 (N_4069,N_1102,N_1895);
and U4070 (N_4070,N_1160,N_1070);
and U4071 (N_4071,N_738,N_2012);
nor U4072 (N_4072,N_109,N_157);
and U4073 (N_4073,N_125,N_1918);
and U4074 (N_4074,N_2036,N_721);
or U4075 (N_4075,N_606,N_440);
nand U4076 (N_4076,N_1023,N_1317);
and U4077 (N_4077,N_2166,N_1209);
or U4078 (N_4078,N_703,N_1559);
nor U4079 (N_4079,N_2411,N_1634);
or U4080 (N_4080,N_1520,N_808);
nor U4081 (N_4081,N_1502,N_1844);
and U4082 (N_4082,N_225,N_1083);
and U4083 (N_4083,N_1263,N_1427);
and U4084 (N_4084,N_25,N_1798);
nor U4085 (N_4085,N_146,N_1746);
and U4086 (N_4086,N_883,N_1480);
nand U4087 (N_4087,N_2380,N_2377);
and U4088 (N_4088,N_1273,N_1564);
nor U4089 (N_4089,N_660,N_1268);
and U4090 (N_4090,N_1126,N_966);
nor U4091 (N_4091,N_2248,N_1103);
or U4092 (N_4092,N_717,N_1423);
or U4093 (N_4093,N_566,N_509);
and U4094 (N_4094,N_2038,N_73);
and U4095 (N_4095,N_1261,N_2252);
and U4096 (N_4096,N_1013,N_138);
or U4097 (N_4097,N_938,N_1878);
nand U4098 (N_4098,N_1203,N_1721);
nor U4099 (N_4099,N_1067,N_531);
nor U4100 (N_4100,N_621,N_1553);
nand U4101 (N_4101,N_1728,N_264);
nor U4102 (N_4102,N_1336,N_1820);
nor U4103 (N_4103,N_1950,N_2161);
and U4104 (N_4104,N_1680,N_189);
nor U4105 (N_4105,N_1179,N_1588);
or U4106 (N_4106,N_1488,N_1237);
nand U4107 (N_4107,N_971,N_2489);
nand U4108 (N_4108,N_221,N_2170);
and U4109 (N_4109,N_2317,N_1682);
nor U4110 (N_4110,N_2086,N_2120);
nor U4111 (N_4111,N_1687,N_1080);
or U4112 (N_4112,N_2486,N_797);
or U4113 (N_4113,N_1200,N_1776);
nand U4114 (N_4114,N_2319,N_810);
nand U4115 (N_4115,N_1527,N_2039);
nand U4116 (N_4116,N_633,N_2170);
nand U4117 (N_4117,N_1556,N_1670);
nor U4118 (N_4118,N_232,N_1252);
and U4119 (N_4119,N_1102,N_747);
and U4120 (N_4120,N_1574,N_796);
nor U4121 (N_4121,N_2347,N_102);
or U4122 (N_4122,N_2486,N_1290);
nor U4123 (N_4123,N_1508,N_2485);
or U4124 (N_4124,N_561,N_418);
and U4125 (N_4125,N_907,N_219);
nand U4126 (N_4126,N_168,N_1008);
and U4127 (N_4127,N_83,N_195);
nand U4128 (N_4128,N_335,N_586);
nor U4129 (N_4129,N_2175,N_1068);
nand U4130 (N_4130,N_335,N_23);
nand U4131 (N_4131,N_1313,N_1762);
nand U4132 (N_4132,N_1778,N_383);
or U4133 (N_4133,N_1953,N_1373);
and U4134 (N_4134,N_65,N_1317);
or U4135 (N_4135,N_1756,N_1165);
nand U4136 (N_4136,N_2356,N_157);
nor U4137 (N_4137,N_1134,N_1142);
and U4138 (N_4138,N_1386,N_551);
and U4139 (N_4139,N_2168,N_1486);
nand U4140 (N_4140,N_1320,N_1297);
nand U4141 (N_4141,N_1884,N_14);
nor U4142 (N_4142,N_711,N_1920);
and U4143 (N_4143,N_467,N_270);
nand U4144 (N_4144,N_1401,N_798);
and U4145 (N_4145,N_1059,N_1326);
nor U4146 (N_4146,N_2063,N_1579);
nand U4147 (N_4147,N_1963,N_1549);
and U4148 (N_4148,N_2128,N_1893);
and U4149 (N_4149,N_2398,N_1915);
and U4150 (N_4150,N_1062,N_1132);
nand U4151 (N_4151,N_1052,N_1123);
xnor U4152 (N_4152,N_1482,N_232);
and U4153 (N_4153,N_636,N_1683);
nor U4154 (N_4154,N_752,N_66);
nand U4155 (N_4155,N_345,N_2285);
nand U4156 (N_4156,N_1782,N_195);
or U4157 (N_4157,N_2118,N_1692);
nand U4158 (N_4158,N_1986,N_2287);
and U4159 (N_4159,N_969,N_2178);
nand U4160 (N_4160,N_1786,N_402);
and U4161 (N_4161,N_120,N_1456);
or U4162 (N_4162,N_405,N_2182);
nor U4163 (N_4163,N_1819,N_1007);
or U4164 (N_4164,N_2016,N_833);
nor U4165 (N_4165,N_1453,N_1262);
or U4166 (N_4166,N_2357,N_606);
and U4167 (N_4167,N_1220,N_2281);
and U4168 (N_4168,N_1497,N_1959);
or U4169 (N_4169,N_2080,N_1429);
nand U4170 (N_4170,N_620,N_2008);
nor U4171 (N_4171,N_1857,N_142);
and U4172 (N_4172,N_1991,N_1822);
and U4173 (N_4173,N_441,N_978);
and U4174 (N_4174,N_875,N_185);
nor U4175 (N_4175,N_613,N_2195);
nand U4176 (N_4176,N_798,N_2265);
nand U4177 (N_4177,N_1781,N_416);
nor U4178 (N_4178,N_947,N_785);
or U4179 (N_4179,N_1784,N_2162);
nor U4180 (N_4180,N_255,N_863);
and U4181 (N_4181,N_1851,N_2490);
nand U4182 (N_4182,N_1533,N_2267);
nor U4183 (N_4183,N_427,N_1449);
nor U4184 (N_4184,N_1387,N_832);
or U4185 (N_4185,N_1131,N_374);
nand U4186 (N_4186,N_1930,N_617);
nand U4187 (N_4187,N_64,N_1396);
nand U4188 (N_4188,N_554,N_1708);
nand U4189 (N_4189,N_1756,N_905);
nor U4190 (N_4190,N_1950,N_936);
or U4191 (N_4191,N_420,N_974);
and U4192 (N_4192,N_1502,N_0);
xnor U4193 (N_4193,N_53,N_1611);
nor U4194 (N_4194,N_53,N_2028);
nor U4195 (N_4195,N_1695,N_2036);
nand U4196 (N_4196,N_856,N_1752);
and U4197 (N_4197,N_804,N_820);
or U4198 (N_4198,N_2367,N_2123);
or U4199 (N_4199,N_1926,N_2021);
and U4200 (N_4200,N_819,N_1538);
nand U4201 (N_4201,N_396,N_344);
or U4202 (N_4202,N_37,N_1347);
nand U4203 (N_4203,N_970,N_1870);
and U4204 (N_4204,N_2030,N_67);
and U4205 (N_4205,N_1913,N_1790);
or U4206 (N_4206,N_1103,N_483);
or U4207 (N_4207,N_2460,N_662);
nand U4208 (N_4208,N_154,N_1598);
or U4209 (N_4209,N_1523,N_1639);
nor U4210 (N_4210,N_436,N_1162);
nor U4211 (N_4211,N_1905,N_620);
or U4212 (N_4212,N_1105,N_1281);
or U4213 (N_4213,N_2443,N_648);
or U4214 (N_4214,N_2043,N_1986);
nand U4215 (N_4215,N_1455,N_198);
and U4216 (N_4216,N_2267,N_2466);
and U4217 (N_4217,N_566,N_987);
nand U4218 (N_4218,N_1697,N_1526);
nor U4219 (N_4219,N_954,N_1110);
nand U4220 (N_4220,N_325,N_165);
and U4221 (N_4221,N_1656,N_19);
nand U4222 (N_4222,N_2458,N_1185);
nor U4223 (N_4223,N_1555,N_1286);
nor U4224 (N_4224,N_2429,N_1847);
or U4225 (N_4225,N_1202,N_1388);
and U4226 (N_4226,N_999,N_2474);
or U4227 (N_4227,N_122,N_2302);
and U4228 (N_4228,N_1080,N_348);
nor U4229 (N_4229,N_549,N_502);
nor U4230 (N_4230,N_1543,N_2129);
or U4231 (N_4231,N_1111,N_2238);
nor U4232 (N_4232,N_1654,N_329);
nor U4233 (N_4233,N_1690,N_910);
or U4234 (N_4234,N_2410,N_1904);
xor U4235 (N_4235,N_1902,N_1924);
and U4236 (N_4236,N_1780,N_943);
xnor U4237 (N_4237,N_202,N_774);
nand U4238 (N_4238,N_1755,N_334);
nor U4239 (N_4239,N_278,N_939);
or U4240 (N_4240,N_1766,N_304);
and U4241 (N_4241,N_225,N_423);
or U4242 (N_4242,N_523,N_862);
nand U4243 (N_4243,N_674,N_25);
and U4244 (N_4244,N_2410,N_287);
or U4245 (N_4245,N_2388,N_1206);
nand U4246 (N_4246,N_881,N_1834);
or U4247 (N_4247,N_236,N_2207);
nand U4248 (N_4248,N_1112,N_2453);
or U4249 (N_4249,N_1709,N_364);
or U4250 (N_4250,N_2133,N_873);
or U4251 (N_4251,N_369,N_1003);
and U4252 (N_4252,N_779,N_635);
nand U4253 (N_4253,N_1397,N_1758);
nand U4254 (N_4254,N_922,N_1101);
nor U4255 (N_4255,N_2033,N_1276);
and U4256 (N_4256,N_153,N_2318);
and U4257 (N_4257,N_2163,N_795);
nand U4258 (N_4258,N_1236,N_2264);
nand U4259 (N_4259,N_2399,N_1473);
nand U4260 (N_4260,N_251,N_676);
nand U4261 (N_4261,N_163,N_2491);
and U4262 (N_4262,N_1583,N_2201);
nand U4263 (N_4263,N_1580,N_205);
and U4264 (N_4264,N_2487,N_1790);
or U4265 (N_4265,N_105,N_1231);
nor U4266 (N_4266,N_2154,N_1379);
nand U4267 (N_4267,N_966,N_245);
or U4268 (N_4268,N_1279,N_541);
or U4269 (N_4269,N_1020,N_1946);
or U4270 (N_4270,N_1515,N_1410);
or U4271 (N_4271,N_1735,N_48);
nor U4272 (N_4272,N_639,N_196);
or U4273 (N_4273,N_1100,N_1215);
nor U4274 (N_4274,N_325,N_2311);
and U4275 (N_4275,N_434,N_807);
nor U4276 (N_4276,N_2470,N_875);
or U4277 (N_4277,N_153,N_359);
and U4278 (N_4278,N_2337,N_1222);
and U4279 (N_4279,N_1640,N_2174);
or U4280 (N_4280,N_1223,N_2291);
and U4281 (N_4281,N_108,N_1);
nand U4282 (N_4282,N_2199,N_2299);
or U4283 (N_4283,N_2060,N_2405);
nand U4284 (N_4284,N_1181,N_1744);
and U4285 (N_4285,N_1279,N_1870);
and U4286 (N_4286,N_526,N_1552);
nor U4287 (N_4287,N_1785,N_298);
nand U4288 (N_4288,N_378,N_1918);
nand U4289 (N_4289,N_205,N_996);
nor U4290 (N_4290,N_1618,N_1951);
nand U4291 (N_4291,N_1954,N_520);
nor U4292 (N_4292,N_1590,N_560);
or U4293 (N_4293,N_669,N_895);
nor U4294 (N_4294,N_1320,N_1046);
nand U4295 (N_4295,N_2067,N_844);
or U4296 (N_4296,N_1554,N_1536);
nand U4297 (N_4297,N_242,N_1903);
and U4298 (N_4298,N_2105,N_1749);
nand U4299 (N_4299,N_1236,N_1021);
or U4300 (N_4300,N_549,N_7);
nand U4301 (N_4301,N_1662,N_2391);
or U4302 (N_4302,N_2367,N_668);
nor U4303 (N_4303,N_1383,N_1660);
and U4304 (N_4304,N_317,N_1565);
nand U4305 (N_4305,N_1906,N_2097);
xnor U4306 (N_4306,N_1658,N_331);
nand U4307 (N_4307,N_2351,N_2467);
nor U4308 (N_4308,N_1014,N_1025);
nand U4309 (N_4309,N_1790,N_1725);
nor U4310 (N_4310,N_249,N_1074);
nand U4311 (N_4311,N_1867,N_943);
or U4312 (N_4312,N_2284,N_1059);
and U4313 (N_4313,N_2391,N_1578);
or U4314 (N_4314,N_2115,N_335);
and U4315 (N_4315,N_1625,N_1301);
or U4316 (N_4316,N_1400,N_221);
nor U4317 (N_4317,N_1855,N_2225);
nor U4318 (N_4318,N_2158,N_564);
and U4319 (N_4319,N_744,N_1787);
nand U4320 (N_4320,N_2042,N_29);
or U4321 (N_4321,N_2125,N_588);
nand U4322 (N_4322,N_1008,N_1855);
nand U4323 (N_4323,N_1274,N_1091);
or U4324 (N_4324,N_854,N_815);
or U4325 (N_4325,N_1110,N_1881);
or U4326 (N_4326,N_139,N_2160);
nor U4327 (N_4327,N_2482,N_1563);
or U4328 (N_4328,N_2457,N_1178);
nand U4329 (N_4329,N_648,N_1958);
nor U4330 (N_4330,N_1138,N_412);
and U4331 (N_4331,N_2129,N_1115);
nor U4332 (N_4332,N_1533,N_1320);
or U4333 (N_4333,N_1274,N_279);
or U4334 (N_4334,N_514,N_2155);
and U4335 (N_4335,N_2011,N_377);
or U4336 (N_4336,N_1917,N_2);
nor U4337 (N_4337,N_2331,N_274);
nand U4338 (N_4338,N_614,N_71);
or U4339 (N_4339,N_1504,N_1758);
nor U4340 (N_4340,N_1715,N_1298);
xnor U4341 (N_4341,N_1329,N_244);
and U4342 (N_4342,N_1755,N_1604);
nand U4343 (N_4343,N_1518,N_1255);
and U4344 (N_4344,N_1576,N_946);
or U4345 (N_4345,N_1490,N_1638);
nor U4346 (N_4346,N_1945,N_1221);
nand U4347 (N_4347,N_716,N_1145);
or U4348 (N_4348,N_1100,N_569);
nor U4349 (N_4349,N_1491,N_1154);
and U4350 (N_4350,N_80,N_77);
or U4351 (N_4351,N_2497,N_1306);
and U4352 (N_4352,N_912,N_1484);
or U4353 (N_4353,N_363,N_395);
or U4354 (N_4354,N_491,N_2175);
nor U4355 (N_4355,N_876,N_700);
and U4356 (N_4356,N_1974,N_105);
or U4357 (N_4357,N_1698,N_1258);
nand U4358 (N_4358,N_1211,N_2230);
nor U4359 (N_4359,N_2295,N_375);
or U4360 (N_4360,N_2497,N_718);
and U4361 (N_4361,N_104,N_2179);
nand U4362 (N_4362,N_649,N_2239);
and U4363 (N_4363,N_1441,N_60);
and U4364 (N_4364,N_335,N_1456);
nor U4365 (N_4365,N_2328,N_1584);
nand U4366 (N_4366,N_1542,N_281);
or U4367 (N_4367,N_1453,N_170);
or U4368 (N_4368,N_932,N_266);
and U4369 (N_4369,N_1291,N_980);
nand U4370 (N_4370,N_767,N_2067);
and U4371 (N_4371,N_409,N_947);
or U4372 (N_4372,N_1496,N_4);
or U4373 (N_4373,N_1740,N_2371);
nor U4374 (N_4374,N_19,N_1856);
or U4375 (N_4375,N_609,N_1039);
nor U4376 (N_4376,N_1510,N_2136);
nand U4377 (N_4377,N_2133,N_1078);
and U4378 (N_4378,N_1463,N_1985);
nand U4379 (N_4379,N_811,N_1483);
xnor U4380 (N_4380,N_1721,N_2223);
nand U4381 (N_4381,N_2445,N_2041);
or U4382 (N_4382,N_855,N_1167);
and U4383 (N_4383,N_2349,N_2095);
or U4384 (N_4384,N_1050,N_1976);
nand U4385 (N_4385,N_2261,N_1083);
xnor U4386 (N_4386,N_613,N_1524);
nor U4387 (N_4387,N_1067,N_558);
or U4388 (N_4388,N_960,N_317);
or U4389 (N_4389,N_1218,N_1203);
nor U4390 (N_4390,N_2306,N_760);
or U4391 (N_4391,N_1667,N_600);
nand U4392 (N_4392,N_1136,N_2166);
and U4393 (N_4393,N_459,N_593);
and U4394 (N_4394,N_1978,N_54);
or U4395 (N_4395,N_134,N_1040);
nor U4396 (N_4396,N_1819,N_922);
nor U4397 (N_4397,N_2196,N_503);
and U4398 (N_4398,N_2172,N_461);
nand U4399 (N_4399,N_2181,N_730);
nand U4400 (N_4400,N_5,N_1826);
or U4401 (N_4401,N_1749,N_296);
nor U4402 (N_4402,N_1905,N_636);
or U4403 (N_4403,N_746,N_2250);
or U4404 (N_4404,N_396,N_1498);
or U4405 (N_4405,N_11,N_185);
nand U4406 (N_4406,N_1832,N_1609);
or U4407 (N_4407,N_1441,N_1737);
or U4408 (N_4408,N_557,N_1765);
nand U4409 (N_4409,N_2207,N_363);
xor U4410 (N_4410,N_970,N_333);
nand U4411 (N_4411,N_1407,N_1658);
and U4412 (N_4412,N_1256,N_2210);
nand U4413 (N_4413,N_1309,N_961);
or U4414 (N_4414,N_462,N_1367);
nand U4415 (N_4415,N_515,N_163);
or U4416 (N_4416,N_2446,N_1676);
nand U4417 (N_4417,N_39,N_1952);
and U4418 (N_4418,N_1805,N_989);
or U4419 (N_4419,N_706,N_1934);
or U4420 (N_4420,N_2487,N_1957);
and U4421 (N_4421,N_667,N_1969);
or U4422 (N_4422,N_2475,N_2103);
nand U4423 (N_4423,N_1558,N_2368);
and U4424 (N_4424,N_631,N_611);
nand U4425 (N_4425,N_467,N_264);
nand U4426 (N_4426,N_565,N_1861);
xnor U4427 (N_4427,N_1464,N_1302);
xor U4428 (N_4428,N_1766,N_1098);
or U4429 (N_4429,N_1550,N_2274);
and U4430 (N_4430,N_2183,N_240);
nor U4431 (N_4431,N_521,N_2323);
nand U4432 (N_4432,N_1809,N_1474);
nor U4433 (N_4433,N_1404,N_338);
nand U4434 (N_4434,N_1844,N_121);
nand U4435 (N_4435,N_276,N_339);
nor U4436 (N_4436,N_531,N_2387);
or U4437 (N_4437,N_1081,N_2175);
nand U4438 (N_4438,N_80,N_1983);
nor U4439 (N_4439,N_302,N_1614);
nand U4440 (N_4440,N_2174,N_952);
nand U4441 (N_4441,N_987,N_1832);
or U4442 (N_4442,N_117,N_550);
or U4443 (N_4443,N_1678,N_1493);
and U4444 (N_4444,N_1416,N_588);
or U4445 (N_4445,N_1027,N_707);
nor U4446 (N_4446,N_814,N_1977);
nor U4447 (N_4447,N_1302,N_351);
nor U4448 (N_4448,N_1858,N_1735);
nor U4449 (N_4449,N_1807,N_2402);
or U4450 (N_4450,N_1573,N_1661);
nand U4451 (N_4451,N_288,N_1561);
or U4452 (N_4452,N_1839,N_2206);
nor U4453 (N_4453,N_280,N_1485);
and U4454 (N_4454,N_466,N_1980);
and U4455 (N_4455,N_0,N_1992);
nor U4456 (N_4456,N_2490,N_621);
and U4457 (N_4457,N_1970,N_435);
nor U4458 (N_4458,N_38,N_2212);
or U4459 (N_4459,N_1506,N_967);
or U4460 (N_4460,N_857,N_1357);
nor U4461 (N_4461,N_417,N_707);
or U4462 (N_4462,N_515,N_1376);
nor U4463 (N_4463,N_598,N_14);
nor U4464 (N_4464,N_1319,N_1964);
nand U4465 (N_4465,N_1056,N_955);
nand U4466 (N_4466,N_1093,N_1336);
nor U4467 (N_4467,N_1038,N_2129);
nor U4468 (N_4468,N_569,N_1278);
nand U4469 (N_4469,N_294,N_1304);
and U4470 (N_4470,N_1129,N_1727);
nor U4471 (N_4471,N_2199,N_946);
nand U4472 (N_4472,N_365,N_132);
nand U4473 (N_4473,N_1626,N_544);
nor U4474 (N_4474,N_1484,N_579);
and U4475 (N_4475,N_293,N_1644);
nor U4476 (N_4476,N_232,N_2139);
or U4477 (N_4477,N_783,N_2326);
nand U4478 (N_4478,N_1070,N_1327);
nand U4479 (N_4479,N_825,N_869);
and U4480 (N_4480,N_1581,N_2289);
nand U4481 (N_4481,N_346,N_2291);
nor U4482 (N_4482,N_1316,N_1351);
nor U4483 (N_4483,N_145,N_1823);
nand U4484 (N_4484,N_335,N_2251);
and U4485 (N_4485,N_722,N_485);
nand U4486 (N_4486,N_138,N_2310);
or U4487 (N_4487,N_2469,N_719);
xor U4488 (N_4488,N_2019,N_893);
nand U4489 (N_4489,N_189,N_1684);
nand U4490 (N_4490,N_1945,N_204);
nand U4491 (N_4491,N_181,N_440);
nand U4492 (N_4492,N_653,N_2434);
nor U4493 (N_4493,N_1303,N_1759);
or U4494 (N_4494,N_1887,N_686);
nor U4495 (N_4495,N_2498,N_551);
or U4496 (N_4496,N_1864,N_236);
nand U4497 (N_4497,N_874,N_2294);
nor U4498 (N_4498,N_936,N_2173);
nor U4499 (N_4499,N_1875,N_1994);
or U4500 (N_4500,N_254,N_365);
nand U4501 (N_4501,N_71,N_2483);
nor U4502 (N_4502,N_1583,N_2242);
nand U4503 (N_4503,N_2448,N_1466);
nor U4504 (N_4504,N_281,N_1831);
nand U4505 (N_4505,N_1786,N_2304);
and U4506 (N_4506,N_1143,N_321);
nor U4507 (N_4507,N_283,N_1725);
nand U4508 (N_4508,N_713,N_1319);
nand U4509 (N_4509,N_1084,N_2077);
and U4510 (N_4510,N_2287,N_1279);
and U4511 (N_4511,N_2128,N_492);
and U4512 (N_4512,N_1808,N_514);
and U4513 (N_4513,N_1959,N_233);
nand U4514 (N_4514,N_1892,N_70);
and U4515 (N_4515,N_1616,N_685);
nor U4516 (N_4516,N_724,N_866);
nand U4517 (N_4517,N_2162,N_2302);
and U4518 (N_4518,N_1941,N_1891);
or U4519 (N_4519,N_35,N_474);
or U4520 (N_4520,N_678,N_490);
nor U4521 (N_4521,N_502,N_2440);
nand U4522 (N_4522,N_2353,N_1267);
nand U4523 (N_4523,N_1105,N_135);
and U4524 (N_4524,N_592,N_1063);
and U4525 (N_4525,N_488,N_852);
or U4526 (N_4526,N_2450,N_2392);
nor U4527 (N_4527,N_497,N_1684);
or U4528 (N_4528,N_1897,N_1296);
nor U4529 (N_4529,N_2214,N_1334);
nor U4530 (N_4530,N_1320,N_629);
and U4531 (N_4531,N_2222,N_2389);
and U4532 (N_4532,N_2044,N_2076);
or U4533 (N_4533,N_2192,N_1690);
nand U4534 (N_4534,N_2340,N_833);
nand U4535 (N_4535,N_944,N_873);
nand U4536 (N_4536,N_972,N_261);
or U4537 (N_4537,N_582,N_2123);
nor U4538 (N_4538,N_67,N_955);
nor U4539 (N_4539,N_846,N_202);
nand U4540 (N_4540,N_242,N_94);
or U4541 (N_4541,N_625,N_2076);
nand U4542 (N_4542,N_1562,N_2083);
or U4543 (N_4543,N_1482,N_1763);
xor U4544 (N_4544,N_2173,N_455);
and U4545 (N_4545,N_874,N_2247);
nor U4546 (N_4546,N_1327,N_1897);
nor U4547 (N_4547,N_1347,N_886);
and U4548 (N_4548,N_305,N_891);
and U4549 (N_4549,N_2177,N_1016);
nor U4550 (N_4550,N_2403,N_1606);
or U4551 (N_4551,N_1580,N_1241);
nand U4552 (N_4552,N_1309,N_801);
and U4553 (N_4553,N_358,N_2471);
or U4554 (N_4554,N_938,N_1492);
nand U4555 (N_4555,N_1775,N_1893);
nand U4556 (N_4556,N_1681,N_329);
and U4557 (N_4557,N_1217,N_92);
nand U4558 (N_4558,N_312,N_1735);
nor U4559 (N_4559,N_1580,N_2443);
nor U4560 (N_4560,N_2077,N_343);
and U4561 (N_4561,N_2335,N_77);
nor U4562 (N_4562,N_1078,N_1522);
and U4563 (N_4563,N_848,N_2073);
nand U4564 (N_4564,N_890,N_960);
or U4565 (N_4565,N_1401,N_636);
nand U4566 (N_4566,N_2009,N_2462);
or U4567 (N_4567,N_1487,N_2289);
nor U4568 (N_4568,N_967,N_1120);
and U4569 (N_4569,N_319,N_198);
nor U4570 (N_4570,N_950,N_1472);
nand U4571 (N_4571,N_1107,N_639);
or U4572 (N_4572,N_2183,N_2448);
nor U4573 (N_4573,N_2325,N_592);
nor U4574 (N_4574,N_2484,N_948);
and U4575 (N_4575,N_2068,N_2387);
nand U4576 (N_4576,N_788,N_1122);
nor U4577 (N_4577,N_1308,N_1267);
or U4578 (N_4578,N_2248,N_1097);
nor U4579 (N_4579,N_2115,N_2002);
nor U4580 (N_4580,N_1130,N_2201);
and U4581 (N_4581,N_1244,N_1204);
nor U4582 (N_4582,N_2025,N_17);
nor U4583 (N_4583,N_1376,N_898);
and U4584 (N_4584,N_1959,N_188);
nand U4585 (N_4585,N_225,N_888);
and U4586 (N_4586,N_601,N_1932);
nand U4587 (N_4587,N_1301,N_83);
or U4588 (N_4588,N_2301,N_539);
and U4589 (N_4589,N_1487,N_2012);
nand U4590 (N_4590,N_726,N_87);
nand U4591 (N_4591,N_2400,N_480);
nor U4592 (N_4592,N_1415,N_2366);
nand U4593 (N_4593,N_2238,N_1672);
nand U4594 (N_4594,N_1448,N_1904);
or U4595 (N_4595,N_554,N_2002);
and U4596 (N_4596,N_1536,N_1663);
or U4597 (N_4597,N_2259,N_650);
and U4598 (N_4598,N_1984,N_1643);
nand U4599 (N_4599,N_720,N_99);
and U4600 (N_4600,N_648,N_1107);
and U4601 (N_4601,N_104,N_386);
nor U4602 (N_4602,N_1608,N_978);
nand U4603 (N_4603,N_1135,N_540);
nor U4604 (N_4604,N_34,N_770);
nor U4605 (N_4605,N_1591,N_1963);
nor U4606 (N_4606,N_1827,N_1775);
nor U4607 (N_4607,N_1331,N_2058);
nand U4608 (N_4608,N_1850,N_2477);
nand U4609 (N_4609,N_2475,N_501);
and U4610 (N_4610,N_42,N_762);
and U4611 (N_4611,N_488,N_2305);
and U4612 (N_4612,N_1943,N_43);
or U4613 (N_4613,N_2221,N_1112);
and U4614 (N_4614,N_1221,N_761);
nor U4615 (N_4615,N_624,N_953);
and U4616 (N_4616,N_259,N_1985);
nor U4617 (N_4617,N_773,N_1579);
nand U4618 (N_4618,N_2297,N_2141);
or U4619 (N_4619,N_1713,N_1145);
nand U4620 (N_4620,N_2355,N_1985);
xor U4621 (N_4621,N_1831,N_651);
nor U4622 (N_4622,N_1931,N_1364);
and U4623 (N_4623,N_1656,N_371);
nor U4624 (N_4624,N_2468,N_1167);
nand U4625 (N_4625,N_232,N_1323);
nor U4626 (N_4626,N_561,N_1574);
and U4627 (N_4627,N_632,N_1330);
nand U4628 (N_4628,N_158,N_307);
nand U4629 (N_4629,N_2456,N_220);
nand U4630 (N_4630,N_2290,N_2408);
nor U4631 (N_4631,N_898,N_2352);
and U4632 (N_4632,N_1973,N_493);
nor U4633 (N_4633,N_1411,N_1739);
xor U4634 (N_4634,N_226,N_727);
nand U4635 (N_4635,N_782,N_1454);
nor U4636 (N_4636,N_814,N_195);
or U4637 (N_4637,N_2004,N_3);
and U4638 (N_4638,N_2306,N_1889);
and U4639 (N_4639,N_1553,N_1301);
nand U4640 (N_4640,N_235,N_2211);
nand U4641 (N_4641,N_2096,N_1979);
or U4642 (N_4642,N_304,N_95);
nand U4643 (N_4643,N_2146,N_1109);
nand U4644 (N_4644,N_1443,N_71);
or U4645 (N_4645,N_1676,N_2383);
nor U4646 (N_4646,N_2166,N_268);
nand U4647 (N_4647,N_770,N_876);
or U4648 (N_4648,N_590,N_1100);
and U4649 (N_4649,N_245,N_676);
nor U4650 (N_4650,N_2288,N_2056);
and U4651 (N_4651,N_778,N_1144);
and U4652 (N_4652,N_140,N_1566);
nand U4653 (N_4653,N_2359,N_1908);
nor U4654 (N_4654,N_1446,N_862);
or U4655 (N_4655,N_1685,N_1353);
or U4656 (N_4656,N_1091,N_604);
nand U4657 (N_4657,N_594,N_696);
or U4658 (N_4658,N_1939,N_297);
nand U4659 (N_4659,N_89,N_1334);
nor U4660 (N_4660,N_1203,N_2386);
and U4661 (N_4661,N_1683,N_1113);
nand U4662 (N_4662,N_2130,N_2297);
nor U4663 (N_4663,N_1285,N_330);
or U4664 (N_4664,N_2323,N_1170);
or U4665 (N_4665,N_853,N_2157);
and U4666 (N_4666,N_1621,N_892);
and U4667 (N_4667,N_1495,N_1128);
nand U4668 (N_4668,N_1551,N_1022);
nand U4669 (N_4669,N_2052,N_1798);
or U4670 (N_4670,N_2029,N_1746);
and U4671 (N_4671,N_1991,N_1120);
and U4672 (N_4672,N_103,N_1395);
or U4673 (N_4673,N_2429,N_1691);
and U4674 (N_4674,N_491,N_1014);
nor U4675 (N_4675,N_1582,N_2308);
or U4676 (N_4676,N_1722,N_1081);
nand U4677 (N_4677,N_1832,N_184);
nand U4678 (N_4678,N_928,N_391);
nor U4679 (N_4679,N_293,N_1823);
nand U4680 (N_4680,N_1051,N_172);
nor U4681 (N_4681,N_944,N_1241);
nand U4682 (N_4682,N_520,N_1530);
or U4683 (N_4683,N_296,N_639);
nor U4684 (N_4684,N_2038,N_2389);
nor U4685 (N_4685,N_1738,N_1734);
nand U4686 (N_4686,N_2197,N_1071);
or U4687 (N_4687,N_61,N_1604);
nand U4688 (N_4688,N_399,N_2332);
nor U4689 (N_4689,N_1068,N_2431);
nand U4690 (N_4690,N_2453,N_1452);
and U4691 (N_4691,N_2396,N_945);
and U4692 (N_4692,N_2249,N_405);
nand U4693 (N_4693,N_4,N_1);
and U4694 (N_4694,N_1115,N_228);
or U4695 (N_4695,N_12,N_856);
and U4696 (N_4696,N_589,N_546);
nand U4697 (N_4697,N_2439,N_1058);
nor U4698 (N_4698,N_891,N_301);
nor U4699 (N_4699,N_642,N_1057);
nand U4700 (N_4700,N_1272,N_454);
nor U4701 (N_4701,N_895,N_1370);
and U4702 (N_4702,N_375,N_457);
and U4703 (N_4703,N_109,N_1772);
or U4704 (N_4704,N_600,N_1813);
nor U4705 (N_4705,N_1246,N_562);
nand U4706 (N_4706,N_1561,N_642);
and U4707 (N_4707,N_385,N_2105);
and U4708 (N_4708,N_1555,N_628);
nor U4709 (N_4709,N_1677,N_1469);
and U4710 (N_4710,N_1299,N_2333);
or U4711 (N_4711,N_2281,N_1191);
and U4712 (N_4712,N_1153,N_2219);
or U4713 (N_4713,N_2070,N_1532);
nand U4714 (N_4714,N_350,N_20);
or U4715 (N_4715,N_2104,N_1355);
xnor U4716 (N_4716,N_874,N_2157);
xor U4717 (N_4717,N_2015,N_1625);
nor U4718 (N_4718,N_2350,N_1195);
or U4719 (N_4719,N_800,N_460);
nand U4720 (N_4720,N_902,N_1171);
and U4721 (N_4721,N_1214,N_1488);
nand U4722 (N_4722,N_1023,N_227);
or U4723 (N_4723,N_1518,N_2404);
and U4724 (N_4724,N_597,N_1413);
or U4725 (N_4725,N_2177,N_2374);
and U4726 (N_4726,N_898,N_274);
nor U4727 (N_4727,N_2199,N_1963);
and U4728 (N_4728,N_2452,N_1767);
nand U4729 (N_4729,N_189,N_1437);
xor U4730 (N_4730,N_1243,N_2026);
and U4731 (N_4731,N_275,N_1706);
nand U4732 (N_4732,N_1573,N_838);
or U4733 (N_4733,N_168,N_2315);
or U4734 (N_4734,N_789,N_781);
and U4735 (N_4735,N_1610,N_2363);
nor U4736 (N_4736,N_143,N_179);
nand U4737 (N_4737,N_1637,N_653);
or U4738 (N_4738,N_1144,N_2203);
and U4739 (N_4739,N_1825,N_927);
and U4740 (N_4740,N_1511,N_2481);
nor U4741 (N_4741,N_1160,N_1050);
and U4742 (N_4742,N_1346,N_2172);
or U4743 (N_4743,N_2445,N_114);
and U4744 (N_4744,N_2095,N_1880);
nand U4745 (N_4745,N_1974,N_1064);
or U4746 (N_4746,N_1377,N_1952);
or U4747 (N_4747,N_62,N_602);
or U4748 (N_4748,N_652,N_2331);
and U4749 (N_4749,N_669,N_1214);
nand U4750 (N_4750,N_2072,N_1747);
nand U4751 (N_4751,N_1239,N_2060);
or U4752 (N_4752,N_1380,N_2271);
nor U4753 (N_4753,N_1047,N_221);
and U4754 (N_4754,N_89,N_255);
nor U4755 (N_4755,N_620,N_1006);
or U4756 (N_4756,N_1558,N_910);
nand U4757 (N_4757,N_157,N_951);
nor U4758 (N_4758,N_223,N_2129);
and U4759 (N_4759,N_1571,N_2077);
or U4760 (N_4760,N_1260,N_1364);
nand U4761 (N_4761,N_26,N_378);
nor U4762 (N_4762,N_1785,N_1512);
nor U4763 (N_4763,N_926,N_2363);
and U4764 (N_4764,N_1511,N_1577);
and U4765 (N_4765,N_2357,N_865);
and U4766 (N_4766,N_643,N_1824);
and U4767 (N_4767,N_2356,N_1216);
or U4768 (N_4768,N_587,N_983);
xnor U4769 (N_4769,N_1959,N_221);
nand U4770 (N_4770,N_452,N_386);
or U4771 (N_4771,N_2408,N_95);
or U4772 (N_4772,N_2453,N_898);
or U4773 (N_4773,N_816,N_2045);
nand U4774 (N_4774,N_2024,N_509);
nand U4775 (N_4775,N_1238,N_1089);
or U4776 (N_4776,N_1619,N_2013);
nor U4777 (N_4777,N_1031,N_767);
or U4778 (N_4778,N_2092,N_1058);
nor U4779 (N_4779,N_883,N_1878);
or U4780 (N_4780,N_413,N_2224);
nand U4781 (N_4781,N_1877,N_2364);
and U4782 (N_4782,N_2340,N_2370);
and U4783 (N_4783,N_1884,N_122);
or U4784 (N_4784,N_1342,N_545);
nand U4785 (N_4785,N_122,N_1794);
or U4786 (N_4786,N_1425,N_124);
nor U4787 (N_4787,N_2200,N_1368);
or U4788 (N_4788,N_1344,N_165);
and U4789 (N_4789,N_2089,N_1614);
nand U4790 (N_4790,N_57,N_913);
or U4791 (N_4791,N_375,N_1016);
nor U4792 (N_4792,N_2158,N_1233);
nand U4793 (N_4793,N_337,N_1844);
and U4794 (N_4794,N_800,N_1067);
nor U4795 (N_4795,N_1840,N_792);
and U4796 (N_4796,N_641,N_2422);
or U4797 (N_4797,N_606,N_2426);
nor U4798 (N_4798,N_435,N_617);
nand U4799 (N_4799,N_110,N_2234);
nand U4800 (N_4800,N_1510,N_1629);
and U4801 (N_4801,N_2262,N_815);
or U4802 (N_4802,N_2120,N_2099);
and U4803 (N_4803,N_995,N_1217);
nor U4804 (N_4804,N_773,N_2278);
and U4805 (N_4805,N_1675,N_2325);
or U4806 (N_4806,N_241,N_1006);
or U4807 (N_4807,N_1777,N_800);
nand U4808 (N_4808,N_648,N_1861);
or U4809 (N_4809,N_1422,N_2027);
xnor U4810 (N_4810,N_2095,N_150);
and U4811 (N_4811,N_2157,N_1831);
or U4812 (N_4812,N_1988,N_32);
nand U4813 (N_4813,N_2283,N_623);
nor U4814 (N_4814,N_1319,N_2064);
nor U4815 (N_4815,N_1544,N_1041);
and U4816 (N_4816,N_122,N_498);
nand U4817 (N_4817,N_561,N_1867);
nand U4818 (N_4818,N_1892,N_1620);
and U4819 (N_4819,N_1118,N_608);
or U4820 (N_4820,N_156,N_1734);
nand U4821 (N_4821,N_1236,N_2310);
nor U4822 (N_4822,N_1141,N_1133);
or U4823 (N_4823,N_2025,N_142);
nand U4824 (N_4824,N_759,N_2076);
or U4825 (N_4825,N_1674,N_2373);
nand U4826 (N_4826,N_525,N_2490);
and U4827 (N_4827,N_2231,N_515);
or U4828 (N_4828,N_955,N_812);
nand U4829 (N_4829,N_349,N_1211);
nand U4830 (N_4830,N_1350,N_1563);
nand U4831 (N_4831,N_696,N_1561);
nand U4832 (N_4832,N_27,N_1677);
nand U4833 (N_4833,N_231,N_2281);
and U4834 (N_4834,N_1184,N_1950);
or U4835 (N_4835,N_318,N_649);
nand U4836 (N_4836,N_1237,N_1738);
nor U4837 (N_4837,N_41,N_2091);
xnor U4838 (N_4838,N_440,N_1007);
and U4839 (N_4839,N_851,N_1314);
and U4840 (N_4840,N_1576,N_643);
or U4841 (N_4841,N_2421,N_890);
and U4842 (N_4842,N_15,N_264);
and U4843 (N_4843,N_1260,N_396);
nand U4844 (N_4844,N_734,N_2016);
xnor U4845 (N_4845,N_58,N_202);
or U4846 (N_4846,N_1748,N_1185);
or U4847 (N_4847,N_2048,N_2000);
or U4848 (N_4848,N_1337,N_1165);
nand U4849 (N_4849,N_608,N_765);
nand U4850 (N_4850,N_2020,N_1256);
nand U4851 (N_4851,N_1377,N_1047);
or U4852 (N_4852,N_1551,N_2130);
nand U4853 (N_4853,N_1810,N_323);
and U4854 (N_4854,N_1129,N_403);
nand U4855 (N_4855,N_958,N_2384);
or U4856 (N_4856,N_2268,N_2010);
nand U4857 (N_4857,N_1438,N_1452);
nand U4858 (N_4858,N_2255,N_154);
nand U4859 (N_4859,N_1249,N_159);
nor U4860 (N_4860,N_39,N_778);
nand U4861 (N_4861,N_1598,N_2165);
and U4862 (N_4862,N_203,N_2345);
or U4863 (N_4863,N_412,N_497);
nor U4864 (N_4864,N_2230,N_1523);
and U4865 (N_4865,N_1054,N_2286);
and U4866 (N_4866,N_401,N_2266);
nor U4867 (N_4867,N_817,N_590);
nand U4868 (N_4868,N_1100,N_2411);
and U4869 (N_4869,N_1864,N_2152);
nand U4870 (N_4870,N_1701,N_594);
nand U4871 (N_4871,N_2322,N_410);
or U4872 (N_4872,N_1063,N_1811);
nor U4873 (N_4873,N_825,N_2486);
nor U4874 (N_4874,N_153,N_366);
nor U4875 (N_4875,N_1385,N_2303);
nand U4876 (N_4876,N_339,N_1625);
nand U4877 (N_4877,N_2378,N_1307);
and U4878 (N_4878,N_1881,N_657);
or U4879 (N_4879,N_1999,N_700);
and U4880 (N_4880,N_440,N_731);
and U4881 (N_4881,N_473,N_2203);
nor U4882 (N_4882,N_752,N_790);
or U4883 (N_4883,N_780,N_2197);
nor U4884 (N_4884,N_74,N_60);
and U4885 (N_4885,N_1146,N_1732);
xor U4886 (N_4886,N_489,N_1659);
nor U4887 (N_4887,N_2352,N_811);
nand U4888 (N_4888,N_1262,N_694);
nor U4889 (N_4889,N_1751,N_166);
nor U4890 (N_4890,N_901,N_912);
and U4891 (N_4891,N_1472,N_2422);
nor U4892 (N_4892,N_1884,N_1548);
or U4893 (N_4893,N_1064,N_1933);
nand U4894 (N_4894,N_1644,N_2458);
xor U4895 (N_4895,N_154,N_1202);
or U4896 (N_4896,N_2331,N_109);
nand U4897 (N_4897,N_561,N_654);
nand U4898 (N_4898,N_1264,N_1455);
nor U4899 (N_4899,N_2355,N_2019);
nor U4900 (N_4900,N_883,N_1484);
nand U4901 (N_4901,N_1020,N_929);
or U4902 (N_4902,N_92,N_1372);
or U4903 (N_4903,N_56,N_2083);
and U4904 (N_4904,N_1167,N_822);
or U4905 (N_4905,N_1218,N_2207);
nor U4906 (N_4906,N_2326,N_1120);
nand U4907 (N_4907,N_1279,N_1024);
or U4908 (N_4908,N_1336,N_168);
and U4909 (N_4909,N_1535,N_2045);
nand U4910 (N_4910,N_1199,N_873);
nand U4911 (N_4911,N_1965,N_139);
nor U4912 (N_4912,N_1970,N_1644);
and U4913 (N_4913,N_820,N_1623);
and U4914 (N_4914,N_2262,N_2284);
or U4915 (N_4915,N_420,N_2220);
or U4916 (N_4916,N_741,N_2280);
or U4917 (N_4917,N_332,N_613);
nand U4918 (N_4918,N_788,N_1235);
and U4919 (N_4919,N_726,N_1443);
or U4920 (N_4920,N_637,N_915);
nor U4921 (N_4921,N_1293,N_807);
nand U4922 (N_4922,N_1007,N_1830);
nor U4923 (N_4923,N_214,N_326);
nor U4924 (N_4924,N_1397,N_1144);
nor U4925 (N_4925,N_1981,N_2438);
or U4926 (N_4926,N_1995,N_1756);
and U4927 (N_4927,N_2112,N_1728);
nor U4928 (N_4928,N_691,N_2161);
nor U4929 (N_4929,N_90,N_903);
nand U4930 (N_4930,N_980,N_1771);
nor U4931 (N_4931,N_2295,N_344);
nand U4932 (N_4932,N_1714,N_239);
nand U4933 (N_4933,N_1408,N_1819);
and U4934 (N_4934,N_920,N_329);
or U4935 (N_4935,N_122,N_1844);
nand U4936 (N_4936,N_2107,N_113);
or U4937 (N_4937,N_929,N_1793);
or U4938 (N_4938,N_2353,N_2178);
and U4939 (N_4939,N_1868,N_520);
nor U4940 (N_4940,N_595,N_988);
and U4941 (N_4941,N_1399,N_125);
or U4942 (N_4942,N_1717,N_461);
and U4943 (N_4943,N_885,N_2401);
or U4944 (N_4944,N_1232,N_561);
nor U4945 (N_4945,N_195,N_210);
or U4946 (N_4946,N_2021,N_2195);
or U4947 (N_4947,N_340,N_1841);
and U4948 (N_4948,N_100,N_1771);
and U4949 (N_4949,N_622,N_895);
nand U4950 (N_4950,N_2205,N_1293);
and U4951 (N_4951,N_1015,N_582);
or U4952 (N_4952,N_374,N_1938);
or U4953 (N_4953,N_2117,N_939);
nor U4954 (N_4954,N_2498,N_1591);
and U4955 (N_4955,N_218,N_2062);
nor U4956 (N_4956,N_1263,N_233);
nor U4957 (N_4957,N_1461,N_742);
and U4958 (N_4958,N_1406,N_600);
and U4959 (N_4959,N_363,N_1799);
nand U4960 (N_4960,N_828,N_1913);
and U4961 (N_4961,N_958,N_1965);
and U4962 (N_4962,N_98,N_89);
nand U4963 (N_4963,N_1301,N_798);
nand U4964 (N_4964,N_2441,N_2424);
and U4965 (N_4965,N_673,N_2367);
nor U4966 (N_4966,N_369,N_1063);
nor U4967 (N_4967,N_666,N_1271);
nor U4968 (N_4968,N_2070,N_2445);
nand U4969 (N_4969,N_158,N_402);
nor U4970 (N_4970,N_1856,N_600);
nor U4971 (N_4971,N_141,N_2286);
or U4972 (N_4972,N_1769,N_507);
nand U4973 (N_4973,N_716,N_2499);
and U4974 (N_4974,N_494,N_2498);
or U4975 (N_4975,N_2376,N_1926);
or U4976 (N_4976,N_1596,N_1073);
nor U4977 (N_4977,N_1498,N_584);
nor U4978 (N_4978,N_2208,N_1155);
nand U4979 (N_4979,N_1004,N_240);
nor U4980 (N_4980,N_835,N_661);
or U4981 (N_4981,N_1339,N_143);
and U4982 (N_4982,N_1978,N_1340);
and U4983 (N_4983,N_1290,N_875);
or U4984 (N_4984,N_2448,N_1408);
or U4985 (N_4985,N_2351,N_1546);
nor U4986 (N_4986,N_117,N_985);
and U4987 (N_4987,N_70,N_2302);
nor U4988 (N_4988,N_1701,N_634);
nand U4989 (N_4989,N_1995,N_2194);
and U4990 (N_4990,N_7,N_477);
or U4991 (N_4991,N_763,N_1252);
or U4992 (N_4992,N_830,N_1520);
nor U4993 (N_4993,N_2452,N_582);
and U4994 (N_4994,N_2069,N_1530);
or U4995 (N_4995,N_922,N_492);
and U4996 (N_4996,N_1365,N_1950);
nor U4997 (N_4997,N_518,N_2339);
or U4998 (N_4998,N_2187,N_476);
and U4999 (N_4999,N_1071,N_48);
nand U5000 (N_5000,N_4160,N_3935);
nor U5001 (N_5001,N_2891,N_3006);
or U5002 (N_5002,N_4824,N_2912);
or U5003 (N_5003,N_4293,N_3863);
nor U5004 (N_5004,N_2639,N_4487);
nor U5005 (N_5005,N_4357,N_3316);
and U5006 (N_5006,N_3434,N_3119);
or U5007 (N_5007,N_4910,N_2704);
nor U5008 (N_5008,N_4673,N_2899);
nand U5009 (N_5009,N_3718,N_3344);
and U5010 (N_5010,N_3491,N_4970);
nand U5011 (N_5011,N_4256,N_3810);
nor U5012 (N_5012,N_4564,N_3276);
or U5013 (N_5013,N_4609,N_3661);
and U5014 (N_5014,N_3297,N_3025);
nand U5015 (N_5015,N_2719,N_3280);
and U5016 (N_5016,N_3027,N_4045);
nor U5017 (N_5017,N_3860,N_2943);
nor U5018 (N_5018,N_4126,N_4375);
nor U5019 (N_5019,N_3263,N_3789);
nand U5020 (N_5020,N_3412,N_4087);
nor U5021 (N_5021,N_4806,N_4592);
and U5022 (N_5022,N_4081,N_4645);
nand U5023 (N_5023,N_3552,N_2625);
and U5024 (N_5024,N_4600,N_3533);
or U5025 (N_5025,N_4103,N_3864);
and U5026 (N_5026,N_3882,N_3506);
or U5027 (N_5027,N_2974,N_4775);
nor U5028 (N_5028,N_4234,N_4577);
nand U5029 (N_5029,N_3107,N_3646);
xor U5030 (N_5030,N_3975,N_3912);
or U5031 (N_5031,N_3854,N_4504);
nand U5032 (N_5032,N_3971,N_3629);
and U5033 (N_5033,N_2699,N_3607);
nor U5034 (N_5034,N_2663,N_4952);
and U5035 (N_5035,N_3139,N_4951);
nor U5036 (N_5036,N_3869,N_4988);
nor U5037 (N_5037,N_3132,N_4248);
nand U5038 (N_5038,N_2695,N_4532);
or U5039 (N_5039,N_2881,N_3505);
or U5040 (N_5040,N_4031,N_4555);
or U5041 (N_5041,N_3560,N_3940);
nand U5042 (N_5042,N_4080,N_4557);
and U5043 (N_5043,N_3362,N_3813);
nor U5044 (N_5044,N_3191,N_2722);
nand U5045 (N_5045,N_4815,N_3787);
nor U5046 (N_5046,N_2817,N_4434);
or U5047 (N_5047,N_4613,N_3063);
and U5048 (N_5048,N_3739,N_2981);
nand U5049 (N_5049,N_3140,N_4595);
nor U5050 (N_5050,N_2933,N_3977);
and U5051 (N_5051,N_3701,N_3488);
and U5052 (N_5052,N_4164,N_3618);
and U5053 (N_5053,N_3407,N_3074);
nor U5054 (N_5054,N_3414,N_3193);
nand U5055 (N_5055,N_3853,N_3990);
and U5056 (N_5056,N_4721,N_3157);
nor U5057 (N_5057,N_3396,N_4314);
nor U5058 (N_5058,N_3167,N_2617);
nand U5059 (N_5059,N_3038,N_2872);
or U5060 (N_5060,N_3928,N_4849);
nor U5061 (N_5061,N_2725,N_3720);
or U5062 (N_5062,N_4127,N_4701);
nand U5063 (N_5063,N_4911,N_3313);
and U5064 (N_5064,N_3921,N_3002);
nand U5065 (N_5065,N_3775,N_3382);
or U5066 (N_5066,N_4455,N_4723);
or U5067 (N_5067,N_3911,N_4887);
nor U5068 (N_5068,N_4593,N_4979);
nand U5069 (N_5069,N_2877,N_4678);
nor U5070 (N_5070,N_4128,N_2917);
nor U5071 (N_5071,N_3965,N_4451);
and U5072 (N_5072,N_4840,N_3647);
or U5073 (N_5073,N_3166,N_4920);
and U5074 (N_5074,N_4236,N_4400);
and U5075 (N_5075,N_2714,N_4744);
and U5076 (N_5076,N_3423,N_4832);
nand U5077 (N_5077,N_4757,N_3530);
nor U5078 (N_5078,N_4756,N_2653);
and U5079 (N_5079,N_3780,N_3648);
or U5080 (N_5080,N_3808,N_4471);
and U5081 (N_5081,N_2800,N_4518);
and U5082 (N_5082,N_2721,N_3405);
and U5083 (N_5083,N_4627,N_4218);
and U5084 (N_5084,N_4318,N_3689);
nor U5085 (N_5085,N_4065,N_2735);
or U5086 (N_5086,N_3746,N_3399);
nand U5087 (N_5087,N_4618,N_3576);
nand U5088 (N_5088,N_3600,N_2772);
and U5089 (N_5089,N_2511,N_2675);
and U5090 (N_5090,N_4215,N_3218);
or U5091 (N_5091,N_2977,N_4221);
and U5092 (N_5092,N_4254,N_4591);
or U5093 (N_5093,N_3814,N_4262);
or U5094 (N_5094,N_4120,N_2835);
nor U5095 (N_5095,N_4583,N_4766);
or U5096 (N_5096,N_3541,N_3499);
nand U5097 (N_5097,N_3080,N_2757);
nand U5098 (N_5098,N_4008,N_4149);
and U5099 (N_5099,N_3788,N_4559);
nor U5100 (N_5100,N_4538,N_4580);
nand U5101 (N_5101,N_3667,N_4790);
nand U5102 (N_5102,N_4829,N_4453);
or U5103 (N_5103,N_3699,N_4855);
nor U5104 (N_5104,N_2765,N_4190);
and U5105 (N_5105,N_4542,N_3807);
and U5106 (N_5106,N_2551,N_2698);
nand U5107 (N_5107,N_4468,N_2586);
or U5108 (N_5108,N_4469,N_3244);
and U5109 (N_5109,N_3302,N_4888);
and U5110 (N_5110,N_3039,N_4093);
nor U5111 (N_5111,N_3142,N_4179);
and U5112 (N_5112,N_2578,N_4977);
and U5113 (N_5113,N_4095,N_2746);
nor U5114 (N_5114,N_3246,N_2686);
nor U5115 (N_5115,N_4937,N_4478);
nor U5116 (N_5116,N_2611,N_3724);
nor U5117 (N_5117,N_3388,N_3816);
and U5118 (N_5118,N_3534,N_3418);
nand U5119 (N_5119,N_2613,N_4411);
or U5120 (N_5120,N_3137,N_4841);
and U5121 (N_5121,N_4116,N_4308);
nand U5122 (N_5122,N_2821,N_4019);
or U5123 (N_5123,N_2650,N_4602);
nor U5124 (N_5124,N_4147,N_3984);
nor U5125 (N_5125,N_2608,N_3351);
nand U5126 (N_5126,N_4989,N_2736);
or U5127 (N_5127,N_4783,N_3563);
and U5128 (N_5128,N_4522,N_3252);
nor U5129 (N_5129,N_4251,N_3215);
or U5130 (N_5130,N_4477,N_3722);
nor U5131 (N_5131,N_3893,N_3517);
nor U5132 (N_5132,N_4519,N_2709);
nand U5133 (N_5133,N_2789,N_3073);
and U5134 (N_5134,N_3035,N_4068);
and U5135 (N_5135,N_3426,N_3852);
nand U5136 (N_5136,N_3374,N_4607);
nand U5137 (N_5137,N_4804,N_4803);
and U5138 (N_5138,N_2681,N_4183);
xor U5139 (N_5139,N_4684,N_2598);
nor U5140 (N_5140,N_4524,N_3309);
and U5141 (N_5141,N_4188,N_4282);
nand U5142 (N_5142,N_2667,N_2702);
or U5143 (N_5143,N_3709,N_4791);
nand U5144 (N_5144,N_3695,N_4596);
nor U5145 (N_5145,N_4525,N_3637);
nor U5146 (N_5146,N_4245,N_2655);
nor U5147 (N_5147,N_3120,N_3470);
nor U5148 (N_5148,N_3029,N_2590);
nand U5149 (N_5149,N_2954,N_3945);
or U5150 (N_5150,N_3992,N_3239);
nand U5151 (N_5151,N_4101,N_3196);
or U5152 (N_5152,N_2979,N_4091);
or U5153 (N_5153,N_4397,N_3105);
or U5154 (N_5154,N_4792,N_3703);
and U5155 (N_5155,N_3043,N_2542);
nand U5156 (N_5156,N_3118,N_2787);
nor U5157 (N_5157,N_3778,N_4422);
and U5158 (N_5158,N_3832,N_2972);
nand U5159 (N_5159,N_3324,N_4007);
or U5160 (N_5160,N_3444,N_3273);
and U5161 (N_5161,N_4482,N_3230);
or U5162 (N_5162,N_4848,N_4754);
nand U5163 (N_5163,N_4717,N_2701);
and U5164 (N_5164,N_4764,N_4612);
nor U5165 (N_5165,N_4125,N_4208);
or U5166 (N_5166,N_4305,N_4941);
nor U5167 (N_5167,N_2514,N_4452);
and U5168 (N_5168,N_3796,N_2993);
nand U5169 (N_5169,N_4294,N_4856);
nand U5170 (N_5170,N_2642,N_3494);
nor U5171 (N_5171,N_3201,N_3512);
or U5172 (N_5172,N_3758,N_3602);
or U5173 (N_5173,N_3500,N_4528);
or U5174 (N_5174,N_3420,N_3985);
nand U5175 (N_5175,N_2875,N_4533);
nor U5176 (N_5176,N_2846,N_4785);
nor U5177 (N_5177,N_4939,N_2637);
nor U5178 (N_5178,N_4996,N_3031);
or U5179 (N_5179,N_4745,N_3266);
nand U5180 (N_5180,N_4277,N_3820);
nand U5181 (N_5181,N_3259,N_2518);
and U5182 (N_5182,N_4074,N_2530);
and U5183 (N_5183,N_4707,N_4635);
nand U5184 (N_5184,N_4648,N_3180);
nor U5185 (N_5185,N_3149,N_4664);
nand U5186 (N_5186,N_3819,N_3200);
nor U5187 (N_5187,N_4644,N_2706);
and U5188 (N_5188,N_3842,N_3152);
nor U5189 (N_5189,N_2873,N_3472);
nand U5190 (N_5190,N_4110,N_3238);
and U5191 (N_5191,N_3123,N_2963);
nor U5192 (N_5192,N_2842,N_3183);
nand U5193 (N_5193,N_3631,N_3906);
nand U5194 (N_5194,N_4017,N_2643);
and U5195 (N_5195,N_3665,N_4874);
xnor U5196 (N_5196,N_3130,N_3584);
nand U5197 (N_5197,N_3331,N_3871);
or U5198 (N_5198,N_2594,N_3765);
or U5199 (N_5199,N_2575,N_4155);
and U5200 (N_5200,N_4315,N_3233);
and U5201 (N_5201,N_3510,N_3656);
nor U5202 (N_5202,N_2726,N_2890);
or U5203 (N_5203,N_3948,N_3059);
and U5204 (N_5204,N_2632,N_2852);
or U5205 (N_5205,N_2671,N_4443);
nor U5206 (N_5206,N_3227,N_3224);
nand U5207 (N_5207,N_2627,N_4051);
and U5208 (N_5208,N_4184,N_3640);
nor U5209 (N_5209,N_3442,N_4746);
nand U5210 (N_5210,N_3855,N_4833);
or U5211 (N_5211,N_2538,N_3705);
or U5212 (N_5212,N_2634,N_3887);
xnor U5213 (N_5213,N_2900,N_2517);
nor U5214 (N_5214,N_4403,N_3897);
and U5215 (N_5215,N_2938,N_3134);
or U5216 (N_5216,N_4092,N_3177);
nor U5217 (N_5217,N_3404,N_4521);
and U5218 (N_5218,N_4381,N_2743);
or U5219 (N_5219,N_2636,N_2922);
or U5220 (N_5220,N_4801,N_2591);
and U5221 (N_5221,N_3587,N_3428);
and U5222 (N_5222,N_3763,N_3170);
nor U5223 (N_5223,N_4346,N_2946);
or U5224 (N_5224,N_3553,N_3683);
nor U5225 (N_5225,N_4048,N_3469);
or U5226 (N_5226,N_3612,N_3391);
nor U5227 (N_5227,N_3686,N_2600);
xor U5228 (N_5228,N_3682,N_2762);
or U5229 (N_5229,N_3354,N_3798);
nor U5230 (N_5230,N_3806,N_2833);
nand U5231 (N_5231,N_4681,N_2868);
nor U5232 (N_5232,N_2557,N_4028);
and U5233 (N_5233,N_3096,N_3131);
nand U5234 (N_5234,N_3779,N_2595);
nor U5235 (N_5235,N_3979,N_3815);
nor U5236 (N_5236,N_2597,N_3202);
nor U5237 (N_5237,N_3700,N_3590);
nor U5238 (N_5238,N_3684,N_2967);
or U5239 (N_5239,N_3734,N_3728);
nand U5240 (N_5240,N_3052,N_3189);
or U5241 (N_5241,N_4949,N_3525);
and U5242 (N_5242,N_2834,N_4408);
nand U5243 (N_5243,N_2660,N_2926);
xor U5244 (N_5244,N_4137,N_3147);
nor U5245 (N_5245,N_3973,N_2715);
and U5246 (N_5246,N_3639,N_3537);
and U5247 (N_5247,N_3311,N_3962);
nor U5248 (N_5248,N_3811,N_4715);
and U5249 (N_5249,N_3085,N_4200);
or U5250 (N_5250,N_4617,N_3794);
nand U5251 (N_5251,N_4235,N_3485);
nand U5252 (N_5252,N_4881,N_4198);
and U5253 (N_5253,N_3457,N_3347);
nor U5254 (N_5254,N_3782,N_4192);
nor U5255 (N_5255,N_3733,N_3148);
or U5256 (N_5256,N_4695,N_3204);
nor U5257 (N_5257,N_3748,N_2690);
or U5258 (N_5258,N_4386,N_2661);
and U5259 (N_5259,N_2662,N_4082);
nor U5260 (N_5260,N_4063,N_3459);
and U5261 (N_5261,N_3799,N_4788);
and U5262 (N_5262,N_4808,N_3019);
or U5263 (N_5263,N_4893,N_2563);
or U5264 (N_5264,N_3994,N_4971);
nor U5265 (N_5265,N_4373,N_4406);
nor U5266 (N_5266,N_2934,N_2674);
and U5267 (N_5267,N_3967,N_4114);
nand U5268 (N_5268,N_4049,N_4420);
xnor U5269 (N_5269,N_3264,N_3918);
nor U5270 (N_5270,N_2969,N_2940);
nand U5271 (N_5271,N_3519,N_4820);
nand U5272 (N_5272,N_4735,N_3922);
and U5273 (N_5273,N_3033,N_2592);
and U5274 (N_5274,N_3509,N_2991);
nand U5275 (N_5275,N_4932,N_2703);
nand U5276 (N_5276,N_4475,N_2871);
and U5277 (N_5277,N_3495,N_2853);
nor U5278 (N_5278,N_3487,N_4143);
nand U5279 (N_5279,N_2570,N_4024);
nand U5280 (N_5280,N_4816,N_2870);
nand U5281 (N_5281,N_4786,N_2945);
nor U5282 (N_5282,N_2893,N_3749);
nand U5283 (N_5283,N_4889,N_4161);
nand U5284 (N_5284,N_3936,N_4614);
nand U5285 (N_5285,N_4676,N_2734);
nand U5286 (N_5286,N_3980,N_4569);
nor U5287 (N_5287,N_2565,N_2519);
or U5288 (N_5288,N_3556,N_3754);
xnor U5289 (N_5289,N_2700,N_4223);
and U5290 (N_5290,N_4604,N_2745);
nor U5291 (N_5291,N_4812,N_4647);
nor U5292 (N_5292,N_4167,N_3927);
and U5293 (N_5293,N_4599,N_3174);
and U5294 (N_5294,N_4740,N_3551);
or U5295 (N_5295,N_4439,N_4146);
nor U5296 (N_5296,N_4005,N_2666);
nor U5297 (N_5297,N_4663,N_2541);
and U5298 (N_5298,N_3524,N_4578);
or U5299 (N_5299,N_2792,N_4148);
and U5300 (N_5300,N_3416,N_3299);
and U5301 (N_5301,N_4864,N_3229);
and U5302 (N_5302,N_4258,N_3178);
nand U5303 (N_5303,N_2811,N_4298);
nor U5304 (N_5304,N_4880,N_2858);
and U5305 (N_5305,N_4969,N_2876);
nand U5306 (N_5306,N_4817,N_4417);
nand U5307 (N_5307,N_4712,N_4997);
nor U5308 (N_5308,N_3672,N_4135);
nor U5309 (N_5309,N_4755,N_3760);
and U5310 (N_5310,N_3714,N_4589);
nand U5311 (N_5311,N_4079,N_4437);
or U5312 (N_5312,N_2626,N_3172);
nor U5313 (N_5313,N_3923,N_3092);
or U5314 (N_5314,N_3471,N_4809);
or U5315 (N_5315,N_3272,N_4145);
and U5316 (N_5316,N_3357,N_3326);
nand U5317 (N_5317,N_4974,N_4180);
nor U5318 (N_5318,N_3360,N_4704);
and U5319 (N_5319,N_4535,N_4446);
nor U5320 (N_5320,N_3070,N_3004);
or U5321 (N_5321,N_4683,N_4153);
and U5322 (N_5322,N_4741,N_3370);
and U5323 (N_5323,N_3339,N_4018);
and U5324 (N_5324,N_2628,N_4526);
nand U5325 (N_5325,N_4432,N_2764);
nor U5326 (N_5326,N_2901,N_2656);
nor U5327 (N_5327,N_4926,N_3046);
and U5328 (N_5328,N_4301,N_3660);
nor U5329 (N_5329,N_3498,N_4123);
nand U5330 (N_5330,N_4558,N_3332);
or U5331 (N_5331,N_3318,N_2673);
or U5332 (N_5332,N_2652,N_2793);
nand U5333 (N_5333,N_2668,N_2659);
nor U5334 (N_5334,N_3678,N_4056);
or U5335 (N_5335,N_3242,N_4767);
and U5336 (N_5336,N_4543,N_2957);
nand U5337 (N_5337,N_3690,N_4990);
nor U5338 (N_5338,N_4270,N_4083);
or U5339 (N_5339,N_3692,N_4486);
nand U5340 (N_5340,N_2553,N_4942);
and U5341 (N_5341,N_4652,N_3659);
nand U5342 (N_5342,N_4985,N_4943);
nor U5343 (N_5343,N_2903,N_3872);
nor U5344 (N_5344,N_4382,N_4546);
and U5345 (N_5345,N_3858,N_4643);
nor U5346 (N_5346,N_3026,N_3969);
and U5347 (N_5347,N_3275,N_3220);
or U5348 (N_5348,N_3100,N_4325);
or U5349 (N_5349,N_3859,N_4623);
and U5350 (N_5350,N_4368,N_4284);
nor U5351 (N_5351,N_2988,N_4389);
or U5352 (N_5352,N_2738,N_2884);
nor U5353 (N_5353,N_3830,N_3574);
nand U5354 (N_5354,N_3436,N_4333);
nand U5355 (N_5355,N_2915,N_3711);
and U5356 (N_5356,N_2732,N_3300);
and U5357 (N_5357,N_3122,N_4700);
and U5358 (N_5358,N_4021,N_4292);
and U5359 (N_5359,N_3312,N_3323);
or U5360 (N_5360,N_2708,N_4772);
nand U5361 (N_5361,N_4899,N_3159);
and U5362 (N_5362,N_2782,N_2646);
or U5363 (N_5363,N_4228,N_2537);
nor U5364 (N_5364,N_3261,N_3450);
xor U5365 (N_5365,N_4042,N_2843);
nor U5366 (N_5366,N_4030,N_3933);
and U5367 (N_5367,N_3539,N_4445);
or U5368 (N_5368,N_3655,N_3065);
and U5369 (N_5369,N_3740,N_3028);
or U5370 (N_5370,N_4497,N_3076);
nor U5371 (N_5371,N_2589,N_3290);
or U5372 (N_5372,N_3968,N_4751);
nor U5373 (N_5373,N_4253,N_2906);
or U5374 (N_5374,N_3448,N_4196);
or U5375 (N_5375,N_4934,N_4510);
nor U5376 (N_5376,N_4399,N_3993);
and U5377 (N_5377,N_4655,N_3557);
and U5378 (N_5378,N_2504,N_3770);
nor U5379 (N_5379,N_3580,N_4793);
or U5380 (N_5380,N_3657,N_4954);
or U5381 (N_5381,N_2855,N_4134);
xor U5382 (N_5382,N_3094,N_4611);
nand U5383 (N_5383,N_2950,N_3032);
or U5384 (N_5384,N_3458,N_4117);
nor U5385 (N_5385,N_2705,N_2664);
nor U5386 (N_5386,N_4930,N_2694);
nor U5387 (N_5387,N_4416,N_3726);
nand U5388 (N_5388,N_4779,N_2524);
and U5389 (N_5389,N_3995,N_3392);
and U5390 (N_5390,N_3425,N_4871);
nor U5391 (N_5391,N_4867,N_3688);
nand U5392 (N_5392,N_3203,N_3205);
nor U5393 (N_5393,N_2506,N_4882);
and U5394 (N_5394,N_4859,N_4115);
nor U5395 (N_5395,N_4845,N_4088);
nor U5396 (N_5396,N_3044,N_3947);
nand U5397 (N_5397,N_3638,N_4693);
or U5398 (N_5398,N_3715,N_4442);
nand U5399 (N_5399,N_4043,N_3235);
or U5400 (N_5400,N_3024,N_3289);
xor U5401 (N_5401,N_3626,N_2549);
and U5402 (N_5402,N_2780,N_4861);
and U5403 (N_5403,N_4335,N_3099);
and U5404 (N_5404,N_3880,N_4199);
nor U5405 (N_5405,N_4720,N_3380);
and U5406 (N_5406,N_3365,N_4873);
nor U5407 (N_5407,N_4433,N_4878);
nand U5408 (N_5408,N_2930,N_3836);
and U5409 (N_5409,N_4255,N_4187);
and U5410 (N_5410,N_4905,N_4973);
nor U5411 (N_5411,N_3579,N_2838);
or U5412 (N_5412,N_2718,N_3125);
nor U5413 (N_5413,N_4448,N_3356);
nand U5414 (N_5414,N_2997,N_3086);
nor U5415 (N_5415,N_4364,N_3831);
nand U5416 (N_5416,N_2526,N_3153);
and U5417 (N_5417,N_4811,N_3862);
nor U5418 (N_5418,N_3848,N_4632);
nor U5419 (N_5419,N_4242,N_4694);
nand U5420 (N_5420,N_2550,N_3710);
and U5421 (N_5421,N_2631,N_4481);
and U5422 (N_5422,N_2802,N_3679);
or U5423 (N_5423,N_2995,N_3211);
nand U5424 (N_5424,N_3126,N_4565);
nand U5425 (N_5425,N_3265,N_3338);
nand U5426 (N_5426,N_4113,N_3691);
nand U5427 (N_5427,N_3588,N_2895);
nand U5428 (N_5428,N_3282,N_4834);
or U5429 (N_5429,N_2798,N_3821);
nor U5430 (N_5430,N_4947,N_4729);
or U5431 (N_5431,N_2808,N_3616);
nand U5432 (N_5432,N_3623,N_4363);
or U5433 (N_5433,N_4240,N_4994);
nand U5434 (N_5434,N_4336,N_3406);
nand U5435 (N_5435,N_3905,N_4554);
or U5436 (N_5436,N_3865,N_2894);
nand U5437 (N_5437,N_4392,N_4619);
or U5438 (N_5438,N_3572,N_2902);
and U5439 (N_5439,N_4870,N_2779);
or U5440 (N_5440,N_3658,N_3934);
nand U5441 (N_5441,N_3468,N_4984);
and U5442 (N_5442,N_4170,N_3173);
and U5443 (N_5443,N_4109,N_2753);
nand U5444 (N_5444,N_2582,N_3617);
and U5445 (N_5445,N_2577,N_3976);
or U5446 (N_5446,N_3735,N_4641);
and U5447 (N_5447,N_2849,N_4239);
or U5448 (N_5448,N_2566,N_3284);
nand U5449 (N_5449,N_4306,N_2928);
or U5450 (N_5450,N_4009,N_3155);
or U5451 (N_5451,N_3846,N_3376);
and U5452 (N_5452,N_3057,N_2889);
nor U5453 (N_5453,N_4545,N_4679);
nor U5454 (N_5454,N_3803,N_4993);
or U5455 (N_5455,N_3090,N_3805);
and U5456 (N_5456,N_3942,N_2845);
and U5457 (N_5457,N_4799,N_2805);
nand U5458 (N_5458,N_4327,N_3628);
nor U5459 (N_5459,N_4274,N_2605);
and U5460 (N_5460,N_3843,N_3645);
nor U5461 (N_5461,N_2588,N_2618);
and U5462 (N_5462,N_3861,N_4868);
nand U5463 (N_5463,N_4860,N_2769);
or U5464 (N_5464,N_3610,N_3827);
and U5465 (N_5465,N_4150,N_3744);
or U5466 (N_5466,N_2841,N_4457);
and U5467 (N_5467,N_4975,N_4296);
and U5468 (N_5468,N_4365,N_3330);
nor U5469 (N_5469,N_4653,N_4897);
nor U5470 (N_5470,N_3719,N_3003);
nor U5471 (N_5471,N_4283,N_3957);
and U5472 (N_5472,N_3012,N_2507);
or U5473 (N_5473,N_4675,N_3340);
and U5474 (N_5474,N_3483,N_4794);
and U5475 (N_5475,N_4541,N_3010);
or U5476 (N_5476,N_3216,N_3000);
nor U5477 (N_5477,N_4033,N_3115);
and U5478 (N_5478,N_4195,N_2622);
nand U5479 (N_5479,N_3081,N_4854);
nand U5480 (N_5480,N_4719,N_4586);
nand U5481 (N_5481,N_2815,N_3164);
nand U5482 (N_5482,N_4393,N_4372);
nand U5483 (N_5483,N_3755,N_2515);
and U5484 (N_5484,N_3687,N_4276);
or U5485 (N_5485,N_3970,N_4011);
or U5486 (N_5486,N_4003,N_4661);
and U5487 (N_5487,N_3054,N_2684);
or U5488 (N_5488,N_2948,N_2741);
nand U5489 (N_5489,N_4178,N_4395);
nand U5490 (N_5490,N_3165,N_3050);
nor U5491 (N_5491,N_3698,N_3219);
nor U5492 (N_5492,N_3267,N_4810);
nand U5493 (N_5493,N_3802,N_4026);
or U5494 (N_5494,N_4991,N_3381);
or U5495 (N_5495,N_3899,N_4072);
and U5496 (N_5496,N_3464,N_2989);
or U5497 (N_5497,N_3088,N_4173);
nor U5498 (N_5498,N_2624,N_3851);
nand U5499 (N_5499,N_4424,N_2545);
or U5500 (N_5500,N_3364,N_4244);
or U5501 (N_5501,N_3274,N_3486);
nor U5502 (N_5502,N_3825,N_4995);
nor U5503 (N_5503,N_4670,N_2990);
and U5504 (N_5504,N_3730,N_2647);
nor U5505 (N_5505,N_4851,N_4193);
and U5506 (N_5506,N_4725,N_3022);
nor U5507 (N_5507,N_3797,N_3915);
nor U5508 (N_5508,N_2904,N_4227);
and U5509 (N_5509,N_2568,N_3966);
and U5510 (N_5510,N_2911,N_4232);
nor U5511 (N_5511,N_4584,N_2837);
nand U5512 (N_5512,N_4523,N_4421);
or U5513 (N_5513,N_3785,N_4831);
nand U5514 (N_5514,N_3327,N_4548);
and U5515 (N_5515,N_3255,N_4300);
or U5516 (N_5516,N_2540,N_2614);
nand U5517 (N_5517,N_4999,N_4686);
nor U5518 (N_5518,N_2697,N_4488);
nand U5519 (N_5519,N_4371,N_3573);
nor U5520 (N_5520,N_3527,N_3542);
nor U5521 (N_5521,N_2862,N_4929);
nand U5522 (N_5522,N_3055,N_3577);
nor U5523 (N_5523,N_2739,N_2784);
and U5524 (N_5524,N_3453,N_3591);
and U5525 (N_5525,N_3475,N_2516);
and U5526 (N_5526,N_2623,N_2774);
nor U5527 (N_5527,N_4847,N_4597);
or U5528 (N_5528,N_3438,N_4650);
and U5529 (N_5529,N_4212,N_2711);
nand U5530 (N_5530,N_4343,N_4582);
nor U5531 (N_5531,N_4731,N_2885);
or U5532 (N_5532,N_4838,N_2796);
xor U5533 (N_5533,N_2500,N_3538);
nand U5534 (N_5534,N_4646,N_4059);
or U5535 (N_5535,N_4960,N_2982);
and U5536 (N_5536,N_4476,N_4722);
nor U5537 (N_5537,N_3839,N_4027);
or U5538 (N_5538,N_4322,N_4561);
or U5539 (N_5539,N_4826,N_2523);
and U5540 (N_5540,N_4534,N_2830);
and U5541 (N_5541,N_4921,N_4111);
nand U5542 (N_5542,N_4405,N_3649);
nor U5543 (N_5543,N_4827,N_2812);
and U5544 (N_5544,N_4503,N_3348);
nand U5545 (N_5545,N_3410,N_4588);
or U5546 (N_5546,N_4289,N_2879);
nor U5547 (N_5547,N_2863,N_3913);
nor U5548 (N_5548,N_2960,N_3098);
or U5549 (N_5549,N_3795,N_4983);
or U5550 (N_5550,N_3889,N_3293);
and U5551 (N_5551,N_3136,N_2939);
and U5552 (N_5552,N_2867,N_2579);
nor U5553 (N_5553,N_2720,N_2850);
and U5554 (N_5554,N_4964,N_4094);
nand U5555 (N_5555,N_4877,N_4098);
nand U5556 (N_5556,N_3358,N_4414);
xnor U5557 (N_5557,N_3384,N_2648);
or U5558 (N_5558,N_3676,N_3725);
nor U5559 (N_5559,N_3570,N_3737);
nor U5560 (N_5560,N_4016,N_2755);
nand U5561 (N_5561,N_3301,N_3181);
and U5562 (N_5562,N_3071,N_3222);
and U5563 (N_5563,N_4271,N_2996);
and U5564 (N_5564,N_4978,N_3061);
nor U5565 (N_5565,N_4461,N_4224);
and U5566 (N_5566,N_2816,N_4514);
nand U5567 (N_5567,N_3402,N_4642);
and U5568 (N_5568,N_2775,N_3040);
nand U5569 (N_5569,N_3001,N_3195);
or U5570 (N_5570,N_4286,N_4191);
nand U5571 (N_5571,N_4402,N_2810);
or U5572 (N_5572,N_3184,N_3190);
nor U5573 (N_5573,N_2730,N_4344);
and U5574 (N_5574,N_4885,N_4099);
or U5575 (N_5575,N_2797,N_4844);
nand U5576 (N_5576,N_4347,N_4321);
or U5577 (N_5577,N_4015,N_4456);
nor U5578 (N_5578,N_2809,N_2543);
and U5579 (N_5579,N_2935,N_4440);
and U5580 (N_5580,N_4903,N_3210);
and U5581 (N_5581,N_4776,N_3281);
nand U5582 (N_5582,N_4260,N_3920);
nor U5583 (N_5583,N_3480,N_3764);
nand U5584 (N_5584,N_4360,N_2503);
or U5585 (N_5585,N_4501,N_4628);
nand U5586 (N_5586,N_4341,N_4064);
nand U5587 (N_5587,N_3435,N_2869);
and U5588 (N_5588,N_2829,N_2710);
or U5589 (N_5589,N_3632,N_2522);
or U5590 (N_5590,N_3513,N_3981);
nor U5591 (N_5591,N_3613,N_4631);
nand U5592 (N_5592,N_3978,N_4458);
nand U5593 (N_5593,N_2962,N_2689);
nand U5594 (N_5594,N_3334,N_4366);
nor U5595 (N_5595,N_3008,N_2827);
nand U5596 (N_5596,N_2564,N_3742);
or U5597 (N_5597,N_3838,N_4288);
nand U5598 (N_5598,N_2851,N_3585);
nor U5599 (N_5599,N_3829,N_3320);
and U5600 (N_5600,N_3622,N_3236);
and U5601 (N_5601,N_2994,N_2947);
nor U5602 (N_5602,N_2583,N_3708);
or U5603 (N_5603,N_4369,N_4485);
nand U5604 (N_5604,N_3756,N_4924);
nand U5605 (N_5605,N_3186,N_3833);
nor U5606 (N_5606,N_3390,N_3361);
nand U5607 (N_5607,N_4129,N_3427);
nand U5608 (N_5608,N_2707,N_4866);
or U5609 (N_5609,N_2773,N_4107);
or U5610 (N_5610,N_3786,N_2641);
and U5611 (N_5611,N_2559,N_3045);
nand U5612 (N_5612,N_2831,N_4000);
nor U5613 (N_5613,N_3609,N_3296);
and U5614 (N_5614,N_3759,N_3804);
and U5615 (N_5615,N_3555,N_4699);
nand U5616 (N_5616,N_4058,N_3212);
nor U5617 (N_5617,N_2733,N_4892);
nor U5618 (N_5618,N_4320,N_2777);
nand U5619 (N_5619,N_3636,N_3596);
nand U5620 (N_5620,N_4062,N_3403);
and U5621 (N_5621,N_3757,N_3697);
or U5622 (N_5622,N_2978,N_3401);
or U5623 (N_5623,N_3784,N_4061);
nand U5624 (N_5624,N_3881,N_3349);
and U5625 (N_5625,N_2505,N_3150);
nor U5626 (N_5626,N_2790,N_2677);
nand U5627 (N_5627,N_3878,N_4918);
nand U5628 (N_5628,N_4912,N_4037);
or U5629 (N_5629,N_3303,N_2786);
nand U5630 (N_5630,N_3800,N_4506);
or U5631 (N_5631,N_4265,N_4281);
nor U5632 (N_5632,N_3066,N_3951);
nor U5633 (N_5633,N_4268,N_4805);
or U5634 (N_5634,N_4630,N_3058);
nor U5635 (N_5635,N_3953,N_3752);
or U5636 (N_5636,N_4186,N_3589);
and U5637 (N_5637,N_2828,N_3393);
nand U5638 (N_5638,N_4036,N_3548);
nand U5639 (N_5639,N_3615,N_3221);
nor U5640 (N_5640,N_4144,N_3129);
or U5641 (N_5641,N_4691,N_4029);
and U5642 (N_5642,N_4001,N_4895);
nand U5643 (N_5643,N_3955,N_3292);
or U5644 (N_5644,N_3194,N_2971);
or U5645 (N_5645,N_3232,N_3305);
nand U5646 (N_5646,N_3262,N_2680);
nor U5647 (N_5647,N_4680,N_4342);
nand U5648 (N_5648,N_3907,N_3879);
and U5649 (N_5649,N_3892,N_3411);
or U5650 (N_5650,N_2937,N_4089);
nand U5651 (N_5651,N_2958,N_3845);
nand U5652 (N_5652,N_3285,N_4494);
nor U5653 (N_5653,N_4210,N_3738);
and U5654 (N_5654,N_4291,N_3398);
and U5655 (N_5655,N_4249,N_4901);
nor U5656 (N_5656,N_4566,N_3528);
nor U5657 (N_5657,N_3231,N_2682);
and U5658 (N_5658,N_4797,N_3566);
and U5659 (N_5659,N_4869,N_4574);
nand U5660 (N_5660,N_3095,N_3250);
nand U5661 (N_5661,N_3089,N_3109);
or U5662 (N_5662,N_4713,N_3917);
nor U5663 (N_5663,N_3564,N_4762);
nor U5664 (N_5664,N_3768,N_4637);
or U5665 (N_5665,N_3474,N_4168);
or U5666 (N_5666,N_3650,N_2791);
and U5667 (N_5667,N_3452,N_4925);
and U5668 (N_5668,N_2751,N_4297);
nand U5669 (N_5669,N_3350,N_3158);
nor U5670 (N_5670,N_3944,N_2910);
or U5671 (N_5671,N_2691,N_3565);
nor U5672 (N_5672,N_2644,N_4972);
or U5673 (N_5673,N_2548,N_2857);
nor U5674 (N_5674,N_3317,N_4705);
nor U5675 (N_5675,N_3844,N_2824);
nor U5676 (N_5676,N_4362,N_3408);
or U5677 (N_5677,N_3877,N_4206);
nor U5678 (N_5678,N_2737,N_3082);
or U5679 (N_5679,N_4359,N_4263);
nor U5680 (N_5680,N_3521,N_4610);
or U5681 (N_5681,N_3996,N_2531);
or U5682 (N_5682,N_4828,N_3531);
and U5683 (N_5683,N_4622,N_3108);
or U5684 (N_5684,N_3257,N_2799);
nor U5685 (N_5685,N_3341,N_4843);
nand U5686 (N_5686,N_4070,N_4053);
nand U5687 (N_5687,N_2688,N_3958);
nand U5688 (N_5688,N_4002,N_2759);
nor U5689 (N_5689,N_3972,N_3062);
and U5690 (N_5690,N_4919,N_3051);
nor U5691 (N_5691,N_4787,N_4916);
and U5692 (N_5692,N_3479,N_3732);
nor U5693 (N_5693,N_2696,N_2813);
or U5694 (N_5694,N_4938,N_4516);
xnor U5695 (N_5695,N_4319,N_4638);
nor U5696 (N_5696,N_3175,N_4697);
nand U5697 (N_5697,N_4324,N_2558);
nor U5698 (N_5698,N_3383,N_2965);
or U5699 (N_5699,N_4138,N_4738);
nand U5700 (N_5700,N_2953,N_4640);
nor U5701 (N_5701,N_4176,N_3651);
xor U5702 (N_5702,N_3582,N_3397);
nand U5703 (N_5703,N_2576,N_3260);
or U5704 (N_5704,N_3849,N_3005);
nor U5705 (N_5705,N_4649,N_4688);
or U5706 (N_5706,N_4330,N_3133);
nor U5707 (N_5707,N_4441,N_2998);
nor U5708 (N_5708,N_3721,N_4447);
and U5709 (N_5709,N_3675,N_3294);
or U5710 (N_5710,N_4658,N_3419);
nand U5711 (N_5711,N_2807,N_4590);
xnor U5712 (N_5712,N_4247,N_4207);
or U5713 (N_5713,N_3288,N_4807);
nand U5714 (N_5714,N_3328,N_3654);
nor U5715 (N_5715,N_3226,N_4950);
nand U5716 (N_5716,N_3298,N_2633);
nor U5717 (N_5717,N_4032,N_4796);
nand U5718 (N_5718,N_4568,N_3241);
or U5719 (N_5719,N_3633,N_4898);
or U5720 (N_5720,N_4777,N_3670);
nand U5721 (N_5721,N_3502,N_4383);
and U5722 (N_5722,N_3578,N_3207);
or U5723 (N_5723,N_4656,N_2554);
and U5724 (N_5724,N_3956,N_3586);
and U5725 (N_5725,N_4222,N_4634);
or U5726 (N_5726,N_3395,N_4310);
or U5727 (N_5727,N_4226,N_3891);
or U5728 (N_5728,N_3619,N_2788);
or U5729 (N_5729,N_3547,N_4380);
and U5730 (N_5730,N_2785,N_2848);
or U5731 (N_5731,N_3777,N_2552);
nand U5732 (N_5732,N_4958,N_4418);
nor U5733 (N_5733,N_3520,N_2898);
and U5734 (N_5734,N_2685,N_4813);
and U5735 (N_5735,N_2854,N_3171);
nor U5736 (N_5736,N_4760,N_4166);
or U5737 (N_5737,N_4909,N_2747);
nand U5738 (N_5738,N_2896,N_2949);
nor U5739 (N_5739,N_4479,N_4967);
or U5740 (N_5740,N_4175,N_2619);
or U5741 (N_5741,N_4884,N_4355);
nand U5742 (N_5742,N_3497,N_4908);
or U5743 (N_5743,N_4105,N_3791);
nor U5744 (N_5744,N_3490,N_2908);
and U5745 (N_5745,N_3960,N_4177);
nor U5746 (N_5746,N_4651,N_2748);
and U5747 (N_5747,N_4278,N_2723);
or U5748 (N_5748,N_3518,N_3850);
or U5749 (N_5749,N_4495,N_4515);
nor U5750 (N_5750,N_3335,N_4931);
and U5751 (N_5751,N_3837,N_3346);
nor U5752 (N_5752,N_4540,N_3372);
nor U5753 (N_5753,N_4483,N_4963);
nor U5754 (N_5754,N_4132,N_3671);
xor U5755 (N_5755,N_4553,N_4378);
nand U5756 (N_5756,N_2866,N_3523);
nand U5757 (N_5757,N_3169,N_4449);
nor U5758 (N_5758,N_4520,N_3745);
and U5759 (N_5759,N_3378,N_4174);
or U5760 (N_5760,N_4626,N_3371);
nand U5761 (N_5761,N_3034,N_3543);
nor U5762 (N_5762,N_3077,N_2731);
nand U5763 (N_5763,N_4621,N_4814);
or U5764 (N_5764,N_4012,N_3128);
nor U5765 (N_5765,N_3417,N_4472);
nand U5766 (N_5766,N_3023,N_3567);
nand U5767 (N_5767,N_3766,N_3141);
or U5768 (N_5768,N_4358,N_2546);
nor U5769 (N_5769,N_4370,N_4213);
and U5770 (N_5770,N_4726,N_4771);
and U5771 (N_5771,N_4667,N_3473);
and U5772 (N_5772,N_2803,N_4084);
and U5773 (N_5773,N_3325,N_3053);
nand U5774 (N_5774,N_3467,N_4835);
and U5775 (N_5775,N_3723,N_3634);
or U5776 (N_5776,N_2860,N_4575);
and U5777 (N_5777,N_4470,N_3824);
and U5778 (N_5778,N_4579,N_3286);
or U5779 (N_5779,N_3677,N_4431);
or U5780 (N_5780,N_4573,N_3741);
or U5781 (N_5781,N_3614,N_4549);
and U5782 (N_5782,N_3106,N_4778);
or U5783 (N_5783,N_4692,N_3822);
and U5784 (N_5784,N_4703,N_4505);
and U5785 (N_5785,N_4955,N_3223);
nand U5786 (N_5786,N_2913,N_4733);
or U5787 (N_5787,N_4872,N_4100);
nand U5788 (N_5788,N_3117,N_4385);
or U5789 (N_5789,N_3443,N_2609);
nand U5790 (N_5790,N_3295,N_4349);
and U5791 (N_5791,N_4830,N_3176);
nand U5792 (N_5792,N_4769,N_4182);
nor U5793 (N_5793,N_3926,N_2970);
nand U5794 (N_5794,N_4736,N_4396);
or U5795 (N_5795,N_2887,N_2533);
nand U5796 (N_5796,N_4077,N_4987);
nand U5797 (N_5797,N_4798,N_2966);
nor U5798 (N_5798,N_3049,N_4992);
nand U5799 (N_5799,N_4118,N_3042);
nor U5800 (N_5800,N_3208,N_3569);
and U5801 (N_5801,N_3353,N_3545);
nor U5802 (N_5802,N_4928,N_3355);
nor U5803 (N_5803,N_3999,N_2819);
nor U5804 (N_5804,N_4780,N_3793);
or U5805 (N_5805,N_3217,N_2999);
or U5806 (N_5806,N_3924,N_3121);
nor U5807 (N_5807,N_3828,N_4165);
and U5808 (N_5808,N_4257,N_2778);
or U5809 (N_5809,N_2729,N_3237);
and U5810 (N_5810,N_3868,N_4784);
and U5811 (N_5811,N_3621,N_4552);
xor U5812 (N_5812,N_3254,N_2916);
and U5813 (N_5813,N_3603,N_3643);
nor U5814 (N_5814,N_3343,N_3549);
or U5815 (N_5815,N_3694,N_4876);
nor U5816 (N_5816,N_3988,N_3198);
or U5817 (N_5817,N_4585,N_3466);
and U5818 (N_5818,N_2602,N_4875);
or U5819 (N_5819,N_3743,N_3641);
or U5820 (N_5820,N_2801,N_3014);
nand U5821 (N_5821,N_4750,N_4492);
or U5822 (N_5822,N_3439,N_3256);
nor U5823 (N_5823,N_4197,N_4853);
xor U5824 (N_5824,N_3624,N_3400);
nand U5825 (N_5825,N_4214,N_3890);
or U5826 (N_5826,N_3941,N_4665);
nand U5827 (N_5827,N_4961,N_4090);
xnor U5828 (N_5828,N_4423,N_4753);
or U5829 (N_5829,N_3900,N_4839);
and U5830 (N_5830,N_3693,N_3319);
nor U5831 (N_5831,N_4900,N_2544);
or U5832 (N_5832,N_4266,N_4435);
nor U5833 (N_5833,N_4246,N_2593);
nor U5834 (N_5834,N_4902,N_3673);
or U5835 (N_5835,N_3605,N_3036);
and U5836 (N_5836,N_2864,N_4217);
nor U5837 (N_5837,N_3461,N_2973);
or U5838 (N_5838,N_3447,N_2758);
nor U5839 (N_5839,N_3883,N_3101);
and U5840 (N_5840,N_4718,N_2754);
nand U5841 (N_5841,N_3593,N_4172);
nand U5842 (N_5842,N_3251,N_3333);
nor U5843 (N_5843,N_4219,N_4022);
and U5844 (N_5844,N_2712,N_4351);
xor U5845 (N_5845,N_2832,N_4537);
and U5846 (N_5846,N_4752,N_3826);
or U5847 (N_5847,N_3950,N_3680);
nand U5848 (N_5848,N_4124,N_2509);
nor U5849 (N_5849,N_3430,N_3873);
and U5850 (N_5850,N_3963,N_3514);
nand U5851 (N_5851,N_3482,N_4428);
nor U5852 (N_5852,N_2596,N_4915);
or U5853 (N_5853,N_3455,N_4444);
nand U5854 (N_5854,N_4211,N_3481);
nor U5855 (N_5855,N_3716,N_4774);
and U5856 (N_5856,N_2676,N_2968);
or U5857 (N_5857,N_4426,N_3501);
and U5858 (N_5858,N_4047,N_4102);
or U5859 (N_5859,N_3366,N_4714);
nor U5860 (N_5860,N_3268,N_3456);
and U5861 (N_5861,N_4616,N_4427);
nor U5862 (N_5862,N_4491,N_3413);
nand U5863 (N_5863,N_4945,N_2536);
nor U5864 (N_5864,N_4544,N_3929);
nor U5865 (N_5865,N_4499,N_4890);
and U5866 (N_5866,N_2924,N_3662);
nor U5867 (N_5867,N_4040,N_4837);
and U5868 (N_5868,N_3363,N_2620);
nor U5869 (N_5869,N_2693,N_4231);
and U5870 (N_5870,N_4136,N_4672);
nand U5871 (N_5871,N_2914,N_2952);
nand U5872 (N_5872,N_3314,N_3949);
or U5873 (N_5873,N_4407,N_2527);
or U5874 (N_5874,N_4374,N_4086);
nor U5875 (N_5875,N_4758,N_4933);
nor U5876 (N_5876,N_4025,N_4387);
and U5877 (N_5877,N_4237,N_4465);
nand U5878 (N_5878,N_3753,N_3068);
and U5879 (N_5879,N_3817,N_4285);
nand U5880 (N_5880,N_2749,N_4334);
nor U5881 (N_5881,N_2861,N_3526);
or U5882 (N_5882,N_3007,N_2992);
or U5883 (N_5883,N_3421,N_4467);
or U5884 (N_5884,N_4957,N_3608);
or U5885 (N_5885,N_2771,N_3377);
or U5886 (N_5886,N_3712,N_4112);
nor U5887 (N_5887,N_4572,N_4295);
and U5888 (N_5888,N_3379,N_3484);
nand U5889 (N_5889,N_3138,N_3635);
nor U5890 (N_5890,N_4238,N_4724);
nand U5891 (N_5891,N_3113,N_3104);
or U5892 (N_5892,N_4013,N_4085);
nand U5893 (N_5893,N_3352,N_2980);
or U5894 (N_5894,N_4233,N_2679);
nand U5895 (N_5895,N_4419,N_3078);
nor U5896 (N_5896,N_4041,N_4205);
nand U5897 (N_5897,N_2923,N_4450);
nand U5898 (N_5898,N_3642,N_2927);
and U5899 (N_5899,N_4010,N_3258);
nor U5900 (N_5900,N_3345,N_4203);
nor U5901 (N_5901,N_2665,N_2844);
nand U5902 (N_5902,N_3310,N_3336);
or U5903 (N_5903,N_3866,N_4530);
nor U5904 (N_5904,N_4716,N_2951);
nor U5905 (N_5905,N_4356,N_3731);
and U5906 (N_5906,N_3368,N_4204);
nand U5907 (N_5907,N_2918,N_2532);
and U5908 (N_5908,N_2744,N_4842);
nor U5909 (N_5909,N_2621,N_3269);
nor U5910 (N_5910,N_4685,N_3931);
and U5911 (N_5911,N_3249,N_3449);
or U5912 (N_5912,N_3707,N_3064);
nor U5913 (N_5913,N_2920,N_4299);
nand U5914 (N_5914,N_4050,N_2859);
xnor U5915 (N_5915,N_4474,N_2584);
and U5916 (N_5916,N_3476,N_4547);
nor U5917 (N_5917,N_2883,N_2919);
or U5918 (N_5918,N_4946,N_2956);
nor U5919 (N_5919,N_4057,N_4956);
nand U5920 (N_5920,N_4038,N_2907);
or U5921 (N_5921,N_4858,N_2678);
nand U5922 (N_5922,N_4581,N_3818);
nor U5923 (N_5923,N_3151,N_4133);
or U5924 (N_5924,N_3225,N_4259);
nand U5925 (N_5925,N_4338,N_4531);
and U5926 (N_5926,N_4763,N_4857);
and U5927 (N_5927,N_2976,N_4404);
nor U5928 (N_5928,N_4825,N_2756);
and U5929 (N_5929,N_4119,N_4158);
or U5930 (N_5930,N_3446,N_2562);
or U5931 (N_5931,N_3932,N_4261);
and U5932 (N_5932,N_3011,N_3781);
or U5933 (N_5933,N_2521,N_3568);
or U5934 (N_5934,N_3595,N_3415);
and U5935 (N_5935,N_2603,N_3792);
nand U5936 (N_5936,N_2804,N_4513);
or U5937 (N_5937,N_4759,N_3463);
and U5938 (N_5938,N_3367,N_3278);
or U5939 (N_5939,N_3017,N_3874);
xnor U5940 (N_5940,N_2654,N_3154);
nor U5941 (N_5941,N_3496,N_2587);
nand U5942 (N_5942,N_4629,N_3598);
nor U5943 (N_5943,N_4674,N_2818);
and U5944 (N_5944,N_3773,N_4055);
nand U5945 (N_5945,N_4654,N_4509);
or U5946 (N_5946,N_3653,N_3898);
and U5947 (N_5947,N_3304,N_2814);
or U5948 (N_5948,N_4862,N_4154);
or U5949 (N_5949,N_3067,N_2683);
nor U5950 (N_5950,N_4739,N_2975);
and U5951 (N_5951,N_2513,N_3991);
nor U5952 (N_5952,N_4709,N_3020);
nand U5953 (N_5953,N_3424,N_4594);
and U5954 (N_5954,N_4398,N_3489);
nand U5955 (N_5955,N_2847,N_3179);
nor U5956 (N_5956,N_2512,N_2892);
nand U5957 (N_5957,N_4906,N_4097);
and U5958 (N_5958,N_3102,N_4982);
nor U5959 (N_5959,N_4948,N_4608);
or U5960 (N_5960,N_2959,N_2717);
nor U5961 (N_5961,N_2763,N_4413);
or U5962 (N_5962,N_2658,N_4303);
nor U5963 (N_5963,N_2806,N_3188);
nand U5964 (N_5964,N_3937,N_3508);
or U5965 (N_5965,N_2713,N_4460);
nand U5966 (N_5966,N_4615,N_4734);
nor U5967 (N_5967,N_4567,N_4230);
nor U5968 (N_5968,N_2692,N_3093);
nand U5969 (N_5969,N_3097,N_4923);
nand U5970 (N_5970,N_3465,N_3432);
xnor U5971 (N_5971,N_3437,N_4331);
nand U5972 (N_5972,N_4313,N_3767);
or U5973 (N_5973,N_2825,N_4836);
or U5974 (N_5974,N_3916,N_2955);
nor U5975 (N_5975,N_2610,N_4689);
or U5976 (N_5976,N_3248,N_4014);
nor U5977 (N_5977,N_2567,N_2501);
or U5978 (N_5978,N_3192,N_3783);
nor U5979 (N_5979,N_2560,N_2638);
nor U5980 (N_5980,N_3493,N_2856);
and U5981 (N_5981,N_4290,N_2882);
or U5982 (N_5982,N_4252,N_4044);
nor U5983 (N_5983,N_4894,N_3060);
nor U5984 (N_5984,N_2599,N_3144);
and U5985 (N_5985,N_2581,N_3454);
or U5986 (N_5986,N_2645,N_4241);
nand U5987 (N_5987,N_4157,N_4463);
nand U5988 (N_5988,N_4659,N_4896);
nor U5989 (N_5989,N_2961,N_4512);
and U5990 (N_5990,N_4312,N_3611);
xor U5991 (N_5991,N_4275,N_3329);
nand U5992 (N_5992,N_4940,N_3247);
and U5993 (N_5993,N_4511,N_3856);
nor U5994 (N_5994,N_3559,N_3902);
nand U5995 (N_5995,N_2942,N_3056);
nand U5996 (N_5996,N_2649,N_3283);
nand U5997 (N_5997,N_4727,N_4078);
or U5998 (N_5998,N_4986,N_2607);
and U5999 (N_5999,N_4430,N_3041);
nor U6000 (N_6000,N_4367,N_3110);
nor U6001 (N_6001,N_3277,N_3013);
nor U6002 (N_6002,N_2740,N_3084);
or U6003 (N_6003,N_4944,N_3771);
or U6004 (N_6004,N_3901,N_2767);
nand U6005 (N_6005,N_4269,N_2629);
nand U6006 (N_6006,N_3253,N_3359);
nand U6007 (N_6007,N_4354,N_3674);
or U6008 (N_6008,N_3315,N_4603);
nor U6009 (N_6009,N_3914,N_4130);
nand U6010 (N_6010,N_4139,N_2601);
or U6011 (N_6011,N_2573,N_4104);
or U6012 (N_6012,N_4917,N_4865);
or U6013 (N_6013,N_4690,N_4846);
nand U6014 (N_6014,N_3103,N_3030);
nor U6015 (N_6015,N_3535,N_2820);
or U6016 (N_6016,N_3187,N_2612);
nand U6017 (N_6017,N_4821,N_3197);
or U6018 (N_6018,N_4879,N_4066);
xnor U6019 (N_6019,N_3909,N_4151);
xor U6020 (N_6020,N_4459,N_3245);
nand U6021 (N_6021,N_4060,N_3717);
nand U6022 (N_6022,N_4682,N_2822);
nor U6023 (N_6023,N_4765,N_4409);
or U6024 (N_6024,N_3532,N_4229);
or U6025 (N_6025,N_4287,N_3422);
nor U6026 (N_6026,N_2615,N_4438);
or U6027 (N_6027,N_4500,N_3373);
nand U6028 (N_6028,N_3515,N_4953);
nor U6029 (N_6029,N_3522,N_3083);
nand U6030 (N_6030,N_4517,N_4480);
nand U6031 (N_6031,N_2556,N_4490);
nor U6032 (N_6032,N_2640,N_3445);
nor U6033 (N_6033,N_3441,N_2635);
and U6034 (N_6034,N_3385,N_4818);
and U6035 (N_6035,N_3581,N_3160);
nor U6036 (N_6036,N_3644,N_4852);
and U6037 (N_6037,N_4749,N_3835);
nand U6038 (N_6038,N_3747,N_4981);
or U6039 (N_6039,N_4415,N_4464);
or U6040 (N_6040,N_4462,N_3954);
or U6041 (N_6041,N_3601,N_3910);
or U6042 (N_6042,N_4601,N_3885);
and U6043 (N_6043,N_2529,N_3685);
nor U6044 (N_6044,N_2520,N_2525);
nor U6045 (N_6045,N_3604,N_4071);
xor U6046 (N_6046,N_3713,N_2547);
or U6047 (N_6047,N_3037,N_4976);
or U6048 (N_6048,N_4907,N_3386);
nor U6049 (N_6049,N_3214,N_3575);
nor U6050 (N_6050,N_4743,N_2750);
nor U6051 (N_6051,N_3069,N_3387);
or U6052 (N_6052,N_4316,N_3998);
nand U6053 (N_6053,N_4225,N_3919);
and U6054 (N_6054,N_4980,N_2555);
nor U6055 (N_6055,N_4728,N_4108);
and U6056 (N_6056,N_3841,N_4737);
nand U6057 (N_6057,N_3243,N_3342);
nor U6058 (N_6058,N_3599,N_4201);
and U6059 (N_6059,N_4054,N_3666);
or U6060 (N_6060,N_2669,N_2826);
or U6061 (N_6061,N_4795,N_4309);
or U6062 (N_6062,N_4927,N_3886);
and U6063 (N_6063,N_3888,N_2657);
and U6064 (N_6064,N_4394,N_3706);
nor U6065 (N_6065,N_2878,N_4863);
nor U6066 (N_6066,N_2727,N_2630);
nor U6067 (N_6067,N_4273,N_4563);
or U6068 (N_6068,N_3213,N_2580);
and U6069 (N_6069,N_2616,N_3143);
and U6070 (N_6070,N_4073,N_4340);
or U6071 (N_6071,N_2984,N_4625);
nor U6072 (N_6072,N_4570,N_3989);
or U6073 (N_6073,N_3477,N_4529);
or U6074 (N_6074,N_4966,N_4156);
and U6075 (N_6075,N_2651,N_2944);
or U6076 (N_6076,N_4498,N_2761);
nor U6077 (N_6077,N_3306,N_4698);
nor U6078 (N_6078,N_4493,N_4307);
and U6079 (N_6079,N_4410,N_2728);
nand U6080 (N_6080,N_3727,N_3114);
or U6081 (N_6081,N_3389,N_3959);
and U6082 (N_6082,N_3939,N_3908);
nor U6083 (N_6083,N_4502,N_3307);
and U6084 (N_6084,N_3492,N_4243);
or U6085 (N_6085,N_4560,N_2569);
nor U6086 (N_6086,N_4730,N_4076);
or U6087 (N_6087,N_3111,N_2964);
nor U6088 (N_6088,N_3087,N_3156);
nand U6089 (N_6089,N_4536,N_3182);
and U6090 (N_6090,N_2535,N_4507);
and U6091 (N_6091,N_3751,N_4998);
nor U6092 (N_6092,N_4163,N_2724);
and U6093 (N_6093,N_4883,N_4189);
or U6094 (N_6094,N_3801,N_2880);
nand U6095 (N_6095,N_4802,N_4696);
xor U6096 (N_6096,N_4353,N_3440);
or U6097 (N_6097,N_3546,N_4636);
nor U6098 (N_6098,N_4121,N_3162);
or U6099 (N_6099,N_4748,N_2836);
nor U6100 (N_6100,N_4302,N_3536);
and U6101 (N_6101,N_4891,N_2768);
or U6102 (N_6102,N_3668,N_2865);
nand U6103 (N_6103,N_4328,N_4122);
nand U6104 (N_6104,N_3681,N_3185);
nor U6105 (N_6105,N_4311,N_4384);
and U6106 (N_6106,N_3630,N_2528);
nand U6107 (N_6107,N_3135,N_4391);
nor U6108 (N_6108,N_4096,N_4209);
nor U6109 (N_6109,N_2985,N_3857);
or U6110 (N_6110,N_3597,N_3964);
nand U6111 (N_6111,N_3228,N_4633);
or U6112 (N_6112,N_4348,N_2886);
nor U6113 (N_6113,N_4605,N_4706);
or U6114 (N_6114,N_4454,N_3943);
nand U6115 (N_6115,N_3146,N_3287);
nor U6116 (N_6116,N_3561,N_3337);
nand U6117 (N_6117,N_4131,N_4527);
nor U6118 (N_6118,N_2986,N_3291);
nand U6119 (N_6119,N_4106,N_4323);
nand U6120 (N_6120,N_2766,N_4202);
nand U6121 (N_6121,N_3652,N_4620);
or U6122 (N_6122,N_3952,N_3625);
xnor U6123 (N_6123,N_3769,N_2672);
or U6124 (N_6124,N_3696,N_3279);
or U6125 (N_6125,N_4761,N_4598);
nor U6126 (N_6126,N_3558,N_4185);
nor U6127 (N_6127,N_4822,N_3750);
nand U6128 (N_6128,N_4550,N_3209);
and U6129 (N_6129,N_4742,N_4159);
nand U6130 (N_6130,N_4339,N_3375);
nand U6131 (N_6131,N_4800,N_4006);
and U6132 (N_6132,N_4959,N_3776);
and U6133 (N_6133,N_3394,N_4484);
nor U6134 (N_6134,N_4708,N_4337);
and U6135 (N_6135,N_2921,N_3451);
or U6136 (N_6136,N_3270,N_2760);
nand U6137 (N_6137,N_3987,N_4539);
and U6138 (N_6138,N_2606,N_2687);
nand U6139 (N_6139,N_2795,N_3168);
or U6140 (N_6140,N_3145,N_2929);
nor U6141 (N_6141,N_2936,N_3834);
or U6142 (N_6142,N_3606,N_4657);
and U6143 (N_6143,N_4304,N_4329);
nor U6144 (N_6144,N_4556,N_3116);
or U6145 (N_6145,N_4429,N_3540);
nor U6146 (N_6146,N_4662,N_4412);
and U6147 (N_6147,N_3091,N_2783);
nand U6148 (N_6148,N_4332,N_3982);
nor U6149 (N_6149,N_3867,N_3946);
or U6150 (N_6150,N_3409,N_4886);
nand U6151 (N_6151,N_3669,N_4023);
nand U6152 (N_6152,N_4576,N_3620);
and U6153 (N_6153,N_2604,N_3562);
nand U6154 (N_6154,N_3161,N_3663);
or U6155 (N_6155,N_4781,N_4326);
nand U6156 (N_6156,N_2510,N_3904);
and U6157 (N_6157,N_4280,N_4401);
and U6158 (N_6158,N_3974,N_4489);
or U6159 (N_6159,N_4035,N_3199);
or U6160 (N_6160,N_2888,N_3240);
and U6161 (N_6161,N_2776,N_2716);
and U6162 (N_6162,N_4850,N_4020);
or U6163 (N_6163,N_4904,N_4069);
or U6164 (N_6164,N_4436,N_4668);
or U6165 (N_6165,N_3529,N_4768);
or U6166 (N_6166,N_3583,N_2571);
or U6167 (N_6167,N_2897,N_4587);
or U6168 (N_6168,N_4264,N_2987);
or U6169 (N_6169,N_4624,N_3938);
nor U6170 (N_6170,N_2781,N_4508);
or U6171 (N_6171,N_3047,N_4711);
nand U6172 (N_6172,N_4152,N_3594);
nor U6173 (N_6173,N_3127,N_3079);
nor U6174 (N_6174,N_3925,N_4562);
nand U6175 (N_6175,N_3847,N_3163);
or U6176 (N_6176,N_2585,N_4250);
or U6177 (N_6177,N_2941,N_3729);
nand U6178 (N_6178,N_2925,N_3986);
nand U6179 (N_6179,N_4046,N_3016);
and U6180 (N_6180,N_4710,N_4936);
or U6181 (N_6181,N_4216,N_3072);
or U6182 (N_6182,N_2931,N_4194);
nor U6183 (N_6183,N_3896,N_2561);
nor U6184 (N_6184,N_4913,N_4352);
nand U6185 (N_6185,N_4473,N_4606);
nand U6186 (N_6186,N_3961,N_4965);
nand U6187 (N_6187,N_3234,N_3462);
nand U6188 (N_6188,N_3015,N_4140);
nor U6189 (N_6189,N_4361,N_4350);
or U6190 (N_6190,N_2932,N_4962);
and U6191 (N_6191,N_3812,N_2572);
nor U6192 (N_6192,N_3809,N_3884);
nor U6193 (N_6193,N_3554,N_4666);
nor U6194 (N_6194,N_4677,N_3516);
nor U6195 (N_6195,N_3429,N_4376);
nand U6196 (N_6196,N_4279,N_4142);
nor U6197 (N_6197,N_4220,N_4770);
and U6198 (N_6198,N_4267,N_2742);
nand U6199 (N_6199,N_2502,N_3048);
nor U6200 (N_6200,N_3075,N_4390);
or U6201 (N_6201,N_4141,N_3478);
and U6202 (N_6202,N_3503,N_2670);
nor U6203 (N_6203,N_4377,N_4819);
and U6204 (N_6204,N_4272,N_3627);
nand U6205 (N_6205,N_2574,N_4935);
nand U6206 (N_6206,N_4782,N_2534);
and U6207 (N_6207,N_2539,N_4345);
nor U6208 (N_6208,N_4687,N_4169);
or U6209 (N_6209,N_3544,N_4425);
and U6210 (N_6210,N_3369,N_4789);
nor U6211 (N_6211,N_4922,N_4067);
nor U6212 (N_6212,N_3460,N_4171);
nor U6213 (N_6213,N_3021,N_3772);
or U6214 (N_6214,N_4571,N_4639);
or U6215 (N_6215,N_4732,N_2840);
nor U6216 (N_6216,N_4039,N_3504);
or U6217 (N_6217,N_4317,N_2752);
or U6218 (N_6218,N_3206,N_4669);
nand U6219 (N_6219,N_4181,N_3997);
and U6220 (N_6220,N_3983,N_3321);
and U6221 (N_6221,N_3511,N_3322);
or U6222 (N_6222,N_2508,N_4388);
and U6223 (N_6223,N_2909,N_3903);
nor U6224 (N_6224,N_3704,N_4466);
and U6225 (N_6225,N_3433,N_4162);
or U6226 (N_6226,N_4379,N_4660);
or U6227 (N_6227,N_3009,N_3736);
nor U6228 (N_6228,N_2874,N_3840);
nor U6229 (N_6229,N_3823,N_3112);
nor U6230 (N_6230,N_4702,N_3876);
nor U6231 (N_6231,N_4496,N_3774);
nor U6232 (N_6232,N_4747,N_3702);
nand U6233 (N_6233,N_2905,N_4052);
and U6234 (N_6234,N_3571,N_3271);
nand U6235 (N_6235,N_4968,N_4551);
or U6236 (N_6236,N_3790,N_3308);
and U6237 (N_6237,N_3018,N_3592);
nand U6238 (N_6238,N_4075,N_2770);
nor U6239 (N_6239,N_3895,N_3431);
or U6240 (N_6240,N_2983,N_3550);
nor U6241 (N_6241,N_4914,N_3930);
or U6242 (N_6242,N_4671,N_2794);
nand U6243 (N_6243,N_3762,N_3124);
nand U6244 (N_6244,N_3894,N_4034);
nand U6245 (N_6245,N_3870,N_3875);
nor U6246 (N_6246,N_2839,N_4004);
nor U6247 (N_6247,N_3664,N_4773);
nand U6248 (N_6248,N_4823,N_3507);
nor U6249 (N_6249,N_3761,N_2823);
and U6250 (N_6250,N_4084,N_3554);
or U6251 (N_6251,N_3715,N_2870);
and U6252 (N_6252,N_2863,N_4536);
and U6253 (N_6253,N_2555,N_4362);
nand U6254 (N_6254,N_3536,N_3210);
and U6255 (N_6255,N_4980,N_4401);
xor U6256 (N_6256,N_3095,N_4523);
nor U6257 (N_6257,N_3212,N_4535);
or U6258 (N_6258,N_2881,N_3242);
nor U6259 (N_6259,N_3746,N_3185);
nand U6260 (N_6260,N_3420,N_3240);
nand U6261 (N_6261,N_2608,N_3888);
nand U6262 (N_6262,N_3331,N_3237);
and U6263 (N_6263,N_3710,N_3295);
nor U6264 (N_6264,N_2786,N_4108);
or U6265 (N_6265,N_3576,N_2524);
and U6266 (N_6266,N_4273,N_3006);
or U6267 (N_6267,N_3526,N_4199);
nand U6268 (N_6268,N_2959,N_3266);
nand U6269 (N_6269,N_2971,N_3784);
nor U6270 (N_6270,N_4290,N_3925);
and U6271 (N_6271,N_4642,N_3958);
nor U6272 (N_6272,N_4844,N_3432);
and U6273 (N_6273,N_4247,N_3019);
and U6274 (N_6274,N_3670,N_2836);
nor U6275 (N_6275,N_4746,N_4139);
nor U6276 (N_6276,N_3537,N_4668);
or U6277 (N_6277,N_4297,N_4161);
xor U6278 (N_6278,N_4225,N_3235);
nand U6279 (N_6279,N_3447,N_2639);
nand U6280 (N_6280,N_3647,N_4320);
nor U6281 (N_6281,N_3216,N_3511);
nand U6282 (N_6282,N_3817,N_3986);
or U6283 (N_6283,N_4642,N_4748);
or U6284 (N_6284,N_3100,N_3503);
nor U6285 (N_6285,N_2661,N_2581);
nand U6286 (N_6286,N_2774,N_2813);
nand U6287 (N_6287,N_2622,N_4535);
or U6288 (N_6288,N_3265,N_4336);
nand U6289 (N_6289,N_3845,N_3734);
nand U6290 (N_6290,N_3837,N_3526);
or U6291 (N_6291,N_4282,N_2584);
and U6292 (N_6292,N_2598,N_3262);
and U6293 (N_6293,N_4181,N_2715);
nand U6294 (N_6294,N_3552,N_2948);
nand U6295 (N_6295,N_3835,N_4330);
nand U6296 (N_6296,N_4595,N_3188);
and U6297 (N_6297,N_2913,N_4679);
nor U6298 (N_6298,N_3421,N_4245);
or U6299 (N_6299,N_3406,N_3950);
nand U6300 (N_6300,N_3583,N_3593);
nor U6301 (N_6301,N_3872,N_3234);
nor U6302 (N_6302,N_4932,N_3924);
or U6303 (N_6303,N_4960,N_4789);
nand U6304 (N_6304,N_4371,N_3024);
nand U6305 (N_6305,N_4560,N_3516);
nor U6306 (N_6306,N_4061,N_4942);
and U6307 (N_6307,N_4521,N_3597);
or U6308 (N_6308,N_4609,N_3266);
nand U6309 (N_6309,N_2607,N_4811);
or U6310 (N_6310,N_4408,N_4024);
nand U6311 (N_6311,N_3122,N_3485);
and U6312 (N_6312,N_3418,N_2548);
nand U6313 (N_6313,N_2755,N_2806);
nand U6314 (N_6314,N_4810,N_3679);
and U6315 (N_6315,N_3046,N_3841);
and U6316 (N_6316,N_2997,N_4252);
nor U6317 (N_6317,N_2691,N_2922);
nor U6318 (N_6318,N_4805,N_3505);
nand U6319 (N_6319,N_4913,N_2648);
and U6320 (N_6320,N_2581,N_4192);
and U6321 (N_6321,N_3413,N_3794);
nand U6322 (N_6322,N_3745,N_4811);
and U6323 (N_6323,N_3250,N_4032);
nand U6324 (N_6324,N_2778,N_3467);
or U6325 (N_6325,N_3497,N_3314);
nand U6326 (N_6326,N_3698,N_3946);
nor U6327 (N_6327,N_2549,N_2705);
or U6328 (N_6328,N_3060,N_2505);
nand U6329 (N_6329,N_4627,N_4110);
and U6330 (N_6330,N_4287,N_2871);
nor U6331 (N_6331,N_4949,N_3185);
nand U6332 (N_6332,N_3453,N_3408);
and U6333 (N_6333,N_2686,N_4148);
nor U6334 (N_6334,N_2698,N_3364);
nor U6335 (N_6335,N_4982,N_4617);
and U6336 (N_6336,N_3659,N_2891);
nand U6337 (N_6337,N_3820,N_4781);
nor U6338 (N_6338,N_2756,N_3929);
nor U6339 (N_6339,N_4691,N_3765);
and U6340 (N_6340,N_4976,N_4527);
and U6341 (N_6341,N_2624,N_3200);
nor U6342 (N_6342,N_4880,N_3300);
nand U6343 (N_6343,N_3837,N_3353);
xor U6344 (N_6344,N_4263,N_4652);
or U6345 (N_6345,N_4834,N_4912);
nand U6346 (N_6346,N_3418,N_3381);
nand U6347 (N_6347,N_3037,N_4873);
and U6348 (N_6348,N_2791,N_4324);
and U6349 (N_6349,N_2613,N_3641);
or U6350 (N_6350,N_3652,N_3323);
nor U6351 (N_6351,N_3824,N_4856);
nand U6352 (N_6352,N_4789,N_4333);
nor U6353 (N_6353,N_3342,N_4874);
or U6354 (N_6354,N_3946,N_3021);
or U6355 (N_6355,N_3214,N_3445);
nor U6356 (N_6356,N_3436,N_4382);
nand U6357 (N_6357,N_2922,N_3139);
or U6358 (N_6358,N_3788,N_3297);
and U6359 (N_6359,N_4993,N_4504);
nand U6360 (N_6360,N_3746,N_2826);
and U6361 (N_6361,N_3707,N_4984);
nand U6362 (N_6362,N_3799,N_3247);
nor U6363 (N_6363,N_3499,N_4641);
nor U6364 (N_6364,N_3862,N_3429);
nor U6365 (N_6365,N_4036,N_4095);
xnor U6366 (N_6366,N_4277,N_2907);
and U6367 (N_6367,N_2629,N_3528);
nor U6368 (N_6368,N_3437,N_4775);
nor U6369 (N_6369,N_2734,N_4896);
or U6370 (N_6370,N_3333,N_3458);
or U6371 (N_6371,N_3344,N_4979);
or U6372 (N_6372,N_3897,N_4530);
and U6373 (N_6373,N_2655,N_3526);
nand U6374 (N_6374,N_2542,N_4691);
nand U6375 (N_6375,N_3355,N_2542);
or U6376 (N_6376,N_3486,N_3642);
and U6377 (N_6377,N_4715,N_2740);
nand U6378 (N_6378,N_3675,N_4950);
or U6379 (N_6379,N_3738,N_2844);
and U6380 (N_6380,N_2725,N_2992);
or U6381 (N_6381,N_3186,N_2590);
nor U6382 (N_6382,N_4683,N_4698);
nor U6383 (N_6383,N_3524,N_3669);
or U6384 (N_6384,N_2955,N_3423);
nand U6385 (N_6385,N_4418,N_3352);
nor U6386 (N_6386,N_2785,N_4097);
nand U6387 (N_6387,N_4227,N_3288);
nor U6388 (N_6388,N_4004,N_4988);
nor U6389 (N_6389,N_4921,N_3364);
xnor U6390 (N_6390,N_2676,N_4013);
nand U6391 (N_6391,N_3653,N_3065);
and U6392 (N_6392,N_3237,N_3343);
and U6393 (N_6393,N_2741,N_3750);
nand U6394 (N_6394,N_3138,N_2666);
nand U6395 (N_6395,N_4816,N_3818);
nor U6396 (N_6396,N_3192,N_2573);
and U6397 (N_6397,N_3854,N_2956);
nand U6398 (N_6398,N_3741,N_2645);
and U6399 (N_6399,N_3068,N_3906);
nand U6400 (N_6400,N_2880,N_3374);
or U6401 (N_6401,N_3748,N_3904);
nor U6402 (N_6402,N_2957,N_4064);
nor U6403 (N_6403,N_3490,N_2512);
nand U6404 (N_6404,N_2525,N_4647);
or U6405 (N_6405,N_3713,N_3343);
nand U6406 (N_6406,N_4418,N_4987);
or U6407 (N_6407,N_4387,N_2685);
nor U6408 (N_6408,N_3068,N_2742);
nand U6409 (N_6409,N_4645,N_3969);
nor U6410 (N_6410,N_3684,N_3849);
nand U6411 (N_6411,N_2837,N_2807);
nor U6412 (N_6412,N_3363,N_3073);
nor U6413 (N_6413,N_2735,N_2703);
and U6414 (N_6414,N_4820,N_3486);
nand U6415 (N_6415,N_4794,N_3081);
nor U6416 (N_6416,N_3479,N_3971);
nand U6417 (N_6417,N_2613,N_3698);
and U6418 (N_6418,N_3013,N_2879);
or U6419 (N_6419,N_4549,N_3547);
nor U6420 (N_6420,N_3328,N_2702);
or U6421 (N_6421,N_4916,N_3464);
nor U6422 (N_6422,N_3108,N_2755);
nor U6423 (N_6423,N_4231,N_3208);
nor U6424 (N_6424,N_4228,N_3357);
and U6425 (N_6425,N_4847,N_4407);
xor U6426 (N_6426,N_3436,N_4989);
nor U6427 (N_6427,N_3969,N_4255);
nand U6428 (N_6428,N_4067,N_3239);
or U6429 (N_6429,N_3095,N_4095);
nand U6430 (N_6430,N_4046,N_4868);
or U6431 (N_6431,N_4796,N_4893);
nand U6432 (N_6432,N_3406,N_4314);
xor U6433 (N_6433,N_3970,N_4447);
and U6434 (N_6434,N_3083,N_3730);
nand U6435 (N_6435,N_3324,N_2599);
and U6436 (N_6436,N_3904,N_4854);
and U6437 (N_6437,N_4758,N_2549);
and U6438 (N_6438,N_2816,N_3909);
or U6439 (N_6439,N_4708,N_3232);
nor U6440 (N_6440,N_2796,N_3345);
and U6441 (N_6441,N_2844,N_3227);
or U6442 (N_6442,N_3199,N_3938);
and U6443 (N_6443,N_3852,N_3609);
nand U6444 (N_6444,N_4520,N_2581);
nand U6445 (N_6445,N_2891,N_2979);
nand U6446 (N_6446,N_4917,N_3401);
and U6447 (N_6447,N_3386,N_4288);
or U6448 (N_6448,N_3227,N_3337);
nor U6449 (N_6449,N_4651,N_3453);
nor U6450 (N_6450,N_4182,N_3488);
nand U6451 (N_6451,N_4591,N_2601);
and U6452 (N_6452,N_3625,N_3856);
or U6453 (N_6453,N_3046,N_2718);
and U6454 (N_6454,N_2608,N_3929);
and U6455 (N_6455,N_2848,N_4018);
or U6456 (N_6456,N_3558,N_3244);
nor U6457 (N_6457,N_4225,N_2862);
nor U6458 (N_6458,N_3170,N_4378);
or U6459 (N_6459,N_3675,N_3433);
and U6460 (N_6460,N_3049,N_4568);
and U6461 (N_6461,N_2542,N_4524);
and U6462 (N_6462,N_3678,N_2961);
or U6463 (N_6463,N_4381,N_4909);
or U6464 (N_6464,N_4144,N_3580);
and U6465 (N_6465,N_3941,N_3106);
and U6466 (N_6466,N_4737,N_3660);
or U6467 (N_6467,N_4000,N_4502);
nand U6468 (N_6468,N_3373,N_4294);
nand U6469 (N_6469,N_4086,N_3584);
nand U6470 (N_6470,N_4270,N_4225);
or U6471 (N_6471,N_3600,N_4903);
nor U6472 (N_6472,N_3924,N_4077);
and U6473 (N_6473,N_4257,N_3824);
or U6474 (N_6474,N_3867,N_4867);
nand U6475 (N_6475,N_4323,N_4569);
nor U6476 (N_6476,N_3852,N_2635);
nor U6477 (N_6477,N_3139,N_3869);
or U6478 (N_6478,N_2846,N_2954);
nand U6479 (N_6479,N_4060,N_4840);
xnor U6480 (N_6480,N_4652,N_3204);
nand U6481 (N_6481,N_3958,N_3870);
or U6482 (N_6482,N_4307,N_4918);
xnor U6483 (N_6483,N_2938,N_3257);
nor U6484 (N_6484,N_2950,N_3759);
nand U6485 (N_6485,N_4840,N_4808);
and U6486 (N_6486,N_3387,N_2519);
nand U6487 (N_6487,N_2951,N_2732);
or U6488 (N_6488,N_4392,N_2774);
or U6489 (N_6489,N_4765,N_4361);
and U6490 (N_6490,N_3149,N_2737);
nand U6491 (N_6491,N_4872,N_3332);
nor U6492 (N_6492,N_2547,N_3086);
or U6493 (N_6493,N_2662,N_4020);
nor U6494 (N_6494,N_4701,N_4130);
and U6495 (N_6495,N_3922,N_3705);
or U6496 (N_6496,N_4413,N_4781);
and U6497 (N_6497,N_4722,N_2909);
nor U6498 (N_6498,N_3609,N_3214);
xor U6499 (N_6499,N_4373,N_4135);
and U6500 (N_6500,N_3728,N_4644);
nand U6501 (N_6501,N_4282,N_3949);
nand U6502 (N_6502,N_2508,N_2853);
or U6503 (N_6503,N_4605,N_3296);
or U6504 (N_6504,N_2739,N_2660);
and U6505 (N_6505,N_4969,N_4870);
and U6506 (N_6506,N_2731,N_3904);
nor U6507 (N_6507,N_4625,N_4282);
or U6508 (N_6508,N_4820,N_3692);
and U6509 (N_6509,N_4171,N_3495);
or U6510 (N_6510,N_4760,N_3197);
and U6511 (N_6511,N_4240,N_4286);
nor U6512 (N_6512,N_3722,N_2725);
nand U6513 (N_6513,N_3440,N_3975);
and U6514 (N_6514,N_4150,N_3851);
nand U6515 (N_6515,N_4552,N_3252);
nand U6516 (N_6516,N_2733,N_3848);
nor U6517 (N_6517,N_3463,N_3159);
nor U6518 (N_6518,N_2730,N_3964);
nand U6519 (N_6519,N_3844,N_3287);
or U6520 (N_6520,N_3719,N_4978);
and U6521 (N_6521,N_3326,N_4687);
nand U6522 (N_6522,N_4516,N_3488);
and U6523 (N_6523,N_4579,N_3879);
nand U6524 (N_6524,N_3093,N_4132);
or U6525 (N_6525,N_2830,N_4012);
and U6526 (N_6526,N_4345,N_3771);
nand U6527 (N_6527,N_3645,N_3266);
nand U6528 (N_6528,N_2732,N_3589);
nor U6529 (N_6529,N_4124,N_4049);
xnor U6530 (N_6530,N_2843,N_3156);
nand U6531 (N_6531,N_4200,N_4689);
nor U6532 (N_6532,N_3561,N_2522);
and U6533 (N_6533,N_2985,N_2765);
nand U6534 (N_6534,N_3776,N_4040);
or U6535 (N_6535,N_3389,N_4353);
or U6536 (N_6536,N_3940,N_3803);
or U6537 (N_6537,N_4865,N_3827);
or U6538 (N_6538,N_2635,N_2989);
nand U6539 (N_6539,N_4229,N_4159);
and U6540 (N_6540,N_4626,N_3555);
or U6541 (N_6541,N_3605,N_4585);
nor U6542 (N_6542,N_4840,N_2696);
nor U6543 (N_6543,N_3257,N_2557);
and U6544 (N_6544,N_4455,N_2939);
nor U6545 (N_6545,N_4298,N_2970);
or U6546 (N_6546,N_4024,N_4532);
nand U6547 (N_6547,N_4895,N_4266);
and U6548 (N_6548,N_4396,N_2789);
and U6549 (N_6549,N_4348,N_2814);
and U6550 (N_6550,N_4338,N_3534);
or U6551 (N_6551,N_4310,N_3655);
nor U6552 (N_6552,N_4033,N_3807);
nand U6553 (N_6553,N_3516,N_3198);
and U6554 (N_6554,N_3295,N_4362);
nand U6555 (N_6555,N_2818,N_3089);
nand U6556 (N_6556,N_4837,N_2572);
nand U6557 (N_6557,N_4935,N_2980);
or U6558 (N_6558,N_3769,N_4459);
nor U6559 (N_6559,N_3690,N_4517);
nor U6560 (N_6560,N_3186,N_2545);
or U6561 (N_6561,N_4978,N_4254);
and U6562 (N_6562,N_3422,N_2673);
nor U6563 (N_6563,N_3517,N_4171);
nor U6564 (N_6564,N_3172,N_4318);
or U6565 (N_6565,N_4403,N_2832);
and U6566 (N_6566,N_4901,N_2545);
and U6567 (N_6567,N_4895,N_4819);
nor U6568 (N_6568,N_4778,N_2716);
nand U6569 (N_6569,N_3070,N_3489);
or U6570 (N_6570,N_4343,N_4333);
or U6571 (N_6571,N_4683,N_4521);
nand U6572 (N_6572,N_3660,N_3562);
nor U6573 (N_6573,N_4621,N_3326);
nand U6574 (N_6574,N_4087,N_4326);
nand U6575 (N_6575,N_2994,N_3995);
nor U6576 (N_6576,N_2707,N_3624);
nand U6577 (N_6577,N_4991,N_3813);
and U6578 (N_6578,N_4433,N_4745);
or U6579 (N_6579,N_3787,N_4585);
or U6580 (N_6580,N_2820,N_2897);
nor U6581 (N_6581,N_3765,N_3446);
and U6582 (N_6582,N_4020,N_4697);
or U6583 (N_6583,N_3500,N_4531);
and U6584 (N_6584,N_2901,N_4762);
and U6585 (N_6585,N_3190,N_3653);
and U6586 (N_6586,N_3542,N_4361);
nand U6587 (N_6587,N_3529,N_4362);
nor U6588 (N_6588,N_3791,N_3076);
nor U6589 (N_6589,N_3366,N_3746);
nor U6590 (N_6590,N_2781,N_4140);
and U6591 (N_6591,N_4270,N_4612);
and U6592 (N_6592,N_2922,N_2717);
nand U6593 (N_6593,N_3153,N_4893);
or U6594 (N_6594,N_4082,N_4260);
xor U6595 (N_6595,N_2821,N_3060);
and U6596 (N_6596,N_2997,N_4274);
nand U6597 (N_6597,N_3585,N_4169);
nand U6598 (N_6598,N_4271,N_2657);
nor U6599 (N_6599,N_4669,N_4499);
and U6600 (N_6600,N_3660,N_3084);
or U6601 (N_6601,N_3342,N_4790);
nor U6602 (N_6602,N_4327,N_3559);
and U6603 (N_6603,N_2916,N_4848);
nor U6604 (N_6604,N_4682,N_2706);
or U6605 (N_6605,N_4585,N_3699);
nor U6606 (N_6606,N_3684,N_3185);
and U6607 (N_6607,N_4403,N_3915);
nand U6608 (N_6608,N_2932,N_2645);
nand U6609 (N_6609,N_4341,N_2708);
and U6610 (N_6610,N_3669,N_3138);
nand U6611 (N_6611,N_4123,N_3317);
and U6612 (N_6612,N_4379,N_3519);
nand U6613 (N_6613,N_3570,N_4297);
nor U6614 (N_6614,N_3286,N_2992);
nand U6615 (N_6615,N_2864,N_4982);
nor U6616 (N_6616,N_2839,N_3333);
nand U6617 (N_6617,N_4530,N_4442);
nor U6618 (N_6618,N_3086,N_3418);
and U6619 (N_6619,N_2801,N_2713);
nor U6620 (N_6620,N_4734,N_3449);
or U6621 (N_6621,N_3032,N_2946);
and U6622 (N_6622,N_4785,N_4586);
nor U6623 (N_6623,N_3406,N_3853);
or U6624 (N_6624,N_4372,N_2851);
nand U6625 (N_6625,N_4994,N_4533);
or U6626 (N_6626,N_3730,N_3554);
nor U6627 (N_6627,N_4618,N_4909);
nand U6628 (N_6628,N_4483,N_2954);
nor U6629 (N_6629,N_4160,N_4775);
nand U6630 (N_6630,N_4327,N_4355);
nor U6631 (N_6631,N_4867,N_3346);
or U6632 (N_6632,N_2939,N_3857);
nand U6633 (N_6633,N_3059,N_4858);
and U6634 (N_6634,N_3280,N_4474);
nand U6635 (N_6635,N_3582,N_2988);
nand U6636 (N_6636,N_4977,N_4840);
or U6637 (N_6637,N_4486,N_2501);
nand U6638 (N_6638,N_4349,N_4926);
nor U6639 (N_6639,N_3987,N_4552);
nand U6640 (N_6640,N_3201,N_2611);
nor U6641 (N_6641,N_4138,N_2849);
and U6642 (N_6642,N_2718,N_2726);
and U6643 (N_6643,N_3761,N_4259);
nor U6644 (N_6644,N_2738,N_4748);
and U6645 (N_6645,N_2886,N_3496);
and U6646 (N_6646,N_4509,N_2989);
and U6647 (N_6647,N_2741,N_3276);
nand U6648 (N_6648,N_4882,N_4875);
nor U6649 (N_6649,N_3941,N_3982);
nor U6650 (N_6650,N_2769,N_3927);
or U6651 (N_6651,N_3332,N_3537);
nand U6652 (N_6652,N_4545,N_3664);
and U6653 (N_6653,N_4632,N_4949);
and U6654 (N_6654,N_4413,N_4021);
and U6655 (N_6655,N_4848,N_3856);
or U6656 (N_6656,N_4842,N_3456);
nor U6657 (N_6657,N_4371,N_4854);
or U6658 (N_6658,N_3586,N_3388);
and U6659 (N_6659,N_4126,N_3239);
nor U6660 (N_6660,N_4634,N_3688);
and U6661 (N_6661,N_3819,N_4848);
nand U6662 (N_6662,N_4160,N_3788);
or U6663 (N_6663,N_3228,N_2737);
nor U6664 (N_6664,N_2879,N_2897);
or U6665 (N_6665,N_2535,N_4555);
nand U6666 (N_6666,N_4691,N_3149);
and U6667 (N_6667,N_4496,N_4082);
or U6668 (N_6668,N_4718,N_4042);
nor U6669 (N_6669,N_3843,N_4624);
nor U6670 (N_6670,N_4075,N_3498);
nand U6671 (N_6671,N_4670,N_2994);
nand U6672 (N_6672,N_4968,N_4772);
and U6673 (N_6673,N_4988,N_4306);
and U6674 (N_6674,N_4873,N_3224);
nor U6675 (N_6675,N_4990,N_2565);
or U6676 (N_6676,N_4160,N_4847);
xnor U6677 (N_6677,N_4678,N_3666);
nor U6678 (N_6678,N_3822,N_2618);
and U6679 (N_6679,N_3197,N_3227);
nand U6680 (N_6680,N_3082,N_3127);
or U6681 (N_6681,N_2946,N_4251);
nand U6682 (N_6682,N_4428,N_3096);
or U6683 (N_6683,N_4254,N_2779);
or U6684 (N_6684,N_3830,N_2519);
nand U6685 (N_6685,N_4987,N_3006);
nand U6686 (N_6686,N_4705,N_3831);
nor U6687 (N_6687,N_4114,N_4555);
and U6688 (N_6688,N_3363,N_3414);
nor U6689 (N_6689,N_3655,N_3238);
and U6690 (N_6690,N_3648,N_4084);
nor U6691 (N_6691,N_4205,N_2643);
nor U6692 (N_6692,N_4291,N_4967);
nand U6693 (N_6693,N_2642,N_4674);
or U6694 (N_6694,N_3030,N_3908);
and U6695 (N_6695,N_3615,N_2625);
or U6696 (N_6696,N_3770,N_4615);
nand U6697 (N_6697,N_2861,N_4559);
and U6698 (N_6698,N_3271,N_2669);
nand U6699 (N_6699,N_3119,N_3484);
nor U6700 (N_6700,N_4304,N_3313);
and U6701 (N_6701,N_3977,N_3483);
nand U6702 (N_6702,N_2665,N_3646);
nand U6703 (N_6703,N_3393,N_3452);
or U6704 (N_6704,N_3473,N_2994);
nor U6705 (N_6705,N_3726,N_4791);
nand U6706 (N_6706,N_4255,N_3597);
nor U6707 (N_6707,N_4930,N_4530);
nand U6708 (N_6708,N_3181,N_3881);
or U6709 (N_6709,N_4559,N_4046);
nor U6710 (N_6710,N_2860,N_4525);
or U6711 (N_6711,N_4421,N_3301);
nand U6712 (N_6712,N_4418,N_4794);
nand U6713 (N_6713,N_2889,N_3363);
nand U6714 (N_6714,N_3811,N_4492);
or U6715 (N_6715,N_2829,N_3073);
or U6716 (N_6716,N_4088,N_4052);
nand U6717 (N_6717,N_3886,N_3749);
and U6718 (N_6718,N_4310,N_4680);
and U6719 (N_6719,N_4290,N_2911);
and U6720 (N_6720,N_2599,N_4828);
or U6721 (N_6721,N_4124,N_4759);
or U6722 (N_6722,N_3213,N_4786);
and U6723 (N_6723,N_2500,N_3247);
and U6724 (N_6724,N_3805,N_3777);
and U6725 (N_6725,N_4947,N_4471);
nand U6726 (N_6726,N_2571,N_4025);
nor U6727 (N_6727,N_2754,N_4206);
nand U6728 (N_6728,N_4866,N_2535);
and U6729 (N_6729,N_4144,N_3636);
or U6730 (N_6730,N_2788,N_3509);
nor U6731 (N_6731,N_2537,N_3314);
nand U6732 (N_6732,N_3976,N_3947);
nand U6733 (N_6733,N_4747,N_2560);
or U6734 (N_6734,N_4171,N_4303);
or U6735 (N_6735,N_3566,N_3087);
or U6736 (N_6736,N_3033,N_4464);
nor U6737 (N_6737,N_3793,N_3745);
nand U6738 (N_6738,N_2716,N_4528);
nor U6739 (N_6739,N_3022,N_3256);
nand U6740 (N_6740,N_3279,N_2633);
or U6741 (N_6741,N_3818,N_3261);
or U6742 (N_6742,N_3741,N_3564);
and U6743 (N_6743,N_3747,N_2830);
and U6744 (N_6744,N_2659,N_4210);
nor U6745 (N_6745,N_2914,N_4694);
nand U6746 (N_6746,N_3789,N_3153);
and U6747 (N_6747,N_3624,N_2595);
or U6748 (N_6748,N_4613,N_3386);
nor U6749 (N_6749,N_3673,N_4609);
or U6750 (N_6750,N_3439,N_4674);
or U6751 (N_6751,N_4200,N_4686);
and U6752 (N_6752,N_3958,N_2718);
or U6753 (N_6753,N_4162,N_2869);
or U6754 (N_6754,N_2539,N_3690);
or U6755 (N_6755,N_2723,N_3041);
nor U6756 (N_6756,N_3068,N_3997);
nand U6757 (N_6757,N_2869,N_3033);
and U6758 (N_6758,N_2750,N_3967);
and U6759 (N_6759,N_4641,N_2583);
nor U6760 (N_6760,N_4262,N_2921);
or U6761 (N_6761,N_4861,N_3452);
and U6762 (N_6762,N_3242,N_4240);
nand U6763 (N_6763,N_3001,N_2558);
or U6764 (N_6764,N_3165,N_4305);
or U6765 (N_6765,N_2804,N_3234);
or U6766 (N_6766,N_3586,N_2604);
nand U6767 (N_6767,N_4648,N_3575);
nand U6768 (N_6768,N_3274,N_2669);
and U6769 (N_6769,N_3686,N_4660);
nand U6770 (N_6770,N_3246,N_2801);
nand U6771 (N_6771,N_4766,N_2740);
nand U6772 (N_6772,N_3335,N_4952);
xnor U6773 (N_6773,N_2812,N_4532);
and U6774 (N_6774,N_4082,N_2698);
nor U6775 (N_6775,N_4268,N_4929);
nand U6776 (N_6776,N_3936,N_3216);
nand U6777 (N_6777,N_4250,N_4247);
and U6778 (N_6778,N_4575,N_4982);
nor U6779 (N_6779,N_4013,N_2647);
or U6780 (N_6780,N_4136,N_3289);
or U6781 (N_6781,N_3393,N_2929);
or U6782 (N_6782,N_3747,N_4150);
xor U6783 (N_6783,N_4448,N_3064);
or U6784 (N_6784,N_2764,N_3220);
nor U6785 (N_6785,N_4930,N_3822);
nand U6786 (N_6786,N_4429,N_2543);
and U6787 (N_6787,N_4394,N_2968);
and U6788 (N_6788,N_3185,N_3432);
nand U6789 (N_6789,N_3136,N_3953);
and U6790 (N_6790,N_3633,N_2586);
nor U6791 (N_6791,N_4399,N_2798);
nand U6792 (N_6792,N_4986,N_2525);
or U6793 (N_6793,N_4730,N_2961);
nand U6794 (N_6794,N_3604,N_4360);
and U6795 (N_6795,N_2761,N_3669);
or U6796 (N_6796,N_4139,N_2773);
or U6797 (N_6797,N_3115,N_4885);
nand U6798 (N_6798,N_2511,N_4120);
nand U6799 (N_6799,N_4263,N_4351);
or U6800 (N_6800,N_2902,N_2941);
or U6801 (N_6801,N_4423,N_4524);
nand U6802 (N_6802,N_2524,N_3465);
or U6803 (N_6803,N_2569,N_4207);
and U6804 (N_6804,N_3732,N_3497);
or U6805 (N_6805,N_4142,N_2901);
or U6806 (N_6806,N_4145,N_4391);
nand U6807 (N_6807,N_4551,N_3929);
nor U6808 (N_6808,N_3461,N_2732);
or U6809 (N_6809,N_4674,N_3953);
or U6810 (N_6810,N_2988,N_4885);
and U6811 (N_6811,N_3341,N_3634);
or U6812 (N_6812,N_2981,N_4200);
and U6813 (N_6813,N_2767,N_4972);
nand U6814 (N_6814,N_3618,N_4716);
nand U6815 (N_6815,N_3542,N_2566);
and U6816 (N_6816,N_3700,N_3496);
nand U6817 (N_6817,N_3457,N_3054);
and U6818 (N_6818,N_3357,N_4515);
or U6819 (N_6819,N_4749,N_3837);
and U6820 (N_6820,N_3263,N_3245);
or U6821 (N_6821,N_3385,N_3831);
and U6822 (N_6822,N_3934,N_4550);
or U6823 (N_6823,N_3237,N_3088);
and U6824 (N_6824,N_3483,N_3539);
or U6825 (N_6825,N_3501,N_4944);
nor U6826 (N_6826,N_4039,N_4281);
nand U6827 (N_6827,N_4941,N_2714);
nand U6828 (N_6828,N_2647,N_3821);
nand U6829 (N_6829,N_2954,N_3176);
or U6830 (N_6830,N_4276,N_3262);
or U6831 (N_6831,N_4255,N_4138);
nor U6832 (N_6832,N_4761,N_3494);
or U6833 (N_6833,N_2505,N_4356);
or U6834 (N_6834,N_2806,N_4425);
or U6835 (N_6835,N_2699,N_4890);
and U6836 (N_6836,N_3856,N_4020);
or U6837 (N_6837,N_2877,N_4897);
nand U6838 (N_6838,N_3452,N_2919);
nand U6839 (N_6839,N_4544,N_4127);
and U6840 (N_6840,N_4122,N_3217);
nand U6841 (N_6841,N_3925,N_2941);
or U6842 (N_6842,N_2514,N_3736);
nand U6843 (N_6843,N_2980,N_3887);
nor U6844 (N_6844,N_2670,N_4868);
nand U6845 (N_6845,N_4703,N_4771);
and U6846 (N_6846,N_3199,N_4371);
nor U6847 (N_6847,N_4516,N_4217);
and U6848 (N_6848,N_3658,N_3910);
and U6849 (N_6849,N_2503,N_4179);
and U6850 (N_6850,N_3718,N_3617);
or U6851 (N_6851,N_3176,N_4086);
or U6852 (N_6852,N_2551,N_4973);
nand U6853 (N_6853,N_4620,N_3278);
and U6854 (N_6854,N_3604,N_4407);
and U6855 (N_6855,N_3281,N_3530);
or U6856 (N_6856,N_4377,N_3788);
nand U6857 (N_6857,N_2975,N_3590);
and U6858 (N_6858,N_4627,N_2762);
and U6859 (N_6859,N_3564,N_4184);
nand U6860 (N_6860,N_2786,N_4642);
and U6861 (N_6861,N_3243,N_4807);
nand U6862 (N_6862,N_4114,N_4303);
or U6863 (N_6863,N_4506,N_3509);
nand U6864 (N_6864,N_2608,N_3162);
and U6865 (N_6865,N_4752,N_3590);
and U6866 (N_6866,N_3147,N_2625);
nand U6867 (N_6867,N_3194,N_2611);
nor U6868 (N_6868,N_4883,N_2538);
or U6869 (N_6869,N_4653,N_2799);
and U6870 (N_6870,N_4709,N_2862);
nor U6871 (N_6871,N_2515,N_3251);
or U6872 (N_6872,N_4969,N_4048);
or U6873 (N_6873,N_3727,N_3827);
or U6874 (N_6874,N_3486,N_3554);
and U6875 (N_6875,N_3455,N_3638);
nand U6876 (N_6876,N_4048,N_3808);
nor U6877 (N_6877,N_2974,N_3528);
or U6878 (N_6878,N_4036,N_4175);
or U6879 (N_6879,N_3664,N_2831);
nor U6880 (N_6880,N_3576,N_2977);
and U6881 (N_6881,N_3015,N_4658);
nor U6882 (N_6882,N_3390,N_4931);
or U6883 (N_6883,N_3584,N_2542);
nor U6884 (N_6884,N_3348,N_4304);
nand U6885 (N_6885,N_3041,N_4256);
nor U6886 (N_6886,N_3532,N_4838);
and U6887 (N_6887,N_4328,N_2841);
and U6888 (N_6888,N_4475,N_3838);
nand U6889 (N_6889,N_3853,N_3770);
nor U6890 (N_6890,N_2621,N_2943);
nand U6891 (N_6891,N_3358,N_4028);
or U6892 (N_6892,N_3311,N_2521);
nor U6893 (N_6893,N_4761,N_4817);
and U6894 (N_6894,N_2975,N_2699);
and U6895 (N_6895,N_3819,N_3459);
and U6896 (N_6896,N_4069,N_4133);
and U6897 (N_6897,N_4537,N_3994);
or U6898 (N_6898,N_3164,N_4419);
nor U6899 (N_6899,N_3273,N_3540);
xnor U6900 (N_6900,N_2562,N_4322);
or U6901 (N_6901,N_2645,N_4564);
and U6902 (N_6902,N_3879,N_4388);
and U6903 (N_6903,N_2762,N_4646);
or U6904 (N_6904,N_4127,N_3255);
nand U6905 (N_6905,N_3352,N_4440);
and U6906 (N_6906,N_3014,N_3486);
or U6907 (N_6907,N_2784,N_3527);
nand U6908 (N_6908,N_2508,N_4373);
or U6909 (N_6909,N_3686,N_3057);
nor U6910 (N_6910,N_4249,N_3172);
nor U6911 (N_6911,N_4239,N_2722);
or U6912 (N_6912,N_3369,N_3078);
xor U6913 (N_6913,N_3149,N_2927);
and U6914 (N_6914,N_3986,N_3555);
nor U6915 (N_6915,N_2894,N_3844);
nor U6916 (N_6916,N_2674,N_2600);
nor U6917 (N_6917,N_4216,N_2573);
nor U6918 (N_6918,N_3686,N_3799);
and U6919 (N_6919,N_4431,N_3170);
and U6920 (N_6920,N_3525,N_4742);
nand U6921 (N_6921,N_4568,N_2820);
or U6922 (N_6922,N_4090,N_4266);
nand U6923 (N_6923,N_3922,N_3874);
nor U6924 (N_6924,N_3899,N_4814);
xor U6925 (N_6925,N_4773,N_4095);
or U6926 (N_6926,N_2984,N_2957);
or U6927 (N_6927,N_2559,N_2650);
or U6928 (N_6928,N_4512,N_3654);
nand U6929 (N_6929,N_4768,N_2549);
nor U6930 (N_6930,N_2944,N_2796);
and U6931 (N_6931,N_4519,N_4291);
or U6932 (N_6932,N_4083,N_2641);
or U6933 (N_6933,N_3999,N_4429);
nor U6934 (N_6934,N_4153,N_4629);
nor U6935 (N_6935,N_4127,N_3144);
nand U6936 (N_6936,N_4099,N_4329);
nor U6937 (N_6937,N_4106,N_4991);
nand U6938 (N_6938,N_3731,N_3982);
nor U6939 (N_6939,N_3450,N_4182);
nor U6940 (N_6940,N_4929,N_3764);
nor U6941 (N_6941,N_4393,N_3111);
or U6942 (N_6942,N_4397,N_3088);
and U6943 (N_6943,N_4627,N_2968);
nor U6944 (N_6944,N_4098,N_4878);
nor U6945 (N_6945,N_4224,N_3574);
nand U6946 (N_6946,N_3665,N_3747);
nor U6947 (N_6947,N_4440,N_3612);
or U6948 (N_6948,N_2716,N_3613);
nand U6949 (N_6949,N_4347,N_3628);
nand U6950 (N_6950,N_4607,N_3577);
nor U6951 (N_6951,N_4408,N_3712);
and U6952 (N_6952,N_3774,N_4905);
xnor U6953 (N_6953,N_3687,N_3029);
and U6954 (N_6954,N_3629,N_4034);
and U6955 (N_6955,N_4876,N_2648);
or U6956 (N_6956,N_3363,N_3784);
nand U6957 (N_6957,N_2697,N_4999);
or U6958 (N_6958,N_3935,N_4324);
nand U6959 (N_6959,N_3951,N_3705);
nor U6960 (N_6960,N_4744,N_4380);
nand U6961 (N_6961,N_2784,N_2707);
or U6962 (N_6962,N_4086,N_3745);
and U6963 (N_6963,N_2760,N_4029);
nor U6964 (N_6964,N_2619,N_3897);
nor U6965 (N_6965,N_3030,N_3312);
or U6966 (N_6966,N_4101,N_2910);
or U6967 (N_6967,N_2777,N_3047);
or U6968 (N_6968,N_4154,N_3445);
nand U6969 (N_6969,N_4933,N_4450);
nand U6970 (N_6970,N_2697,N_3943);
and U6971 (N_6971,N_4012,N_2670);
or U6972 (N_6972,N_2552,N_4204);
nand U6973 (N_6973,N_4684,N_4716);
and U6974 (N_6974,N_4945,N_4205);
and U6975 (N_6975,N_3004,N_4044);
nand U6976 (N_6976,N_3376,N_2799);
nand U6977 (N_6977,N_4639,N_3372);
nand U6978 (N_6978,N_4161,N_4652);
and U6979 (N_6979,N_2861,N_3051);
nand U6980 (N_6980,N_4506,N_2849);
and U6981 (N_6981,N_3743,N_3261);
and U6982 (N_6982,N_4683,N_2987);
or U6983 (N_6983,N_3297,N_4901);
and U6984 (N_6984,N_3607,N_4618);
nor U6985 (N_6985,N_2583,N_2606);
or U6986 (N_6986,N_4758,N_2571);
or U6987 (N_6987,N_4965,N_3782);
or U6988 (N_6988,N_4725,N_3108);
and U6989 (N_6989,N_4583,N_4725);
or U6990 (N_6990,N_4727,N_3904);
nand U6991 (N_6991,N_3989,N_4195);
nor U6992 (N_6992,N_4179,N_2729);
nor U6993 (N_6993,N_3439,N_3950);
or U6994 (N_6994,N_2584,N_3475);
nand U6995 (N_6995,N_2519,N_4762);
nor U6996 (N_6996,N_4951,N_2550);
nand U6997 (N_6997,N_3112,N_4399);
nand U6998 (N_6998,N_4379,N_3864);
nand U6999 (N_6999,N_2848,N_3206);
nand U7000 (N_7000,N_4735,N_3880);
nor U7001 (N_7001,N_3207,N_3004);
nor U7002 (N_7002,N_4394,N_2783);
nand U7003 (N_7003,N_4433,N_4427);
and U7004 (N_7004,N_4484,N_4679);
and U7005 (N_7005,N_4870,N_2950);
or U7006 (N_7006,N_3903,N_3209);
and U7007 (N_7007,N_2954,N_4645);
nand U7008 (N_7008,N_4914,N_3578);
nand U7009 (N_7009,N_3834,N_4162);
nor U7010 (N_7010,N_3584,N_3664);
nor U7011 (N_7011,N_3977,N_3857);
and U7012 (N_7012,N_3267,N_4920);
and U7013 (N_7013,N_3941,N_4678);
nor U7014 (N_7014,N_2685,N_3597);
nor U7015 (N_7015,N_4782,N_4130);
or U7016 (N_7016,N_3189,N_4664);
and U7017 (N_7017,N_3341,N_4056);
nor U7018 (N_7018,N_3681,N_3230);
nand U7019 (N_7019,N_4381,N_4290);
nand U7020 (N_7020,N_2987,N_4674);
and U7021 (N_7021,N_2998,N_2857);
and U7022 (N_7022,N_4545,N_3350);
and U7023 (N_7023,N_3186,N_3173);
and U7024 (N_7024,N_4390,N_3279);
and U7025 (N_7025,N_3709,N_3511);
nor U7026 (N_7026,N_3344,N_3057);
or U7027 (N_7027,N_4187,N_3700);
nor U7028 (N_7028,N_3744,N_3860);
and U7029 (N_7029,N_4871,N_3451);
nor U7030 (N_7030,N_2500,N_3423);
nor U7031 (N_7031,N_2972,N_4441);
nor U7032 (N_7032,N_4458,N_3595);
and U7033 (N_7033,N_3356,N_3693);
nor U7034 (N_7034,N_4139,N_4909);
nor U7035 (N_7035,N_3983,N_4607);
or U7036 (N_7036,N_4903,N_4288);
or U7037 (N_7037,N_4279,N_4299);
nor U7038 (N_7038,N_2745,N_3300);
and U7039 (N_7039,N_4701,N_3543);
nor U7040 (N_7040,N_4905,N_3723);
and U7041 (N_7041,N_4662,N_3487);
nor U7042 (N_7042,N_4348,N_3953);
and U7043 (N_7043,N_4861,N_4410);
nand U7044 (N_7044,N_4004,N_3506);
and U7045 (N_7045,N_4365,N_4210);
nor U7046 (N_7046,N_3396,N_2627);
or U7047 (N_7047,N_4693,N_4444);
nand U7048 (N_7048,N_4590,N_4605);
nand U7049 (N_7049,N_2613,N_3384);
nor U7050 (N_7050,N_4898,N_4333);
and U7051 (N_7051,N_4926,N_3303);
and U7052 (N_7052,N_3274,N_3670);
and U7053 (N_7053,N_4532,N_4323);
or U7054 (N_7054,N_2644,N_2640);
nor U7055 (N_7055,N_4346,N_3346);
nand U7056 (N_7056,N_4474,N_3412);
and U7057 (N_7057,N_4437,N_3662);
nand U7058 (N_7058,N_3039,N_4535);
nor U7059 (N_7059,N_2863,N_2827);
or U7060 (N_7060,N_3668,N_4568);
and U7061 (N_7061,N_4422,N_2911);
nand U7062 (N_7062,N_2864,N_3105);
or U7063 (N_7063,N_2986,N_3121);
nand U7064 (N_7064,N_3921,N_4522);
nor U7065 (N_7065,N_3205,N_3517);
and U7066 (N_7066,N_4229,N_3538);
or U7067 (N_7067,N_3779,N_2548);
or U7068 (N_7068,N_4484,N_4432);
or U7069 (N_7069,N_3270,N_4916);
or U7070 (N_7070,N_4623,N_4469);
nand U7071 (N_7071,N_3808,N_2660);
nand U7072 (N_7072,N_3181,N_4588);
nand U7073 (N_7073,N_3552,N_3080);
or U7074 (N_7074,N_3667,N_2526);
or U7075 (N_7075,N_2802,N_2952);
or U7076 (N_7076,N_3242,N_2830);
and U7077 (N_7077,N_4353,N_4516);
or U7078 (N_7078,N_2851,N_4127);
nor U7079 (N_7079,N_3760,N_4502);
or U7080 (N_7080,N_2852,N_3856);
or U7081 (N_7081,N_4594,N_4410);
nand U7082 (N_7082,N_4686,N_4727);
nand U7083 (N_7083,N_3045,N_4622);
nor U7084 (N_7084,N_3753,N_2677);
nand U7085 (N_7085,N_4864,N_2706);
nor U7086 (N_7086,N_4435,N_2801);
or U7087 (N_7087,N_3168,N_4904);
or U7088 (N_7088,N_4166,N_4347);
nand U7089 (N_7089,N_4494,N_4261);
and U7090 (N_7090,N_3960,N_3401);
or U7091 (N_7091,N_2624,N_4472);
and U7092 (N_7092,N_4883,N_3698);
nand U7093 (N_7093,N_3321,N_4323);
nor U7094 (N_7094,N_3331,N_3596);
nor U7095 (N_7095,N_3338,N_4112);
or U7096 (N_7096,N_3605,N_4052);
or U7097 (N_7097,N_2556,N_3542);
nand U7098 (N_7098,N_3413,N_3751);
and U7099 (N_7099,N_4654,N_4763);
and U7100 (N_7100,N_3943,N_4940);
or U7101 (N_7101,N_3945,N_2789);
or U7102 (N_7102,N_3966,N_3512);
or U7103 (N_7103,N_2716,N_2880);
nand U7104 (N_7104,N_4676,N_3533);
and U7105 (N_7105,N_4443,N_2995);
nand U7106 (N_7106,N_3704,N_3088);
nor U7107 (N_7107,N_3521,N_3176);
xnor U7108 (N_7108,N_4248,N_4205);
nor U7109 (N_7109,N_3308,N_4463);
nand U7110 (N_7110,N_2928,N_2906);
nand U7111 (N_7111,N_4374,N_3147);
and U7112 (N_7112,N_4887,N_3481);
nand U7113 (N_7113,N_2929,N_4050);
or U7114 (N_7114,N_4875,N_2973);
nor U7115 (N_7115,N_4478,N_2594);
or U7116 (N_7116,N_4247,N_3193);
and U7117 (N_7117,N_2677,N_2848);
and U7118 (N_7118,N_3968,N_2966);
or U7119 (N_7119,N_4236,N_2791);
or U7120 (N_7120,N_3246,N_3063);
or U7121 (N_7121,N_3990,N_2802);
and U7122 (N_7122,N_3371,N_4791);
or U7123 (N_7123,N_2673,N_3986);
nand U7124 (N_7124,N_4023,N_3166);
and U7125 (N_7125,N_3536,N_4007);
or U7126 (N_7126,N_3902,N_3277);
nand U7127 (N_7127,N_4304,N_3069);
nand U7128 (N_7128,N_4948,N_4417);
and U7129 (N_7129,N_3598,N_3981);
nor U7130 (N_7130,N_4719,N_3325);
or U7131 (N_7131,N_4149,N_3503);
and U7132 (N_7132,N_4460,N_2611);
nand U7133 (N_7133,N_4963,N_3160);
nand U7134 (N_7134,N_3906,N_3406);
nand U7135 (N_7135,N_3769,N_3693);
nor U7136 (N_7136,N_3269,N_4637);
nor U7137 (N_7137,N_3471,N_4867);
and U7138 (N_7138,N_4536,N_2959);
or U7139 (N_7139,N_3499,N_4501);
nor U7140 (N_7140,N_4671,N_4228);
nor U7141 (N_7141,N_2803,N_4930);
and U7142 (N_7142,N_2616,N_2927);
nor U7143 (N_7143,N_4715,N_4760);
and U7144 (N_7144,N_2903,N_3607);
nor U7145 (N_7145,N_3462,N_4892);
nand U7146 (N_7146,N_4701,N_2741);
and U7147 (N_7147,N_4843,N_3215);
or U7148 (N_7148,N_3418,N_2876);
and U7149 (N_7149,N_3967,N_3943);
or U7150 (N_7150,N_4528,N_2683);
or U7151 (N_7151,N_2834,N_4052);
or U7152 (N_7152,N_4047,N_2767);
and U7153 (N_7153,N_4017,N_3052);
nor U7154 (N_7154,N_4206,N_3287);
or U7155 (N_7155,N_3348,N_4144);
nand U7156 (N_7156,N_4219,N_3254);
and U7157 (N_7157,N_4809,N_4487);
nor U7158 (N_7158,N_4000,N_3545);
and U7159 (N_7159,N_2940,N_4469);
nand U7160 (N_7160,N_4858,N_3612);
and U7161 (N_7161,N_4945,N_3922);
nand U7162 (N_7162,N_2573,N_4421);
or U7163 (N_7163,N_2674,N_3450);
nand U7164 (N_7164,N_3683,N_4850);
nand U7165 (N_7165,N_3285,N_4272);
or U7166 (N_7166,N_4938,N_3847);
and U7167 (N_7167,N_3304,N_3864);
nand U7168 (N_7168,N_4837,N_4191);
and U7169 (N_7169,N_3229,N_2828);
and U7170 (N_7170,N_4388,N_4537);
and U7171 (N_7171,N_3801,N_2621);
or U7172 (N_7172,N_4456,N_3677);
nor U7173 (N_7173,N_3499,N_3211);
nand U7174 (N_7174,N_3815,N_3031);
nor U7175 (N_7175,N_4236,N_4564);
and U7176 (N_7176,N_4385,N_3938);
nor U7177 (N_7177,N_4260,N_3100);
or U7178 (N_7178,N_3027,N_4357);
or U7179 (N_7179,N_3718,N_2678);
and U7180 (N_7180,N_2553,N_4257);
nand U7181 (N_7181,N_3396,N_4490);
or U7182 (N_7182,N_3135,N_3081);
or U7183 (N_7183,N_3995,N_4263);
and U7184 (N_7184,N_3047,N_4559);
or U7185 (N_7185,N_4692,N_3444);
and U7186 (N_7186,N_3724,N_2648);
and U7187 (N_7187,N_2721,N_3733);
nand U7188 (N_7188,N_3546,N_4181);
and U7189 (N_7189,N_4403,N_2590);
nand U7190 (N_7190,N_3984,N_3004);
and U7191 (N_7191,N_4717,N_3249);
nand U7192 (N_7192,N_4349,N_3558);
and U7193 (N_7193,N_4023,N_2658);
or U7194 (N_7194,N_4243,N_3775);
nand U7195 (N_7195,N_3489,N_4646);
and U7196 (N_7196,N_3108,N_2985);
nand U7197 (N_7197,N_3083,N_3137);
and U7198 (N_7198,N_3330,N_2748);
or U7199 (N_7199,N_3011,N_4949);
nand U7200 (N_7200,N_4880,N_4174);
and U7201 (N_7201,N_3253,N_3655);
nand U7202 (N_7202,N_4113,N_3682);
nor U7203 (N_7203,N_4297,N_3827);
and U7204 (N_7204,N_3297,N_3205);
or U7205 (N_7205,N_3833,N_4310);
nand U7206 (N_7206,N_3822,N_4908);
and U7207 (N_7207,N_4586,N_4849);
and U7208 (N_7208,N_3387,N_4490);
and U7209 (N_7209,N_2807,N_4427);
and U7210 (N_7210,N_3126,N_2917);
and U7211 (N_7211,N_3389,N_3970);
or U7212 (N_7212,N_4488,N_2524);
and U7213 (N_7213,N_3543,N_2779);
and U7214 (N_7214,N_4047,N_2949);
nand U7215 (N_7215,N_3030,N_4714);
nor U7216 (N_7216,N_3108,N_2894);
or U7217 (N_7217,N_4883,N_3791);
or U7218 (N_7218,N_4481,N_4031);
or U7219 (N_7219,N_3475,N_3535);
and U7220 (N_7220,N_3982,N_4213);
nor U7221 (N_7221,N_3560,N_2671);
nand U7222 (N_7222,N_3407,N_2502);
and U7223 (N_7223,N_4390,N_3288);
or U7224 (N_7224,N_2966,N_4055);
or U7225 (N_7225,N_3235,N_4463);
and U7226 (N_7226,N_3244,N_3109);
nor U7227 (N_7227,N_4333,N_3348);
nor U7228 (N_7228,N_4390,N_3899);
nand U7229 (N_7229,N_3707,N_3991);
nor U7230 (N_7230,N_4877,N_4646);
nand U7231 (N_7231,N_2590,N_4852);
and U7232 (N_7232,N_3273,N_3371);
nor U7233 (N_7233,N_3104,N_4145);
or U7234 (N_7234,N_2804,N_2991);
nand U7235 (N_7235,N_3090,N_2935);
nor U7236 (N_7236,N_2600,N_4243);
or U7237 (N_7237,N_4283,N_3421);
nor U7238 (N_7238,N_3054,N_4585);
nand U7239 (N_7239,N_3064,N_3038);
nor U7240 (N_7240,N_2850,N_3836);
nor U7241 (N_7241,N_4084,N_3384);
and U7242 (N_7242,N_4280,N_3206);
nor U7243 (N_7243,N_3622,N_3769);
nor U7244 (N_7244,N_3258,N_4418);
or U7245 (N_7245,N_2852,N_3222);
or U7246 (N_7246,N_4904,N_4651);
or U7247 (N_7247,N_4046,N_4252);
nor U7248 (N_7248,N_4607,N_4011);
nand U7249 (N_7249,N_3435,N_2793);
nand U7250 (N_7250,N_4720,N_3204);
and U7251 (N_7251,N_4354,N_3592);
nand U7252 (N_7252,N_4034,N_4358);
nand U7253 (N_7253,N_3064,N_4252);
nand U7254 (N_7254,N_4438,N_4196);
and U7255 (N_7255,N_4077,N_3386);
nand U7256 (N_7256,N_3460,N_3109);
or U7257 (N_7257,N_4238,N_2578);
and U7258 (N_7258,N_3251,N_3580);
or U7259 (N_7259,N_3542,N_2713);
and U7260 (N_7260,N_3264,N_2865);
or U7261 (N_7261,N_3716,N_4372);
nor U7262 (N_7262,N_4478,N_2555);
or U7263 (N_7263,N_2898,N_3156);
and U7264 (N_7264,N_4821,N_4801);
nand U7265 (N_7265,N_2816,N_4518);
nand U7266 (N_7266,N_4004,N_3461);
and U7267 (N_7267,N_3343,N_4878);
nand U7268 (N_7268,N_4645,N_3144);
or U7269 (N_7269,N_4420,N_4329);
nor U7270 (N_7270,N_4130,N_3274);
nand U7271 (N_7271,N_3292,N_2930);
nor U7272 (N_7272,N_2634,N_4611);
nand U7273 (N_7273,N_4567,N_4885);
and U7274 (N_7274,N_3686,N_4016);
nor U7275 (N_7275,N_3123,N_3444);
nor U7276 (N_7276,N_4257,N_4427);
nand U7277 (N_7277,N_4177,N_3882);
xor U7278 (N_7278,N_2551,N_4884);
or U7279 (N_7279,N_3638,N_3233);
nand U7280 (N_7280,N_4510,N_3490);
nor U7281 (N_7281,N_2706,N_4853);
or U7282 (N_7282,N_2950,N_3880);
nand U7283 (N_7283,N_4163,N_4611);
and U7284 (N_7284,N_4462,N_3237);
nor U7285 (N_7285,N_2652,N_3120);
and U7286 (N_7286,N_2941,N_3763);
nand U7287 (N_7287,N_2619,N_3595);
nand U7288 (N_7288,N_4461,N_3056);
and U7289 (N_7289,N_3871,N_3863);
or U7290 (N_7290,N_3422,N_2806);
nor U7291 (N_7291,N_4935,N_3306);
or U7292 (N_7292,N_2538,N_3824);
or U7293 (N_7293,N_3604,N_3878);
xor U7294 (N_7294,N_4766,N_3960);
nor U7295 (N_7295,N_4816,N_4411);
nand U7296 (N_7296,N_4617,N_3497);
or U7297 (N_7297,N_4301,N_2512);
nand U7298 (N_7298,N_4151,N_4777);
or U7299 (N_7299,N_2797,N_2697);
and U7300 (N_7300,N_3818,N_4344);
nor U7301 (N_7301,N_3210,N_3163);
or U7302 (N_7302,N_3971,N_4097);
xnor U7303 (N_7303,N_4666,N_4906);
and U7304 (N_7304,N_2587,N_2605);
or U7305 (N_7305,N_2680,N_3454);
nor U7306 (N_7306,N_4270,N_4916);
nand U7307 (N_7307,N_2740,N_3975);
nand U7308 (N_7308,N_4420,N_4237);
or U7309 (N_7309,N_2970,N_2597);
and U7310 (N_7310,N_3609,N_3271);
or U7311 (N_7311,N_4548,N_4327);
nor U7312 (N_7312,N_4992,N_2712);
or U7313 (N_7313,N_2872,N_4579);
nor U7314 (N_7314,N_4090,N_3713);
nand U7315 (N_7315,N_3491,N_4191);
nor U7316 (N_7316,N_3770,N_4476);
or U7317 (N_7317,N_3807,N_4630);
and U7318 (N_7318,N_4810,N_3856);
nand U7319 (N_7319,N_4318,N_4795);
or U7320 (N_7320,N_3834,N_2733);
nor U7321 (N_7321,N_4621,N_3149);
nand U7322 (N_7322,N_2509,N_3112);
or U7323 (N_7323,N_2931,N_4239);
nand U7324 (N_7324,N_3275,N_2784);
and U7325 (N_7325,N_2878,N_3228);
and U7326 (N_7326,N_4455,N_3294);
nor U7327 (N_7327,N_4623,N_3588);
or U7328 (N_7328,N_3397,N_4507);
nor U7329 (N_7329,N_4268,N_3164);
and U7330 (N_7330,N_4250,N_4585);
nor U7331 (N_7331,N_3133,N_2574);
nand U7332 (N_7332,N_3154,N_3706);
or U7333 (N_7333,N_3012,N_4919);
nor U7334 (N_7334,N_2681,N_4159);
or U7335 (N_7335,N_2770,N_3828);
and U7336 (N_7336,N_4161,N_3795);
or U7337 (N_7337,N_4191,N_3158);
or U7338 (N_7338,N_3795,N_4541);
or U7339 (N_7339,N_3884,N_3171);
nand U7340 (N_7340,N_4693,N_3073);
nand U7341 (N_7341,N_4065,N_4325);
nor U7342 (N_7342,N_3908,N_2762);
nor U7343 (N_7343,N_3132,N_3352);
nor U7344 (N_7344,N_3357,N_2511);
nor U7345 (N_7345,N_4397,N_4351);
or U7346 (N_7346,N_4657,N_4775);
nand U7347 (N_7347,N_2945,N_3329);
nand U7348 (N_7348,N_4836,N_3545);
nand U7349 (N_7349,N_4959,N_4920);
nand U7350 (N_7350,N_2787,N_4184);
or U7351 (N_7351,N_3740,N_4240);
and U7352 (N_7352,N_3975,N_3421);
or U7353 (N_7353,N_4855,N_4175);
and U7354 (N_7354,N_3189,N_2671);
and U7355 (N_7355,N_4203,N_3208);
or U7356 (N_7356,N_3248,N_4727);
and U7357 (N_7357,N_4229,N_4064);
nor U7358 (N_7358,N_3180,N_3850);
nor U7359 (N_7359,N_3184,N_3524);
nand U7360 (N_7360,N_4845,N_3403);
nand U7361 (N_7361,N_4788,N_4337);
and U7362 (N_7362,N_4835,N_3406);
nor U7363 (N_7363,N_4400,N_2647);
and U7364 (N_7364,N_3941,N_3605);
nor U7365 (N_7365,N_2842,N_3342);
nand U7366 (N_7366,N_2622,N_4923);
nand U7367 (N_7367,N_2975,N_2717);
nand U7368 (N_7368,N_3713,N_3579);
and U7369 (N_7369,N_3727,N_4996);
or U7370 (N_7370,N_2595,N_3199);
nor U7371 (N_7371,N_3435,N_3965);
or U7372 (N_7372,N_3466,N_3222);
nor U7373 (N_7373,N_4828,N_4253);
or U7374 (N_7374,N_3036,N_4290);
and U7375 (N_7375,N_4169,N_4125);
and U7376 (N_7376,N_3824,N_4137);
nor U7377 (N_7377,N_2875,N_2948);
nand U7378 (N_7378,N_3775,N_4873);
nor U7379 (N_7379,N_4832,N_4121);
nand U7380 (N_7380,N_3796,N_4111);
nand U7381 (N_7381,N_4877,N_2623);
nand U7382 (N_7382,N_4906,N_3279);
and U7383 (N_7383,N_2509,N_3043);
and U7384 (N_7384,N_3441,N_3263);
nand U7385 (N_7385,N_3147,N_4376);
and U7386 (N_7386,N_2711,N_2543);
nand U7387 (N_7387,N_3945,N_3338);
nand U7388 (N_7388,N_4958,N_3024);
nand U7389 (N_7389,N_3507,N_4939);
and U7390 (N_7390,N_4667,N_3764);
and U7391 (N_7391,N_3057,N_4726);
and U7392 (N_7392,N_4169,N_4579);
and U7393 (N_7393,N_2522,N_3994);
nand U7394 (N_7394,N_3558,N_4782);
nor U7395 (N_7395,N_3085,N_3695);
nor U7396 (N_7396,N_3455,N_3370);
nor U7397 (N_7397,N_3432,N_3662);
and U7398 (N_7398,N_3532,N_2584);
and U7399 (N_7399,N_4487,N_3960);
nand U7400 (N_7400,N_3613,N_3615);
and U7401 (N_7401,N_3716,N_2749);
and U7402 (N_7402,N_4473,N_2544);
and U7403 (N_7403,N_3275,N_3427);
nand U7404 (N_7404,N_2634,N_3196);
nand U7405 (N_7405,N_3664,N_4534);
and U7406 (N_7406,N_3059,N_3100);
and U7407 (N_7407,N_4885,N_2932);
nand U7408 (N_7408,N_2530,N_4150);
and U7409 (N_7409,N_4566,N_4041);
and U7410 (N_7410,N_4390,N_4415);
nor U7411 (N_7411,N_3012,N_3642);
or U7412 (N_7412,N_2836,N_3198);
and U7413 (N_7413,N_2507,N_4505);
nand U7414 (N_7414,N_3036,N_2733);
and U7415 (N_7415,N_2529,N_4928);
and U7416 (N_7416,N_3916,N_2764);
nand U7417 (N_7417,N_3935,N_4933);
or U7418 (N_7418,N_4781,N_3668);
nand U7419 (N_7419,N_3989,N_2721);
nand U7420 (N_7420,N_3878,N_4955);
nand U7421 (N_7421,N_4190,N_4337);
or U7422 (N_7422,N_3757,N_3432);
nor U7423 (N_7423,N_4559,N_3039);
nor U7424 (N_7424,N_4385,N_3976);
nand U7425 (N_7425,N_4436,N_4820);
or U7426 (N_7426,N_4993,N_3656);
nor U7427 (N_7427,N_3841,N_2979);
nor U7428 (N_7428,N_3203,N_3705);
nand U7429 (N_7429,N_3090,N_4479);
nor U7430 (N_7430,N_2977,N_3379);
nor U7431 (N_7431,N_2716,N_2640);
xor U7432 (N_7432,N_4671,N_4469);
and U7433 (N_7433,N_3180,N_2533);
nand U7434 (N_7434,N_3834,N_3418);
and U7435 (N_7435,N_3933,N_4633);
nor U7436 (N_7436,N_3656,N_3021);
and U7437 (N_7437,N_3810,N_4030);
nor U7438 (N_7438,N_3469,N_4751);
or U7439 (N_7439,N_3336,N_4792);
or U7440 (N_7440,N_3401,N_3547);
or U7441 (N_7441,N_4084,N_3670);
nor U7442 (N_7442,N_4859,N_3982);
nor U7443 (N_7443,N_2569,N_4293);
nand U7444 (N_7444,N_2667,N_4594);
nor U7445 (N_7445,N_4155,N_2977);
and U7446 (N_7446,N_3241,N_3030);
and U7447 (N_7447,N_2500,N_2868);
nor U7448 (N_7448,N_2673,N_4528);
xnor U7449 (N_7449,N_3271,N_4513);
nor U7450 (N_7450,N_3636,N_4412);
or U7451 (N_7451,N_2769,N_4855);
and U7452 (N_7452,N_2504,N_4501);
and U7453 (N_7453,N_3416,N_4378);
and U7454 (N_7454,N_3045,N_3699);
and U7455 (N_7455,N_2606,N_2642);
nor U7456 (N_7456,N_2774,N_4843);
and U7457 (N_7457,N_4050,N_3678);
and U7458 (N_7458,N_4463,N_4037);
and U7459 (N_7459,N_4660,N_4706);
nor U7460 (N_7460,N_3181,N_3025);
and U7461 (N_7461,N_4926,N_4270);
or U7462 (N_7462,N_4589,N_3752);
or U7463 (N_7463,N_4617,N_4257);
or U7464 (N_7464,N_4826,N_2747);
or U7465 (N_7465,N_4349,N_2508);
xor U7466 (N_7466,N_3169,N_3115);
nand U7467 (N_7467,N_2759,N_3731);
nor U7468 (N_7468,N_2981,N_3876);
nand U7469 (N_7469,N_4615,N_4570);
and U7470 (N_7470,N_4704,N_4177);
nand U7471 (N_7471,N_3933,N_3294);
nor U7472 (N_7472,N_4179,N_2701);
nor U7473 (N_7473,N_2697,N_2632);
or U7474 (N_7474,N_3282,N_3063);
nor U7475 (N_7475,N_4114,N_2537);
and U7476 (N_7476,N_3927,N_4172);
and U7477 (N_7477,N_2986,N_3364);
nor U7478 (N_7478,N_4865,N_4028);
or U7479 (N_7479,N_3308,N_3832);
nand U7480 (N_7480,N_4319,N_2922);
nor U7481 (N_7481,N_3139,N_4094);
nor U7482 (N_7482,N_3497,N_2577);
or U7483 (N_7483,N_3454,N_4433);
nor U7484 (N_7484,N_3305,N_3464);
xnor U7485 (N_7485,N_3385,N_3063);
nor U7486 (N_7486,N_3548,N_4218);
nand U7487 (N_7487,N_4766,N_3527);
nand U7488 (N_7488,N_3953,N_3692);
or U7489 (N_7489,N_4664,N_3840);
and U7490 (N_7490,N_4249,N_3466);
nand U7491 (N_7491,N_4540,N_3023);
nor U7492 (N_7492,N_4762,N_4977);
nand U7493 (N_7493,N_3024,N_4891);
nor U7494 (N_7494,N_4768,N_2902);
nor U7495 (N_7495,N_3554,N_2617);
nor U7496 (N_7496,N_4170,N_2669);
nand U7497 (N_7497,N_2856,N_3972);
nor U7498 (N_7498,N_2758,N_4662);
nor U7499 (N_7499,N_4256,N_3483);
or U7500 (N_7500,N_5679,N_5562);
xnor U7501 (N_7501,N_5678,N_7217);
or U7502 (N_7502,N_5600,N_7362);
nand U7503 (N_7503,N_6980,N_7113);
or U7504 (N_7504,N_7162,N_5023);
and U7505 (N_7505,N_7059,N_5959);
or U7506 (N_7506,N_6407,N_7248);
and U7507 (N_7507,N_6520,N_5418);
and U7508 (N_7508,N_5828,N_5355);
xnor U7509 (N_7509,N_5712,N_5097);
or U7510 (N_7510,N_5033,N_5560);
and U7511 (N_7511,N_6059,N_5024);
and U7512 (N_7512,N_6434,N_5886);
and U7513 (N_7513,N_6217,N_5128);
nor U7514 (N_7514,N_7137,N_6202);
nand U7515 (N_7515,N_6421,N_7377);
nand U7516 (N_7516,N_6963,N_6997);
and U7517 (N_7517,N_7039,N_6351);
nand U7518 (N_7518,N_6218,N_6086);
nand U7519 (N_7519,N_6853,N_6797);
nand U7520 (N_7520,N_7483,N_5360);
nand U7521 (N_7521,N_6388,N_6064);
nand U7522 (N_7522,N_6163,N_5518);
or U7523 (N_7523,N_5867,N_5935);
nor U7524 (N_7524,N_6174,N_6899);
nand U7525 (N_7525,N_7041,N_6277);
or U7526 (N_7526,N_6114,N_6026);
nand U7527 (N_7527,N_5158,N_5747);
or U7528 (N_7528,N_6286,N_6385);
nor U7529 (N_7529,N_6964,N_7357);
and U7530 (N_7530,N_5055,N_6832);
and U7531 (N_7531,N_5166,N_5126);
and U7532 (N_7532,N_6012,N_6358);
nor U7533 (N_7533,N_7388,N_6786);
nand U7534 (N_7534,N_5784,N_5841);
or U7535 (N_7535,N_6413,N_5339);
nor U7536 (N_7536,N_5569,N_7364);
nor U7537 (N_7537,N_7087,N_5929);
nand U7538 (N_7538,N_6606,N_5022);
or U7539 (N_7539,N_5471,N_6659);
nand U7540 (N_7540,N_5016,N_6770);
and U7541 (N_7541,N_5373,N_6763);
nand U7542 (N_7542,N_6562,N_5982);
nand U7543 (N_7543,N_7212,N_5907);
and U7544 (N_7544,N_6144,N_6554);
nor U7545 (N_7545,N_6664,N_5842);
nor U7546 (N_7546,N_6690,N_6519);
nor U7547 (N_7547,N_5881,N_7480);
or U7548 (N_7548,N_7214,N_6037);
or U7549 (N_7549,N_5082,N_5833);
nor U7550 (N_7550,N_5541,N_5150);
nand U7551 (N_7551,N_6005,N_5141);
or U7552 (N_7552,N_6641,N_6447);
and U7553 (N_7553,N_5244,N_5405);
and U7554 (N_7554,N_6563,N_5762);
or U7555 (N_7555,N_5919,N_5465);
nor U7556 (N_7556,N_5791,N_6632);
or U7557 (N_7557,N_5401,N_5845);
or U7558 (N_7558,N_5273,N_6992);
and U7559 (N_7559,N_6045,N_5334);
nor U7560 (N_7560,N_6576,N_6183);
and U7561 (N_7561,N_6881,N_6192);
nand U7562 (N_7562,N_6120,N_5351);
nor U7563 (N_7563,N_5636,N_5194);
or U7564 (N_7564,N_7126,N_6707);
and U7565 (N_7565,N_5298,N_7481);
or U7566 (N_7566,N_7308,N_7276);
nand U7567 (N_7567,N_5192,N_7218);
and U7568 (N_7568,N_6715,N_5756);
nor U7569 (N_7569,N_6834,N_5065);
and U7570 (N_7570,N_6542,N_6527);
nor U7571 (N_7571,N_6041,N_5502);
and U7572 (N_7572,N_5299,N_6986);
nand U7573 (N_7573,N_5080,N_5875);
nor U7574 (N_7574,N_5611,N_7210);
nand U7575 (N_7575,N_6231,N_5314);
nor U7576 (N_7576,N_6541,N_5794);
and U7577 (N_7577,N_5731,N_5153);
and U7578 (N_7578,N_6851,N_5409);
nor U7579 (N_7579,N_7190,N_5889);
and U7580 (N_7580,N_5795,N_6315);
nand U7581 (N_7581,N_6386,N_5849);
or U7582 (N_7582,N_5127,N_7426);
nand U7583 (N_7583,N_6210,N_6160);
nor U7584 (N_7584,N_5102,N_6206);
nand U7585 (N_7585,N_6904,N_6816);
nor U7586 (N_7586,N_6106,N_5478);
or U7587 (N_7587,N_5764,N_6538);
nor U7588 (N_7588,N_5744,N_5480);
nor U7589 (N_7589,N_5948,N_6984);
nand U7590 (N_7590,N_7149,N_6034);
or U7591 (N_7591,N_6586,N_6995);
nor U7592 (N_7592,N_6536,N_5695);
nand U7593 (N_7593,N_7492,N_5258);
nor U7594 (N_7594,N_6234,N_5680);
nor U7595 (N_7595,N_7375,N_7057);
nand U7596 (N_7596,N_6165,N_6254);
nand U7597 (N_7597,N_5508,N_5301);
or U7598 (N_7598,N_5533,N_6304);
or U7599 (N_7599,N_6172,N_6877);
nand U7600 (N_7600,N_5343,N_5709);
and U7601 (N_7601,N_5321,N_6621);
or U7602 (N_7602,N_6622,N_6485);
and U7603 (N_7603,N_6173,N_6177);
nor U7604 (N_7604,N_5821,N_6883);
or U7605 (N_7605,N_6199,N_7222);
nor U7606 (N_7606,N_5608,N_5383);
nand U7607 (N_7607,N_6938,N_6249);
and U7608 (N_7608,N_5655,N_5340);
or U7609 (N_7609,N_5977,N_6808);
or U7610 (N_7610,N_5835,N_7200);
nor U7611 (N_7611,N_5345,N_6750);
nor U7612 (N_7612,N_5958,N_5840);
and U7613 (N_7613,N_7437,N_6467);
nor U7614 (N_7614,N_6945,N_5199);
or U7615 (N_7615,N_5838,N_6241);
or U7616 (N_7616,N_6500,N_5701);
nor U7617 (N_7617,N_7441,N_7233);
and U7618 (N_7618,N_6108,N_7453);
or U7619 (N_7619,N_5281,N_5399);
and U7620 (N_7620,N_5124,N_5090);
nor U7621 (N_7621,N_7229,N_6435);
and U7622 (N_7622,N_7431,N_5063);
nand U7623 (N_7623,N_5937,N_6164);
nand U7624 (N_7624,N_6783,N_7455);
and U7625 (N_7625,N_5243,N_5939);
nor U7626 (N_7626,N_6533,N_6637);
and U7627 (N_7627,N_7472,N_5610);
nor U7628 (N_7628,N_6625,N_5514);
nand U7629 (N_7629,N_6593,N_6999);
and U7630 (N_7630,N_5598,N_6932);
and U7631 (N_7631,N_7077,N_6374);
and U7632 (N_7632,N_6159,N_7345);
and U7633 (N_7633,N_5564,N_5619);
or U7634 (N_7634,N_7342,N_7312);
and U7635 (N_7635,N_5002,N_6560);
nor U7636 (N_7636,N_6867,N_6776);
nor U7637 (N_7637,N_5675,N_6968);
and U7638 (N_7638,N_5285,N_7489);
or U7639 (N_7639,N_6511,N_7167);
or U7640 (N_7640,N_5966,N_5164);
nand U7641 (N_7641,N_6640,N_5924);
and U7642 (N_7642,N_6966,N_7242);
or U7643 (N_7643,N_6890,N_7280);
and U7644 (N_7644,N_5513,N_7287);
and U7645 (N_7645,N_7022,N_6870);
nor U7646 (N_7646,N_7114,N_7000);
and U7647 (N_7647,N_6534,N_5808);
nand U7648 (N_7648,N_7407,N_6901);
and U7649 (N_7649,N_5705,N_5653);
nor U7650 (N_7650,N_7452,N_7465);
nor U7651 (N_7651,N_7095,N_5635);
and U7652 (N_7652,N_5499,N_6452);
nor U7653 (N_7653,N_5358,N_5210);
nor U7654 (N_7654,N_5446,N_6155);
nand U7655 (N_7655,N_5894,N_5910);
nor U7656 (N_7656,N_5738,N_7320);
nand U7657 (N_7657,N_5839,N_6491);
nand U7658 (N_7658,N_6761,N_6322);
nand U7659 (N_7659,N_7098,N_6395);
nand U7660 (N_7660,N_5672,N_5238);
nor U7661 (N_7661,N_6729,N_6962);
nand U7662 (N_7662,N_5879,N_7406);
or U7663 (N_7663,N_6913,N_5818);
nor U7664 (N_7664,N_6660,N_5187);
nor U7665 (N_7665,N_5404,N_5230);
or U7666 (N_7666,N_6893,N_5615);
and U7667 (N_7667,N_5017,N_5219);
nand U7668 (N_7668,N_5282,N_6492);
or U7669 (N_7669,N_6055,N_6833);
nand U7670 (N_7670,N_6117,N_6926);
nand U7671 (N_7671,N_6198,N_5092);
nor U7672 (N_7672,N_5753,N_7050);
or U7673 (N_7673,N_6824,N_7428);
and U7674 (N_7674,N_6830,N_6800);
or U7675 (N_7675,N_6376,N_5522);
nand U7676 (N_7676,N_5944,N_7111);
nor U7677 (N_7677,N_5980,N_5684);
or U7678 (N_7678,N_6673,N_7354);
and U7679 (N_7679,N_7230,N_5294);
nor U7680 (N_7680,N_6835,N_6071);
nand U7681 (N_7681,N_5946,N_5938);
and U7682 (N_7682,N_6720,N_6047);
and U7683 (N_7683,N_6810,N_6356);
or U7684 (N_7684,N_6123,N_7238);
and U7685 (N_7685,N_5912,N_7378);
nand U7686 (N_7686,N_6112,N_6687);
nand U7687 (N_7687,N_5084,N_5716);
or U7688 (N_7688,N_5323,N_5302);
or U7689 (N_7689,N_5999,N_6317);
and U7690 (N_7690,N_6787,N_6662);
or U7691 (N_7691,N_6567,N_6344);
nand U7692 (N_7692,N_6179,N_6171);
or U7693 (N_7693,N_6359,N_6517);
nand U7694 (N_7694,N_6128,N_5226);
nand U7695 (N_7695,N_6521,N_6205);
nor U7696 (N_7696,N_6247,N_6608);
nand U7697 (N_7697,N_6424,N_7156);
nand U7698 (N_7698,N_6397,N_5379);
and U7699 (N_7699,N_7062,N_5066);
or U7700 (N_7700,N_6296,N_6748);
nand U7701 (N_7701,N_5832,N_5677);
nor U7702 (N_7702,N_7414,N_6175);
nor U7703 (N_7703,N_5783,N_5754);
and U7704 (N_7704,N_6765,N_6955);
nand U7705 (N_7705,N_6250,N_6242);
and U7706 (N_7706,N_5468,N_6595);
or U7707 (N_7707,N_6915,N_5030);
nor U7708 (N_7708,N_6185,N_5311);
and U7709 (N_7709,N_6818,N_6384);
nand U7710 (N_7710,N_5687,N_7495);
nand U7711 (N_7711,N_5654,N_6569);
nor U7712 (N_7712,N_5272,N_5426);
nor U7713 (N_7713,N_6178,N_6590);
nor U7714 (N_7714,N_5917,N_5139);
nand U7715 (N_7715,N_6746,N_5739);
or U7716 (N_7716,N_7031,N_6594);
or U7717 (N_7717,N_6767,N_5632);
nand U7718 (N_7718,N_6456,N_7145);
nor U7719 (N_7719,N_5457,N_6483);
nand U7720 (N_7720,N_6880,N_6489);
or U7721 (N_7721,N_6739,N_5553);
nand U7722 (N_7722,N_5018,N_5700);
nor U7723 (N_7723,N_6345,N_5901);
or U7724 (N_7724,N_5666,N_6579);
nor U7725 (N_7725,N_6826,N_6737);
xor U7726 (N_7726,N_7189,N_6000);
and U7727 (N_7727,N_7464,N_5807);
nor U7728 (N_7728,N_6961,N_6067);
nand U7729 (N_7729,N_6855,N_6602);
or U7730 (N_7730,N_6793,N_5361);
nand U7731 (N_7731,N_6781,N_5740);
and U7732 (N_7732,N_5231,N_5526);
and U7733 (N_7733,N_6098,N_6268);
nand U7734 (N_7734,N_5202,N_6136);
and U7735 (N_7735,N_6119,N_7366);
nor U7736 (N_7736,N_6546,N_5941);
and U7737 (N_7737,N_6142,N_6036);
xor U7738 (N_7738,N_6558,N_6646);
nor U7739 (N_7739,N_5888,N_7326);
nand U7740 (N_7740,N_6667,N_5147);
nor U7741 (N_7741,N_7344,N_5543);
nor U7742 (N_7742,N_7123,N_7301);
or U7743 (N_7743,N_5736,N_5656);
nor U7744 (N_7744,N_6592,N_6382);
nor U7745 (N_7745,N_7392,N_5032);
nand U7746 (N_7746,N_5184,N_5670);
nor U7747 (N_7747,N_5035,N_7102);
nor U7748 (N_7748,N_5289,N_6956);
nand U7749 (N_7749,N_5162,N_5115);
and U7750 (N_7750,N_5581,N_5971);
and U7751 (N_7751,N_6878,N_5782);
nor U7752 (N_7752,N_5330,N_6862);
nand U7753 (N_7753,N_5693,N_7278);
nand U7754 (N_7754,N_7066,N_5934);
nor U7755 (N_7755,N_6292,N_5490);
nand U7756 (N_7756,N_5384,N_5182);
and U7757 (N_7757,N_6158,N_5211);
and U7758 (N_7758,N_6285,N_6188);
nand U7759 (N_7759,N_7139,N_6768);
xor U7760 (N_7760,N_7467,N_7361);
and U7761 (N_7761,N_6400,N_5037);
and U7762 (N_7762,N_6011,N_6203);
or U7763 (N_7763,N_6008,N_6967);
nand U7764 (N_7764,N_5039,N_6223);
nor U7765 (N_7765,N_5583,N_5786);
or U7766 (N_7766,N_5613,N_5352);
or U7767 (N_7767,N_7018,N_6204);
nor U7768 (N_7768,N_6807,N_7376);
and U7769 (N_7769,N_6013,N_5930);
and U7770 (N_7770,N_6745,N_7420);
or U7771 (N_7771,N_6742,N_6639);
nand U7772 (N_7772,N_5427,N_5824);
nand U7773 (N_7773,N_6912,N_7255);
nand U7774 (N_7774,N_5453,N_5223);
nand U7775 (N_7775,N_6327,N_6137);
or U7776 (N_7776,N_5998,N_7448);
or U7777 (N_7777,N_7067,N_5987);
or U7778 (N_7778,N_6216,N_5572);
nor U7779 (N_7779,N_6419,N_6338);
nand U7780 (N_7780,N_5500,N_7380);
nor U7781 (N_7781,N_7083,N_7013);
nand U7782 (N_7782,N_7252,N_7429);
and U7783 (N_7783,N_6732,N_5725);
nand U7784 (N_7784,N_5758,N_6676);
and U7785 (N_7785,N_5617,N_6403);
or U7786 (N_7786,N_5530,N_6050);
nor U7787 (N_7787,N_5057,N_5891);
and U7788 (N_7788,N_5317,N_5266);
or U7789 (N_7789,N_5129,N_7314);
nand U7790 (N_7790,N_7418,N_6460);
and U7791 (N_7791,N_6256,N_7140);
nand U7792 (N_7792,N_6649,N_5606);
nor U7793 (N_7793,N_7239,N_6815);
and U7794 (N_7794,N_5232,N_6596);
nand U7795 (N_7795,N_6156,N_7129);
and U7796 (N_7796,N_7413,N_5324);
and U7797 (N_7797,N_7417,N_5646);
or U7798 (N_7798,N_5131,N_5096);
nor U7799 (N_7799,N_7215,N_6484);
or U7800 (N_7800,N_6110,N_7141);
nand U7801 (N_7801,N_5292,N_6414);
nand U7802 (N_7802,N_7109,N_5048);
and U7803 (N_7803,N_5699,N_6430);
or U7804 (N_7804,N_7091,N_6230);
nand U7805 (N_7805,N_6196,N_5088);
nor U7806 (N_7806,N_6614,N_7183);
nor U7807 (N_7807,N_5704,N_5138);
and U7808 (N_7808,N_7168,N_6598);
nand U7809 (N_7809,N_5075,N_5819);
and U7810 (N_7810,N_6528,N_5239);
nand U7811 (N_7811,N_6105,N_6604);
nand U7812 (N_7812,N_6154,N_6948);
nor U7813 (N_7813,N_6982,N_6871);
nor U7814 (N_7814,N_6147,N_6891);
and U7815 (N_7815,N_7164,N_6708);
nor U7816 (N_7816,N_5013,N_6033);
or U7817 (N_7817,N_6021,N_5437);
nand U7818 (N_7818,N_7463,N_5058);
and U7819 (N_7819,N_6918,N_5026);
or U7820 (N_7820,N_5227,N_5969);
and U7821 (N_7821,N_6258,N_7339);
nor U7822 (N_7822,N_6073,N_6752);
and U7823 (N_7823,N_6087,N_5641);
nand U7824 (N_7824,N_6193,N_6700);
nand U7825 (N_7825,N_5949,N_6079);
and U7826 (N_7826,N_7135,N_5902);
or U7827 (N_7827,N_7277,N_5940);
nand U7828 (N_7828,N_5261,N_7147);
or U7829 (N_7829,N_5588,N_5325);
or U7830 (N_7830,N_6896,N_7082);
or U7831 (N_7831,N_5594,N_7103);
nor U7832 (N_7832,N_5054,N_5719);
nand U7833 (N_7833,N_6184,N_5010);
or U7834 (N_7834,N_7370,N_5196);
or U7835 (N_7835,N_5111,N_6780);
nor U7836 (N_7836,N_6642,N_7004);
and U7837 (N_7837,N_6548,N_6812);
nor U7838 (N_7838,N_7052,N_6052);
and U7839 (N_7839,N_6979,N_5309);
nor U7840 (N_7840,N_6272,N_5714);
and U7841 (N_7841,N_6279,N_5750);
or U7842 (N_7842,N_5884,N_6138);
nor U7843 (N_7843,N_7254,N_6333);
or U7844 (N_7844,N_5485,N_6378);
and U7845 (N_7845,N_6189,N_5393);
nand U7846 (N_7846,N_5883,N_6283);
nand U7847 (N_7847,N_5348,N_6907);
nand U7848 (N_7848,N_6126,N_5920);
nand U7849 (N_7849,N_6131,N_7471);
and U7850 (N_7850,N_6436,N_5876);
nor U7851 (N_7851,N_6450,N_7038);
nand U7852 (N_7852,N_6772,N_7346);
or U7853 (N_7853,N_6619,N_6991);
nor U7854 (N_7854,N_6577,N_5354);
nand U7855 (N_7855,N_5246,N_6349);
and U7856 (N_7856,N_5118,N_7115);
and U7857 (N_7857,N_5320,N_5439);
and U7858 (N_7858,N_6473,N_5060);
nor U7859 (N_7859,N_5040,N_5277);
xor U7860 (N_7860,N_5625,N_6451);
or U7861 (N_7861,N_6207,N_6253);
nor U7862 (N_7862,N_7462,N_7488);
nor U7863 (N_7863,N_6457,N_6028);
nand U7864 (N_7864,N_5943,N_5378);
nor U7865 (N_7865,N_7296,N_5205);
and U7866 (N_7866,N_6943,N_5767);
and U7867 (N_7867,N_6262,N_5178);
nand U7868 (N_7868,N_6412,N_5052);
nand U7869 (N_7869,N_6898,N_6774);
and U7870 (N_7870,N_5322,N_6464);
xor U7871 (N_7871,N_6100,N_6820);
nand U7872 (N_7872,N_6522,N_5603);
or U7873 (N_7873,N_5132,N_5217);
nand U7874 (N_7874,N_5270,N_6080);
and U7875 (N_7875,N_5267,N_7390);
nor U7876 (N_7876,N_6251,N_5357);
nand U7877 (N_7877,N_5776,N_5724);
and U7878 (N_7878,N_5640,N_7011);
and U7879 (N_7879,N_5637,N_6391);
and U7880 (N_7880,N_7244,N_6042);
or U7881 (N_7881,N_5950,N_5715);
nand U7882 (N_7882,N_6805,N_6214);
or U7883 (N_7883,N_5955,N_5604);
nand U7884 (N_7884,N_5781,N_7369);
nand U7885 (N_7885,N_5592,N_6257);
and U7886 (N_7886,N_6738,N_7476);
nor U7887 (N_7887,N_5326,N_6297);
nand U7888 (N_7888,N_6307,N_6718);
nand U7889 (N_7889,N_5547,N_6273);
nand U7890 (N_7890,N_6631,N_5095);
nand U7891 (N_7891,N_5371,N_6053);
and U7892 (N_7892,N_5593,N_5444);
and U7893 (N_7893,N_5804,N_5722);
or U7894 (N_7894,N_6377,N_5899);
nor U7895 (N_7895,N_5253,N_5411);
nor U7896 (N_7896,N_5336,N_7384);
or U7897 (N_7897,N_7024,N_7397);
nand U7898 (N_7898,N_6298,N_5046);
nor U7899 (N_7899,N_5788,N_7173);
or U7900 (N_7900,N_5820,N_5488);
nand U7901 (N_7901,N_5616,N_5119);
or U7902 (N_7902,N_7386,N_5844);
nand U7903 (N_7903,N_7268,N_5774);
nand U7904 (N_7904,N_6446,N_6440);
and U7905 (N_7905,N_5951,N_6766);
or U7906 (N_7906,N_5586,N_5053);
nor U7907 (N_7907,N_6837,N_7374);
nand U7908 (N_7908,N_6624,N_6083);
nand U7909 (N_7909,N_7184,N_5104);
or U7910 (N_7910,N_6396,N_6725);
and U7911 (N_7911,N_6044,N_6906);
and U7912 (N_7912,N_6782,N_7090);
and U7913 (N_7913,N_6726,N_6404);
nand U7914 (N_7914,N_6681,N_7125);
or U7915 (N_7915,N_6688,N_5374);
or U7916 (N_7916,N_6628,N_5109);
nand U7917 (N_7917,N_6654,N_5407);
or U7918 (N_7918,N_6167,N_5531);
or U7919 (N_7919,N_5525,N_5051);
nor U7920 (N_7920,N_7457,N_6872);
and U7921 (N_7921,N_5293,N_6441);
nor U7922 (N_7922,N_5609,N_6854);
or U7923 (N_7923,N_6024,N_7089);
or U7924 (N_7924,N_5093,N_6613);
or U7925 (N_7925,N_5516,N_7026);
or U7926 (N_7926,N_5529,N_6466);
nor U7927 (N_7927,N_5003,N_7043);
nand U7928 (N_7928,N_6074,N_7385);
nand U7929 (N_7929,N_5275,N_5861);
and U7930 (N_7930,N_6553,N_5450);
nor U7931 (N_7931,N_6462,N_5652);
nand U7932 (N_7932,N_6838,N_6882);
or U7933 (N_7933,N_7267,N_7450);
or U7934 (N_7934,N_6672,N_7466);
and U7935 (N_7935,N_6109,N_5208);
and U7936 (N_7936,N_6523,N_6507);
nor U7937 (N_7937,N_7061,N_5662);
or U7938 (N_7938,N_6305,N_6107);
and U7939 (N_7939,N_5155,N_6121);
nor U7940 (N_7940,N_5857,N_5831);
nor U7941 (N_7941,N_6705,N_5172);
nor U7942 (N_7942,N_6438,N_5491);
nor U7943 (N_7943,N_7181,N_5300);
and U7944 (N_7944,N_5268,N_6796);
and U7945 (N_7945,N_5858,N_6601);
and U7946 (N_7946,N_7042,N_5785);
or U7947 (N_7947,N_7270,N_6002);
and U7948 (N_7948,N_5436,N_6844);
and U7949 (N_7949,N_5766,N_5658);
and U7950 (N_7950,N_5843,N_6879);
nor U7951 (N_7951,N_5318,N_7211);
nand U7952 (N_7952,N_6375,N_7161);
nor U7953 (N_7953,N_7275,N_5790);
or U7954 (N_7954,N_7063,N_5906);
nor U7955 (N_7955,N_5872,N_5771);
nor U7956 (N_7956,N_6515,N_7227);
xor U7957 (N_7957,N_6971,N_6030);
and U7958 (N_7958,N_6010,N_6994);
and U7959 (N_7959,N_6468,N_7092);
or U7960 (N_7960,N_5346,N_6860);
nand U7961 (N_7961,N_6009,N_6482);
or U7962 (N_7962,N_6146,N_5618);
nor U7963 (N_7963,N_7319,N_5100);
nor U7964 (N_7964,N_6727,N_6617);
and U7965 (N_7965,N_7408,N_7148);
and U7966 (N_7966,N_6070,N_6627);
or U7967 (N_7967,N_6609,N_5419);
nor U7968 (N_7968,N_7228,N_6828);
and U7969 (N_7969,N_5686,N_6319);
nand U7970 (N_7970,N_7056,N_6556);
nor U7971 (N_7971,N_6827,N_6209);
nor U7972 (N_7972,N_7434,N_6916);
or U7973 (N_7973,N_5925,N_5333);
and U7974 (N_7974,N_5769,N_5799);
nor U7975 (N_7975,N_6266,N_5041);
nand U7976 (N_7976,N_6381,N_6111);
xor U7977 (N_7977,N_7309,N_5422);
or U7978 (N_7978,N_5535,N_6389);
nor U7979 (N_7979,N_7444,N_5554);
and U7980 (N_7980,N_5923,N_6734);
or U7981 (N_7981,N_7197,N_6347);
nand U7982 (N_7982,N_5537,N_6884);
or U7983 (N_7983,N_7101,N_6993);
or U7984 (N_7984,N_7298,N_6288);
or U7985 (N_7985,N_7100,N_6263);
or U7986 (N_7986,N_5911,N_6928);
and U7987 (N_7987,N_5143,N_7093);
or U7988 (N_7988,N_5663,N_5170);
or U7989 (N_7989,N_7006,N_6565);
nand U7990 (N_7990,N_6859,N_7220);
nor U7991 (N_7991,N_5551,N_7293);
and U7992 (N_7992,N_5792,N_6866);
or U7993 (N_7993,N_5430,N_5620);
nor U7994 (N_7994,N_7247,N_5628);
or U7995 (N_7995,N_7338,N_5174);
or U7996 (N_7996,N_6362,N_5234);
nor U7997 (N_7997,N_7021,N_6588);
or U7998 (N_7998,N_5027,N_7236);
nand U7999 (N_7999,N_6847,N_7080);
nor U8000 (N_8000,N_6721,N_6633);
and U8001 (N_8001,N_7106,N_5347);
or U8002 (N_8002,N_5218,N_5315);
and U8003 (N_8003,N_6201,N_6023);
xor U8004 (N_8004,N_6863,N_5681);
nor U8005 (N_8005,N_5846,N_5733);
nor U8006 (N_8006,N_5524,N_6244);
and U8007 (N_8007,N_6150,N_7016);
nor U8008 (N_8008,N_6427,N_5389);
or U8009 (N_8009,N_6448,N_7235);
nand U8010 (N_8010,N_6326,N_6924);
nor U8011 (N_8011,N_6299,N_6379);
or U8012 (N_8012,N_5248,N_6061);
nand U8013 (N_8013,N_5896,N_6324);
or U8014 (N_8014,N_7195,N_6743);
and U8015 (N_8015,N_6399,N_6494);
nor U8016 (N_8016,N_6089,N_5428);
nand U8017 (N_8017,N_7482,N_5802);
nor U8018 (N_8018,N_5986,N_7353);
and U8019 (N_8019,N_7435,N_5176);
nand U8020 (N_8020,N_7142,N_7279);
nor U8021 (N_8021,N_6846,N_5648);
and U8022 (N_8022,N_6006,N_5319);
and U8023 (N_8023,N_6246,N_5449);
and U8024 (N_8024,N_7349,N_5429);
or U8025 (N_8025,N_5121,N_5448);
nand U8026 (N_8026,N_6689,N_6278);
nand U8027 (N_8027,N_5413,N_6040);
nor U8028 (N_8028,N_6211,N_6751);
and U8029 (N_8029,N_6488,N_7330);
nand U8030 (N_8030,N_6845,N_6227);
or U8031 (N_8031,N_7201,N_5214);
or U8032 (N_8032,N_5312,N_7474);
and U8033 (N_8033,N_6157,N_6383);
or U8034 (N_8034,N_5869,N_5112);
or U8035 (N_8035,N_6368,N_7485);
nand U8036 (N_8036,N_5649,N_7216);
nand U8037 (N_8037,N_6289,N_5789);
and U8038 (N_8038,N_6417,N_6169);
or U8039 (N_8039,N_6096,N_5956);
or U8040 (N_8040,N_5942,N_6771);
nor U8041 (N_8041,N_7323,N_6795);
nand U8042 (N_8042,N_5854,N_6303);
or U8043 (N_8043,N_7405,N_6367);
xor U8044 (N_8044,N_6550,N_6501);
nand U8045 (N_8045,N_5650,N_6996);
nor U8046 (N_8046,N_6019,N_5735);
and U8047 (N_8047,N_5059,N_6764);
or U8048 (N_8048,N_6583,N_6530);
nand U8049 (N_8049,N_6735,N_5689);
or U8050 (N_8050,N_6537,N_6741);
or U8051 (N_8051,N_6927,N_5101);
and U8052 (N_8052,N_6544,N_6566);
nor U8053 (N_8053,N_7005,N_5953);
nand U8054 (N_8054,N_5414,N_7134);
nand U8055 (N_8055,N_5988,N_6187);
or U8056 (N_8056,N_6293,N_6392);
nand U8057 (N_8057,N_5287,N_5555);
nand U8058 (N_8058,N_5741,N_5577);
and U8059 (N_8059,N_6573,N_6671);
nand U8060 (N_8060,N_5149,N_5534);
nand U8061 (N_8061,N_7447,N_6698);
nand U8062 (N_8062,N_5501,N_6480);
nand U8063 (N_8063,N_6954,N_6804);
or U8064 (N_8064,N_5812,N_5660);
and U8065 (N_8065,N_6161,N_6477);
and U8066 (N_8066,N_6524,N_5417);
nand U8067 (N_8067,N_7411,N_7107);
and U8068 (N_8068,N_6271,N_5931);
and U8069 (N_8069,N_6133,N_5262);
or U8070 (N_8070,N_6166,N_5370);
or U8071 (N_8071,N_6364,N_6406);
nor U8072 (N_8072,N_7079,N_5344);
and U8073 (N_8073,N_5201,N_6775);
and U8074 (N_8074,N_5497,N_7243);
or U8075 (N_8075,N_6295,N_6437);
nor U8076 (N_8076,N_7198,N_6060);
nand U8077 (N_8077,N_5580,N_7153);
and U8078 (N_8078,N_7415,N_7170);
nand U8079 (N_8079,N_5834,N_7014);
xnor U8080 (N_8080,N_5203,N_6151);
nor U8081 (N_8081,N_7251,N_5175);
xnor U8082 (N_8082,N_5241,N_6235);
or U8083 (N_8083,N_6723,N_5589);
nand U8084 (N_8084,N_5042,N_7105);
or U8085 (N_8085,N_5866,N_6340);
nand U8086 (N_8086,N_5797,N_5265);
nand U8087 (N_8087,N_6426,N_5154);
nor U8088 (N_8088,N_7117,N_6069);
or U8089 (N_8089,N_5880,N_7347);
or U8090 (N_8090,N_6529,N_7324);
and U8091 (N_8091,N_7012,N_5623);
nor U8092 (N_8092,N_6029,N_5970);
or U8093 (N_8093,N_7340,N_7421);
nor U8094 (N_8094,N_7305,N_5064);
and U8095 (N_8095,N_5163,N_5512);
or U8096 (N_8096,N_5932,N_5895);
and U8097 (N_8097,N_5009,N_6703);
or U8098 (N_8098,N_6587,N_5968);
or U8099 (N_8099,N_7128,N_7350);
and U8100 (N_8100,N_5160,N_6267);
nand U8101 (N_8101,N_5091,N_6497);
or U8102 (N_8102,N_7023,N_6091);
or U8103 (N_8103,N_6420,N_6090);
and U8104 (N_8104,N_7300,N_5721);
nand U8105 (N_8105,N_6197,N_7071);
or U8106 (N_8106,N_6471,N_7193);
nor U8107 (N_8107,N_6243,N_6001);
or U8108 (N_8108,N_5447,N_7295);
nand U8109 (N_8109,N_6652,N_6035);
nor U8110 (N_8110,N_6942,N_5976);
nor U8111 (N_8111,N_5368,N_6094);
and U8112 (N_8112,N_5992,N_6894);
and U8113 (N_8113,N_7253,N_7172);
nand U8114 (N_8114,N_6219,N_6868);
and U8115 (N_8115,N_6516,N_7076);
or U8116 (N_8116,N_6095,N_5366);
and U8117 (N_8117,N_6714,N_6819);
nor U8118 (N_8118,N_7202,N_7015);
or U8119 (N_8119,N_5410,N_5183);
and U8120 (N_8120,N_6481,N_6978);
nor U8121 (N_8121,N_5233,N_5979);
and U8122 (N_8122,N_6848,N_6153);
and U8123 (N_8123,N_7150,N_6331);
xnor U8124 (N_8124,N_7240,N_5078);
and U8125 (N_8125,N_6897,N_7290);
nor U8126 (N_8126,N_7379,N_5469);
or U8127 (N_8127,N_5916,N_6811);
nand U8128 (N_8128,N_5952,N_5487);
nand U8129 (N_8129,N_6004,N_6320);
and U8130 (N_8130,N_7175,N_5983);
nand U8131 (N_8131,N_5106,N_7269);
or U8132 (N_8132,N_6465,N_7332);
and U8133 (N_8133,N_5596,N_6401);
nor U8134 (N_8134,N_6355,N_5981);
or U8135 (N_8135,N_6335,N_7281);
or U8136 (N_8136,N_6754,N_6518);
or U8137 (N_8137,N_5926,N_5255);
nand U8138 (N_8138,N_5467,N_7365);
nor U8139 (N_8139,N_5161,N_6168);
nor U8140 (N_8140,N_6616,N_5591);
nor U8141 (N_8141,N_5280,N_7316);
or U8142 (N_8142,N_5552,N_6309);
nand U8143 (N_8143,N_5136,N_5728);
and U8144 (N_8144,N_6139,N_5836);
or U8145 (N_8145,N_6603,N_6970);
and U8146 (N_8146,N_7163,N_7283);
nand U8147 (N_8147,N_6665,N_6498);
nand U8148 (N_8148,N_6017,N_6803);
and U8149 (N_8149,N_5290,N_5156);
or U8150 (N_8150,N_6935,N_5067);
nand U8151 (N_8151,N_7325,N_7249);
nand U8152 (N_8152,N_6929,N_5729);
or U8153 (N_8153,N_7321,N_6762);
nor U8154 (N_8154,N_6459,N_5375);
nand U8155 (N_8155,N_7404,N_6865);
nor U8156 (N_8156,N_6103,N_6618);
nor U8157 (N_8157,N_5228,N_5308);
nand U8158 (N_8158,N_6370,N_7151);
nor U8159 (N_8159,N_6900,N_5751);
nor U8160 (N_8160,N_6976,N_5362);
nand U8161 (N_8161,N_5582,N_6115);
xnor U8162 (N_8162,N_7402,N_6509);
and U8163 (N_8163,N_6032,N_5859);
or U8164 (N_8164,N_6557,N_7373);
and U8165 (N_8165,N_7058,N_5961);
nor U8166 (N_8166,N_7393,N_5813);
nand U8167 (N_8167,N_5456,N_6600);
nor U8168 (N_8168,N_6983,N_6792);
or U8169 (N_8169,N_6232,N_5737);
or U8170 (N_8170,N_5645,N_6549);
nand U8171 (N_8171,N_5928,N_5683);
or U8172 (N_8172,N_6535,N_6007);
nor U8173 (N_8173,N_6213,N_5387);
nor U8174 (N_8174,N_6113,N_6057);
or U8175 (N_8175,N_5964,N_6949);
or U8176 (N_8176,N_5338,N_5558);
nor U8177 (N_8177,N_5350,N_7017);
and U8178 (N_8178,N_6821,N_6236);
or U8179 (N_8179,N_5856,N_5517);
or U8180 (N_8180,N_5098,N_5984);
nand U8181 (N_8181,N_6260,N_6712);
nand U8182 (N_8182,N_7136,N_5775);
and U8183 (N_8183,N_7449,N_5278);
nor U8184 (N_8184,N_5873,N_6409);
or U8185 (N_8185,N_5890,N_5878);
nand U8186 (N_8186,N_6056,N_5523);
nor U8187 (N_8187,N_5481,N_6152);
or U8188 (N_8188,N_6065,N_5642);
or U8189 (N_8189,N_5622,N_6873);
nand U8190 (N_8190,N_5044,N_5458);
nor U8191 (N_8191,N_6051,N_6081);
or U8192 (N_8192,N_6686,N_5676);
nand U8193 (N_8193,N_6410,N_5587);
nand U8194 (N_8194,N_6747,N_6675);
and U8195 (N_8195,N_5800,N_5103);
nor U8196 (N_8196,N_5474,N_6334);
and U8197 (N_8197,N_5305,N_6361);
xnor U8198 (N_8198,N_5151,N_5908);
nor U8199 (N_8199,N_5536,N_5359);
and U8200 (N_8200,N_5108,N_5778);
or U8201 (N_8201,N_6025,N_5197);
nand U8202 (N_8202,N_5990,N_5688);
nor U8203 (N_8203,N_6886,N_5204);
nand U8204 (N_8204,N_5452,N_6387);
nor U8205 (N_8205,N_7359,N_6788);
or U8206 (N_8206,N_6802,N_6323);
nor U8207 (N_8207,N_7034,N_7360);
nor U8208 (N_8208,N_7473,N_7469);
nor U8209 (N_8209,N_5036,N_6981);
nand U8210 (N_8210,N_5420,N_6532);
or U8211 (N_8211,N_6789,N_6291);
nand U8212 (N_8212,N_5216,N_5123);
or U8213 (N_8213,N_6908,N_6181);
nand U8214 (N_8214,N_6239,N_5975);
or U8215 (N_8215,N_5263,N_7208);
or U8216 (N_8216,N_6229,N_5546);
and U8217 (N_8217,N_7122,N_5624);
xor U8218 (N_8218,N_7313,N_7046);
nand U8219 (N_8219,N_6063,N_7029);
nor U8220 (N_8220,N_7131,N_7055);
nor U8221 (N_8221,N_5544,N_6914);
and U8222 (N_8222,N_7118,N_5424);
nor U8223 (N_8223,N_5825,N_6082);
nand U8224 (N_8224,N_7394,N_6043);
nor U8225 (N_8225,N_5329,N_5973);
or U8226 (N_8226,N_6031,N_7258);
nor U8227 (N_8227,N_5435,N_5763);
and U8228 (N_8228,N_5260,N_7297);
nand U8229 (N_8229,N_5047,N_5798);
nand U8230 (N_8230,N_6731,N_7331);
nor U8231 (N_8231,N_7490,N_6237);
nor U8232 (N_8232,N_6393,N_7182);
nor U8233 (N_8233,N_5627,N_6225);
nor U8234 (N_8234,N_7419,N_5264);
nor U8235 (N_8235,N_5113,N_5475);
and U8236 (N_8236,N_6905,N_7037);
or U8237 (N_8237,N_6077,N_6597);
and U8238 (N_8238,N_6337,N_5690);
or U8239 (N_8239,N_5179,N_5692);
nand U8240 (N_8240,N_6540,N_6778);
nand U8241 (N_8241,N_6559,N_7265);
or U8242 (N_8242,N_6280,N_6143);
nor U8243 (N_8243,N_6858,N_5638);
and U8244 (N_8244,N_7094,N_7231);
and U8245 (N_8245,N_6486,N_6127);
nor U8246 (N_8246,N_5585,N_5229);
nand U8247 (N_8247,N_6443,N_6444);
and U8248 (N_8248,N_5107,N_5073);
or U8249 (N_8249,N_5459,N_6390);
and U8250 (N_8250,N_7306,N_7358);
and U8251 (N_8251,N_6724,N_7019);
or U8252 (N_8252,N_7110,N_5094);
nor U8253 (N_8253,N_6940,N_7351);
nor U8254 (N_8254,N_6773,N_7245);
or U8255 (N_8255,N_5303,N_6850);
or U8256 (N_8256,N_5237,N_7400);
nor U8257 (N_8257,N_6301,N_7264);
nor U8258 (N_8258,N_7032,N_5074);
nor U8259 (N_8259,N_7329,N_5365);
or U8260 (N_8260,N_5130,N_6791);
nor U8261 (N_8261,N_6572,N_5723);
or U8262 (N_8262,N_6655,N_7237);
nor U8263 (N_8263,N_7097,N_7396);
and U8264 (N_8264,N_5643,N_6799);
nand U8265 (N_8265,N_5994,N_5657);
nor U8266 (N_8266,N_6933,N_7068);
or U8267 (N_8267,N_6885,N_6849);
or U8268 (N_8268,N_5019,N_7436);
or U8269 (N_8269,N_6611,N_6701);
or U8270 (N_8270,N_5960,N_5159);
nand U8271 (N_8271,N_6864,N_5331);
nor U8272 (N_8272,N_6829,N_6702);
and U8273 (N_8273,N_6958,N_5691);
or U8274 (N_8274,N_7285,N_7064);
nor U8275 (N_8275,N_5696,N_7088);
nand U8276 (N_8276,N_5133,N_6503);
nor U8277 (N_8277,N_5484,N_5703);
or U8278 (N_8278,N_5671,N_6944);
nand U8279 (N_8279,N_6222,N_5431);
nand U8280 (N_8280,N_6325,N_7121);
and U8281 (N_8281,N_5313,N_6694);
nand U8282 (N_8282,N_5198,N_7256);
nor U8283 (N_8283,N_6591,N_5466);
nand U8284 (N_8284,N_7383,N_5561);
nor U8285 (N_8285,N_6014,N_6479);
or U8286 (N_8286,N_5726,N_6744);
nand U8287 (N_8287,N_5482,N_6454);
nand U8288 (N_8288,N_5406,N_6921);
nor U8289 (N_8289,N_5829,N_5962);
and U8290 (N_8290,N_7044,N_6920);
nand U8291 (N_8291,N_5757,N_5386);
nor U8292 (N_8292,N_6046,N_7234);
nor U8293 (N_8293,N_7025,N_6332);
nor U8294 (N_8294,N_6215,N_5773);
nand U8295 (N_8295,N_6668,N_6910);
nand U8296 (N_8296,N_5887,N_7176);
nor U8297 (N_8297,N_5250,N_6398);
nor U8298 (N_8298,N_5621,N_6431);
nand U8299 (N_8299,N_5506,N_5089);
and U8300 (N_8300,N_5996,N_5905);
nand U8301 (N_8301,N_5711,N_7232);
nor U8302 (N_8302,N_6841,N_5742);
nor U8303 (N_8303,N_5827,N_6977);
nand U8304 (N_8304,N_7124,N_5460);
or U8305 (N_8305,N_5815,N_5882);
nor U8306 (N_8306,N_7196,N_7219);
and U8307 (N_8307,N_5985,N_7335);
or U8308 (N_8308,N_7497,N_6950);
and U8309 (N_8309,N_6194,N_7322);
nand U8310 (N_8310,N_6823,N_7372);
nor U8311 (N_8311,N_6371,N_7440);
and U8312 (N_8312,N_6129,N_6252);
nor U8313 (N_8313,N_6623,N_5086);
or U8314 (N_8314,N_6817,N_5215);
nor U8315 (N_8315,N_5408,N_6814);
nand U8316 (N_8316,N_5904,N_5025);
or U8317 (N_8317,N_6212,N_5085);
nor U8318 (N_8318,N_5341,N_6224);
nor U8319 (N_8319,N_6990,N_7030);
or U8320 (N_8320,N_7348,N_5473);
nand U8321 (N_8321,N_5306,N_6959);
and U8322 (N_8322,N_6248,N_5076);
or U8323 (N_8323,N_6469,N_6526);
and U8324 (N_8324,N_7007,N_5768);
and U8325 (N_8325,N_7274,N_5493);
nand U8326 (N_8326,N_5476,N_7398);
nor U8327 (N_8327,N_5664,N_6552);
and U8328 (N_8328,N_5441,N_6876);
or U8329 (N_8329,N_5388,N_5125);
nor U8330 (N_8330,N_5122,N_5963);
and U8331 (N_8331,N_6947,N_5507);
or U8332 (N_8332,N_7207,N_6974);
nand U8333 (N_8333,N_6342,N_6936);
or U8334 (N_8334,N_6049,N_6843);
nor U8335 (N_8335,N_7119,N_5443);
nand U8336 (N_8336,N_6415,N_5367);
and U8337 (N_8337,N_7143,N_7166);
or U8338 (N_8338,N_6736,N_5532);
or U8339 (N_8339,N_6180,N_7104);
nor U8340 (N_8340,N_5116,N_6394);
or U8341 (N_8341,N_7070,N_5043);
or U8342 (N_8342,N_5492,N_7060);
nor U8343 (N_8343,N_6941,N_5954);
nor U8344 (N_8344,N_5915,N_6221);
and U8345 (N_8345,N_6240,N_5240);
and U8346 (N_8346,N_7146,N_7263);
nand U8347 (N_8347,N_6429,N_7371);
and U8348 (N_8348,N_7499,N_7291);
xor U8349 (N_8349,N_7299,N_5945);
nand U8350 (N_8350,N_7099,N_5631);
or U8351 (N_8351,N_6270,N_6969);
nand U8352 (N_8352,N_5576,N_5402);
xnor U8353 (N_8353,N_7461,N_6650);
nand U8354 (N_8354,N_5542,N_5195);
nand U8355 (N_8355,N_5708,N_5803);
nor U8356 (N_8356,N_5913,N_6998);
or U8357 (N_8357,N_7284,N_5779);
nand U8358 (N_8358,N_5008,N_7053);
or U8359 (N_8359,N_6909,N_5674);
nand U8360 (N_8360,N_7468,N_6670);
or U8361 (N_8361,N_5442,N_5189);
and U8362 (N_8362,N_6822,N_7224);
nand U8363 (N_8363,N_5072,N_7010);
or U8364 (N_8364,N_5570,N_5070);
or U8365 (N_8365,N_6545,N_7327);
and U8366 (N_8366,N_6066,N_7363);
or U8367 (N_8367,N_6200,N_5259);
and U8368 (N_8368,N_6951,N_5029);
or U8369 (N_8369,N_5396,N_5114);
nor U8370 (N_8370,N_6809,N_5947);
nor U8371 (N_8371,N_7033,N_7432);
and U8372 (N_8372,N_7294,N_6836);
or U8373 (N_8373,N_5909,N_6755);
nor U8374 (N_8374,N_5579,N_6084);
nor U8375 (N_8375,N_7171,N_6048);
nor U8376 (N_8376,N_5847,N_6027);
or U8377 (N_8377,N_6228,N_6461);
or U8378 (N_8378,N_5575,N_6306);
or U8379 (N_8379,N_5848,N_5573);
and U8380 (N_8380,N_7310,N_6704);
and U8381 (N_8381,N_7425,N_5634);
nor U8382 (N_8382,N_6312,N_5297);
nor U8383 (N_8383,N_5830,N_6952);
or U8384 (N_8384,N_6615,N_6476);
and U8385 (N_8385,N_6629,N_5918);
nor U8386 (N_8386,N_6571,N_5257);
or U8387 (N_8387,N_5605,N_7205);
and U8388 (N_8388,N_5746,N_5380);
nor U8389 (N_8389,N_5432,N_7442);
nor U8390 (N_8390,N_6294,N_5081);
nand U8391 (N_8391,N_5364,N_5342);
nand U8392 (N_8392,N_5972,N_5451);
nor U8393 (N_8393,N_5682,N_5548);
nand U8394 (N_8394,N_6078,N_5897);
nor U8395 (N_8395,N_6960,N_6930);
or U8396 (N_8396,N_6405,N_5400);
nand U8397 (N_8397,N_5403,N_7424);
nand U8398 (N_8398,N_6104,N_6648);
nand U8399 (N_8399,N_5892,N_6785);
nand U8400 (N_8400,N_6656,N_6794);
nand U8401 (N_8401,N_6190,N_5463);
nor U8402 (N_8402,N_5021,N_5868);
nand U8403 (N_8403,N_7009,N_6380);
nand U8404 (N_8404,N_6578,N_5087);
or U8405 (N_8405,N_6842,N_6682);
and U8406 (N_8406,N_7381,N_5519);
nand U8407 (N_8407,N_7333,N_6825);
nand U8408 (N_8408,N_5180,N_7049);
and U8409 (N_8409,N_5557,N_6372);
or U8410 (N_8410,N_5455,N_7075);
nor U8411 (N_8411,N_5269,N_7204);
nand U8412 (N_8412,N_5120,N_6749);
nand U8413 (N_8413,N_7487,N_6985);
nand U8414 (N_8414,N_6075,N_6697);
or U8415 (N_8415,N_6506,N_6874);
nand U8416 (N_8416,N_5793,N_6348);
nand U8417 (N_8417,N_5957,N_6195);
nand U8418 (N_8418,N_5852,N_5796);
and U8419 (N_8419,N_6965,N_7223);
or U8420 (N_8420,N_5221,N_7246);
and U8421 (N_8421,N_7288,N_5006);
or U8422 (N_8422,N_5145,N_7477);
nand U8423 (N_8423,N_5801,N_5707);
nand U8424 (N_8424,N_7470,N_7048);
and U8425 (N_8425,N_6287,N_7086);
and U8426 (N_8426,N_7003,N_7416);
and U8427 (N_8427,N_6274,N_7282);
nor U8428 (N_8428,N_7303,N_6892);
and U8429 (N_8429,N_6363,N_5140);
nor U8430 (N_8430,N_7475,N_5743);
or U8431 (N_8431,N_7307,N_5335);
and U8432 (N_8432,N_7159,N_7133);
nand U8433 (N_8433,N_5668,N_5727);
nor U8434 (N_8434,N_6302,N_5031);
or U8435 (N_8435,N_5612,N_7085);
nand U8436 (N_8436,N_7439,N_6411);
nor U8437 (N_8437,N_5826,N_6493);
nor U8438 (N_8438,N_6308,N_5382);
nor U8439 (N_8439,N_5556,N_6972);
nand U8440 (N_8440,N_6719,N_7259);
and U8441 (N_8441,N_7213,N_5877);
and U8442 (N_8442,N_6182,N_6685);
nor U8443 (N_8443,N_5855,N_5167);
nor U8444 (N_8444,N_5732,N_5356);
nor U8445 (N_8445,N_5316,N_5412);
nand U8446 (N_8446,N_5220,N_7194);
and U8447 (N_8447,N_5236,N_5185);
nor U8448 (N_8448,N_7199,N_5853);
nand U8449 (N_8449,N_5809,N_7001);
nand U8450 (N_8450,N_5822,N_7289);
and U8451 (N_8451,N_6445,N_5991);
nor U8452 (N_8452,N_7069,N_5434);
or U8453 (N_8453,N_7454,N_5271);
nor U8454 (N_8454,N_6663,N_6699);
nand U8455 (N_8455,N_6695,N_5274);
or U8456 (N_8456,N_6857,N_5206);
or U8457 (N_8457,N_5717,N_6313);
and U8458 (N_8458,N_5978,N_7028);
nor U8459 (N_8459,N_5381,N_6245);
nand U8460 (N_8460,N_7250,N_6226);
nor U8461 (N_8461,N_7498,N_6455);
and U8462 (N_8462,N_6269,N_5698);
nor U8463 (N_8463,N_6300,N_5421);
nand U8464 (N_8464,N_6911,N_5000);
and U8465 (N_8465,N_5083,N_7036);
nand U8466 (N_8466,N_6505,N_7399);
nor U8467 (N_8467,N_6097,N_6134);
nor U8468 (N_8468,N_5135,N_6869);
or U8469 (N_8469,N_7409,N_5965);
or U8470 (N_8470,N_7020,N_7096);
nor U8471 (N_8471,N_5805,N_5563);
nand U8472 (N_8472,N_6321,N_7304);
and U8473 (N_8473,N_5193,N_5283);
nor U8474 (N_8474,N_5020,N_6630);
nor U8475 (N_8475,N_6265,N_5505);
nand U8476 (N_8476,N_5304,N_5157);
and U8477 (N_8477,N_5288,N_6259);
or U8478 (N_8478,N_6408,N_5870);
or U8479 (N_8479,N_5550,N_6923);
nor U8480 (N_8480,N_6922,N_5933);
or U8481 (N_8481,N_5479,N_6238);
or U8482 (N_8482,N_5337,N_5377);
nand U8483 (N_8483,N_5353,N_5415);
nor U8484 (N_8484,N_5590,N_6442);
or U8485 (N_8485,N_6551,N_7486);
or U8486 (N_8486,N_5068,N_7257);
xnor U8487 (N_8487,N_6653,N_5077);
or U8488 (N_8488,N_5477,N_6088);
nand U8489 (N_8489,N_6678,N_7132);
and U8490 (N_8490,N_6740,N_7318);
nor U8491 (N_8491,N_7165,N_6988);
nor U8492 (N_8492,N_6439,N_7073);
or U8493 (N_8493,N_7185,N_7427);
and U8494 (N_8494,N_6693,N_6643);
or U8495 (N_8495,N_6525,N_7262);
and U8496 (N_8496,N_5105,N_6176);
or U8497 (N_8497,N_5860,N_6946);
nand U8498 (N_8498,N_6402,N_7138);
nand U8499 (N_8499,N_6463,N_7225);
nand U8500 (N_8500,N_5489,N_6539);
nand U8501 (N_8501,N_6580,N_5276);
nand U8502 (N_8502,N_6102,N_7160);
nor U8503 (N_8503,N_5045,N_6474);
and U8504 (N_8504,N_7008,N_5772);
and U8505 (N_8505,N_5565,N_6666);
xor U8506 (N_8506,N_6038,N_6472);
nor U8507 (N_8507,N_5639,N_5647);
nor U8508 (N_8508,N_5921,N_7177);
nand U8509 (N_8509,N_5509,N_6638);
and U8510 (N_8510,N_7328,N_7261);
nand U8511 (N_8511,N_6709,N_7065);
nor U8512 (N_8512,N_6692,N_6130);
nor U8513 (N_8513,N_6116,N_6852);
and U8514 (N_8514,N_5398,N_7266);
nor U8515 (N_8515,N_7081,N_7302);
nor U8516 (N_8516,N_5997,N_5349);
nor U8517 (N_8517,N_7209,N_5438);
nand U8518 (N_8518,N_6124,N_6547);
nor U8519 (N_8519,N_6581,N_5863);
nor U8520 (N_8520,N_6889,N_6626);
nand U8521 (N_8521,N_6584,N_5416);
nand U8522 (N_8522,N_6661,N_6759);
nor U8523 (N_8523,N_6636,N_5599);
and U8524 (N_8524,N_5597,N_6339);
nand U8525 (N_8525,N_6276,N_6919);
nor U8526 (N_8526,N_7035,N_7074);
and U8527 (N_8527,N_5862,N_6856);
and U8528 (N_8528,N_6760,N_5146);
nor U8529 (N_8529,N_5574,N_7158);
and U8530 (N_8530,N_6003,N_5363);
and U8531 (N_8531,N_5014,N_6564);
and U8532 (N_8532,N_6264,N_5584);
nor U8533 (N_8533,N_6366,N_7403);
or U8534 (N_8534,N_5936,N_7187);
nand U8535 (N_8535,N_6341,N_5539);
nor U8536 (N_8536,N_7315,N_5099);
nand U8537 (N_8537,N_6076,N_6316);
and U8538 (N_8538,N_7174,N_6706);
nand U8539 (N_8539,N_5284,N_5190);
nand U8540 (N_8540,N_7478,N_7144);
and U8541 (N_8541,N_7260,N_6233);
nor U8542 (N_8542,N_5390,N_6149);
or U8543 (N_8543,N_5486,N_5212);
nor U8544 (N_8544,N_6917,N_5814);
or U8545 (N_8545,N_6953,N_6208);
or U8546 (N_8546,N_5601,N_5568);
nand U8547 (N_8547,N_7343,N_5659);
and U8548 (N_8548,N_5864,N_5254);
or U8549 (N_8549,N_6634,N_7192);
nor U8550 (N_8550,N_6575,N_6496);
and U8551 (N_8551,N_6016,N_7446);
and U8552 (N_8552,N_6510,N_5222);
or U8553 (N_8553,N_5079,N_6658);
and U8554 (N_8554,N_7226,N_6677);
and U8555 (N_8555,N_5296,N_5495);
nand U8556 (N_8556,N_7367,N_6099);
or U8557 (N_8557,N_5007,N_7311);
and U8558 (N_8558,N_6635,N_6039);
xor U8559 (N_8559,N_7433,N_5510);
nor U8560 (N_8560,N_6328,N_5900);
xor U8561 (N_8561,N_6568,N_5630);
or U8562 (N_8562,N_7395,N_5702);
or U8563 (N_8563,N_6645,N_5871);
or U8564 (N_8564,N_5749,N_7179);
or U8565 (N_8565,N_5394,N_6784);
nand U8566 (N_8566,N_5759,N_6514);
nand U8567 (N_8567,N_6989,N_5559);
nand U8568 (N_8568,N_5765,N_6612);
nor U8569 (N_8569,N_5188,N_5472);
nor U8570 (N_8570,N_5327,N_5310);
and U8571 (N_8571,N_5651,N_5967);
nand U8572 (N_8572,N_6135,N_6831);
nor U8573 (N_8573,N_5171,N_7292);
and U8574 (N_8574,N_6433,N_6887);
or U8575 (N_8575,N_6022,N_5445);
or U8576 (N_8576,N_6020,N_6683);
nand U8577 (N_8577,N_5395,N_6806);
and U8578 (N_8578,N_5134,N_5307);
and U8579 (N_8579,N_6499,N_6186);
nand U8580 (N_8580,N_7116,N_5332);
nand U8581 (N_8581,N_6585,N_5011);
nand U8582 (N_8582,N_6487,N_7120);
and U8583 (N_8583,N_6669,N_5454);
nand U8584 (N_8584,N_5001,N_6903);
and U8585 (N_8585,N_5816,N_7221);
nor U8586 (N_8586,N_5391,N_5181);
or U8587 (N_8587,N_5498,N_5567);
nand U8588 (N_8588,N_7336,N_7241);
and U8589 (N_8589,N_6798,N_6284);
nand U8590 (N_8590,N_6508,N_6502);
or U8591 (N_8591,N_5165,N_6148);
nand U8592 (N_8592,N_7155,N_5669);
and U8593 (N_8593,N_5462,N_6684);
and U8594 (N_8594,N_7337,N_6311);
nand U8595 (N_8595,N_6310,N_5710);
nor U8596 (N_8596,N_5470,N_6343);
or U8597 (N_8597,N_6281,N_6769);
or U8598 (N_8598,N_6068,N_5748);
nand U8599 (N_8599,N_5152,N_5440);
nand U8600 (N_8600,N_5496,N_5249);
or U8601 (N_8601,N_5734,N_5494);
nand U8602 (N_8602,N_5144,N_6125);
and U8603 (N_8603,N_6925,N_6644);
or U8604 (N_8604,N_7169,N_5810);
nand U8605 (N_8605,N_5528,N_5464);
and U8606 (N_8606,N_6132,N_6346);
and U8607 (N_8607,N_5665,N_7401);
and U8608 (N_8608,N_6813,N_5279);
nand U8609 (N_8609,N_7112,N_7054);
or U8610 (N_8610,N_5760,N_6691);
nor U8611 (N_8611,N_5661,N_6973);
or U8612 (N_8612,N_5213,N_6162);
or U8613 (N_8613,N_5521,N_5974);
nor U8614 (N_8614,N_5186,N_7002);
and U8615 (N_8615,N_7078,N_6730);
and U8616 (N_8616,N_5989,N_7334);
nand U8617 (N_8617,N_5993,N_5874);
nand U8618 (N_8618,N_6934,N_5069);
and U8619 (N_8619,N_5761,N_6145);
nand U8620 (N_8620,N_5511,N_5644);
nand U8621 (N_8621,N_6365,N_5520);
and U8622 (N_8622,N_6018,N_6453);
nor U8623 (N_8623,N_6543,N_6101);
and U8624 (N_8624,N_6458,N_7154);
nor U8625 (N_8625,N_6902,N_5369);
and U8626 (N_8626,N_7387,N_7186);
and U8627 (N_8627,N_7479,N_5251);
nand U8628 (N_8628,N_5752,N_5173);
and U8629 (N_8629,N_7273,N_6570);
or U8630 (N_8630,N_6753,N_5851);
nand U8631 (N_8631,N_5922,N_7459);
nor U8632 (N_8632,N_5177,N_6758);
or U8633 (N_8633,N_5549,N_6757);
nor U8634 (N_8634,N_6875,N_6733);
and U8635 (N_8635,N_5168,N_6722);
and U8636 (N_8636,N_6713,N_5817);
and U8637 (N_8637,N_5245,N_6373);
or U8638 (N_8638,N_5012,N_5005);
nor U8639 (N_8639,N_7382,N_5667);
and U8640 (N_8640,N_5209,N_7494);
nor U8641 (N_8641,N_6728,N_5697);
nor U8642 (N_8642,N_5137,N_5004);
nand U8643 (N_8643,N_5483,N_5515);
nor U8644 (N_8644,N_7127,N_5614);
nor U8645 (N_8645,N_5061,N_7045);
nand U8646 (N_8646,N_6582,N_5629);
nor U8647 (N_8647,N_6336,N_7443);
xor U8648 (N_8648,N_5034,N_7389);
or U8649 (N_8649,N_6957,N_6987);
or U8650 (N_8650,N_6428,N_5425);
and U8651 (N_8651,N_6058,N_5423);
or U8652 (N_8652,N_6975,N_7445);
nor U8653 (N_8653,N_7438,N_6092);
and U8654 (N_8654,N_6072,N_6937);
and U8655 (N_8655,N_5607,N_6470);
and U8656 (N_8656,N_6779,N_7410);
and U8657 (N_8657,N_5633,N_6801);
or U8658 (N_8658,N_7412,N_5117);
or U8659 (N_8659,N_6141,N_6432);
nand U8660 (N_8660,N_5062,N_7152);
nand U8661 (N_8661,N_7458,N_5885);
and U8662 (N_8662,N_5038,N_5169);
nor U8663 (N_8663,N_6696,N_6314);
and U8664 (N_8664,N_6352,N_5673);
and U8665 (N_8665,N_7206,N_5256);
and U8666 (N_8666,N_6716,N_6790);
nor U8667 (N_8667,N_5865,N_6555);
and U8668 (N_8668,N_5755,N_7203);
nor U8669 (N_8669,N_6416,N_6895);
nor U8670 (N_8670,N_6777,N_6191);
or U8671 (N_8671,N_7493,N_6495);
nor U8672 (N_8672,N_6085,N_5110);
and U8673 (N_8673,N_7272,N_7108);
or U8674 (N_8674,N_5385,N_6651);
nand U8675 (N_8675,N_5713,N_7422);
and U8676 (N_8676,N_7391,N_5503);
nor U8677 (N_8677,N_5780,N_6354);
nor U8678 (N_8678,N_5142,N_6369);
nor U8679 (N_8679,N_6140,N_5235);
nor U8680 (N_8680,N_5376,N_6170);
nand U8681 (N_8681,N_7191,N_7286);
or U8682 (N_8682,N_5927,N_5706);
nor U8683 (N_8683,N_7180,N_7341);
and U8684 (N_8684,N_6679,N_5397);
and U8685 (N_8685,N_5787,N_5392);
or U8686 (N_8686,N_5694,N_6931);
nand U8687 (N_8687,N_5538,N_7496);
nand U8688 (N_8688,N_6710,N_6620);
nor U8689 (N_8689,N_6647,N_7355);
and U8690 (N_8690,N_6674,N_6513);
nand U8691 (N_8691,N_6478,N_6504);
nand U8692 (N_8692,N_6574,N_6093);
xor U8693 (N_8693,N_6360,N_6290);
and U8694 (N_8694,N_6490,N_5247);
or U8695 (N_8695,N_6122,N_5685);
nor U8696 (N_8696,N_5540,N_6717);
and U8697 (N_8697,N_7027,N_6422);
and U8698 (N_8698,N_6512,N_5770);
nor U8699 (N_8699,N_6423,N_7460);
and U8700 (N_8700,N_6054,N_5207);
nor U8701 (N_8701,N_5806,N_7130);
nand U8702 (N_8702,N_7356,N_6015);
or U8703 (N_8703,N_5602,N_6531);
nor U8704 (N_8704,N_5777,N_6939);
nand U8705 (N_8705,N_5071,N_5720);
or U8706 (N_8706,N_5995,N_7484);
nor U8707 (N_8707,N_6711,N_5893);
or U8708 (N_8708,N_7423,N_5191);
nand U8709 (N_8709,N_5504,N_5571);
nand U8710 (N_8710,N_5433,N_5224);
nand U8711 (N_8711,N_5718,N_6275);
nand U8712 (N_8712,N_7271,N_5372);
nor U8713 (N_8713,N_5850,N_5252);
nand U8714 (N_8714,N_5200,N_6255);
and U8715 (N_8715,N_6599,N_5898);
and U8716 (N_8716,N_5049,N_5566);
or U8717 (N_8717,N_6350,N_7352);
xnor U8718 (N_8718,N_7084,N_5148);
or U8719 (N_8719,N_5578,N_7491);
nand U8720 (N_8720,N_6449,N_6840);
nor U8721 (N_8721,N_7317,N_7072);
nand U8722 (N_8722,N_6418,N_6839);
nor U8723 (N_8723,N_6425,N_7178);
and U8724 (N_8724,N_6282,N_5811);
nand U8725 (N_8725,N_7430,N_6062);
nor U8726 (N_8726,N_5015,N_5545);
and U8727 (N_8727,N_7451,N_6657);
or U8728 (N_8728,N_5295,N_6680);
nor U8729 (N_8729,N_5745,N_6357);
and U8730 (N_8730,N_5730,N_5823);
nor U8731 (N_8731,N_6610,N_5527);
nand U8732 (N_8732,N_6589,N_5291);
and U8733 (N_8733,N_6261,N_5837);
or U8734 (N_8734,N_6330,N_7456);
and U8735 (N_8735,N_5286,N_6329);
nor U8736 (N_8736,N_7040,N_5328);
nor U8737 (N_8737,N_6353,N_6756);
nand U8738 (N_8738,N_5914,N_6220);
and U8739 (N_8739,N_5903,N_7157);
or U8740 (N_8740,N_6605,N_5626);
nand U8741 (N_8741,N_5056,N_5242);
or U8742 (N_8742,N_6475,N_6318);
nand U8743 (N_8743,N_5461,N_7188);
or U8744 (N_8744,N_6607,N_6888);
or U8745 (N_8745,N_6561,N_6861);
nor U8746 (N_8746,N_7368,N_7051);
nand U8747 (N_8747,N_6118,N_5595);
nand U8748 (N_8748,N_5225,N_5050);
nand U8749 (N_8749,N_5028,N_7047);
and U8750 (N_8750,N_6623,N_6600);
or U8751 (N_8751,N_5403,N_6062);
nand U8752 (N_8752,N_6666,N_6964);
and U8753 (N_8753,N_6584,N_6827);
nor U8754 (N_8754,N_6950,N_5537);
nor U8755 (N_8755,N_6925,N_6910);
nor U8756 (N_8756,N_5689,N_5744);
nor U8757 (N_8757,N_5280,N_7377);
nor U8758 (N_8758,N_5603,N_6999);
nor U8759 (N_8759,N_5944,N_5395);
and U8760 (N_8760,N_7080,N_5066);
nand U8761 (N_8761,N_5269,N_6431);
nor U8762 (N_8762,N_7169,N_7285);
nand U8763 (N_8763,N_6241,N_7178);
nand U8764 (N_8764,N_5682,N_6371);
and U8765 (N_8765,N_5318,N_6641);
and U8766 (N_8766,N_5468,N_6783);
nand U8767 (N_8767,N_5982,N_6231);
or U8768 (N_8768,N_5198,N_5450);
nor U8769 (N_8769,N_5110,N_5857);
and U8770 (N_8770,N_5803,N_7292);
nand U8771 (N_8771,N_5417,N_7267);
and U8772 (N_8772,N_5960,N_5697);
and U8773 (N_8773,N_5883,N_5742);
and U8774 (N_8774,N_6998,N_6562);
and U8775 (N_8775,N_5177,N_6608);
nand U8776 (N_8776,N_6956,N_7428);
or U8777 (N_8777,N_5176,N_6500);
and U8778 (N_8778,N_7419,N_7288);
nand U8779 (N_8779,N_7185,N_5865);
nand U8780 (N_8780,N_5330,N_5286);
and U8781 (N_8781,N_5126,N_5814);
or U8782 (N_8782,N_6103,N_6333);
and U8783 (N_8783,N_6156,N_5063);
nand U8784 (N_8784,N_5243,N_5116);
nor U8785 (N_8785,N_6806,N_5517);
and U8786 (N_8786,N_7115,N_5692);
nor U8787 (N_8787,N_5738,N_6770);
and U8788 (N_8788,N_6839,N_5266);
nand U8789 (N_8789,N_6938,N_5945);
and U8790 (N_8790,N_5837,N_7359);
or U8791 (N_8791,N_7164,N_7496);
and U8792 (N_8792,N_7455,N_5884);
nor U8793 (N_8793,N_6702,N_5478);
nand U8794 (N_8794,N_5365,N_6824);
or U8795 (N_8795,N_7005,N_5814);
or U8796 (N_8796,N_6400,N_6255);
nor U8797 (N_8797,N_6201,N_6551);
or U8798 (N_8798,N_7480,N_5597);
nand U8799 (N_8799,N_5067,N_7138);
nand U8800 (N_8800,N_6104,N_6879);
nor U8801 (N_8801,N_5807,N_7314);
or U8802 (N_8802,N_6734,N_6386);
and U8803 (N_8803,N_5106,N_5988);
nor U8804 (N_8804,N_5508,N_7231);
or U8805 (N_8805,N_7148,N_7079);
nor U8806 (N_8806,N_5666,N_5619);
or U8807 (N_8807,N_6052,N_5516);
and U8808 (N_8808,N_6034,N_5163);
nand U8809 (N_8809,N_6714,N_5035);
or U8810 (N_8810,N_6630,N_7273);
and U8811 (N_8811,N_6602,N_6930);
nand U8812 (N_8812,N_5172,N_5315);
nand U8813 (N_8813,N_6108,N_7323);
and U8814 (N_8814,N_5170,N_6429);
nor U8815 (N_8815,N_6031,N_6129);
nor U8816 (N_8816,N_5258,N_5118);
or U8817 (N_8817,N_7137,N_5814);
nor U8818 (N_8818,N_5347,N_6434);
nor U8819 (N_8819,N_6649,N_7017);
and U8820 (N_8820,N_6509,N_6889);
or U8821 (N_8821,N_6177,N_5208);
nand U8822 (N_8822,N_5838,N_6334);
nor U8823 (N_8823,N_6688,N_6317);
or U8824 (N_8824,N_7343,N_5523);
nor U8825 (N_8825,N_5668,N_5688);
and U8826 (N_8826,N_6571,N_5469);
nor U8827 (N_8827,N_6171,N_7401);
xor U8828 (N_8828,N_6917,N_6134);
nand U8829 (N_8829,N_7287,N_6251);
nor U8830 (N_8830,N_5918,N_6505);
nor U8831 (N_8831,N_7091,N_6250);
and U8832 (N_8832,N_5390,N_6255);
and U8833 (N_8833,N_5788,N_7191);
nor U8834 (N_8834,N_6747,N_5619);
nor U8835 (N_8835,N_5861,N_7243);
and U8836 (N_8836,N_6717,N_5954);
nor U8837 (N_8837,N_7367,N_6118);
or U8838 (N_8838,N_7140,N_7112);
nor U8839 (N_8839,N_6454,N_6640);
nor U8840 (N_8840,N_5431,N_6314);
or U8841 (N_8841,N_5141,N_6041);
nor U8842 (N_8842,N_5431,N_5093);
nand U8843 (N_8843,N_6598,N_6574);
or U8844 (N_8844,N_7290,N_6509);
or U8845 (N_8845,N_6585,N_5825);
nor U8846 (N_8846,N_6943,N_6400);
and U8847 (N_8847,N_7165,N_6006);
nor U8848 (N_8848,N_7374,N_6996);
xnor U8849 (N_8849,N_5685,N_6111);
and U8850 (N_8850,N_6413,N_6911);
or U8851 (N_8851,N_5590,N_6558);
nand U8852 (N_8852,N_5367,N_5592);
and U8853 (N_8853,N_6641,N_5573);
or U8854 (N_8854,N_5492,N_6421);
nand U8855 (N_8855,N_5731,N_5879);
or U8856 (N_8856,N_5336,N_6770);
or U8857 (N_8857,N_5159,N_7119);
or U8858 (N_8858,N_7022,N_7250);
nor U8859 (N_8859,N_5939,N_6479);
and U8860 (N_8860,N_6270,N_5311);
and U8861 (N_8861,N_7148,N_5347);
nor U8862 (N_8862,N_5556,N_6732);
and U8863 (N_8863,N_5062,N_5558);
nor U8864 (N_8864,N_5535,N_6217);
nor U8865 (N_8865,N_6091,N_6218);
or U8866 (N_8866,N_6108,N_7463);
or U8867 (N_8867,N_7274,N_6363);
xnor U8868 (N_8868,N_6592,N_7439);
nand U8869 (N_8869,N_5355,N_5812);
nor U8870 (N_8870,N_5312,N_6597);
and U8871 (N_8871,N_7408,N_5133);
nor U8872 (N_8872,N_5410,N_5343);
or U8873 (N_8873,N_6350,N_6630);
nor U8874 (N_8874,N_5407,N_7108);
nor U8875 (N_8875,N_6758,N_6504);
and U8876 (N_8876,N_6359,N_6386);
and U8877 (N_8877,N_5256,N_5091);
and U8878 (N_8878,N_6910,N_6623);
or U8879 (N_8879,N_5843,N_5316);
or U8880 (N_8880,N_5792,N_6771);
nor U8881 (N_8881,N_5589,N_7367);
and U8882 (N_8882,N_5257,N_5135);
nor U8883 (N_8883,N_5798,N_7491);
nor U8884 (N_8884,N_6288,N_6471);
or U8885 (N_8885,N_6362,N_6454);
nand U8886 (N_8886,N_6240,N_7181);
nand U8887 (N_8887,N_7425,N_5600);
or U8888 (N_8888,N_7105,N_6024);
and U8889 (N_8889,N_7148,N_6961);
or U8890 (N_8890,N_7493,N_5108);
or U8891 (N_8891,N_6324,N_7068);
nor U8892 (N_8892,N_5039,N_7227);
nor U8893 (N_8893,N_5837,N_5536);
nor U8894 (N_8894,N_7286,N_5723);
nand U8895 (N_8895,N_6987,N_5216);
nor U8896 (N_8896,N_7030,N_7458);
nand U8897 (N_8897,N_5477,N_7215);
nor U8898 (N_8898,N_5269,N_6944);
nand U8899 (N_8899,N_5869,N_5059);
and U8900 (N_8900,N_7258,N_6279);
and U8901 (N_8901,N_7139,N_5759);
nor U8902 (N_8902,N_6777,N_5009);
or U8903 (N_8903,N_6559,N_5171);
or U8904 (N_8904,N_5020,N_5381);
nand U8905 (N_8905,N_7370,N_6610);
nor U8906 (N_8906,N_6214,N_6745);
nand U8907 (N_8907,N_7106,N_5291);
or U8908 (N_8908,N_5409,N_7462);
nor U8909 (N_8909,N_5519,N_6340);
or U8910 (N_8910,N_5268,N_5658);
xor U8911 (N_8911,N_7169,N_6937);
and U8912 (N_8912,N_6347,N_6786);
or U8913 (N_8913,N_6544,N_7402);
or U8914 (N_8914,N_5555,N_6493);
or U8915 (N_8915,N_5377,N_5720);
nor U8916 (N_8916,N_6551,N_6138);
or U8917 (N_8917,N_6825,N_5234);
and U8918 (N_8918,N_5259,N_5020);
or U8919 (N_8919,N_6373,N_6038);
and U8920 (N_8920,N_5556,N_6576);
nor U8921 (N_8921,N_7080,N_5443);
or U8922 (N_8922,N_7381,N_5295);
nand U8923 (N_8923,N_6871,N_7310);
or U8924 (N_8924,N_6405,N_6299);
and U8925 (N_8925,N_5152,N_6398);
and U8926 (N_8926,N_6286,N_5004);
and U8927 (N_8927,N_5477,N_5098);
and U8928 (N_8928,N_7160,N_7223);
nor U8929 (N_8929,N_6548,N_5111);
nor U8930 (N_8930,N_6034,N_5197);
or U8931 (N_8931,N_7058,N_7037);
nor U8932 (N_8932,N_5659,N_5545);
nand U8933 (N_8933,N_6571,N_5106);
nor U8934 (N_8934,N_6916,N_5523);
or U8935 (N_8935,N_5479,N_6120);
nand U8936 (N_8936,N_6734,N_6499);
nand U8937 (N_8937,N_6732,N_7266);
and U8938 (N_8938,N_6298,N_7070);
nand U8939 (N_8939,N_5677,N_6549);
and U8940 (N_8940,N_5422,N_5323);
nor U8941 (N_8941,N_7228,N_6050);
nand U8942 (N_8942,N_5140,N_6425);
nand U8943 (N_8943,N_6542,N_7448);
or U8944 (N_8944,N_5829,N_6123);
nor U8945 (N_8945,N_6219,N_6988);
nand U8946 (N_8946,N_6993,N_5516);
nand U8947 (N_8947,N_6854,N_6400);
and U8948 (N_8948,N_5090,N_6969);
nand U8949 (N_8949,N_7145,N_5768);
and U8950 (N_8950,N_6317,N_5896);
nor U8951 (N_8951,N_7118,N_5602);
and U8952 (N_8952,N_6486,N_5486);
nor U8953 (N_8953,N_6058,N_6875);
nand U8954 (N_8954,N_7189,N_6236);
nand U8955 (N_8955,N_5553,N_6547);
or U8956 (N_8956,N_5440,N_5580);
nand U8957 (N_8957,N_6218,N_6674);
nor U8958 (N_8958,N_5016,N_6267);
nand U8959 (N_8959,N_5729,N_7215);
nand U8960 (N_8960,N_6745,N_7119);
nand U8961 (N_8961,N_6469,N_5745);
nand U8962 (N_8962,N_6860,N_6915);
nand U8963 (N_8963,N_6697,N_7036);
or U8964 (N_8964,N_5738,N_6706);
nor U8965 (N_8965,N_7343,N_6970);
nand U8966 (N_8966,N_6068,N_5160);
nand U8967 (N_8967,N_5351,N_6970);
or U8968 (N_8968,N_5963,N_5336);
or U8969 (N_8969,N_5806,N_6811);
nand U8970 (N_8970,N_6560,N_6720);
nand U8971 (N_8971,N_5773,N_5945);
and U8972 (N_8972,N_6267,N_5089);
nand U8973 (N_8973,N_5326,N_6340);
and U8974 (N_8974,N_6625,N_6324);
or U8975 (N_8975,N_5016,N_5163);
or U8976 (N_8976,N_6008,N_7053);
and U8977 (N_8977,N_7342,N_5885);
or U8978 (N_8978,N_6519,N_5720);
nand U8979 (N_8979,N_7313,N_5370);
or U8980 (N_8980,N_5492,N_5783);
and U8981 (N_8981,N_5723,N_7467);
or U8982 (N_8982,N_5532,N_7186);
or U8983 (N_8983,N_5890,N_5269);
and U8984 (N_8984,N_6603,N_6001);
and U8985 (N_8985,N_6737,N_5947);
nand U8986 (N_8986,N_5834,N_6980);
nand U8987 (N_8987,N_5321,N_7410);
and U8988 (N_8988,N_6684,N_5617);
nor U8989 (N_8989,N_6181,N_5504);
and U8990 (N_8990,N_5522,N_5986);
nor U8991 (N_8991,N_6989,N_5021);
nor U8992 (N_8992,N_5983,N_6542);
or U8993 (N_8993,N_5885,N_7092);
and U8994 (N_8994,N_6105,N_7343);
nand U8995 (N_8995,N_6259,N_5256);
and U8996 (N_8996,N_7387,N_7111);
or U8997 (N_8997,N_5665,N_6175);
and U8998 (N_8998,N_7403,N_5320);
and U8999 (N_8999,N_6843,N_5587);
and U9000 (N_9000,N_5962,N_6627);
or U9001 (N_9001,N_6278,N_7367);
or U9002 (N_9002,N_6450,N_5543);
nor U9003 (N_9003,N_6473,N_5022);
nor U9004 (N_9004,N_6096,N_6826);
and U9005 (N_9005,N_5911,N_5736);
or U9006 (N_9006,N_7466,N_7214);
nor U9007 (N_9007,N_6840,N_5125);
and U9008 (N_9008,N_5713,N_5831);
or U9009 (N_9009,N_5652,N_6102);
nor U9010 (N_9010,N_6202,N_7150);
nor U9011 (N_9011,N_7485,N_6742);
nor U9012 (N_9012,N_5522,N_6377);
or U9013 (N_9013,N_5344,N_7381);
nand U9014 (N_9014,N_5486,N_6793);
nand U9015 (N_9015,N_7475,N_6768);
or U9016 (N_9016,N_5179,N_7091);
and U9017 (N_9017,N_6092,N_7105);
nor U9018 (N_9018,N_6627,N_5446);
or U9019 (N_9019,N_6113,N_6834);
nand U9020 (N_9020,N_5953,N_5756);
or U9021 (N_9021,N_6711,N_6085);
or U9022 (N_9022,N_6083,N_5896);
nor U9023 (N_9023,N_5530,N_6544);
or U9024 (N_9024,N_6666,N_6359);
or U9025 (N_9025,N_5997,N_5909);
nand U9026 (N_9026,N_6957,N_6794);
or U9027 (N_9027,N_5030,N_7117);
or U9028 (N_9028,N_6493,N_5056);
or U9029 (N_9029,N_7004,N_5361);
nor U9030 (N_9030,N_6555,N_6480);
and U9031 (N_9031,N_6827,N_7173);
nor U9032 (N_9032,N_6059,N_7246);
nand U9033 (N_9033,N_7401,N_7074);
nor U9034 (N_9034,N_6866,N_5956);
nand U9035 (N_9035,N_7235,N_5864);
and U9036 (N_9036,N_5157,N_5855);
nand U9037 (N_9037,N_6005,N_5260);
nand U9038 (N_9038,N_6174,N_6562);
nand U9039 (N_9039,N_6346,N_7457);
or U9040 (N_9040,N_5912,N_5614);
nand U9041 (N_9041,N_5330,N_5110);
or U9042 (N_9042,N_6603,N_6153);
nor U9043 (N_9043,N_6843,N_6659);
nor U9044 (N_9044,N_7238,N_5061);
or U9045 (N_9045,N_6632,N_6186);
nand U9046 (N_9046,N_5553,N_5027);
nand U9047 (N_9047,N_6658,N_7412);
or U9048 (N_9048,N_5985,N_7056);
and U9049 (N_9049,N_6203,N_7049);
nor U9050 (N_9050,N_7155,N_6729);
nand U9051 (N_9051,N_6825,N_7408);
nor U9052 (N_9052,N_5510,N_6999);
or U9053 (N_9053,N_6166,N_5358);
nand U9054 (N_9054,N_7313,N_7489);
nor U9055 (N_9055,N_7287,N_6225);
nand U9056 (N_9056,N_6262,N_7476);
nand U9057 (N_9057,N_5940,N_6654);
nor U9058 (N_9058,N_7028,N_6449);
nand U9059 (N_9059,N_5206,N_5530);
nor U9060 (N_9060,N_6856,N_7325);
nor U9061 (N_9061,N_5371,N_6067);
nand U9062 (N_9062,N_5344,N_6029);
and U9063 (N_9063,N_7175,N_6927);
or U9064 (N_9064,N_6960,N_6317);
xor U9065 (N_9065,N_6033,N_5654);
and U9066 (N_9066,N_5166,N_6731);
or U9067 (N_9067,N_6527,N_6311);
nor U9068 (N_9068,N_7245,N_6149);
nand U9069 (N_9069,N_5482,N_6144);
or U9070 (N_9070,N_5090,N_6594);
nand U9071 (N_9071,N_5574,N_5804);
nand U9072 (N_9072,N_6104,N_5563);
nand U9073 (N_9073,N_5513,N_7489);
nor U9074 (N_9074,N_5326,N_7438);
nand U9075 (N_9075,N_5653,N_5773);
or U9076 (N_9076,N_5303,N_6368);
or U9077 (N_9077,N_5512,N_6408);
nand U9078 (N_9078,N_5613,N_6923);
nand U9079 (N_9079,N_6112,N_7076);
and U9080 (N_9080,N_5924,N_5349);
nor U9081 (N_9081,N_5836,N_7249);
nand U9082 (N_9082,N_5075,N_5921);
and U9083 (N_9083,N_5606,N_7124);
and U9084 (N_9084,N_7316,N_5734);
or U9085 (N_9085,N_6436,N_7315);
or U9086 (N_9086,N_5209,N_6837);
nor U9087 (N_9087,N_7073,N_6240);
nand U9088 (N_9088,N_5137,N_6363);
nor U9089 (N_9089,N_7062,N_7414);
nor U9090 (N_9090,N_6176,N_5842);
and U9091 (N_9091,N_5429,N_6351);
or U9092 (N_9092,N_7220,N_6335);
nand U9093 (N_9093,N_5455,N_5391);
or U9094 (N_9094,N_5446,N_5289);
nand U9095 (N_9095,N_6914,N_6161);
xor U9096 (N_9096,N_5717,N_5808);
nor U9097 (N_9097,N_5169,N_6626);
nand U9098 (N_9098,N_5174,N_6490);
nor U9099 (N_9099,N_7093,N_5326);
nor U9100 (N_9100,N_6697,N_7451);
and U9101 (N_9101,N_7350,N_6083);
or U9102 (N_9102,N_5181,N_6958);
and U9103 (N_9103,N_5723,N_5981);
and U9104 (N_9104,N_5357,N_5276);
or U9105 (N_9105,N_6675,N_5729);
or U9106 (N_9106,N_7204,N_5778);
and U9107 (N_9107,N_7459,N_7051);
nand U9108 (N_9108,N_6957,N_7406);
or U9109 (N_9109,N_6188,N_6251);
nand U9110 (N_9110,N_7004,N_7106);
or U9111 (N_9111,N_6835,N_6412);
and U9112 (N_9112,N_6907,N_7237);
xnor U9113 (N_9113,N_7401,N_5173);
xnor U9114 (N_9114,N_5179,N_7477);
nand U9115 (N_9115,N_5984,N_5044);
nand U9116 (N_9116,N_5768,N_5043);
and U9117 (N_9117,N_6230,N_6441);
and U9118 (N_9118,N_5684,N_5915);
or U9119 (N_9119,N_7359,N_5676);
nand U9120 (N_9120,N_6754,N_6932);
or U9121 (N_9121,N_6791,N_6290);
nand U9122 (N_9122,N_6800,N_5999);
nand U9123 (N_9123,N_5310,N_6375);
nand U9124 (N_9124,N_6470,N_5375);
and U9125 (N_9125,N_5031,N_5057);
nand U9126 (N_9126,N_6647,N_6724);
nor U9127 (N_9127,N_5843,N_7407);
nand U9128 (N_9128,N_7072,N_6561);
nor U9129 (N_9129,N_6893,N_5764);
nor U9130 (N_9130,N_6226,N_5628);
or U9131 (N_9131,N_5121,N_5369);
nand U9132 (N_9132,N_7230,N_7353);
and U9133 (N_9133,N_5824,N_5338);
nor U9134 (N_9134,N_6354,N_7051);
or U9135 (N_9135,N_5908,N_7303);
nand U9136 (N_9136,N_6550,N_6942);
and U9137 (N_9137,N_7283,N_5667);
nand U9138 (N_9138,N_5217,N_5087);
and U9139 (N_9139,N_5342,N_5059);
nor U9140 (N_9140,N_7076,N_5825);
nor U9141 (N_9141,N_5333,N_7309);
nor U9142 (N_9142,N_5890,N_6708);
and U9143 (N_9143,N_5116,N_5841);
nor U9144 (N_9144,N_5518,N_6365);
or U9145 (N_9145,N_7108,N_6968);
and U9146 (N_9146,N_6396,N_5960);
or U9147 (N_9147,N_5037,N_6122);
nand U9148 (N_9148,N_5617,N_6754);
and U9149 (N_9149,N_5017,N_6601);
nor U9150 (N_9150,N_6434,N_5664);
nor U9151 (N_9151,N_7134,N_5602);
nand U9152 (N_9152,N_7024,N_6504);
or U9153 (N_9153,N_5169,N_7056);
nand U9154 (N_9154,N_6073,N_6366);
nor U9155 (N_9155,N_5862,N_7447);
and U9156 (N_9156,N_7396,N_7128);
nor U9157 (N_9157,N_5760,N_6763);
and U9158 (N_9158,N_6264,N_5809);
nor U9159 (N_9159,N_7060,N_6971);
nand U9160 (N_9160,N_6916,N_5604);
nand U9161 (N_9161,N_7169,N_6340);
and U9162 (N_9162,N_6116,N_6429);
or U9163 (N_9163,N_6899,N_6180);
or U9164 (N_9164,N_5135,N_7367);
and U9165 (N_9165,N_5634,N_5316);
nor U9166 (N_9166,N_7244,N_6646);
and U9167 (N_9167,N_6431,N_7359);
xnor U9168 (N_9168,N_5254,N_6572);
and U9169 (N_9169,N_5905,N_5480);
nor U9170 (N_9170,N_6195,N_5254);
and U9171 (N_9171,N_5621,N_6005);
or U9172 (N_9172,N_6022,N_5204);
nand U9173 (N_9173,N_7065,N_5929);
nand U9174 (N_9174,N_6685,N_5977);
or U9175 (N_9175,N_6782,N_6088);
nor U9176 (N_9176,N_6501,N_7207);
nor U9177 (N_9177,N_5964,N_7473);
and U9178 (N_9178,N_6401,N_6312);
nor U9179 (N_9179,N_6868,N_5833);
nand U9180 (N_9180,N_6348,N_7004);
nor U9181 (N_9181,N_5402,N_6560);
or U9182 (N_9182,N_7147,N_5063);
and U9183 (N_9183,N_5139,N_5715);
nor U9184 (N_9184,N_6693,N_6299);
and U9185 (N_9185,N_5858,N_6622);
nor U9186 (N_9186,N_5857,N_5279);
and U9187 (N_9187,N_5342,N_5812);
nand U9188 (N_9188,N_6806,N_7397);
xor U9189 (N_9189,N_6543,N_6232);
nand U9190 (N_9190,N_5046,N_5542);
nand U9191 (N_9191,N_5342,N_6523);
or U9192 (N_9192,N_6557,N_6228);
nand U9193 (N_9193,N_7373,N_7155);
nand U9194 (N_9194,N_6677,N_6682);
or U9195 (N_9195,N_6205,N_5443);
nand U9196 (N_9196,N_7261,N_5615);
nand U9197 (N_9197,N_6373,N_6184);
and U9198 (N_9198,N_5941,N_7000);
and U9199 (N_9199,N_7183,N_7409);
nand U9200 (N_9200,N_5785,N_7215);
nor U9201 (N_9201,N_5360,N_5552);
or U9202 (N_9202,N_5582,N_5314);
nand U9203 (N_9203,N_5621,N_5194);
nand U9204 (N_9204,N_7335,N_5701);
nand U9205 (N_9205,N_5410,N_5579);
and U9206 (N_9206,N_6867,N_5971);
and U9207 (N_9207,N_6024,N_6147);
nor U9208 (N_9208,N_5081,N_5599);
or U9209 (N_9209,N_5040,N_5022);
nor U9210 (N_9210,N_6262,N_6357);
nor U9211 (N_9211,N_7491,N_6617);
nor U9212 (N_9212,N_6772,N_5315);
and U9213 (N_9213,N_7245,N_7310);
or U9214 (N_9214,N_6644,N_5292);
and U9215 (N_9215,N_6730,N_6940);
and U9216 (N_9216,N_6975,N_7106);
and U9217 (N_9217,N_5919,N_5371);
and U9218 (N_9218,N_5749,N_7408);
and U9219 (N_9219,N_7307,N_6825);
or U9220 (N_9220,N_7007,N_7434);
nor U9221 (N_9221,N_7202,N_7496);
or U9222 (N_9222,N_6816,N_5633);
nand U9223 (N_9223,N_5032,N_5382);
nor U9224 (N_9224,N_5887,N_6766);
and U9225 (N_9225,N_6119,N_5946);
nand U9226 (N_9226,N_6914,N_7084);
or U9227 (N_9227,N_6188,N_5688);
and U9228 (N_9228,N_5321,N_5860);
nand U9229 (N_9229,N_7200,N_6894);
and U9230 (N_9230,N_6625,N_7079);
or U9231 (N_9231,N_6965,N_5734);
or U9232 (N_9232,N_6902,N_5884);
nor U9233 (N_9233,N_6777,N_7303);
nand U9234 (N_9234,N_5575,N_7337);
and U9235 (N_9235,N_5118,N_6130);
nor U9236 (N_9236,N_5205,N_6826);
or U9237 (N_9237,N_7104,N_6059);
or U9238 (N_9238,N_6952,N_6457);
or U9239 (N_9239,N_7048,N_7184);
nor U9240 (N_9240,N_6100,N_7399);
and U9241 (N_9241,N_6822,N_5607);
and U9242 (N_9242,N_6487,N_5317);
and U9243 (N_9243,N_6107,N_5408);
nand U9244 (N_9244,N_5379,N_6939);
nor U9245 (N_9245,N_6158,N_5512);
nand U9246 (N_9246,N_5131,N_5218);
xor U9247 (N_9247,N_6754,N_5392);
nor U9248 (N_9248,N_6994,N_5826);
nand U9249 (N_9249,N_5876,N_6748);
and U9250 (N_9250,N_7064,N_5893);
nand U9251 (N_9251,N_7119,N_6906);
and U9252 (N_9252,N_5205,N_6702);
or U9253 (N_9253,N_5832,N_6760);
and U9254 (N_9254,N_7351,N_7052);
or U9255 (N_9255,N_6211,N_7432);
or U9256 (N_9256,N_6750,N_6912);
nand U9257 (N_9257,N_5470,N_7111);
and U9258 (N_9258,N_7326,N_7371);
nand U9259 (N_9259,N_7343,N_6930);
nor U9260 (N_9260,N_5436,N_7463);
nor U9261 (N_9261,N_6143,N_6739);
or U9262 (N_9262,N_5378,N_5658);
nand U9263 (N_9263,N_6641,N_5546);
or U9264 (N_9264,N_6905,N_6848);
nand U9265 (N_9265,N_6321,N_5657);
or U9266 (N_9266,N_7055,N_7304);
nor U9267 (N_9267,N_6632,N_5598);
and U9268 (N_9268,N_6713,N_5057);
or U9269 (N_9269,N_5627,N_7317);
nand U9270 (N_9270,N_6614,N_5216);
nor U9271 (N_9271,N_7204,N_7149);
and U9272 (N_9272,N_6153,N_5481);
or U9273 (N_9273,N_5591,N_5214);
nor U9274 (N_9274,N_6046,N_6855);
and U9275 (N_9275,N_5955,N_6058);
and U9276 (N_9276,N_5675,N_6879);
nor U9277 (N_9277,N_5392,N_6768);
nand U9278 (N_9278,N_6123,N_7320);
or U9279 (N_9279,N_6199,N_6718);
nor U9280 (N_9280,N_5310,N_5156);
nand U9281 (N_9281,N_7303,N_5985);
nor U9282 (N_9282,N_5579,N_6842);
or U9283 (N_9283,N_6904,N_6441);
and U9284 (N_9284,N_6297,N_5025);
and U9285 (N_9285,N_6660,N_5721);
nand U9286 (N_9286,N_6685,N_6902);
nor U9287 (N_9287,N_6372,N_6484);
and U9288 (N_9288,N_5166,N_5176);
nor U9289 (N_9289,N_5696,N_7050);
nor U9290 (N_9290,N_7127,N_5505);
or U9291 (N_9291,N_6542,N_5596);
or U9292 (N_9292,N_7467,N_6554);
or U9293 (N_9293,N_5588,N_7458);
or U9294 (N_9294,N_7148,N_6929);
and U9295 (N_9295,N_7144,N_5651);
nand U9296 (N_9296,N_7264,N_6608);
nand U9297 (N_9297,N_6718,N_6867);
nand U9298 (N_9298,N_7405,N_5580);
nand U9299 (N_9299,N_5135,N_5413);
nand U9300 (N_9300,N_6932,N_6268);
or U9301 (N_9301,N_6623,N_5119);
nand U9302 (N_9302,N_6746,N_7120);
nand U9303 (N_9303,N_6418,N_7190);
or U9304 (N_9304,N_6503,N_7392);
and U9305 (N_9305,N_6053,N_5767);
and U9306 (N_9306,N_5970,N_7256);
or U9307 (N_9307,N_6217,N_6067);
nor U9308 (N_9308,N_6576,N_5493);
and U9309 (N_9309,N_5628,N_5125);
and U9310 (N_9310,N_6773,N_7024);
and U9311 (N_9311,N_7316,N_5736);
or U9312 (N_9312,N_5637,N_7215);
or U9313 (N_9313,N_5990,N_6178);
nand U9314 (N_9314,N_7266,N_6086);
and U9315 (N_9315,N_5163,N_5542);
nand U9316 (N_9316,N_6669,N_6082);
nand U9317 (N_9317,N_7151,N_6876);
xor U9318 (N_9318,N_6203,N_5922);
nor U9319 (N_9319,N_6865,N_5705);
nor U9320 (N_9320,N_6511,N_6529);
or U9321 (N_9321,N_6895,N_5075);
and U9322 (N_9322,N_7188,N_5790);
and U9323 (N_9323,N_6479,N_7083);
or U9324 (N_9324,N_7270,N_7188);
or U9325 (N_9325,N_5905,N_5226);
nand U9326 (N_9326,N_7217,N_6814);
and U9327 (N_9327,N_7228,N_5103);
nand U9328 (N_9328,N_6477,N_6027);
nor U9329 (N_9329,N_5332,N_6755);
nor U9330 (N_9330,N_6945,N_7308);
and U9331 (N_9331,N_5141,N_6378);
or U9332 (N_9332,N_6177,N_7280);
or U9333 (N_9333,N_6637,N_5872);
or U9334 (N_9334,N_5638,N_7279);
nor U9335 (N_9335,N_5604,N_6466);
nand U9336 (N_9336,N_5293,N_5635);
or U9337 (N_9337,N_6709,N_7337);
nor U9338 (N_9338,N_7295,N_7360);
nand U9339 (N_9339,N_7001,N_5054);
and U9340 (N_9340,N_6518,N_5350);
nor U9341 (N_9341,N_6191,N_5083);
and U9342 (N_9342,N_6148,N_5619);
nand U9343 (N_9343,N_6579,N_5688);
or U9344 (N_9344,N_5758,N_7354);
nand U9345 (N_9345,N_6901,N_5013);
nor U9346 (N_9346,N_6694,N_6138);
nor U9347 (N_9347,N_5930,N_5495);
nor U9348 (N_9348,N_5844,N_6348);
and U9349 (N_9349,N_5590,N_6828);
nor U9350 (N_9350,N_6884,N_6965);
nand U9351 (N_9351,N_7484,N_5917);
nor U9352 (N_9352,N_5840,N_5924);
or U9353 (N_9353,N_6894,N_6954);
nor U9354 (N_9354,N_5882,N_5192);
nor U9355 (N_9355,N_6051,N_5438);
or U9356 (N_9356,N_5021,N_5979);
and U9357 (N_9357,N_7015,N_5432);
or U9358 (N_9358,N_5598,N_6968);
nor U9359 (N_9359,N_7021,N_5527);
nor U9360 (N_9360,N_5727,N_6177);
nor U9361 (N_9361,N_7469,N_7498);
nand U9362 (N_9362,N_7488,N_7411);
nor U9363 (N_9363,N_7330,N_7217);
or U9364 (N_9364,N_7157,N_6644);
nand U9365 (N_9365,N_6620,N_7422);
nor U9366 (N_9366,N_7209,N_5948);
nand U9367 (N_9367,N_6297,N_5041);
or U9368 (N_9368,N_5138,N_6352);
or U9369 (N_9369,N_5570,N_5102);
nor U9370 (N_9370,N_7072,N_7171);
nor U9371 (N_9371,N_6241,N_7338);
nor U9372 (N_9372,N_6556,N_6539);
nand U9373 (N_9373,N_6416,N_7406);
or U9374 (N_9374,N_6938,N_5419);
and U9375 (N_9375,N_5354,N_6550);
and U9376 (N_9376,N_6684,N_5006);
nor U9377 (N_9377,N_5753,N_6983);
and U9378 (N_9378,N_7352,N_6465);
nand U9379 (N_9379,N_6463,N_6036);
nand U9380 (N_9380,N_5144,N_6951);
or U9381 (N_9381,N_5364,N_6239);
nor U9382 (N_9382,N_7044,N_5592);
nor U9383 (N_9383,N_7133,N_5025);
and U9384 (N_9384,N_5297,N_6596);
or U9385 (N_9385,N_5121,N_5123);
or U9386 (N_9386,N_6881,N_6358);
and U9387 (N_9387,N_6692,N_5021);
nand U9388 (N_9388,N_7340,N_6787);
nand U9389 (N_9389,N_6100,N_7431);
and U9390 (N_9390,N_5054,N_6149);
nand U9391 (N_9391,N_6408,N_5571);
and U9392 (N_9392,N_7312,N_6276);
nand U9393 (N_9393,N_6502,N_5091);
nand U9394 (N_9394,N_7256,N_6275);
nand U9395 (N_9395,N_6700,N_5756);
or U9396 (N_9396,N_5459,N_7148);
and U9397 (N_9397,N_5218,N_5406);
or U9398 (N_9398,N_5681,N_6673);
and U9399 (N_9399,N_6097,N_7494);
nand U9400 (N_9400,N_7340,N_5401);
nand U9401 (N_9401,N_5962,N_6388);
nand U9402 (N_9402,N_5639,N_5853);
nand U9403 (N_9403,N_6638,N_5234);
or U9404 (N_9404,N_6830,N_6723);
and U9405 (N_9405,N_5909,N_6292);
nor U9406 (N_9406,N_6195,N_5195);
and U9407 (N_9407,N_6427,N_5525);
nand U9408 (N_9408,N_7019,N_6361);
nor U9409 (N_9409,N_5798,N_5198);
nand U9410 (N_9410,N_6153,N_6097);
or U9411 (N_9411,N_7045,N_5401);
and U9412 (N_9412,N_6121,N_7458);
and U9413 (N_9413,N_5865,N_6802);
and U9414 (N_9414,N_5226,N_6766);
nor U9415 (N_9415,N_6480,N_6244);
nand U9416 (N_9416,N_5835,N_5617);
and U9417 (N_9417,N_7490,N_5486);
nor U9418 (N_9418,N_5086,N_5601);
nand U9419 (N_9419,N_5632,N_5045);
nor U9420 (N_9420,N_6878,N_6787);
nand U9421 (N_9421,N_5345,N_6058);
nor U9422 (N_9422,N_5300,N_6241);
or U9423 (N_9423,N_6537,N_5017);
nor U9424 (N_9424,N_5416,N_5156);
nand U9425 (N_9425,N_6657,N_5345);
and U9426 (N_9426,N_6564,N_5261);
nor U9427 (N_9427,N_6163,N_6008);
or U9428 (N_9428,N_5032,N_5678);
and U9429 (N_9429,N_6369,N_5502);
nor U9430 (N_9430,N_6598,N_5112);
or U9431 (N_9431,N_7123,N_7028);
nand U9432 (N_9432,N_6286,N_6096);
nor U9433 (N_9433,N_6708,N_6063);
and U9434 (N_9434,N_5071,N_6792);
or U9435 (N_9435,N_5187,N_6467);
nor U9436 (N_9436,N_5064,N_5553);
nor U9437 (N_9437,N_5323,N_5875);
or U9438 (N_9438,N_6225,N_5186);
and U9439 (N_9439,N_5843,N_5480);
nand U9440 (N_9440,N_5729,N_5680);
and U9441 (N_9441,N_6260,N_5397);
or U9442 (N_9442,N_7330,N_6298);
and U9443 (N_9443,N_5430,N_5930);
nor U9444 (N_9444,N_5446,N_7468);
nand U9445 (N_9445,N_7499,N_5535);
and U9446 (N_9446,N_5776,N_5133);
or U9447 (N_9447,N_5067,N_7257);
and U9448 (N_9448,N_5554,N_7319);
or U9449 (N_9449,N_5269,N_7198);
or U9450 (N_9450,N_5267,N_6014);
nor U9451 (N_9451,N_6082,N_5709);
and U9452 (N_9452,N_6129,N_5095);
and U9453 (N_9453,N_5263,N_6198);
nor U9454 (N_9454,N_5277,N_5045);
or U9455 (N_9455,N_5926,N_6973);
or U9456 (N_9456,N_7198,N_5391);
nor U9457 (N_9457,N_5088,N_6619);
nor U9458 (N_9458,N_6060,N_7164);
and U9459 (N_9459,N_6944,N_5381);
nand U9460 (N_9460,N_5980,N_5588);
nor U9461 (N_9461,N_6044,N_5429);
and U9462 (N_9462,N_6112,N_6717);
and U9463 (N_9463,N_5108,N_6417);
and U9464 (N_9464,N_6643,N_6216);
nand U9465 (N_9465,N_5318,N_6383);
and U9466 (N_9466,N_6126,N_6106);
nand U9467 (N_9467,N_6368,N_5439);
nor U9468 (N_9468,N_7416,N_6716);
nor U9469 (N_9469,N_6025,N_6778);
and U9470 (N_9470,N_5882,N_7323);
or U9471 (N_9471,N_6000,N_7100);
nor U9472 (N_9472,N_6011,N_5855);
and U9473 (N_9473,N_5891,N_5727);
nand U9474 (N_9474,N_6502,N_5357);
nor U9475 (N_9475,N_6269,N_6149);
nor U9476 (N_9476,N_5871,N_7297);
nor U9477 (N_9477,N_5597,N_6259);
and U9478 (N_9478,N_7076,N_6802);
nand U9479 (N_9479,N_5217,N_5875);
or U9480 (N_9480,N_6648,N_6432);
nor U9481 (N_9481,N_7045,N_5150);
nor U9482 (N_9482,N_6048,N_5237);
nand U9483 (N_9483,N_5769,N_5138);
and U9484 (N_9484,N_7484,N_6358);
and U9485 (N_9485,N_6516,N_5192);
nor U9486 (N_9486,N_6805,N_6220);
or U9487 (N_9487,N_7232,N_7243);
and U9488 (N_9488,N_6010,N_7408);
nor U9489 (N_9489,N_7377,N_6174);
nand U9490 (N_9490,N_5857,N_5476);
nor U9491 (N_9491,N_5874,N_6788);
nand U9492 (N_9492,N_6014,N_5600);
and U9493 (N_9493,N_6310,N_5228);
nor U9494 (N_9494,N_5939,N_6415);
and U9495 (N_9495,N_5884,N_6598);
and U9496 (N_9496,N_6618,N_7150);
and U9497 (N_9497,N_6415,N_5209);
and U9498 (N_9498,N_6015,N_6353);
nor U9499 (N_9499,N_6339,N_6783);
nor U9500 (N_9500,N_6390,N_7066);
nor U9501 (N_9501,N_6426,N_6987);
and U9502 (N_9502,N_7336,N_5333);
nand U9503 (N_9503,N_5225,N_6525);
or U9504 (N_9504,N_6015,N_5973);
nand U9505 (N_9505,N_6508,N_6339);
nand U9506 (N_9506,N_6664,N_7445);
nand U9507 (N_9507,N_7422,N_5488);
nand U9508 (N_9508,N_6595,N_5521);
and U9509 (N_9509,N_7227,N_6643);
or U9510 (N_9510,N_6132,N_5153);
nor U9511 (N_9511,N_5287,N_6827);
nor U9512 (N_9512,N_5890,N_5678);
and U9513 (N_9513,N_5011,N_6964);
nand U9514 (N_9514,N_5565,N_6896);
nor U9515 (N_9515,N_6556,N_5229);
and U9516 (N_9516,N_7389,N_7134);
nand U9517 (N_9517,N_5278,N_5214);
nand U9518 (N_9518,N_6375,N_7145);
or U9519 (N_9519,N_5268,N_6401);
and U9520 (N_9520,N_5907,N_7127);
nor U9521 (N_9521,N_6242,N_6381);
or U9522 (N_9522,N_6631,N_5898);
or U9523 (N_9523,N_6970,N_5940);
or U9524 (N_9524,N_5544,N_6834);
or U9525 (N_9525,N_5716,N_7216);
or U9526 (N_9526,N_5924,N_6164);
nand U9527 (N_9527,N_6570,N_6690);
nand U9528 (N_9528,N_6316,N_5712);
and U9529 (N_9529,N_5589,N_6457);
and U9530 (N_9530,N_6495,N_6697);
or U9531 (N_9531,N_7187,N_6694);
nand U9532 (N_9532,N_6964,N_5693);
or U9533 (N_9533,N_5619,N_7061);
or U9534 (N_9534,N_6168,N_6349);
xor U9535 (N_9535,N_7364,N_5886);
nand U9536 (N_9536,N_5073,N_7090);
nor U9537 (N_9537,N_5486,N_5817);
nand U9538 (N_9538,N_6810,N_5843);
and U9539 (N_9539,N_5251,N_6555);
nor U9540 (N_9540,N_6080,N_5945);
nor U9541 (N_9541,N_5773,N_7454);
and U9542 (N_9542,N_5513,N_5272);
and U9543 (N_9543,N_5334,N_7099);
and U9544 (N_9544,N_7493,N_7146);
nand U9545 (N_9545,N_5125,N_5245);
xnor U9546 (N_9546,N_5106,N_5557);
nand U9547 (N_9547,N_5136,N_6444);
nor U9548 (N_9548,N_5576,N_5364);
nand U9549 (N_9549,N_5263,N_6719);
or U9550 (N_9550,N_6840,N_6525);
and U9551 (N_9551,N_6760,N_7480);
nand U9552 (N_9552,N_5866,N_5604);
nand U9553 (N_9553,N_6083,N_7077);
nand U9554 (N_9554,N_6934,N_5062);
nand U9555 (N_9555,N_6968,N_6573);
nand U9556 (N_9556,N_6078,N_6350);
or U9557 (N_9557,N_7109,N_5859);
nand U9558 (N_9558,N_7206,N_5021);
or U9559 (N_9559,N_6421,N_6760);
nor U9560 (N_9560,N_5775,N_5492);
nor U9561 (N_9561,N_7161,N_6300);
nand U9562 (N_9562,N_5319,N_7477);
and U9563 (N_9563,N_5875,N_6925);
or U9564 (N_9564,N_5940,N_5340);
nand U9565 (N_9565,N_6575,N_5103);
nor U9566 (N_9566,N_5351,N_6561);
nand U9567 (N_9567,N_6713,N_6478);
or U9568 (N_9568,N_5561,N_7448);
nand U9569 (N_9569,N_6128,N_7412);
or U9570 (N_9570,N_6111,N_5022);
nand U9571 (N_9571,N_5496,N_6970);
or U9572 (N_9572,N_7117,N_7346);
and U9573 (N_9573,N_5043,N_6822);
nand U9574 (N_9574,N_5141,N_7145);
and U9575 (N_9575,N_5275,N_5192);
or U9576 (N_9576,N_7034,N_6655);
and U9577 (N_9577,N_6277,N_6321);
and U9578 (N_9578,N_7490,N_5288);
nand U9579 (N_9579,N_6402,N_5474);
or U9580 (N_9580,N_5358,N_5178);
nand U9581 (N_9581,N_5831,N_5333);
and U9582 (N_9582,N_6049,N_7365);
and U9583 (N_9583,N_7202,N_7285);
and U9584 (N_9584,N_6724,N_6210);
or U9585 (N_9585,N_5429,N_7296);
and U9586 (N_9586,N_6344,N_7156);
or U9587 (N_9587,N_7101,N_7447);
or U9588 (N_9588,N_5393,N_5294);
nor U9589 (N_9589,N_7026,N_6671);
and U9590 (N_9590,N_5523,N_6488);
nor U9591 (N_9591,N_6448,N_6083);
and U9592 (N_9592,N_5317,N_6274);
and U9593 (N_9593,N_6711,N_6428);
and U9594 (N_9594,N_7126,N_6225);
nand U9595 (N_9595,N_6238,N_7016);
or U9596 (N_9596,N_6271,N_5107);
nor U9597 (N_9597,N_5211,N_6334);
nand U9598 (N_9598,N_6021,N_5060);
or U9599 (N_9599,N_5726,N_5832);
and U9600 (N_9600,N_6208,N_6957);
and U9601 (N_9601,N_6033,N_6089);
nor U9602 (N_9602,N_5680,N_5461);
nand U9603 (N_9603,N_5102,N_7405);
and U9604 (N_9604,N_7036,N_6019);
nor U9605 (N_9605,N_6178,N_7307);
or U9606 (N_9606,N_5604,N_6107);
or U9607 (N_9607,N_5739,N_7298);
and U9608 (N_9608,N_7320,N_5363);
and U9609 (N_9609,N_7317,N_5238);
nand U9610 (N_9610,N_5521,N_7296);
and U9611 (N_9611,N_6882,N_5850);
or U9612 (N_9612,N_7057,N_7152);
or U9613 (N_9613,N_6977,N_7044);
or U9614 (N_9614,N_7135,N_5383);
nand U9615 (N_9615,N_5635,N_5370);
nand U9616 (N_9616,N_5238,N_6180);
nor U9617 (N_9617,N_6863,N_6412);
or U9618 (N_9618,N_5713,N_6317);
and U9619 (N_9619,N_6436,N_7013);
nor U9620 (N_9620,N_6581,N_6931);
nor U9621 (N_9621,N_7425,N_6782);
and U9622 (N_9622,N_7251,N_5709);
nand U9623 (N_9623,N_6042,N_7151);
and U9624 (N_9624,N_6178,N_5575);
and U9625 (N_9625,N_5630,N_6546);
or U9626 (N_9626,N_5871,N_6603);
nor U9627 (N_9627,N_6820,N_5510);
nand U9628 (N_9628,N_6856,N_6025);
and U9629 (N_9629,N_6552,N_6267);
or U9630 (N_9630,N_7161,N_6051);
or U9631 (N_9631,N_6098,N_5113);
nand U9632 (N_9632,N_5631,N_5017);
nand U9633 (N_9633,N_7010,N_5544);
and U9634 (N_9634,N_6912,N_6531);
and U9635 (N_9635,N_5610,N_7299);
and U9636 (N_9636,N_6473,N_5506);
or U9637 (N_9637,N_6390,N_5342);
or U9638 (N_9638,N_5657,N_7116);
nor U9639 (N_9639,N_5630,N_5861);
nand U9640 (N_9640,N_5143,N_6946);
nand U9641 (N_9641,N_6243,N_6664);
nor U9642 (N_9642,N_7205,N_5801);
and U9643 (N_9643,N_5096,N_5085);
nand U9644 (N_9644,N_7350,N_6662);
nand U9645 (N_9645,N_7349,N_7079);
nand U9646 (N_9646,N_6693,N_6758);
nand U9647 (N_9647,N_7230,N_5473);
nor U9648 (N_9648,N_5331,N_6981);
nor U9649 (N_9649,N_5035,N_6998);
nor U9650 (N_9650,N_7430,N_6049);
nor U9651 (N_9651,N_7470,N_5374);
nand U9652 (N_9652,N_5641,N_7127);
and U9653 (N_9653,N_6183,N_5037);
and U9654 (N_9654,N_5058,N_5190);
or U9655 (N_9655,N_5880,N_7430);
xor U9656 (N_9656,N_5510,N_7256);
nand U9657 (N_9657,N_7007,N_5861);
nand U9658 (N_9658,N_6351,N_6508);
nand U9659 (N_9659,N_6895,N_7075);
nand U9660 (N_9660,N_6674,N_5189);
or U9661 (N_9661,N_7435,N_6540);
nor U9662 (N_9662,N_6590,N_5073);
nor U9663 (N_9663,N_6250,N_7155);
nor U9664 (N_9664,N_7479,N_5876);
and U9665 (N_9665,N_6331,N_5852);
nor U9666 (N_9666,N_7040,N_6536);
or U9667 (N_9667,N_6737,N_5221);
or U9668 (N_9668,N_6507,N_7261);
nor U9669 (N_9669,N_5519,N_6696);
xnor U9670 (N_9670,N_6190,N_6387);
nand U9671 (N_9671,N_7426,N_5248);
nor U9672 (N_9672,N_7120,N_6102);
and U9673 (N_9673,N_7437,N_7045);
nand U9674 (N_9674,N_6038,N_5049);
or U9675 (N_9675,N_5552,N_7286);
nor U9676 (N_9676,N_6954,N_6730);
nand U9677 (N_9677,N_5957,N_5253);
nor U9678 (N_9678,N_6901,N_6050);
nand U9679 (N_9679,N_6783,N_5069);
or U9680 (N_9680,N_5847,N_5047);
or U9681 (N_9681,N_6896,N_7111);
and U9682 (N_9682,N_6093,N_6144);
or U9683 (N_9683,N_5052,N_5066);
nand U9684 (N_9684,N_5750,N_7168);
nor U9685 (N_9685,N_5733,N_5023);
nor U9686 (N_9686,N_5232,N_6214);
nor U9687 (N_9687,N_5740,N_5192);
and U9688 (N_9688,N_5088,N_6398);
nor U9689 (N_9689,N_6148,N_7282);
nand U9690 (N_9690,N_6111,N_7016);
nand U9691 (N_9691,N_6186,N_7433);
or U9692 (N_9692,N_6397,N_6411);
or U9693 (N_9693,N_5103,N_5532);
nor U9694 (N_9694,N_5165,N_6650);
nand U9695 (N_9695,N_6789,N_7448);
nor U9696 (N_9696,N_6925,N_5877);
and U9697 (N_9697,N_5413,N_6447);
nand U9698 (N_9698,N_6140,N_6652);
nor U9699 (N_9699,N_7049,N_5033);
nand U9700 (N_9700,N_5151,N_7297);
or U9701 (N_9701,N_6507,N_5499);
nor U9702 (N_9702,N_7465,N_6377);
nor U9703 (N_9703,N_6017,N_5174);
nand U9704 (N_9704,N_5207,N_6058);
nand U9705 (N_9705,N_5522,N_5888);
nand U9706 (N_9706,N_7452,N_6350);
and U9707 (N_9707,N_6545,N_6781);
nand U9708 (N_9708,N_7190,N_5733);
nand U9709 (N_9709,N_5580,N_6807);
nand U9710 (N_9710,N_7299,N_7493);
nor U9711 (N_9711,N_5847,N_7497);
xor U9712 (N_9712,N_5164,N_7430);
nand U9713 (N_9713,N_5547,N_7441);
and U9714 (N_9714,N_7369,N_5199);
nand U9715 (N_9715,N_5072,N_5261);
or U9716 (N_9716,N_6456,N_5673);
or U9717 (N_9717,N_6332,N_7376);
or U9718 (N_9718,N_7020,N_6090);
nor U9719 (N_9719,N_6600,N_6116);
or U9720 (N_9720,N_5734,N_5816);
nand U9721 (N_9721,N_6721,N_5644);
nand U9722 (N_9722,N_6575,N_6790);
xnor U9723 (N_9723,N_5362,N_5037);
or U9724 (N_9724,N_6357,N_5685);
xnor U9725 (N_9725,N_6998,N_5434);
and U9726 (N_9726,N_6776,N_6208);
nand U9727 (N_9727,N_6105,N_6298);
or U9728 (N_9728,N_6914,N_6880);
nand U9729 (N_9729,N_7172,N_5940);
nor U9730 (N_9730,N_6790,N_7104);
nand U9731 (N_9731,N_6493,N_7324);
or U9732 (N_9732,N_5309,N_6815);
and U9733 (N_9733,N_5655,N_6056);
or U9734 (N_9734,N_7470,N_5423);
nand U9735 (N_9735,N_5352,N_5853);
and U9736 (N_9736,N_6893,N_6569);
nor U9737 (N_9737,N_5863,N_6860);
and U9738 (N_9738,N_6377,N_5664);
nor U9739 (N_9739,N_6384,N_6931);
and U9740 (N_9740,N_7497,N_5466);
and U9741 (N_9741,N_7238,N_5446);
nand U9742 (N_9742,N_5190,N_6174);
and U9743 (N_9743,N_7377,N_7297);
or U9744 (N_9744,N_5612,N_7113);
nor U9745 (N_9745,N_5614,N_5618);
nand U9746 (N_9746,N_7304,N_5185);
nand U9747 (N_9747,N_5942,N_5725);
or U9748 (N_9748,N_5817,N_6102);
or U9749 (N_9749,N_5073,N_5025);
or U9750 (N_9750,N_5606,N_5209);
or U9751 (N_9751,N_5251,N_6046);
or U9752 (N_9752,N_6341,N_6902);
and U9753 (N_9753,N_5519,N_7111);
nor U9754 (N_9754,N_6100,N_5754);
nand U9755 (N_9755,N_6705,N_6915);
and U9756 (N_9756,N_7242,N_6397);
or U9757 (N_9757,N_6823,N_6881);
nor U9758 (N_9758,N_7239,N_5345);
nand U9759 (N_9759,N_6205,N_5498);
nor U9760 (N_9760,N_6513,N_5318);
and U9761 (N_9761,N_5428,N_6557);
nand U9762 (N_9762,N_5883,N_7238);
and U9763 (N_9763,N_5121,N_7389);
or U9764 (N_9764,N_6356,N_7434);
and U9765 (N_9765,N_7302,N_6790);
nand U9766 (N_9766,N_5813,N_5203);
or U9767 (N_9767,N_6338,N_5251);
and U9768 (N_9768,N_5219,N_6498);
nand U9769 (N_9769,N_6522,N_6734);
nor U9770 (N_9770,N_6632,N_6435);
or U9771 (N_9771,N_5330,N_6688);
and U9772 (N_9772,N_7398,N_6000);
nand U9773 (N_9773,N_5719,N_7331);
or U9774 (N_9774,N_7082,N_7027);
nor U9775 (N_9775,N_5060,N_5225);
or U9776 (N_9776,N_7312,N_5939);
and U9777 (N_9777,N_6721,N_6703);
or U9778 (N_9778,N_7241,N_7162);
or U9779 (N_9779,N_6580,N_7212);
or U9780 (N_9780,N_7468,N_6335);
nor U9781 (N_9781,N_6604,N_6974);
and U9782 (N_9782,N_5810,N_5767);
nor U9783 (N_9783,N_5155,N_7285);
nor U9784 (N_9784,N_5150,N_5900);
or U9785 (N_9785,N_6085,N_5141);
nor U9786 (N_9786,N_7115,N_6559);
nand U9787 (N_9787,N_7462,N_5560);
or U9788 (N_9788,N_6976,N_6829);
nor U9789 (N_9789,N_5186,N_6934);
or U9790 (N_9790,N_7428,N_5961);
nor U9791 (N_9791,N_5404,N_5233);
nor U9792 (N_9792,N_5797,N_5196);
and U9793 (N_9793,N_7080,N_5713);
xnor U9794 (N_9794,N_6290,N_7201);
or U9795 (N_9795,N_5673,N_5298);
nor U9796 (N_9796,N_7116,N_7249);
nand U9797 (N_9797,N_6508,N_6865);
or U9798 (N_9798,N_5512,N_5527);
nor U9799 (N_9799,N_5749,N_5421);
nor U9800 (N_9800,N_6550,N_5801);
or U9801 (N_9801,N_7495,N_7188);
or U9802 (N_9802,N_7077,N_5111);
or U9803 (N_9803,N_6628,N_5213);
and U9804 (N_9804,N_6235,N_5322);
nor U9805 (N_9805,N_5422,N_5775);
xor U9806 (N_9806,N_6340,N_7003);
nand U9807 (N_9807,N_7357,N_7042);
and U9808 (N_9808,N_6530,N_6168);
and U9809 (N_9809,N_6870,N_6906);
or U9810 (N_9810,N_6618,N_5355);
or U9811 (N_9811,N_5561,N_6970);
or U9812 (N_9812,N_6631,N_5836);
or U9813 (N_9813,N_5812,N_6809);
and U9814 (N_9814,N_6638,N_6031);
or U9815 (N_9815,N_5242,N_6581);
and U9816 (N_9816,N_6139,N_6787);
or U9817 (N_9817,N_7230,N_6308);
or U9818 (N_9818,N_5014,N_5349);
and U9819 (N_9819,N_7038,N_7298);
nor U9820 (N_9820,N_6150,N_5371);
nand U9821 (N_9821,N_6081,N_5799);
and U9822 (N_9822,N_7127,N_7022);
and U9823 (N_9823,N_6228,N_6548);
or U9824 (N_9824,N_6748,N_6783);
or U9825 (N_9825,N_7243,N_6778);
nand U9826 (N_9826,N_6021,N_6918);
nor U9827 (N_9827,N_7405,N_5429);
or U9828 (N_9828,N_7171,N_7350);
nand U9829 (N_9829,N_6593,N_7281);
nand U9830 (N_9830,N_7275,N_5482);
and U9831 (N_9831,N_6397,N_5077);
nand U9832 (N_9832,N_5951,N_7456);
or U9833 (N_9833,N_5719,N_7011);
nor U9834 (N_9834,N_6826,N_5662);
nand U9835 (N_9835,N_5157,N_6146);
nor U9836 (N_9836,N_6606,N_6275);
nor U9837 (N_9837,N_5494,N_7133);
nand U9838 (N_9838,N_7223,N_7323);
nand U9839 (N_9839,N_6421,N_5929);
nand U9840 (N_9840,N_5219,N_7316);
and U9841 (N_9841,N_7136,N_7240);
and U9842 (N_9842,N_7152,N_6202);
nand U9843 (N_9843,N_6916,N_5152);
or U9844 (N_9844,N_6375,N_6320);
nor U9845 (N_9845,N_6499,N_5290);
and U9846 (N_9846,N_5608,N_5105);
and U9847 (N_9847,N_7309,N_7498);
nand U9848 (N_9848,N_5200,N_5750);
nand U9849 (N_9849,N_5915,N_5044);
or U9850 (N_9850,N_5746,N_6702);
nor U9851 (N_9851,N_5074,N_6629);
nor U9852 (N_9852,N_6175,N_6406);
nand U9853 (N_9853,N_6883,N_6681);
xor U9854 (N_9854,N_6863,N_6229);
or U9855 (N_9855,N_6362,N_7088);
and U9856 (N_9856,N_6783,N_6900);
nand U9857 (N_9857,N_6164,N_7102);
or U9858 (N_9858,N_7481,N_7381);
nor U9859 (N_9859,N_5453,N_5630);
or U9860 (N_9860,N_6731,N_5189);
and U9861 (N_9861,N_5039,N_6334);
or U9862 (N_9862,N_6398,N_6025);
and U9863 (N_9863,N_7081,N_6398);
and U9864 (N_9864,N_6529,N_5383);
nand U9865 (N_9865,N_6934,N_7443);
nand U9866 (N_9866,N_6235,N_5041);
nand U9867 (N_9867,N_5776,N_5935);
or U9868 (N_9868,N_6978,N_6861);
nand U9869 (N_9869,N_5781,N_6658);
or U9870 (N_9870,N_5791,N_6687);
nor U9871 (N_9871,N_5392,N_5570);
and U9872 (N_9872,N_5173,N_5166);
nor U9873 (N_9873,N_6435,N_7257);
nand U9874 (N_9874,N_6051,N_6503);
or U9875 (N_9875,N_5433,N_6901);
nor U9876 (N_9876,N_6430,N_7116);
or U9877 (N_9877,N_5804,N_5403);
or U9878 (N_9878,N_6763,N_5987);
and U9879 (N_9879,N_6065,N_7143);
nor U9880 (N_9880,N_6266,N_7463);
or U9881 (N_9881,N_6700,N_5088);
nor U9882 (N_9882,N_5871,N_5108);
nor U9883 (N_9883,N_6662,N_6555);
nand U9884 (N_9884,N_5825,N_7269);
nand U9885 (N_9885,N_5053,N_5202);
and U9886 (N_9886,N_6186,N_7277);
nor U9887 (N_9887,N_5924,N_6101);
or U9888 (N_9888,N_6592,N_5659);
and U9889 (N_9889,N_5937,N_5559);
nand U9890 (N_9890,N_6168,N_6499);
nand U9891 (N_9891,N_6631,N_6947);
nand U9892 (N_9892,N_5622,N_5231);
nand U9893 (N_9893,N_7052,N_5199);
nor U9894 (N_9894,N_5696,N_6006);
or U9895 (N_9895,N_5141,N_6568);
and U9896 (N_9896,N_5835,N_5674);
or U9897 (N_9897,N_5733,N_7387);
or U9898 (N_9898,N_7164,N_7192);
and U9899 (N_9899,N_7156,N_7227);
nand U9900 (N_9900,N_5776,N_6666);
nand U9901 (N_9901,N_6344,N_6891);
nand U9902 (N_9902,N_5298,N_5536);
and U9903 (N_9903,N_7100,N_5423);
or U9904 (N_9904,N_7063,N_6419);
nor U9905 (N_9905,N_7008,N_6650);
or U9906 (N_9906,N_6710,N_6150);
nor U9907 (N_9907,N_5189,N_6622);
or U9908 (N_9908,N_7346,N_5939);
and U9909 (N_9909,N_5092,N_5722);
and U9910 (N_9910,N_5455,N_5177);
or U9911 (N_9911,N_5687,N_5253);
or U9912 (N_9912,N_5338,N_6970);
nor U9913 (N_9913,N_6425,N_7498);
or U9914 (N_9914,N_7470,N_5411);
or U9915 (N_9915,N_7091,N_7080);
or U9916 (N_9916,N_6974,N_5075);
or U9917 (N_9917,N_5873,N_6172);
or U9918 (N_9918,N_6630,N_6550);
nor U9919 (N_9919,N_5675,N_7499);
nand U9920 (N_9920,N_5707,N_5982);
or U9921 (N_9921,N_5810,N_5632);
nand U9922 (N_9922,N_6432,N_6800);
nor U9923 (N_9923,N_5484,N_6236);
nor U9924 (N_9924,N_7486,N_6375);
nor U9925 (N_9925,N_6529,N_5918);
nor U9926 (N_9926,N_7177,N_7173);
nand U9927 (N_9927,N_6511,N_6281);
or U9928 (N_9928,N_6915,N_5032);
or U9929 (N_9929,N_7427,N_7031);
nor U9930 (N_9930,N_5332,N_5415);
and U9931 (N_9931,N_6575,N_5887);
nor U9932 (N_9932,N_6777,N_5604);
and U9933 (N_9933,N_6694,N_5575);
nand U9934 (N_9934,N_5030,N_6991);
and U9935 (N_9935,N_5823,N_7124);
nor U9936 (N_9936,N_5096,N_5352);
and U9937 (N_9937,N_5213,N_5865);
or U9938 (N_9938,N_5171,N_7320);
or U9939 (N_9939,N_5823,N_7175);
nor U9940 (N_9940,N_5097,N_5734);
or U9941 (N_9941,N_7251,N_6397);
nor U9942 (N_9942,N_6898,N_7249);
and U9943 (N_9943,N_6600,N_6283);
and U9944 (N_9944,N_5900,N_6606);
nand U9945 (N_9945,N_6749,N_7270);
nor U9946 (N_9946,N_6906,N_5645);
nand U9947 (N_9947,N_6412,N_5063);
nand U9948 (N_9948,N_6896,N_6820);
nand U9949 (N_9949,N_6570,N_6278);
and U9950 (N_9950,N_6610,N_5983);
or U9951 (N_9951,N_6285,N_5828);
nor U9952 (N_9952,N_6084,N_6530);
or U9953 (N_9953,N_7426,N_5222);
or U9954 (N_9954,N_7124,N_5703);
nand U9955 (N_9955,N_6799,N_5030);
or U9956 (N_9956,N_5043,N_6857);
nand U9957 (N_9957,N_5209,N_6414);
nor U9958 (N_9958,N_7048,N_6886);
or U9959 (N_9959,N_6533,N_6917);
or U9960 (N_9960,N_7348,N_5213);
nor U9961 (N_9961,N_6340,N_6727);
and U9962 (N_9962,N_5906,N_7494);
or U9963 (N_9963,N_7107,N_7217);
nor U9964 (N_9964,N_5482,N_7078);
or U9965 (N_9965,N_7148,N_6572);
and U9966 (N_9966,N_7247,N_7147);
and U9967 (N_9967,N_6619,N_7119);
nand U9968 (N_9968,N_7088,N_5258);
nor U9969 (N_9969,N_5415,N_6327);
nand U9970 (N_9970,N_5361,N_5475);
and U9971 (N_9971,N_5799,N_6235);
and U9972 (N_9972,N_5977,N_6922);
and U9973 (N_9973,N_5853,N_6920);
and U9974 (N_9974,N_6189,N_6305);
nand U9975 (N_9975,N_6652,N_5271);
or U9976 (N_9976,N_5993,N_5301);
and U9977 (N_9977,N_5818,N_6853);
nor U9978 (N_9978,N_5017,N_7438);
nand U9979 (N_9979,N_7117,N_5501);
and U9980 (N_9980,N_5590,N_5628);
nor U9981 (N_9981,N_5899,N_6009);
or U9982 (N_9982,N_5427,N_6446);
and U9983 (N_9983,N_5113,N_6762);
and U9984 (N_9984,N_5722,N_6035);
or U9985 (N_9985,N_7475,N_5308);
and U9986 (N_9986,N_7033,N_7227);
nand U9987 (N_9987,N_6845,N_5399);
or U9988 (N_9988,N_7146,N_6192);
or U9989 (N_9989,N_7452,N_5451);
and U9990 (N_9990,N_5754,N_5160);
nor U9991 (N_9991,N_6290,N_7196);
nand U9992 (N_9992,N_7307,N_5881);
nand U9993 (N_9993,N_5110,N_6934);
nor U9994 (N_9994,N_7102,N_5419);
nand U9995 (N_9995,N_6662,N_6453);
and U9996 (N_9996,N_6040,N_6638);
nand U9997 (N_9997,N_5296,N_7456);
nand U9998 (N_9998,N_5056,N_6027);
or U9999 (N_9999,N_5908,N_7432);
and UO_0 (O_0,N_8462,N_7903);
or UO_1 (O_1,N_8161,N_7736);
or UO_2 (O_2,N_7884,N_8792);
nand UO_3 (O_3,N_9099,N_9273);
nand UO_4 (O_4,N_7857,N_8014);
nor UO_5 (O_5,N_9937,N_8882);
nor UO_6 (O_6,N_8076,N_9342);
or UO_7 (O_7,N_9927,N_7983);
nor UO_8 (O_8,N_8901,N_9746);
nor UO_9 (O_9,N_9195,N_7862);
xor UO_10 (O_10,N_9851,N_8690);
and UO_11 (O_11,N_9052,N_7721);
xor UO_12 (O_12,N_9874,N_9568);
nor UO_13 (O_13,N_9967,N_9347);
nor UO_14 (O_14,N_7569,N_9436);
nor UO_15 (O_15,N_9857,N_9644);
or UO_16 (O_16,N_9421,N_8750);
or UO_17 (O_17,N_8235,N_8022);
nor UO_18 (O_18,N_7770,N_7952);
and UO_19 (O_19,N_8639,N_7558);
and UO_20 (O_20,N_7960,N_9480);
and UO_21 (O_21,N_9507,N_8840);
or UO_22 (O_22,N_9727,N_9003);
nor UO_23 (O_23,N_9009,N_8715);
nand UO_24 (O_24,N_7723,N_8706);
and UO_25 (O_25,N_7518,N_8164);
nor UO_26 (O_26,N_7689,N_8024);
nor UO_27 (O_27,N_7729,N_8531);
nand UO_28 (O_28,N_9543,N_7988);
nand UO_29 (O_29,N_8342,N_9864);
and UO_30 (O_30,N_8511,N_8737);
nor UO_31 (O_31,N_9961,N_8598);
and UO_32 (O_32,N_8207,N_7882);
and UO_33 (O_33,N_7767,N_7662);
and UO_34 (O_34,N_9128,N_9056);
and UO_35 (O_35,N_8606,N_8732);
and UO_36 (O_36,N_8368,N_9910);
nor UO_37 (O_37,N_7758,N_8218);
nand UO_38 (O_38,N_9596,N_9968);
xor UO_39 (O_39,N_8234,N_7941);
nand UO_40 (O_40,N_9115,N_8058);
and UO_41 (O_41,N_8516,N_9267);
or UO_42 (O_42,N_9245,N_8809);
and UO_43 (O_43,N_9084,N_8766);
nand UO_44 (O_44,N_7938,N_8382);
or UO_45 (O_45,N_9385,N_8028);
or UO_46 (O_46,N_9881,N_8470);
or UO_47 (O_47,N_7820,N_8265);
nand UO_48 (O_48,N_7691,N_9379);
nand UO_49 (O_49,N_8284,N_9884);
and UO_50 (O_50,N_8093,N_8204);
or UO_51 (O_51,N_9808,N_8434);
or UO_52 (O_52,N_7972,N_8187);
or UO_53 (O_53,N_9268,N_8930);
xnor UO_54 (O_54,N_7711,N_9562);
or UO_55 (O_55,N_8186,N_8959);
nand UO_56 (O_56,N_8893,N_8729);
nor UO_57 (O_57,N_8733,N_9757);
nor UO_58 (O_58,N_8271,N_8576);
or UO_59 (O_59,N_7587,N_7567);
nand UO_60 (O_60,N_9139,N_7502);
and UO_61 (O_61,N_9711,N_8042);
and UO_62 (O_62,N_9623,N_8736);
nor UO_63 (O_63,N_8743,N_7744);
and UO_64 (O_64,N_8222,N_8769);
nor UO_65 (O_65,N_8900,N_7838);
nand UO_66 (O_66,N_7638,N_9241);
nand UO_67 (O_67,N_8712,N_8481);
nor UO_68 (O_68,N_9166,N_9984);
nand UO_69 (O_69,N_9331,N_8804);
or UO_70 (O_70,N_8634,N_7605);
nor UO_71 (O_71,N_8334,N_8723);
or UO_72 (O_72,N_8389,N_9903);
nor UO_73 (O_73,N_8077,N_7777);
nor UO_74 (O_74,N_8998,N_9057);
and UO_75 (O_75,N_8594,N_9229);
nor UO_76 (O_76,N_8274,N_8623);
nor UO_77 (O_77,N_8564,N_8622);
nand UO_78 (O_78,N_7986,N_9875);
nor UO_79 (O_79,N_8181,N_8902);
xor UO_80 (O_80,N_8927,N_8009);
or UO_81 (O_81,N_9610,N_8018);
nand UO_82 (O_82,N_9200,N_7977);
and UO_83 (O_83,N_7676,N_8475);
or UO_84 (O_84,N_9716,N_9947);
nor UO_85 (O_85,N_8864,N_9849);
nor UO_86 (O_86,N_9174,N_9791);
or UO_87 (O_87,N_9244,N_9476);
nor UO_88 (O_88,N_9395,N_9497);
nor UO_89 (O_89,N_8433,N_8524);
nand UO_90 (O_90,N_9451,N_9304);
nand UO_91 (O_91,N_9614,N_9521);
and UO_92 (O_92,N_7548,N_9813);
and UO_93 (O_93,N_7612,N_9856);
nand UO_94 (O_94,N_8986,N_7867);
xor UO_95 (O_95,N_9198,N_8242);
nand UO_96 (O_96,N_8169,N_8089);
nor UO_97 (O_97,N_8418,N_9558);
or UO_98 (O_98,N_8851,N_9809);
nand UO_99 (O_99,N_9738,N_9688);
nand UO_100 (O_100,N_7993,N_9122);
nor UO_101 (O_101,N_8638,N_9876);
nor UO_102 (O_102,N_9647,N_9587);
nor UO_103 (O_103,N_8507,N_7955);
nor UO_104 (O_104,N_9093,N_9569);
nor UO_105 (O_105,N_8289,N_8579);
and UO_106 (O_106,N_9165,N_8315);
and UO_107 (O_107,N_7851,N_9310);
and UO_108 (O_108,N_8086,N_7534);
or UO_109 (O_109,N_9210,N_8198);
nand UO_110 (O_110,N_8976,N_9770);
nor UO_111 (O_111,N_9134,N_8275);
nand UO_112 (O_112,N_8513,N_9088);
nand UO_113 (O_113,N_9905,N_7979);
nand UO_114 (O_114,N_7841,N_9613);
or UO_115 (O_115,N_9818,N_8735);
or UO_116 (O_116,N_9706,N_9433);
or UO_117 (O_117,N_8057,N_8149);
nand UO_118 (O_118,N_8728,N_9277);
or UO_119 (O_119,N_9110,N_8045);
nor UO_120 (O_120,N_7728,N_8779);
nand UO_121 (O_121,N_9887,N_8473);
or UO_122 (O_122,N_7812,N_7682);
and UO_123 (O_123,N_7763,N_9503);
nor UO_124 (O_124,N_9748,N_9296);
nor UO_125 (O_125,N_9519,N_9589);
and UO_126 (O_126,N_9042,N_8081);
and UO_127 (O_127,N_9760,N_9831);
or UO_128 (O_128,N_8810,N_9799);
nor UO_129 (O_129,N_7526,N_8548);
nand UO_130 (O_130,N_9798,N_9676);
nand UO_131 (O_131,N_8788,N_8938);
or UO_132 (O_132,N_9089,N_8359);
nand UO_133 (O_133,N_8801,N_7818);
and UO_134 (O_134,N_8694,N_7775);
or UO_135 (O_135,N_8569,N_8329);
and UO_136 (O_136,N_7814,N_9971);
and UO_137 (O_137,N_9917,N_7883);
and UO_138 (O_138,N_8353,N_9982);
or UO_139 (O_139,N_9812,N_9202);
or UO_140 (O_140,N_9130,N_9733);
or UO_141 (O_141,N_9516,N_7781);
nor UO_142 (O_142,N_8451,N_8378);
and UO_143 (O_143,N_7858,N_8328);
nor UO_144 (O_144,N_9540,N_9272);
nor UO_145 (O_145,N_8146,N_8410);
nand UO_146 (O_146,N_9499,N_9445);
or UO_147 (O_147,N_8912,N_7627);
and UO_148 (O_148,N_9450,N_9429);
or UO_149 (O_149,N_8923,N_8637);
and UO_150 (O_150,N_8709,N_8246);
or UO_151 (O_151,N_9280,N_9209);
and UO_152 (O_152,N_9566,N_8617);
or UO_153 (O_153,N_8904,N_9745);
nor UO_154 (O_154,N_9888,N_8270);
xnor UO_155 (O_155,N_8961,N_8859);
and UO_156 (O_156,N_9021,N_8727);
nor UO_157 (O_157,N_9619,N_8427);
nand UO_158 (O_158,N_7906,N_9140);
or UO_159 (O_159,N_8701,N_9156);
or UO_160 (O_160,N_8114,N_7732);
or UO_161 (O_161,N_9981,N_9144);
nand UO_162 (O_162,N_9010,N_9635);
nor UO_163 (O_163,N_8095,N_7875);
and UO_164 (O_164,N_7507,N_9742);
nand UO_165 (O_165,N_8425,N_7871);
and UO_166 (O_166,N_8600,N_9517);
and UO_167 (O_167,N_8768,N_8011);
and UO_168 (O_168,N_8957,N_9087);
nand UO_169 (O_169,N_9208,N_8170);
or UO_170 (O_170,N_9270,N_8488);
or UO_171 (O_171,N_7920,N_8110);
nand UO_172 (O_172,N_8316,N_9324);
nand UO_173 (O_173,N_9816,N_7512);
or UO_174 (O_174,N_8363,N_9292);
nand UO_175 (O_175,N_9825,N_8245);
and UO_176 (O_176,N_9150,N_9051);
and UO_177 (O_177,N_7800,N_9205);
nand UO_178 (O_178,N_7730,N_8978);
and UO_179 (O_179,N_7779,N_8082);
and UO_180 (O_180,N_8633,N_9348);
and UO_181 (O_181,N_7553,N_8442);
nor UO_182 (O_182,N_7821,N_8565);
and UO_183 (O_183,N_8400,N_7734);
nor UO_184 (O_184,N_7663,N_9253);
nand UO_185 (O_185,N_9625,N_9269);
nor UO_186 (O_186,N_9151,N_7590);
nor UO_187 (O_187,N_8458,N_8312);
nand UO_188 (O_188,N_9697,N_9882);
and UO_189 (O_189,N_8966,N_8763);
or UO_190 (O_190,N_9337,N_8260);
nand UO_191 (O_191,N_7674,N_9576);
or UO_192 (O_192,N_8604,N_7896);
and UO_193 (O_193,N_9175,N_9390);
nand UO_194 (O_194,N_8681,N_8361);
nor UO_195 (O_195,N_8950,N_8500);
nor UO_196 (O_196,N_9537,N_8483);
nand UO_197 (O_197,N_8940,N_9283);
nor UO_198 (O_198,N_7540,N_9452);
and UO_199 (O_199,N_7611,N_9242);
and UO_200 (O_200,N_9732,N_9854);
nor UO_201 (O_201,N_7551,N_7600);
nand UO_202 (O_202,N_9233,N_8339);
and UO_203 (O_203,N_8918,N_9877);
or UO_204 (O_204,N_9034,N_9621);
nand UO_205 (O_205,N_7580,N_9370);
or UO_206 (O_206,N_9701,N_9369);
nand UO_207 (O_207,N_9815,N_7788);
nand UO_208 (O_208,N_9050,N_9317);
xnor UO_209 (O_209,N_8281,N_8338);
nand UO_210 (O_210,N_8373,N_9496);
or UO_211 (O_211,N_9548,N_8999);
nand UO_212 (O_212,N_9758,N_8515);
nor UO_213 (O_213,N_9456,N_8408);
nor UO_214 (O_214,N_8443,N_7887);
nor UO_215 (O_215,N_9472,N_9731);
nor UO_216 (O_216,N_7704,N_9237);
or UO_217 (O_217,N_9408,N_8017);
and UO_218 (O_218,N_9194,N_8040);
or UO_219 (O_219,N_9800,N_8798);
and UO_220 (O_220,N_7660,N_9129);
or UO_221 (O_221,N_9495,N_9402);
or UO_222 (O_222,N_7618,N_8455);
nand UO_223 (O_223,N_7850,N_8630);
nor UO_224 (O_224,N_8835,N_9207);
or UO_225 (O_225,N_8941,N_8143);
nor UO_226 (O_226,N_9406,N_7520);
nor UO_227 (O_227,N_9931,N_7584);
nor UO_228 (O_228,N_9991,N_9158);
or UO_229 (O_229,N_8060,N_9249);
nand UO_230 (O_230,N_7668,N_7702);
nor UO_231 (O_231,N_8306,N_8535);
nor UO_232 (O_232,N_8725,N_7586);
nor UO_233 (O_233,N_8925,N_8330);
or UO_234 (O_234,N_8908,N_9639);
and UO_235 (O_235,N_8583,N_9899);
nor UO_236 (O_236,N_7630,N_8348);
and UO_237 (O_237,N_9817,N_9567);
nor UO_238 (O_238,N_7500,N_9303);
or UO_239 (O_239,N_9040,N_8273);
nor UO_240 (O_240,N_7523,N_8230);
and UO_241 (O_241,N_8787,N_8526);
and UO_242 (O_242,N_8296,N_7692);
or UO_243 (O_243,N_9399,N_8573);
nor UO_244 (O_244,N_9527,N_9065);
nor UO_245 (O_245,N_8943,N_8991);
or UO_246 (O_246,N_9988,N_9330);
or UO_247 (O_247,N_8030,N_9352);
nor UO_248 (O_248,N_7697,N_9414);
and UO_249 (O_249,N_9952,N_9775);
nand UO_250 (O_250,N_8984,N_8069);
and UO_251 (O_251,N_8173,N_8080);
and UO_252 (O_252,N_7560,N_9400);
nor UO_253 (O_253,N_9354,N_8720);
and UO_254 (O_254,N_9327,N_9943);
and UO_255 (O_255,N_8447,N_9845);
and UO_256 (O_256,N_9764,N_8213);
nand UO_257 (O_257,N_8355,N_8233);
nand UO_258 (O_258,N_7950,N_7591);
nand UO_259 (O_259,N_9391,N_9939);
and UO_260 (O_260,N_8770,N_9542);
or UO_261 (O_261,N_9940,N_8716);
xor UO_262 (O_262,N_8942,N_8759);
and UO_263 (O_263,N_8752,N_9538);
and UO_264 (O_264,N_8783,N_9046);
nand UO_265 (O_265,N_8003,N_9434);
or UO_266 (O_266,N_7637,N_9013);
and UO_267 (O_267,N_8160,N_7672);
nand UO_268 (O_268,N_9178,N_9419);
nand UO_269 (O_269,N_9344,N_7823);
nand UO_270 (O_270,N_9058,N_8512);
nor UO_271 (O_271,N_9524,N_9275);
nand UO_272 (O_272,N_9989,N_8200);
and UO_273 (O_273,N_9980,N_8349);
and UO_274 (O_274,N_8292,N_9918);
and UO_275 (O_275,N_9228,N_8054);
and UO_276 (O_276,N_8297,N_8140);
and UO_277 (O_277,N_9231,N_9855);
and UO_278 (O_278,N_7588,N_9141);
and UO_279 (O_279,N_9047,N_8553);
and UO_280 (O_280,N_7984,N_7936);
nand UO_281 (O_281,N_8175,N_9031);
nand UO_282 (O_282,N_9541,N_9563);
xnor UO_283 (O_283,N_8889,N_8440);
nand UO_284 (O_284,N_9776,N_9997);
nor UO_285 (O_285,N_7846,N_7870);
nor UO_286 (O_286,N_9622,N_7865);
or UO_287 (O_287,N_9907,N_8877);
nand UO_288 (O_288,N_8407,N_9276);
and UO_289 (O_289,N_9546,N_9750);
nand UO_290 (O_290,N_8791,N_9708);
nand UO_291 (O_291,N_8038,N_8112);
and UO_292 (O_292,N_9753,N_8130);
or UO_293 (O_293,N_7552,N_8257);
nand UO_294 (O_294,N_8672,N_9754);
and UO_295 (O_295,N_9819,N_9023);
nor UO_296 (O_296,N_7978,N_8308);
and UO_297 (O_297,N_9838,N_8561);
nor UO_298 (O_298,N_9502,N_9357);
and UO_299 (O_299,N_9384,N_9301);
nor UO_300 (O_300,N_8087,N_9858);
nand UO_301 (O_301,N_9983,N_7546);
or UO_302 (O_302,N_9630,N_9409);
nor UO_303 (O_303,N_8421,N_7621);
and UO_304 (O_304,N_8761,N_9343);
and UO_305 (O_305,N_8029,N_7532);
nor UO_306 (O_306,N_9702,N_9609);
and UO_307 (O_307,N_7976,N_8746);
nand UO_308 (O_308,N_9498,N_7954);
and UO_309 (O_309,N_7886,N_9972);
nor UO_310 (O_310,N_8674,N_7749);
nor UO_311 (O_311,N_8873,N_9945);
or UO_312 (O_312,N_8300,N_9137);
nor UO_313 (O_313,N_8241,N_7971);
or UO_314 (O_314,N_7571,N_9778);
or UO_315 (O_315,N_8201,N_8294);
nand UO_316 (O_316,N_7733,N_7636);
or UO_317 (O_317,N_9740,N_8466);
and UO_318 (O_318,N_7869,N_9650);
or UO_319 (O_319,N_7908,N_7650);
nor UO_320 (O_320,N_8336,N_8302);
and UO_321 (O_321,N_9618,N_8664);
nor UO_322 (O_322,N_9119,N_8874);
and UO_323 (O_323,N_8062,N_7911);
or UO_324 (O_324,N_8523,N_7610);
or UO_325 (O_325,N_8879,N_7828);
nand UO_326 (O_326,N_9802,N_9728);
nand UO_327 (O_327,N_9915,N_9801);
nor UO_328 (O_328,N_7687,N_8663);
nor UO_329 (O_329,N_8493,N_8747);
nor UO_330 (O_330,N_9019,N_8960);
or UO_331 (O_331,N_9147,N_9374);
or UO_332 (O_332,N_9360,N_7585);
nor UO_333 (O_333,N_8267,N_8128);
nand UO_334 (O_334,N_8963,N_8650);
and UO_335 (O_335,N_9975,N_8450);
nor UO_336 (O_336,N_8730,N_7918);
and UO_337 (O_337,N_9167,N_9190);
or UO_338 (O_338,N_9594,N_9687);
or UO_339 (O_339,N_8365,N_8215);
xnor UO_340 (O_340,N_8061,N_9302);
xnor UO_341 (O_341,N_9788,N_7774);
nor UO_342 (O_342,N_8574,N_8394);
nand UO_343 (O_343,N_8980,N_9001);
and UO_344 (O_344,N_7998,N_9085);
and UO_345 (O_345,N_8608,N_9216);
and UO_346 (O_346,N_9413,N_8206);
nand UO_347 (O_347,N_7557,N_9365);
nand UO_348 (O_348,N_7945,N_8482);
nand UO_349 (O_349,N_8449,N_8092);
nand UO_350 (O_350,N_7959,N_8805);
and UO_351 (O_351,N_7745,N_8514);
and UO_352 (O_352,N_8745,N_8479);
nand UO_353 (O_353,N_8262,N_7652);
or UO_354 (O_354,N_7822,N_7522);
or UO_355 (O_355,N_9912,N_9787);
or UO_356 (O_356,N_8367,N_8148);
nor UO_357 (O_357,N_9323,N_8607);
nor UO_358 (O_358,N_9512,N_9934);
nor UO_359 (O_359,N_8700,N_8007);
nor UO_360 (O_360,N_7686,N_9847);
nand UO_361 (O_361,N_7608,N_9559);
nor UO_362 (O_362,N_9694,N_8417);
nand UO_363 (O_363,N_8891,N_8609);
nor UO_364 (O_364,N_8824,N_8718);
nand UO_365 (O_365,N_8452,N_8865);
nor UO_366 (O_366,N_9112,N_7695);
nor UO_367 (O_367,N_9018,N_9116);
and UO_368 (O_368,N_8456,N_8955);
nor UO_369 (O_369,N_8020,N_7815);
nand UO_370 (O_370,N_8166,N_9326);
and UO_371 (O_371,N_9284,N_7521);
and UO_372 (O_372,N_8127,N_7835);
nand UO_373 (O_373,N_8277,N_9904);
nand UO_374 (O_374,N_8554,N_7578);
and UO_375 (O_375,N_8176,N_9785);
or UO_376 (O_376,N_7773,N_7914);
and UO_377 (O_377,N_9552,N_8832);
nor UO_378 (O_378,N_8897,N_9295);
nand UO_379 (O_379,N_9640,N_7963);
and UO_380 (O_380,N_8678,N_8845);
nand UO_381 (O_381,N_8108,N_8320);
and UO_382 (O_382,N_9938,N_8740);
nor UO_383 (O_383,N_8282,N_9059);
and UO_384 (O_384,N_7910,N_7659);
nand UO_385 (O_385,N_8705,N_9328);
or UO_386 (O_386,N_9107,N_9751);
nand UO_387 (O_387,N_8340,N_7826);
nor UO_388 (O_388,N_8614,N_8734);
or UO_389 (O_389,N_8046,N_7949);
nor UO_390 (O_390,N_8540,N_8100);
or UO_391 (O_391,N_7836,N_8806);
or UO_392 (O_392,N_8974,N_9773);
or UO_393 (O_393,N_7975,N_8304);
nor UO_394 (O_394,N_8887,N_8439);
or UO_395 (O_395,N_8863,N_7525);
nand UO_396 (O_396,N_9090,N_7603);
and UO_397 (O_397,N_8151,N_9699);
or UO_398 (O_398,N_9029,N_8590);
and UO_399 (O_399,N_8305,N_8875);
and UO_400 (O_400,N_8670,N_9339);
nor UO_401 (O_401,N_7593,N_8357);
or UO_402 (O_402,N_9243,N_8319);
or UO_403 (O_403,N_7604,N_7802);
or UO_404 (O_404,N_8362,N_7505);
or UO_405 (O_405,N_9737,N_9823);
nand UO_406 (O_406,N_7899,N_8065);
or UO_407 (O_407,N_7542,N_9712);
or UO_408 (O_408,N_9325,N_8613);
or UO_409 (O_409,N_9747,N_7684);
nor UO_410 (O_410,N_9525,N_7916);
and UO_411 (O_411,N_9710,N_9215);
nand UO_412 (O_412,N_8921,N_9836);
and UO_413 (O_413,N_9841,N_9157);
and UO_414 (O_414,N_9765,N_8929);
and UO_415 (O_415,N_8915,N_9582);
and UO_416 (O_416,N_8254,N_9677);
nand UO_417 (O_417,N_9792,N_9772);
and UO_418 (O_418,N_8838,N_9033);
nand UO_419 (O_419,N_9951,N_8621);
and UO_420 (O_420,N_9062,N_9479);
nor UO_421 (O_421,N_8432,N_9182);
nor UO_422 (O_422,N_9911,N_8861);
and UO_423 (O_423,N_9306,N_7933);
nor UO_424 (O_424,N_8188,N_9936);
nor UO_425 (O_425,N_7649,N_7602);
and UO_426 (O_426,N_9769,N_9811);
and UO_427 (O_427,N_9236,N_7880);
nand UO_428 (O_428,N_8822,N_9477);
and UO_429 (O_429,N_8404,N_8880);
nor UO_430 (O_430,N_7698,N_9045);
or UO_431 (O_431,N_7693,N_8220);
nor UO_432 (O_432,N_9183,N_9196);
or UO_433 (O_433,N_8125,N_7996);
or UO_434 (O_434,N_7623,N_7819);
and UO_435 (O_435,N_9070,N_7844);
nor UO_436 (O_436,N_9455,N_8631);
or UO_437 (O_437,N_8209,N_9474);
or UO_438 (O_438,N_7705,N_9313);
and UO_439 (O_439,N_9960,N_8947);
or UO_440 (O_440,N_7619,N_8474);
and UO_441 (O_441,N_9724,N_9532);
nand UO_442 (O_442,N_8210,N_7696);
and UO_443 (O_443,N_8559,N_9591);
xor UO_444 (O_444,N_8800,N_7940);
and UO_445 (O_445,N_7997,N_7853);
and UO_446 (O_446,N_8468,N_7973);
or UO_447 (O_447,N_8934,N_8172);
and UO_448 (O_448,N_8385,N_7508);
or UO_449 (O_449,N_8506,N_8505);
nor UO_450 (O_450,N_9382,N_9553);
or UO_451 (O_451,N_9660,N_8096);
and UO_452 (O_452,N_8666,N_8495);
and UO_453 (O_453,N_9528,N_7943);
or UO_454 (O_454,N_7824,N_8909);
nor UO_455 (O_455,N_9493,N_9916);
or UO_456 (O_456,N_8437,N_9213);
or UO_457 (O_457,N_9255,N_9104);
or UO_458 (O_458,N_7985,N_8646);
or UO_459 (O_459,N_8123,N_8883);
nor UO_460 (O_460,N_9970,N_9136);
nor UO_461 (O_461,N_7524,N_9766);
nand UO_462 (O_462,N_8118,N_8823);
nor UO_463 (O_463,N_8120,N_7861);
and UO_464 (O_464,N_9868,N_7632);
or UO_465 (O_465,N_7948,N_8147);
or UO_466 (O_466,N_9920,N_8985);
nor UO_467 (O_467,N_9017,N_7568);
and UO_468 (O_468,N_9022,N_7885);
and UO_469 (O_469,N_9696,N_7554);
or UO_470 (O_470,N_7889,N_9626);
and UO_471 (O_471,N_9080,N_8104);
nand UO_472 (O_472,N_7995,N_9431);
and UO_473 (O_473,N_9892,N_9319);
nand UO_474 (O_474,N_8826,N_8344);
and UO_475 (O_475,N_9248,N_9844);
or UO_476 (O_476,N_8472,N_9771);
and UO_477 (O_477,N_7566,N_9491);
nand UO_478 (O_478,N_8406,N_8541);
and UO_479 (O_479,N_9329,N_8677);
or UO_480 (O_480,N_9185,N_8388);
nand UO_481 (O_481,N_8227,N_9529);
and UO_482 (O_482,N_8828,N_7628);
or UO_483 (O_483,N_8064,N_8714);
xor UO_484 (O_484,N_9297,N_9860);
nor UO_485 (O_485,N_9761,N_7629);
or UO_486 (O_486,N_7708,N_7656);
or UO_487 (O_487,N_9473,N_9469);
and UO_488 (O_488,N_7783,N_8871);
and UO_489 (O_489,N_8726,N_8221);
nor UO_490 (O_490,N_9393,N_8989);
nand UO_491 (O_491,N_8847,N_7596);
nor UO_492 (O_492,N_8758,N_8286);
and UO_493 (O_493,N_8272,N_8298);
or UO_494 (O_494,N_8471,N_7913);
or UO_495 (O_495,N_8928,N_9834);
and UO_496 (O_496,N_7719,N_8549);
nor UO_497 (O_497,N_9651,N_8223);
nand UO_498 (O_498,N_9173,N_9336);
and UO_499 (O_499,N_8786,N_7595);
and UO_500 (O_500,N_8454,N_8981);
or UO_501 (O_501,N_7657,N_8131);
and UO_502 (O_502,N_9935,N_7701);
or UO_503 (O_503,N_9102,N_9779);
nor UO_504 (O_504,N_8926,N_9079);
and UO_505 (O_505,N_8906,N_8337);
nor UO_506 (O_506,N_8776,N_8580);
nor UO_507 (O_507,N_9279,N_8441);
nand UO_508 (O_508,N_7925,N_8962);
and UO_509 (O_509,N_9986,N_7527);
and UO_510 (O_510,N_9902,N_9925);
and UO_511 (O_511,N_8232,N_9883);
or UO_512 (O_512,N_8424,N_9155);
nor UO_513 (O_513,N_9189,N_8135);
and UO_514 (O_514,N_9867,N_8136);
and UO_515 (O_515,N_7699,N_8692);
nand UO_516 (O_516,N_7756,N_8852);
or UO_517 (O_517,N_7785,N_9486);
and UO_518 (O_518,N_9420,N_8510);
and UO_519 (O_519,N_8675,N_8560);
nor UO_520 (O_520,N_8476,N_9933);
or UO_521 (O_521,N_9488,N_8066);
or UO_522 (O_522,N_9259,N_9634);
or UO_523 (O_523,N_9736,N_8612);
nor UO_524 (O_524,N_8465,N_7641);
nor UO_525 (O_525,N_9544,N_8099);
and UO_526 (O_526,N_8317,N_7556);
or UO_527 (O_527,N_9187,N_8171);
or UO_528 (O_528,N_9002,N_9741);
or UO_529 (O_529,N_9394,N_9305);
nand UO_530 (O_530,N_8008,N_7535);
and UO_531 (O_531,N_9163,N_8333);
and UO_532 (O_532,N_7811,N_9036);
nor UO_533 (O_533,N_9759,N_9969);
nand UO_534 (O_534,N_8687,N_8738);
and UO_535 (O_535,N_8521,N_9181);
nor UO_536 (O_536,N_8619,N_9929);
or UO_537 (O_537,N_9028,N_8689);
nor UO_538 (O_538,N_8830,N_9274);
nand UO_539 (O_539,N_8982,N_7747);
nand UO_540 (O_540,N_8191,N_9246);
and UO_541 (O_541,N_9432,N_7864);
nand UO_542 (O_542,N_9359,N_9153);
or UO_543 (O_543,N_9581,N_9777);
or UO_544 (O_544,N_9695,N_8152);
and UO_545 (O_545,N_9879,N_8652);
xnor UO_546 (O_546,N_7961,N_9999);
or UO_547 (O_547,N_8428,N_9992);
or UO_548 (O_548,N_8821,N_8053);
nor UO_549 (O_549,N_7583,N_8844);
nand UO_550 (O_550,N_7877,N_8402);
and UO_551 (O_551,N_8343,N_8537);
nor UO_552 (O_552,N_9232,N_8990);
and UO_553 (O_553,N_7965,N_8074);
or UO_554 (O_554,N_7562,N_9846);
nor UO_555 (O_555,N_9422,N_8203);
nor UO_556 (O_556,N_9962,N_9224);
and UO_557 (O_557,N_7873,N_9332);
nor UO_558 (O_558,N_8935,N_9922);
and UO_559 (O_559,N_7968,N_8250);
nand UO_560 (O_560,N_8291,N_9333);
and UO_561 (O_561,N_8183,N_9781);
or UO_562 (O_562,N_9570,N_9286);
nor UO_563 (O_563,N_8953,N_7561);
and UO_564 (O_564,N_9355,N_9689);
nor UO_565 (O_565,N_7804,N_9160);
and UO_566 (O_566,N_8698,N_7926);
nand UO_567 (O_567,N_7991,N_8279);
nand UO_568 (O_568,N_8647,N_8139);
nor UO_569 (O_569,N_9315,N_7924);
nand UO_570 (O_570,N_8979,N_9238);
nand UO_571 (O_571,N_9900,N_8858);
and UO_572 (O_572,N_8036,N_8811);
nand UO_573 (O_573,N_7670,N_8952);
and UO_574 (O_574,N_9501,N_7741);
or UO_575 (O_575,N_9560,N_9222);
and UO_576 (O_576,N_8448,N_7958);
or UO_577 (O_577,N_9392,N_9535);
and UO_578 (O_578,N_8413,N_8395);
nor UO_579 (O_579,N_7653,N_8094);
and UO_580 (O_580,N_8542,N_9478);
or UO_581 (O_581,N_7690,N_9557);
nand UO_582 (O_582,N_7654,N_9835);
nor UO_583 (O_583,N_8760,N_9271);
or UO_584 (O_584,N_8657,N_9842);
nand UO_585 (O_585,N_7712,N_8293);
nor UO_586 (O_586,N_9605,N_7541);
or UO_587 (O_587,N_9014,N_8582);
nor UO_588 (O_588,N_9523,N_8593);
and UO_589 (O_589,N_9954,N_9471);
and UO_590 (O_590,N_8295,N_9005);
nor UO_591 (O_591,N_8419,N_9744);
nand UO_592 (O_592,N_7727,N_9261);
or UO_593 (O_593,N_9449,N_9025);
and UO_594 (O_594,N_9631,N_8162);
and UO_595 (O_595,N_8544,N_9941);
nand UO_596 (O_596,N_8816,N_9448);
and UO_597 (O_597,N_8556,N_8144);
nor UO_598 (O_598,N_8263,N_8494);
or UO_599 (O_599,N_8551,N_9511);
nand UO_600 (O_600,N_7651,N_9703);
nand UO_601 (O_601,N_9597,N_7805);
and UO_602 (O_602,N_9361,N_9906);
or UO_603 (O_603,N_8174,N_7620);
nor UO_604 (O_604,N_8645,N_9247);
and UO_605 (O_605,N_8749,N_9797);
nand UO_606 (O_606,N_8679,N_9211);
or UO_607 (O_607,N_9515,N_9837);
or UO_608 (O_608,N_8850,N_7946);
or UO_609 (O_609,N_9611,N_7707);
nand UO_610 (O_610,N_8754,N_8596);
nor UO_611 (O_611,N_7716,N_9805);
or UO_612 (O_612,N_8285,N_9561);
nand UO_613 (O_613,N_8477,N_9913);
nand UO_614 (O_614,N_8919,N_8004);
nand UO_615 (O_615,N_8686,N_8973);
and UO_616 (O_616,N_9092,N_9586);
or UO_617 (O_617,N_9682,N_9679);
and UO_618 (O_618,N_9607,N_8155);
or UO_619 (O_619,N_8485,N_8228);
nor UO_620 (O_620,N_9668,N_7813);
nand UO_621 (O_621,N_8971,N_9681);
nand UO_622 (O_622,N_8327,N_8031);
nor UO_623 (O_623,N_8669,N_8802);
and UO_624 (O_624,N_8356,N_9024);
nand UO_625 (O_625,N_8892,N_9948);
nor UO_626 (O_626,N_7776,N_8696);
nor UO_627 (O_627,N_8519,N_9076);
xnor UO_628 (O_628,N_7685,N_8266);
and UO_629 (O_629,N_7762,N_8192);
nand UO_630 (O_630,N_8499,N_9467);
nor UO_631 (O_631,N_7513,N_8438);
and UO_632 (O_632,N_9633,N_9974);
nor UO_633 (O_633,N_7793,N_9852);
nand UO_634 (O_634,N_7759,N_9299);
nor UO_635 (O_635,N_9755,N_7982);
nand UO_636 (O_636,N_8489,N_9894);
and UO_637 (O_637,N_9671,N_9234);
and UO_638 (O_638,N_9719,N_8585);
or UO_639 (O_639,N_7563,N_7750);
and UO_640 (O_640,N_7607,N_9990);
nor UO_641 (O_641,N_9015,N_8380);
and UO_642 (O_642,N_9850,N_7766);
nor UO_643 (O_643,N_7932,N_9086);
nand UO_644 (O_644,N_8050,N_7791);
nor UO_645 (O_645,N_8314,N_9113);
nor UO_646 (O_646,N_7859,N_9097);
and UO_647 (O_647,N_7742,N_7509);
and UO_648 (O_648,N_8016,N_8211);
and UO_649 (O_649,N_8193,N_9179);
nor UO_650 (O_650,N_7953,N_8951);
nand UO_651 (O_651,N_9843,N_8924);
and UO_652 (O_652,N_8497,N_9726);
nand UO_653 (O_653,N_9520,N_8097);
and UO_654 (O_654,N_7909,N_9389);
or UO_655 (O_655,N_8808,N_8185);
and UO_656 (O_656,N_7631,N_8253);
nand UO_657 (O_657,N_8570,N_8577);
nor UO_658 (O_658,N_9341,N_9599);
nor UO_659 (O_659,N_9683,N_7739);
and UO_660 (O_660,N_9547,N_8673);
nor UO_661 (O_661,N_8849,N_8422);
nand UO_662 (O_662,N_9522,N_8699);
nand UO_663 (O_663,N_9729,N_8435);
and UO_664 (O_664,N_9898,N_9412);
nor UO_665 (O_665,N_9822,N_9756);
and UO_666 (O_666,N_9308,N_7680);
or UO_667 (O_667,N_7679,N_8522);
and UO_668 (O_668,N_9206,N_8572);
or UO_669 (O_669,N_7967,N_7570);
nor UO_670 (O_670,N_7888,N_9862);
and UO_671 (O_671,N_9461,N_8001);
xnor UO_672 (O_672,N_9896,N_7669);
or UO_673 (O_673,N_7942,N_9309);
and UO_674 (O_674,N_8771,N_7917);
nand UO_675 (O_675,N_9578,N_7825);
and UO_676 (O_676,N_9509,N_8997);
nand UO_677 (O_677,N_9592,N_7832);
nor UO_678 (O_678,N_9993,N_9201);
nor UO_679 (O_679,N_8529,N_8085);
nor UO_680 (O_680,N_8231,N_9583);
or UO_681 (O_681,N_8248,N_8068);
or UO_682 (O_682,N_7878,N_9351);
nand UO_683 (O_683,N_9571,N_8857);
nand UO_684 (O_684,N_9585,N_9264);
and UO_685 (O_685,N_9680,N_8545);
nand UO_686 (O_686,N_9998,N_8178);
or UO_687 (O_687,N_9949,N_8225);
nand UO_688 (O_688,N_8122,N_9869);
and UO_689 (O_689,N_7989,N_7681);
or UO_690 (O_690,N_9666,N_7987);
or UO_691 (O_691,N_9440,N_9789);
nand UO_692 (O_692,N_8954,N_8351);
or UO_693 (O_693,N_9691,N_8629);
nand UO_694 (O_694,N_9437,N_8133);
xnor UO_695 (O_695,N_8731,N_8525);
or UO_696 (O_696,N_8492,N_9663);
or UO_697 (O_697,N_8051,N_7752);
and UO_698 (O_698,N_9577,N_9117);
nor UO_699 (O_699,N_8091,N_8399);
nand UO_700 (O_700,N_9055,N_8083);
and UO_701 (O_701,N_8199,N_9262);
nor UO_702 (O_702,N_9530,N_8557);
or UO_703 (O_703,N_9453,N_9749);
nand UO_704 (O_704,N_9987,N_8364);
or UO_705 (O_705,N_8948,N_8970);
and UO_706 (O_706,N_8431,N_7848);
nand UO_707 (O_707,N_9794,N_9909);
nand UO_708 (O_708,N_9282,N_8599);
and UO_709 (O_709,N_9793,N_9958);
nor UO_710 (O_710,N_8323,N_9533);
xor UO_711 (O_711,N_9642,N_8555);
nand UO_712 (O_712,N_7661,N_8387);
or UO_713 (O_713,N_9152,N_9398);
nor UO_714 (O_714,N_8581,N_9020);
or UO_715 (O_715,N_9774,N_8026);
and UO_716 (O_716,N_8781,N_7688);
nand UO_717 (O_717,N_8744,N_9314);
nor UO_718 (O_718,N_7529,N_9686);
and UO_719 (O_719,N_9481,N_9700);
or UO_720 (O_720,N_7845,N_9979);
nand UO_721 (O_721,N_8134,N_8911);
or UO_722 (O_722,N_9848,N_7829);
or UO_723 (O_723,N_7648,N_9054);
nand UO_724 (O_724,N_8167,N_7514);
and UO_725 (O_725,N_9725,N_8719);
nand UO_726 (O_726,N_8992,N_8785);
and UO_727 (O_727,N_8643,N_9996);
nor UO_728 (O_728,N_9346,N_7757);
or UO_729 (O_729,N_8707,N_9871);
nand UO_730 (O_730,N_9604,N_8655);
and UO_731 (O_731,N_8168,N_7582);
nor UO_732 (O_732,N_9485,N_8710);
nand UO_733 (O_733,N_8189,N_7720);
nor UO_734 (O_734,N_9072,N_9923);
or UO_735 (O_735,N_9784,N_9281);
nand UO_736 (O_736,N_9069,N_8249);
nand UO_737 (O_737,N_9565,N_8774);
nor UO_738 (O_738,N_8420,N_7852);
or UO_739 (O_739,N_9752,N_9489);
and UO_740 (O_740,N_9397,N_8722);
or UO_741 (O_741,N_7606,N_8480);
nor UO_742 (O_742,N_7703,N_9221);
or UO_743 (O_743,N_9180,N_8753);
nor UO_744 (O_744,N_7706,N_7576);
and UO_745 (O_745,N_9470,N_8177);
nor UO_746 (O_746,N_7544,N_9767);
nor UO_747 (O_747,N_8803,N_7579);
or UO_748 (O_748,N_9227,N_8163);
or UO_749 (O_749,N_8405,N_9298);
nor UO_750 (O_750,N_8287,N_8243);
and UO_751 (O_751,N_7574,N_9803);
and UO_752 (O_752,N_8142,N_8377);
or UO_753 (O_753,N_9891,N_8695);
nor UO_754 (O_754,N_7622,N_8866);
and UO_755 (O_755,N_9007,N_8661);
nor UO_756 (O_756,N_7503,N_7683);
or UO_757 (O_757,N_7992,N_9114);
nand UO_758 (O_758,N_9721,N_9575);
nand UO_759 (O_759,N_8756,N_7782);
nand UO_760 (O_760,N_9338,N_8656);
or UO_761 (O_761,N_8777,N_9465);
or UO_762 (O_762,N_9239,N_7738);
nor UO_763 (O_763,N_7787,N_8078);
nor UO_764 (O_764,N_8815,N_9588);
nand UO_765 (O_765,N_7724,N_8374);
or UO_766 (O_766,N_9572,N_9287);
and UO_767 (O_767,N_8518,N_9366);
and UO_768 (O_768,N_8591,N_7614);
nand UO_769 (O_769,N_9257,N_8605);
or UO_770 (O_770,N_8782,N_7860);
and UO_771 (O_771,N_7543,N_9307);
nor UO_772 (O_772,N_9120,N_7931);
nor UO_773 (O_773,N_9839,N_8595);
or UO_774 (O_774,N_9670,N_8592);
or UO_775 (O_775,N_9126,N_8616);
nor UO_776 (O_776,N_9417,N_8212);
and UO_777 (O_777,N_9381,N_8264);
nand UO_778 (O_778,N_8584,N_8255);
and UO_779 (O_779,N_8528,N_8224);
nand UO_780 (O_780,N_8651,N_8032);
nor UO_781 (O_781,N_9545,N_9146);
nand UO_782 (O_782,N_9386,N_9928);
or UO_783 (O_783,N_8252,N_8890);
and UO_784 (O_784,N_8238,N_8813);
nand UO_785 (O_785,N_9447,N_8048);
nor UO_786 (O_786,N_8278,N_8208);
or UO_787 (O_787,N_7531,N_9349);
or UO_788 (O_788,N_8831,N_8044);
or UO_789 (O_789,N_9377,N_9459);
nand UO_790 (O_790,N_7900,N_9859);
and UO_791 (O_791,N_8713,N_9030);
or UO_792 (O_792,N_7890,N_9885);
nand UO_793 (O_793,N_8153,N_9217);
or UO_794 (O_794,N_9043,N_9713);
nor UO_795 (O_795,N_7827,N_8641);
and UO_796 (O_796,N_8817,N_8739);
nand UO_797 (O_797,N_9795,N_8236);
nand UO_798 (O_798,N_9693,N_9441);
nor UO_799 (O_799,N_8194,N_9435);
or UO_800 (O_800,N_9371,N_8626);
nand UO_801 (O_801,N_9484,N_9704);
nor UO_802 (O_802,N_9536,N_8288);
or UO_803 (O_803,N_8905,N_9138);
or UO_804 (O_804,N_7798,N_8156);
and UO_805 (O_805,N_8446,N_9258);
nor UO_806 (O_806,N_8876,N_7981);
nor UO_807 (O_807,N_7646,N_9468);
nand UO_808 (O_808,N_7726,N_9926);
nor UO_809 (O_809,N_9656,N_9454);
and UO_810 (O_810,N_9690,N_8668);
nand UO_811 (O_811,N_9291,N_9285);
nand UO_812 (O_812,N_8575,N_8550);
nor UO_813 (O_813,N_7581,N_9439);
and UO_814 (O_814,N_8881,N_8226);
or UO_815 (O_815,N_9866,N_8415);
nor UO_816 (O_816,N_7671,N_8269);
or UO_817 (O_817,N_8855,N_9720);
nor UO_818 (O_818,N_8461,N_9118);
and UO_819 (O_819,N_9985,N_9100);
and UO_820 (O_820,N_9403,N_7849);
or UO_821 (O_821,N_7572,N_8662);
nand UO_822 (O_822,N_9171,N_9105);
nor UO_823 (O_823,N_9220,N_9782);
nor UO_824 (O_824,N_8765,N_9378);
nand UO_825 (O_825,N_9345,N_9584);
and UO_826 (O_826,N_9598,N_9293);
or UO_827 (O_827,N_7594,N_8945);
nor UO_828 (O_828,N_8307,N_7645);
or UO_829 (O_829,N_7609,N_9500);
and UO_830 (O_830,N_8383,N_8795);
nor UO_831 (O_831,N_7939,N_7642);
xnor UO_832 (O_832,N_8393,N_9730);
nor UO_833 (O_833,N_9197,N_8075);
nand UO_834 (O_834,N_8070,N_7807);
or UO_835 (O_835,N_9762,N_8392);
or UO_836 (O_836,N_9460,N_7904);
nand UO_837 (O_837,N_9573,N_7919);
and UO_838 (O_838,N_8137,N_9199);
nor UO_839 (O_839,N_7537,N_9492);
and UO_840 (O_840,N_9290,N_9438);
nand UO_841 (O_841,N_7601,N_7547);
nand UO_842 (O_842,N_8784,N_7847);
and UO_843 (O_843,N_8610,N_8688);
nor UO_844 (O_844,N_9124,N_9049);
or UO_845 (O_845,N_7803,N_7644);
and UO_846 (O_846,N_7855,N_8478);
nor UO_847 (O_847,N_9678,N_9164);
nor UO_848 (O_848,N_8751,N_8501);
or UO_849 (O_849,N_9895,N_9387);
nor UO_850 (O_850,N_9288,N_7592);
or UO_851 (O_851,N_8067,N_9804);
or UO_852 (O_852,N_9278,N_7673);
nand UO_853 (O_853,N_7735,N_7768);
nand UO_854 (O_854,N_7895,N_8534);
nand UO_855 (O_855,N_9096,N_9383);
nand UO_856 (O_856,N_9035,N_8469);
xor UO_857 (O_857,N_9464,N_7510);
and UO_858 (O_858,N_8794,N_7575);
nand UO_859 (O_859,N_7639,N_8390);
and UO_860 (O_860,N_7634,N_8618);
nand UO_861 (O_861,N_8214,N_9410);
nor UO_862 (O_862,N_7599,N_9396);
or UO_863 (O_863,N_9722,N_9615);
nor UO_864 (O_864,N_9672,N_8708);
and UO_865 (O_865,N_8021,N_8508);
nand UO_866 (O_866,N_8988,N_7999);
and UO_867 (O_867,N_8933,N_8742);
nand UO_868 (O_868,N_8635,N_8632);
or UO_869 (O_869,N_7874,N_7778);
or UO_870 (O_870,N_9192,N_8423);
nor UO_871 (O_871,N_9921,N_9654);
nor UO_872 (O_872,N_9641,N_9824);
nand UO_873 (O_873,N_8247,N_8322);
nand UO_874 (O_874,N_8098,N_7792);
nand UO_875 (O_875,N_8101,N_8539);
nand UO_876 (O_876,N_9901,N_8366);
or UO_877 (O_877,N_8975,N_9482);
nor UO_878 (O_878,N_8346,N_7856);
or UO_879 (O_879,N_9657,N_7528);
and UO_880 (O_880,N_9665,N_9083);
nand UO_881 (O_881,N_9424,N_9698);
or UO_882 (O_882,N_9863,N_7816);
and UO_883 (O_883,N_9780,N_9457);
nand UO_884 (O_884,N_7725,N_8755);
nor UO_885 (O_885,N_8190,N_7927);
and UO_886 (O_886,N_7831,N_9204);
and UO_887 (O_887,N_7837,N_9123);
and UO_888 (O_888,N_8872,N_8280);
xnor UO_889 (O_889,N_8848,N_8119);
nor UO_890 (O_890,N_8611,N_9964);
nand UO_891 (O_891,N_8019,N_8903);
or UO_892 (O_892,N_8566,N_8775);
and UO_893 (O_893,N_9807,N_8797);
and UO_894 (O_894,N_8996,N_8109);
nand UO_895 (O_895,N_8052,N_7937);
nor UO_896 (O_896,N_8910,N_9966);
and UO_897 (O_897,N_9311,N_8697);
nand UO_898 (O_898,N_8102,N_9490);
and UO_899 (O_899,N_8259,N_9796);
and UO_900 (O_900,N_9148,N_8290);
and UO_901 (O_901,N_8391,N_9717);
and UO_902 (O_902,N_8457,N_7789);
or UO_903 (O_903,N_8807,N_7617);
nor UO_904 (O_904,N_9786,N_9662);
nor UO_905 (O_905,N_9684,N_8276);
and UO_906 (O_906,N_9600,N_9994);
or UO_907 (O_907,N_8762,N_7536);
and UO_908 (O_908,N_9707,N_8034);
or UO_909 (O_909,N_8870,N_9709);
or UO_910 (O_910,N_8240,N_8013);
nor UO_911 (O_911,N_8202,N_7717);
and UO_912 (O_912,N_8159,N_8814);
or UO_913 (O_913,N_9149,N_8682);
nor UO_914 (O_914,N_7667,N_8888);
nor UO_915 (O_915,N_8517,N_7990);
and UO_916 (O_916,N_7947,N_8121);
nor UO_917 (O_917,N_8055,N_7589);
nor UO_918 (O_918,N_9645,N_9101);
and UO_919 (O_919,N_8854,N_7901);
or UO_920 (O_920,N_7780,N_7615);
nand UO_921 (O_921,N_8116,N_7748);
or UO_922 (O_922,N_9963,N_9334);
or UO_923 (O_923,N_7897,N_7740);
nor UO_924 (O_924,N_9827,N_9405);
and UO_925 (O_925,N_8691,N_8603);
nor UO_926 (O_926,N_7935,N_7957);
nor UO_927 (O_927,N_9318,N_8318);
or UO_928 (O_928,N_8358,N_8219);
or UO_929 (O_929,N_8640,N_8113);
and UO_930 (O_930,N_7795,N_8341);
nor UO_931 (O_931,N_9423,N_7516);
nor UO_932 (O_932,N_9320,N_8158);
or UO_933 (O_933,N_7891,N_9193);
nand UO_934 (O_934,N_7731,N_8426);
nor UO_935 (O_935,N_9783,N_8530);
nand UO_936 (O_936,N_8703,N_9425);
or UO_937 (O_937,N_7951,N_9427);
and UO_938 (O_938,N_8429,N_8244);
and UO_939 (O_939,N_7863,N_9531);
nor UO_940 (O_940,N_8773,N_8825);
and UO_941 (O_941,N_9924,N_7840);
nor UO_942 (O_942,N_8680,N_7616);
nand UO_943 (O_943,N_9601,N_7854);
nor UO_944 (O_944,N_9000,N_8588);
nand UO_945 (O_945,N_9494,N_9212);
or UO_946 (O_946,N_7625,N_8693);
and UO_947 (O_947,N_9513,N_9620);
and UO_948 (O_948,N_7994,N_9692);
and UO_949 (O_949,N_8311,N_9430);
nor UO_950 (O_950,N_9184,N_8748);
and UO_951 (O_951,N_9580,N_7635);
nor UO_952 (O_952,N_8372,N_8653);
and UO_953 (O_953,N_9006,N_8299);
and UO_954 (O_954,N_8589,N_7506);
nand UO_955 (O_955,N_8563,N_9214);
or UO_956 (O_956,N_8899,N_7809);
or UO_957 (O_957,N_7624,N_8310);
and UO_958 (O_958,N_7577,N_8049);
nand UO_959 (O_959,N_8345,N_8862);
or UO_960 (O_960,N_8490,N_8936);
nand UO_961 (O_961,N_9829,N_8676);
nor UO_962 (O_962,N_8504,N_9188);
nand UO_963 (O_963,N_8412,N_7830);
or UO_964 (O_964,N_8430,N_9016);
nand UO_965 (O_965,N_7753,N_7833);
and UO_966 (O_966,N_8180,N_9340);
nor UO_967 (O_967,N_9627,N_9930);
nor UO_968 (O_968,N_9428,N_8010);
or UO_969 (O_969,N_8757,N_8552);
or UO_970 (O_970,N_8403,N_8460);
nor UO_971 (O_971,N_7944,N_9098);
and UO_972 (O_972,N_7765,N_7713);
or UO_973 (O_973,N_8628,N_8946);
and UO_974 (O_974,N_9978,N_8683);
or UO_975 (O_975,N_8268,N_9853);
and UO_976 (O_976,N_8636,N_9300);
or UO_977 (O_977,N_9458,N_9820);
or UO_978 (O_978,N_8376,N_9555);
nor UO_979 (O_979,N_9048,N_8088);
nor UO_980 (O_980,N_8126,N_9550);
nor UO_981 (O_981,N_7817,N_7658);
nor UO_982 (O_982,N_8371,N_8313);
or UO_983 (O_983,N_7647,N_8833);
nand UO_984 (O_984,N_8827,N_9705);
nor UO_985 (O_985,N_9008,N_8411);
nor UO_986 (O_986,N_8527,N_8922);
and UO_987 (O_987,N_9932,N_8587);
and UO_988 (O_988,N_8836,N_9081);
nand UO_989 (O_989,N_8111,N_7872);
nand UO_990 (O_990,N_8958,N_8005);
nor UO_991 (O_991,N_9995,N_8886);
or UO_992 (O_992,N_9127,N_9675);
or UO_993 (O_993,N_8648,N_8436);
and UO_994 (O_994,N_8624,N_8196);
nand UO_995 (O_995,N_9810,N_8350);
nand UO_996 (O_996,N_8665,N_9442);
nor UO_997 (O_997,N_9861,N_9335);
nor UO_998 (O_998,N_8917,N_9177);
and UO_999 (O_999,N_7771,N_9514);
nor UO_1000 (O_1000,N_7665,N_9889);
or UO_1001 (O_1001,N_9289,N_9388);
nor UO_1002 (O_1002,N_8654,N_7921);
and UO_1003 (O_1003,N_8667,N_8414);
nand UO_1004 (O_1004,N_9067,N_9826);
nand UO_1005 (O_1005,N_7834,N_7786);
and UO_1006 (O_1006,N_9956,N_8132);
nand UO_1007 (O_1007,N_8913,N_9132);
nand UO_1008 (O_1008,N_9830,N_8025);
or UO_1009 (O_1009,N_7677,N_7504);
nor UO_1010 (O_1010,N_9172,N_9739);
or UO_1011 (O_1011,N_9890,N_8047);
and UO_1012 (O_1012,N_8702,N_9897);
nor UO_1013 (O_1013,N_8401,N_9077);
nor UO_1014 (O_1014,N_8129,N_8597);
or UO_1015 (O_1015,N_9044,N_7956);
xnor UO_1016 (O_1016,N_8106,N_9832);
nor UO_1017 (O_1017,N_8995,N_9061);
nand UO_1018 (O_1018,N_9880,N_7879);
or UO_1019 (O_1019,N_7754,N_9316);
nand UO_1020 (O_1020,N_9944,N_9353);
and UO_1021 (O_1021,N_9091,N_8195);
nor UO_1022 (O_1022,N_8154,N_9977);
and UO_1023 (O_1023,N_7806,N_8084);
nand UO_1024 (O_1024,N_8829,N_8023);
nor UO_1025 (O_1025,N_8586,N_9475);
or UO_1026 (O_1026,N_9415,N_9593);
nand UO_1027 (O_1027,N_9094,N_9554);
nor UO_1028 (O_1028,N_8352,N_8039);
nand UO_1029 (O_1029,N_7597,N_9556);
or UO_1030 (O_1030,N_9735,N_8453);
or UO_1031 (O_1031,N_9606,N_8837);
and UO_1032 (O_1032,N_9223,N_9407);
or UO_1033 (O_1033,N_8642,N_8027);
or UO_1034 (O_1034,N_9368,N_9661);
nand UO_1035 (O_1035,N_9715,N_7555);
nor UO_1036 (O_1036,N_7930,N_8324);
nand UO_1037 (O_1037,N_9976,N_9643);
nor UO_1038 (O_1038,N_8627,N_9263);
nor UO_1039 (O_1039,N_9053,N_9169);
nor UO_1040 (O_1040,N_8546,N_8834);
nand UO_1041 (O_1041,N_8326,N_8843);
and UO_1042 (O_1042,N_7573,N_8949);
and UO_1043 (O_1043,N_9870,N_9251);
or UO_1044 (O_1044,N_9108,N_7626);
nand UO_1045 (O_1045,N_9714,N_7912);
nor UO_1046 (O_1046,N_8625,N_8964);
nor UO_1047 (O_1047,N_8498,N_8409);
xnor UO_1048 (O_1048,N_8090,N_9176);
and UO_1049 (O_1049,N_9872,N_8856);
nand UO_1050 (O_1050,N_8671,N_9653);
xor UO_1051 (O_1051,N_9664,N_7894);
and UO_1052 (O_1052,N_9027,N_9121);
and UO_1053 (O_1053,N_8660,N_9230);
and UO_1054 (O_1054,N_8987,N_8532);
or UO_1055 (O_1055,N_9648,N_9376);
nand UO_1056 (O_1056,N_8772,N_9878);
nand UO_1057 (O_1057,N_8347,N_9446);
nor UO_1058 (O_1058,N_8538,N_9950);
or UO_1059 (O_1059,N_8033,N_8818);
nor UO_1060 (O_1060,N_8043,N_8229);
nand UO_1061 (O_1061,N_8567,N_8939);
nor UO_1062 (O_1062,N_7790,N_8150);
nor UO_1063 (O_1063,N_9060,N_9364);
nor UO_1064 (O_1064,N_7655,N_8217);
nand UO_1065 (O_1065,N_9483,N_7545);
nand UO_1066 (O_1066,N_7970,N_9579);
nand UO_1067 (O_1067,N_8914,N_8486);
nor UO_1068 (O_1068,N_8812,N_9064);
or UO_1069 (O_1069,N_8396,N_8141);
nand UO_1070 (O_1070,N_8309,N_8820);
and UO_1071 (O_1071,N_7709,N_7769);
or UO_1072 (O_1072,N_9965,N_7714);
and UO_1073 (O_1073,N_8920,N_8321);
and UO_1074 (O_1074,N_9131,N_8063);
nor UO_1075 (O_1075,N_7980,N_8256);
nor UO_1076 (O_1076,N_9063,N_7715);
or UO_1077 (O_1077,N_8558,N_9685);
nand UO_1078 (O_1078,N_8578,N_8568);
nor UO_1079 (O_1079,N_8386,N_9226);
and UO_1080 (O_1080,N_9252,N_7907);
or UO_1081 (O_1081,N_9106,N_8107);
nor UO_1082 (O_1082,N_8867,N_9908);
and UO_1083 (O_1083,N_7550,N_9462);
nand UO_1084 (O_1084,N_8853,N_7868);
nand UO_1085 (O_1085,N_9669,N_8615);
or UO_1086 (O_1086,N_9125,N_7761);
or UO_1087 (O_1087,N_8379,N_9356);
nand UO_1088 (O_1088,N_8983,N_8283);
nand UO_1089 (O_1089,N_9367,N_8932);
nand UO_1090 (O_1090,N_7694,N_9375);
xor UO_1091 (O_1091,N_8543,N_9768);
nand UO_1092 (O_1092,N_8487,N_8944);
nor UO_1093 (O_1093,N_8117,N_9574);
or UO_1094 (O_1094,N_8496,N_8684);
nand UO_1095 (O_1095,N_7964,N_9959);
and UO_1096 (O_1096,N_8796,N_9037);
or UO_1097 (O_1097,N_9636,N_8931);
and UO_1098 (O_1098,N_9632,N_8620);
and UO_1099 (O_1099,N_7515,N_9628);
and UO_1100 (O_1100,N_7517,N_9667);
nor UO_1101 (O_1101,N_9534,N_7801);
nor UO_1102 (O_1102,N_8059,N_9743);
and UO_1103 (O_1103,N_7892,N_9191);
and UO_1104 (O_1104,N_8894,N_8397);
nor UO_1105 (O_1105,N_7796,N_9790);
nor UO_1106 (O_1106,N_9886,N_7722);
and UO_1107 (O_1107,N_7923,N_9508);
or UO_1108 (O_1108,N_9973,N_7666);
or UO_1109 (O_1109,N_8398,N_8416);
nor UO_1110 (O_1110,N_8778,N_8138);
and UO_1111 (O_1111,N_9350,N_7743);
or UO_1112 (O_1112,N_9159,N_8381);
nand UO_1113 (O_1113,N_8717,N_8360);
or UO_1114 (O_1114,N_9763,N_7969);
or UO_1115 (O_1115,N_8644,N_7613);
nor UO_1116 (O_1116,N_8965,N_8896);
or UO_1117 (O_1117,N_8601,N_9652);
and UO_1118 (O_1118,N_8459,N_7915);
nor UO_1119 (O_1119,N_8972,N_9840);
nand UO_1120 (O_1120,N_8037,N_7737);
or UO_1121 (O_1121,N_9373,N_9161);
nand UO_1122 (O_1122,N_7922,N_8711);
nand UO_1123 (O_1123,N_8685,N_8533);
nand UO_1124 (O_1124,N_8491,N_7530);
nor UO_1125 (O_1125,N_9362,N_9539);
nor UO_1126 (O_1126,N_9821,N_8115);
nor UO_1127 (O_1127,N_9294,N_8520);
nor UO_1128 (O_1128,N_7565,N_9658);
nand UO_1129 (O_1129,N_8967,N_9111);
or UO_1130 (O_1130,N_9095,N_8547);
or UO_1131 (O_1131,N_7898,N_7718);
and UO_1132 (O_1132,N_8895,N_7501);
or UO_1133 (O_1133,N_8354,N_9074);
nor UO_1134 (O_1134,N_9602,N_8602);
or UO_1135 (O_1135,N_9637,N_7810);
or UO_1136 (O_1136,N_7675,N_9186);
nor UO_1137 (O_1137,N_7843,N_8571);
xnor UO_1138 (O_1138,N_9723,N_8002);
and UO_1139 (O_1139,N_8724,N_8103);
or UO_1140 (O_1140,N_8916,N_9444);
and UO_1141 (O_1141,N_8072,N_8041);
and UO_1142 (O_1142,N_9404,N_9143);
xnor UO_1143 (O_1143,N_7700,N_8464);
and UO_1144 (O_1144,N_9142,N_7905);
and UO_1145 (O_1145,N_7764,N_7929);
nor UO_1146 (O_1146,N_7808,N_8790);
and UO_1147 (O_1147,N_9957,N_8325);
nor UO_1148 (O_1148,N_8384,N_8562);
xor UO_1149 (O_1149,N_8331,N_9590);
or UO_1150 (O_1150,N_9655,N_8704);
and UO_1151 (O_1151,N_9265,N_9073);
nand UO_1152 (O_1152,N_8969,N_9219);
and UO_1153 (O_1153,N_9372,N_9946);
or UO_1154 (O_1154,N_8956,N_9011);
nor UO_1155 (O_1155,N_7934,N_9463);
and UO_1156 (O_1156,N_9380,N_8509);
and UO_1157 (O_1157,N_8444,N_8105);
nand UO_1158 (O_1158,N_9041,N_8780);
or UO_1159 (O_1159,N_8868,N_9401);
nor UO_1160 (O_1160,N_7751,N_8884);
or UO_1161 (O_1161,N_9646,N_8907);
or UO_1162 (O_1162,N_8157,N_8237);
and UO_1163 (O_1163,N_9133,N_8239);
and UO_1164 (O_1164,N_9321,N_7966);
or UO_1165 (O_1165,N_9411,N_8124);
or UO_1166 (O_1166,N_8659,N_7842);
and UO_1167 (O_1167,N_7839,N_9814);
or UO_1168 (O_1168,N_7564,N_9416);
or UO_1169 (O_1169,N_9082,N_7549);
or UO_1170 (O_1170,N_7760,N_8056);
and UO_1171 (O_1171,N_9718,N_8502);
nor UO_1172 (O_1172,N_9608,N_9833);
or UO_1173 (O_1173,N_9487,N_9919);
nand UO_1174 (O_1174,N_8370,N_7640);
nor UO_1175 (O_1175,N_7539,N_9734);
nand UO_1176 (O_1176,N_7962,N_9638);
and UO_1177 (O_1177,N_8819,N_9806);
or UO_1178 (O_1178,N_9260,N_7799);
or UO_1179 (O_1179,N_8860,N_8767);
and UO_1180 (O_1180,N_8073,N_8079);
and UO_1181 (O_1181,N_8006,N_8375);
nor UO_1182 (O_1182,N_9955,N_9673);
and UO_1183 (O_1183,N_9418,N_9953);
and UO_1184 (O_1184,N_8841,N_9266);
or UO_1185 (O_1185,N_7974,N_9068);
or UO_1186 (O_1186,N_9358,N_9551);
and UO_1187 (O_1187,N_8536,N_8258);
nand UO_1188 (O_1188,N_8145,N_8261);
and UO_1189 (O_1189,N_9254,N_9873);
nand UO_1190 (O_1190,N_9914,N_8445);
or UO_1191 (O_1191,N_8937,N_9616);
or UO_1192 (O_1192,N_8484,N_7755);
or UO_1193 (O_1193,N_7772,N_8839);
and UO_1194 (O_1194,N_9109,N_7797);
or UO_1195 (O_1195,N_8764,N_8184);
and UO_1196 (O_1196,N_9674,N_9235);
or UO_1197 (O_1197,N_7893,N_9865);
nor UO_1198 (O_1198,N_8015,N_8842);
or UO_1199 (O_1199,N_9256,N_8012);
or UO_1200 (O_1200,N_8000,N_9526);
nand UO_1201 (O_1201,N_8165,N_7881);
or UO_1202 (O_1202,N_7538,N_8179);
or UO_1203 (O_1203,N_8335,N_7678);
and UO_1204 (O_1204,N_9225,N_8898);
or UO_1205 (O_1205,N_9162,N_7902);
nor UO_1206 (O_1206,N_8205,N_8649);
or UO_1207 (O_1207,N_9549,N_9426);
nand UO_1208 (O_1208,N_8789,N_9075);
or UO_1209 (O_1209,N_8197,N_9518);
nand UO_1210 (O_1210,N_7643,N_9893);
nor UO_1211 (O_1211,N_8869,N_8658);
and UO_1212 (O_1212,N_7511,N_9145);
or UO_1213 (O_1213,N_8799,N_7928);
and UO_1214 (O_1214,N_7876,N_9649);
nand UO_1215 (O_1215,N_9466,N_8035);
or UO_1216 (O_1216,N_9026,N_9828);
nor UO_1217 (O_1217,N_7710,N_9039);
and UO_1218 (O_1218,N_9012,N_8994);
and UO_1219 (O_1219,N_8885,N_9603);
nand UO_1220 (O_1220,N_8993,N_9203);
nand UO_1221 (O_1221,N_7559,N_7746);
nor UO_1222 (O_1222,N_8301,N_9505);
and UO_1223 (O_1223,N_8467,N_9564);
and UO_1224 (O_1224,N_9168,N_8182);
nand UO_1225 (O_1225,N_8741,N_9510);
or UO_1226 (O_1226,N_8793,N_9612);
nand UO_1227 (O_1227,N_7664,N_8332);
nand UO_1228 (O_1228,N_9322,N_8369);
nor UO_1229 (O_1229,N_8878,N_8721);
nand UO_1230 (O_1230,N_9071,N_8503);
or UO_1231 (O_1231,N_8846,N_9624);
nand UO_1232 (O_1232,N_7519,N_9506);
and UO_1233 (O_1233,N_8463,N_7533);
or UO_1234 (O_1234,N_9363,N_7794);
and UO_1235 (O_1235,N_9038,N_7866);
or UO_1236 (O_1236,N_8071,N_9629);
nand UO_1237 (O_1237,N_9154,N_8968);
nand UO_1238 (O_1238,N_7633,N_9170);
nand UO_1239 (O_1239,N_9595,N_9443);
or UO_1240 (O_1240,N_9659,N_9942);
nor UO_1241 (O_1241,N_9312,N_9004);
nor UO_1242 (O_1242,N_9066,N_8303);
xnor UO_1243 (O_1243,N_8251,N_9218);
nand UO_1244 (O_1244,N_8216,N_7784);
nand UO_1245 (O_1245,N_9135,N_9250);
and UO_1246 (O_1246,N_9504,N_9240);
or UO_1247 (O_1247,N_9032,N_7598);
or UO_1248 (O_1248,N_9103,N_9617);
or UO_1249 (O_1249,N_8977,N_9078);
or UO_1250 (O_1250,N_9633,N_8238);
or UO_1251 (O_1251,N_9509,N_9309);
nand UO_1252 (O_1252,N_9446,N_8695);
nand UO_1253 (O_1253,N_8204,N_9710);
or UO_1254 (O_1254,N_8372,N_7587);
nand UO_1255 (O_1255,N_9181,N_8892);
nor UO_1256 (O_1256,N_7727,N_8546);
or UO_1257 (O_1257,N_9544,N_9830);
and UO_1258 (O_1258,N_9438,N_9220);
nand UO_1259 (O_1259,N_7943,N_8573);
or UO_1260 (O_1260,N_9651,N_7743);
and UO_1261 (O_1261,N_7788,N_8774);
nor UO_1262 (O_1262,N_7958,N_9008);
nand UO_1263 (O_1263,N_9720,N_8828);
nand UO_1264 (O_1264,N_8135,N_7898);
nand UO_1265 (O_1265,N_9177,N_7835);
nor UO_1266 (O_1266,N_9016,N_7628);
and UO_1267 (O_1267,N_9513,N_9285);
and UO_1268 (O_1268,N_8743,N_9070);
or UO_1269 (O_1269,N_8339,N_9762);
and UO_1270 (O_1270,N_9867,N_8342);
or UO_1271 (O_1271,N_9336,N_8764);
and UO_1272 (O_1272,N_9900,N_8288);
nand UO_1273 (O_1273,N_9595,N_9666);
and UO_1274 (O_1274,N_8644,N_7595);
xor UO_1275 (O_1275,N_9732,N_9696);
nor UO_1276 (O_1276,N_7532,N_8388);
nand UO_1277 (O_1277,N_9285,N_9122);
and UO_1278 (O_1278,N_8307,N_8373);
and UO_1279 (O_1279,N_7512,N_8190);
nand UO_1280 (O_1280,N_7680,N_8296);
nand UO_1281 (O_1281,N_7605,N_8110);
nand UO_1282 (O_1282,N_8875,N_8133);
nor UO_1283 (O_1283,N_7585,N_9766);
nand UO_1284 (O_1284,N_7553,N_9622);
and UO_1285 (O_1285,N_9203,N_9783);
nand UO_1286 (O_1286,N_8315,N_9603);
and UO_1287 (O_1287,N_7571,N_9062);
nand UO_1288 (O_1288,N_8007,N_8760);
and UO_1289 (O_1289,N_8526,N_9238);
or UO_1290 (O_1290,N_9268,N_9670);
nor UO_1291 (O_1291,N_9647,N_9309);
or UO_1292 (O_1292,N_8510,N_8312);
xor UO_1293 (O_1293,N_8730,N_9395);
nor UO_1294 (O_1294,N_8727,N_8951);
or UO_1295 (O_1295,N_9494,N_9841);
nand UO_1296 (O_1296,N_9938,N_9620);
or UO_1297 (O_1297,N_9578,N_9493);
and UO_1298 (O_1298,N_9011,N_8415);
nor UO_1299 (O_1299,N_8701,N_8934);
or UO_1300 (O_1300,N_8705,N_8101);
nand UO_1301 (O_1301,N_9698,N_8741);
or UO_1302 (O_1302,N_7995,N_9863);
nor UO_1303 (O_1303,N_8861,N_9232);
or UO_1304 (O_1304,N_7577,N_9708);
and UO_1305 (O_1305,N_9675,N_8013);
or UO_1306 (O_1306,N_7672,N_8232);
nand UO_1307 (O_1307,N_8903,N_8922);
and UO_1308 (O_1308,N_9445,N_7929);
nor UO_1309 (O_1309,N_9951,N_8775);
nor UO_1310 (O_1310,N_8610,N_9512);
nor UO_1311 (O_1311,N_9270,N_8166);
nand UO_1312 (O_1312,N_8968,N_9704);
and UO_1313 (O_1313,N_9443,N_8966);
nand UO_1314 (O_1314,N_8867,N_9274);
and UO_1315 (O_1315,N_7632,N_9396);
or UO_1316 (O_1316,N_7916,N_9993);
nor UO_1317 (O_1317,N_7576,N_8269);
or UO_1318 (O_1318,N_7793,N_8099);
nor UO_1319 (O_1319,N_8351,N_8473);
or UO_1320 (O_1320,N_9135,N_9384);
nor UO_1321 (O_1321,N_9537,N_8044);
and UO_1322 (O_1322,N_8364,N_9266);
or UO_1323 (O_1323,N_8507,N_8636);
nor UO_1324 (O_1324,N_8716,N_9000);
or UO_1325 (O_1325,N_9376,N_8068);
nand UO_1326 (O_1326,N_7866,N_9944);
nand UO_1327 (O_1327,N_7573,N_8248);
nand UO_1328 (O_1328,N_9576,N_9134);
and UO_1329 (O_1329,N_7704,N_7703);
or UO_1330 (O_1330,N_7929,N_7848);
and UO_1331 (O_1331,N_8888,N_7752);
and UO_1332 (O_1332,N_8415,N_9791);
nand UO_1333 (O_1333,N_9539,N_7829);
nor UO_1334 (O_1334,N_9075,N_8174);
and UO_1335 (O_1335,N_9972,N_9345);
nor UO_1336 (O_1336,N_9159,N_9622);
or UO_1337 (O_1337,N_7750,N_7911);
nor UO_1338 (O_1338,N_7748,N_8858);
nor UO_1339 (O_1339,N_8632,N_7678);
and UO_1340 (O_1340,N_8928,N_7626);
and UO_1341 (O_1341,N_9499,N_9124);
and UO_1342 (O_1342,N_7544,N_8019);
or UO_1343 (O_1343,N_9352,N_8873);
or UO_1344 (O_1344,N_8506,N_8901);
or UO_1345 (O_1345,N_9551,N_8173);
or UO_1346 (O_1346,N_9125,N_9263);
nor UO_1347 (O_1347,N_9707,N_8300);
or UO_1348 (O_1348,N_9163,N_9476);
nand UO_1349 (O_1349,N_8716,N_7844);
or UO_1350 (O_1350,N_8206,N_8871);
nor UO_1351 (O_1351,N_7856,N_8079);
or UO_1352 (O_1352,N_7809,N_7845);
and UO_1353 (O_1353,N_9917,N_7827);
nand UO_1354 (O_1354,N_9490,N_7837);
nor UO_1355 (O_1355,N_8930,N_9091);
nor UO_1356 (O_1356,N_8475,N_8386);
and UO_1357 (O_1357,N_7592,N_7869);
nand UO_1358 (O_1358,N_8741,N_9710);
and UO_1359 (O_1359,N_7916,N_8167);
or UO_1360 (O_1360,N_8979,N_9103);
nand UO_1361 (O_1361,N_8296,N_9477);
and UO_1362 (O_1362,N_7759,N_9940);
nand UO_1363 (O_1363,N_9536,N_9592);
or UO_1364 (O_1364,N_8763,N_8743);
and UO_1365 (O_1365,N_8722,N_8192);
nor UO_1366 (O_1366,N_9626,N_7843);
nand UO_1367 (O_1367,N_7624,N_8894);
or UO_1368 (O_1368,N_9835,N_9469);
and UO_1369 (O_1369,N_9817,N_9980);
and UO_1370 (O_1370,N_9823,N_9593);
and UO_1371 (O_1371,N_7577,N_8608);
nor UO_1372 (O_1372,N_9622,N_7837);
nor UO_1373 (O_1373,N_9708,N_9145);
and UO_1374 (O_1374,N_8708,N_8771);
and UO_1375 (O_1375,N_7853,N_9861);
nor UO_1376 (O_1376,N_7795,N_9723);
nand UO_1377 (O_1377,N_9887,N_9175);
nor UO_1378 (O_1378,N_9650,N_8624);
or UO_1379 (O_1379,N_8839,N_7726);
nor UO_1380 (O_1380,N_8551,N_9635);
nor UO_1381 (O_1381,N_8206,N_9920);
nand UO_1382 (O_1382,N_9478,N_8042);
and UO_1383 (O_1383,N_7619,N_9410);
and UO_1384 (O_1384,N_8909,N_8539);
or UO_1385 (O_1385,N_9547,N_8652);
nand UO_1386 (O_1386,N_8428,N_8941);
and UO_1387 (O_1387,N_9756,N_9678);
nand UO_1388 (O_1388,N_8707,N_8440);
or UO_1389 (O_1389,N_8913,N_8398);
nand UO_1390 (O_1390,N_8609,N_8950);
or UO_1391 (O_1391,N_8296,N_9484);
and UO_1392 (O_1392,N_9650,N_8642);
or UO_1393 (O_1393,N_9497,N_8424);
xnor UO_1394 (O_1394,N_9569,N_7785);
and UO_1395 (O_1395,N_8561,N_8128);
and UO_1396 (O_1396,N_8867,N_9545);
nor UO_1397 (O_1397,N_7712,N_8243);
or UO_1398 (O_1398,N_9408,N_9178);
nor UO_1399 (O_1399,N_9433,N_9111);
nor UO_1400 (O_1400,N_7850,N_8469);
nor UO_1401 (O_1401,N_9467,N_9746);
nor UO_1402 (O_1402,N_8102,N_7662);
or UO_1403 (O_1403,N_8933,N_7520);
nor UO_1404 (O_1404,N_8622,N_9350);
nor UO_1405 (O_1405,N_7610,N_8393);
and UO_1406 (O_1406,N_8198,N_7636);
and UO_1407 (O_1407,N_7991,N_9183);
and UO_1408 (O_1408,N_8935,N_8754);
nor UO_1409 (O_1409,N_9664,N_7864);
nand UO_1410 (O_1410,N_9440,N_9612);
nor UO_1411 (O_1411,N_7746,N_8989);
nand UO_1412 (O_1412,N_7649,N_9342);
and UO_1413 (O_1413,N_9432,N_8601);
xor UO_1414 (O_1414,N_9829,N_8451);
or UO_1415 (O_1415,N_7877,N_8176);
and UO_1416 (O_1416,N_9539,N_7876);
and UO_1417 (O_1417,N_7718,N_9680);
nand UO_1418 (O_1418,N_9810,N_9870);
and UO_1419 (O_1419,N_9963,N_8736);
nand UO_1420 (O_1420,N_9174,N_7580);
and UO_1421 (O_1421,N_8810,N_9793);
nand UO_1422 (O_1422,N_7520,N_7783);
xor UO_1423 (O_1423,N_8487,N_7711);
and UO_1424 (O_1424,N_8996,N_9092);
or UO_1425 (O_1425,N_9809,N_9701);
nand UO_1426 (O_1426,N_9257,N_8160);
nor UO_1427 (O_1427,N_9734,N_8952);
and UO_1428 (O_1428,N_8225,N_7767);
or UO_1429 (O_1429,N_9296,N_7683);
or UO_1430 (O_1430,N_9413,N_8981);
or UO_1431 (O_1431,N_7770,N_9312);
nor UO_1432 (O_1432,N_7739,N_8768);
nor UO_1433 (O_1433,N_8667,N_7566);
and UO_1434 (O_1434,N_8743,N_7946);
nor UO_1435 (O_1435,N_8759,N_9585);
nor UO_1436 (O_1436,N_8569,N_8760);
or UO_1437 (O_1437,N_7707,N_8120);
nand UO_1438 (O_1438,N_8655,N_7873);
nor UO_1439 (O_1439,N_9976,N_9150);
nand UO_1440 (O_1440,N_9504,N_9264);
nand UO_1441 (O_1441,N_7959,N_9039);
nor UO_1442 (O_1442,N_8281,N_8915);
or UO_1443 (O_1443,N_8475,N_9287);
or UO_1444 (O_1444,N_9397,N_8053);
or UO_1445 (O_1445,N_9424,N_8186);
or UO_1446 (O_1446,N_9448,N_8701);
nor UO_1447 (O_1447,N_9620,N_9411);
or UO_1448 (O_1448,N_9632,N_9313);
and UO_1449 (O_1449,N_7706,N_9842);
nor UO_1450 (O_1450,N_7569,N_9126);
or UO_1451 (O_1451,N_9157,N_9078);
and UO_1452 (O_1452,N_8672,N_9104);
nand UO_1453 (O_1453,N_8848,N_9639);
and UO_1454 (O_1454,N_7910,N_9127);
nor UO_1455 (O_1455,N_8136,N_9695);
and UO_1456 (O_1456,N_9376,N_8814);
or UO_1457 (O_1457,N_8382,N_8100);
nand UO_1458 (O_1458,N_9655,N_7826);
nand UO_1459 (O_1459,N_9310,N_8076);
or UO_1460 (O_1460,N_8316,N_9204);
nor UO_1461 (O_1461,N_8565,N_9629);
and UO_1462 (O_1462,N_8281,N_9626);
or UO_1463 (O_1463,N_8197,N_7507);
nor UO_1464 (O_1464,N_8415,N_8267);
nand UO_1465 (O_1465,N_7780,N_9897);
and UO_1466 (O_1466,N_7536,N_9902);
nor UO_1467 (O_1467,N_9492,N_7870);
and UO_1468 (O_1468,N_9851,N_8492);
or UO_1469 (O_1469,N_9939,N_9509);
nand UO_1470 (O_1470,N_9007,N_8957);
nor UO_1471 (O_1471,N_8398,N_8087);
nand UO_1472 (O_1472,N_8979,N_8942);
and UO_1473 (O_1473,N_8061,N_9068);
and UO_1474 (O_1474,N_9276,N_8097);
or UO_1475 (O_1475,N_8347,N_8112);
nor UO_1476 (O_1476,N_9396,N_9541);
and UO_1477 (O_1477,N_9409,N_9694);
or UO_1478 (O_1478,N_8613,N_7640);
nand UO_1479 (O_1479,N_8127,N_9411);
nor UO_1480 (O_1480,N_7796,N_8057);
nor UO_1481 (O_1481,N_8209,N_9918);
nand UO_1482 (O_1482,N_9847,N_7723);
and UO_1483 (O_1483,N_9260,N_9174);
nor UO_1484 (O_1484,N_8176,N_9186);
and UO_1485 (O_1485,N_8756,N_9352);
nor UO_1486 (O_1486,N_9450,N_8258);
or UO_1487 (O_1487,N_8692,N_9595);
nor UO_1488 (O_1488,N_8516,N_9028);
and UO_1489 (O_1489,N_8333,N_9051);
or UO_1490 (O_1490,N_7767,N_8916);
nor UO_1491 (O_1491,N_8487,N_9106);
and UO_1492 (O_1492,N_9524,N_8657);
nand UO_1493 (O_1493,N_9409,N_8994);
nor UO_1494 (O_1494,N_8049,N_7946);
nor UO_1495 (O_1495,N_7642,N_9822);
and UO_1496 (O_1496,N_9564,N_7599);
nand UO_1497 (O_1497,N_8632,N_8499);
and UO_1498 (O_1498,N_9609,N_7960);
and UO_1499 (O_1499,N_8387,N_9005);
endmodule