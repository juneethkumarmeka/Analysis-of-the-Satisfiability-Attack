module basic_1000_10000_1500_2_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5006,N_5007,N_5008,N_5009,N_5013,N_5015,N_5016,N_5019,N_5021,N_5022,N_5023,N_5024,N_5025,N_5029,N_5030,N_5035,N_5036,N_5040,N_5041,N_5043,N_5044,N_5046,N_5049,N_5052,N_5053,N_5054,N_5056,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5065,N_5067,N_5068,N_5069,N_5073,N_5074,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5084,N_5085,N_5086,N_5088,N_5089,N_5095,N_5096,N_5097,N_5101,N_5103,N_5105,N_5106,N_5109,N_5110,N_5112,N_5114,N_5117,N_5118,N_5119,N_5120,N_5122,N_5123,N_5124,N_5125,N_5128,N_5131,N_5132,N_5133,N_5135,N_5136,N_5138,N_5139,N_5142,N_5143,N_5145,N_5146,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5158,N_5161,N_5163,N_5164,N_5165,N_5166,N_5172,N_5174,N_5176,N_5177,N_5178,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5189,N_5190,N_5191,N_5193,N_5194,N_5196,N_5197,N_5199,N_5201,N_5202,N_5203,N_5205,N_5206,N_5208,N_5209,N_5211,N_5213,N_5215,N_5216,N_5217,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5227,N_5228,N_5229,N_5230,N_5231,N_5233,N_5234,N_5235,N_5236,N_5238,N_5239,N_5241,N_5242,N_5244,N_5247,N_5248,N_5249,N_5255,N_5258,N_5260,N_5261,N_5263,N_5264,N_5265,N_5267,N_5269,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5278,N_5281,N_5282,N_5283,N_5287,N_5289,N_5291,N_5293,N_5295,N_5296,N_5298,N_5300,N_5303,N_5306,N_5307,N_5309,N_5310,N_5312,N_5314,N_5315,N_5317,N_5319,N_5320,N_5322,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5332,N_5335,N_5337,N_5339,N_5340,N_5341,N_5342,N_5345,N_5347,N_5349,N_5351,N_5352,N_5353,N_5355,N_5357,N_5359,N_5360,N_5361,N_5363,N_5365,N_5366,N_5368,N_5371,N_5372,N_5373,N_5374,N_5377,N_5378,N_5379,N_5381,N_5382,N_5384,N_5385,N_5387,N_5389,N_5390,N_5391,N_5393,N_5394,N_5395,N_5396,N_5397,N_5399,N_5401,N_5405,N_5406,N_5407,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5419,N_5422,N_5424,N_5425,N_5426,N_5429,N_5430,N_5433,N_5435,N_5436,N_5438,N_5440,N_5441,N_5442,N_5445,N_5446,N_5447,N_5450,N_5454,N_5455,N_5457,N_5458,N_5459,N_5461,N_5465,N_5466,N_5467,N_5470,N_5472,N_5473,N_5475,N_5477,N_5479,N_5480,N_5481,N_5482,N_5483,N_5485,N_5486,N_5487,N_5489,N_5490,N_5491,N_5492,N_5495,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5505,N_5506,N_5508,N_5510,N_5511,N_5514,N_5515,N_5516,N_5517,N_5519,N_5521,N_5524,N_5527,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5548,N_5551,N_5552,N_5555,N_5557,N_5559,N_5562,N_5563,N_5566,N_5567,N_5569,N_5572,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5594,N_5596,N_5598,N_5599,N_5600,N_5602,N_5604,N_5606,N_5607,N_5608,N_5609,N_5612,N_5613,N_5614,N_5615,N_5618,N_5619,N_5620,N_5622,N_5625,N_5627,N_5631,N_5635,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5646,N_5647,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5657,N_5658,N_5661,N_5667,N_5668,N_5670,N_5671,N_5672,N_5673,N_5676,N_5677,N_5679,N_5681,N_5683,N_5684,N_5685,N_5686,N_5690,N_5691,N_5693,N_5694,N_5696,N_5702,N_5703,N_5705,N_5707,N_5708,N_5710,N_5711,N_5714,N_5715,N_5716,N_5718,N_5719,N_5720,N_5724,N_5725,N_5726,N_5729,N_5731,N_5733,N_5734,N_5735,N_5739,N_5741,N_5743,N_5744,N_5746,N_5747,N_5749,N_5751,N_5752,N_5753,N_5755,N_5756,N_5757,N_5758,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5775,N_5776,N_5777,N_5779,N_5780,N_5782,N_5783,N_5785,N_5786,N_5787,N_5788,N_5790,N_5795,N_5796,N_5797,N_5798,N_5799,N_5802,N_5803,N_5804,N_5805,N_5806,N_5808,N_5810,N_5811,N_5816,N_5819,N_5821,N_5822,N_5823,N_5825,N_5826,N_5827,N_5828,N_5829,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5838,N_5839,N_5840,N_5842,N_5843,N_5844,N_5845,N_5846,N_5848,N_5849,N_5853,N_5859,N_5860,N_5861,N_5863,N_5864,N_5865,N_5866,N_5869,N_5870,N_5871,N_5872,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5883,N_5884,N_5885,N_5888,N_5891,N_5892,N_5894,N_5896,N_5898,N_5899,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5918,N_5921,N_5923,N_5924,N_5926,N_5929,N_5930,N_5931,N_5932,N_5934,N_5935,N_5936,N_5937,N_5938,N_5940,N_5942,N_5943,N_5944,N_5945,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5955,N_5957,N_5960,N_5961,N_5963,N_5965,N_5966,N_5967,N_5968,N_5969,N_5971,N_5972,N_5973,N_5977,N_5978,N_5979,N_5980,N_5981,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6009,N_6010,N_6014,N_6015,N_6016,N_6017,N_6020,N_6021,N_6022,N_6023,N_6026,N_6027,N_6028,N_6029,N_6031,N_6032,N_6033,N_6036,N_6037,N_6038,N_6040,N_6041,N_6043,N_6044,N_6047,N_6048,N_6049,N_6050,N_6051,N_6053,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6068,N_6069,N_6072,N_6073,N_6076,N_6077,N_6081,N_6082,N_6083,N_6086,N_6087,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6103,N_6105,N_6108,N_6109,N_6110,N_6111,N_6112,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6123,N_6125,N_6126,N_6127,N_6128,N_6129,N_6134,N_6136,N_6139,N_6141,N_6144,N_6145,N_6147,N_6148,N_6149,N_6150,N_6153,N_6154,N_6157,N_6158,N_6161,N_6162,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6177,N_6178,N_6180,N_6182,N_6184,N_6188,N_6189,N_6191,N_6193,N_6194,N_6195,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6206,N_6208,N_6209,N_6210,N_6212,N_6214,N_6216,N_6217,N_6218,N_6219,N_6221,N_6222,N_6223,N_6228,N_6229,N_6230,N_6231,N_6233,N_6234,N_6237,N_6241,N_6243,N_6244,N_6246,N_6247,N_6248,N_6251,N_6252,N_6253,N_6256,N_6260,N_6261,N_6262,N_6264,N_6265,N_6267,N_6269,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6281,N_6283,N_6284,N_6287,N_6288,N_6289,N_6291,N_6292,N_6293,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6309,N_6312,N_6313,N_6315,N_6316,N_6318,N_6319,N_6320,N_6322,N_6324,N_6325,N_6326,N_6327,N_6328,N_6331,N_6334,N_6335,N_6337,N_6339,N_6340,N_6342,N_6343,N_6345,N_6347,N_6349,N_6350,N_6351,N_6352,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6370,N_6371,N_6373,N_6375,N_6376,N_6385,N_6386,N_6388,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6400,N_6401,N_6402,N_6404,N_6406,N_6408,N_6409,N_6410,N_6411,N_6412,N_6414,N_6416,N_6417,N_6418,N_6421,N_6423,N_6425,N_6430,N_6432,N_6435,N_6436,N_6439,N_6441,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6451,N_6453,N_6454,N_6458,N_6459,N_6460,N_6461,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6472,N_6474,N_6476,N_6477,N_6479,N_6480,N_6482,N_6483,N_6484,N_6486,N_6487,N_6490,N_6492,N_6493,N_6497,N_6498,N_6500,N_6502,N_6503,N_6504,N_6506,N_6507,N_6508,N_6509,N_6510,N_6512,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6524,N_6526,N_6528,N_6529,N_6531,N_6532,N_6533,N_6541,N_6542,N_6543,N_6544,N_6547,N_6548,N_6549,N_6552,N_6554,N_6555,N_6556,N_6557,N_6560,N_6561,N_6562,N_6564,N_6565,N_6567,N_6569,N_6570,N_6571,N_6573,N_6574,N_6576,N_6579,N_6580,N_6581,N_6583,N_6584,N_6585,N_6587,N_6589,N_6590,N_6591,N_6595,N_6597,N_6598,N_6599,N_6602,N_6605,N_6607,N_6608,N_6610,N_6612,N_6613,N_6614,N_6615,N_6617,N_6619,N_6624,N_6626,N_6627,N_6628,N_6629,N_6630,N_6633,N_6635,N_6636,N_6637,N_6642,N_6644,N_6646,N_6647,N_6648,N_6649,N_6653,N_6654,N_6655,N_6656,N_6657,N_6659,N_6660,N_6663,N_6664,N_6667,N_6668,N_6671,N_6672,N_6674,N_6677,N_6679,N_6680,N_6681,N_6682,N_6684,N_6687,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6699,N_6700,N_6701,N_6704,N_6707,N_6709,N_6711,N_6712,N_6713,N_6716,N_6717,N_6718,N_6723,N_6724,N_6725,N_6726,N_6728,N_6729,N_6731,N_6732,N_6735,N_6736,N_6737,N_6738,N_6739,N_6742,N_6744,N_6746,N_6747,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6757,N_6758,N_6761,N_6763,N_6764,N_6766,N_6767,N_6769,N_6770,N_6775,N_6776,N_6777,N_6780,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6789,N_6790,N_6791,N_6792,N_6794,N_6798,N_6799,N_6800,N_6804,N_6805,N_6806,N_6807,N_6809,N_6810,N_6811,N_6813,N_6814,N_6815,N_6816,N_6818,N_6820,N_6821,N_6823,N_6824,N_6826,N_6827,N_6829,N_6831,N_6832,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6842,N_6843,N_6844,N_6846,N_6847,N_6848,N_6850,N_6851,N_6852,N_6856,N_6857,N_6859,N_6860,N_6861,N_6864,N_6866,N_6867,N_6868,N_6870,N_6871,N_6873,N_6874,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6883,N_6885,N_6886,N_6887,N_6891,N_6892,N_6896,N_6898,N_6899,N_6901,N_6902,N_6906,N_6907,N_6908,N_6910,N_6911,N_6913,N_6916,N_6917,N_6918,N_6921,N_6922,N_6926,N_6929,N_6931,N_6932,N_6933,N_6934,N_6936,N_6941,N_6944,N_6948,N_6949,N_6951,N_6952,N_6954,N_6955,N_6956,N_6960,N_6962,N_6963,N_6965,N_6966,N_6969,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6981,N_6982,N_6983,N_6986,N_6988,N_6990,N_6991,N_6993,N_6996,N_6997,N_6998,N_6999,N_7001,N_7004,N_7007,N_7008,N_7009,N_7010,N_7012,N_7013,N_7017,N_7018,N_7019,N_7020,N_7023,N_7024,N_7025,N_7026,N_7028,N_7029,N_7030,N_7031,N_7032,N_7039,N_7040,N_7041,N_7043,N_7044,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7056,N_7058,N_7059,N_7064,N_7065,N_7066,N_7068,N_7072,N_7073,N_7074,N_7078,N_7079,N_7080,N_7081,N_7083,N_7086,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7097,N_7100,N_7101,N_7102,N_7103,N_7104,N_7108,N_7109,N_7112,N_7113,N_7115,N_7116,N_7118,N_7119,N_7121,N_7122,N_7123,N_7125,N_7126,N_7127,N_7128,N_7129,N_7131,N_7132,N_7133,N_7137,N_7138,N_7140,N_7143,N_7144,N_7145,N_7147,N_7148,N_7150,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7164,N_7165,N_7167,N_7169,N_7170,N_7171,N_7172,N_7174,N_7175,N_7177,N_7180,N_7182,N_7184,N_7185,N_7186,N_7189,N_7195,N_7196,N_7197,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7211,N_7212,N_7215,N_7217,N_7218,N_7219,N_7224,N_7225,N_7226,N_7227,N_7230,N_7234,N_7236,N_7237,N_7238,N_7240,N_7241,N_7242,N_7243,N_7244,N_7246,N_7248,N_7249,N_7250,N_7253,N_7255,N_7257,N_7259,N_7260,N_7261,N_7262,N_7263,N_7265,N_7266,N_7267,N_7269,N_7272,N_7273,N_7274,N_7276,N_7278,N_7281,N_7282,N_7283,N_7284,N_7286,N_7287,N_7288,N_7289,N_7290,N_7292,N_7297,N_7299,N_7302,N_7303,N_7305,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7322,N_7324,N_7326,N_7329,N_7330,N_7332,N_7334,N_7336,N_7337,N_7338,N_7340,N_7342,N_7344,N_7345,N_7346,N_7347,N_7348,N_7353,N_7354,N_7355,N_7357,N_7358,N_7359,N_7360,N_7361,N_7363,N_7364,N_7367,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7378,N_7380,N_7382,N_7383,N_7384,N_7385,N_7387,N_7389,N_7390,N_7391,N_7392,N_7393,N_7397,N_7398,N_7399,N_7400,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7412,N_7413,N_7420,N_7421,N_7423,N_7425,N_7430,N_7432,N_7433,N_7434,N_7436,N_7437,N_7438,N_7439,N_7442,N_7443,N_7445,N_7446,N_7447,N_7448,N_7449,N_7452,N_7455,N_7457,N_7458,N_7459,N_7461,N_7464,N_7467,N_7468,N_7469,N_7470,N_7473,N_7475,N_7476,N_7478,N_7479,N_7481,N_7483,N_7484,N_7487,N_7489,N_7491,N_7492,N_7493,N_7494,N_7496,N_7500,N_7502,N_7504,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7514,N_7517,N_7523,N_7528,N_7529,N_7531,N_7534,N_7539,N_7541,N_7542,N_7545,N_7546,N_7548,N_7549,N_7551,N_7552,N_7554,N_7555,N_7556,N_7559,N_7561,N_7562,N_7565,N_7567,N_7568,N_7570,N_7571,N_7572,N_7573,N_7574,N_7576,N_7577,N_7581,N_7585,N_7589,N_7592,N_7593,N_7594,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7603,N_7604,N_7607,N_7609,N_7613,N_7615,N_7621,N_7622,N_7626,N_7627,N_7628,N_7632,N_7633,N_7636,N_7637,N_7638,N_7641,N_7642,N_7643,N_7644,N_7647,N_7649,N_7650,N_7652,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7662,N_7663,N_7664,N_7666,N_7667,N_7668,N_7669,N_7672,N_7675,N_7676,N_7677,N_7679,N_7680,N_7681,N_7685,N_7688,N_7690,N_7692,N_7694,N_7695,N_7696,N_7699,N_7700,N_7701,N_7702,N_7703,N_7707,N_7709,N_7710,N_7712,N_7714,N_7715,N_7717,N_7718,N_7719,N_7720,N_7721,N_7723,N_7726,N_7727,N_7728,N_7729,N_7733,N_7735,N_7737,N_7741,N_7745,N_7746,N_7747,N_7748,N_7750,N_7751,N_7752,N_7756,N_7759,N_7760,N_7762,N_7766,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7779,N_7784,N_7785,N_7786,N_7787,N_7791,N_7792,N_7793,N_7795,N_7796,N_7797,N_7799,N_7801,N_7802,N_7803,N_7804,N_7807,N_7808,N_7810,N_7811,N_7813,N_7814,N_7815,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7825,N_7826,N_7827,N_7828,N_7830,N_7832,N_7835,N_7837,N_7838,N_7839,N_7841,N_7843,N_7844,N_7846,N_7851,N_7853,N_7855,N_7856,N_7857,N_7862,N_7863,N_7865,N_7868,N_7869,N_7872,N_7873,N_7877,N_7879,N_7881,N_7882,N_7884,N_7887,N_7891,N_7896,N_7897,N_7898,N_7901,N_7903,N_7905,N_7906,N_7907,N_7909,N_7911,N_7913,N_7914,N_7917,N_7918,N_7922,N_7924,N_7925,N_7926,N_7927,N_7929,N_7937,N_7941,N_7943,N_7945,N_7946,N_7947,N_7952,N_7953,N_7954,N_7958,N_7959,N_7960,N_7964,N_7965,N_7967,N_7968,N_7969,N_7970,N_7971,N_7974,N_7975,N_7979,N_7983,N_7984,N_7985,N_7986,N_7989,N_7992,N_7993,N_7994,N_7996,N_7997,N_7998,N_7999,N_8000,N_8002,N_8003,N_8006,N_8008,N_8009,N_8011,N_8012,N_8014,N_8015,N_8016,N_8018,N_8020,N_8021,N_8022,N_8024,N_8025,N_8026,N_8027,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8037,N_8038,N_8039,N_8041,N_8042,N_8043,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8053,N_8057,N_8058,N_8061,N_8062,N_8063,N_8064,N_8066,N_8068,N_8074,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8084,N_8085,N_8086,N_8087,N_8089,N_8091,N_8093,N_8096,N_8097,N_8098,N_8101,N_8102,N_8104,N_8105,N_8106,N_8107,N_8118,N_8122,N_8124,N_8126,N_8128,N_8130,N_8134,N_8135,N_8136,N_8138,N_8141,N_8142,N_8145,N_8147,N_8149,N_8150,N_8151,N_8152,N_8153,N_8155,N_8157,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8173,N_8177,N_8178,N_8180,N_8181,N_8182,N_8185,N_8186,N_8188,N_8189,N_8190,N_8191,N_8193,N_8195,N_8198,N_8199,N_8200,N_8201,N_8202,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8214,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8237,N_8240,N_8241,N_8242,N_8243,N_8244,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8253,N_8254,N_8255,N_8257,N_8258,N_8259,N_8260,N_8261,N_8263,N_8264,N_8268,N_8269,N_8275,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8284,N_8289,N_8290,N_8291,N_8293,N_8296,N_8297,N_8301,N_8302,N_8305,N_8306,N_8311,N_8313,N_8314,N_8315,N_8316,N_8317,N_8319,N_8322,N_8323,N_8324,N_8327,N_8331,N_8332,N_8333,N_8335,N_8336,N_8337,N_8338,N_8340,N_8342,N_8343,N_8347,N_8348,N_8349,N_8351,N_8354,N_8355,N_8357,N_8361,N_8362,N_8364,N_8366,N_8367,N_8368,N_8369,N_8371,N_8372,N_8374,N_8375,N_8376,N_8377,N_8378,N_8381,N_8384,N_8386,N_8387,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8397,N_8399,N_8400,N_8402,N_8404,N_8405,N_8406,N_8408,N_8413,N_8417,N_8418,N_8419,N_8420,N_8421,N_8423,N_8424,N_8425,N_8426,N_8430,N_8433,N_8435,N_8437,N_8438,N_8440,N_8441,N_8442,N_8443,N_8445,N_8446,N_8448,N_8449,N_8453,N_8454,N_8457,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8472,N_8474,N_8475,N_8477,N_8478,N_8482,N_8485,N_8488,N_8490,N_8491,N_8495,N_8496,N_8497,N_8498,N_8499,N_8504,N_8505,N_8509,N_8511,N_8514,N_8515,N_8516,N_8518,N_8519,N_8520,N_8522,N_8524,N_8526,N_8527,N_8528,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8541,N_8542,N_8543,N_8545,N_8546,N_8548,N_8549,N_8550,N_8551,N_8552,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8563,N_8565,N_8566,N_8568,N_8572,N_8573,N_8574,N_8578,N_8579,N_8581,N_8582,N_8585,N_8586,N_8587,N_8588,N_8590,N_8591,N_8594,N_8595,N_8597,N_8598,N_8599,N_8601,N_8602,N_8604,N_8606,N_8608,N_8609,N_8614,N_8618,N_8620,N_8621,N_8624,N_8627,N_8628,N_8629,N_8630,N_8633,N_8635,N_8639,N_8640,N_8641,N_8642,N_8644,N_8645,N_8646,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8659,N_8660,N_8662,N_8663,N_8664,N_8666,N_8670,N_8671,N_8672,N_8675,N_8678,N_8681,N_8683,N_8684,N_8685,N_8687,N_8689,N_8690,N_8692,N_8694,N_8695,N_8697,N_8698,N_8699,N_8700,N_8701,N_8707,N_8710,N_8712,N_8713,N_8715,N_8716,N_8717,N_8718,N_8722,N_8723,N_8724,N_8726,N_8728,N_8730,N_8731,N_8732,N_8734,N_8737,N_8738,N_8740,N_8741,N_8742,N_8744,N_8745,N_8749,N_8751,N_8752,N_8753,N_8756,N_8758,N_8760,N_8761,N_8763,N_8764,N_8765,N_8767,N_8769,N_8770,N_8772,N_8773,N_8774,N_8775,N_8776,N_8778,N_8779,N_8780,N_8783,N_8784,N_8786,N_8787,N_8788,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8802,N_8803,N_8804,N_8806,N_8808,N_8809,N_8810,N_8811,N_8812,N_8815,N_8816,N_8819,N_8820,N_8822,N_8823,N_8825,N_8826,N_8827,N_8832,N_8833,N_8838,N_8839,N_8841,N_8843,N_8844,N_8845,N_8846,N_8848,N_8849,N_8851,N_8852,N_8853,N_8855,N_8856,N_8857,N_8859,N_8860,N_8861,N_8862,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8873,N_8874,N_8875,N_8876,N_8877,N_8879,N_8880,N_8881,N_8884,N_8885,N_8887,N_8888,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8898,N_8899,N_8900,N_8902,N_8906,N_8908,N_8910,N_8913,N_8916,N_8917,N_8921,N_8922,N_8923,N_8924,N_8925,N_8929,N_8930,N_8932,N_8934,N_8937,N_8938,N_8939,N_8940,N_8941,N_8945,N_8948,N_8949,N_8951,N_8953,N_8955,N_8956,N_8957,N_8959,N_8961,N_8962,N_8964,N_8966,N_8968,N_8969,N_8971,N_8972,N_8974,N_8975,N_8976,N_8977,N_8978,N_8987,N_8990,N_8991,N_8992,N_8993,N_8998,N_8999,N_9000,N_9001,N_9002,N_9004,N_9005,N_9009,N_9010,N_9011,N_9012,N_9014,N_9015,N_9017,N_9018,N_9019,N_9020,N_9022,N_9027,N_9030,N_9032,N_9033,N_9034,N_9036,N_9043,N_9045,N_9046,N_9052,N_9054,N_9056,N_9057,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9066,N_9069,N_9071,N_9075,N_9076,N_9077,N_9079,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9094,N_9096,N_9099,N_9102,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9113,N_9114,N_9116,N_9118,N_9119,N_9120,N_9123,N_9125,N_9127,N_9128,N_9129,N_9131,N_9133,N_9135,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9145,N_9146,N_9147,N_9149,N_9153,N_9154,N_9156,N_9157,N_9158,N_9160,N_9161,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9172,N_9173,N_9174,N_9176,N_9178,N_9179,N_9180,N_9183,N_9184,N_9185,N_9186,N_9187,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9196,N_9198,N_9201,N_9202,N_9203,N_9205,N_9207,N_9208,N_9210,N_9211,N_9213,N_9217,N_9218,N_9220,N_9223,N_9224,N_9227,N_9228,N_9230,N_9231,N_9232,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9241,N_9242,N_9244,N_9245,N_9246,N_9247,N_9249,N_9250,N_9252,N_9255,N_9256,N_9257,N_9261,N_9263,N_9265,N_9266,N_9267,N_9270,N_9273,N_9276,N_9277,N_9278,N_9279,N_9281,N_9284,N_9285,N_9286,N_9287,N_9289,N_9291,N_9293,N_9294,N_9296,N_9303,N_9304,N_9305,N_9307,N_9308,N_9311,N_9313,N_9315,N_9316,N_9318,N_9319,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9328,N_9329,N_9331,N_9333,N_9336,N_9338,N_9340,N_9341,N_9342,N_9344,N_9346,N_9347,N_9348,N_9349,N_9352,N_9355,N_9356,N_9357,N_9358,N_9359,N_9361,N_9363,N_9364,N_9366,N_9367,N_9368,N_9369,N_9372,N_9373,N_9375,N_9376,N_9377,N_9379,N_9381,N_9382,N_9384,N_9386,N_9389,N_9390,N_9395,N_9397,N_9398,N_9399,N_9400,N_9403,N_9404,N_9405,N_9406,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9416,N_9419,N_9421,N_9426,N_9427,N_9428,N_9430,N_9433,N_9435,N_9439,N_9440,N_9441,N_9442,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9452,N_9454,N_9455,N_9456,N_9457,N_9458,N_9461,N_9463,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9475,N_9476,N_9478,N_9480,N_9481,N_9485,N_9486,N_9489,N_9490,N_9491,N_9492,N_9493,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9507,N_9508,N_9510,N_9512,N_9513,N_9514,N_9517,N_9519,N_9522,N_9524,N_9525,N_9526,N_9527,N_9529,N_9530,N_9533,N_9534,N_9535,N_9536,N_9538,N_9539,N_9540,N_9541,N_9542,N_9544,N_9546,N_9547,N_9548,N_9549,N_9551,N_9552,N_9553,N_9554,N_9556,N_9557,N_9562,N_9563,N_9564,N_9565,N_9566,N_9569,N_9572,N_9573,N_9574,N_9575,N_9579,N_9581,N_9584,N_9585,N_9588,N_9589,N_9590,N_9591,N_9593,N_9594,N_9595,N_9596,N_9600,N_9601,N_9602,N_9605,N_9607,N_9608,N_9609,N_9610,N_9614,N_9615,N_9616,N_9617,N_9620,N_9621,N_9626,N_9627,N_9628,N_9629,N_9631,N_9632,N_9633,N_9634,N_9635,N_9637,N_9638,N_9639,N_9641,N_9642,N_9643,N_9646,N_9648,N_9649,N_9651,N_9652,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9663,N_9664,N_9668,N_9669,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9678,N_9679,N_9680,N_9681,N_9684,N_9685,N_9686,N_9687,N_9689,N_9691,N_9694,N_9698,N_9699,N_9700,N_9702,N_9703,N_9704,N_9705,N_9708,N_9711,N_9712,N_9713,N_9716,N_9717,N_9721,N_9724,N_9725,N_9726,N_9727,N_9730,N_9733,N_9735,N_9740,N_9742,N_9744,N_9745,N_9747,N_9748,N_9751,N_9752,N_9755,N_9756,N_9757,N_9758,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9770,N_9774,N_9775,N_9777,N_9778,N_9779,N_9782,N_9783,N_9784,N_9787,N_9791,N_9792,N_9794,N_9795,N_9796,N_9797,N_9798,N_9800,N_9801,N_9805,N_9806,N_9807,N_9810,N_9812,N_9813,N_9814,N_9815,N_9816,N_9818,N_9819,N_9823,N_9824,N_9827,N_9829,N_9830,N_9832,N_9833,N_9835,N_9836,N_9838,N_9840,N_9842,N_9843,N_9845,N_9850,N_9851,N_9852,N_9853,N_9854,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9865,N_9866,N_9868,N_9869,N_9870,N_9872,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9886,N_9887,N_9888,N_9889,N_9891,N_9892,N_9896,N_9898,N_9900,N_9903,N_9906,N_9907,N_9908,N_9910,N_9911,N_9916,N_9917,N_9918,N_9919,N_9921,N_9922,N_9923,N_9924,N_9926,N_9929,N_9931,N_9932,N_9934,N_9936,N_9937,N_9938,N_9939,N_9940,N_9942,N_9946,N_9947,N_9949,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9967,N_9968,N_9970,N_9973,N_9974,N_9976,N_9979,N_9980,N_9981,N_9982,N_9984,N_9986,N_9987,N_9989,N_9990,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_513,In_230);
nor U1 (N_1,In_323,In_625);
nand U2 (N_2,In_550,In_413);
and U3 (N_3,In_375,In_443);
nand U4 (N_4,In_414,In_901);
xnor U5 (N_5,In_336,In_491);
and U6 (N_6,In_638,In_80);
nand U7 (N_7,In_907,In_433);
xor U8 (N_8,In_37,In_938);
xor U9 (N_9,In_205,In_537);
or U10 (N_10,In_632,In_244);
nand U11 (N_11,In_646,In_580);
xor U12 (N_12,In_419,In_3);
and U13 (N_13,In_998,In_502);
nor U14 (N_14,In_705,In_430);
or U15 (N_15,In_78,In_933);
or U16 (N_16,In_824,In_819);
nand U17 (N_17,In_146,In_424);
xnor U18 (N_18,In_755,In_578);
nor U19 (N_19,In_975,In_963);
nor U20 (N_20,In_772,In_354);
and U21 (N_21,In_461,In_607);
xnor U22 (N_22,In_792,In_741);
and U23 (N_23,In_355,In_62);
xnor U24 (N_24,In_642,In_435);
nand U25 (N_25,In_5,In_46);
xnor U26 (N_26,In_978,In_690);
and U27 (N_27,In_965,In_340);
or U28 (N_28,In_591,In_608);
and U29 (N_29,In_472,In_116);
xor U30 (N_30,In_226,In_282);
and U31 (N_31,In_503,In_620);
and U32 (N_32,In_319,In_330);
nor U33 (N_33,In_402,In_379);
xor U34 (N_34,In_884,In_781);
xnor U35 (N_35,In_121,In_889);
or U36 (N_36,In_429,In_717);
or U37 (N_37,In_664,In_564);
nor U38 (N_38,In_799,In_416);
or U39 (N_39,In_233,In_91);
or U40 (N_40,In_881,In_953);
nand U41 (N_41,In_158,In_453);
and U42 (N_42,In_125,In_868);
or U43 (N_43,In_8,In_639);
and U44 (N_44,In_830,In_57);
nor U45 (N_45,In_460,In_659);
nor U46 (N_46,In_65,In_179);
xnor U47 (N_47,In_696,In_411);
xnor U48 (N_48,In_18,In_571);
nor U49 (N_49,In_869,In_95);
nor U50 (N_50,In_152,In_213);
nor U51 (N_51,In_627,In_342);
and U52 (N_52,In_816,In_444);
nand U53 (N_53,In_805,In_315);
and U54 (N_54,In_609,In_959);
xor U55 (N_55,In_641,In_787);
nor U56 (N_56,In_900,In_676);
nand U57 (N_57,In_814,In_692);
xor U58 (N_58,In_228,In_196);
nor U59 (N_59,In_759,In_955);
nand U60 (N_60,In_581,In_716);
nor U61 (N_61,In_990,In_878);
or U62 (N_62,In_221,In_986);
xnor U63 (N_63,In_480,In_989);
nor U64 (N_64,In_55,In_155);
and U65 (N_65,In_268,In_619);
nor U66 (N_66,In_421,In_410);
nor U67 (N_67,In_310,In_668);
xor U68 (N_68,In_209,In_590);
xnor U69 (N_69,In_241,In_86);
nor U70 (N_70,In_64,In_616);
or U71 (N_71,In_686,In_101);
nand U72 (N_72,In_321,In_593);
xnor U73 (N_73,In_111,In_718);
nor U74 (N_74,In_45,In_273);
xnor U75 (N_75,In_836,In_594);
nor U76 (N_76,In_850,In_967);
nand U77 (N_77,In_396,In_937);
nor U78 (N_78,In_4,In_184);
nor U79 (N_79,In_687,In_750);
or U80 (N_80,In_795,In_286);
or U81 (N_81,In_266,In_229);
and U82 (N_82,In_710,In_909);
and U83 (N_83,In_538,In_165);
xor U84 (N_84,In_497,In_366);
nand U85 (N_85,In_259,In_761);
nand U86 (N_86,In_255,In_441);
or U87 (N_87,In_711,In_398);
nand U88 (N_88,In_918,In_670);
or U89 (N_89,In_793,In_983);
or U90 (N_90,In_575,In_631);
or U91 (N_91,In_139,In_349);
and U92 (N_92,In_399,In_964);
nor U93 (N_93,In_358,In_450);
or U94 (N_94,In_370,In_700);
nand U95 (N_95,In_432,In_307);
or U96 (N_96,In_911,In_299);
nor U97 (N_97,In_614,In_389);
or U98 (N_98,In_623,In_777);
nand U99 (N_99,In_23,In_505);
or U100 (N_100,In_512,In_767);
nand U101 (N_101,In_903,In_455);
nand U102 (N_102,In_932,In_465);
nor U103 (N_103,In_574,In_372);
and U104 (N_104,In_504,In_547);
or U105 (N_105,In_689,In_477);
nand U106 (N_106,In_70,In_364);
nand U107 (N_107,In_464,In_498);
nand U108 (N_108,In_207,In_138);
and U109 (N_109,In_22,In_770);
nand U110 (N_110,In_506,In_846);
and U111 (N_111,In_753,In_493);
xor U112 (N_112,In_265,In_913);
xnor U113 (N_113,In_854,In_720);
xnor U114 (N_114,In_954,In_874);
nor U115 (N_115,In_764,In_507);
nor U116 (N_116,In_866,In_181);
xor U117 (N_117,In_611,In_855);
nand U118 (N_118,In_906,In_841);
nor U119 (N_119,In_448,In_300);
or U120 (N_120,In_335,In_79);
or U121 (N_121,In_883,In_54);
or U122 (N_122,In_806,In_789);
or U123 (N_123,In_579,In_756);
nor U124 (N_124,In_308,In_157);
or U125 (N_125,In_539,In_40);
or U126 (N_126,In_865,In_30);
nand U127 (N_127,In_762,In_356);
nand U128 (N_128,In_626,In_114);
nor U129 (N_129,In_980,In_813);
or U130 (N_130,In_663,In_261);
or U131 (N_131,In_985,In_133);
nand U132 (N_132,In_677,In_597);
xor U133 (N_133,In_469,In_104);
nor U134 (N_134,In_306,In_407);
and U135 (N_135,In_13,In_148);
nor U136 (N_136,In_405,In_263);
xnor U137 (N_137,In_406,In_856);
nand U138 (N_138,In_691,In_739);
and U139 (N_139,In_956,In_712);
nor U140 (N_140,In_979,In_784);
nand U141 (N_141,In_377,In_549);
xnor U142 (N_142,In_298,In_216);
nor U143 (N_143,In_724,In_729);
and U144 (N_144,In_942,In_757);
and U145 (N_145,In_17,In_797);
nor U146 (N_146,In_288,In_815);
nor U147 (N_147,In_48,In_170);
nor U148 (N_148,In_327,In_829);
nand U149 (N_149,In_409,In_891);
and U150 (N_150,In_988,In_678);
nor U151 (N_151,In_615,In_16);
and U152 (N_152,In_371,In_749);
and U153 (N_153,In_339,In_754);
and U154 (N_154,In_490,In_807);
nand U155 (N_155,In_38,In_621);
nand U156 (N_156,In_383,In_143);
xor U157 (N_157,In_658,In_803);
nor U158 (N_158,In_332,In_177);
nand U159 (N_159,In_508,In_224);
nor U160 (N_160,In_285,In_195);
nand U161 (N_161,In_704,In_534);
or U162 (N_162,In_861,In_565);
nor U163 (N_163,In_217,In_599);
nor U164 (N_164,In_888,In_128);
nand U165 (N_165,In_301,In_950);
xnor U166 (N_166,In_996,In_630);
and U167 (N_167,In_47,In_701);
and U168 (N_168,In_730,In_648);
nor U169 (N_169,In_246,In_183);
and U170 (N_170,In_434,In_334);
nor U171 (N_171,In_337,In_931);
nand U172 (N_172,In_949,In_360);
nand U173 (N_173,In_873,In_722);
nand U174 (N_174,In_624,In_236);
xor U175 (N_175,In_896,In_20);
nand U176 (N_176,In_408,In_431);
and U177 (N_177,In_773,In_218);
xnor U178 (N_178,In_766,In_516);
nand U179 (N_179,In_733,In_316);
nor U180 (N_180,In_129,In_890);
xnor U181 (N_181,In_857,In_837);
nor U182 (N_182,In_636,In_500);
nand U183 (N_183,In_166,In_665);
or U184 (N_184,In_87,In_7);
nor U185 (N_185,In_518,In_769);
nand U186 (N_186,In_482,In_295);
and U187 (N_187,In_920,In_528);
or U188 (N_188,In_187,In_917);
and U189 (N_189,In_731,In_26);
nor U190 (N_190,In_583,In_847);
or U191 (N_191,In_708,In_737);
or U192 (N_192,In_788,In_897);
xor U193 (N_193,In_400,In_763);
nand U194 (N_194,In_73,In_289);
nand U195 (N_195,In_810,In_385);
and U196 (N_196,In_10,In_489);
and U197 (N_197,In_771,In_804);
and U198 (N_198,In_457,In_381);
nor U199 (N_199,In_163,In_256);
or U200 (N_200,In_248,In_275);
or U201 (N_201,In_557,In_826);
or U202 (N_202,In_351,In_479);
and U203 (N_203,In_290,In_693);
xnor U204 (N_204,In_452,In_2);
nand U205 (N_205,In_403,In_296);
and U206 (N_206,In_966,In_572);
nor U207 (N_207,In_219,In_499);
xnor U208 (N_208,In_728,In_476);
nand U209 (N_209,In_532,In_74);
nand U210 (N_210,In_347,In_438);
and U211 (N_211,In_343,In_936);
or U212 (N_212,In_556,In_56);
or U213 (N_213,In_192,In_660);
xnor U214 (N_214,In_801,In_178);
xnor U215 (N_215,In_530,In_982);
and U216 (N_216,In_67,In_223);
or U217 (N_217,In_214,In_113);
and U218 (N_218,In_822,In_484);
and U219 (N_219,In_117,In_735);
nand U220 (N_220,In_600,In_811);
nand U221 (N_221,In_254,In_291);
nand U222 (N_222,In_833,In_501);
nand U223 (N_223,In_543,In_662);
or U224 (N_224,In_899,In_232);
or U225 (N_225,In_652,In_515);
or U226 (N_226,In_32,In_919);
nor U227 (N_227,In_924,In_736);
xnor U228 (N_228,In_531,In_82);
nor U229 (N_229,In_456,In_12);
and U230 (N_230,In_76,In_27);
and U231 (N_231,In_552,In_258);
or U232 (N_232,In_523,In_270);
or U233 (N_233,In_628,In_544);
xnor U234 (N_234,In_415,In_470);
and U235 (N_235,In_359,In_210);
and U236 (N_236,In_649,In_215);
or U237 (N_237,In_613,In_486);
nand U238 (N_238,In_401,In_58);
and U239 (N_239,In_34,In_667);
or U240 (N_240,In_249,In_318);
nor U241 (N_241,In_368,In_303);
and U242 (N_242,In_987,In_118);
or U243 (N_243,In_951,In_108);
or U244 (N_244,In_605,In_595);
or U245 (N_245,In_317,In_776);
xor U246 (N_246,In_220,In_640);
xnor U247 (N_247,In_545,In_863);
or U248 (N_248,In_714,In_601);
and U249 (N_249,In_175,In_94);
and U250 (N_250,In_783,In_203);
nand U251 (N_251,In_535,In_968);
nand U252 (N_252,In_361,In_130);
and U253 (N_253,In_774,In_972);
nand U254 (N_254,In_393,In_747);
or U255 (N_255,In_684,In_876);
nand U256 (N_256,In_832,In_934);
nor U257 (N_257,In_382,In_387);
or U258 (N_258,In_345,In_109);
nor U259 (N_259,In_939,In_732);
and U260 (N_260,In_893,In_748);
xor U261 (N_261,In_420,In_313);
nand U262 (N_262,In_98,In_745);
nand U263 (N_263,In_743,In_193);
nor U264 (N_264,In_997,In_751);
or U265 (N_265,In_53,In_474);
nor U266 (N_266,In_162,In_522);
and U267 (N_267,In_568,In_160);
xor U268 (N_268,In_782,In_439);
and U269 (N_269,In_706,In_851);
and U270 (N_270,In_365,In_488);
nor U271 (N_271,In_656,In_943);
nor U272 (N_272,In_558,In_471);
or U273 (N_273,In_481,In_147);
and U274 (N_274,In_634,In_765);
nand U275 (N_275,In_200,In_309);
or U276 (N_276,In_463,In_569);
nand U277 (N_277,In_596,In_312);
or U278 (N_278,In_981,In_752);
and U279 (N_279,In_825,In_586);
or U280 (N_280,In_51,In_872);
xnor U281 (N_281,In_362,In_190);
or U282 (N_282,In_645,In_925);
nor U283 (N_283,In_135,In_848);
nand U284 (N_284,In_796,In_529);
nor U285 (N_285,In_322,In_703);
nand U286 (N_286,In_237,In_324);
nor U287 (N_287,In_151,In_390);
nor U288 (N_288,In_827,In_992);
and U289 (N_289,In_929,In_820);
or U290 (N_290,In_467,In_50);
and U291 (N_291,In_940,In_127);
nor U292 (N_292,In_388,In_519);
xor U293 (N_293,In_239,In_885);
nor U294 (N_294,In_898,In_274);
or U295 (N_295,In_587,In_852);
and U296 (N_296,In_606,In_436);
nor U297 (N_297,In_140,In_446);
nand U298 (N_298,In_740,In_576);
xnor U299 (N_299,In_675,In_331);
or U300 (N_300,In_485,In_122);
nor U301 (N_301,In_257,In_914);
and U302 (N_302,In_688,In_926);
xnor U303 (N_303,In_853,In_923);
and U304 (N_304,In_786,In_842);
or U305 (N_305,In_902,In_877);
nor U306 (N_306,In_245,In_397);
xor U307 (N_307,In_746,In_29);
nor U308 (N_308,In_39,In_858);
or U309 (N_309,In_993,In_650);
and U310 (N_310,In_945,In_267);
xnor U311 (N_311,In_928,In_887);
nor U312 (N_312,In_839,In_768);
or U313 (N_313,In_36,In_328);
and U314 (N_314,In_72,In_566);
and U315 (N_315,In_437,In_991);
or U316 (N_316,In_644,In_584);
or U317 (N_317,In_1,In_791);
nor U318 (N_318,In_598,In_844);
nand U319 (N_319,In_352,In_41);
nand U320 (N_320,In_592,In_277);
and U321 (N_321,In_798,In_487);
nand U322 (N_322,In_24,In_554);
xnor U323 (N_323,In_176,In_211);
or U324 (N_324,In_618,In_418);
xor U325 (N_325,In_995,In_617);
or U326 (N_326,In_142,In_633);
nand U327 (N_327,In_510,In_201);
or U328 (N_328,In_679,In_559);
nand U329 (N_329,In_260,In_449);
xor U330 (N_330,In_567,In_159);
or U331 (N_331,In_392,In_81);
or U332 (N_332,In_19,In_653);
or U333 (N_333,In_647,In_694);
and U334 (N_334,In_42,In_191);
and U335 (N_335,In_871,In_831);
nand U336 (N_336,In_131,In_673);
or U337 (N_337,In_90,In_380);
or U338 (N_338,In_802,In_102);
or U339 (N_339,In_671,In_106);
and U340 (N_340,In_188,In_404);
or U341 (N_341,In_304,In_280);
or U342 (N_342,In_553,In_651);
or U343 (N_343,In_173,In_394);
xnor U344 (N_344,In_744,In_97);
nand U345 (N_345,In_373,In_657);
nor U346 (N_346,In_948,In_520);
or U347 (N_347,In_517,In_194);
or U348 (N_348,In_120,In_325);
or U349 (N_349,In_346,In_669);
and U350 (N_350,In_561,In_944);
xnor U351 (N_351,In_725,In_952);
xor U352 (N_352,In_112,In_680);
and U353 (N_353,In_511,In_199);
and U354 (N_354,In_186,In_103);
and U355 (N_355,In_459,In_971);
nor U356 (N_356,In_338,In_521);
xor U357 (N_357,In_843,In_845);
nor U358 (N_358,In_43,In_719);
or U359 (N_359,In_182,In_250);
nor U360 (N_360,In_93,In_234);
or U361 (N_361,In_367,In_661);
xnor U362 (N_362,In_126,In_760);
nor U363 (N_363,In_875,In_137);
xnor U364 (N_364,In_682,In_483);
nand U365 (N_365,In_941,In_14);
nand U366 (N_366,In_478,In_68);
and U367 (N_367,In_738,In_818);
nand U368 (N_368,In_808,In_302);
xnor U369 (N_369,In_252,In_417);
nand U370 (N_370,In_134,In_727);
or U371 (N_371,In_994,In_353);
nand U372 (N_372,In_603,In_473);
nand U373 (N_373,In_425,In_734);
and U374 (N_374,In_107,In_333);
nand U375 (N_375,In_52,In_75);
nor U376 (N_376,In_524,In_150);
nor U377 (N_377,In_915,In_976);
xor U378 (N_378,In_458,In_172);
nor U379 (N_379,In_541,In_59);
xnor U380 (N_380,In_440,In_314);
or U381 (N_381,In_536,In_812);
xnor U382 (N_382,In_683,In_442);
xnor U383 (N_383,In_726,In_573);
nand U384 (N_384,In_61,In_492);
or U385 (N_385,In_879,In_238);
and U386 (N_386,In_376,In_123);
nor U387 (N_387,In_622,In_124);
xnor U388 (N_388,In_284,In_281);
and U389 (N_389,In_922,In_231);
and U390 (N_390,In_862,In_961);
nand U391 (N_391,In_235,In_9);
xor U392 (N_392,In_422,In_984);
or U393 (N_393,In_655,In_629);
xor U394 (N_394,In_742,In_156);
nor U395 (N_395,In_495,In_835);
and U396 (N_396,In_369,In_63);
and U397 (N_397,In_350,In_202);
or U398 (N_398,In_269,In_695);
nand U399 (N_399,In_189,In_864);
nand U400 (N_400,In_702,In_169);
xor U401 (N_401,In_119,In_60);
nand U402 (N_402,In_49,In_582);
nand U403 (N_403,In_311,In_180);
or U404 (N_404,In_612,In_821);
and U405 (N_405,In_840,In_96);
or U406 (N_406,In_905,In_882);
and U407 (N_407,In_794,In_198);
or U408 (N_408,In_962,In_880);
xor U409 (N_409,In_208,In_699);
and U410 (N_410,In_697,In_886);
nor U411 (N_411,In_800,In_916);
and U412 (N_412,In_447,In_363);
or U413 (N_413,In_870,In_715);
and U414 (N_414,In_533,In_859);
xor U415 (N_415,In_88,In_144);
or U416 (N_416,In_391,In_264);
or U417 (N_417,In_698,In_386);
and U418 (N_418,In_935,In_320);
nand U419 (N_419,In_348,In_279);
nor U420 (N_420,In_970,In_153);
or U421 (N_421,In_892,In_610);
nor U422 (N_422,In_560,In_253);
or U423 (N_423,In_15,In_908);
and U424 (N_424,In_240,In_654);
nor U425 (N_425,In_31,In_115);
and U426 (N_426,In_287,In_21);
and U427 (N_427,In_514,In_171);
or U428 (N_428,In_570,In_602);
or U429 (N_429,In_555,In_930);
nor U430 (N_430,In_974,In_164);
and U431 (N_431,In_977,In_604);
xor U432 (N_432,In_85,In_378);
nand U433 (N_433,In_384,In_283);
nand U434 (N_434,In_973,In_785);
nor U435 (N_435,In_721,In_685);
or U436 (N_436,In_585,In_25);
or U437 (N_437,In_723,In_0);
xor U438 (N_438,In_834,In_666);
nand U439 (N_439,In_895,In_779);
and U440 (N_440,In_423,In_357);
nand U441 (N_441,In_509,In_969);
xnor U442 (N_442,In_672,In_293);
nand U443 (N_443,In_161,In_526);
nor U444 (N_444,In_132,In_149);
nand U445 (N_445,In_77,In_958);
and U446 (N_446,In_525,In_412);
nor U447 (N_447,In_242,In_775);
or U448 (N_448,In_894,In_11);
and U449 (N_449,In_790,In_35);
nor U450 (N_450,In_44,In_957);
nor U451 (N_451,In_713,In_527);
or U452 (N_452,In_204,In_99);
or U453 (N_453,In_462,In_946);
nand U454 (N_454,In_197,In_92);
nand U455 (N_455,In_838,In_849);
nor U456 (N_456,In_276,In_344);
nor U457 (N_457,In_428,In_921);
or U458 (N_458,In_71,In_145);
nand U459 (N_459,In_562,In_251);
and U460 (N_460,In_206,In_395);
nor U461 (N_461,In_912,In_947);
or U462 (N_462,In_546,In_867);
xor U463 (N_463,In_66,In_294);
nand U464 (N_464,In_222,In_105);
nor U465 (N_465,In_681,In_329);
or U466 (N_466,In_271,In_185);
or U467 (N_467,In_292,In_272);
xor U468 (N_468,In_305,In_707);
or U469 (N_469,In_100,In_278);
or U470 (N_470,In_643,In_69);
nand U471 (N_471,In_960,In_828);
and U472 (N_472,In_674,In_817);
nand U473 (N_473,In_778,In_860);
and U474 (N_474,In_168,In_426);
nor U475 (N_475,In_326,In_904);
nand U476 (N_476,In_637,In_475);
and U477 (N_477,In_225,In_588);
nor U478 (N_478,In_243,In_927);
nor U479 (N_479,In_154,In_551);
and U480 (N_480,In_910,In_466);
xnor U481 (N_481,In_6,In_110);
xor U482 (N_482,In_136,In_374);
and U483 (N_483,In_427,In_548);
nor U484 (N_484,In_83,In_589);
nand U485 (N_485,In_141,In_999);
nor U486 (N_486,In_577,In_167);
xor U487 (N_487,In_454,In_174);
nand U488 (N_488,In_227,In_823);
and U489 (N_489,In_262,In_563);
xnor U490 (N_490,In_451,In_468);
nand U491 (N_491,In_809,In_33);
nand U492 (N_492,In_247,In_84);
and U493 (N_493,In_542,In_758);
nand U494 (N_494,In_445,In_212);
or U495 (N_495,In_297,In_89);
xnor U496 (N_496,In_780,In_28);
or U497 (N_497,In_341,In_709);
or U498 (N_498,In_540,In_494);
or U499 (N_499,In_496,In_635);
xnor U500 (N_500,In_138,In_1);
nor U501 (N_501,In_289,In_683);
nor U502 (N_502,In_450,In_355);
nand U503 (N_503,In_83,In_439);
or U504 (N_504,In_255,In_860);
or U505 (N_505,In_377,In_788);
and U506 (N_506,In_883,In_932);
and U507 (N_507,In_937,In_175);
or U508 (N_508,In_631,In_994);
nand U509 (N_509,In_801,In_863);
nor U510 (N_510,In_911,In_60);
and U511 (N_511,In_991,In_154);
xnor U512 (N_512,In_325,In_664);
and U513 (N_513,In_694,In_539);
and U514 (N_514,In_827,In_976);
nand U515 (N_515,In_841,In_958);
nand U516 (N_516,In_114,In_75);
nor U517 (N_517,In_657,In_499);
and U518 (N_518,In_949,In_235);
and U519 (N_519,In_738,In_717);
or U520 (N_520,In_498,In_314);
nor U521 (N_521,In_547,In_879);
and U522 (N_522,In_924,In_294);
nor U523 (N_523,In_706,In_958);
xnor U524 (N_524,In_142,In_6);
and U525 (N_525,In_144,In_551);
and U526 (N_526,In_10,In_49);
or U527 (N_527,In_714,In_974);
or U528 (N_528,In_414,In_274);
nand U529 (N_529,In_132,In_798);
and U530 (N_530,In_613,In_322);
xnor U531 (N_531,In_157,In_98);
and U532 (N_532,In_826,In_894);
nand U533 (N_533,In_660,In_411);
nand U534 (N_534,In_99,In_254);
or U535 (N_535,In_774,In_318);
nand U536 (N_536,In_890,In_907);
xor U537 (N_537,In_217,In_775);
xnor U538 (N_538,In_971,In_604);
nor U539 (N_539,In_879,In_888);
or U540 (N_540,In_811,In_37);
nor U541 (N_541,In_474,In_839);
nand U542 (N_542,In_400,In_151);
or U543 (N_543,In_216,In_972);
xor U544 (N_544,In_757,In_989);
or U545 (N_545,In_529,In_172);
xor U546 (N_546,In_56,In_95);
nand U547 (N_547,In_559,In_658);
xor U548 (N_548,In_623,In_266);
and U549 (N_549,In_967,In_504);
nor U550 (N_550,In_902,In_675);
xor U551 (N_551,In_833,In_227);
nor U552 (N_552,In_667,In_195);
xor U553 (N_553,In_223,In_984);
xnor U554 (N_554,In_144,In_495);
nand U555 (N_555,In_393,In_866);
and U556 (N_556,In_623,In_511);
xnor U557 (N_557,In_274,In_433);
nand U558 (N_558,In_952,In_421);
and U559 (N_559,In_15,In_279);
or U560 (N_560,In_380,In_976);
and U561 (N_561,In_563,In_470);
and U562 (N_562,In_694,In_459);
nor U563 (N_563,In_136,In_833);
or U564 (N_564,In_839,In_729);
xnor U565 (N_565,In_823,In_768);
and U566 (N_566,In_754,In_651);
xor U567 (N_567,In_522,In_573);
nand U568 (N_568,In_270,In_371);
nor U569 (N_569,In_740,In_749);
nand U570 (N_570,In_712,In_847);
or U571 (N_571,In_748,In_204);
and U572 (N_572,In_632,In_988);
nor U573 (N_573,In_291,In_267);
and U574 (N_574,In_484,In_222);
or U575 (N_575,In_643,In_134);
nor U576 (N_576,In_7,In_756);
xnor U577 (N_577,In_867,In_28);
nand U578 (N_578,In_766,In_756);
and U579 (N_579,In_301,In_480);
and U580 (N_580,In_511,In_285);
nand U581 (N_581,In_176,In_791);
xnor U582 (N_582,In_100,In_670);
nand U583 (N_583,In_392,In_791);
and U584 (N_584,In_822,In_225);
nor U585 (N_585,In_52,In_265);
nor U586 (N_586,In_745,In_292);
xor U587 (N_587,In_41,In_347);
and U588 (N_588,In_431,In_919);
nor U589 (N_589,In_628,In_246);
and U590 (N_590,In_849,In_991);
nand U591 (N_591,In_707,In_570);
xnor U592 (N_592,In_781,In_33);
nand U593 (N_593,In_640,In_569);
nor U594 (N_594,In_749,In_656);
and U595 (N_595,In_77,In_297);
and U596 (N_596,In_491,In_908);
or U597 (N_597,In_212,In_321);
nand U598 (N_598,In_545,In_760);
nand U599 (N_599,In_271,In_549);
or U600 (N_600,In_804,In_658);
and U601 (N_601,In_162,In_965);
and U602 (N_602,In_785,In_437);
nand U603 (N_603,In_83,In_834);
xnor U604 (N_604,In_693,In_770);
nor U605 (N_605,In_82,In_389);
and U606 (N_606,In_652,In_456);
nand U607 (N_607,In_657,In_7);
and U608 (N_608,In_385,In_731);
and U609 (N_609,In_546,In_55);
nor U610 (N_610,In_424,In_153);
nor U611 (N_611,In_253,In_672);
nand U612 (N_612,In_133,In_794);
xor U613 (N_613,In_10,In_163);
or U614 (N_614,In_223,In_513);
nand U615 (N_615,In_385,In_248);
nor U616 (N_616,In_158,In_703);
or U617 (N_617,In_91,In_578);
nand U618 (N_618,In_276,In_742);
nor U619 (N_619,In_99,In_213);
nor U620 (N_620,In_323,In_904);
nor U621 (N_621,In_98,In_686);
nor U622 (N_622,In_685,In_571);
and U623 (N_623,In_803,In_656);
xnor U624 (N_624,In_878,In_300);
xnor U625 (N_625,In_721,In_972);
nor U626 (N_626,In_339,In_178);
nor U627 (N_627,In_185,In_574);
xor U628 (N_628,In_197,In_448);
and U629 (N_629,In_25,In_514);
nand U630 (N_630,In_350,In_77);
and U631 (N_631,In_160,In_562);
and U632 (N_632,In_763,In_175);
nand U633 (N_633,In_283,In_554);
nand U634 (N_634,In_307,In_397);
xnor U635 (N_635,In_471,In_392);
or U636 (N_636,In_899,In_814);
nor U637 (N_637,In_215,In_750);
and U638 (N_638,In_131,In_103);
and U639 (N_639,In_193,In_762);
nor U640 (N_640,In_363,In_102);
xnor U641 (N_641,In_852,In_316);
or U642 (N_642,In_629,In_841);
nor U643 (N_643,In_877,In_778);
or U644 (N_644,In_611,In_261);
nor U645 (N_645,In_170,In_609);
and U646 (N_646,In_738,In_353);
and U647 (N_647,In_791,In_345);
xnor U648 (N_648,In_651,In_881);
nor U649 (N_649,In_684,In_11);
or U650 (N_650,In_94,In_792);
nand U651 (N_651,In_871,In_253);
or U652 (N_652,In_832,In_735);
and U653 (N_653,In_614,In_554);
xor U654 (N_654,In_138,In_35);
or U655 (N_655,In_758,In_29);
nand U656 (N_656,In_81,In_71);
xor U657 (N_657,In_198,In_613);
nand U658 (N_658,In_94,In_364);
nor U659 (N_659,In_618,In_594);
or U660 (N_660,In_354,In_518);
nand U661 (N_661,In_478,In_473);
nand U662 (N_662,In_151,In_757);
xnor U663 (N_663,In_68,In_992);
and U664 (N_664,In_381,In_739);
nand U665 (N_665,In_587,In_35);
nor U666 (N_666,In_756,In_602);
nor U667 (N_667,In_936,In_674);
nor U668 (N_668,In_97,In_730);
and U669 (N_669,In_35,In_401);
and U670 (N_670,In_285,In_186);
nor U671 (N_671,In_956,In_26);
nand U672 (N_672,In_928,In_306);
nor U673 (N_673,In_557,In_852);
nor U674 (N_674,In_391,In_159);
and U675 (N_675,In_219,In_960);
nand U676 (N_676,In_430,In_422);
or U677 (N_677,In_752,In_87);
nor U678 (N_678,In_351,In_90);
nor U679 (N_679,In_932,In_760);
or U680 (N_680,In_127,In_156);
xor U681 (N_681,In_861,In_993);
nand U682 (N_682,In_271,In_547);
nand U683 (N_683,In_554,In_820);
nor U684 (N_684,In_176,In_566);
and U685 (N_685,In_6,In_378);
and U686 (N_686,In_910,In_552);
nor U687 (N_687,In_59,In_712);
xor U688 (N_688,In_696,In_38);
xnor U689 (N_689,In_603,In_412);
nor U690 (N_690,In_758,In_903);
xnor U691 (N_691,In_626,In_687);
nor U692 (N_692,In_884,In_358);
nor U693 (N_693,In_292,In_459);
and U694 (N_694,In_491,In_639);
xnor U695 (N_695,In_991,In_579);
xor U696 (N_696,In_824,In_284);
xnor U697 (N_697,In_671,In_730);
xnor U698 (N_698,In_648,In_346);
and U699 (N_699,In_507,In_620);
and U700 (N_700,In_562,In_630);
or U701 (N_701,In_718,In_962);
xnor U702 (N_702,In_102,In_765);
nor U703 (N_703,In_533,In_808);
and U704 (N_704,In_334,In_801);
nor U705 (N_705,In_798,In_596);
and U706 (N_706,In_133,In_846);
nand U707 (N_707,In_559,In_16);
nor U708 (N_708,In_703,In_225);
nor U709 (N_709,In_849,In_833);
and U710 (N_710,In_721,In_122);
and U711 (N_711,In_439,In_424);
nor U712 (N_712,In_956,In_649);
xnor U713 (N_713,In_161,In_982);
xor U714 (N_714,In_739,In_201);
or U715 (N_715,In_277,In_910);
nand U716 (N_716,In_84,In_357);
nor U717 (N_717,In_399,In_449);
nand U718 (N_718,In_437,In_548);
nor U719 (N_719,In_190,In_48);
nand U720 (N_720,In_775,In_102);
and U721 (N_721,In_507,In_964);
xor U722 (N_722,In_39,In_334);
nand U723 (N_723,In_165,In_595);
xnor U724 (N_724,In_929,In_82);
or U725 (N_725,In_208,In_206);
xnor U726 (N_726,In_448,In_900);
nand U727 (N_727,In_143,In_850);
nand U728 (N_728,In_311,In_316);
and U729 (N_729,In_154,In_379);
nand U730 (N_730,In_903,In_975);
nand U731 (N_731,In_910,In_558);
nand U732 (N_732,In_538,In_273);
nor U733 (N_733,In_709,In_291);
xnor U734 (N_734,In_690,In_461);
and U735 (N_735,In_887,In_643);
and U736 (N_736,In_104,In_357);
nand U737 (N_737,In_194,In_211);
and U738 (N_738,In_627,In_830);
or U739 (N_739,In_514,In_103);
or U740 (N_740,In_565,In_48);
or U741 (N_741,In_891,In_662);
xor U742 (N_742,In_937,In_371);
nand U743 (N_743,In_592,In_470);
nand U744 (N_744,In_589,In_345);
xnor U745 (N_745,In_703,In_924);
xnor U746 (N_746,In_546,In_970);
nor U747 (N_747,In_288,In_651);
or U748 (N_748,In_150,In_703);
xnor U749 (N_749,In_228,In_142);
or U750 (N_750,In_374,In_148);
xor U751 (N_751,In_134,In_857);
or U752 (N_752,In_352,In_525);
nor U753 (N_753,In_298,In_807);
nor U754 (N_754,In_790,In_142);
xor U755 (N_755,In_522,In_209);
and U756 (N_756,In_859,In_468);
xor U757 (N_757,In_894,In_604);
or U758 (N_758,In_658,In_938);
xor U759 (N_759,In_142,In_920);
and U760 (N_760,In_372,In_607);
nand U761 (N_761,In_801,In_715);
xor U762 (N_762,In_189,In_22);
nor U763 (N_763,In_730,In_652);
and U764 (N_764,In_269,In_615);
nand U765 (N_765,In_319,In_698);
nor U766 (N_766,In_834,In_305);
nand U767 (N_767,In_456,In_880);
nand U768 (N_768,In_977,In_334);
or U769 (N_769,In_699,In_613);
and U770 (N_770,In_897,In_802);
nand U771 (N_771,In_294,In_779);
xor U772 (N_772,In_545,In_500);
nor U773 (N_773,In_687,In_783);
xor U774 (N_774,In_39,In_831);
xnor U775 (N_775,In_480,In_14);
nand U776 (N_776,In_242,In_327);
xor U777 (N_777,In_854,In_837);
nand U778 (N_778,In_1,In_525);
xnor U779 (N_779,In_196,In_426);
or U780 (N_780,In_513,In_987);
nor U781 (N_781,In_124,In_378);
and U782 (N_782,In_587,In_801);
nor U783 (N_783,In_304,In_45);
nor U784 (N_784,In_254,In_173);
and U785 (N_785,In_10,In_404);
xnor U786 (N_786,In_122,In_935);
and U787 (N_787,In_641,In_420);
or U788 (N_788,In_708,In_718);
nor U789 (N_789,In_813,In_412);
nand U790 (N_790,In_848,In_434);
nor U791 (N_791,In_326,In_906);
and U792 (N_792,In_287,In_821);
and U793 (N_793,In_650,In_375);
or U794 (N_794,In_862,In_353);
xor U795 (N_795,In_67,In_288);
or U796 (N_796,In_834,In_220);
nor U797 (N_797,In_345,In_92);
xnor U798 (N_798,In_479,In_806);
nand U799 (N_799,In_116,In_796);
and U800 (N_800,In_864,In_872);
or U801 (N_801,In_611,In_811);
or U802 (N_802,In_714,In_493);
nor U803 (N_803,In_913,In_909);
xor U804 (N_804,In_356,In_700);
and U805 (N_805,In_267,In_574);
and U806 (N_806,In_337,In_520);
and U807 (N_807,In_586,In_463);
xnor U808 (N_808,In_84,In_696);
and U809 (N_809,In_688,In_204);
or U810 (N_810,In_306,In_942);
and U811 (N_811,In_862,In_344);
nand U812 (N_812,In_653,In_159);
or U813 (N_813,In_863,In_137);
nor U814 (N_814,In_71,In_434);
or U815 (N_815,In_461,In_448);
xor U816 (N_816,In_895,In_387);
nand U817 (N_817,In_918,In_608);
nor U818 (N_818,In_107,In_512);
or U819 (N_819,In_700,In_540);
or U820 (N_820,In_252,In_74);
xor U821 (N_821,In_39,In_824);
nand U822 (N_822,In_488,In_417);
nor U823 (N_823,In_292,In_885);
or U824 (N_824,In_546,In_451);
or U825 (N_825,In_553,In_328);
nor U826 (N_826,In_740,In_823);
xnor U827 (N_827,In_101,In_221);
and U828 (N_828,In_553,In_816);
xnor U829 (N_829,In_430,In_605);
or U830 (N_830,In_117,In_321);
xor U831 (N_831,In_87,In_217);
nor U832 (N_832,In_955,In_814);
or U833 (N_833,In_613,In_829);
or U834 (N_834,In_102,In_565);
or U835 (N_835,In_915,In_887);
and U836 (N_836,In_991,In_929);
xnor U837 (N_837,In_146,In_678);
nor U838 (N_838,In_853,In_200);
nand U839 (N_839,In_398,In_232);
or U840 (N_840,In_335,In_104);
nor U841 (N_841,In_512,In_717);
or U842 (N_842,In_885,In_419);
or U843 (N_843,In_98,In_806);
and U844 (N_844,In_441,In_419);
xor U845 (N_845,In_69,In_558);
or U846 (N_846,In_450,In_796);
and U847 (N_847,In_48,In_961);
xnor U848 (N_848,In_506,In_996);
or U849 (N_849,In_733,In_520);
xnor U850 (N_850,In_768,In_561);
nor U851 (N_851,In_983,In_838);
or U852 (N_852,In_891,In_304);
xor U853 (N_853,In_126,In_328);
nor U854 (N_854,In_489,In_20);
nor U855 (N_855,In_673,In_326);
nor U856 (N_856,In_902,In_152);
xor U857 (N_857,In_194,In_39);
nor U858 (N_858,In_360,In_851);
nand U859 (N_859,In_831,In_311);
and U860 (N_860,In_351,In_921);
or U861 (N_861,In_299,In_5);
xor U862 (N_862,In_477,In_685);
nor U863 (N_863,In_941,In_166);
or U864 (N_864,In_688,In_641);
nor U865 (N_865,In_509,In_380);
nor U866 (N_866,In_79,In_147);
xor U867 (N_867,In_200,In_791);
nand U868 (N_868,In_38,In_812);
nor U869 (N_869,In_644,In_994);
xor U870 (N_870,In_533,In_316);
or U871 (N_871,In_320,In_587);
xnor U872 (N_872,In_346,In_795);
nand U873 (N_873,In_779,In_244);
nor U874 (N_874,In_91,In_707);
or U875 (N_875,In_335,In_582);
xnor U876 (N_876,In_157,In_797);
nor U877 (N_877,In_833,In_284);
xnor U878 (N_878,In_603,In_472);
or U879 (N_879,In_727,In_669);
or U880 (N_880,In_601,In_133);
xnor U881 (N_881,In_301,In_374);
nand U882 (N_882,In_881,In_920);
and U883 (N_883,In_104,In_216);
xor U884 (N_884,In_408,In_656);
and U885 (N_885,In_19,In_889);
nand U886 (N_886,In_847,In_532);
and U887 (N_887,In_901,In_141);
and U888 (N_888,In_36,In_402);
or U889 (N_889,In_913,In_728);
nand U890 (N_890,In_612,In_978);
nand U891 (N_891,In_340,In_990);
and U892 (N_892,In_762,In_918);
or U893 (N_893,In_769,In_575);
nand U894 (N_894,In_781,In_382);
or U895 (N_895,In_208,In_534);
and U896 (N_896,In_257,In_851);
nand U897 (N_897,In_913,In_24);
nand U898 (N_898,In_212,In_640);
nor U899 (N_899,In_756,In_116);
nor U900 (N_900,In_628,In_701);
nand U901 (N_901,In_226,In_511);
or U902 (N_902,In_473,In_286);
xnor U903 (N_903,In_390,In_255);
xor U904 (N_904,In_952,In_436);
nand U905 (N_905,In_566,In_898);
nor U906 (N_906,In_32,In_653);
nand U907 (N_907,In_768,In_412);
nor U908 (N_908,In_13,In_202);
or U909 (N_909,In_613,In_924);
xnor U910 (N_910,In_507,In_807);
and U911 (N_911,In_535,In_462);
nor U912 (N_912,In_413,In_802);
nand U913 (N_913,In_838,In_766);
and U914 (N_914,In_80,In_982);
or U915 (N_915,In_907,In_806);
nand U916 (N_916,In_982,In_91);
nor U917 (N_917,In_717,In_870);
or U918 (N_918,In_808,In_570);
xor U919 (N_919,In_188,In_377);
nand U920 (N_920,In_13,In_509);
nor U921 (N_921,In_415,In_75);
nor U922 (N_922,In_106,In_338);
nor U923 (N_923,In_294,In_791);
and U924 (N_924,In_470,In_600);
and U925 (N_925,In_438,In_345);
nor U926 (N_926,In_431,In_508);
xnor U927 (N_927,In_133,In_359);
xor U928 (N_928,In_228,In_668);
and U929 (N_929,In_710,In_386);
and U930 (N_930,In_206,In_268);
and U931 (N_931,In_911,In_789);
or U932 (N_932,In_610,In_596);
or U933 (N_933,In_110,In_197);
xor U934 (N_934,In_594,In_664);
xnor U935 (N_935,In_467,In_929);
nand U936 (N_936,In_54,In_352);
or U937 (N_937,In_544,In_81);
or U938 (N_938,In_884,In_545);
and U939 (N_939,In_164,In_742);
nor U940 (N_940,In_376,In_908);
nand U941 (N_941,In_29,In_984);
and U942 (N_942,In_629,In_21);
nor U943 (N_943,In_863,In_477);
and U944 (N_944,In_666,In_641);
or U945 (N_945,In_877,In_298);
and U946 (N_946,In_477,In_201);
nor U947 (N_947,In_91,In_669);
nor U948 (N_948,In_808,In_573);
nand U949 (N_949,In_430,In_862);
and U950 (N_950,In_191,In_672);
nor U951 (N_951,In_739,In_141);
and U952 (N_952,In_293,In_333);
or U953 (N_953,In_894,In_321);
and U954 (N_954,In_887,In_691);
and U955 (N_955,In_522,In_849);
xor U956 (N_956,In_415,In_249);
or U957 (N_957,In_348,In_473);
nor U958 (N_958,In_626,In_917);
or U959 (N_959,In_226,In_308);
or U960 (N_960,In_26,In_872);
xor U961 (N_961,In_561,In_989);
nand U962 (N_962,In_566,In_885);
xor U963 (N_963,In_278,In_223);
nand U964 (N_964,In_363,In_549);
and U965 (N_965,In_601,In_791);
nand U966 (N_966,In_662,In_525);
and U967 (N_967,In_853,In_89);
xnor U968 (N_968,In_180,In_387);
nand U969 (N_969,In_155,In_499);
or U970 (N_970,In_159,In_411);
nor U971 (N_971,In_791,In_521);
or U972 (N_972,In_806,In_117);
nor U973 (N_973,In_445,In_397);
nor U974 (N_974,In_901,In_568);
and U975 (N_975,In_428,In_845);
nor U976 (N_976,In_158,In_743);
nand U977 (N_977,In_674,In_709);
xor U978 (N_978,In_43,In_858);
xnor U979 (N_979,In_397,In_1);
xnor U980 (N_980,In_908,In_776);
nand U981 (N_981,In_363,In_109);
nand U982 (N_982,In_122,In_296);
xnor U983 (N_983,In_610,In_186);
xor U984 (N_984,In_55,In_920);
nor U985 (N_985,In_774,In_870);
nor U986 (N_986,In_94,In_655);
or U987 (N_987,In_229,In_69);
xnor U988 (N_988,In_994,In_960);
xnor U989 (N_989,In_386,In_415);
and U990 (N_990,In_145,In_152);
or U991 (N_991,In_63,In_190);
and U992 (N_992,In_184,In_273);
nand U993 (N_993,In_971,In_202);
or U994 (N_994,In_584,In_859);
nor U995 (N_995,In_238,In_48);
and U996 (N_996,In_724,In_332);
nand U997 (N_997,In_124,In_732);
or U998 (N_998,In_374,In_720);
nand U999 (N_999,In_832,In_146);
nand U1000 (N_1000,In_515,In_806);
or U1001 (N_1001,In_914,In_373);
xor U1002 (N_1002,In_241,In_56);
nor U1003 (N_1003,In_848,In_716);
and U1004 (N_1004,In_593,In_288);
or U1005 (N_1005,In_220,In_922);
or U1006 (N_1006,In_125,In_272);
or U1007 (N_1007,In_339,In_869);
and U1008 (N_1008,In_162,In_459);
or U1009 (N_1009,In_938,In_206);
or U1010 (N_1010,In_625,In_76);
or U1011 (N_1011,In_279,In_703);
nand U1012 (N_1012,In_487,In_772);
or U1013 (N_1013,In_530,In_575);
and U1014 (N_1014,In_447,In_750);
or U1015 (N_1015,In_211,In_133);
and U1016 (N_1016,In_216,In_959);
or U1017 (N_1017,In_287,In_540);
or U1018 (N_1018,In_103,In_613);
or U1019 (N_1019,In_534,In_825);
or U1020 (N_1020,In_520,In_344);
nand U1021 (N_1021,In_143,In_322);
nand U1022 (N_1022,In_312,In_710);
xor U1023 (N_1023,In_875,In_26);
xor U1024 (N_1024,In_827,In_194);
and U1025 (N_1025,In_562,In_264);
xnor U1026 (N_1026,In_82,In_373);
or U1027 (N_1027,In_141,In_121);
xor U1028 (N_1028,In_654,In_398);
nand U1029 (N_1029,In_299,In_200);
nor U1030 (N_1030,In_425,In_205);
and U1031 (N_1031,In_899,In_709);
or U1032 (N_1032,In_208,In_758);
xnor U1033 (N_1033,In_372,In_157);
nand U1034 (N_1034,In_456,In_857);
nor U1035 (N_1035,In_56,In_274);
xor U1036 (N_1036,In_627,In_868);
nor U1037 (N_1037,In_814,In_94);
nand U1038 (N_1038,In_724,In_345);
or U1039 (N_1039,In_47,In_536);
or U1040 (N_1040,In_592,In_746);
nand U1041 (N_1041,In_544,In_908);
nor U1042 (N_1042,In_814,In_448);
and U1043 (N_1043,In_37,In_360);
nand U1044 (N_1044,In_332,In_776);
or U1045 (N_1045,In_780,In_510);
nand U1046 (N_1046,In_171,In_142);
and U1047 (N_1047,In_407,In_547);
nor U1048 (N_1048,In_515,In_110);
or U1049 (N_1049,In_575,In_44);
xnor U1050 (N_1050,In_33,In_62);
nor U1051 (N_1051,In_478,In_633);
nand U1052 (N_1052,In_255,In_811);
or U1053 (N_1053,In_785,In_922);
xor U1054 (N_1054,In_875,In_550);
xnor U1055 (N_1055,In_881,In_412);
xnor U1056 (N_1056,In_961,In_361);
or U1057 (N_1057,In_966,In_275);
nor U1058 (N_1058,In_489,In_101);
or U1059 (N_1059,In_562,In_417);
xnor U1060 (N_1060,In_203,In_882);
nor U1061 (N_1061,In_539,In_426);
and U1062 (N_1062,In_891,In_452);
xnor U1063 (N_1063,In_268,In_477);
nor U1064 (N_1064,In_944,In_821);
or U1065 (N_1065,In_421,In_726);
nand U1066 (N_1066,In_701,In_472);
and U1067 (N_1067,In_625,In_444);
nor U1068 (N_1068,In_159,In_155);
nor U1069 (N_1069,In_777,In_561);
and U1070 (N_1070,In_442,In_161);
nand U1071 (N_1071,In_61,In_295);
or U1072 (N_1072,In_174,In_665);
nand U1073 (N_1073,In_501,In_404);
nand U1074 (N_1074,In_368,In_613);
nor U1075 (N_1075,In_187,In_160);
and U1076 (N_1076,In_95,In_268);
xor U1077 (N_1077,In_363,In_226);
and U1078 (N_1078,In_556,In_483);
nor U1079 (N_1079,In_694,In_831);
nand U1080 (N_1080,In_43,In_226);
xor U1081 (N_1081,In_615,In_95);
and U1082 (N_1082,In_654,In_59);
nor U1083 (N_1083,In_113,In_896);
and U1084 (N_1084,In_632,In_556);
or U1085 (N_1085,In_750,In_348);
xor U1086 (N_1086,In_13,In_451);
nand U1087 (N_1087,In_167,In_46);
and U1088 (N_1088,In_682,In_544);
or U1089 (N_1089,In_839,In_83);
and U1090 (N_1090,In_355,In_642);
or U1091 (N_1091,In_913,In_259);
nor U1092 (N_1092,In_527,In_127);
or U1093 (N_1093,In_593,In_860);
or U1094 (N_1094,In_363,In_665);
or U1095 (N_1095,In_954,In_733);
nor U1096 (N_1096,In_149,In_768);
nor U1097 (N_1097,In_88,In_840);
nand U1098 (N_1098,In_90,In_489);
xor U1099 (N_1099,In_330,In_553);
nor U1100 (N_1100,In_412,In_171);
and U1101 (N_1101,In_264,In_563);
nor U1102 (N_1102,In_641,In_876);
or U1103 (N_1103,In_367,In_658);
and U1104 (N_1104,In_205,In_524);
nor U1105 (N_1105,In_635,In_525);
xor U1106 (N_1106,In_459,In_97);
nand U1107 (N_1107,In_560,In_913);
and U1108 (N_1108,In_743,In_469);
xnor U1109 (N_1109,In_430,In_916);
nand U1110 (N_1110,In_57,In_293);
or U1111 (N_1111,In_922,In_672);
and U1112 (N_1112,In_74,In_438);
nand U1113 (N_1113,In_741,In_200);
nand U1114 (N_1114,In_505,In_237);
or U1115 (N_1115,In_663,In_67);
nand U1116 (N_1116,In_923,In_355);
xor U1117 (N_1117,In_675,In_756);
or U1118 (N_1118,In_747,In_993);
or U1119 (N_1119,In_892,In_120);
nor U1120 (N_1120,In_287,In_526);
nand U1121 (N_1121,In_725,In_514);
and U1122 (N_1122,In_38,In_673);
nor U1123 (N_1123,In_247,In_757);
xnor U1124 (N_1124,In_824,In_906);
xor U1125 (N_1125,In_810,In_160);
xor U1126 (N_1126,In_779,In_259);
or U1127 (N_1127,In_131,In_58);
nor U1128 (N_1128,In_394,In_552);
or U1129 (N_1129,In_762,In_572);
or U1130 (N_1130,In_907,In_551);
or U1131 (N_1131,In_289,In_503);
and U1132 (N_1132,In_658,In_333);
xor U1133 (N_1133,In_185,In_93);
or U1134 (N_1134,In_284,In_337);
nand U1135 (N_1135,In_742,In_799);
xor U1136 (N_1136,In_830,In_814);
xnor U1137 (N_1137,In_890,In_214);
nor U1138 (N_1138,In_170,In_625);
nor U1139 (N_1139,In_864,In_422);
and U1140 (N_1140,In_471,In_719);
nand U1141 (N_1141,In_582,In_631);
or U1142 (N_1142,In_166,In_330);
and U1143 (N_1143,In_540,In_285);
or U1144 (N_1144,In_574,In_649);
and U1145 (N_1145,In_100,In_947);
and U1146 (N_1146,In_645,In_970);
nand U1147 (N_1147,In_339,In_878);
nand U1148 (N_1148,In_450,In_673);
and U1149 (N_1149,In_196,In_736);
xor U1150 (N_1150,In_144,In_964);
or U1151 (N_1151,In_191,In_305);
nor U1152 (N_1152,In_883,In_846);
or U1153 (N_1153,In_578,In_296);
nand U1154 (N_1154,In_9,In_744);
nand U1155 (N_1155,In_899,In_760);
and U1156 (N_1156,In_858,In_114);
and U1157 (N_1157,In_630,In_53);
and U1158 (N_1158,In_871,In_218);
and U1159 (N_1159,In_816,In_775);
xor U1160 (N_1160,In_395,In_545);
or U1161 (N_1161,In_521,In_568);
nand U1162 (N_1162,In_97,In_747);
nand U1163 (N_1163,In_749,In_829);
xor U1164 (N_1164,In_189,In_196);
and U1165 (N_1165,In_93,In_676);
and U1166 (N_1166,In_584,In_858);
xnor U1167 (N_1167,In_267,In_628);
nor U1168 (N_1168,In_858,In_933);
nand U1169 (N_1169,In_746,In_155);
or U1170 (N_1170,In_779,In_339);
nor U1171 (N_1171,In_831,In_994);
or U1172 (N_1172,In_731,In_375);
or U1173 (N_1173,In_298,In_895);
xor U1174 (N_1174,In_524,In_943);
and U1175 (N_1175,In_952,In_343);
nand U1176 (N_1176,In_171,In_202);
xor U1177 (N_1177,In_663,In_516);
and U1178 (N_1178,In_353,In_156);
nor U1179 (N_1179,In_31,In_51);
nand U1180 (N_1180,In_622,In_980);
xor U1181 (N_1181,In_367,In_279);
or U1182 (N_1182,In_55,In_75);
nor U1183 (N_1183,In_282,In_453);
and U1184 (N_1184,In_89,In_280);
nor U1185 (N_1185,In_922,In_764);
and U1186 (N_1186,In_322,In_956);
and U1187 (N_1187,In_808,In_180);
xor U1188 (N_1188,In_420,In_430);
xor U1189 (N_1189,In_981,In_114);
and U1190 (N_1190,In_332,In_82);
xor U1191 (N_1191,In_698,In_9);
and U1192 (N_1192,In_543,In_445);
nand U1193 (N_1193,In_128,In_137);
nand U1194 (N_1194,In_204,In_413);
nand U1195 (N_1195,In_230,In_819);
nand U1196 (N_1196,In_936,In_399);
nor U1197 (N_1197,In_345,In_487);
xor U1198 (N_1198,In_566,In_586);
and U1199 (N_1199,In_544,In_889);
or U1200 (N_1200,In_451,In_737);
and U1201 (N_1201,In_162,In_848);
nand U1202 (N_1202,In_501,In_418);
nand U1203 (N_1203,In_485,In_178);
nand U1204 (N_1204,In_774,In_717);
nor U1205 (N_1205,In_788,In_968);
nand U1206 (N_1206,In_915,In_622);
and U1207 (N_1207,In_7,In_846);
nor U1208 (N_1208,In_867,In_954);
or U1209 (N_1209,In_382,In_73);
nor U1210 (N_1210,In_383,In_559);
or U1211 (N_1211,In_25,In_982);
nand U1212 (N_1212,In_49,In_166);
or U1213 (N_1213,In_467,In_666);
nor U1214 (N_1214,In_371,In_0);
or U1215 (N_1215,In_869,In_419);
xor U1216 (N_1216,In_834,In_731);
xnor U1217 (N_1217,In_242,In_925);
xnor U1218 (N_1218,In_732,In_191);
xnor U1219 (N_1219,In_598,In_141);
nor U1220 (N_1220,In_325,In_903);
xnor U1221 (N_1221,In_90,In_427);
nor U1222 (N_1222,In_71,In_299);
nor U1223 (N_1223,In_623,In_668);
and U1224 (N_1224,In_56,In_922);
and U1225 (N_1225,In_72,In_514);
xnor U1226 (N_1226,In_48,In_631);
or U1227 (N_1227,In_388,In_91);
and U1228 (N_1228,In_972,In_882);
nor U1229 (N_1229,In_539,In_244);
nor U1230 (N_1230,In_907,In_437);
or U1231 (N_1231,In_235,In_597);
and U1232 (N_1232,In_703,In_817);
xnor U1233 (N_1233,In_860,In_67);
nor U1234 (N_1234,In_175,In_558);
nand U1235 (N_1235,In_20,In_759);
or U1236 (N_1236,In_202,In_655);
nor U1237 (N_1237,In_623,In_480);
or U1238 (N_1238,In_652,In_957);
xnor U1239 (N_1239,In_871,In_402);
nor U1240 (N_1240,In_671,In_160);
nand U1241 (N_1241,In_217,In_365);
nand U1242 (N_1242,In_647,In_953);
and U1243 (N_1243,In_81,In_28);
nor U1244 (N_1244,In_455,In_355);
nand U1245 (N_1245,In_305,In_718);
or U1246 (N_1246,In_34,In_3);
and U1247 (N_1247,In_601,In_746);
nor U1248 (N_1248,In_963,In_718);
nor U1249 (N_1249,In_111,In_788);
xnor U1250 (N_1250,In_334,In_382);
and U1251 (N_1251,In_346,In_400);
or U1252 (N_1252,In_661,In_156);
nand U1253 (N_1253,In_71,In_876);
or U1254 (N_1254,In_539,In_189);
nand U1255 (N_1255,In_356,In_569);
and U1256 (N_1256,In_591,In_962);
and U1257 (N_1257,In_666,In_608);
and U1258 (N_1258,In_774,In_537);
or U1259 (N_1259,In_142,In_992);
nand U1260 (N_1260,In_211,In_86);
xnor U1261 (N_1261,In_738,In_864);
or U1262 (N_1262,In_670,In_479);
or U1263 (N_1263,In_984,In_842);
or U1264 (N_1264,In_572,In_839);
or U1265 (N_1265,In_618,In_530);
and U1266 (N_1266,In_92,In_209);
nor U1267 (N_1267,In_986,In_403);
xor U1268 (N_1268,In_376,In_681);
xnor U1269 (N_1269,In_988,In_292);
nand U1270 (N_1270,In_83,In_504);
nand U1271 (N_1271,In_221,In_384);
nand U1272 (N_1272,In_832,In_948);
nand U1273 (N_1273,In_502,In_899);
xor U1274 (N_1274,In_665,In_857);
xnor U1275 (N_1275,In_104,In_484);
or U1276 (N_1276,In_525,In_953);
and U1277 (N_1277,In_323,In_352);
nand U1278 (N_1278,In_151,In_693);
or U1279 (N_1279,In_192,In_255);
nand U1280 (N_1280,In_467,In_179);
nand U1281 (N_1281,In_29,In_389);
xnor U1282 (N_1282,In_331,In_258);
nor U1283 (N_1283,In_324,In_38);
and U1284 (N_1284,In_510,In_257);
nand U1285 (N_1285,In_780,In_639);
xnor U1286 (N_1286,In_222,In_201);
nand U1287 (N_1287,In_285,In_323);
nor U1288 (N_1288,In_814,In_191);
and U1289 (N_1289,In_270,In_540);
nand U1290 (N_1290,In_704,In_354);
xnor U1291 (N_1291,In_963,In_379);
nand U1292 (N_1292,In_286,In_99);
xor U1293 (N_1293,In_605,In_65);
or U1294 (N_1294,In_101,In_814);
nand U1295 (N_1295,In_918,In_936);
or U1296 (N_1296,In_413,In_466);
nor U1297 (N_1297,In_822,In_424);
xor U1298 (N_1298,In_790,In_795);
and U1299 (N_1299,In_749,In_354);
nand U1300 (N_1300,In_880,In_887);
nand U1301 (N_1301,In_560,In_73);
nand U1302 (N_1302,In_673,In_961);
nor U1303 (N_1303,In_941,In_608);
nand U1304 (N_1304,In_830,In_578);
xnor U1305 (N_1305,In_121,In_510);
or U1306 (N_1306,In_202,In_684);
xor U1307 (N_1307,In_184,In_24);
nor U1308 (N_1308,In_816,In_954);
nand U1309 (N_1309,In_526,In_185);
xor U1310 (N_1310,In_458,In_554);
or U1311 (N_1311,In_485,In_435);
and U1312 (N_1312,In_816,In_866);
nor U1313 (N_1313,In_986,In_326);
or U1314 (N_1314,In_815,In_74);
nand U1315 (N_1315,In_246,In_577);
and U1316 (N_1316,In_242,In_236);
xor U1317 (N_1317,In_819,In_925);
nor U1318 (N_1318,In_476,In_968);
or U1319 (N_1319,In_148,In_74);
or U1320 (N_1320,In_349,In_160);
and U1321 (N_1321,In_734,In_782);
nor U1322 (N_1322,In_519,In_319);
and U1323 (N_1323,In_883,In_720);
and U1324 (N_1324,In_557,In_444);
and U1325 (N_1325,In_357,In_838);
nand U1326 (N_1326,In_270,In_106);
nand U1327 (N_1327,In_701,In_22);
nor U1328 (N_1328,In_934,In_472);
xor U1329 (N_1329,In_935,In_984);
nand U1330 (N_1330,In_246,In_651);
nand U1331 (N_1331,In_54,In_459);
or U1332 (N_1332,In_762,In_652);
nor U1333 (N_1333,In_930,In_855);
xnor U1334 (N_1334,In_625,In_715);
xnor U1335 (N_1335,In_223,In_41);
and U1336 (N_1336,In_136,In_803);
nor U1337 (N_1337,In_729,In_243);
and U1338 (N_1338,In_774,In_593);
nor U1339 (N_1339,In_583,In_809);
nand U1340 (N_1340,In_940,In_540);
and U1341 (N_1341,In_141,In_85);
or U1342 (N_1342,In_508,In_524);
and U1343 (N_1343,In_617,In_191);
and U1344 (N_1344,In_666,In_490);
nand U1345 (N_1345,In_614,In_106);
nand U1346 (N_1346,In_847,In_264);
nor U1347 (N_1347,In_369,In_818);
nor U1348 (N_1348,In_991,In_27);
nor U1349 (N_1349,In_643,In_390);
nor U1350 (N_1350,In_913,In_609);
xor U1351 (N_1351,In_118,In_840);
nand U1352 (N_1352,In_417,In_622);
and U1353 (N_1353,In_184,In_962);
xor U1354 (N_1354,In_167,In_142);
nand U1355 (N_1355,In_675,In_989);
xor U1356 (N_1356,In_412,In_336);
xor U1357 (N_1357,In_9,In_332);
nand U1358 (N_1358,In_617,In_749);
nor U1359 (N_1359,In_541,In_682);
xor U1360 (N_1360,In_189,In_424);
nand U1361 (N_1361,In_359,In_949);
or U1362 (N_1362,In_146,In_129);
nand U1363 (N_1363,In_67,In_821);
nor U1364 (N_1364,In_547,In_507);
and U1365 (N_1365,In_81,In_578);
and U1366 (N_1366,In_306,In_980);
xnor U1367 (N_1367,In_156,In_22);
nor U1368 (N_1368,In_474,In_199);
nor U1369 (N_1369,In_957,In_936);
xnor U1370 (N_1370,In_158,In_282);
and U1371 (N_1371,In_389,In_949);
or U1372 (N_1372,In_940,In_653);
nor U1373 (N_1373,In_137,In_805);
nand U1374 (N_1374,In_54,In_722);
or U1375 (N_1375,In_408,In_362);
or U1376 (N_1376,In_275,In_572);
and U1377 (N_1377,In_10,In_678);
or U1378 (N_1378,In_50,In_641);
or U1379 (N_1379,In_618,In_152);
xor U1380 (N_1380,In_979,In_890);
xnor U1381 (N_1381,In_616,In_909);
and U1382 (N_1382,In_468,In_85);
xor U1383 (N_1383,In_673,In_302);
xor U1384 (N_1384,In_420,In_144);
and U1385 (N_1385,In_99,In_344);
or U1386 (N_1386,In_310,In_928);
nand U1387 (N_1387,In_155,In_883);
and U1388 (N_1388,In_858,In_739);
nand U1389 (N_1389,In_926,In_546);
xor U1390 (N_1390,In_124,In_924);
and U1391 (N_1391,In_543,In_943);
nand U1392 (N_1392,In_766,In_221);
nor U1393 (N_1393,In_410,In_666);
nand U1394 (N_1394,In_972,In_580);
nand U1395 (N_1395,In_878,In_827);
or U1396 (N_1396,In_55,In_942);
nor U1397 (N_1397,In_10,In_849);
or U1398 (N_1398,In_231,In_610);
and U1399 (N_1399,In_673,In_180);
xnor U1400 (N_1400,In_136,In_161);
nand U1401 (N_1401,In_464,In_13);
xor U1402 (N_1402,In_923,In_492);
nor U1403 (N_1403,In_619,In_329);
or U1404 (N_1404,In_781,In_616);
nand U1405 (N_1405,In_907,In_970);
xnor U1406 (N_1406,In_926,In_818);
and U1407 (N_1407,In_94,In_217);
or U1408 (N_1408,In_507,In_474);
and U1409 (N_1409,In_100,In_538);
and U1410 (N_1410,In_278,In_902);
nor U1411 (N_1411,In_795,In_379);
nand U1412 (N_1412,In_499,In_229);
nand U1413 (N_1413,In_115,In_417);
xor U1414 (N_1414,In_839,In_643);
nor U1415 (N_1415,In_757,In_311);
nand U1416 (N_1416,In_7,In_615);
or U1417 (N_1417,In_150,In_922);
and U1418 (N_1418,In_694,In_857);
and U1419 (N_1419,In_448,In_87);
xor U1420 (N_1420,In_568,In_345);
or U1421 (N_1421,In_161,In_531);
or U1422 (N_1422,In_843,In_329);
and U1423 (N_1423,In_993,In_532);
xor U1424 (N_1424,In_129,In_528);
xnor U1425 (N_1425,In_102,In_487);
xnor U1426 (N_1426,In_869,In_381);
or U1427 (N_1427,In_566,In_997);
and U1428 (N_1428,In_256,In_893);
nand U1429 (N_1429,In_534,In_807);
or U1430 (N_1430,In_983,In_981);
nor U1431 (N_1431,In_506,In_166);
or U1432 (N_1432,In_78,In_350);
nand U1433 (N_1433,In_193,In_931);
nand U1434 (N_1434,In_431,In_312);
and U1435 (N_1435,In_225,In_853);
nand U1436 (N_1436,In_25,In_659);
or U1437 (N_1437,In_543,In_577);
and U1438 (N_1438,In_92,In_970);
nor U1439 (N_1439,In_464,In_615);
or U1440 (N_1440,In_863,In_531);
and U1441 (N_1441,In_249,In_220);
xnor U1442 (N_1442,In_518,In_425);
or U1443 (N_1443,In_499,In_335);
or U1444 (N_1444,In_165,In_556);
or U1445 (N_1445,In_584,In_665);
or U1446 (N_1446,In_514,In_301);
nand U1447 (N_1447,In_336,In_769);
xor U1448 (N_1448,In_541,In_851);
nor U1449 (N_1449,In_623,In_889);
and U1450 (N_1450,In_816,In_959);
and U1451 (N_1451,In_365,In_611);
nand U1452 (N_1452,In_770,In_120);
or U1453 (N_1453,In_243,In_441);
and U1454 (N_1454,In_907,In_393);
or U1455 (N_1455,In_334,In_52);
xor U1456 (N_1456,In_105,In_240);
nand U1457 (N_1457,In_416,In_875);
nand U1458 (N_1458,In_362,In_22);
nor U1459 (N_1459,In_760,In_880);
nor U1460 (N_1460,In_396,In_234);
or U1461 (N_1461,In_426,In_354);
or U1462 (N_1462,In_410,In_29);
nor U1463 (N_1463,In_339,In_505);
xor U1464 (N_1464,In_880,In_941);
nor U1465 (N_1465,In_372,In_267);
nand U1466 (N_1466,In_394,In_850);
xnor U1467 (N_1467,In_942,In_369);
nand U1468 (N_1468,In_764,In_431);
and U1469 (N_1469,In_278,In_594);
xor U1470 (N_1470,In_313,In_953);
xnor U1471 (N_1471,In_600,In_554);
and U1472 (N_1472,In_419,In_649);
nand U1473 (N_1473,In_250,In_916);
or U1474 (N_1474,In_504,In_17);
and U1475 (N_1475,In_643,In_603);
or U1476 (N_1476,In_580,In_921);
nor U1477 (N_1477,In_33,In_416);
nand U1478 (N_1478,In_793,In_495);
nor U1479 (N_1479,In_551,In_290);
xor U1480 (N_1480,In_567,In_60);
or U1481 (N_1481,In_626,In_511);
xnor U1482 (N_1482,In_541,In_237);
or U1483 (N_1483,In_128,In_439);
xor U1484 (N_1484,In_495,In_772);
or U1485 (N_1485,In_35,In_340);
and U1486 (N_1486,In_546,In_68);
and U1487 (N_1487,In_955,In_469);
nor U1488 (N_1488,In_662,In_954);
nand U1489 (N_1489,In_988,In_420);
or U1490 (N_1490,In_667,In_498);
or U1491 (N_1491,In_501,In_805);
xor U1492 (N_1492,In_776,In_549);
or U1493 (N_1493,In_601,In_859);
xnor U1494 (N_1494,In_453,In_884);
xor U1495 (N_1495,In_249,In_629);
or U1496 (N_1496,In_33,In_478);
xor U1497 (N_1497,In_0,In_331);
xor U1498 (N_1498,In_554,In_779);
xnor U1499 (N_1499,In_578,In_315);
nor U1500 (N_1500,In_898,In_299);
xnor U1501 (N_1501,In_508,In_584);
nand U1502 (N_1502,In_266,In_12);
and U1503 (N_1503,In_857,In_383);
and U1504 (N_1504,In_762,In_400);
nand U1505 (N_1505,In_254,In_599);
nand U1506 (N_1506,In_842,In_729);
nand U1507 (N_1507,In_187,In_753);
nor U1508 (N_1508,In_298,In_879);
nand U1509 (N_1509,In_694,In_377);
and U1510 (N_1510,In_100,In_245);
xor U1511 (N_1511,In_319,In_754);
and U1512 (N_1512,In_134,In_744);
xnor U1513 (N_1513,In_524,In_411);
xnor U1514 (N_1514,In_759,In_83);
nand U1515 (N_1515,In_904,In_866);
or U1516 (N_1516,In_941,In_699);
nor U1517 (N_1517,In_758,In_224);
and U1518 (N_1518,In_175,In_143);
or U1519 (N_1519,In_38,In_752);
nor U1520 (N_1520,In_536,In_306);
or U1521 (N_1521,In_544,In_360);
or U1522 (N_1522,In_117,In_588);
and U1523 (N_1523,In_449,In_691);
nand U1524 (N_1524,In_109,In_273);
nor U1525 (N_1525,In_128,In_321);
xnor U1526 (N_1526,In_186,In_309);
xnor U1527 (N_1527,In_216,In_400);
and U1528 (N_1528,In_962,In_459);
xor U1529 (N_1529,In_808,In_10);
nor U1530 (N_1530,In_244,In_570);
nand U1531 (N_1531,In_885,In_722);
nand U1532 (N_1532,In_903,In_386);
or U1533 (N_1533,In_293,In_176);
xnor U1534 (N_1534,In_556,In_135);
nand U1535 (N_1535,In_272,In_456);
nand U1536 (N_1536,In_347,In_11);
xor U1537 (N_1537,In_537,In_942);
or U1538 (N_1538,In_878,In_831);
nand U1539 (N_1539,In_400,In_770);
or U1540 (N_1540,In_202,In_132);
or U1541 (N_1541,In_208,In_663);
and U1542 (N_1542,In_806,In_387);
nand U1543 (N_1543,In_646,In_442);
or U1544 (N_1544,In_409,In_286);
or U1545 (N_1545,In_229,In_576);
nand U1546 (N_1546,In_881,In_61);
nand U1547 (N_1547,In_186,In_166);
nand U1548 (N_1548,In_708,In_276);
xnor U1549 (N_1549,In_407,In_628);
xnor U1550 (N_1550,In_775,In_206);
nand U1551 (N_1551,In_14,In_433);
xnor U1552 (N_1552,In_58,In_307);
or U1553 (N_1553,In_741,In_640);
nor U1554 (N_1554,In_444,In_692);
nor U1555 (N_1555,In_584,In_235);
or U1556 (N_1556,In_737,In_484);
or U1557 (N_1557,In_161,In_568);
nor U1558 (N_1558,In_195,In_248);
and U1559 (N_1559,In_355,In_82);
nand U1560 (N_1560,In_144,In_455);
and U1561 (N_1561,In_890,In_872);
or U1562 (N_1562,In_258,In_863);
xor U1563 (N_1563,In_637,In_762);
and U1564 (N_1564,In_965,In_241);
xnor U1565 (N_1565,In_430,In_358);
nand U1566 (N_1566,In_78,In_681);
xnor U1567 (N_1567,In_72,In_669);
nor U1568 (N_1568,In_209,In_144);
xor U1569 (N_1569,In_175,In_859);
and U1570 (N_1570,In_879,In_70);
and U1571 (N_1571,In_311,In_192);
xnor U1572 (N_1572,In_317,In_673);
xor U1573 (N_1573,In_599,In_474);
or U1574 (N_1574,In_551,In_850);
nand U1575 (N_1575,In_533,In_122);
or U1576 (N_1576,In_462,In_47);
xor U1577 (N_1577,In_129,In_633);
xnor U1578 (N_1578,In_290,In_604);
and U1579 (N_1579,In_703,In_937);
nor U1580 (N_1580,In_575,In_661);
and U1581 (N_1581,In_384,In_951);
and U1582 (N_1582,In_961,In_976);
xor U1583 (N_1583,In_971,In_603);
xnor U1584 (N_1584,In_856,In_713);
nor U1585 (N_1585,In_957,In_648);
nor U1586 (N_1586,In_160,In_63);
and U1587 (N_1587,In_950,In_411);
nand U1588 (N_1588,In_583,In_195);
xnor U1589 (N_1589,In_734,In_318);
nor U1590 (N_1590,In_161,In_25);
or U1591 (N_1591,In_415,In_252);
and U1592 (N_1592,In_908,In_100);
nor U1593 (N_1593,In_766,In_914);
nand U1594 (N_1594,In_371,In_314);
xor U1595 (N_1595,In_641,In_307);
nor U1596 (N_1596,In_467,In_324);
nand U1597 (N_1597,In_87,In_919);
nor U1598 (N_1598,In_900,In_952);
nor U1599 (N_1599,In_63,In_213);
and U1600 (N_1600,In_255,In_105);
nor U1601 (N_1601,In_811,In_993);
and U1602 (N_1602,In_750,In_448);
or U1603 (N_1603,In_991,In_752);
xor U1604 (N_1604,In_542,In_280);
or U1605 (N_1605,In_493,In_211);
xor U1606 (N_1606,In_748,In_168);
nand U1607 (N_1607,In_157,In_508);
and U1608 (N_1608,In_706,In_478);
nor U1609 (N_1609,In_978,In_353);
nand U1610 (N_1610,In_841,In_43);
nor U1611 (N_1611,In_805,In_362);
nor U1612 (N_1612,In_506,In_165);
nand U1613 (N_1613,In_98,In_529);
and U1614 (N_1614,In_532,In_624);
or U1615 (N_1615,In_981,In_558);
and U1616 (N_1616,In_173,In_398);
or U1617 (N_1617,In_573,In_319);
xnor U1618 (N_1618,In_156,In_264);
nand U1619 (N_1619,In_150,In_583);
and U1620 (N_1620,In_202,In_244);
xor U1621 (N_1621,In_632,In_992);
or U1622 (N_1622,In_213,In_47);
nor U1623 (N_1623,In_714,In_487);
xor U1624 (N_1624,In_530,In_558);
or U1625 (N_1625,In_303,In_972);
xor U1626 (N_1626,In_571,In_768);
nor U1627 (N_1627,In_985,In_195);
or U1628 (N_1628,In_290,In_375);
nand U1629 (N_1629,In_87,In_106);
xor U1630 (N_1630,In_711,In_376);
nand U1631 (N_1631,In_964,In_819);
nor U1632 (N_1632,In_282,In_917);
and U1633 (N_1633,In_956,In_711);
and U1634 (N_1634,In_921,In_36);
nand U1635 (N_1635,In_145,In_169);
or U1636 (N_1636,In_385,In_395);
nand U1637 (N_1637,In_982,In_601);
nor U1638 (N_1638,In_227,In_676);
and U1639 (N_1639,In_629,In_939);
xnor U1640 (N_1640,In_439,In_930);
nor U1641 (N_1641,In_787,In_884);
or U1642 (N_1642,In_219,In_423);
or U1643 (N_1643,In_116,In_811);
nor U1644 (N_1644,In_233,In_787);
and U1645 (N_1645,In_895,In_570);
nand U1646 (N_1646,In_527,In_919);
and U1647 (N_1647,In_598,In_762);
nor U1648 (N_1648,In_557,In_610);
xor U1649 (N_1649,In_952,In_664);
nor U1650 (N_1650,In_180,In_851);
xnor U1651 (N_1651,In_589,In_926);
xor U1652 (N_1652,In_55,In_460);
and U1653 (N_1653,In_673,In_273);
nor U1654 (N_1654,In_943,In_775);
nor U1655 (N_1655,In_896,In_617);
or U1656 (N_1656,In_466,In_715);
nor U1657 (N_1657,In_250,In_831);
nand U1658 (N_1658,In_424,In_914);
nor U1659 (N_1659,In_980,In_295);
nand U1660 (N_1660,In_663,In_17);
nor U1661 (N_1661,In_481,In_955);
nand U1662 (N_1662,In_844,In_202);
or U1663 (N_1663,In_304,In_11);
nand U1664 (N_1664,In_198,In_52);
nand U1665 (N_1665,In_987,In_276);
nor U1666 (N_1666,In_290,In_107);
and U1667 (N_1667,In_639,In_527);
nor U1668 (N_1668,In_499,In_692);
xor U1669 (N_1669,In_171,In_55);
nor U1670 (N_1670,In_939,In_974);
xor U1671 (N_1671,In_750,In_638);
and U1672 (N_1672,In_563,In_422);
or U1673 (N_1673,In_675,In_171);
and U1674 (N_1674,In_551,In_345);
and U1675 (N_1675,In_305,In_69);
or U1676 (N_1676,In_374,In_822);
nor U1677 (N_1677,In_224,In_143);
nand U1678 (N_1678,In_922,In_870);
or U1679 (N_1679,In_590,In_773);
or U1680 (N_1680,In_129,In_645);
nor U1681 (N_1681,In_564,In_580);
xor U1682 (N_1682,In_941,In_661);
nor U1683 (N_1683,In_448,In_263);
and U1684 (N_1684,In_869,In_627);
nor U1685 (N_1685,In_981,In_273);
nor U1686 (N_1686,In_689,In_13);
xor U1687 (N_1687,In_683,In_385);
nand U1688 (N_1688,In_231,In_740);
or U1689 (N_1689,In_157,In_3);
or U1690 (N_1690,In_741,In_755);
nand U1691 (N_1691,In_821,In_597);
nor U1692 (N_1692,In_138,In_2);
nand U1693 (N_1693,In_911,In_971);
and U1694 (N_1694,In_813,In_962);
and U1695 (N_1695,In_894,In_892);
nor U1696 (N_1696,In_331,In_52);
nor U1697 (N_1697,In_713,In_469);
or U1698 (N_1698,In_249,In_630);
and U1699 (N_1699,In_221,In_63);
and U1700 (N_1700,In_634,In_762);
and U1701 (N_1701,In_172,In_951);
nand U1702 (N_1702,In_234,In_236);
and U1703 (N_1703,In_467,In_925);
xor U1704 (N_1704,In_78,In_374);
nand U1705 (N_1705,In_868,In_202);
or U1706 (N_1706,In_770,In_278);
or U1707 (N_1707,In_231,In_237);
xnor U1708 (N_1708,In_355,In_599);
or U1709 (N_1709,In_603,In_402);
and U1710 (N_1710,In_48,In_200);
nor U1711 (N_1711,In_70,In_801);
and U1712 (N_1712,In_657,In_250);
and U1713 (N_1713,In_566,In_528);
and U1714 (N_1714,In_904,In_375);
xnor U1715 (N_1715,In_570,In_683);
nor U1716 (N_1716,In_578,In_884);
nor U1717 (N_1717,In_432,In_403);
xnor U1718 (N_1718,In_311,In_992);
nor U1719 (N_1719,In_725,In_163);
or U1720 (N_1720,In_118,In_12);
and U1721 (N_1721,In_374,In_626);
or U1722 (N_1722,In_288,In_934);
xnor U1723 (N_1723,In_164,In_32);
and U1724 (N_1724,In_840,In_724);
and U1725 (N_1725,In_588,In_446);
xor U1726 (N_1726,In_208,In_164);
xnor U1727 (N_1727,In_163,In_284);
nor U1728 (N_1728,In_639,In_274);
and U1729 (N_1729,In_546,In_879);
xor U1730 (N_1730,In_872,In_152);
and U1731 (N_1731,In_527,In_611);
xnor U1732 (N_1732,In_453,In_866);
or U1733 (N_1733,In_929,In_23);
nand U1734 (N_1734,In_170,In_583);
or U1735 (N_1735,In_249,In_143);
nor U1736 (N_1736,In_92,In_421);
or U1737 (N_1737,In_0,In_727);
xnor U1738 (N_1738,In_837,In_480);
nor U1739 (N_1739,In_401,In_935);
or U1740 (N_1740,In_131,In_285);
nand U1741 (N_1741,In_865,In_196);
nand U1742 (N_1742,In_258,In_432);
nand U1743 (N_1743,In_10,In_384);
nor U1744 (N_1744,In_235,In_243);
and U1745 (N_1745,In_381,In_32);
nand U1746 (N_1746,In_409,In_266);
and U1747 (N_1747,In_782,In_340);
nand U1748 (N_1748,In_219,In_833);
nand U1749 (N_1749,In_845,In_893);
xnor U1750 (N_1750,In_343,In_643);
xor U1751 (N_1751,In_826,In_376);
nor U1752 (N_1752,In_174,In_67);
xnor U1753 (N_1753,In_277,In_402);
or U1754 (N_1754,In_679,In_392);
or U1755 (N_1755,In_967,In_344);
or U1756 (N_1756,In_926,In_520);
nor U1757 (N_1757,In_673,In_796);
or U1758 (N_1758,In_600,In_165);
nor U1759 (N_1759,In_555,In_120);
or U1760 (N_1760,In_690,In_447);
nor U1761 (N_1761,In_398,In_602);
or U1762 (N_1762,In_110,In_755);
and U1763 (N_1763,In_605,In_304);
xor U1764 (N_1764,In_849,In_434);
and U1765 (N_1765,In_270,In_65);
and U1766 (N_1766,In_143,In_166);
xnor U1767 (N_1767,In_776,In_279);
and U1768 (N_1768,In_767,In_342);
or U1769 (N_1769,In_156,In_710);
nand U1770 (N_1770,In_734,In_56);
and U1771 (N_1771,In_155,In_825);
nand U1772 (N_1772,In_478,In_895);
xnor U1773 (N_1773,In_375,In_589);
xor U1774 (N_1774,In_572,In_358);
xor U1775 (N_1775,In_557,In_183);
nand U1776 (N_1776,In_224,In_341);
nand U1777 (N_1777,In_551,In_497);
nand U1778 (N_1778,In_99,In_873);
nor U1779 (N_1779,In_375,In_567);
nor U1780 (N_1780,In_542,In_390);
nor U1781 (N_1781,In_581,In_233);
or U1782 (N_1782,In_107,In_67);
and U1783 (N_1783,In_405,In_675);
and U1784 (N_1784,In_983,In_598);
nor U1785 (N_1785,In_245,In_471);
nand U1786 (N_1786,In_663,In_553);
and U1787 (N_1787,In_922,In_133);
or U1788 (N_1788,In_904,In_433);
nor U1789 (N_1789,In_553,In_961);
and U1790 (N_1790,In_81,In_418);
nand U1791 (N_1791,In_548,In_254);
or U1792 (N_1792,In_552,In_923);
nor U1793 (N_1793,In_127,In_473);
nor U1794 (N_1794,In_1,In_662);
nand U1795 (N_1795,In_716,In_799);
nand U1796 (N_1796,In_509,In_497);
and U1797 (N_1797,In_106,In_287);
or U1798 (N_1798,In_633,In_120);
and U1799 (N_1799,In_138,In_65);
xor U1800 (N_1800,In_129,In_281);
nand U1801 (N_1801,In_864,In_180);
and U1802 (N_1802,In_902,In_96);
or U1803 (N_1803,In_285,In_674);
or U1804 (N_1804,In_489,In_842);
and U1805 (N_1805,In_277,In_664);
xnor U1806 (N_1806,In_867,In_82);
nor U1807 (N_1807,In_359,In_723);
nand U1808 (N_1808,In_385,In_944);
and U1809 (N_1809,In_220,In_537);
nand U1810 (N_1810,In_150,In_287);
nand U1811 (N_1811,In_188,In_154);
nor U1812 (N_1812,In_717,In_530);
nor U1813 (N_1813,In_37,In_928);
and U1814 (N_1814,In_624,In_578);
xor U1815 (N_1815,In_49,In_242);
nor U1816 (N_1816,In_430,In_535);
or U1817 (N_1817,In_71,In_415);
and U1818 (N_1818,In_664,In_45);
nand U1819 (N_1819,In_992,In_961);
nor U1820 (N_1820,In_282,In_360);
or U1821 (N_1821,In_453,In_24);
xor U1822 (N_1822,In_185,In_476);
nand U1823 (N_1823,In_655,In_722);
or U1824 (N_1824,In_275,In_806);
or U1825 (N_1825,In_63,In_316);
and U1826 (N_1826,In_468,In_530);
and U1827 (N_1827,In_660,In_841);
and U1828 (N_1828,In_24,In_500);
xor U1829 (N_1829,In_210,In_895);
xnor U1830 (N_1830,In_538,In_631);
or U1831 (N_1831,In_374,In_157);
xnor U1832 (N_1832,In_73,In_256);
or U1833 (N_1833,In_181,In_161);
or U1834 (N_1834,In_780,In_835);
nand U1835 (N_1835,In_698,In_664);
xor U1836 (N_1836,In_456,In_688);
or U1837 (N_1837,In_522,In_585);
xor U1838 (N_1838,In_173,In_704);
nor U1839 (N_1839,In_387,In_23);
xnor U1840 (N_1840,In_632,In_383);
nand U1841 (N_1841,In_79,In_538);
nand U1842 (N_1842,In_938,In_16);
xnor U1843 (N_1843,In_104,In_126);
and U1844 (N_1844,In_955,In_143);
xor U1845 (N_1845,In_624,In_906);
nor U1846 (N_1846,In_404,In_326);
and U1847 (N_1847,In_222,In_614);
xnor U1848 (N_1848,In_22,In_708);
or U1849 (N_1849,In_335,In_796);
nand U1850 (N_1850,In_239,In_468);
xor U1851 (N_1851,In_541,In_278);
nor U1852 (N_1852,In_955,In_769);
and U1853 (N_1853,In_889,In_594);
nor U1854 (N_1854,In_405,In_384);
xnor U1855 (N_1855,In_129,In_678);
nand U1856 (N_1856,In_172,In_797);
and U1857 (N_1857,In_940,In_93);
or U1858 (N_1858,In_175,In_161);
and U1859 (N_1859,In_647,In_121);
xor U1860 (N_1860,In_982,In_367);
xnor U1861 (N_1861,In_984,In_611);
nor U1862 (N_1862,In_302,In_430);
and U1863 (N_1863,In_420,In_583);
nor U1864 (N_1864,In_143,In_167);
xnor U1865 (N_1865,In_186,In_924);
and U1866 (N_1866,In_899,In_100);
or U1867 (N_1867,In_350,In_120);
nand U1868 (N_1868,In_704,In_959);
or U1869 (N_1869,In_893,In_179);
nor U1870 (N_1870,In_542,In_144);
nor U1871 (N_1871,In_702,In_528);
and U1872 (N_1872,In_709,In_206);
and U1873 (N_1873,In_488,In_252);
nor U1874 (N_1874,In_373,In_65);
or U1875 (N_1875,In_191,In_300);
nor U1876 (N_1876,In_802,In_553);
xnor U1877 (N_1877,In_9,In_176);
or U1878 (N_1878,In_289,In_155);
nor U1879 (N_1879,In_169,In_916);
nor U1880 (N_1880,In_61,In_504);
xor U1881 (N_1881,In_745,In_584);
nor U1882 (N_1882,In_710,In_975);
nand U1883 (N_1883,In_448,In_797);
nor U1884 (N_1884,In_254,In_575);
nand U1885 (N_1885,In_819,In_969);
nand U1886 (N_1886,In_914,In_859);
and U1887 (N_1887,In_426,In_709);
or U1888 (N_1888,In_193,In_590);
nand U1889 (N_1889,In_959,In_514);
and U1890 (N_1890,In_212,In_149);
and U1891 (N_1891,In_259,In_496);
nand U1892 (N_1892,In_368,In_98);
nor U1893 (N_1893,In_149,In_671);
nand U1894 (N_1894,In_273,In_545);
and U1895 (N_1895,In_456,In_757);
and U1896 (N_1896,In_533,In_308);
xor U1897 (N_1897,In_184,In_390);
nor U1898 (N_1898,In_662,In_166);
xnor U1899 (N_1899,In_49,In_699);
or U1900 (N_1900,In_149,In_268);
and U1901 (N_1901,In_495,In_242);
nand U1902 (N_1902,In_685,In_273);
or U1903 (N_1903,In_437,In_511);
or U1904 (N_1904,In_463,In_766);
xnor U1905 (N_1905,In_177,In_716);
nand U1906 (N_1906,In_67,In_282);
nor U1907 (N_1907,In_867,In_617);
nand U1908 (N_1908,In_18,In_476);
nor U1909 (N_1909,In_14,In_859);
nor U1910 (N_1910,In_507,In_192);
nand U1911 (N_1911,In_458,In_173);
nand U1912 (N_1912,In_942,In_155);
nand U1913 (N_1913,In_815,In_169);
and U1914 (N_1914,In_384,In_124);
and U1915 (N_1915,In_857,In_191);
nor U1916 (N_1916,In_340,In_758);
or U1917 (N_1917,In_565,In_378);
nand U1918 (N_1918,In_471,In_434);
and U1919 (N_1919,In_49,In_42);
nand U1920 (N_1920,In_903,In_308);
xnor U1921 (N_1921,In_980,In_716);
or U1922 (N_1922,In_344,In_141);
nand U1923 (N_1923,In_265,In_287);
and U1924 (N_1924,In_8,In_994);
xor U1925 (N_1925,In_361,In_140);
xnor U1926 (N_1926,In_341,In_782);
nand U1927 (N_1927,In_424,In_186);
xor U1928 (N_1928,In_279,In_861);
or U1929 (N_1929,In_168,In_362);
xnor U1930 (N_1930,In_77,In_647);
or U1931 (N_1931,In_410,In_324);
nand U1932 (N_1932,In_396,In_277);
or U1933 (N_1933,In_530,In_342);
nand U1934 (N_1934,In_824,In_814);
nand U1935 (N_1935,In_442,In_985);
or U1936 (N_1936,In_625,In_392);
nor U1937 (N_1937,In_569,In_67);
nand U1938 (N_1938,In_909,In_939);
nand U1939 (N_1939,In_63,In_951);
nand U1940 (N_1940,In_339,In_60);
nor U1941 (N_1941,In_102,In_331);
xor U1942 (N_1942,In_470,In_171);
or U1943 (N_1943,In_86,In_444);
xor U1944 (N_1944,In_508,In_756);
and U1945 (N_1945,In_805,In_290);
nor U1946 (N_1946,In_101,In_329);
nand U1947 (N_1947,In_855,In_276);
nand U1948 (N_1948,In_391,In_45);
nor U1949 (N_1949,In_83,In_64);
xnor U1950 (N_1950,In_816,In_407);
and U1951 (N_1951,In_862,In_529);
xor U1952 (N_1952,In_866,In_560);
xnor U1953 (N_1953,In_690,In_503);
nor U1954 (N_1954,In_10,In_763);
nor U1955 (N_1955,In_419,In_877);
or U1956 (N_1956,In_455,In_423);
nor U1957 (N_1957,In_260,In_416);
nand U1958 (N_1958,In_432,In_469);
nor U1959 (N_1959,In_372,In_965);
and U1960 (N_1960,In_251,In_856);
or U1961 (N_1961,In_56,In_516);
nor U1962 (N_1962,In_73,In_587);
or U1963 (N_1963,In_511,In_952);
or U1964 (N_1964,In_88,In_256);
nand U1965 (N_1965,In_498,In_765);
and U1966 (N_1966,In_915,In_752);
nand U1967 (N_1967,In_271,In_316);
xnor U1968 (N_1968,In_653,In_196);
xnor U1969 (N_1969,In_988,In_894);
nand U1970 (N_1970,In_875,In_842);
nor U1971 (N_1971,In_115,In_524);
xor U1972 (N_1972,In_467,In_792);
nand U1973 (N_1973,In_74,In_395);
or U1974 (N_1974,In_804,In_256);
xnor U1975 (N_1975,In_785,In_834);
nor U1976 (N_1976,In_343,In_868);
or U1977 (N_1977,In_148,In_813);
or U1978 (N_1978,In_468,In_956);
or U1979 (N_1979,In_370,In_316);
nand U1980 (N_1980,In_239,In_263);
nor U1981 (N_1981,In_213,In_722);
xor U1982 (N_1982,In_695,In_324);
nand U1983 (N_1983,In_388,In_39);
and U1984 (N_1984,In_134,In_971);
nand U1985 (N_1985,In_671,In_524);
xnor U1986 (N_1986,In_839,In_604);
or U1987 (N_1987,In_725,In_206);
xor U1988 (N_1988,In_868,In_330);
nor U1989 (N_1989,In_85,In_683);
nand U1990 (N_1990,In_267,In_209);
nor U1991 (N_1991,In_340,In_135);
nor U1992 (N_1992,In_343,In_369);
or U1993 (N_1993,In_931,In_108);
xnor U1994 (N_1994,In_690,In_301);
or U1995 (N_1995,In_286,In_628);
or U1996 (N_1996,In_553,In_297);
or U1997 (N_1997,In_12,In_4);
and U1998 (N_1998,In_235,In_875);
and U1999 (N_1999,In_257,In_85);
nand U2000 (N_2000,In_976,In_129);
xor U2001 (N_2001,In_623,In_492);
nor U2002 (N_2002,In_299,In_820);
nor U2003 (N_2003,In_122,In_621);
nand U2004 (N_2004,In_221,In_852);
xnor U2005 (N_2005,In_377,In_572);
nand U2006 (N_2006,In_64,In_344);
nand U2007 (N_2007,In_450,In_192);
or U2008 (N_2008,In_266,In_46);
xnor U2009 (N_2009,In_856,In_583);
and U2010 (N_2010,In_401,In_234);
nor U2011 (N_2011,In_168,In_881);
xnor U2012 (N_2012,In_477,In_320);
nor U2013 (N_2013,In_746,In_502);
xor U2014 (N_2014,In_387,In_918);
nand U2015 (N_2015,In_399,In_226);
and U2016 (N_2016,In_573,In_261);
nor U2017 (N_2017,In_103,In_100);
xor U2018 (N_2018,In_915,In_603);
and U2019 (N_2019,In_699,In_494);
nor U2020 (N_2020,In_982,In_834);
xor U2021 (N_2021,In_507,In_763);
and U2022 (N_2022,In_291,In_309);
nand U2023 (N_2023,In_593,In_786);
nand U2024 (N_2024,In_575,In_799);
or U2025 (N_2025,In_84,In_765);
or U2026 (N_2026,In_74,In_119);
nor U2027 (N_2027,In_211,In_954);
nand U2028 (N_2028,In_888,In_173);
nand U2029 (N_2029,In_402,In_360);
xor U2030 (N_2030,In_251,In_152);
nand U2031 (N_2031,In_636,In_889);
nand U2032 (N_2032,In_241,In_951);
and U2033 (N_2033,In_161,In_343);
or U2034 (N_2034,In_76,In_753);
and U2035 (N_2035,In_189,In_929);
or U2036 (N_2036,In_81,In_123);
and U2037 (N_2037,In_571,In_259);
and U2038 (N_2038,In_269,In_74);
nor U2039 (N_2039,In_608,In_319);
nand U2040 (N_2040,In_361,In_803);
and U2041 (N_2041,In_168,In_490);
nor U2042 (N_2042,In_234,In_237);
xor U2043 (N_2043,In_977,In_197);
xnor U2044 (N_2044,In_42,In_65);
and U2045 (N_2045,In_151,In_835);
xor U2046 (N_2046,In_705,In_472);
nand U2047 (N_2047,In_701,In_423);
xor U2048 (N_2048,In_556,In_827);
and U2049 (N_2049,In_208,In_358);
or U2050 (N_2050,In_932,In_661);
nand U2051 (N_2051,In_960,In_669);
nor U2052 (N_2052,In_956,In_746);
xnor U2053 (N_2053,In_478,In_540);
and U2054 (N_2054,In_829,In_254);
nand U2055 (N_2055,In_183,In_702);
nand U2056 (N_2056,In_982,In_479);
xor U2057 (N_2057,In_573,In_58);
or U2058 (N_2058,In_744,In_894);
or U2059 (N_2059,In_466,In_742);
or U2060 (N_2060,In_975,In_861);
nor U2061 (N_2061,In_275,In_594);
nor U2062 (N_2062,In_997,In_518);
nor U2063 (N_2063,In_673,In_428);
and U2064 (N_2064,In_95,In_433);
or U2065 (N_2065,In_214,In_534);
nand U2066 (N_2066,In_392,In_383);
nor U2067 (N_2067,In_385,In_561);
and U2068 (N_2068,In_420,In_452);
nor U2069 (N_2069,In_418,In_215);
nor U2070 (N_2070,In_901,In_238);
or U2071 (N_2071,In_189,In_938);
and U2072 (N_2072,In_275,In_499);
nor U2073 (N_2073,In_16,In_950);
nand U2074 (N_2074,In_7,In_395);
xnor U2075 (N_2075,In_870,In_67);
nand U2076 (N_2076,In_987,In_627);
nor U2077 (N_2077,In_818,In_594);
and U2078 (N_2078,In_669,In_238);
nand U2079 (N_2079,In_717,In_98);
xor U2080 (N_2080,In_160,In_317);
and U2081 (N_2081,In_333,In_193);
nor U2082 (N_2082,In_287,In_882);
nand U2083 (N_2083,In_916,In_838);
nand U2084 (N_2084,In_118,In_825);
xor U2085 (N_2085,In_545,In_677);
xnor U2086 (N_2086,In_573,In_153);
or U2087 (N_2087,In_201,In_137);
xnor U2088 (N_2088,In_75,In_320);
or U2089 (N_2089,In_494,In_602);
xor U2090 (N_2090,In_284,In_426);
or U2091 (N_2091,In_779,In_905);
or U2092 (N_2092,In_245,In_945);
nand U2093 (N_2093,In_718,In_94);
xnor U2094 (N_2094,In_498,In_622);
nor U2095 (N_2095,In_126,In_41);
xnor U2096 (N_2096,In_19,In_238);
or U2097 (N_2097,In_655,In_162);
nand U2098 (N_2098,In_560,In_58);
xnor U2099 (N_2099,In_401,In_597);
xor U2100 (N_2100,In_507,In_813);
xnor U2101 (N_2101,In_820,In_108);
nor U2102 (N_2102,In_800,In_862);
and U2103 (N_2103,In_777,In_580);
nand U2104 (N_2104,In_903,In_34);
or U2105 (N_2105,In_194,In_521);
and U2106 (N_2106,In_957,In_263);
xnor U2107 (N_2107,In_966,In_424);
nor U2108 (N_2108,In_964,In_376);
nor U2109 (N_2109,In_330,In_931);
xnor U2110 (N_2110,In_550,In_958);
xor U2111 (N_2111,In_892,In_674);
nor U2112 (N_2112,In_927,In_707);
xor U2113 (N_2113,In_91,In_812);
and U2114 (N_2114,In_54,In_525);
xnor U2115 (N_2115,In_454,In_330);
nand U2116 (N_2116,In_388,In_701);
xnor U2117 (N_2117,In_228,In_47);
and U2118 (N_2118,In_360,In_387);
or U2119 (N_2119,In_196,In_430);
or U2120 (N_2120,In_742,In_498);
and U2121 (N_2121,In_333,In_229);
and U2122 (N_2122,In_733,In_843);
xor U2123 (N_2123,In_427,In_949);
nand U2124 (N_2124,In_469,In_205);
or U2125 (N_2125,In_451,In_160);
xor U2126 (N_2126,In_425,In_515);
nor U2127 (N_2127,In_795,In_443);
nand U2128 (N_2128,In_602,In_725);
and U2129 (N_2129,In_457,In_62);
nor U2130 (N_2130,In_22,In_4);
xor U2131 (N_2131,In_474,In_861);
and U2132 (N_2132,In_80,In_204);
and U2133 (N_2133,In_594,In_74);
xnor U2134 (N_2134,In_228,In_869);
or U2135 (N_2135,In_196,In_243);
and U2136 (N_2136,In_384,In_694);
xor U2137 (N_2137,In_230,In_456);
and U2138 (N_2138,In_66,In_977);
and U2139 (N_2139,In_747,In_908);
nand U2140 (N_2140,In_898,In_113);
nor U2141 (N_2141,In_252,In_348);
nor U2142 (N_2142,In_28,In_559);
or U2143 (N_2143,In_226,In_854);
and U2144 (N_2144,In_736,In_844);
nor U2145 (N_2145,In_191,In_868);
and U2146 (N_2146,In_130,In_53);
nand U2147 (N_2147,In_436,In_201);
or U2148 (N_2148,In_546,In_392);
or U2149 (N_2149,In_918,In_76);
and U2150 (N_2150,In_306,In_272);
xor U2151 (N_2151,In_408,In_202);
or U2152 (N_2152,In_64,In_383);
nand U2153 (N_2153,In_389,In_295);
nand U2154 (N_2154,In_960,In_677);
and U2155 (N_2155,In_918,In_952);
nand U2156 (N_2156,In_780,In_163);
xnor U2157 (N_2157,In_128,In_978);
xnor U2158 (N_2158,In_633,In_51);
xnor U2159 (N_2159,In_348,In_518);
and U2160 (N_2160,In_616,In_739);
nand U2161 (N_2161,In_834,In_739);
nor U2162 (N_2162,In_157,In_839);
xnor U2163 (N_2163,In_806,In_585);
or U2164 (N_2164,In_940,In_330);
nor U2165 (N_2165,In_995,In_406);
nor U2166 (N_2166,In_982,In_207);
nand U2167 (N_2167,In_66,In_407);
and U2168 (N_2168,In_789,In_268);
or U2169 (N_2169,In_995,In_683);
nand U2170 (N_2170,In_16,In_886);
nor U2171 (N_2171,In_635,In_357);
xor U2172 (N_2172,In_895,In_247);
xor U2173 (N_2173,In_486,In_819);
nor U2174 (N_2174,In_366,In_49);
or U2175 (N_2175,In_713,In_793);
nor U2176 (N_2176,In_480,In_821);
xnor U2177 (N_2177,In_212,In_818);
xor U2178 (N_2178,In_777,In_665);
nor U2179 (N_2179,In_260,In_542);
nand U2180 (N_2180,In_191,In_534);
or U2181 (N_2181,In_209,In_342);
and U2182 (N_2182,In_585,In_147);
or U2183 (N_2183,In_237,In_716);
nor U2184 (N_2184,In_486,In_313);
xor U2185 (N_2185,In_948,In_973);
and U2186 (N_2186,In_67,In_533);
nand U2187 (N_2187,In_252,In_386);
nor U2188 (N_2188,In_826,In_215);
nor U2189 (N_2189,In_508,In_674);
and U2190 (N_2190,In_20,In_855);
nor U2191 (N_2191,In_53,In_125);
nand U2192 (N_2192,In_421,In_127);
nor U2193 (N_2193,In_845,In_450);
xor U2194 (N_2194,In_696,In_971);
or U2195 (N_2195,In_735,In_96);
nor U2196 (N_2196,In_901,In_719);
nand U2197 (N_2197,In_238,In_273);
nand U2198 (N_2198,In_250,In_346);
and U2199 (N_2199,In_328,In_63);
and U2200 (N_2200,In_570,In_218);
nand U2201 (N_2201,In_334,In_677);
xor U2202 (N_2202,In_518,In_38);
or U2203 (N_2203,In_750,In_77);
xor U2204 (N_2204,In_323,In_943);
nor U2205 (N_2205,In_560,In_245);
and U2206 (N_2206,In_531,In_136);
or U2207 (N_2207,In_232,In_31);
nor U2208 (N_2208,In_665,In_332);
xnor U2209 (N_2209,In_766,In_971);
and U2210 (N_2210,In_479,In_12);
and U2211 (N_2211,In_30,In_782);
nor U2212 (N_2212,In_125,In_605);
nor U2213 (N_2213,In_823,In_228);
or U2214 (N_2214,In_355,In_264);
or U2215 (N_2215,In_219,In_999);
nand U2216 (N_2216,In_410,In_317);
xor U2217 (N_2217,In_837,In_741);
or U2218 (N_2218,In_620,In_375);
nor U2219 (N_2219,In_219,In_799);
nand U2220 (N_2220,In_818,In_14);
or U2221 (N_2221,In_670,In_826);
or U2222 (N_2222,In_788,In_547);
xnor U2223 (N_2223,In_444,In_749);
or U2224 (N_2224,In_579,In_49);
nor U2225 (N_2225,In_823,In_695);
nor U2226 (N_2226,In_791,In_822);
nand U2227 (N_2227,In_557,In_692);
xnor U2228 (N_2228,In_295,In_622);
and U2229 (N_2229,In_170,In_498);
and U2230 (N_2230,In_674,In_245);
nor U2231 (N_2231,In_102,In_127);
nor U2232 (N_2232,In_296,In_745);
nor U2233 (N_2233,In_589,In_936);
nor U2234 (N_2234,In_155,In_32);
and U2235 (N_2235,In_607,In_626);
or U2236 (N_2236,In_594,In_401);
nor U2237 (N_2237,In_761,In_974);
nor U2238 (N_2238,In_81,In_627);
nand U2239 (N_2239,In_637,In_474);
nor U2240 (N_2240,In_747,In_4);
or U2241 (N_2241,In_70,In_669);
xnor U2242 (N_2242,In_231,In_65);
nor U2243 (N_2243,In_901,In_30);
and U2244 (N_2244,In_96,In_342);
nor U2245 (N_2245,In_826,In_350);
xnor U2246 (N_2246,In_577,In_429);
nor U2247 (N_2247,In_258,In_435);
and U2248 (N_2248,In_785,In_68);
nand U2249 (N_2249,In_428,In_68);
nor U2250 (N_2250,In_171,In_555);
nor U2251 (N_2251,In_666,In_891);
or U2252 (N_2252,In_366,In_976);
nand U2253 (N_2253,In_47,In_439);
and U2254 (N_2254,In_239,In_131);
nor U2255 (N_2255,In_610,In_425);
xor U2256 (N_2256,In_447,In_770);
xor U2257 (N_2257,In_820,In_878);
nand U2258 (N_2258,In_402,In_367);
or U2259 (N_2259,In_663,In_815);
nand U2260 (N_2260,In_869,In_247);
or U2261 (N_2261,In_614,In_560);
nor U2262 (N_2262,In_795,In_588);
nand U2263 (N_2263,In_316,In_646);
or U2264 (N_2264,In_350,In_158);
nand U2265 (N_2265,In_683,In_396);
and U2266 (N_2266,In_943,In_756);
nor U2267 (N_2267,In_239,In_366);
nor U2268 (N_2268,In_82,In_182);
or U2269 (N_2269,In_12,In_259);
xnor U2270 (N_2270,In_278,In_539);
or U2271 (N_2271,In_284,In_105);
or U2272 (N_2272,In_274,In_412);
nand U2273 (N_2273,In_517,In_281);
and U2274 (N_2274,In_450,In_377);
or U2275 (N_2275,In_561,In_727);
or U2276 (N_2276,In_679,In_318);
nor U2277 (N_2277,In_783,In_531);
xnor U2278 (N_2278,In_20,In_353);
and U2279 (N_2279,In_158,In_375);
and U2280 (N_2280,In_768,In_800);
and U2281 (N_2281,In_313,In_183);
nor U2282 (N_2282,In_51,In_225);
or U2283 (N_2283,In_949,In_324);
xnor U2284 (N_2284,In_447,In_686);
and U2285 (N_2285,In_52,In_769);
nand U2286 (N_2286,In_280,In_110);
nor U2287 (N_2287,In_984,In_325);
nor U2288 (N_2288,In_857,In_52);
xnor U2289 (N_2289,In_664,In_829);
nor U2290 (N_2290,In_542,In_152);
xnor U2291 (N_2291,In_93,In_835);
nand U2292 (N_2292,In_364,In_172);
and U2293 (N_2293,In_322,In_194);
nand U2294 (N_2294,In_19,In_394);
xnor U2295 (N_2295,In_712,In_844);
and U2296 (N_2296,In_854,In_18);
nor U2297 (N_2297,In_46,In_756);
and U2298 (N_2298,In_886,In_769);
nand U2299 (N_2299,In_874,In_366);
nor U2300 (N_2300,In_532,In_454);
and U2301 (N_2301,In_548,In_128);
and U2302 (N_2302,In_483,In_836);
and U2303 (N_2303,In_295,In_770);
or U2304 (N_2304,In_908,In_39);
and U2305 (N_2305,In_45,In_58);
nand U2306 (N_2306,In_955,In_215);
and U2307 (N_2307,In_274,In_352);
and U2308 (N_2308,In_543,In_88);
and U2309 (N_2309,In_799,In_871);
xnor U2310 (N_2310,In_200,In_954);
xor U2311 (N_2311,In_964,In_591);
xor U2312 (N_2312,In_226,In_595);
and U2313 (N_2313,In_64,In_233);
xnor U2314 (N_2314,In_114,In_426);
nor U2315 (N_2315,In_893,In_369);
or U2316 (N_2316,In_62,In_678);
or U2317 (N_2317,In_380,In_119);
nand U2318 (N_2318,In_484,In_361);
nand U2319 (N_2319,In_255,In_523);
and U2320 (N_2320,In_939,In_762);
nor U2321 (N_2321,In_791,In_994);
xor U2322 (N_2322,In_599,In_175);
nand U2323 (N_2323,In_535,In_75);
xnor U2324 (N_2324,In_20,In_977);
xnor U2325 (N_2325,In_307,In_819);
nand U2326 (N_2326,In_724,In_492);
and U2327 (N_2327,In_960,In_588);
xor U2328 (N_2328,In_972,In_466);
and U2329 (N_2329,In_916,In_367);
xnor U2330 (N_2330,In_745,In_719);
nor U2331 (N_2331,In_712,In_690);
nand U2332 (N_2332,In_926,In_586);
and U2333 (N_2333,In_90,In_895);
xor U2334 (N_2334,In_798,In_898);
nand U2335 (N_2335,In_975,In_383);
nor U2336 (N_2336,In_869,In_227);
nand U2337 (N_2337,In_129,In_619);
nor U2338 (N_2338,In_456,In_460);
or U2339 (N_2339,In_97,In_190);
or U2340 (N_2340,In_930,In_73);
nand U2341 (N_2341,In_967,In_432);
and U2342 (N_2342,In_977,In_304);
or U2343 (N_2343,In_843,In_694);
xor U2344 (N_2344,In_387,In_352);
nor U2345 (N_2345,In_971,In_524);
xor U2346 (N_2346,In_692,In_556);
and U2347 (N_2347,In_338,In_875);
xor U2348 (N_2348,In_987,In_529);
or U2349 (N_2349,In_711,In_358);
nor U2350 (N_2350,In_328,In_62);
nor U2351 (N_2351,In_608,In_714);
nor U2352 (N_2352,In_891,In_972);
and U2353 (N_2353,In_567,In_420);
or U2354 (N_2354,In_412,In_101);
and U2355 (N_2355,In_820,In_481);
xor U2356 (N_2356,In_119,In_837);
or U2357 (N_2357,In_279,In_73);
nor U2358 (N_2358,In_539,In_195);
xnor U2359 (N_2359,In_803,In_269);
nor U2360 (N_2360,In_869,In_569);
and U2361 (N_2361,In_864,In_785);
nor U2362 (N_2362,In_93,In_46);
nor U2363 (N_2363,In_484,In_196);
or U2364 (N_2364,In_124,In_185);
xor U2365 (N_2365,In_530,In_718);
nand U2366 (N_2366,In_750,In_999);
nand U2367 (N_2367,In_60,In_789);
nand U2368 (N_2368,In_302,In_116);
and U2369 (N_2369,In_71,In_523);
nand U2370 (N_2370,In_192,In_864);
and U2371 (N_2371,In_732,In_722);
xor U2372 (N_2372,In_129,In_382);
and U2373 (N_2373,In_425,In_359);
xor U2374 (N_2374,In_261,In_646);
nor U2375 (N_2375,In_122,In_370);
or U2376 (N_2376,In_520,In_687);
xnor U2377 (N_2377,In_795,In_963);
xnor U2378 (N_2378,In_30,In_777);
and U2379 (N_2379,In_204,In_541);
xnor U2380 (N_2380,In_582,In_750);
nand U2381 (N_2381,In_784,In_877);
nand U2382 (N_2382,In_590,In_604);
nor U2383 (N_2383,In_678,In_955);
nand U2384 (N_2384,In_169,In_49);
nor U2385 (N_2385,In_893,In_488);
or U2386 (N_2386,In_518,In_740);
nor U2387 (N_2387,In_832,In_220);
nor U2388 (N_2388,In_243,In_507);
or U2389 (N_2389,In_972,In_154);
nor U2390 (N_2390,In_719,In_678);
xor U2391 (N_2391,In_757,In_373);
nand U2392 (N_2392,In_236,In_469);
nand U2393 (N_2393,In_497,In_912);
nand U2394 (N_2394,In_947,In_209);
and U2395 (N_2395,In_129,In_917);
or U2396 (N_2396,In_808,In_829);
xor U2397 (N_2397,In_572,In_182);
nand U2398 (N_2398,In_231,In_802);
nand U2399 (N_2399,In_947,In_13);
nand U2400 (N_2400,In_25,In_396);
and U2401 (N_2401,In_565,In_160);
and U2402 (N_2402,In_106,In_518);
and U2403 (N_2403,In_664,In_520);
and U2404 (N_2404,In_73,In_873);
or U2405 (N_2405,In_299,In_551);
xor U2406 (N_2406,In_278,In_137);
xor U2407 (N_2407,In_436,In_755);
xnor U2408 (N_2408,In_959,In_374);
and U2409 (N_2409,In_963,In_757);
or U2410 (N_2410,In_564,In_603);
nor U2411 (N_2411,In_968,In_797);
nand U2412 (N_2412,In_322,In_901);
and U2413 (N_2413,In_910,In_871);
and U2414 (N_2414,In_547,In_386);
and U2415 (N_2415,In_15,In_444);
nand U2416 (N_2416,In_990,In_324);
nor U2417 (N_2417,In_135,In_704);
nor U2418 (N_2418,In_535,In_397);
or U2419 (N_2419,In_121,In_651);
or U2420 (N_2420,In_670,In_69);
nor U2421 (N_2421,In_650,In_822);
xnor U2422 (N_2422,In_903,In_237);
nand U2423 (N_2423,In_870,In_881);
and U2424 (N_2424,In_28,In_706);
nand U2425 (N_2425,In_184,In_560);
nor U2426 (N_2426,In_421,In_758);
nand U2427 (N_2427,In_702,In_942);
xor U2428 (N_2428,In_140,In_675);
and U2429 (N_2429,In_202,In_923);
xnor U2430 (N_2430,In_49,In_764);
and U2431 (N_2431,In_518,In_676);
or U2432 (N_2432,In_219,In_11);
xnor U2433 (N_2433,In_598,In_795);
nor U2434 (N_2434,In_453,In_784);
and U2435 (N_2435,In_983,In_119);
nor U2436 (N_2436,In_133,In_761);
nor U2437 (N_2437,In_690,In_146);
and U2438 (N_2438,In_45,In_801);
and U2439 (N_2439,In_319,In_643);
xor U2440 (N_2440,In_367,In_892);
and U2441 (N_2441,In_744,In_498);
nor U2442 (N_2442,In_48,In_33);
or U2443 (N_2443,In_58,In_628);
xnor U2444 (N_2444,In_115,In_277);
xor U2445 (N_2445,In_190,In_157);
nor U2446 (N_2446,In_152,In_318);
nand U2447 (N_2447,In_990,In_557);
or U2448 (N_2448,In_875,In_180);
nor U2449 (N_2449,In_925,In_76);
or U2450 (N_2450,In_560,In_869);
and U2451 (N_2451,In_315,In_179);
xnor U2452 (N_2452,In_660,In_218);
or U2453 (N_2453,In_622,In_160);
or U2454 (N_2454,In_338,In_497);
or U2455 (N_2455,In_366,In_72);
and U2456 (N_2456,In_649,In_553);
xor U2457 (N_2457,In_67,In_43);
nand U2458 (N_2458,In_768,In_471);
and U2459 (N_2459,In_590,In_482);
or U2460 (N_2460,In_52,In_799);
xnor U2461 (N_2461,In_83,In_384);
nand U2462 (N_2462,In_14,In_275);
xnor U2463 (N_2463,In_36,In_64);
nand U2464 (N_2464,In_464,In_778);
nor U2465 (N_2465,In_846,In_933);
or U2466 (N_2466,In_414,In_593);
or U2467 (N_2467,In_510,In_677);
or U2468 (N_2468,In_949,In_710);
nor U2469 (N_2469,In_439,In_223);
or U2470 (N_2470,In_696,In_991);
or U2471 (N_2471,In_625,In_75);
or U2472 (N_2472,In_230,In_572);
or U2473 (N_2473,In_835,In_82);
or U2474 (N_2474,In_178,In_747);
nand U2475 (N_2475,In_193,In_58);
nand U2476 (N_2476,In_484,In_442);
nand U2477 (N_2477,In_384,In_292);
xor U2478 (N_2478,In_923,In_218);
nand U2479 (N_2479,In_199,In_470);
nand U2480 (N_2480,In_879,In_553);
nand U2481 (N_2481,In_884,In_925);
nor U2482 (N_2482,In_660,In_193);
or U2483 (N_2483,In_968,In_287);
and U2484 (N_2484,In_77,In_430);
nor U2485 (N_2485,In_669,In_662);
and U2486 (N_2486,In_414,In_452);
or U2487 (N_2487,In_374,In_981);
nand U2488 (N_2488,In_783,In_507);
xnor U2489 (N_2489,In_821,In_138);
and U2490 (N_2490,In_198,In_559);
and U2491 (N_2491,In_797,In_807);
and U2492 (N_2492,In_976,In_632);
nand U2493 (N_2493,In_110,In_691);
nand U2494 (N_2494,In_318,In_272);
and U2495 (N_2495,In_836,In_42);
and U2496 (N_2496,In_437,In_176);
nand U2497 (N_2497,In_589,In_461);
or U2498 (N_2498,In_845,In_944);
nor U2499 (N_2499,In_421,In_272);
or U2500 (N_2500,In_605,In_845);
or U2501 (N_2501,In_472,In_449);
xnor U2502 (N_2502,In_969,In_361);
and U2503 (N_2503,In_982,In_958);
nand U2504 (N_2504,In_167,In_47);
and U2505 (N_2505,In_652,In_747);
xor U2506 (N_2506,In_139,In_862);
nor U2507 (N_2507,In_80,In_25);
nand U2508 (N_2508,In_87,In_928);
nor U2509 (N_2509,In_651,In_103);
xnor U2510 (N_2510,In_583,In_775);
nand U2511 (N_2511,In_776,In_127);
nor U2512 (N_2512,In_600,In_232);
xnor U2513 (N_2513,In_567,In_572);
nand U2514 (N_2514,In_335,In_808);
nor U2515 (N_2515,In_941,In_795);
nor U2516 (N_2516,In_701,In_878);
or U2517 (N_2517,In_850,In_219);
nor U2518 (N_2518,In_659,In_88);
nor U2519 (N_2519,In_815,In_616);
or U2520 (N_2520,In_192,In_349);
nand U2521 (N_2521,In_409,In_546);
or U2522 (N_2522,In_355,In_797);
nand U2523 (N_2523,In_202,In_257);
or U2524 (N_2524,In_171,In_123);
nand U2525 (N_2525,In_91,In_532);
or U2526 (N_2526,In_273,In_343);
nor U2527 (N_2527,In_370,In_340);
xnor U2528 (N_2528,In_837,In_469);
and U2529 (N_2529,In_122,In_440);
nor U2530 (N_2530,In_5,In_241);
and U2531 (N_2531,In_767,In_322);
xor U2532 (N_2532,In_758,In_211);
or U2533 (N_2533,In_476,In_620);
or U2534 (N_2534,In_45,In_459);
and U2535 (N_2535,In_816,In_508);
nor U2536 (N_2536,In_892,In_895);
xnor U2537 (N_2537,In_123,In_899);
xnor U2538 (N_2538,In_395,In_611);
xnor U2539 (N_2539,In_170,In_858);
nor U2540 (N_2540,In_584,In_245);
xnor U2541 (N_2541,In_348,In_289);
xnor U2542 (N_2542,In_108,In_514);
and U2543 (N_2543,In_173,In_332);
xor U2544 (N_2544,In_64,In_204);
nand U2545 (N_2545,In_71,In_520);
and U2546 (N_2546,In_559,In_511);
nor U2547 (N_2547,In_141,In_245);
or U2548 (N_2548,In_152,In_598);
xnor U2549 (N_2549,In_330,In_930);
xnor U2550 (N_2550,In_955,In_571);
nor U2551 (N_2551,In_17,In_919);
nand U2552 (N_2552,In_504,In_58);
nor U2553 (N_2553,In_583,In_24);
nor U2554 (N_2554,In_215,In_692);
or U2555 (N_2555,In_100,In_550);
and U2556 (N_2556,In_770,In_741);
nor U2557 (N_2557,In_419,In_404);
nor U2558 (N_2558,In_846,In_268);
xor U2559 (N_2559,In_867,In_726);
nand U2560 (N_2560,In_293,In_633);
xnor U2561 (N_2561,In_961,In_148);
nand U2562 (N_2562,In_561,In_360);
and U2563 (N_2563,In_744,In_219);
nor U2564 (N_2564,In_864,In_176);
and U2565 (N_2565,In_104,In_502);
xor U2566 (N_2566,In_257,In_477);
nand U2567 (N_2567,In_492,In_450);
nand U2568 (N_2568,In_547,In_766);
nor U2569 (N_2569,In_433,In_343);
nor U2570 (N_2570,In_779,In_715);
xnor U2571 (N_2571,In_523,In_380);
and U2572 (N_2572,In_916,In_707);
nor U2573 (N_2573,In_373,In_110);
nand U2574 (N_2574,In_1,In_333);
and U2575 (N_2575,In_968,In_256);
nand U2576 (N_2576,In_883,In_809);
and U2577 (N_2577,In_39,In_671);
nand U2578 (N_2578,In_936,In_647);
or U2579 (N_2579,In_354,In_53);
nand U2580 (N_2580,In_692,In_545);
and U2581 (N_2581,In_549,In_886);
xnor U2582 (N_2582,In_323,In_149);
or U2583 (N_2583,In_413,In_903);
nor U2584 (N_2584,In_137,In_733);
xnor U2585 (N_2585,In_240,In_788);
nor U2586 (N_2586,In_98,In_28);
and U2587 (N_2587,In_812,In_563);
and U2588 (N_2588,In_889,In_191);
and U2589 (N_2589,In_556,In_796);
nand U2590 (N_2590,In_343,In_368);
nand U2591 (N_2591,In_21,In_895);
or U2592 (N_2592,In_740,In_457);
nand U2593 (N_2593,In_291,In_364);
nor U2594 (N_2594,In_379,In_357);
xnor U2595 (N_2595,In_508,In_483);
nor U2596 (N_2596,In_897,In_378);
xor U2597 (N_2597,In_772,In_233);
nor U2598 (N_2598,In_786,In_495);
nand U2599 (N_2599,In_642,In_637);
or U2600 (N_2600,In_43,In_714);
nand U2601 (N_2601,In_776,In_983);
nor U2602 (N_2602,In_358,In_767);
nand U2603 (N_2603,In_246,In_542);
nand U2604 (N_2604,In_286,In_465);
and U2605 (N_2605,In_58,In_361);
xor U2606 (N_2606,In_714,In_642);
nand U2607 (N_2607,In_711,In_101);
and U2608 (N_2608,In_529,In_417);
nor U2609 (N_2609,In_95,In_759);
nand U2610 (N_2610,In_92,In_486);
or U2611 (N_2611,In_229,In_441);
and U2612 (N_2612,In_930,In_63);
or U2613 (N_2613,In_312,In_28);
or U2614 (N_2614,In_8,In_217);
or U2615 (N_2615,In_875,In_499);
nand U2616 (N_2616,In_99,In_723);
nand U2617 (N_2617,In_664,In_997);
nor U2618 (N_2618,In_281,In_702);
xnor U2619 (N_2619,In_91,In_159);
nor U2620 (N_2620,In_304,In_700);
xor U2621 (N_2621,In_115,In_901);
nand U2622 (N_2622,In_322,In_999);
xnor U2623 (N_2623,In_501,In_742);
nand U2624 (N_2624,In_651,In_438);
xor U2625 (N_2625,In_187,In_967);
xnor U2626 (N_2626,In_8,In_589);
xor U2627 (N_2627,In_33,In_765);
or U2628 (N_2628,In_701,In_616);
or U2629 (N_2629,In_283,In_128);
xnor U2630 (N_2630,In_70,In_17);
nor U2631 (N_2631,In_873,In_721);
and U2632 (N_2632,In_434,In_203);
and U2633 (N_2633,In_459,In_993);
nor U2634 (N_2634,In_769,In_854);
or U2635 (N_2635,In_427,In_96);
xor U2636 (N_2636,In_618,In_889);
nor U2637 (N_2637,In_911,In_308);
nand U2638 (N_2638,In_797,In_98);
nor U2639 (N_2639,In_490,In_341);
nand U2640 (N_2640,In_804,In_38);
or U2641 (N_2641,In_261,In_947);
and U2642 (N_2642,In_458,In_813);
and U2643 (N_2643,In_211,In_129);
nor U2644 (N_2644,In_776,In_477);
or U2645 (N_2645,In_268,In_389);
xor U2646 (N_2646,In_160,In_557);
xnor U2647 (N_2647,In_511,In_96);
nor U2648 (N_2648,In_366,In_862);
or U2649 (N_2649,In_817,In_18);
or U2650 (N_2650,In_270,In_140);
nand U2651 (N_2651,In_683,In_559);
nand U2652 (N_2652,In_104,In_163);
or U2653 (N_2653,In_235,In_998);
and U2654 (N_2654,In_487,In_660);
xor U2655 (N_2655,In_429,In_774);
xnor U2656 (N_2656,In_647,In_870);
or U2657 (N_2657,In_361,In_341);
nor U2658 (N_2658,In_356,In_301);
nand U2659 (N_2659,In_689,In_664);
nand U2660 (N_2660,In_775,In_65);
nor U2661 (N_2661,In_566,In_410);
nand U2662 (N_2662,In_409,In_951);
or U2663 (N_2663,In_59,In_997);
or U2664 (N_2664,In_188,In_603);
or U2665 (N_2665,In_468,In_143);
or U2666 (N_2666,In_473,In_64);
and U2667 (N_2667,In_876,In_560);
nor U2668 (N_2668,In_163,In_646);
nand U2669 (N_2669,In_105,In_760);
nand U2670 (N_2670,In_133,In_851);
nand U2671 (N_2671,In_101,In_100);
nand U2672 (N_2672,In_148,In_356);
nand U2673 (N_2673,In_846,In_33);
nand U2674 (N_2674,In_16,In_352);
xor U2675 (N_2675,In_37,In_899);
or U2676 (N_2676,In_648,In_67);
and U2677 (N_2677,In_347,In_609);
nand U2678 (N_2678,In_400,In_342);
nand U2679 (N_2679,In_801,In_330);
nand U2680 (N_2680,In_447,In_790);
xnor U2681 (N_2681,In_929,In_352);
or U2682 (N_2682,In_837,In_159);
or U2683 (N_2683,In_949,In_465);
or U2684 (N_2684,In_814,In_6);
xor U2685 (N_2685,In_383,In_72);
and U2686 (N_2686,In_258,In_726);
and U2687 (N_2687,In_388,In_984);
nor U2688 (N_2688,In_158,In_214);
nand U2689 (N_2689,In_603,In_196);
nand U2690 (N_2690,In_23,In_572);
xor U2691 (N_2691,In_204,In_936);
xor U2692 (N_2692,In_803,In_772);
xor U2693 (N_2693,In_727,In_492);
or U2694 (N_2694,In_962,In_422);
nand U2695 (N_2695,In_914,In_175);
or U2696 (N_2696,In_734,In_436);
and U2697 (N_2697,In_635,In_306);
nand U2698 (N_2698,In_357,In_1);
nor U2699 (N_2699,In_235,In_937);
xnor U2700 (N_2700,In_955,In_854);
nor U2701 (N_2701,In_343,In_367);
and U2702 (N_2702,In_659,In_103);
xnor U2703 (N_2703,In_237,In_741);
and U2704 (N_2704,In_168,In_17);
or U2705 (N_2705,In_300,In_239);
nand U2706 (N_2706,In_288,In_123);
nor U2707 (N_2707,In_41,In_553);
or U2708 (N_2708,In_373,In_260);
xnor U2709 (N_2709,In_895,In_748);
xnor U2710 (N_2710,In_263,In_14);
xor U2711 (N_2711,In_376,In_5);
nor U2712 (N_2712,In_785,In_262);
or U2713 (N_2713,In_319,In_477);
nor U2714 (N_2714,In_851,In_20);
nor U2715 (N_2715,In_182,In_799);
xor U2716 (N_2716,In_709,In_806);
and U2717 (N_2717,In_712,In_168);
and U2718 (N_2718,In_535,In_532);
or U2719 (N_2719,In_130,In_475);
or U2720 (N_2720,In_58,In_880);
or U2721 (N_2721,In_771,In_46);
or U2722 (N_2722,In_220,In_992);
nand U2723 (N_2723,In_66,In_28);
or U2724 (N_2724,In_820,In_244);
nor U2725 (N_2725,In_745,In_631);
xnor U2726 (N_2726,In_576,In_970);
xnor U2727 (N_2727,In_168,In_30);
xnor U2728 (N_2728,In_247,In_434);
xnor U2729 (N_2729,In_597,In_241);
and U2730 (N_2730,In_158,In_227);
and U2731 (N_2731,In_155,In_921);
nand U2732 (N_2732,In_635,In_294);
or U2733 (N_2733,In_270,In_520);
nand U2734 (N_2734,In_775,In_307);
or U2735 (N_2735,In_513,In_343);
nor U2736 (N_2736,In_441,In_699);
nand U2737 (N_2737,In_309,In_526);
and U2738 (N_2738,In_700,In_104);
nor U2739 (N_2739,In_419,In_15);
nand U2740 (N_2740,In_956,In_952);
nand U2741 (N_2741,In_772,In_384);
or U2742 (N_2742,In_313,In_594);
nor U2743 (N_2743,In_87,In_192);
and U2744 (N_2744,In_325,In_494);
and U2745 (N_2745,In_777,In_955);
and U2746 (N_2746,In_496,In_793);
nand U2747 (N_2747,In_167,In_164);
or U2748 (N_2748,In_658,In_736);
and U2749 (N_2749,In_422,In_813);
xnor U2750 (N_2750,In_197,In_757);
and U2751 (N_2751,In_614,In_935);
nand U2752 (N_2752,In_178,In_862);
nor U2753 (N_2753,In_327,In_964);
or U2754 (N_2754,In_641,In_783);
xor U2755 (N_2755,In_880,In_145);
or U2756 (N_2756,In_550,In_375);
nor U2757 (N_2757,In_545,In_842);
nand U2758 (N_2758,In_104,In_177);
and U2759 (N_2759,In_103,In_273);
nor U2760 (N_2760,In_163,In_463);
xnor U2761 (N_2761,In_615,In_339);
and U2762 (N_2762,In_749,In_879);
nor U2763 (N_2763,In_736,In_879);
xor U2764 (N_2764,In_869,In_967);
nand U2765 (N_2765,In_648,In_287);
and U2766 (N_2766,In_647,In_635);
xor U2767 (N_2767,In_283,In_577);
nor U2768 (N_2768,In_830,In_7);
nand U2769 (N_2769,In_790,In_976);
nand U2770 (N_2770,In_953,In_686);
xor U2771 (N_2771,In_412,In_894);
or U2772 (N_2772,In_782,In_118);
or U2773 (N_2773,In_939,In_118);
or U2774 (N_2774,In_110,In_697);
nor U2775 (N_2775,In_810,In_509);
or U2776 (N_2776,In_403,In_446);
nand U2777 (N_2777,In_217,In_354);
xor U2778 (N_2778,In_465,In_9);
xnor U2779 (N_2779,In_3,In_434);
and U2780 (N_2780,In_831,In_147);
or U2781 (N_2781,In_257,In_633);
or U2782 (N_2782,In_34,In_780);
xnor U2783 (N_2783,In_988,In_708);
xnor U2784 (N_2784,In_826,In_994);
nor U2785 (N_2785,In_455,In_534);
nor U2786 (N_2786,In_355,In_769);
nor U2787 (N_2787,In_337,In_690);
xnor U2788 (N_2788,In_858,In_662);
xnor U2789 (N_2789,In_611,In_47);
nor U2790 (N_2790,In_492,In_766);
and U2791 (N_2791,In_721,In_223);
or U2792 (N_2792,In_109,In_378);
nor U2793 (N_2793,In_143,In_169);
nor U2794 (N_2794,In_716,In_545);
nor U2795 (N_2795,In_612,In_328);
nand U2796 (N_2796,In_570,In_359);
nor U2797 (N_2797,In_404,In_566);
and U2798 (N_2798,In_209,In_366);
nor U2799 (N_2799,In_257,In_111);
nor U2800 (N_2800,In_298,In_837);
nor U2801 (N_2801,In_318,In_788);
and U2802 (N_2802,In_432,In_682);
or U2803 (N_2803,In_873,In_288);
and U2804 (N_2804,In_184,In_540);
nor U2805 (N_2805,In_485,In_84);
or U2806 (N_2806,In_603,In_869);
nand U2807 (N_2807,In_743,In_28);
and U2808 (N_2808,In_584,In_976);
nand U2809 (N_2809,In_973,In_823);
xnor U2810 (N_2810,In_778,In_756);
nor U2811 (N_2811,In_914,In_917);
xor U2812 (N_2812,In_698,In_939);
xor U2813 (N_2813,In_942,In_771);
xor U2814 (N_2814,In_469,In_892);
nand U2815 (N_2815,In_871,In_176);
nand U2816 (N_2816,In_506,In_380);
nor U2817 (N_2817,In_371,In_96);
or U2818 (N_2818,In_55,In_138);
xnor U2819 (N_2819,In_343,In_27);
or U2820 (N_2820,In_512,In_427);
nor U2821 (N_2821,In_149,In_614);
nand U2822 (N_2822,In_388,In_276);
and U2823 (N_2823,In_254,In_737);
and U2824 (N_2824,In_798,In_478);
nand U2825 (N_2825,In_529,In_293);
nand U2826 (N_2826,In_783,In_659);
nor U2827 (N_2827,In_612,In_460);
nand U2828 (N_2828,In_139,In_121);
xnor U2829 (N_2829,In_396,In_77);
or U2830 (N_2830,In_931,In_5);
nand U2831 (N_2831,In_329,In_883);
nor U2832 (N_2832,In_743,In_579);
or U2833 (N_2833,In_106,In_530);
nand U2834 (N_2834,In_501,In_641);
nor U2835 (N_2835,In_466,In_647);
nor U2836 (N_2836,In_68,In_554);
or U2837 (N_2837,In_708,In_328);
xnor U2838 (N_2838,In_759,In_33);
xnor U2839 (N_2839,In_489,In_627);
or U2840 (N_2840,In_864,In_257);
nand U2841 (N_2841,In_715,In_144);
and U2842 (N_2842,In_215,In_625);
or U2843 (N_2843,In_393,In_29);
and U2844 (N_2844,In_194,In_965);
xnor U2845 (N_2845,In_125,In_656);
and U2846 (N_2846,In_723,In_804);
or U2847 (N_2847,In_416,In_854);
nand U2848 (N_2848,In_56,In_553);
and U2849 (N_2849,In_92,In_686);
and U2850 (N_2850,In_397,In_201);
nand U2851 (N_2851,In_365,In_257);
nor U2852 (N_2852,In_981,In_842);
or U2853 (N_2853,In_785,In_939);
and U2854 (N_2854,In_376,In_829);
xor U2855 (N_2855,In_48,In_780);
and U2856 (N_2856,In_750,In_854);
xnor U2857 (N_2857,In_855,In_373);
and U2858 (N_2858,In_530,In_244);
nor U2859 (N_2859,In_130,In_855);
or U2860 (N_2860,In_232,In_929);
and U2861 (N_2861,In_294,In_657);
xor U2862 (N_2862,In_255,In_362);
and U2863 (N_2863,In_458,In_290);
and U2864 (N_2864,In_739,In_998);
xor U2865 (N_2865,In_7,In_651);
xnor U2866 (N_2866,In_413,In_659);
nor U2867 (N_2867,In_972,In_766);
xor U2868 (N_2868,In_76,In_684);
xor U2869 (N_2869,In_0,In_483);
nor U2870 (N_2870,In_53,In_10);
or U2871 (N_2871,In_480,In_512);
nand U2872 (N_2872,In_785,In_380);
nand U2873 (N_2873,In_499,In_153);
nand U2874 (N_2874,In_363,In_562);
nand U2875 (N_2875,In_446,In_492);
nor U2876 (N_2876,In_994,In_589);
and U2877 (N_2877,In_676,In_44);
nor U2878 (N_2878,In_690,In_908);
and U2879 (N_2879,In_902,In_488);
and U2880 (N_2880,In_890,In_556);
xnor U2881 (N_2881,In_898,In_806);
nand U2882 (N_2882,In_858,In_794);
nand U2883 (N_2883,In_513,In_478);
nand U2884 (N_2884,In_86,In_228);
nor U2885 (N_2885,In_326,In_930);
nor U2886 (N_2886,In_53,In_22);
and U2887 (N_2887,In_68,In_155);
or U2888 (N_2888,In_620,In_630);
and U2889 (N_2889,In_422,In_665);
or U2890 (N_2890,In_181,In_541);
and U2891 (N_2891,In_676,In_149);
nand U2892 (N_2892,In_380,In_350);
and U2893 (N_2893,In_391,In_356);
nor U2894 (N_2894,In_186,In_216);
xnor U2895 (N_2895,In_937,In_230);
nor U2896 (N_2896,In_595,In_996);
nand U2897 (N_2897,In_277,In_933);
nor U2898 (N_2898,In_784,In_605);
xnor U2899 (N_2899,In_265,In_22);
or U2900 (N_2900,In_138,In_153);
nand U2901 (N_2901,In_295,In_546);
nor U2902 (N_2902,In_697,In_842);
and U2903 (N_2903,In_496,In_191);
or U2904 (N_2904,In_414,In_94);
nand U2905 (N_2905,In_368,In_799);
and U2906 (N_2906,In_184,In_954);
nand U2907 (N_2907,In_995,In_919);
xor U2908 (N_2908,In_60,In_301);
or U2909 (N_2909,In_704,In_827);
nand U2910 (N_2910,In_209,In_126);
or U2911 (N_2911,In_199,In_493);
nor U2912 (N_2912,In_122,In_924);
and U2913 (N_2913,In_789,In_867);
nand U2914 (N_2914,In_459,In_859);
and U2915 (N_2915,In_273,In_682);
nor U2916 (N_2916,In_254,In_567);
nand U2917 (N_2917,In_661,In_81);
and U2918 (N_2918,In_554,In_628);
xnor U2919 (N_2919,In_212,In_380);
xnor U2920 (N_2920,In_28,In_282);
nand U2921 (N_2921,In_107,In_645);
and U2922 (N_2922,In_159,In_211);
nor U2923 (N_2923,In_967,In_61);
or U2924 (N_2924,In_757,In_556);
xnor U2925 (N_2925,In_185,In_287);
and U2926 (N_2926,In_248,In_619);
or U2927 (N_2927,In_722,In_284);
nor U2928 (N_2928,In_695,In_81);
xnor U2929 (N_2929,In_69,In_739);
nand U2930 (N_2930,In_395,In_398);
nor U2931 (N_2931,In_970,In_306);
nand U2932 (N_2932,In_855,In_534);
xnor U2933 (N_2933,In_49,In_777);
or U2934 (N_2934,In_784,In_695);
and U2935 (N_2935,In_658,In_111);
xnor U2936 (N_2936,In_386,In_339);
nor U2937 (N_2937,In_388,In_267);
or U2938 (N_2938,In_531,In_810);
and U2939 (N_2939,In_885,In_486);
or U2940 (N_2940,In_379,In_485);
nand U2941 (N_2941,In_662,In_818);
or U2942 (N_2942,In_75,In_299);
nand U2943 (N_2943,In_354,In_907);
and U2944 (N_2944,In_551,In_2);
and U2945 (N_2945,In_665,In_396);
nor U2946 (N_2946,In_511,In_205);
and U2947 (N_2947,In_64,In_910);
or U2948 (N_2948,In_83,In_711);
xnor U2949 (N_2949,In_211,In_11);
or U2950 (N_2950,In_852,In_613);
nand U2951 (N_2951,In_229,In_433);
nor U2952 (N_2952,In_152,In_940);
nand U2953 (N_2953,In_957,In_202);
nor U2954 (N_2954,In_526,In_138);
or U2955 (N_2955,In_619,In_925);
xor U2956 (N_2956,In_156,In_421);
and U2957 (N_2957,In_299,In_768);
or U2958 (N_2958,In_411,In_668);
and U2959 (N_2959,In_708,In_625);
nor U2960 (N_2960,In_868,In_362);
and U2961 (N_2961,In_549,In_36);
nand U2962 (N_2962,In_116,In_201);
or U2963 (N_2963,In_280,In_464);
xnor U2964 (N_2964,In_824,In_222);
or U2965 (N_2965,In_746,In_715);
nand U2966 (N_2966,In_889,In_655);
nor U2967 (N_2967,In_563,In_313);
or U2968 (N_2968,In_392,In_43);
nand U2969 (N_2969,In_110,In_628);
nor U2970 (N_2970,In_558,In_707);
and U2971 (N_2971,In_221,In_305);
or U2972 (N_2972,In_601,In_555);
or U2973 (N_2973,In_254,In_223);
nor U2974 (N_2974,In_108,In_917);
and U2975 (N_2975,In_949,In_889);
and U2976 (N_2976,In_420,In_889);
xnor U2977 (N_2977,In_121,In_850);
nand U2978 (N_2978,In_290,In_995);
and U2979 (N_2979,In_58,In_982);
xor U2980 (N_2980,In_71,In_802);
or U2981 (N_2981,In_69,In_134);
xor U2982 (N_2982,In_251,In_354);
nor U2983 (N_2983,In_212,In_368);
xnor U2984 (N_2984,In_218,In_653);
nand U2985 (N_2985,In_559,In_648);
and U2986 (N_2986,In_209,In_915);
nand U2987 (N_2987,In_404,In_791);
nor U2988 (N_2988,In_881,In_763);
nand U2989 (N_2989,In_877,In_738);
or U2990 (N_2990,In_529,In_801);
nand U2991 (N_2991,In_336,In_341);
and U2992 (N_2992,In_382,In_309);
nor U2993 (N_2993,In_763,In_493);
and U2994 (N_2994,In_523,In_29);
nand U2995 (N_2995,In_124,In_861);
nand U2996 (N_2996,In_829,In_510);
or U2997 (N_2997,In_132,In_950);
nor U2998 (N_2998,In_119,In_255);
or U2999 (N_2999,In_803,In_853);
or U3000 (N_3000,In_692,In_408);
or U3001 (N_3001,In_237,In_292);
nor U3002 (N_3002,In_434,In_667);
nand U3003 (N_3003,In_393,In_676);
nand U3004 (N_3004,In_221,In_375);
and U3005 (N_3005,In_102,In_342);
or U3006 (N_3006,In_948,In_736);
and U3007 (N_3007,In_82,In_899);
nand U3008 (N_3008,In_34,In_267);
or U3009 (N_3009,In_659,In_870);
or U3010 (N_3010,In_504,In_372);
nor U3011 (N_3011,In_813,In_497);
and U3012 (N_3012,In_43,In_208);
nand U3013 (N_3013,In_633,In_40);
or U3014 (N_3014,In_762,In_502);
nor U3015 (N_3015,In_254,In_6);
xnor U3016 (N_3016,In_627,In_119);
and U3017 (N_3017,In_671,In_439);
xor U3018 (N_3018,In_755,In_444);
and U3019 (N_3019,In_513,In_477);
and U3020 (N_3020,In_712,In_301);
nand U3021 (N_3021,In_664,In_915);
nand U3022 (N_3022,In_507,In_442);
nand U3023 (N_3023,In_24,In_910);
xor U3024 (N_3024,In_221,In_754);
xor U3025 (N_3025,In_975,In_539);
xnor U3026 (N_3026,In_749,In_713);
nand U3027 (N_3027,In_490,In_783);
nand U3028 (N_3028,In_215,In_323);
xnor U3029 (N_3029,In_602,In_480);
nand U3030 (N_3030,In_466,In_264);
nor U3031 (N_3031,In_858,In_888);
xnor U3032 (N_3032,In_175,In_59);
xor U3033 (N_3033,In_197,In_556);
and U3034 (N_3034,In_858,In_549);
nand U3035 (N_3035,In_161,In_851);
and U3036 (N_3036,In_905,In_152);
xor U3037 (N_3037,In_759,In_226);
nor U3038 (N_3038,In_583,In_83);
xnor U3039 (N_3039,In_437,In_116);
nor U3040 (N_3040,In_70,In_419);
xnor U3041 (N_3041,In_372,In_390);
nor U3042 (N_3042,In_12,In_982);
or U3043 (N_3043,In_346,In_131);
nand U3044 (N_3044,In_661,In_187);
nand U3045 (N_3045,In_841,In_850);
and U3046 (N_3046,In_677,In_739);
nor U3047 (N_3047,In_331,In_297);
nor U3048 (N_3048,In_63,In_831);
nor U3049 (N_3049,In_606,In_910);
nor U3050 (N_3050,In_46,In_599);
or U3051 (N_3051,In_60,In_906);
xnor U3052 (N_3052,In_446,In_879);
nor U3053 (N_3053,In_872,In_517);
nand U3054 (N_3054,In_706,In_716);
or U3055 (N_3055,In_32,In_158);
nand U3056 (N_3056,In_368,In_606);
and U3057 (N_3057,In_120,In_580);
nor U3058 (N_3058,In_566,In_439);
xnor U3059 (N_3059,In_163,In_258);
nor U3060 (N_3060,In_793,In_799);
or U3061 (N_3061,In_918,In_934);
xnor U3062 (N_3062,In_305,In_223);
or U3063 (N_3063,In_508,In_313);
nand U3064 (N_3064,In_231,In_2);
xor U3065 (N_3065,In_708,In_11);
and U3066 (N_3066,In_402,In_328);
and U3067 (N_3067,In_297,In_473);
and U3068 (N_3068,In_232,In_859);
nor U3069 (N_3069,In_998,In_253);
and U3070 (N_3070,In_736,In_257);
and U3071 (N_3071,In_916,In_418);
xor U3072 (N_3072,In_437,In_239);
xnor U3073 (N_3073,In_936,In_565);
nand U3074 (N_3074,In_833,In_566);
nor U3075 (N_3075,In_885,In_644);
nor U3076 (N_3076,In_34,In_1);
nor U3077 (N_3077,In_580,In_813);
nand U3078 (N_3078,In_351,In_340);
nor U3079 (N_3079,In_286,In_348);
and U3080 (N_3080,In_365,In_366);
nand U3081 (N_3081,In_194,In_787);
nand U3082 (N_3082,In_398,In_866);
xor U3083 (N_3083,In_392,In_213);
and U3084 (N_3084,In_171,In_824);
nand U3085 (N_3085,In_321,In_943);
nand U3086 (N_3086,In_98,In_698);
or U3087 (N_3087,In_479,In_35);
nand U3088 (N_3088,In_556,In_510);
and U3089 (N_3089,In_457,In_4);
nand U3090 (N_3090,In_840,In_260);
xnor U3091 (N_3091,In_67,In_254);
and U3092 (N_3092,In_743,In_554);
and U3093 (N_3093,In_326,In_881);
xor U3094 (N_3094,In_267,In_328);
nand U3095 (N_3095,In_396,In_219);
xnor U3096 (N_3096,In_77,In_162);
and U3097 (N_3097,In_739,In_730);
xor U3098 (N_3098,In_757,In_477);
xnor U3099 (N_3099,In_111,In_108);
or U3100 (N_3100,In_341,In_260);
nor U3101 (N_3101,In_271,In_108);
and U3102 (N_3102,In_879,In_450);
or U3103 (N_3103,In_493,In_515);
or U3104 (N_3104,In_302,In_305);
nor U3105 (N_3105,In_377,In_114);
nor U3106 (N_3106,In_701,In_745);
and U3107 (N_3107,In_595,In_797);
xnor U3108 (N_3108,In_128,In_204);
nand U3109 (N_3109,In_20,In_650);
nand U3110 (N_3110,In_398,In_303);
and U3111 (N_3111,In_332,In_35);
and U3112 (N_3112,In_123,In_271);
and U3113 (N_3113,In_893,In_272);
xnor U3114 (N_3114,In_677,In_870);
or U3115 (N_3115,In_322,In_915);
and U3116 (N_3116,In_504,In_535);
xor U3117 (N_3117,In_826,In_52);
xor U3118 (N_3118,In_741,In_191);
xor U3119 (N_3119,In_338,In_162);
xor U3120 (N_3120,In_935,In_748);
nor U3121 (N_3121,In_655,In_262);
and U3122 (N_3122,In_383,In_795);
or U3123 (N_3123,In_665,In_530);
nor U3124 (N_3124,In_472,In_652);
nor U3125 (N_3125,In_756,In_959);
nand U3126 (N_3126,In_441,In_582);
xnor U3127 (N_3127,In_18,In_622);
and U3128 (N_3128,In_658,In_777);
or U3129 (N_3129,In_158,In_257);
nor U3130 (N_3130,In_409,In_837);
or U3131 (N_3131,In_384,In_947);
nand U3132 (N_3132,In_453,In_664);
nand U3133 (N_3133,In_20,In_839);
xor U3134 (N_3134,In_630,In_385);
nand U3135 (N_3135,In_64,In_876);
and U3136 (N_3136,In_849,In_665);
nand U3137 (N_3137,In_671,In_749);
or U3138 (N_3138,In_269,In_642);
or U3139 (N_3139,In_133,In_435);
or U3140 (N_3140,In_847,In_684);
nor U3141 (N_3141,In_287,In_166);
xnor U3142 (N_3142,In_321,In_293);
nand U3143 (N_3143,In_925,In_131);
or U3144 (N_3144,In_234,In_552);
nor U3145 (N_3145,In_366,In_711);
and U3146 (N_3146,In_670,In_113);
and U3147 (N_3147,In_610,In_861);
and U3148 (N_3148,In_365,In_644);
nand U3149 (N_3149,In_569,In_192);
xnor U3150 (N_3150,In_32,In_298);
nand U3151 (N_3151,In_928,In_789);
and U3152 (N_3152,In_856,In_500);
or U3153 (N_3153,In_943,In_414);
nand U3154 (N_3154,In_590,In_961);
nor U3155 (N_3155,In_173,In_790);
nor U3156 (N_3156,In_917,In_40);
xnor U3157 (N_3157,In_322,In_895);
nand U3158 (N_3158,In_624,In_665);
nand U3159 (N_3159,In_973,In_906);
nor U3160 (N_3160,In_178,In_415);
nand U3161 (N_3161,In_990,In_801);
and U3162 (N_3162,In_173,In_419);
xor U3163 (N_3163,In_261,In_338);
or U3164 (N_3164,In_216,In_289);
nand U3165 (N_3165,In_907,In_585);
xnor U3166 (N_3166,In_960,In_444);
nor U3167 (N_3167,In_878,In_82);
and U3168 (N_3168,In_488,In_526);
nor U3169 (N_3169,In_114,In_585);
nand U3170 (N_3170,In_852,In_63);
nor U3171 (N_3171,In_673,In_393);
nor U3172 (N_3172,In_461,In_24);
or U3173 (N_3173,In_325,In_912);
nor U3174 (N_3174,In_202,In_656);
and U3175 (N_3175,In_652,In_254);
nand U3176 (N_3176,In_907,In_997);
or U3177 (N_3177,In_629,In_772);
nor U3178 (N_3178,In_869,In_625);
nand U3179 (N_3179,In_183,In_689);
and U3180 (N_3180,In_437,In_943);
and U3181 (N_3181,In_264,In_117);
or U3182 (N_3182,In_907,In_232);
or U3183 (N_3183,In_156,In_241);
nor U3184 (N_3184,In_327,In_939);
nand U3185 (N_3185,In_235,In_43);
or U3186 (N_3186,In_132,In_262);
xor U3187 (N_3187,In_933,In_718);
or U3188 (N_3188,In_879,In_401);
xnor U3189 (N_3189,In_958,In_117);
nand U3190 (N_3190,In_674,In_778);
xnor U3191 (N_3191,In_103,In_243);
nor U3192 (N_3192,In_374,In_186);
nor U3193 (N_3193,In_788,In_174);
nand U3194 (N_3194,In_313,In_418);
or U3195 (N_3195,In_640,In_181);
xor U3196 (N_3196,In_813,In_819);
and U3197 (N_3197,In_632,In_163);
xnor U3198 (N_3198,In_629,In_984);
or U3199 (N_3199,In_888,In_92);
nand U3200 (N_3200,In_680,In_717);
xnor U3201 (N_3201,In_322,In_209);
xor U3202 (N_3202,In_461,In_932);
nand U3203 (N_3203,In_278,In_196);
nand U3204 (N_3204,In_76,In_889);
nand U3205 (N_3205,In_798,In_544);
nor U3206 (N_3206,In_612,In_875);
xnor U3207 (N_3207,In_372,In_0);
xnor U3208 (N_3208,In_48,In_915);
xor U3209 (N_3209,In_335,In_922);
xnor U3210 (N_3210,In_967,In_58);
and U3211 (N_3211,In_588,In_40);
nand U3212 (N_3212,In_578,In_320);
xnor U3213 (N_3213,In_809,In_723);
nand U3214 (N_3214,In_351,In_764);
xnor U3215 (N_3215,In_558,In_634);
and U3216 (N_3216,In_314,In_939);
or U3217 (N_3217,In_223,In_585);
nand U3218 (N_3218,In_386,In_356);
xor U3219 (N_3219,In_648,In_518);
xnor U3220 (N_3220,In_897,In_778);
xor U3221 (N_3221,In_124,In_728);
xnor U3222 (N_3222,In_812,In_43);
and U3223 (N_3223,In_14,In_176);
nand U3224 (N_3224,In_841,In_381);
or U3225 (N_3225,In_627,In_696);
xnor U3226 (N_3226,In_2,In_981);
xnor U3227 (N_3227,In_501,In_390);
nor U3228 (N_3228,In_470,In_889);
xor U3229 (N_3229,In_478,In_681);
and U3230 (N_3230,In_826,In_291);
or U3231 (N_3231,In_176,In_458);
xnor U3232 (N_3232,In_366,In_718);
xnor U3233 (N_3233,In_854,In_140);
or U3234 (N_3234,In_293,In_369);
xor U3235 (N_3235,In_224,In_112);
or U3236 (N_3236,In_922,In_188);
nand U3237 (N_3237,In_242,In_157);
xnor U3238 (N_3238,In_740,In_729);
and U3239 (N_3239,In_64,In_520);
xor U3240 (N_3240,In_493,In_695);
xor U3241 (N_3241,In_573,In_2);
nor U3242 (N_3242,In_134,In_114);
nand U3243 (N_3243,In_899,In_322);
and U3244 (N_3244,In_799,In_752);
nand U3245 (N_3245,In_144,In_947);
or U3246 (N_3246,In_911,In_994);
or U3247 (N_3247,In_688,In_815);
nor U3248 (N_3248,In_648,In_238);
and U3249 (N_3249,In_34,In_161);
and U3250 (N_3250,In_112,In_792);
nand U3251 (N_3251,In_981,In_105);
nor U3252 (N_3252,In_869,In_836);
nor U3253 (N_3253,In_552,In_328);
xnor U3254 (N_3254,In_111,In_748);
or U3255 (N_3255,In_927,In_837);
or U3256 (N_3256,In_595,In_280);
nor U3257 (N_3257,In_213,In_338);
nor U3258 (N_3258,In_610,In_379);
xor U3259 (N_3259,In_626,In_549);
xnor U3260 (N_3260,In_796,In_65);
nor U3261 (N_3261,In_119,In_742);
nand U3262 (N_3262,In_228,In_59);
nor U3263 (N_3263,In_210,In_805);
nor U3264 (N_3264,In_485,In_877);
xor U3265 (N_3265,In_970,In_42);
nor U3266 (N_3266,In_92,In_559);
or U3267 (N_3267,In_623,In_750);
nor U3268 (N_3268,In_228,In_600);
and U3269 (N_3269,In_759,In_855);
xor U3270 (N_3270,In_421,In_340);
xor U3271 (N_3271,In_48,In_527);
xor U3272 (N_3272,In_353,In_556);
nand U3273 (N_3273,In_32,In_367);
nand U3274 (N_3274,In_947,In_788);
xnor U3275 (N_3275,In_478,In_880);
nor U3276 (N_3276,In_34,In_546);
or U3277 (N_3277,In_715,In_858);
or U3278 (N_3278,In_575,In_26);
or U3279 (N_3279,In_461,In_43);
or U3280 (N_3280,In_322,In_116);
nand U3281 (N_3281,In_9,In_1);
or U3282 (N_3282,In_941,In_409);
nor U3283 (N_3283,In_737,In_622);
or U3284 (N_3284,In_361,In_117);
nor U3285 (N_3285,In_358,In_911);
and U3286 (N_3286,In_305,In_950);
and U3287 (N_3287,In_147,In_974);
nor U3288 (N_3288,In_93,In_291);
or U3289 (N_3289,In_454,In_519);
xor U3290 (N_3290,In_349,In_128);
nand U3291 (N_3291,In_941,In_324);
xor U3292 (N_3292,In_353,In_564);
xor U3293 (N_3293,In_44,In_297);
or U3294 (N_3294,In_456,In_568);
and U3295 (N_3295,In_940,In_596);
and U3296 (N_3296,In_267,In_542);
xnor U3297 (N_3297,In_910,In_890);
or U3298 (N_3298,In_197,In_746);
or U3299 (N_3299,In_594,In_792);
nand U3300 (N_3300,In_953,In_207);
or U3301 (N_3301,In_951,In_968);
nand U3302 (N_3302,In_427,In_307);
and U3303 (N_3303,In_775,In_291);
nor U3304 (N_3304,In_999,In_761);
nor U3305 (N_3305,In_2,In_751);
nand U3306 (N_3306,In_776,In_496);
and U3307 (N_3307,In_858,In_103);
and U3308 (N_3308,In_943,In_311);
or U3309 (N_3309,In_426,In_398);
nor U3310 (N_3310,In_467,In_79);
xnor U3311 (N_3311,In_933,In_73);
nor U3312 (N_3312,In_605,In_140);
nor U3313 (N_3313,In_705,In_835);
or U3314 (N_3314,In_611,In_890);
nor U3315 (N_3315,In_239,In_592);
or U3316 (N_3316,In_24,In_978);
nor U3317 (N_3317,In_461,In_661);
nor U3318 (N_3318,In_913,In_354);
nor U3319 (N_3319,In_823,In_625);
or U3320 (N_3320,In_976,In_537);
and U3321 (N_3321,In_714,In_684);
or U3322 (N_3322,In_837,In_177);
and U3323 (N_3323,In_570,In_913);
xnor U3324 (N_3324,In_517,In_472);
nor U3325 (N_3325,In_410,In_463);
nand U3326 (N_3326,In_110,In_720);
xnor U3327 (N_3327,In_45,In_464);
and U3328 (N_3328,In_426,In_331);
xor U3329 (N_3329,In_799,In_883);
or U3330 (N_3330,In_916,In_679);
or U3331 (N_3331,In_344,In_794);
nor U3332 (N_3332,In_320,In_787);
nand U3333 (N_3333,In_61,In_162);
xor U3334 (N_3334,In_612,In_229);
nor U3335 (N_3335,In_703,In_760);
or U3336 (N_3336,In_523,In_603);
nand U3337 (N_3337,In_153,In_119);
nand U3338 (N_3338,In_222,In_804);
or U3339 (N_3339,In_186,In_201);
and U3340 (N_3340,In_343,In_475);
and U3341 (N_3341,In_749,In_833);
nand U3342 (N_3342,In_320,In_442);
nand U3343 (N_3343,In_19,In_654);
xor U3344 (N_3344,In_353,In_771);
xnor U3345 (N_3345,In_508,In_213);
and U3346 (N_3346,In_298,In_931);
or U3347 (N_3347,In_514,In_244);
and U3348 (N_3348,In_649,In_39);
nor U3349 (N_3349,In_454,In_735);
and U3350 (N_3350,In_149,In_437);
nor U3351 (N_3351,In_644,In_737);
or U3352 (N_3352,In_247,In_410);
nand U3353 (N_3353,In_780,In_142);
nor U3354 (N_3354,In_892,In_483);
nand U3355 (N_3355,In_269,In_879);
or U3356 (N_3356,In_640,In_482);
nand U3357 (N_3357,In_946,In_253);
or U3358 (N_3358,In_261,In_614);
or U3359 (N_3359,In_932,In_328);
and U3360 (N_3360,In_86,In_649);
nor U3361 (N_3361,In_244,In_556);
or U3362 (N_3362,In_416,In_370);
nand U3363 (N_3363,In_364,In_565);
xnor U3364 (N_3364,In_562,In_713);
nor U3365 (N_3365,In_474,In_591);
nand U3366 (N_3366,In_495,In_124);
nand U3367 (N_3367,In_491,In_271);
nor U3368 (N_3368,In_833,In_570);
or U3369 (N_3369,In_63,In_465);
or U3370 (N_3370,In_972,In_394);
xnor U3371 (N_3371,In_51,In_893);
nand U3372 (N_3372,In_652,In_740);
xnor U3373 (N_3373,In_124,In_660);
nor U3374 (N_3374,In_505,In_607);
nor U3375 (N_3375,In_522,In_798);
or U3376 (N_3376,In_491,In_355);
xor U3377 (N_3377,In_571,In_266);
nand U3378 (N_3378,In_13,In_472);
xnor U3379 (N_3379,In_698,In_878);
xnor U3380 (N_3380,In_519,In_125);
or U3381 (N_3381,In_23,In_839);
xnor U3382 (N_3382,In_387,In_809);
or U3383 (N_3383,In_532,In_657);
nand U3384 (N_3384,In_243,In_833);
nor U3385 (N_3385,In_545,In_546);
and U3386 (N_3386,In_880,In_959);
and U3387 (N_3387,In_881,In_880);
xor U3388 (N_3388,In_963,In_102);
nor U3389 (N_3389,In_45,In_400);
and U3390 (N_3390,In_139,In_670);
and U3391 (N_3391,In_407,In_898);
or U3392 (N_3392,In_857,In_719);
or U3393 (N_3393,In_205,In_842);
and U3394 (N_3394,In_257,In_540);
or U3395 (N_3395,In_25,In_637);
nor U3396 (N_3396,In_329,In_662);
nor U3397 (N_3397,In_332,In_816);
or U3398 (N_3398,In_91,In_625);
nor U3399 (N_3399,In_121,In_215);
nor U3400 (N_3400,In_124,In_613);
xor U3401 (N_3401,In_908,In_496);
and U3402 (N_3402,In_384,In_615);
nor U3403 (N_3403,In_674,In_220);
nand U3404 (N_3404,In_80,In_243);
nor U3405 (N_3405,In_871,In_44);
and U3406 (N_3406,In_795,In_206);
nand U3407 (N_3407,In_20,In_711);
nor U3408 (N_3408,In_343,In_305);
nand U3409 (N_3409,In_599,In_327);
or U3410 (N_3410,In_104,In_283);
nor U3411 (N_3411,In_216,In_481);
or U3412 (N_3412,In_643,In_301);
xor U3413 (N_3413,In_355,In_423);
nand U3414 (N_3414,In_104,In_950);
or U3415 (N_3415,In_527,In_88);
or U3416 (N_3416,In_945,In_823);
and U3417 (N_3417,In_147,In_471);
nor U3418 (N_3418,In_992,In_213);
or U3419 (N_3419,In_97,In_232);
nand U3420 (N_3420,In_982,In_420);
or U3421 (N_3421,In_132,In_926);
xor U3422 (N_3422,In_451,In_842);
nand U3423 (N_3423,In_109,In_581);
nor U3424 (N_3424,In_946,In_703);
and U3425 (N_3425,In_885,In_978);
nand U3426 (N_3426,In_889,In_755);
nor U3427 (N_3427,In_667,In_70);
and U3428 (N_3428,In_153,In_695);
and U3429 (N_3429,In_80,In_749);
and U3430 (N_3430,In_507,In_745);
or U3431 (N_3431,In_426,In_746);
and U3432 (N_3432,In_704,In_264);
and U3433 (N_3433,In_45,In_175);
and U3434 (N_3434,In_764,In_282);
xnor U3435 (N_3435,In_65,In_56);
or U3436 (N_3436,In_434,In_430);
nor U3437 (N_3437,In_939,In_89);
nor U3438 (N_3438,In_539,In_474);
or U3439 (N_3439,In_844,In_858);
xor U3440 (N_3440,In_660,In_848);
xnor U3441 (N_3441,In_768,In_352);
and U3442 (N_3442,In_465,In_460);
or U3443 (N_3443,In_447,In_263);
or U3444 (N_3444,In_516,In_270);
nor U3445 (N_3445,In_779,In_477);
or U3446 (N_3446,In_479,In_32);
nor U3447 (N_3447,In_325,In_840);
nand U3448 (N_3448,In_456,In_279);
nand U3449 (N_3449,In_86,In_756);
xnor U3450 (N_3450,In_258,In_828);
and U3451 (N_3451,In_702,In_216);
and U3452 (N_3452,In_598,In_610);
nor U3453 (N_3453,In_533,In_351);
nor U3454 (N_3454,In_66,In_272);
nand U3455 (N_3455,In_100,In_696);
xor U3456 (N_3456,In_85,In_229);
nor U3457 (N_3457,In_954,In_224);
or U3458 (N_3458,In_179,In_520);
nor U3459 (N_3459,In_983,In_918);
nor U3460 (N_3460,In_201,In_700);
xor U3461 (N_3461,In_669,In_961);
xnor U3462 (N_3462,In_67,In_27);
nor U3463 (N_3463,In_912,In_896);
and U3464 (N_3464,In_342,In_254);
nor U3465 (N_3465,In_191,In_706);
or U3466 (N_3466,In_559,In_430);
and U3467 (N_3467,In_582,In_68);
xor U3468 (N_3468,In_512,In_581);
nor U3469 (N_3469,In_537,In_374);
xor U3470 (N_3470,In_699,In_808);
nand U3471 (N_3471,In_64,In_138);
nand U3472 (N_3472,In_100,In_228);
xor U3473 (N_3473,In_139,In_167);
and U3474 (N_3474,In_84,In_275);
xor U3475 (N_3475,In_799,In_581);
xnor U3476 (N_3476,In_420,In_276);
nor U3477 (N_3477,In_639,In_599);
or U3478 (N_3478,In_483,In_605);
xnor U3479 (N_3479,In_627,In_324);
or U3480 (N_3480,In_577,In_42);
xnor U3481 (N_3481,In_388,In_789);
and U3482 (N_3482,In_72,In_140);
xnor U3483 (N_3483,In_21,In_859);
nand U3484 (N_3484,In_231,In_166);
nor U3485 (N_3485,In_149,In_360);
nor U3486 (N_3486,In_821,In_615);
or U3487 (N_3487,In_989,In_369);
and U3488 (N_3488,In_242,In_293);
nor U3489 (N_3489,In_875,In_858);
nor U3490 (N_3490,In_46,In_179);
nand U3491 (N_3491,In_618,In_673);
and U3492 (N_3492,In_920,In_947);
or U3493 (N_3493,In_713,In_903);
xor U3494 (N_3494,In_802,In_787);
or U3495 (N_3495,In_676,In_80);
xnor U3496 (N_3496,In_707,In_459);
or U3497 (N_3497,In_228,In_12);
nand U3498 (N_3498,In_127,In_48);
nand U3499 (N_3499,In_764,In_171);
nand U3500 (N_3500,In_117,In_176);
nand U3501 (N_3501,In_530,In_817);
xnor U3502 (N_3502,In_590,In_779);
nand U3503 (N_3503,In_117,In_392);
nor U3504 (N_3504,In_942,In_752);
xor U3505 (N_3505,In_834,In_226);
xor U3506 (N_3506,In_942,In_517);
and U3507 (N_3507,In_824,In_163);
nor U3508 (N_3508,In_810,In_934);
and U3509 (N_3509,In_354,In_19);
or U3510 (N_3510,In_700,In_369);
nand U3511 (N_3511,In_121,In_191);
xnor U3512 (N_3512,In_931,In_267);
or U3513 (N_3513,In_56,In_254);
xor U3514 (N_3514,In_236,In_166);
xnor U3515 (N_3515,In_461,In_301);
nand U3516 (N_3516,In_661,In_915);
nand U3517 (N_3517,In_140,In_607);
nor U3518 (N_3518,In_768,In_150);
and U3519 (N_3519,In_117,In_144);
and U3520 (N_3520,In_979,In_297);
and U3521 (N_3521,In_938,In_803);
and U3522 (N_3522,In_315,In_760);
nand U3523 (N_3523,In_810,In_585);
and U3524 (N_3524,In_537,In_686);
or U3525 (N_3525,In_777,In_753);
nor U3526 (N_3526,In_324,In_689);
nand U3527 (N_3527,In_650,In_114);
and U3528 (N_3528,In_952,In_654);
or U3529 (N_3529,In_462,In_499);
or U3530 (N_3530,In_771,In_909);
nand U3531 (N_3531,In_654,In_679);
nand U3532 (N_3532,In_103,In_221);
or U3533 (N_3533,In_68,In_404);
nor U3534 (N_3534,In_455,In_889);
and U3535 (N_3535,In_449,In_826);
nor U3536 (N_3536,In_632,In_43);
nand U3537 (N_3537,In_721,In_799);
or U3538 (N_3538,In_76,In_678);
or U3539 (N_3539,In_213,In_548);
nand U3540 (N_3540,In_735,In_430);
xnor U3541 (N_3541,In_233,In_612);
nand U3542 (N_3542,In_683,In_504);
nand U3543 (N_3543,In_424,In_504);
or U3544 (N_3544,In_516,In_57);
nand U3545 (N_3545,In_81,In_307);
xnor U3546 (N_3546,In_38,In_759);
nor U3547 (N_3547,In_461,In_267);
and U3548 (N_3548,In_965,In_670);
and U3549 (N_3549,In_568,In_720);
and U3550 (N_3550,In_556,In_808);
or U3551 (N_3551,In_927,In_390);
nor U3552 (N_3552,In_368,In_355);
xor U3553 (N_3553,In_758,In_3);
nand U3554 (N_3554,In_231,In_35);
xnor U3555 (N_3555,In_520,In_427);
and U3556 (N_3556,In_348,In_495);
and U3557 (N_3557,In_208,In_969);
or U3558 (N_3558,In_947,In_66);
xor U3559 (N_3559,In_761,In_411);
nor U3560 (N_3560,In_341,In_610);
xor U3561 (N_3561,In_238,In_834);
nor U3562 (N_3562,In_502,In_675);
or U3563 (N_3563,In_740,In_956);
or U3564 (N_3564,In_610,In_756);
and U3565 (N_3565,In_309,In_626);
nor U3566 (N_3566,In_127,In_59);
or U3567 (N_3567,In_445,In_417);
nand U3568 (N_3568,In_771,In_26);
or U3569 (N_3569,In_615,In_317);
xor U3570 (N_3570,In_995,In_834);
xor U3571 (N_3571,In_539,In_840);
nor U3572 (N_3572,In_64,In_737);
xor U3573 (N_3573,In_146,In_72);
nand U3574 (N_3574,In_95,In_263);
nor U3575 (N_3575,In_151,In_644);
xnor U3576 (N_3576,In_799,In_507);
or U3577 (N_3577,In_820,In_239);
nor U3578 (N_3578,In_550,In_315);
or U3579 (N_3579,In_767,In_520);
xor U3580 (N_3580,In_244,In_594);
and U3581 (N_3581,In_948,In_743);
nand U3582 (N_3582,In_260,In_55);
nor U3583 (N_3583,In_69,In_230);
xnor U3584 (N_3584,In_968,In_427);
and U3585 (N_3585,In_973,In_414);
xnor U3586 (N_3586,In_667,In_210);
or U3587 (N_3587,In_869,In_316);
nor U3588 (N_3588,In_116,In_513);
nor U3589 (N_3589,In_612,In_401);
nor U3590 (N_3590,In_258,In_946);
nor U3591 (N_3591,In_241,In_945);
xnor U3592 (N_3592,In_630,In_980);
and U3593 (N_3593,In_191,In_269);
and U3594 (N_3594,In_832,In_238);
and U3595 (N_3595,In_647,In_105);
or U3596 (N_3596,In_665,In_278);
nand U3597 (N_3597,In_745,In_400);
or U3598 (N_3598,In_124,In_621);
and U3599 (N_3599,In_431,In_257);
nor U3600 (N_3600,In_863,In_550);
or U3601 (N_3601,In_920,In_340);
or U3602 (N_3602,In_975,In_899);
nor U3603 (N_3603,In_948,In_49);
nor U3604 (N_3604,In_355,In_385);
xor U3605 (N_3605,In_623,In_366);
nor U3606 (N_3606,In_569,In_999);
xnor U3607 (N_3607,In_406,In_96);
nand U3608 (N_3608,In_312,In_429);
nor U3609 (N_3609,In_706,In_564);
nand U3610 (N_3610,In_172,In_69);
nor U3611 (N_3611,In_366,In_811);
and U3612 (N_3612,In_468,In_777);
and U3613 (N_3613,In_354,In_560);
or U3614 (N_3614,In_852,In_712);
nand U3615 (N_3615,In_585,In_323);
nor U3616 (N_3616,In_69,In_952);
xor U3617 (N_3617,In_909,In_787);
nor U3618 (N_3618,In_326,In_74);
xnor U3619 (N_3619,In_746,In_989);
nand U3620 (N_3620,In_540,In_619);
nand U3621 (N_3621,In_865,In_177);
nor U3622 (N_3622,In_155,In_329);
nor U3623 (N_3623,In_540,In_582);
nand U3624 (N_3624,In_683,In_941);
or U3625 (N_3625,In_288,In_605);
and U3626 (N_3626,In_629,In_482);
xor U3627 (N_3627,In_751,In_783);
nor U3628 (N_3628,In_126,In_935);
nand U3629 (N_3629,In_591,In_72);
and U3630 (N_3630,In_718,In_487);
or U3631 (N_3631,In_664,In_29);
and U3632 (N_3632,In_953,In_344);
nand U3633 (N_3633,In_270,In_515);
or U3634 (N_3634,In_840,In_580);
or U3635 (N_3635,In_755,In_76);
or U3636 (N_3636,In_747,In_166);
xnor U3637 (N_3637,In_615,In_859);
nor U3638 (N_3638,In_937,In_200);
and U3639 (N_3639,In_329,In_285);
or U3640 (N_3640,In_762,In_822);
nor U3641 (N_3641,In_270,In_529);
and U3642 (N_3642,In_518,In_697);
nor U3643 (N_3643,In_589,In_38);
or U3644 (N_3644,In_98,In_818);
and U3645 (N_3645,In_201,In_214);
xnor U3646 (N_3646,In_244,In_391);
nor U3647 (N_3647,In_143,In_680);
nand U3648 (N_3648,In_64,In_578);
nor U3649 (N_3649,In_197,In_516);
nor U3650 (N_3650,In_961,In_436);
nand U3651 (N_3651,In_56,In_768);
and U3652 (N_3652,In_513,In_474);
or U3653 (N_3653,In_845,In_970);
and U3654 (N_3654,In_555,In_331);
nor U3655 (N_3655,In_648,In_603);
and U3656 (N_3656,In_688,In_490);
nand U3657 (N_3657,In_351,In_549);
xnor U3658 (N_3658,In_530,In_215);
or U3659 (N_3659,In_777,In_134);
and U3660 (N_3660,In_366,In_806);
xor U3661 (N_3661,In_494,In_965);
nand U3662 (N_3662,In_297,In_232);
or U3663 (N_3663,In_845,In_68);
and U3664 (N_3664,In_557,In_50);
nor U3665 (N_3665,In_450,In_488);
or U3666 (N_3666,In_162,In_618);
nand U3667 (N_3667,In_832,In_331);
nand U3668 (N_3668,In_971,In_219);
or U3669 (N_3669,In_643,In_687);
and U3670 (N_3670,In_634,In_894);
nor U3671 (N_3671,In_710,In_727);
nor U3672 (N_3672,In_220,In_883);
or U3673 (N_3673,In_635,In_833);
xnor U3674 (N_3674,In_688,In_288);
and U3675 (N_3675,In_235,In_723);
xor U3676 (N_3676,In_503,In_661);
xnor U3677 (N_3677,In_229,In_194);
xnor U3678 (N_3678,In_511,In_214);
nand U3679 (N_3679,In_630,In_890);
or U3680 (N_3680,In_946,In_373);
xor U3681 (N_3681,In_21,In_928);
and U3682 (N_3682,In_617,In_659);
nor U3683 (N_3683,In_956,In_477);
and U3684 (N_3684,In_899,In_278);
xor U3685 (N_3685,In_744,In_87);
nor U3686 (N_3686,In_771,In_298);
nand U3687 (N_3687,In_762,In_375);
or U3688 (N_3688,In_599,In_191);
and U3689 (N_3689,In_704,In_14);
and U3690 (N_3690,In_955,In_507);
xnor U3691 (N_3691,In_713,In_28);
or U3692 (N_3692,In_901,In_856);
nand U3693 (N_3693,In_255,In_407);
nor U3694 (N_3694,In_346,In_382);
nand U3695 (N_3695,In_518,In_826);
or U3696 (N_3696,In_869,In_960);
nand U3697 (N_3697,In_722,In_782);
nor U3698 (N_3698,In_336,In_153);
or U3699 (N_3699,In_575,In_503);
nor U3700 (N_3700,In_245,In_752);
nor U3701 (N_3701,In_175,In_708);
or U3702 (N_3702,In_608,In_392);
and U3703 (N_3703,In_233,In_670);
and U3704 (N_3704,In_10,In_90);
nand U3705 (N_3705,In_590,In_106);
and U3706 (N_3706,In_572,In_338);
or U3707 (N_3707,In_111,In_305);
xnor U3708 (N_3708,In_171,In_27);
nand U3709 (N_3709,In_132,In_811);
xor U3710 (N_3710,In_578,In_812);
xnor U3711 (N_3711,In_658,In_815);
nor U3712 (N_3712,In_490,In_804);
or U3713 (N_3713,In_128,In_876);
and U3714 (N_3714,In_698,In_551);
or U3715 (N_3715,In_770,In_96);
nand U3716 (N_3716,In_238,In_557);
nand U3717 (N_3717,In_933,In_659);
and U3718 (N_3718,In_756,In_145);
xor U3719 (N_3719,In_29,In_990);
nand U3720 (N_3720,In_100,In_847);
xnor U3721 (N_3721,In_217,In_12);
or U3722 (N_3722,In_628,In_126);
xnor U3723 (N_3723,In_363,In_151);
and U3724 (N_3724,In_530,In_520);
or U3725 (N_3725,In_616,In_755);
or U3726 (N_3726,In_556,In_767);
xor U3727 (N_3727,In_736,In_825);
or U3728 (N_3728,In_693,In_466);
and U3729 (N_3729,In_910,In_81);
or U3730 (N_3730,In_867,In_753);
and U3731 (N_3731,In_71,In_707);
or U3732 (N_3732,In_427,In_973);
and U3733 (N_3733,In_354,In_159);
nor U3734 (N_3734,In_378,In_781);
nand U3735 (N_3735,In_54,In_425);
or U3736 (N_3736,In_482,In_504);
or U3737 (N_3737,In_31,In_462);
nor U3738 (N_3738,In_543,In_249);
or U3739 (N_3739,In_328,In_407);
or U3740 (N_3740,In_712,In_611);
nor U3741 (N_3741,In_527,In_871);
xor U3742 (N_3742,In_572,In_887);
nor U3743 (N_3743,In_830,In_367);
or U3744 (N_3744,In_272,In_975);
or U3745 (N_3745,In_449,In_442);
nor U3746 (N_3746,In_383,In_205);
xor U3747 (N_3747,In_393,In_581);
and U3748 (N_3748,In_987,In_180);
nor U3749 (N_3749,In_216,In_574);
and U3750 (N_3750,In_516,In_765);
and U3751 (N_3751,In_916,In_100);
and U3752 (N_3752,In_409,In_402);
and U3753 (N_3753,In_126,In_136);
and U3754 (N_3754,In_798,In_880);
and U3755 (N_3755,In_418,In_944);
or U3756 (N_3756,In_916,In_587);
and U3757 (N_3757,In_673,In_704);
nand U3758 (N_3758,In_427,In_796);
or U3759 (N_3759,In_488,In_7);
nor U3760 (N_3760,In_66,In_573);
xnor U3761 (N_3761,In_0,In_367);
nor U3762 (N_3762,In_824,In_494);
and U3763 (N_3763,In_576,In_560);
and U3764 (N_3764,In_959,In_422);
and U3765 (N_3765,In_683,In_930);
xor U3766 (N_3766,In_921,In_919);
nor U3767 (N_3767,In_50,In_542);
xor U3768 (N_3768,In_953,In_291);
xor U3769 (N_3769,In_645,In_896);
nor U3770 (N_3770,In_499,In_614);
xnor U3771 (N_3771,In_512,In_20);
and U3772 (N_3772,In_96,In_407);
nor U3773 (N_3773,In_181,In_371);
or U3774 (N_3774,In_325,In_204);
nand U3775 (N_3775,In_513,In_718);
nand U3776 (N_3776,In_337,In_302);
or U3777 (N_3777,In_187,In_380);
and U3778 (N_3778,In_889,In_551);
or U3779 (N_3779,In_221,In_651);
nor U3780 (N_3780,In_671,In_602);
nand U3781 (N_3781,In_575,In_915);
xor U3782 (N_3782,In_646,In_193);
or U3783 (N_3783,In_435,In_907);
or U3784 (N_3784,In_764,In_60);
or U3785 (N_3785,In_214,In_669);
nand U3786 (N_3786,In_556,In_921);
nor U3787 (N_3787,In_706,In_253);
xor U3788 (N_3788,In_14,In_940);
nand U3789 (N_3789,In_510,In_5);
or U3790 (N_3790,In_296,In_603);
and U3791 (N_3791,In_980,In_921);
nor U3792 (N_3792,In_147,In_121);
nor U3793 (N_3793,In_822,In_31);
or U3794 (N_3794,In_557,In_47);
or U3795 (N_3795,In_981,In_87);
nand U3796 (N_3796,In_198,In_310);
nand U3797 (N_3797,In_239,In_810);
nand U3798 (N_3798,In_428,In_45);
and U3799 (N_3799,In_774,In_128);
and U3800 (N_3800,In_779,In_745);
or U3801 (N_3801,In_577,In_766);
or U3802 (N_3802,In_899,In_467);
and U3803 (N_3803,In_177,In_600);
and U3804 (N_3804,In_308,In_542);
nor U3805 (N_3805,In_394,In_295);
and U3806 (N_3806,In_817,In_785);
xnor U3807 (N_3807,In_394,In_476);
nand U3808 (N_3808,In_710,In_560);
or U3809 (N_3809,In_654,In_670);
or U3810 (N_3810,In_728,In_732);
and U3811 (N_3811,In_465,In_866);
or U3812 (N_3812,In_319,In_68);
or U3813 (N_3813,In_863,In_420);
nor U3814 (N_3814,In_385,In_353);
or U3815 (N_3815,In_495,In_40);
and U3816 (N_3816,In_436,In_862);
xnor U3817 (N_3817,In_640,In_13);
nor U3818 (N_3818,In_197,In_572);
and U3819 (N_3819,In_391,In_635);
nand U3820 (N_3820,In_508,In_650);
nor U3821 (N_3821,In_28,In_971);
nor U3822 (N_3822,In_56,In_728);
nand U3823 (N_3823,In_311,In_693);
xnor U3824 (N_3824,In_733,In_213);
and U3825 (N_3825,In_177,In_475);
xor U3826 (N_3826,In_648,In_582);
xnor U3827 (N_3827,In_714,In_90);
nand U3828 (N_3828,In_646,In_502);
or U3829 (N_3829,In_575,In_126);
and U3830 (N_3830,In_447,In_208);
and U3831 (N_3831,In_811,In_570);
nor U3832 (N_3832,In_886,In_692);
nor U3833 (N_3833,In_354,In_178);
nor U3834 (N_3834,In_738,In_379);
xnor U3835 (N_3835,In_258,In_603);
nand U3836 (N_3836,In_790,In_803);
nor U3837 (N_3837,In_833,In_213);
and U3838 (N_3838,In_292,In_278);
xnor U3839 (N_3839,In_20,In_790);
xnor U3840 (N_3840,In_864,In_899);
xor U3841 (N_3841,In_342,In_891);
and U3842 (N_3842,In_670,In_910);
or U3843 (N_3843,In_465,In_114);
nor U3844 (N_3844,In_967,In_100);
and U3845 (N_3845,In_33,In_89);
or U3846 (N_3846,In_878,In_750);
or U3847 (N_3847,In_911,In_351);
and U3848 (N_3848,In_243,In_860);
and U3849 (N_3849,In_181,In_208);
and U3850 (N_3850,In_361,In_703);
or U3851 (N_3851,In_706,In_580);
xor U3852 (N_3852,In_320,In_214);
or U3853 (N_3853,In_599,In_34);
nand U3854 (N_3854,In_846,In_276);
nor U3855 (N_3855,In_601,In_478);
nand U3856 (N_3856,In_697,In_352);
nor U3857 (N_3857,In_646,In_451);
xnor U3858 (N_3858,In_468,In_984);
or U3859 (N_3859,In_820,In_727);
nand U3860 (N_3860,In_397,In_189);
nand U3861 (N_3861,In_501,In_324);
and U3862 (N_3862,In_79,In_314);
and U3863 (N_3863,In_141,In_125);
nor U3864 (N_3864,In_26,In_398);
nand U3865 (N_3865,In_904,In_48);
and U3866 (N_3866,In_107,In_11);
or U3867 (N_3867,In_379,In_338);
xnor U3868 (N_3868,In_8,In_693);
xor U3869 (N_3869,In_619,In_907);
and U3870 (N_3870,In_45,In_79);
and U3871 (N_3871,In_908,In_915);
or U3872 (N_3872,In_486,In_78);
nor U3873 (N_3873,In_518,In_131);
xor U3874 (N_3874,In_98,In_649);
or U3875 (N_3875,In_912,In_652);
and U3876 (N_3876,In_888,In_568);
and U3877 (N_3877,In_611,In_931);
xnor U3878 (N_3878,In_134,In_355);
or U3879 (N_3879,In_103,In_486);
xnor U3880 (N_3880,In_627,In_326);
nor U3881 (N_3881,In_263,In_108);
nor U3882 (N_3882,In_500,In_963);
or U3883 (N_3883,In_615,In_929);
nor U3884 (N_3884,In_715,In_623);
nor U3885 (N_3885,In_201,In_289);
and U3886 (N_3886,In_441,In_731);
nor U3887 (N_3887,In_717,In_448);
xor U3888 (N_3888,In_355,In_724);
or U3889 (N_3889,In_338,In_27);
nand U3890 (N_3890,In_220,In_22);
or U3891 (N_3891,In_813,In_439);
xnor U3892 (N_3892,In_419,In_689);
and U3893 (N_3893,In_869,In_663);
xor U3894 (N_3894,In_668,In_481);
nor U3895 (N_3895,In_967,In_173);
and U3896 (N_3896,In_640,In_514);
or U3897 (N_3897,In_653,In_64);
and U3898 (N_3898,In_510,In_570);
and U3899 (N_3899,In_59,In_216);
nand U3900 (N_3900,In_212,In_71);
and U3901 (N_3901,In_974,In_254);
xor U3902 (N_3902,In_738,In_168);
xnor U3903 (N_3903,In_220,In_798);
nor U3904 (N_3904,In_682,In_394);
or U3905 (N_3905,In_604,In_618);
nand U3906 (N_3906,In_620,In_555);
xnor U3907 (N_3907,In_489,In_800);
nor U3908 (N_3908,In_498,In_909);
nand U3909 (N_3909,In_760,In_292);
nand U3910 (N_3910,In_199,In_908);
or U3911 (N_3911,In_770,In_912);
nand U3912 (N_3912,In_520,In_834);
nand U3913 (N_3913,In_432,In_77);
nand U3914 (N_3914,In_864,In_465);
nor U3915 (N_3915,In_675,In_132);
nand U3916 (N_3916,In_544,In_510);
xor U3917 (N_3917,In_115,In_861);
nand U3918 (N_3918,In_968,In_816);
nor U3919 (N_3919,In_264,In_547);
nand U3920 (N_3920,In_238,In_176);
nor U3921 (N_3921,In_528,In_396);
and U3922 (N_3922,In_922,In_809);
xor U3923 (N_3923,In_703,In_530);
and U3924 (N_3924,In_844,In_146);
xnor U3925 (N_3925,In_168,In_228);
or U3926 (N_3926,In_944,In_449);
or U3927 (N_3927,In_480,In_118);
nand U3928 (N_3928,In_335,In_242);
xnor U3929 (N_3929,In_336,In_812);
nor U3930 (N_3930,In_379,In_584);
nand U3931 (N_3931,In_492,In_55);
xnor U3932 (N_3932,In_433,In_512);
nor U3933 (N_3933,In_909,In_218);
nor U3934 (N_3934,In_304,In_446);
xnor U3935 (N_3935,In_624,In_178);
xor U3936 (N_3936,In_859,In_190);
nand U3937 (N_3937,In_735,In_389);
and U3938 (N_3938,In_638,In_176);
and U3939 (N_3939,In_995,In_743);
xor U3940 (N_3940,In_617,In_507);
and U3941 (N_3941,In_442,In_670);
xnor U3942 (N_3942,In_370,In_335);
or U3943 (N_3943,In_594,In_393);
and U3944 (N_3944,In_154,In_849);
and U3945 (N_3945,In_74,In_510);
and U3946 (N_3946,In_70,In_713);
nand U3947 (N_3947,In_210,In_223);
xor U3948 (N_3948,In_16,In_555);
nor U3949 (N_3949,In_440,In_802);
or U3950 (N_3950,In_645,In_893);
and U3951 (N_3951,In_568,In_548);
nand U3952 (N_3952,In_612,In_533);
nor U3953 (N_3953,In_953,In_3);
nor U3954 (N_3954,In_433,In_683);
nand U3955 (N_3955,In_982,In_239);
or U3956 (N_3956,In_603,In_349);
nor U3957 (N_3957,In_298,In_276);
nor U3958 (N_3958,In_593,In_406);
xnor U3959 (N_3959,In_464,In_102);
nand U3960 (N_3960,In_291,In_237);
and U3961 (N_3961,In_650,In_586);
nor U3962 (N_3962,In_534,In_316);
and U3963 (N_3963,In_166,In_548);
nand U3964 (N_3964,In_160,In_918);
or U3965 (N_3965,In_346,In_24);
or U3966 (N_3966,In_387,In_781);
nor U3967 (N_3967,In_321,In_525);
nand U3968 (N_3968,In_585,In_403);
nor U3969 (N_3969,In_585,In_804);
or U3970 (N_3970,In_884,In_115);
xnor U3971 (N_3971,In_106,In_187);
or U3972 (N_3972,In_627,In_86);
and U3973 (N_3973,In_276,In_380);
nor U3974 (N_3974,In_40,In_50);
nor U3975 (N_3975,In_72,In_45);
or U3976 (N_3976,In_484,In_784);
nand U3977 (N_3977,In_924,In_212);
or U3978 (N_3978,In_276,In_2);
xnor U3979 (N_3979,In_911,In_781);
nand U3980 (N_3980,In_567,In_779);
nor U3981 (N_3981,In_156,In_959);
nor U3982 (N_3982,In_980,In_255);
xor U3983 (N_3983,In_502,In_842);
nor U3984 (N_3984,In_332,In_491);
and U3985 (N_3985,In_583,In_277);
xnor U3986 (N_3986,In_867,In_64);
xnor U3987 (N_3987,In_894,In_511);
or U3988 (N_3988,In_941,In_490);
nand U3989 (N_3989,In_771,In_599);
and U3990 (N_3990,In_880,In_266);
nor U3991 (N_3991,In_94,In_207);
and U3992 (N_3992,In_976,In_96);
xor U3993 (N_3993,In_217,In_622);
nor U3994 (N_3994,In_727,In_75);
nand U3995 (N_3995,In_753,In_597);
nor U3996 (N_3996,In_983,In_254);
or U3997 (N_3997,In_374,In_716);
xor U3998 (N_3998,In_185,In_385);
nand U3999 (N_3999,In_161,In_544);
nor U4000 (N_4000,In_438,In_916);
xor U4001 (N_4001,In_976,In_593);
or U4002 (N_4002,In_48,In_369);
or U4003 (N_4003,In_29,In_435);
or U4004 (N_4004,In_48,In_218);
and U4005 (N_4005,In_643,In_497);
and U4006 (N_4006,In_684,In_393);
or U4007 (N_4007,In_562,In_574);
or U4008 (N_4008,In_790,In_257);
nor U4009 (N_4009,In_33,In_936);
xnor U4010 (N_4010,In_504,In_152);
nor U4011 (N_4011,In_407,In_65);
nor U4012 (N_4012,In_760,In_907);
nand U4013 (N_4013,In_3,In_759);
and U4014 (N_4014,In_436,In_319);
and U4015 (N_4015,In_727,In_239);
and U4016 (N_4016,In_167,In_930);
xor U4017 (N_4017,In_146,In_707);
xor U4018 (N_4018,In_857,In_907);
nor U4019 (N_4019,In_232,In_670);
or U4020 (N_4020,In_476,In_944);
xnor U4021 (N_4021,In_612,In_500);
nand U4022 (N_4022,In_413,In_836);
xor U4023 (N_4023,In_319,In_287);
nor U4024 (N_4024,In_426,In_345);
or U4025 (N_4025,In_676,In_624);
nand U4026 (N_4026,In_865,In_181);
nand U4027 (N_4027,In_179,In_326);
or U4028 (N_4028,In_362,In_308);
xnor U4029 (N_4029,In_660,In_320);
nand U4030 (N_4030,In_664,In_47);
and U4031 (N_4031,In_947,In_655);
nand U4032 (N_4032,In_266,In_301);
nand U4033 (N_4033,In_56,In_749);
nand U4034 (N_4034,In_772,In_783);
xnor U4035 (N_4035,In_180,In_470);
or U4036 (N_4036,In_759,In_288);
and U4037 (N_4037,In_813,In_523);
or U4038 (N_4038,In_132,In_197);
or U4039 (N_4039,In_449,In_37);
and U4040 (N_4040,In_70,In_687);
nor U4041 (N_4041,In_366,In_514);
nand U4042 (N_4042,In_107,In_153);
and U4043 (N_4043,In_309,In_377);
nor U4044 (N_4044,In_618,In_508);
xnor U4045 (N_4045,In_700,In_489);
nor U4046 (N_4046,In_959,In_192);
xor U4047 (N_4047,In_292,In_351);
nand U4048 (N_4048,In_992,In_592);
nor U4049 (N_4049,In_750,In_747);
nor U4050 (N_4050,In_332,In_447);
or U4051 (N_4051,In_830,In_519);
or U4052 (N_4052,In_49,In_282);
or U4053 (N_4053,In_156,In_408);
nor U4054 (N_4054,In_174,In_641);
or U4055 (N_4055,In_37,In_929);
and U4056 (N_4056,In_212,In_326);
nor U4057 (N_4057,In_597,In_290);
nor U4058 (N_4058,In_872,In_774);
nor U4059 (N_4059,In_791,In_347);
xnor U4060 (N_4060,In_436,In_820);
or U4061 (N_4061,In_954,In_769);
nor U4062 (N_4062,In_373,In_682);
xor U4063 (N_4063,In_484,In_333);
xor U4064 (N_4064,In_546,In_264);
xnor U4065 (N_4065,In_506,In_177);
xnor U4066 (N_4066,In_507,In_865);
and U4067 (N_4067,In_254,In_488);
and U4068 (N_4068,In_792,In_129);
nor U4069 (N_4069,In_283,In_75);
or U4070 (N_4070,In_955,In_839);
nor U4071 (N_4071,In_844,In_924);
nand U4072 (N_4072,In_570,In_666);
xnor U4073 (N_4073,In_364,In_674);
or U4074 (N_4074,In_993,In_974);
nor U4075 (N_4075,In_494,In_870);
nand U4076 (N_4076,In_780,In_32);
nor U4077 (N_4077,In_851,In_326);
or U4078 (N_4078,In_411,In_462);
xnor U4079 (N_4079,In_53,In_405);
and U4080 (N_4080,In_921,In_67);
nor U4081 (N_4081,In_598,In_261);
nand U4082 (N_4082,In_180,In_751);
and U4083 (N_4083,In_743,In_897);
nor U4084 (N_4084,In_701,In_869);
nor U4085 (N_4085,In_66,In_619);
nand U4086 (N_4086,In_262,In_425);
and U4087 (N_4087,In_286,In_779);
xor U4088 (N_4088,In_246,In_171);
or U4089 (N_4089,In_665,In_154);
nor U4090 (N_4090,In_591,In_849);
nand U4091 (N_4091,In_426,In_361);
nand U4092 (N_4092,In_908,In_279);
xor U4093 (N_4093,In_609,In_488);
and U4094 (N_4094,In_874,In_891);
nand U4095 (N_4095,In_623,In_582);
xor U4096 (N_4096,In_66,In_895);
and U4097 (N_4097,In_145,In_46);
xnor U4098 (N_4098,In_129,In_268);
or U4099 (N_4099,In_313,In_935);
and U4100 (N_4100,In_220,In_233);
or U4101 (N_4101,In_162,In_966);
and U4102 (N_4102,In_939,In_467);
and U4103 (N_4103,In_671,In_865);
and U4104 (N_4104,In_640,In_133);
nor U4105 (N_4105,In_936,In_417);
or U4106 (N_4106,In_478,In_223);
or U4107 (N_4107,In_905,In_785);
nor U4108 (N_4108,In_513,In_938);
xor U4109 (N_4109,In_245,In_691);
nand U4110 (N_4110,In_893,In_400);
xor U4111 (N_4111,In_935,In_97);
and U4112 (N_4112,In_944,In_113);
or U4113 (N_4113,In_172,In_758);
nand U4114 (N_4114,In_891,In_592);
xor U4115 (N_4115,In_930,In_678);
and U4116 (N_4116,In_789,In_129);
nor U4117 (N_4117,In_564,In_592);
or U4118 (N_4118,In_65,In_102);
xor U4119 (N_4119,In_701,In_487);
nor U4120 (N_4120,In_359,In_803);
xnor U4121 (N_4121,In_943,In_515);
nor U4122 (N_4122,In_447,In_0);
xnor U4123 (N_4123,In_30,In_763);
nand U4124 (N_4124,In_434,In_891);
nand U4125 (N_4125,In_650,In_713);
nand U4126 (N_4126,In_480,In_738);
or U4127 (N_4127,In_42,In_477);
nand U4128 (N_4128,In_645,In_575);
xnor U4129 (N_4129,In_522,In_304);
nand U4130 (N_4130,In_830,In_193);
and U4131 (N_4131,In_9,In_943);
nor U4132 (N_4132,In_800,In_652);
nand U4133 (N_4133,In_794,In_978);
and U4134 (N_4134,In_455,In_372);
xnor U4135 (N_4135,In_44,In_668);
and U4136 (N_4136,In_444,In_170);
xor U4137 (N_4137,In_927,In_648);
and U4138 (N_4138,In_151,In_29);
nor U4139 (N_4139,In_331,In_878);
and U4140 (N_4140,In_39,In_464);
or U4141 (N_4141,In_252,In_690);
xnor U4142 (N_4142,In_533,In_489);
and U4143 (N_4143,In_431,In_472);
or U4144 (N_4144,In_224,In_609);
and U4145 (N_4145,In_308,In_281);
nand U4146 (N_4146,In_986,In_997);
nor U4147 (N_4147,In_746,In_891);
or U4148 (N_4148,In_200,In_662);
nand U4149 (N_4149,In_490,In_113);
xnor U4150 (N_4150,In_375,In_12);
and U4151 (N_4151,In_442,In_883);
or U4152 (N_4152,In_126,In_68);
nor U4153 (N_4153,In_561,In_812);
and U4154 (N_4154,In_973,In_534);
or U4155 (N_4155,In_993,In_221);
or U4156 (N_4156,In_689,In_658);
or U4157 (N_4157,In_479,In_570);
nor U4158 (N_4158,In_317,In_684);
or U4159 (N_4159,In_964,In_185);
and U4160 (N_4160,In_533,In_416);
xor U4161 (N_4161,In_934,In_594);
and U4162 (N_4162,In_417,In_729);
and U4163 (N_4163,In_460,In_204);
xnor U4164 (N_4164,In_853,In_735);
and U4165 (N_4165,In_173,In_330);
and U4166 (N_4166,In_333,In_3);
nand U4167 (N_4167,In_363,In_634);
or U4168 (N_4168,In_86,In_711);
xor U4169 (N_4169,In_888,In_855);
xor U4170 (N_4170,In_497,In_291);
or U4171 (N_4171,In_970,In_498);
xnor U4172 (N_4172,In_103,In_885);
xor U4173 (N_4173,In_319,In_788);
nand U4174 (N_4174,In_666,In_303);
xor U4175 (N_4175,In_603,In_624);
nor U4176 (N_4176,In_508,In_759);
nor U4177 (N_4177,In_62,In_632);
nor U4178 (N_4178,In_127,In_979);
or U4179 (N_4179,In_656,In_359);
or U4180 (N_4180,In_559,In_20);
xnor U4181 (N_4181,In_510,In_711);
xor U4182 (N_4182,In_234,In_813);
and U4183 (N_4183,In_396,In_269);
and U4184 (N_4184,In_493,In_987);
nand U4185 (N_4185,In_327,In_792);
xnor U4186 (N_4186,In_706,In_828);
xor U4187 (N_4187,In_590,In_571);
and U4188 (N_4188,In_565,In_324);
nand U4189 (N_4189,In_520,In_656);
and U4190 (N_4190,In_614,In_111);
xor U4191 (N_4191,In_820,In_532);
xor U4192 (N_4192,In_189,In_810);
or U4193 (N_4193,In_543,In_811);
and U4194 (N_4194,In_837,In_887);
or U4195 (N_4195,In_225,In_54);
nor U4196 (N_4196,In_996,In_931);
nor U4197 (N_4197,In_55,In_629);
nor U4198 (N_4198,In_871,In_474);
nor U4199 (N_4199,In_558,In_941);
nand U4200 (N_4200,In_51,In_19);
nor U4201 (N_4201,In_15,In_297);
or U4202 (N_4202,In_200,In_574);
nor U4203 (N_4203,In_327,In_114);
xor U4204 (N_4204,In_22,In_91);
or U4205 (N_4205,In_473,In_124);
nand U4206 (N_4206,In_216,In_118);
xnor U4207 (N_4207,In_812,In_681);
nor U4208 (N_4208,In_434,In_88);
nand U4209 (N_4209,In_774,In_402);
xor U4210 (N_4210,In_671,In_547);
nor U4211 (N_4211,In_651,In_907);
xor U4212 (N_4212,In_389,In_474);
nor U4213 (N_4213,In_947,In_333);
nand U4214 (N_4214,In_102,In_283);
nand U4215 (N_4215,In_707,In_980);
nor U4216 (N_4216,In_747,In_336);
xnor U4217 (N_4217,In_429,In_118);
nor U4218 (N_4218,In_194,In_835);
nand U4219 (N_4219,In_69,In_743);
and U4220 (N_4220,In_936,In_511);
or U4221 (N_4221,In_180,In_615);
and U4222 (N_4222,In_168,In_928);
nand U4223 (N_4223,In_759,In_325);
and U4224 (N_4224,In_911,In_646);
xnor U4225 (N_4225,In_328,In_79);
or U4226 (N_4226,In_360,In_829);
nor U4227 (N_4227,In_766,In_179);
nor U4228 (N_4228,In_36,In_952);
nand U4229 (N_4229,In_827,In_51);
xnor U4230 (N_4230,In_755,In_189);
and U4231 (N_4231,In_316,In_851);
nor U4232 (N_4232,In_374,In_467);
xor U4233 (N_4233,In_837,In_727);
and U4234 (N_4234,In_489,In_369);
or U4235 (N_4235,In_888,In_350);
or U4236 (N_4236,In_202,In_529);
xor U4237 (N_4237,In_235,In_360);
nor U4238 (N_4238,In_258,In_518);
nand U4239 (N_4239,In_951,In_231);
nand U4240 (N_4240,In_104,In_56);
or U4241 (N_4241,In_500,In_955);
and U4242 (N_4242,In_157,In_418);
nor U4243 (N_4243,In_669,In_440);
xor U4244 (N_4244,In_178,In_468);
or U4245 (N_4245,In_72,In_769);
nor U4246 (N_4246,In_426,In_37);
xor U4247 (N_4247,In_98,In_805);
xnor U4248 (N_4248,In_962,In_879);
nor U4249 (N_4249,In_164,In_538);
xnor U4250 (N_4250,In_656,In_889);
nor U4251 (N_4251,In_540,In_300);
nand U4252 (N_4252,In_592,In_242);
nand U4253 (N_4253,In_879,In_891);
nor U4254 (N_4254,In_495,In_592);
or U4255 (N_4255,In_278,In_397);
nand U4256 (N_4256,In_393,In_881);
nand U4257 (N_4257,In_648,In_961);
nor U4258 (N_4258,In_693,In_175);
or U4259 (N_4259,In_212,In_900);
nand U4260 (N_4260,In_465,In_954);
nor U4261 (N_4261,In_448,In_686);
nand U4262 (N_4262,In_489,In_632);
and U4263 (N_4263,In_914,In_36);
or U4264 (N_4264,In_410,In_414);
nand U4265 (N_4265,In_971,In_750);
nand U4266 (N_4266,In_316,In_230);
nor U4267 (N_4267,In_894,In_728);
nand U4268 (N_4268,In_141,In_684);
and U4269 (N_4269,In_907,In_139);
or U4270 (N_4270,In_441,In_738);
nand U4271 (N_4271,In_602,In_328);
or U4272 (N_4272,In_434,In_935);
nand U4273 (N_4273,In_639,In_260);
or U4274 (N_4274,In_965,In_32);
and U4275 (N_4275,In_111,In_298);
and U4276 (N_4276,In_710,In_464);
nand U4277 (N_4277,In_237,In_893);
xor U4278 (N_4278,In_538,In_883);
and U4279 (N_4279,In_141,In_156);
xor U4280 (N_4280,In_929,In_455);
nor U4281 (N_4281,In_248,In_527);
nor U4282 (N_4282,In_154,In_388);
or U4283 (N_4283,In_322,In_215);
nor U4284 (N_4284,In_806,In_608);
nand U4285 (N_4285,In_690,In_999);
and U4286 (N_4286,In_262,In_761);
and U4287 (N_4287,In_101,In_568);
nor U4288 (N_4288,In_626,In_311);
xor U4289 (N_4289,In_883,In_848);
xnor U4290 (N_4290,In_646,In_698);
or U4291 (N_4291,In_991,In_976);
nand U4292 (N_4292,In_124,In_692);
and U4293 (N_4293,In_222,In_48);
nand U4294 (N_4294,In_887,In_537);
and U4295 (N_4295,In_604,In_472);
xor U4296 (N_4296,In_795,In_271);
nor U4297 (N_4297,In_853,In_832);
or U4298 (N_4298,In_308,In_834);
or U4299 (N_4299,In_782,In_621);
and U4300 (N_4300,In_456,In_67);
nor U4301 (N_4301,In_168,In_137);
xnor U4302 (N_4302,In_975,In_831);
or U4303 (N_4303,In_313,In_570);
or U4304 (N_4304,In_333,In_532);
or U4305 (N_4305,In_315,In_878);
or U4306 (N_4306,In_895,In_442);
nand U4307 (N_4307,In_164,In_836);
or U4308 (N_4308,In_792,In_876);
xnor U4309 (N_4309,In_8,In_411);
nor U4310 (N_4310,In_605,In_743);
or U4311 (N_4311,In_472,In_689);
and U4312 (N_4312,In_558,In_494);
xnor U4313 (N_4313,In_752,In_33);
or U4314 (N_4314,In_417,In_791);
and U4315 (N_4315,In_579,In_262);
nor U4316 (N_4316,In_909,In_288);
nor U4317 (N_4317,In_594,In_812);
nand U4318 (N_4318,In_105,In_938);
nand U4319 (N_4319,In_326,In_98);
nand U4320 (N_4320,In_188,In_961);
xor U4321 (N_4321,In_530,In_747);
nor U4322 (N_4322,In_777,In_8);
or U4323 (N_4323,In_827,In_171);
nor U4324 (N_4324,In_324,In_729);
and U4325 (N_4325,In_822,In_381);
and U4326 (N_4326,In_556,In_177);
and U4327 (N_4327,In_342,In_496);
nand U4328 (N_4328,In_658,In_387);
or U4329 (N_4329,In_674,In_807);
xor U4330 (N_4330,In_237,In_988);
or U4331 (N_4331,In_807,In_418);
nor U4332 (N_4332,In_8,In_597);
xnor U4333 (N_4333,In_47,In_491);
nor U4334 (N_4334,In_449,In_625);
or U4335 (N_4335,In_958,In_219);
and U4336 (N_4336,In_828,In_471);
nor U4337 (N_4337,In_192,In_113);
xnor U4338 (N_4338,In_100,In_270);
nor U4339 (N_4339,In_79,In_330);
and U4340 (N_4340,In_867,In_347);
and U4341 (N_4341,In_838,In_786);
nand U4342 (N_4342,In_371,In_31);
xnor U4343 (N_4343,In_540,In_747);
nor U4344 (N_4344,In_324,In_549);
xnor U4345 (N_4345,In_877,In_101);
xor U4346 (N_4346,In_935,In_463);
nor U4347 (N_4347,In_221,In_929);
xnor U4348 (N_4348,In_391,In_709);
or U4349 (N_4349,In_655,In_125);
nand U4350 (N_4350,In_711,In_480);
or U4351 (N_4351,In_699,In_549);
xnor U4352 (N_4352,In_208,In_400);
or U4353 (N_4353,In_58,In_129);
or U4354 (N_4354,In_516,In_959);
nand U4355 (N_4355,In_297,In_516);
xnor U4356 (N_4356,In_337,In_887);
nor U4357 (N_4357,In_588,In_548);
and U4358 (N_4358,In_8,In_661);
nor U4359 (N_4359,In_717,In_358);
xnor U4360 (N_4360,In_333,In_106);
nor U4361 (N_4361,In_168,In_541);
and U4362 (N_4362,In_636,In_479);
nand U4363 (N_4363,In_523,In_44);
and U4364 (N_4364,In_990,In_602);
or U4365 (N_4365,In_706,In_523);
and U4366 (N_4366,In_651,In_811);
and U4367 (N_4367,In_890,In_0);
nand U4368 (N_4368,In_94,In_479);
xor U4369 (N_4369,In_65,In_448);
nand U4370 (N_4370,In_825,In_99);
nor U4371 (N_4371,In_224,In_518);
nand U4372 (N_4372,In_517,In_966);
and U4373 (N_4373,In_852,In_716);
nand U4374 (N_4374,In_850,In_672);
nor U4375 (N_4375,In_955,In_919);
or U4376 (N_4376,In_497,In_373);
xor U4377 (N_4377,In_110,In_672);
and U4378 (N_4378,In_434,In_139);
xor U4379 (N_4379,In_168,In_63);
nor U4380 (N_4380,In_940,In_10);
or U4381 (N_4381,In_161,In_696);
and U4382 (N_4382,In_374,In_277);
nand U4383 (N_4383,In_863,In_542);
nor U4384 (N_4384,In_233,In_989);
xnor U4385 (N_4385,In_904,In_877);
nor U4386 (N_4386,In_549,In_239);
or U4387 (N_4387,In_484,In_237);
and U4388 (N_4388,In_304,In_444);
xnor U4389 (N_4389,In_871,In_310);
or U4390 (N_4390,In_988,In_688);
or U4391 (N_4391,In_361,In_165);
nand U4392 (N_4392,In_826,In_210);
nand U4393 (N_4393,In_999,In_851);
or U4394 (N_4394,In_321,In_318);
nand U4395 (N_4395,In_495,In_949);
nand U4396 (N_4396,In_738,In_970);
and U4397 (N_4397,In_118,In_170);
and U4398 (N_4398,In_754,In_435);
nand U4399 (N_4399,In_884,In_890);
nand U4400 (N_4400,In_28,In_212);
and U4401 (N_4401,In_926,In_458);
nor U4402 (N_4402,In_988,In_797);
or U4403 (N_4403,In_129,In_105);
xor U4404 (N_4404,In_658,In_286);
or U4405 (N_4405,In_873,In_626);
nand U4406 (N_4406,In_289,In_516);
nand U4407 (N_4407,In_30,In_147);
xnor U4408 (N_4408,In_602,In_646);
xnor U4409 (N_4409,In_446,In_300);
and U4410 (N_4410,In_159,In_543);
or U4411 (N_4411,In_386,In_860);
xnor U4412 (N_4412,In_284,In_326);
nand U4413 (N_4413,In_618,In_708);
or U4414 (N_4414,In_439,In_985);
nand U4415 (N_4415,In_778,In_195);
and U4416 (N_4416,In_130,In_656);
nand U4417 (N_4417,In_814,In_823);
nor U4418 (N_4418,In_787,In_257);
xnor U4419 (N_4419,In_986,In_988);
nor U4420 (N_4420,In_811,In_323);
or U4421 (N_4421,In_858,In_568);
or U4422 (N_4422,In_495,In_202);
or U4423 (N_4423,In_97,In_934);
xnor U4424 (N_4424,In_946,In_721);
xnor U4425 (N_4425,In_497,In_364);
or U4426 (N_4426,In_559,In_139);
or U4427 (N_4427,In_102,In_421);
xor U4428 (N_4428,In_449,In_411);
nand U4429 (N_4429,In_600,In_103);
xnor U4430 (N_4430,In_822,In_363);
or U4431 (N_4431,In_783,In_9);
or U4432 (N_4432,In_74,In_494);
xor U4433 (N_4433,In_483,In_419);
nor U4434 (N_4434,In_649,In_543);
nor U4435 (N_4435,In_164,In_725);
xnor U4436 (N_4436,In_870,In_267);
nor U4437 (N_4437,In_672,In_63);
nand U4438 (N_4438,In_884,In_933);
and U4439 (N_4439,In_728,In_554);
and U4440 (N_4440,In_757,In_497);
nand U4441 (N_4441,In_486,In_62);
and U4442 (N_4442,In_464,In_779);
nand U4443 (N_4443,In_701,In_450);
xnor U4444 (N_4444,In_68,In_966);
nand U4445 (N_4445,In_332,In_719);
nor U4446 (N_4446,In_822,In_891);
nand U4447 (N_4447,In_779,In_855);
or U4448 (N_4448,In_792,In_659);
and U4449 (N_4449,In_649,In_748);
nor U4450 (N_4450,In_552,In_767);
or U4451 (N_4451,In_687,In_157);
nand U4452 (N_4452,In_580,In_318);
nand U4453 (N_4453,In_390,In_694);
nand U4454 (N_4454,In_107,In_631);
and U4455 (N_4455,In_791,In_893);
nand U4456 (N_4456,In_137,In_680);
and U4457 (N_4457,In_175,In_595);
or U4458 (N_4458,In_773,In_354);
nor U4459 (N_4459,In_877,In_942);
and U4460 (N_4460,In_194,In_11);
and U4461 (N_4461,In_378,In_420);
xnor U4462 (N_4462,In_11,In_982);
or U4463 (N_4463,In_619,In_197);
or U4464 (N_4464,In_619,In_84);
or U4465 (N_4465,In_123,In_883);
and U4466 (N_4466,In_114,In_69);
nor U4467 (N_4467,In_6,In_892);
xor U4468 (N_4468,In_410,In_213);
nor U4469 (N_4469,In_212,In_172);
and U4470 (N_4470,In_331,In_55);
nor U4471 (N_4471,In_899,In_143);
xnor U4472 (N_4472,In_658,In_273);
nand U4473 (N_4473,In_776,In_781);
nor U4474 (N_4474,In_891,In_599);
or U4475 (N_4475,In_912,In_95);
and U4476 (N_4476,In_950,In_76);
or U4477 (N_4477,In_412,In_361);
nand U4478 (N_4478,In_203,In_732);
or U4479 (N_4479,In_841,In_815);
nor U4480 (N_4480,In_598,In_70);
and U4481 (N_4481,In_651,In_45);
and U4482 (N_4482,In_905,In_780);
nor U4483 (N_4483,In_213,In_867);
nand U4484 (N_4484,In_674,In_432);
nand U4485 (N_4485,In_760,In_132);
and U4486 (N_4486,In_985,In_880);
or U4487 (N_4487,In_394,In_516);
nand U4488 (N_4488,In_124,In_195);
or U4489 (N_4489,In_239,In_257);
or U4490 (N_4490,In_107,In_545);
xnor U4491 (N_4491,In_766,In_263);
or U4492 (N_4492,In_907,In_420);
or U4493 (N_4493,In_609,In_974);
and U4494 (N_4494,In_948,In_876);
or U4495 (N_4495,In_307,In_753);
nor U4496 (N_4496,In_839,In_927);
xor U4497 (N_4497,In_539,In_351);
nand U4498 (N_4498,In_693,In_168);
nor U4499 (N_4499,In_630,In_770);
nand U4500 (N_4500,In_570,In_51);
nor U4501 (N_4501,In_399,In_895);
nor U4502 (N_4502,In_778,In_644);
nor U4503 (N_4503,In_738,In_367);
or U4504 (N_4504,In_869,In_164);
nor U4505 (N_4505,In_117,In_423);
nand U4506 (N_4506,In_717,In_733);
nor U4507 (N_4507,In_121,In_941);
nand U4508 (N_4508,In_799,In_932);
nand U4509 (N_4509,In_592,In_280);
xor U4510 (N_4510,In_566,In_87);
nor U4511 (N_4511,In_534,In_337);
and U4512 (N_4512,In_267,In_785);
and U4513 (N_4513,In_809,In_649);
nor U4514 (N_4514,In_408,In_207);
and U4515 (N_4515,In_302,In_772);
and U4516 (N_4516,In_228,In_720);
nand U4517 (N_4517,In_125,In_138);
xnor U4518 (N_4518,In_361,In_938);
or U4519 (N_4519,In_943,In_208);
xor U4520 (N_4520,In_877,In_790);
or U4521 (N_4521,In_644,In_922);
nand U4522 (N_4522,In_685,In_699);
xor U4523 (N_4523,In_128,In_46);
and U4524 (N_4524,In_678,In_178);
nor U4525 (N_4525,In_29,In_404);
or U4526 (N_4526,In_761,In_184);
and U4527 (N_4527,In_301,In_484);
or U4528 (N_4528,In_727,In_269);
xnor U4529 (N_4529,In_266,In_440);
and U4530 (N_4530,In_884,In_749);
nor U4531 (N_4531,In_834,In_802);
xnor U4532 (N_4532,In_512,In_554);
and U4533 (N_4533,In_33,In_326);
nor U4534 (N_4534,In_52,In_703);
or U4535 (N_4535,In_329,In_40);
or U4536 (N_4536,In_755,In_104);
and U4537 (N_4537,In_204,In_757);
nor U4538 (N_4538,In_763,In_698);
nor U4539 (N_4539,In_331,In_130);
nor U4540 (N_4540,In_586,In_103);
nand U4541 (N_4541,In_754,In_751);
or U4542 (N_4542,In_695,In_919);
or U4543 (N_4543,In_441,In_162);
nand U4544 (N_4544,In_40,In_516);
nand U4545 (N_4545,In_625,In_725);
and U4546 (N_4546,In_844,In_207);
nor U4547 (N_4547,In_816,In_813);
or U4548 (N_4548,In_600,In_716);
and U4549 (N_4549,In_371,In_216);
nand U4550 (N_4550,In_699,In_169);
or U4551 (N_4551,In_953,In_799);
xnor U4552 (N_4552,In_481,In_387);
and U4553 (N_4553,In_541,In_516);
nand U4554 (N_4554,In_428,In_35);
xor U4555 (N_4555,In_500,In_604);
nor U4556 (N_4556,In_448,In_82);
xnor U4557 (N_4557,In_238,In_228);
nand U4558 (N_4558,In_502,In_947);
or U4559 (N_4559,In_752,In_270);
or U4560 (N_4560,In_103,In_616);
and U4561 (N_4561,In_247,In_455);
nor U4562 (N_4562,In_829,In_56);
or U4563 (N_4563,In_197,In_934);
and U4564 (N_4564,In_409,In_655);
nand U4565 (N_4565,In_525,In_385);
xnor U4566 (N_4566,In_421,In_966);
or U4567 (N_4567,In_57,In_524);
xor U4568 (N_4568,In_420,In_217);
nand U4569 (N_4569,In_102,In_600);
xnor U4570 (N_4570,In_249,In_165);
nor U4571 (N_4571,In_897,In_208);
or U4572 (N_4572,In_80,In_416);
xor U4573 (N_4573,In_470,In_719);
xor U4574 (N_4574,In_353,In_945);
nor U4575 (N_4575,In_760,In_273);
and U4576 (N_4576,In_527,In_891);
or U4577 (N_4577,In_508,In_547);
or U4578 (N_4578,In_907,In_842);
and U4579 (N_4579,In_436,In_484);
nor U4580 (N_4580,In_664,In_927);
or U4581 (N_4581,In_401,In_927);
or U4582 (N_4582,In_811,In_793);
nand U4583 (N_4583,In_53,In_424);
and U4584 (N_4584,In_29,In_982);
nand U4585 (N_4585,In_347,In_655);
nor U4586 (N_4586,In_576,In_487);
or U4587 (N_4587,In_409,In_177);
and U4588 (N_4588,In_537,In_470);
nor U4589 (N_4589,In_334,In_30);
nor U4590 (N_4590,In_552,In_184);
nand U4591 (N_4591,In_280,In_371);
nand U4592 (N_4592,In_295,In_162);
nor U4593 (N_4593,In_905,In_487);
nor U4594 (N_4594,In_840,In_851);
xor U4595 (N_4595,In_140,In_554);
xnor U4596 (N_4596,In_706,In_324);
and U4597 (N_4597,In_532,In_774);
nor U4598 (N_4598,In_445,In_199);
nor U4599 (N_4599,In_581,In_757);
nand U4600 (N_4600,In_176,In_6);
xnor U4601 (N_4601,In_284,In_488);
xnor U4602 (N_4602,In_660,In_802);
nor U4603 (N_4603,In_866,In_166);
or U4604 (N_4604,In_845,In_940);
nor U4605 (N_4605,In_749,In_838);
or U4606 (N_4606,In_789,In_954);
xnor U4607 (N_4607,In_306,In_424);
nand U4608 (N_4608,In_52,In_737);
or U4609 (N_4609,In_494,In_953);
nor U4610 (N_4610,In_555,In_591);
or U4611 (N_4611,In_833,In_975);
nand U4612 (N_4612,In_383,In_210);
nand U4613 (N_4613,In_400,In_326);
or U4614 (N_4614,In_999,In_968);
and U4615 (N_4615,In_408,In_461);
nand U4616 (N_4616,In_3,In_809);
xor U4617 (N_4617,In_422,In_645);
nor U4618 (N_4618,In_97,In_618);
and U4619 (N_4619,In_869,In_700);
xor U4620 (N_4620,In_906,In_650);
xnor U4621 (N_4621,In_598,In_803);
and U4622 (N_4622,In_616,In_908);
or U4623 (N_4623,In_749,In_346);
or U4624 (N_4624,In_7,In_264);
xor U4625 (N_4625,In_361,In_386);
nand U4626 (N_4626,In_220,In_994);
nand U4627 (N_4627,In_518,In_779);
nand U4628 (N_4628,In_386,In_322);
xor U4629 (N_4629,In_765,In_967);
xnor U4630 (N_4630,In_796,In_184);
nor U4631 (N_4631,In_666,In_324);
xor U4632 (N_4632,In_787,In_847);
and U4633 (N_4633,In_733,In_348);
xnor U4634 (N_4634,In_489,In_39);
or U4635 (N_4635,In_393,In_531);
xnor U4636 (N_4636,In_625,In_636);
nand U4637 (N_4637,In_227,In_872);
xnor U4638 (N_4638,In_237,In_677);
xnor U4639 (N_4639,In_422,In_47);
and U4640 (N_4640,In_566,In_544);
or U4641 (N_4641,In_284,In_17);
xnor U4642 (N_4642,In_328,In_249);
and U4643 (N_4643,In_46,In_48);
and U4644 (N_4644,In_154,In_382);
and U4645 (N_4645,In_384,In_909);
and U4646 (N_4646,In_621,In_588);
nor U4647 (N_4647,In_29,In_792);
nand U4648 (N_4648,In_953,In_185);
and U4649 (N_4649,In_359,In_976);
and U4650 (N_4650,In_24,In_75);
nand U4651 (N_4651,In_539,In_188);
and U4652 (N_4652,In_963,In_764);
and U4653 (N_4653,In_520,In_832);
xnor U4654 (N_4654,In_562,In_598);
and U4655 (N_4655,In_735,In_622);
and U4656 (N_4656,In_73,In_620);
or U4657 (N_4657,In_162,In_985);
or U4658 (N_4658,In_327,In_437);
nand U4659 (N_4659,In_996,In_708);
or U4660 (N_4660,In_186,In_534);
or U4661 (N_4661,In_632,In_505);
xnor U4662 (N_4662,In_758,In_343);
nand U4663 (N_4663,In_243,In_834);
nor U4664 (N_4664,In_79,In_309);
xor U4665 (N_4665,In_488,In_104);
xnor U4666 (N_4666,In_352,In_172);
nand U4667 (N_4667,In_198,In_451);
nor U4668 (N_4668,In_806,In_864);
xor U4669 (N_4669,In_506,In_776);
xnor U4670 (N_4670,In_444,In_676);
and U4671 (N_4671,In_790,In_711);
xor U4672 (N_4672,In_599,In_376);
nor U4673 (N_4673,In_57,In_79);
xnor U4674 (N_4674,In_608,In_719);
xor U4675 (N_4675,In_620,In_910);
nand U4676 (N_4676,In_361,In_399);
nand U4677 (N_4677,In_715,In_859);
and U4678 (N_4678,In_369,In_170);
nand U4679 (N_4679,In_319,In_595);
nand U4680 (N_4680,In_829,In_439);
or U4681 (N_4681,In_467,In_945);
nand U4682 (N_4682,In_284,In_577);
nand U4683 (N_4683,In_959,In_916);
or U4684 (N_4684,In_542,In_629);
and U4685 (N_4685,In_70,In_381);
or U4686 (N_4686,In_15,In_138);
or U4687 (N_4687,In_708,In_194);
or U4688 (N_4688,In_527,In_349);
and U4689 (N_4689,In_498,In_40);
xnor U4690 (N_4690,In_98,In_999);
nand U4691 (N_4691,In_447,In_560);
nor U4692 (N_4692,In_588,In_606);
and U4693 (N_4693,In_282,In_225);
and U4694 (N_4694,In_273,In_952);
or U4695 (N_4695,In_547,In_477);
nor U4696 (N_4696,In_626,In_215);
or U4697 (N_4697,In_649,In_875);
xnor U4698 (N_4698,In_444,In_834);
nor U4699 (N_4699,In_667,In_937);
and U4700 (N_4700,In_249,In_942);
nand U4701 (N_4701,In_503,In_410);
xor U4702 (N_4702,In_174,In_18);
and U4703 (N_4703,In_724,In_978);
xnor U4704 (N_4704,In_440,In_504);
and U4705 (N_4705,In_114,In_60);
or U4706 (N_4706,In_317,In_346);
xor U4707 (N_4707,In_505,In_375);
nand U4708 (N_4708,In_600,In_483);
or U4709 (N_4709,In_87,In_660);
nand U4710 (N_4710,In_353,In_886);
nor U4711 (N_4711,In_553,In_558);
nand U4712 (N_4712,In_469,In_581);
or U4713 (N_4713,In_145,In_206);
and U4714 (N_4714,In_674,In_325);
and U4715 (N_4715,In_282,In_189);
xor U4716 (N_4716,In_170,In_594);
nor U4717 (N_4717,In_600,In_15);
and U4718 (N_4718,In_95,In_351);
or U4719 (N_4719,In_487,In_583);
or U4720 (N_4720,In_259,In_363);
xnor U4721 (N_4721,In_902,In_867);
nand U4722 (N_4722,In_102,In_892);
and U4723 (N_4723,In_484,In_868);
or U4724 (N_4724,In_735,In_94);
and U4725 (N_4725,In_624,In_196);
nand U4726 (N_4726,In_14,In_81);
and U4727 (N_4727,In_392,In_772);
xor U4728 (N_4728,In_93,In_448);
xnor U4729 (N_4729,In_860,In_529);
or U4730 (N_4730,In_34,In_507);
nand U4731 (N_4731,In_603,In_450);
nor U4732 (N_4732,In_369,In_347);
nor U4733 (N_4733,In_565,In_723);
or U4734 (N_4734,In_369,In_951);
nor U4735 (N_4735,In_748,In_387);
nor U4736 (N_4736,In_211,In_327);
or U4737 (N_4737,In_822,In_167);
xnor U4738 (N_4738,In_0,In_691);
and U4739 (N_4739,In_441,In_439);
or U4740 (N_4740,In_580,In_227);
nand U4741 (N_4741,In_30,In_174);
nand U4742 (N_4742,In_473,In_743);
nand U4743 (N_4743,In_929,In_691);
and U4744 (N_4744,In_50,In_330);
nor U4745 (N_4745,In_239,In_477);
xnor U4746 (N_4746,In_273,In_139);
nand U4747 (N_4747,In_879,In_675);
xnor U4748 (N_4748,In_652,In_660);
or U4749 (N_4749,In_7,In_346);
nor U4750 (N_4750,In_42,In_500);
and U4751 (N_4751,In_176,In_424);
and U4752 (N_4752,In_967,In_877);
nand U4753 (N_4753,In_230,In_707);
nor U4754 (N_4754,In_946,In_796);
nand U4755 (N_4755,In_238,In_356);
nor U4756 (N_4756,In_613,In_786);
and U4757 (N_4757,In_68,In_414);
or U4758 (N_4758,In_893,In_7);
nand U4759 (N_4759,In_145,In_389);
or U4760 (N_4760,In_934,In_542);
nand U4761 (N_4761,In_942,In_395);
or U4762 (N_4762,In_266,In_587);
xor U4763 (N_4763,In_503,In_310);
nand U4764 (N_4764,In_333,In_400);
nand U4765 (N_4765,In_439,In_39);
and U4766 (N_4766,In_638,In_159);
nor U4767 (N_4767,In_258,In_346);
and U4768 (N_4768,In_156,In_99);
and U4769 (N_4769,In_419,In_870);
nand U4770 (N_4770,In_424,In_536);
nor U4771 (N_4771,In_458,In_449);
nand U4772 (N_4772,In_579,In_961);
and U4773 (N_4773,In_703,In_466);
and U4774 (N_4774,In_208,In_407);
nand U4775 (N_4775,In_712,In_302);
nor U4776 (N_4776,In_807,In_707);
xor U4777 (N_4777,In_740,In_307);
or U4778 (N_4778,In_715,In_472);
nor U4779 (N_4779,In_903,In_752);
xor U4780 (N_4780,In_205,In_16);
or U4781 (N_4781,In_22,In_34);
nor U4782 (N_4782,In_423,In_101);
xor U4783 (N_4783,In_665,In_670);
nor U4784 (N_4784,In_707,In_677);
nand U4785 (N_4785,In_428,In_289);
xor U4786 (N_4786,In_436,In_10);
and U4787 (N_4787,In_296,In_717);
or U4788 (N_4788,In_818,In_543);
nand U4789 (N_4789,In_485,In_417);
xor U4790 (N_4790,In_229,In_769);
nand U4791 (N_4791,In_175,In_303);
nand U4792 (N_4792,In_987,In_51);
and U4793 (N_4793,In_161,In_853);
nor U4794 (N_4794,In_496,In_816);
nor U4795 (N_4795,In_323,In_829);
xnor U4796 (N_4796,In_329,In_727);
and U4797 (N_4797,In_242,In_226);
xnor U4798 (N_4798,In_592,In_956);
xnor U4799 (N_4799,In_427,In_10);
or U4800 (N_4800,In_793,In_31);
or U4801 (N_4801,In_962,In_684);
nand U4802 (N_4802,In_242,In_619);
nor U4803 (N_4803,In_108,In_513);
nand U4804 (N_4804,In_226,In_680);
nand U4805 (N_4805,In_528,In_324);
or U4806 (N_4806,In_218,In_530);
nor U4807 (N_4807,In_202,In_98);
or U4808 (N_4808,In_135,In_161);
and U4809 (N_4809,In_348,In_439);
xnor U4810 (N_4810,In_589,In_810);
or U4811 (N_4811,In_551,In_662);
nand U4812 (N_4812,In_552,In_656);
nor U4813 (N_4813,In_569,In_444);
nand U4814 (N_4814,In_773,In_96);
nand U4815 (N_4815,In_176,In_910);
and U4816 (N_4816,In_31,In_611);
nand U4817 (N_4817,In_924,In_437);
nand U4818 (N_4818,In_231,In_379);
or U4819 (N_4819,In_875,In_79);
and U4820 (N_4820,In_241,In_901);
and U4821 (N_4821,In_750,In_499);
nor U4822 (N_4822,In_663,In_382);
nand U4823 (N_4823,In_781,In_348);
nor U4824 (N_4824,In_653,In_813);
and U4825 (N_4825,In_568,In_383);
and U4826 (N_4826,In_632,In_777);
or U4827 (N_4827,In_322,In_839);
nor U4828 (N_4828,In_851,In_922);
and U4829 (N_4829,In_209,In_567);
xnor U4830 (N_4830,In_835,In_628);
xor U4831 (N_4831,In_48,In_121);
nor U4832 (N_4832,In_50,In_406);
xor U4833 (N_4833,In_635,In_522);
nor U4834 (N_4834,In_998,In_884);
nand U4835 (N_4835,In_591,In_415);
nor U4836 (N_4836,In_924,In_170);
and U4837 (N_4837,In_804,In_986);
nand U4838 (N_4838,In_276,In_444);
nand U4839 (N_4839,In_74,In_476);
xor U4840 (N_4840,In_641,In_842);
nor U4841 (N_4841,In_224,In_564);
xnor U4842 (N_4842,In_246,In_736);
and U4843 (N_4843,In_873,In_161);
xor U4844 (N_4844,In_591,In_84);
nor U4845 (N_4845,In_861,In_604);
nand U4846 (N_4846,In_99,In_298);
nor U4847 (N_4847,In_507,In_568);
and U4848 (N_4848,In_527,In_370);
or U4849 (N_4849,In_983,In_920);
and U4850 (N_4850,In_976,In_26);
or U4851 (N_4851,In_350,In_565);
nor U4852 (N_4852,In_612,In_336);
nor U4853 (N_4853,In_607,In_389);
xor U4854 (N_4854,In_735,In_892);
nand U4855 (N_4855,In_725,In_115);
nor U4856 (N_4856,In_747,In_560);
xnor U4857 (N_4857,In_179,In_210);
nand U4858 (N_4858,In_268,In_63);
xor U4859 (N_4859,In_815,In_943);
and U4860 (N_4860,In_113,In_29);
xnor U4861 (N_4861,In_105,In_286);
xor U4862 (N_4862,In_262,In_846);
or U4863 (N_4863,In_323,In_348);
or U4864 (N_4864,In_135,In_741);
nor U4865 (N_4865,In_636,In_418);
nor U4866 (N_4866,In_700,In_562);
and U4867 (N_4867,In_997,In_930);
and U4868 (N_4868,In_169,In_457);
nand U4869 (N_4869,In_709,In_600);
nand U4870 (N_4870,In_768,In_583);
nand U4871 (N_4871,In_14,In_718);
and U4872 (N_4872,In_584,In_27);
nor U4873 (N_4873,In_956,In_490);
or U4874 (N_4874,In_957,In_716);
nor U4875 (N_4875,In_626,In_825);
nand U4876 (N_4876,In_292,In_274);
or U4877 (N_4877,In_563,In_207);
nand U4878 (N_4878,In_376,In_993);
and U4879 (N_4879,In_716,In_75);
nor U4880 (N_4880,In_706,In_926);
and U4881 (N_4881,In_527,In_971);
xor U4882 (N_4882,In_659,In_355);
xor U4883 (N_4883,In_687,In_214);
nor U4884 (N_4884,In_49,In_726);
and U4885 (N_4885,In_10,In_918);
nand U4886 (N_4886,In_104,In_882);
nand U4887 (N_4887,In_987,In_8);
or U4888 (N_4888,In_656,In_636);
nor U4889 (N_4889,In_947,In_641);
and U4890 (N_4890,In_738,In_660);
nor U4891 (N_4891,In_398,In_250);
or U4892 (N_4892,In_316,In_799);
and U4893 (N_4893,In_501,In_177);
nor U4894 (N_4894,In_115,In_696);
nor U4895 (N_4895,In_693,In_485);
nor U4896 (N_4896,In_176,In_983);
and U4897 (N_4897,In_945,In_259);
nor U4898 (N_4898,In_937,In_866);
nand U4899 (N_4899,In_752,In_754);
nand U4900 (N_4900,In_623,In_404);
nand U4901 (N_4901,In_530,In_108);
nand U4902 (N_4902,In_314,In_993);
nand U4903 (N_4903,In_661,In_721);
xor U4904 (N_4904,In_198,In_710);
or U4905 (N_4905,In_2,In_330);
xor U4906 (N_4906,In_302,In_301);
nor U4907 (N_4907,In_416,In_502);
nor U4908 (N_4908,In_820,In_782);
or U4909 (N_4909,In_780,In_27);
nand U4910 (N_4910,In_621,In_120);
nand U4911 (N_4911,In_509,In_128);
xor U4912 (N_4912,In_228,In_206);
xor U4913 (N_4913,In_7,In_409);
nor U4914 (N_4914,In_596,In_961);
nor U4915 (N_4915,In_878,In_148);
nand U4916 (N_4916,In_769,In_81);
and U4917 (N_4917,In_908,In_811);
nand U4918 (N_4918,In_588,In_190);
nor U4919 (N_4919,In_779,In_230);
nand U4920 (N_4920,In_621,In_134);
nor U4921 (N_4921,In_871,In_593);
nor U4922 (N_4922,In_121,In_541);
nor U4923 (N_4923,In_97,In_769);
or U4924 (N_4924,In_769,In_252);
and U4925 (N_4925,In_897,In_715);
nor U4926 (N_4926,In_566,In_916);
nor U4927 (N_4927,In_44,In_549);
or U4928 (N_4928,In_152,In_295);
xnor U4929 (N_4929,In_237,In_882);
nor U4930 (N_4930,In_271,In_431);
and U4931 (N_4931,In_801,In_975);
nor U4932 (N_4932,In_878,In_695);
and U4933 (N_4933,In_479,In_308);
and U4934 (N_4934,In_340,In_821);
and U4935 (N_4935,In_691,In_753);
or U4936 (N_4936,In_550,In_394);
nand U4937 (N_4937,In_331,In_600);
nand U4938 (N_4938,In_74,In_470);
xor U4939 (N_4939,In_524,In_879);
nand U4940 (N_4940,In_360,In_257);
nand U4941 (N_4941,In_62,In_129);
xor U4942 (N_4942,In_124,In_935);
xor U4943 (N_4943,In_47,In_732);
xnor U4944 (N_4944,In_362,In_497);
or U4945 (N_4945,In_795,In_870);
or U4946 (N_4946,In_9,In_276);
nand U4947 (N_4947,In_746,In_876);
xnor U4948 (N_4948,In_77,In_82);
and U4949 (N_4949,In_511,In_135);
xnor U4950 (N_4950,In_504,In_354);
or U4951 (N_4951,In_663,In_299);
or U4952 (N_4952,In_466,In_549);
and U4953 (N_4953,In_14,In_885);
nor U4954 (N_4954,In_704,In_258);
nand U4955 (N_4955,In_5,In_306);
and U4956 (N_4956,In_371,In_512);
and U4957 (N_4957,In_265,In_527);
or U4958 (N_4958,In_780,In_650);
xnor U4959 (N_4959,In_657,In_709);
or U4960 (N_4960,In_485,In_560);
xor U4961 (N_4961,In_589,In_772);
and U4962 (N_4962,In_812,In_286);
and U4963 (N_4963,In_338,In_737);
nand U4964 (N_4964,In_55,In_417);
and U4965 (N_4965,In_712,In_997);
nand U4966 (N_4966,In_130,In_990);
or U4967 (N_4967,In_609,In_921);
nand U4968 (N_4968,In_245,In_963);
xor U4969 (N_4969,In_56,In_852);
or U4970 (N_4970,In_975,In_944);
nor U4971 (N_4971,In_464,In_261);
and U4972 (N_4972,In_1,In_245);
nor U4973 (N_4973,In_208,In_155);
or U4974 (N_4974,In_926,In_166);
xnor U4975 (N_4975,In_941,In_228);
or U4976 (N_4976,In_970,In_37);
nor U4977 (N_4977,In_805,In_112);
xor U4978 (N_4978,In_337,In_535);
xor U4979 (N_4979,In_823,In_872);
or U4980 (N_4980,In_966,In_501);
and U4981 (N_4981,In_732,In_849);
and U4982 (N_4982,In_731,In_577);
xnor U4983 (N_4983,In_320,In_449);
nand U4984 (N_4984,In_49,In_158);
and U4985 (N_4985,In_457,In_263);
and U4986 (N_4986,In_275,In_522);
nor U4987 (N_4987,In_926,In_347);
nor U4988 (N_4988,In_267,In_394);
or U4989 (N_4989,In_591,In_315);
xor U4990 (N_4990,In_396,In_132);
nor U4991 (N_4991,In_815,In_165);
or U4992 (N_4992,In_292,In_911);
xnor U4993 (N_4993,In_425,In_257);
nand U4994 (N_4994,In_592,In_967);
and U4995 (N_4995,In_234,In_493);
nand U4996 (N_4996,In_661,In_939);
and U4997 (N_4997,In_26,In_896);
xor U4998 (N_4998,In_640,In_151);
xor U4999 (N_4999,In_447,In_968);
and U5000 (N_5000,N_404,N_1306);
xor U5001 (N_5001,N_3634,N_4630);
and U5002 (N_5002,N_1850,N_618);
xnor U5003 (N_5003,N_539,N_2380);
xnor U5004 (N_5004,N_2168,N_2983);
or U5005 (N_5005,N_2172,N_4478);
nor U5006 (N_5006,N_4923,N_4715);
or U5007 (N_5007,N_1980,N_859);
nor U5008 (N_5008,N_4955,N_1780);
and U5009 (N_5009,N_1958,N_2578);
nor U5010 (N_5010,N_2857,N_1370);
nor U5011 (N_5011,N_413,N_24);
and U5012 (N_5012,N_2126,N_4263);
xor U5013 (N_5013,N_4689,N_3066);
or U5014 (N_5014,N_4585,N_2193);
and U5015 (N_5015,N_3992,N_2307);
xor U5016 (N_5016,N_4175,N_2903);
xnor U5017 (N_5017,N_306,N_3905);
xnor U5018 (N_5018,N_4842,N_311);
xnor U5019 (N_5019,N_3844,N_3647);
nor U5020 (N_5020,N_1545,N_683);
or U5021 (N_5021,N_4363,N_3358);
nor U5022 (N_5022,N_2460,N_4623);
nand U5023 (N_5023,N_4265,N_3530);
nor U5024 (N_5024,N_3230,N_4277);
nand U5025 (N_5025,N_361,N_743);
xor U5026 (N_5026,N_2496,N_1792);
or U5027 (N_5027,N_511,N_3696);
or U5028 (N_5028,N_1194,N_3328);
xor U5029 (N_5029,N_1090,N_1726);
nor U5030 (N_5030,N_2033,N_4801);
and U5031 (N_5031,N_3497,N_2544);
and U5032 (N_5032,N_2194,N_2000);
xor U5033 (N_5033,N_3729,N_398);
nand U5034 (N_5034,N_3330,N_1427);
and U5035 (N_5035,N_1063,N_4687);
nand U5036 (N_5036,N_2199,N_386);
or U5037 (N_5037,N_3372,N_2760);
or U5038 (N_5038,N_4077,N_3478);
nand U5039 (N_5039,N_1614,N_2407);
nor U5040 (N_5040,N_2830,N_2090);
or U5041 (N_5041,N_2438,N_3891);
and U5042 (N_5042,N_2395,N_3040);
nor U5043 (N_5043,N_4112,N_4144);
xor U5044 (N_5044,N_610,N_1616);
and U5045 (N_5045,N_1151,N_2015);
nor U5046 (N_5046,N_1952,N_4587);
nand U5047 (N_5047,N_1812,N_1831);
nor U5048 (N_5048,N_3990,N_476);
nor U5049 (N_5049,N_1525,N_2612);
and U5050 (N_5050,N_4578,N_4927);
or U5051 (N_5051,N_796,N_3265);
xnor U5052 (N_5052,N_556,N_3746);
xor U5053 (N_5053,N_4481,N_3979);
nor U5054 (N_5054,N_3940,N_2315);
nor U5055 (N_5055,N_2519,N_4004);
or U5056 (N_5056,N_200,N_2243);
xnor U5057 (N_5057,N_1155,N_1429);
nand U5058 (N_5058,N_3913,N_2252);
and U5059 (N_5059,N_693,N_604);
and U5060 (N_5060,N_4752,N_4371);
nand U5061 (N_5061,N_1786,N_67);
nor U5062 (N_5062,N_347,N_3097);
nor U5063 (N_5063,N_4453,N_4061);
xor U5064 (N_5064,N_1512,N_4659);
nor U5065 (N_5065,N_2351,N_498);
xor U5066 (N_5066,N_1891,N_3752);
xor U5067 (N_5067,N_3459,N_852);
nand U5068 (N_5068,N_3870,N_2258);
nor U5069 (N_5069,N_1297,N_1269);
xnor U5070 (N_5070,N_553,N_1230);
and U5071 (N_5071,N_210,N_4919);
nor U5072 (N_5072,N_3189,N_1499);
or U5073 (N_5073,N_1927,N_2353);
and U5074 (N_5074,N_1048,N_3117);
nand U5075 (N_5075,N_4704,N_1560);
or U5076 (N_5076,N_3254,N_4023);
or U5077 (N_5077,N_472,N_3334);
or U5078 (N_5078,N_794,N_4522);
nand U5079 (N_5079,N_3597,N_238);
nor U5080 (N_5080,N_977,N_3878);
nand U5081 (N_5081,N_3717,N_1332);
nand U5082 (N_5082,N_1642,N_2248);
or U5083 (N_5083,N_401,N_4465);
xor U5084 (N_5084,N_4768,N_1790);
nand U5085 (N_5085,N_862,N_2652);
and U5086 (N_5086,N_2056,N_3383);
xnor U5087 (N_5087,N_2817,N_4504);
nor U5088 (N_5088,N_2308,N_1347);
xnor U5089 (N_5089,N_854,N_2456);
xnor U5090 (N_5090,N_951,N_2229);
nor U5091 (N_5091,N_3939,N_3397);
and U5092 (N_5092,N_3047,N_2616);
and U5093 (N_5093,N_2179,N_1915);
and U5094 (N_5094,N_2222,N_4290);
xnor U5095 (N_5095,N_3734,N_113);
xor U5096 (N_5096,N_509,N_2533);
xor U5097 (N_5097,N_301,N_4967);
xor U5098 (N_5098,N_1083,N_2709);
and U5099 (N_5099,N_307,N_2672);
and U5100 (N_5100,N_3103,N_4408);
or U5101 (N_5101,N_4648,N_1648);
and U5102 (N_5102,N_265,N_3831);
or U5103 (N_5103,N_1121,N_997);
and U5104 (N_5104,N_3392,N_4025);
xor U5105 (N_5105,N_1870,N_450);
xor U5106 (N_5106,N_4428,N_3957);
and U5107 (N_5107,N_237,N_1920);
xor U5108 (N_5108,N_4382,N_798);
nor U5109 (N_5109,N_12,N_4078);
nor U5110 (N_5110,N_4940,N_581);
or U5111 (N_5111,N_2052,N_2543);
or U5112 (N_5112,N_2355,N_276);
and U5113 (N_5113,N_3260,N_1233);
or U5114 (N_5114,N_4951,N_3731);
and U5115 (N_5115,N_146,N_1774);
and U5116 (N_5116,N_3196,N_37);
nor U5117 (N_5117,N_4507,N_4596);
nand U5118 (N_5118,N_3069,N_4232);
and U5119 (N_5119,N_4091,N_2350);
xnor U5120 (N_5120,N_1342,N_3185);
or U5121 (N_5121,N_4270,N_3379);
nand U5122 (N_5122,N_2928,N_78);
and U5123 (N_5123,N_737,N_4423);
xnor U5124 (N_5124,N_1341,N_428);
nor U5125 (N_5125,N_4526,N_2918);
nor U5126 (N_5126,N_272,N_3811);
nand U5127 (N_5127,N_4145,N_2539);
or U5128 (N_5128,N_205,N_2439);
or U5129 (N_5129,N_2484,N_1491);
xor U5130 (N_5130,N_4062,N_1842);
xnor U5131 (N_5131,N_3823,N_1629);
nand U5132 (N_5132,N_4664,N_2964);
nand U5133 (N_5133,N_3853,N_4284);
or U5134 (N_5134,N_954,N_4421);
and U5135 (N_5135,N_4295,N_152);
xor U5136 (N_5136,N_1945,N_2171);
nor U5137 (N_5137,N_1054,N_4093);
nor U5138 (N_5138,N_706,N_584);
nor U5139 (N_5139,N_3516,N_4647);
nand U5140 (N_5140,N_4088,N_1730);
nor U5141 (N_5141,N_679,N_4095);
nand U5142 (N_5142,N_1882,N_3310);
nor U5143 (N_5143,N_461,N_1771);
xor U5144 (N_5144,N_1623,N_4652);
nand U5145 (N_5145,N_2626,N_2869);
xnor U5146 (N_5146,N_362,N_3055);
nor U5147 (N_5147,N_1075,N_1888);
or U5148 (N_5148,N_2664,N_3596);
nand U5149 (N_5149,N_3958,N_625);
nor U5150 (N_5150,N_4656,N_1047);
nand U5151 (N_5151,N_3956,N_1702);
xor U5152 (N_5152,N_2769,N_633);
and U5153 (N_5153,N_3413,N_264);
nand U5154 (N_5154,N_2149,N_3114);
and U5155 (N_5155,N_4928,N_1025);
and U5156 (N_5156,N_4282,N_1459);
nand U5157 (N_5157,N_3449,N_545);
and U5158 (N_5158,N_2134,N_3872);
xor U5159 (N_5159,N_10,N_742);
or U5160 (N_5160,N_491,N_1807);
or U5161 (N_5161,N_920,N_1638);
xnor U5162 (N_5162,N_196,N_363);
nand U5163 (N_5163,N_3214,N_3626);
and U5164 (N_5164,N_3663,N_1365);
nor U5165 (N_5165,N_2992,N_1191);
xnor U5166 (N_5166,N_3266,N_2599);
nand U5167 (N_5167,N_4355,N_2389);
or U5168 (N_5168,N_2982,N_1367);
nor U5169 (N_5169,N_3085,N_534);
nor U5170 (N_5170,N_3165,N_3445);
nand U5171 (N_5171,N_2553,N_4399);
or U5172 (N_5172,N_782,N_4267);
and U5173 (N_5173,N_1637,N_203);
or U5174 (N_5174,N_2795,N_139);
nor U5175 (N_5175,N_1383,N_4356);
or U5176 (N_5176,N_4384,N_3946);
or U5177 (N_5177,N_4931,N_3876);
or U5178 (N_5178,N_3549,N_3246);
and U5179 (N_5179,N_120,N_4783);
nor U5180 (N_5180,N_43,N_4729);
xnor U5181 (N_5181,N_1304,N_3513);
xnor U5182 (N_5182,N_2595,N_436);
nor U5183 (N_5183,N_890,N_4024);
xnor U5184 (N_5184,N_577,N_1716);
xnor U5185 (N_5185,N_3728,N_1506);
nand U5186 (N_5186,N_790,N_3666);
nor U5187 (N_5187,N_1896,N_1044);
nand U5188 (N_5188,N_2705,N_620);
nor U5189 (N_5189,N_3491,N_844);
or U5190 (N_5190,N_3226,N_1772);
and U5191 (N_5191,N_1229,N_2949);
nand U5192 (N_5192,N_4431,N_4863);
and U5193 (N_5193,N_395,N_516);
or U5194 (N_5194,N_151,N_135);
nor U5195 (N_5195,N_3381,N_686);
xnor U5196 (N_5196,N_2494,N_2382);
nor U5197 (N_5197,N_376,N_2192);
nand U5198 (N_5198,N_2343,N_3178);
xnor U5199 (N_5199,N_628,N_142);
xor U5200 (N_5200,N_3465,N_1785);
and U5201 (N_5201,N_2835,N_4926);
or U5202 (N_5202,N_3309,N_4694);
and U5203 (N_5203,N_2984,N_3276);
nor U5204 (N_5204,N_4812,N_3423);
nor U5205 (N_5205,N_1886,N_4747);
and U5206 (N_5206,N_2666,N_2790);
and U5207 (N_5207,N_1813,N_2966);
or U5208 (N_5208,N_1213,N_317);
nand U5209 (N_5209,N_967,N_1169);
and U5210 (N_5210,N_4369,N_247);
and U5211 (N_5211,N_328,N_864);
nand U5212 (N_5212,N_338,N_4543);
nor U5213 (N_5213,N_2403,N_4167);
xor U5214 (N_5214,N_2721,N_3518);
xnor U5215 (N_5215,N_4242,N_636);
or U5216 (N_5216,N_1029,N_290);
and U5217 (N_5217,N_174,N_674);
nor U5218 (N_5218,N_4550,N_2772);
nand U5219 (N_5219,N_144,N_3152);
and U5220 (N_5220,N_297,N_4847);
nand U5221 (N_5221,N_1941,N_2914);
xor U5222 (N_5222,N_1892,N_1251);
nand U5223 (N_5223,N_2281,N_3593);
or U5224 (N_5224,N_3616,N_3754);
or U5225 (N_5225,N_2782,N_3279);
nand U5226 (N_5226,N_2880,N_1996);
nand U5227 (N_5227,N_2723,N_3953);
and U5228 (N_5228,N_3164,N_195);
nand U5229 (N_5229,N_3719,N_849);
nor U5230 (N_5230,N_3959,N_3598);
and U5231 (N_5231,N_3716,N_74);
or U5232 (N_5232,N_1284,N_2681);
xnor U5233 (N_5233,N_3357,N_3702);
xor U5234 (N_5234,N_3573,N_3089);
nand U5235 (N_5235,N_2216,N_4096);
xor U5236 (N_5236,N_54,N_3700);
or U5237 (N_5237,N_1398,N_957);
and U5238 (N_5238,N_2839,N_3830);
and U5239 (N_5239,N_4915,N_3076);
or U5240 (N_5240,N_751,N_3863);
or U5241 (N_5241,N_860,N_2718);
and U5242 (N_5242,N_1405,N_4162);
and U5243 (N_5243,N_1042,N_694);
and U5244 (N_5244,N_3555,N_2700);
nor U5245 (N_5245,N_172,N_1215);
nor U5246 (N_5246,N_3553,N_1744);
or U5247 (N_5247,N_4865,N_3690);
and U5248 (N_5248,N_2923,N_764);
xor U5249 (N_5249,N_3967,N_2);
and U5250 (N_5250,N_788,N_1680);
nor U5251 (N_5251,N_382,N_2017);
xor U5252 (N_5252,N_1404,N_1632);
xnor U5253 (N_5253,N_1684,N_2627);
nor U5254 (N_5254,N_1705,N_3221);
and U5255 (N_5255,N_4047,N_3390);
and U5256 (N_5256,N_3481,N_1281);
or U5257 (N_5257,N_687,N_853);
xor U5258 (N_5258,N_3858,N_2195);
nor U5259 (N_5259,N_2062,N_3348);
nor U5260 (N_5260,N_2853,N_2895);
and U5261 (N_5261,N_3452,N_1561);
or U5262 (N_5262,N_4612,N_3949);
xor U5263 (N_5263,N_2478,N_1337);
nand U5264 (N_5264,N_153,N_115);
nand U5265 (N_5265,N_2094,N_4850);
nand U5266 (N_5266,N_1556,N_4495);
xor U5267 (N_5267,N_2204,N_591);
nor U5268 (N_5268,N_2596,N_3715);
and U5269 (N_5269,N_2971,N_4691);
nor U5270 (N_5270,N_4040,N_1312);
xnor U5271 (N_5271,N_2811,N_3817);
and U5272 (N_5272,N_1816,N_4236);
xnor U5273 (N_5273,N_1052,N_3337);
xnor U5274 (N_5274,N_2943,N_279);
nor U5275 (N_5275,N_2297,N_622);
xnor U5276 (N_5276,N_3936,N_1140);
nor U5277 (N_5277,N_1817,N_2941);
nand U5278 (N_5278,N_2485,N_702);
nor U5279 (N_5279,N_3453,N_1656);
xor U5280 (N_5280,N_938,N_729);
nor U5281 (N_5281,N_564,N_3346);
xor U5282 (N_5282,N_4224,N_3378);
xnor U5283 (N_5283,N_191,N_2648);
xnor U5284 (N_5284,N_2487,N_3400);
nor U5285 (N_5285,N_3336,N_3096);
and U5286 (N_5286,N_2729,N_927);
and U5287 (N_5287,N_2799,N_4828);
xnor U5288 (N_5288,N_1302,N_3755);
nor U5289 (N_5289,N_4539,N_906);
nand U5290 (N_5290,N_598,N_1551);
nor U5291 (N_5291,N_262,N_3180);
nand U5292 (N_5292,N_433,N_4509);
and U5293 (N_5293,N_2255,N_4468);
and U5294 (N_5294,N_3768,N_632);
nand U5295 (N_5295,N_4151,N_1541);
nor U5296 (N_5296,N_3283,N_2261);
nor U5297 (N_5297,N_2574,N_2099);
nor U5298 (N_5298,N_2774,N_1372);
or U5299 (N_5299,N_1620,N_4698);
nand U5300 (N_5300,N_910,N_2414);
and U5301 (N_5301,N_3366,N_4633);
or U5302 (N_5302,N_4721,N_4442);
or U5303 (N_5303,N_4143,N_4100);
nor U5304 (N_5304,N_4855,N_3763);
and U5305 (N_5305,N_3241,N_3082);
or U5306 (N_5306,N_2463,N_4903);
nor U5307 (N_5307,N_242,N_3901);
or U5308 (N_5308,N_1818,N_70);
nor U5309 (N_5309,N_1708,N_903);
nand U5310 (N_5310,N_340,N_64);
and U5311 (N_5311,N_2112,N_2091);
or U5312 (N_5312,N_3539,N_3461);
nor U5313 (N_5313,N_2898,N_358);
nor U5314 (N_5314,N_4517,N_1657);
or U5315 (N_5315,N_1206,N_421);
nand U5316 (N_5316,N_3438,N_2613);
or U5317 (N_5317,N_924,N_2958);
nand U5318 (N_5318,N_356,N_409);
nor U5319 (N_5319,N_992,N_2735);
xnor U5320 (N_5320,N_2997,N_3910);
or U5321 (N_5321,N_4849,N_2232);
or U5322 (N_5322,N_1704,N_1250);
nand U5323 (N_5323,N_93,N_1550);
nand U5324 (N_5324,N_698,N_2571);
and U5325 (N_5325,N_2715,N_2980);
xnor U5326 (N_5326,N_2783,N_4213);
or U5327 (N_5327,N_2634,N_2186);
or U5328 (N_5328,N_89,N_4204);
or U5329 (N_5329,N_1921,N_3933);
or U5330 (N_5330,N_2738,N_394);
and U5331 (N_5331,N_4124,N_865);
nand U5332 (N_5332,N_3506,N_4046);
nand U5333 (N_5333,N_1410,N_2884);
nor U5334 (N_5334,N_4942,N_3380);
and U5335 (N_5335,N_1701,N_4748);
nor U5336 (N_5336,N_4965,N_3159);
or U5337 (N_5337,N_3224,N_4310);
and U5338 (N_5338,N_4693,N_2486);
or U5339 (N_5339,N_2200,N_1674);
nand U5340 (N_5340,N_3407,N_3249);
and U5341 (N_5341,N_1880,N_774);
nor U5342 (N_5342,N_2098,N_3437);
or U5343 (N_5343,N_1755,N_2588);
nor U5344 (N_5344,N_998,N_4475);
nor U5345 (N_5345,N_650,N_4299);
nor U5346 (N_5346,N_2538,N_3988);
or U5347 (N_5347,N_1500,N_3815);
and U5348 (N_5348,N_1388,N_4383);
xor U5349 (N_5349,N_4220,N_3471);
nand U5350 (N_5350,N_3501,N_4339);
xnor U5351 (N_5351,N_2785,N_800);
nor U5352 (N_5352,N_4774,N_712);
nor U5353 (N_5353,N_3802,N_3801);
xnor U5354 (N_5354,N_3744,N_3883);
nor U5355 (N_5355,N_4595,N_425);
nand U5356 (N_5356,N_593,N_4785);
and U5357 (N_5357,N_730,N_3673);
nor U5358 (N_5358,N_2654,N_1908);
nand U5359 (N_5359,N_2967,N_2837);
nor U5360 (N_5360,N_2237,N_204);
xnor U5361 (N_5361,N_2908,N_2051);
nand U5362 (N_5362,N_3977,N_1977);
xnor U5363 (N_5363,N_1677,N_3208);
and U5364 (N_5364,N_3125,N_3730);
nor U5365 (N_5365,N_2739,N_3764);
xnor U5366 (N_5366,N_2922,N_1204);
or U5367 (N_5367,N_911,N_983);
nor U5368 (N_5368,N_3251,N_2111);
xnor U5369 (N_5369,N_3895,N_3790);
xor U5370 (N_5370,N_3295,N_785);
or U5371 (N_5371,N_4780,N_733);
xor U5372 (N_5372,N_4745,N_1455);
nor U5373 (N_5373,N_122,N_2568);
and U5374 (N_5374,N_1411,N_3482);
nand U5375 (N_5375,N_805,N_2130);
or U5376 (N_5376,N_1962,N_1861);
xnor U5377 (N_5377,N_4060,N_1067);
nor U5378 (N_5378,N_4619,N_4896);
and U5379 (N_5379,N_1027,N_4616);
and U5380 (N_5380,N_3948,N_579);
nand U5381 (N_5381,N_1382,N_348);
or U5382 (N_5382,N_937,N_1456);
nor U5383 (N_5383,N_3252,N_4337);
nor U5384 (N_5384,N_2674,N_4920);
nand U5385 (N_5385,N_2174,N_568);
nor U5386 (N_5386,N_2671,N_3410);
xor U5387 (N_5387,N_573,N_2934);
or U5388 (N_5388,N_1999,N_657);
and U5389 (N_5389,N_2066,N_3982);
and U5390 (N_5390,N_4169,N_1722);
nand U5391 (N_5391,N_1476,N_4479);
and U5392 (N_5392,N_3470,N_415);
nand U5393 (N_5393,N_7,N_2313);
xnor U5394 (N_5394,N_1033,N_4982);
and U5395 (N_5395,N_2896,N_4400);
nor U5396 (N_5396,N_4971,N_2239);
nand U5397 (N_5397,N_1147,N_1205);
or U5398 (N_5398,N_918,N_4448);
and U5399 (N_5399,N_2608,N_3842);
nand U5400 (N_5400,N_2931,N_4571);
xor U5401 (N_5401,N_4520,N_3091);
or U5402 (N_5402,N_1254,N_1112);
nor U5403 (N_5403,N_128,N_4076);
nand U5404 (N_5404,N_1686,N_2888);
or U5405 (N_5405,N_2184,N_3919);
and U5406 (N_5406,N_4233,N_876);
xor U5407 (N_5407,N_4196,N_2552);
or U5408 (N_5408,N_4870,N_3025);
xnor U5409 (N_5409,N_2013,N_3727);
xor U5410 (N_5410,N_1466,N_4358);
xor U5411 (N_5411,N_1914,N_2491);
nor U5412 (N_5412,N_2766,N_3443);
and U5413 (N_5413,N_4699,N_2357);
and U5414 (N_5414,N_4191,N_17);
nor U5415 (N_5415,N_669,N_529);
nor U5416 (N_5416,N_4878,N_1403);
nand U5417 (N_5417,N_2527,N_2950);
nand U5418 (N_5418,N_837,N_1397);
xnor U5419 (N_5419,N_2773,N_4872);
or U5420 (N_5420,N_381,N_3139);
or U5421 (N_5421,N_3485,N_4063);
xnor U5422 (N_5422,N_776,N_3638);
and U5423 (N_5423,N_3405,N_935);
or U5424 (N_5424,N_1271,N_2041);
xor U5425 (N_5425,N_2002,N_652);
and U5426 (N_5426,N_119,N_1485);
and U5427 (N_5427,N_3981,N_707);
xor U5428 (N_5428,N_2363,N_4523);
nor U5429 (N_5429,N_4327,N_23);
and U5430 (N_5430,N_4746,N_1146);
xnor U5431 (N_5431,N_2048,N_4795);
and U5432 (N_5432,N_892,N_771);
or U5433 (N_5433,N_3333,N_1673);
nor U5434 (N_5434,N_4493,N_1462);
and U5435 (N_5435,N_228,N_4009);
nand U5436 (N_5436,N_3402,N_3054);
nor U5437 (N_5437,N_3079,N_1399);
xnor U5438 (N_5438,N_391,N_1448);
xnor U5439 (N_5439,N_4483,N_3431);
or U5440 (N_5440,N_4029,N_3050);
nor U5441 (N_5441,N_2336,N_4244);
xor U5442 (N_5442,N_1059,N_2637);
or U5443 (N_5443,N_1401,N_2159);
nor U5444 (N_5444,N_576,N_4451);
and U5445 (N_5445,N_4129,N_4807);
nand U5446 (N_5446,N_2489,N_664);
or U5447 (N_5447,N_3281,N_4621);
or U5448 (N_5448,N_4978,N_3363);
and U5449 (N_5449,N_2140,N_821);
nand U5450 (N_5450,N_4153,N_791);
xor U5451 (N_5451,N_2849,N_1948);
nand U5452 (N_5452,N_4271,N_1292);
nor U5453 (N_5453,N_4788,N_2752);
or U5454 (N_5454,N_4172,N_11);
xor U5455 (N_5455,N_761,N_4203);
nand U5456 (N_5456,N_367,N_840);
xnor U5457 (N_5457,N_1672,N_4357);
xnor U5458 (N_5458,N_1148,N_1574);
nand U5459 (N_5459,N_1103,N_4929);
and U5460 (N_5460,N_4871,N_1473);
and U5461 (N_5461,N_922,N_1081);
nor U5462 (N_5462,N_3899,N_3551);
nor U5463 (N_5463,N_804,N_4713);
or U5464 (N_5464,N_1978,N_299);
and U5465 (N_5465,N_3862,N_1894);
xor U5466 (N_5466,N_692,N_2832);
nor U5467 (N_5467,N_4794,N_4246);
or U5468 (N_5468,N_4097,N_4973);
xnor U5469 (N_5469,N_1264,N_4851);
xor U5470 (N_5470,N_4590,N_1009);
nand U5471 (N_5471,N_3109,N_4617);
and U5472 (N_5472,N_1859,N_1161);
nand U5473 (N_5473,N_2361,N_3170);
nand U5474 (N_5474,N_4341,N_2871);
nand U5475 (N_5475,N_4456,N_2713);
or U5476 (N_5476,N_2046,N_2584);
nand U5477 (N_5477,N_2287,N_4737);
nand U5478 (N_5478,N_169,N_4222);
xnor U5479 (N_5479,N_3502,N_2935);
xor U5480 (N_5480,N_540,N_646);
or U5481 (N_5481,N_240,N_2665);
xnor U5482 (N_5482,N_536,N_201);
nand U5483 (N_5483,N_3664,N_1502);
nand U5484 (N_5484,N_1699,N_3589);
nand U5485 (N_5485,N_2632,N_647);
and U5486 (N_5486,N_4818,N_2082);
nand U5487 (N_5487,N_3387,N_4071);
nor U5488 (N_5488,N_735,N_250);
xor U5489 (N_5489,N_4255,N_1320);
nand U5490 (N_5490,N_101,N_2285);
or U5491 (N_5491,N_2408,N_2989);
nand U5492 (N_5492,N_1323,N_2619);
nor U5493 (N_5493,N_2573,N_2886);
nand U5494 (N_5494,N_359,N_1910);
nand U5495 (N_5495,N_324,N_2702);
or U5496 (N_5496,N_2084,N_407);
nand U5497 (N_5497,N_3195,N_147);
or U5498 (N_5498,N_663,N_230);
nor U5499 (N_5499,N_684,N_1728);
or U5500 (N_5500,N_2188,N_1336);
nand U5501 (N_5501,N_2236,N_480);
nand U5502 (N_5502,N_3784,N_3001);
and U5503 (N_5503,N_4391,N_2712);
nand U5504 (N_5504,N_2183,N_2717);
nand U5505 (N_5505,N_3356,N_4755);
or U5506 (N_5506,N_4909,N_3163);
nand U5507 (N_5507,N_4489,N_1606);
and U5508 (N_5508,N_1643,N_3659);
xor U5509 (N_5509,N_4345,N_1417);
and U5510 (N_5510,N_149,N_2656);
nand U5511 (N_5511,N_3263,N_3197);
nand U5512 (N_5512,N_2165,N_3841);
nor U5513 (N_5513,N_945,N_3242);
nor U5514 (N_5514,N_2579,N_4986);
nor U5515 (N_5515,N_1335,N_2120);
and U5516 (N_5516,N_457,N_3723);
xor U5517 (N_5517,N_1596,N_1706);
nor U5518 (N_5518,N_4485,N_2268);
or U5519 (N_5519,N_489,N_944);
xor U5520 (N_5520,N_1330,N_4054);
or U5521 (N_5521,N_2844,N_2796);
xnor U5522 (N_5522,N_2322,N_4413);
xnor U5523 (N_5523,N_907,N_3329);
nor U5524 (N_5524,N_1055,N_1554);
nand U5525 (N_5525,N_2367,N_2018);
xnor U5526 (N_5526,N_3256,N_4728);
xor U5527 (N_5527,N_1354,N_597);
or U5528 (N_5528,N_1107,N_1428);
nand U5529 (N_5529,N_4065,N_1353);
nor U5530 (N_5530,N_4226,N_4300);
and U5531 (N_5531,N_158,N_3030);
nand U5532 (N_5532,N_2556,N_4174);
xnor U5533 (N_5533,N_1781,N_0);
and U5534 (N_5534,N_4274,N_2375);
nand U5535 (N_5535,N_3519,N_690);
and U5536 (N_5536,N_2187,N_1068);
or U5537 (N_5537,N_1835,N_95);
and U5538 (N_5538,N_2461,N_2387);
xnor U5539 (N_5539,N_1765,N_3115);
nor U5540 (N_5540,N_4505,N_3800);
or U5541 (N_5541,N_1150,N_308);
and U5542 (N_5542,N_1858,N_8);
xor U5543 (N_5543,N_1022,N_1235);
and U5544 (N_5544,N_4666,N_1950);
and U5545 (N_5545,N_1767,N_2865);
nand U5546 (N_5546,N_475,N_423);
or U5547 (N_5547,N_2549,N_2330);
nor U5548 (N_5548,N_4135,N_1217);
nand U5549 (N_5549,N_2025,N_827);
or U5550 (N_5550,N_127,N_4538);
and U5551 (N_5551,N_448,N_4389);
nand U5552 (N_5552,N_1819,N_1294);
xor U5553 (N_5553,N_2970,N_3099);
or U5554 (N_5554,N_2876,N_2761);
xnor U5555 (N_5555,N_184,N_2532);
or U5556 (N_5556,N_4702,N_3860);
xor U5557 (N_5557,N_2981,N_2282);
nor U5558 (N_5558,N_1414,N_4503);
and U5559 (N_5559,N_365,N_4880);
or U5560 (N_5560,N_3247,N_3672);
xnor U5561 (N_5561,N_81,N_1757);
nor U5562 (N_5562,N_2039,N_700);
and U5563 (N_5563,N_3104,N_4979);
nand U5564 (N_5564,N_2913,N_4217);
or U5565 (N_5565,N_1588,N_4525);
xnor U5566 (N_5566,N_2021,N_4375);
and U5567 (N_5567,N_2581,N_3012);
xnor U5568 (N_5568,N_1753,N_2128);
and U5569 (N_5569,N_384,N_3877);
and U5570 (N_5570,N_3218,N_4886);
xor U5571 (N_5571,N_3315,N_4335);
xnor U5572 (N_5572,N_1939,N_2698);
or U5573 (N_5573,N_1795,N_2298);
xor U5574 (N_5574,N_1998,N_20);
and U5575 (N_5575,N_1308,N_3859);
or U5576 (N_5576,N_4042,N_3918);
or U5577 (N_5577,N_1532,N_2905);
nor U5578 (N_5578,N_244,N_33);
xor U5579 (N_5579,N_4639,N_1985);
and U5580 (N_5580,N_1837,N_1547);
or U5581 (N_5581,N_4320,N_1801);
or U5582 (N_5582,N_1208,N_949);
xor U5583 (N_5583,N_4305,N_2262);
xor U5584 (N_5584,N_2242,N_2932);
nor U5585 (N_5585,N_1814,N_1319);
xnor U5586 (N_5586,N_1970,N_3278);
and U5587 (N_5587,N_3167,N_812);
nor U5588 (N_5588,N_283,N_2863);
and U5589 (N_5589,N_3866,N_3439);
nor U5590 (N_5590,N_3962,N_4147);
nand U5591 (N_5591,N_2119,N_2814);
and U5592 (N_5592,N_1625,N_3289);
xor U5593 (N_5593,N_1695,N_3533);
nor U5594 (N_5594,N_77,N_4614);
xor U5595 (N_5595,N_3492,N_4642);
xor U5596 (N_5596,N_4336,N_956);
nor U5597 (N_5597,N_835,N_166);
nand U5598 (N_5598,N_4048,N_3833);
or U5599 (N_5599,N_4466,N_4458);
xor U5600 (N_5600,N_756,N_769);
xnor U5601 (N_5601,N_1222,N_1587);
or U5602 (N_5602,N_4532,N_1460);
nand U5603 (N_5603,N_1483,N_4582);
or U5604 (N_5604,N_3839,N_3614);
nor U5605 (N_5605,N_575,N_1199);
nor U5606 (N_5606,N_1543,N_1768);
and U5607 (N_5607,N_3521,N_4852);
nand U5608 (N_5608,N_1128,N_4223);
or U5609 (N_5609,N_2479,N_270);
xnor U5610 (N_5610,N_1855,N_1438);
and U5611 (N_5611,N_3846,N_2009);
and U5612 (N_5612,N_2337,N_1393);
or U5613 (N_5613,N_3585,N_2708);
or U5614 (N_5614,N_3743,N_1391);
xnor U5615 (N_5615,N_2816,N_1508);
and U5616 (N_5616,N_92,N_548);
nand U5617 (N_5617,N_132,N_3709);
or U5618 (N_5618,N_1988,N_2741);
and U5619 (N_5619,N_4997,N_4548);
and U5620 (N_5620,N_1899,N_2939);
xnor U5621 (N_5621,N_4899,N_4700);
and U5622 (N_5622,N_3023,N_2955);
or U5623 (N_5623,N_4820,N_2314);
nand U5624 (N_5624,N_3134,N_4956);
nor U5625 (N_5625,N_4117,N_1902);
nor U5626 (N_5626,N_1869,N_2645);
or U5627 (N_5627,N_755,N_2900);
xnor U5628 (N_5628,N_4106,N_3075);
and U5629 (N_5629,N_4195,N_4516);
nor U5630 (N_5630,N_3753,N_298);
xnor U5631 (N_5631,N_1360,N_1469);
or U5632 (N_5632,N_4118,N_4449);
and U5633 (N_5633,N_2275,N_1177);
xnor U5634 (N_5634,N_3951,N_1533);
and U5635 (N_5635,N_1349,N_2824);
and U5636 (N_5636,N_3433,N_3684);
xnor U5637 (N_5637,N_1856,N_710);
nor U5638 (N_5638,N_3147,N_993);
xnor U5639 (N_5639,N_2798,N_1474);
and U5640 (N_5640,N_3885,N_3712);
nor U5641 (N_5641,N_3984,N_2466);
nor U5642 (N_5642,N_2373,N_3311);
nand U5643 (N_5643,N_1515,N_4922);
xor U5644 (N_5644,N_2758,N_1723);
and U5645 (N_5645,N_2661,N_437);
and U5646 (N_5646,N_2077,N_3536);
xor U5647 (N_5647,N_1446,N_3261);
nand U5648 (N_5648,N_1756,N_2088);
xnor U5649 (N_5649,N_3880,N_341);
or U5650 (N_5650,N_4989,N_970);
or U5651 (N_5651,N_3124,N_4146);
nand U5652 (N_5652,N_2951,N_1020);
or U5653 (N_5653,N_2166,N_2362);
nand U5654 (N_5654,N_1513,N_344);
or U5655 (N_5655,N_985,N_3287);
nand U5656 (N_5656,N_4467,N_3917);
nor U5657 (N_5657,N_4398,N_4089);
and U5658 (N_5658,N_866,N_2050);
or U5659 (N_5659,N_818,N_253);
and U5660 (N_5660,N_4716,N_1839);
and U5661 (N_5661,N_4188,N_2873);
nor U5662 (N_5662,N_4501,N_1418);
and U5663 (N_5663,N_4212,N_4317);
nor U5664 (N_5664,N_3004,N_3600);
nor U5665 (N_5665,N_2415,N_3016);
xor U5666 (N_5666,N_1080,N_1881);
or U5667 (N_5667,N_1170,N_65);
xor U5668 (N_5668,N_1558,N_524);
or U5669 (N_5669,N_2711,N_4193);
and U5670 (N_5670,N_1761,N_3697);
nor U5671 (N_5671,N_3789,N_2043);
or U5672 (N_5672,N_483,N_2245);
nand U5673 (N_5673,N_520,N_1750);
xor U5674 (N_5674,N_767,N_4658);
and U5675 (N_5675,N_1218,N_3554);
and U5676 (N_5676,N_1071,N_3794);
nand U5677 (N_5677,N_1933,N_2818);
and U5678 (N_5678,N_3365,N_2442);
nor U5679 (N_5679,N_3851,N_2004);
or U5680 (N_5680,N_3546,N_4786);
nor U5681 (N_5681,N_2081,N_4683);
xnor U5682 (N_5682,N_2153,N_3002);
nor U5683 (N_5683,N_190,N_4627);
nor U5684 (N_5684,N_4286,N_4808);
and U5685 (N_5685,N_624,N_3654);
xnor U5686 (N_5686,N_2576,N_1764);
nor U5687 (N_5687,N_2152,N_3179);
nor U5688 (N_5688,N_3624,N_4083);
nand U5689 (N_5689,N_3774,N_1694);
or U5690 (N_5690,N_1598,N_3522);
nand U5691 (N_5691,N_4977,N_4092);
nand U5692 (N_5692,N_1621,N_4309);
or U5693 (N_5693,N_170,N_3113);
and U5694 (N_5694,N_2190,N_474);
nor U5695 (N_5695,N_3509,N_3474);
or U5696 (N_5696,N_3759,N_1890);
nor U5697 (N_5697,N_4278,N_1030);
xnor U5698 (N_5698,N_3897,N_3270);
nor U5699 (N_5699,N_2942,N_2291);
nor U5700 (N_5700,N_59,N_3169);
nor U5701 (N_5701,N_4816,N_2856);
or U5702 (N_5702,N_2724,N_2477);
and U5703 (N_5703,N_2504,N_102);
and U5704 (N_5704,N_1564,N_4645);
xnor U5705 (N_5705,N_4497,N_266);
or U5706 (N_5706,N_1176,N_259);
or U5707 (N_5707,N_4688,N_4376);
or U5708 (N_5708,N_1573,N_916);
nor U5709 (N_5709,N_930,N_1135);
or U5710 (N_5710,N_1452,N_4695);
nand U5711 (N_5711,N_4321,N_4730);
nor U5712 (N_5712,N_3520,N_4273);
and U5713 (N_5713,N_287,N_874);
or U5714 (N_5714,N_3112,N_1073);
xor U5715 (N_5715,N_4447,N_3486);
nor U5716 (N_5716,N_1493,N_3401);
xnor U5717 (N_5717,N_4665,N_902);
or U5718 (N_5718,N_1865,N_2516);
nand U5719 (N_5719,N_3623,N_1143);
nor U5720 (N_5720,N_1965,N_1782);
or U5721 (N_5721,N_49,N_2118);
xnor U5722 (N_5722,N_2215,N_4727);
xnor U5723 (N_5723,N_2335,N_1182);
nor U5724 (N_5724,N_2224,N_4996);
or U5725 (N_5725,N_4459,N_3943);
nand U5726 (N_5726,N_3106,N_611);
xnor U5727 (N_5727,N_2850,N_1791);
and U5728 (N_5728,N_1955,N_3203);
nor U5729 (N_5729,N_4120,N_4308);
nor U5730 (N_5730,N_3564,N_53);
and U5731 (N_5731,N_3489,N_3909);
nor U5732 (N_5732,N_4090,N_1386);
nor U5733 (N_5733,N_3010,N_2745);
xor U5734 (N_5734,N_4953,N_3008);
and U5735 (N_5735,N_326,N_3704);
nand U5736 (N_5736,N_1557,N_2176);
or U5737 (N_5737,N_4393,N_410);
nor U5738 (N_5738,N_1118,N_4844);
nand U5739 (N_5739,N_3020,N_1671);
and U5740 (N_5740,N_1285,N_609);
and U5741 (N_5741,N_2392,N_1334);
nor U5742 (N_5742,N_2093,N_3175);
xor U5743 (N_5743,N_339,N_608);
nor U5744 (N_5744,N_1461,N_4790);
nand U5745 (N_5745,N_3669,N_3151);
nor U5746 (N_5746,N_2907,N_1944);
and U5747 (N_5747,N_2945,N_4856);
and U5748 (N_5748,N_4676,N_807);
and U5749 (N_5749,N_1195,N_1225);
and U5750 (N_5750,N_3168,N_4600);
or U5751 (N_5751,N_1576,N_4013);
nor U5752 (N_5752,N_1087,N_1242);
nand U5753 (N_5753,N_3932,N_4625);
xnor U5754 (N_5754,N_2601,N_1871);
or U5755 (N_5755,N_3136,N_3326);
and U5756 (N_5756,N_3291,N_2116);
xnor U5757 (N_5757,N_1644,N_345);
or U5758 (N_5758,N_4370,N_2059);
nor U5759 (N_5759,N_3976,N_4551);
nand U5760 (N_5760,N_2106,N_1082);
and U5761 (N_5761,N_4628,N_858);
or U5762 (N_5762,N_1331,N_2154);
nand U5763 (N_5763,N_2288,N_3524);
nor U5764 (N_5764,N_3619,N_1937);
and U5765 (N_5765,N_211,N_3240);
nor U5766 (N_5766,N_2728,N_2586);
or U5767 (N_5767,N_3544,N_2299);
nand U5768 (N_5768,N_1198,N_950);
xor U5769 (N_5769,N_987,N_2957);
nor U5770 (N_5770,N_3633,N_3761);
nand U5771 (N_5771,N_225,N_2756);
and U5772 (N_5772,N_3590,N_3393);
or U5773 (N_5773,N_3757,N_1338);
or U5774 (N_5774,N_1187,N_4779);
nor U5775 (N_5775,N_1188,N_4266);
nand U5776 (N_5776,N_4420,N_1355);
or U5777 (N_5777,N_1203,N_440);
and U5778 (N_5778,N_3559,N_453);
or U5779 (N_5779,N_3925,N_4677);
or U5780 (N_5780,N_1392,N_62);
xor U5781 (N_5781,N_600,N_2220);
or U5782 (N_5782,N_209,N_1321);
nor U5783 (N_5783,N_4480,N_3297);
and U5784 (N_5784,N_22,N_2334);
nor U5785 (N_5785,N_4432,N_4427);
or U5786 (N_5786,N_3828,N_3223);
xnor U5787 (N_5787,N_2289,N_2383);
nor U5788 (N_5788,N_588,N_678);
nand U5789 (N_5789,N_519,N_2457);
and U5790 (N_5790,N_2686,N_1803);
nand U5791 (N_5791,N_2937,N_4958);
xnor U5792 (N_5792,N_2620,N_1906);
or U5793 (N_5793,N_2095,N_4834);
xor U5794 (N_5794,N_1883,N_2842);
or U5795 (N_5795,N_3837,N_2131);
nor U5796 (N_5796,N_4570,N_537);
nor U5797 (N_5797,N_708,N_1976);
and U5798 (N_5798,N_1599,N_3300);
and U5799 (N_5799,N_526,N_3662);
xor U5800 (N_5800,N_2606,N_2536);
and U5801 (N_5801,N_831,N_731);
and U5802 (N_5802,N_594,N_2453);
xnor U5803 (N_5803,N_4331,N_3698);
and U5804 (N_5804,N_4670,N_3692);
and U5805 (N_5805,N_3205,N_2845);
or U5806 (N_5806,N_3907,N_2240);
nor U5807 (N_5807,N_312,N_1719);
nor U5808 (N_5808,N_1211,N_4074);
xor U5809 (N_5809,N_4564,N_2506);
nor U5810 (N_5810,N_4874,N_4515);
or U5811 (N_5811,N_3921,N_2294);
or U5812 (N_5812,N_4036,N_757);
or U5813 (N_5813,N_4739,N_248);
or U5814 (N_5814,N_1441,N_3377);
or U5815 (N_5815,N_3345,N_235);
nand U5816 (N_5816,N_3578,N_1484);
nand U5817 (N_5817,N_2379,N_227);
or U5818 (N_5818,N_4961,N_1024);
nor U5819 (N_5819,N_4051,N_1692);
nand U5820 (N_5820,N_4803,N_4771);
nand U5821 (N_5821,N_1162,N_335);
xor U5822 (N_5822,N_3072,N_1925);
xnor U5823 (N_5823,N_4474,N_4875);
xnor U5824 (N_5824,N_3711,N_2467);
or U5825 (N_5825,N_3780,N_1986);
and U5826 (N_5826,N_346,N_4791);
and U5827 (N_5827,N_2820,N_561);
and U5828 (N_5828,N_778,N_1581);
nand U5829 (N_5829,N_4668,N_2029);
nand U5830 (N_5830,N_2743,N_1811);
and U5831 (N_5831,N_2454,N_672);
and U5832 (N_5832,N_197,N_4165);
xnor U5833 (N_5833,N_1065,N_4976);
and U5834 (N_5834,N_4749,N_2247);
xor U5835 (N_5835,N_2906,N_251);
or U5836 (N_5836,N_3024,N_383);
and U5837 (N_5837,N_3887,N_2765);
xor U5838 (N_5838,N_1734,N_1276);
or U5839 (N_5839,N_4778,N_670);
xnor U5840 (N_5840,N_982,N_4889);
nor U5841 (N_5841,N_1174,N_84);
nand U5842 (N_5842,N_4650,N_467);
or U5843 (N_5843,N_3523,N_3319);
nor U5844 (N_5844,N_3088,N_2019);
and U5845 (N_5845,N_867,N_4643);
or U5846 (N_5846,N_4939,N_470);
xor U5847 (N_5847,N_403,N_1380);
or U5848 (N_5848,N_114,N_720);
and U5849 (N_5849,N_2902,N_3605);
and U5850 (N_5850,N_284,N_3972);
or U5851 (N_5851,N_1139,N_4450);
xor U5852 (N_5852,N_366,N_2501);
nand U5853 (N_5853,N_773,N_3678);
xor U5854 (N_5854,N_3615,N_4759);
and U5855 (N_5855,N_1193,N_2764);
nor U5856 (N_5856,N_4114,N_4910);
and U5857 (N_5857,N_4669,N_4140);
nand U5858 (N_5858,N_4898,N_2707);
nand U5859 (N_5859,N_1742,N_3508);
or U5860 (N_5860,N_789,N_3991);
nand U5861 (N_5861,N_3118,N_294);
xor U5862 (N_5862,N_4777,N_3576);
or U5863 (N_5863,N_878,N_1345);
nand U5864 (N_5864,N_2846,N_4527);
nand U5865 (N_5865,N_4726,N_1773);
xnor U5866 (N_5866,N_2493,N_4839);
or U5867 (N_5867,N_79,N_3586);
or U5868 (N_5868,N_468,N_1729);
or U5869 (N_5869,N_4935,N_621);
and U5870 (N_5870,N_3144,N_850);
xor U5871 (N_5871,N_1829,N_4050);
or U5872 (N_5872,N_3234,N_4058);
nor U5873 (N_5873,N_4123,N_3639);
nand U5874 (N_5874,N_4241,N_2685);
or U5875 (N_5875,N_2978,N_964);
xor U5876 (N_5876,N_4086,N_171);
or U5877 (N_5877,N_4708,N_676);
xnor U5878 (N_5878,N_4680,N_14);
or U5879 (N_5879,N_3107,N_3849);
or U5880 (N_5880,N_2593,N_1521);
or U5881 (N_5881,N_435,N_1580);
or U5882 (N_5882,N_419,N_3090);
nand U5883 (N_5883,N_1327,N_3490);
xnor U5884 (N_5884,N_1307,N_108);
xnor U5885 (N_5885,N_4422,N_557);
nand U5886 (N_5886,N_1400,N_3320);
nor U5887 (N_5887,N_2901,N_4772);
nand U5888 (N_5888,N_39,N_165);
nand U5889 (N_5889,N_1932,N_4164);
xnor U5890 (N_5890,N_1357,N_68);
xor U5891 (N_5891,N_1972,N_952);
or U5892 (N_5892,N_3994,N_4049);
nor U5893 (N_5893,N_538,N_380);
nand U5894 (N_5894,N_1536,N_2864);
or U5895 (N_5895,N_3884,N_3235);
nand U5896 (N_5896,N_2663,N_2668);
nand U5897 (N_5897,N_1069,N_1612);
nor U5898 (N_5898,N_4462,N_2450);
or U5899 (N_5899,N_2569,N_2792);
nand U5900 (N_5900,N_643,N_4646);
or U5901 (N_5901,N_3355,N_1175);
nor U5902 (N_5902,N_217,N_4269);
nand U5903 (N_5903,N_1465,N_1209);
nor U5904 (N_5904,N_1096,N_4276);
xor U5905 (N_5905,N_656,N_377);
nand U5906 (N_5906,N_4249,N_231);
or U5907 (N_5907,N_959,N_4814);
nor U5908 (N_5908,N_2378,N_3132);
and U5909 (N_5909,N_3537,N_898);
nor U5910 (N_5910,N_249,N_112);
xnor U5911 (N_5911,N_4436,N_869);
nor U5912 (N_5912,N_502,N_1434);
nand U5913 (N_5913,N_905,N_3855);
nor U5914 (N_5914,N_3670,N_2722);
and U5915 (N_5915,N_278,N_3928);
xor U5916 (N_5916,N_291,N_1093);
xor U5917 (N_5917,N_3645,N_966);
nor U5918 (N_5918,N_3468,N_1072);
or U5919 (N_5919,N_2803,N_1261);
and U5920 (N_5920,N_3561,N_2329);
or U5921 (N_5921,N_357,N_1237);
nand U5922 (N_5922,N_1210,N_989);
nand U5923 (N_5923,N_1124,N_3649);
xor U5924 (N_5924,N_4662,N_2411);
or U5925 (N_5925,N_3538,N_329);
and U5926 (N_5926,N_216,N_1415);
and U5927 (N_5927,N_4268,N_1339);
nor U5928 (N_5928,N_4081,N_50);
or U5929 (N_5929,N_2727,N_2144);
and U5930 (N_5930,N_3488,N_770);
nor U5931 (N_5931,N_4945,N_1732);
xor U5932 (N_5932,N_4288,N_2049);
nand U5933 (N_5933,N_1990,N_4157);
or U5934 (N_5934,N_4001,N_1116);
or U5935 (N_5935,N_3915,N_1102);
xnor U5936 (N_5936,N_1433,N_4201);
nand U5937 (N_5937,N_2182,N_3171);
or U5938 (N_5938,N_2067,N_1464);
xor U5939 (N_5939,N_550,N_559);
xor U5940 (N_5940,N_3603,N_1662);
or U5941 (N_5941,N_2936,N_517);
nor U5942 (N_5942,N_2812,N_2296);
xnor U5943 (N_5943,N_506,N_3382);
nand U5944 (N_5944,N_1325,N_1769);
xnor U5945 (N_5945,N_1717,N_3324);
xnor U5946 (N_5946,N_2113,N_2339);
nand U5947 (N_5947,N_104,N_4180);
xnor U5948 (N_5948,N_2063,N_4230);
or U5949 (N_5949,N_1074,N_3059);
nor U5950 (N_5950,N_26,N_3960);
and U5951 (N_5951,N_4597,N_2554);
and U5952 (N_5952,N_1179,N_716);
or U5953 (N_5953,N_4964,N_3816);
nand U5954 (N_5954,N_1681,N_2271);
nand U5955 (N_5955,N_1156,N_2629);
xnor U5956 (N_5956,N_3775,N_879);
and U5957 (N_5957,N_3033,N_2778);
nor U5958 (N_5958,N_3788,N_3017);
xor U5959 (N_5959,N_333,N_3495);
and U5960 (N_5960,N_212,N_296);
xnor U5961 (N_5961,N_125,N_269);
xnor U5962 (N_5962,N_2781,N_4411);
nand U5963 (N_5963,N_194,N_31);
and U5964 (N_5964,N_51,N_2680);
nand U5965 (N_5965,N_471,N_232);
and U5966 (N_5966,N_1636,N_2572);
and U5967 (N_5967,N_3011,N_3272);
nor U5968 (N_5968,N_1333,N_3202);
nand U5969 (N_5969,N_4127,N_3044);
xnor U5970 (N_5970,N_2499,N_2409);
nand U5971 (N_5971,N_1981,N_4657);
or U5972 (N_5972,N_3848,N_1492);
nor U5973 (N_5973,N_4392,N_1439);
and U5974 (N_5974,N_1594,N_168);
xnor U5975 (N_5975,N_4245,N_449);
or U5976 (N_5976,N_3813,N_2517);
or U5977 (N_5977,N_1008,N_2667);
and U5978 (N_5978,N_330,N_4492);
nor U5979 (N_5979,N_1275,N_3307);
and U5980 (N_5980,N_1245,N_4718);
xnor U5981 (N_5981,N_1092,N_833);
or U5982 (N_5982,N_451,N_3042);
or U5983 (N_5983,N_3172,N_3013);
and U5984 (N_5984,N_2162,N_4104);
xnor U5985 (N_5985,N_3695,N_3557);
or U5986 (N_5986,N_1348,N_4601);
xor U5987 (N_5987,N_1967,N_350);
nand U5988 (N_5988,N_4806,N_4035);
nand U5989 (N_5989,N_4496,N_2570);
or U5990 (N_5990,N_4014,N_2038);
nor U5991 (N_5991,N_1478,N_1424);
and U5992 (N_5992,N_830,N_4206);
nor U5993 (N_5993,N_2223,N_4615);
and U5994 (N_5994,N_3681,N_1346);
nand U5995 (N_5995,N_4589,N_4592);
nand U5996 (N_5996,N_1326,N_136);
and U5997 (N_5997,N_4351,N_552);
or U5998 (N_5998,N_3869,N_1741);
or U5999 (N_5999,N_839,N_173);
or U6000 (N_6000,N_4325,N_4705);
nor U6001 (N_6001,N_4883,N_343);
or U6002 (N_6002,N_75,N_4530);
nand U6003 (N_6003,N_2930,N_3983);
nand U6004 (N_6004,N_3512,N_793);
and U6005 (N_6005,N_3741,N_1595);
and U6006 (N_6006,N_1862,N_106);
xnor U6007 (N_6007,N_2219,N_2622);
nand U6008 (N_6008,N_4476,N_1572);
or U6009 (N_6009,N_1149,N_1278);
xnor U6010 (N_6010,N_3083,N_3222);
xor U6011 (N_6011,N_2737,N_1749);
nor U6012 (N_6012,N_1004,N_932);
or U6013 (N_6013,N_4488,N_1013);
nor U6014 (N_6014,N_4149,N_1141);
nand U6015 (N_6015,N_375,N_4843);
nand U6016 (N_6016,N_3804,N_4486);
nand U6017 (N_6017,N_1668,N_1823);
nand U6018 (N_6018,N_2202,N_1759);
or U6019 (N_6019,N_703,N_429);
xnor U6020 (N_6020,N_736,N_3095);
nand U6021 (N_6021,N_2374,N_3835);
and U6022 (N_6022,N_2283,N_2428);
nand U6023 (N_6023,N_4087,N_1665);
or U6024 (N_6024,N_4412,N_4018);
or U6025 (N_6025,N_711,N_631);
nand U6026 (N_6026,N_2843,N_3399);
nor U6027 (N_6027,N_4758,N_1738);
nand U6028 (N_6028,N_3874,N_1216);
nand U6029 (N_6029,N_2926,N_1364);
xor U6030 (N_6030,N_4610,N_47);
nor U6031 (N_6031,N_1196,N_1688);
and U6032 (N_6032,N_1266,N_456);
and U6033 (N_6033,N_1608,N_4198);
nor U6034 (N_6034,N_3836,N_3212);
nand U6035 (N_6035,N_2488,N_3123);
nand U6036 (N_6036,N_2731,N_1202);
nor U6037 (N_6037,N_497,N_3807);
xor U6038 (N_6038,N_2061,N_843);
xor U6039 (N_6039,N_4799,N_1046);
and U6040 (N_6040,N_3782,N_3053);
xnor U6041 (N_6041,N_2354,N_1984);
xor U6042 (N_6042,N_4122,N_4832);
and U6043 (N_6043,N_3353,N_3483);
nand U6044 (N_6044,N_3475,N_4921);
nor U6045 (N_6045,N_3073,N_1496);
xnor U6046 (N_6046,N_4275,N_2398);
xnor U6047 (N_6047,N_252,N_3535);
and U6048 (N_6048,N_1389,N_4161);
or U6049 (N_6049,N_2114,N_2070);
xnor U6050 (N_6050,N_2520,N_3778);
or U6051 (N_6051,N_4372,N_4836);
and U6052 (N_6052,N_3707,N_3916);
nor U6053 (N_6053,N_3865,N_1799);
xor U6054 (N_6054,N_781,N_2776);
xnor U6055 (N_6055,N_2892,N_1420);
xor U6056 (N_6056,N_2016,N_562);
xor U6057 (N_6057,N_3302,N_4629);
nand U6058 (N_6058,N_2618,N_1995);
nor U6059 (N_6059,N_1947,N_1482);
and U6060 (N_6060,N_3350,N_243);
nor U6061 (N_6061,N_2604,N_3679);
nand U6062 (N_6062,N_1351,N_406);
and U6063 (N_6063,N_4901,N_3022);
nor U6064 (N_6064,N_1510,N_3233);
nor U6065 (N_6065,N_1003,N_2103);
nor U6066 (N_6066,N_2441,N_1132);
nand U6067 (N_6067,N_2794,N_3504);
xnor U6068 (N_6068,N_4379,N_3429);
nor U6069 (N_6069,N_442,N_2904);
xnor U6070 (N_6070,N_352,N_4037);
nand U6071 (N_6071,N_4916,N_2225);
nand U6072 (N_6072,N_3154,N_4334);
nor U6073 (N_6073,N_2511,N_1436);
xnor U6074 (N_6074,N_1698,N_3787);
and U6075 (N_6075,N_4173,N_426);
or U6076 (N_6076,N_4022,N_1804);
and U6077 (N_6077,N_1916,N_1703);
or U6078 (N_6078,N_2163,N_4353);
and U6079 (N_6079,N_4215,N_2976);
or U6080 (N_6080,N_4069,N_1794);
or U6081 (N_6081,N_167,N_2560);
and U6082 (N_6082,N_4663,N_4963);
and U6083 (N_6083,N_1851,N_2924);
nand U6084 (N_6084,N_857,N_2413);
nor U6085 (N_6085,N_3068,N_286);
or U6086 (N_6086,N_3852,N_4966);
nand U6087 (N_6087,N_2915,N_2651);
nand U6088 (N_6088,N_2558,N_4228);
and U6089 (N_6089,N_3738,N_1877);
xnor U6090 (N_6090,N_893,N_601);
nand U6091 (N_6091,N_3652,N_486);
nor U6092 (N_6092,N_763,N_1633);
xor U6093 (N_6093,N_4374,N_4329);
or U6094 (N_6094,N_680,N_3100);
and U6095 (N_6095,N_3867,N_2129);
nor U6096 (N_6096,N_1645,N_1089);
nor U6097 (N_6097,N_1241,N_3067);
or U6098 (N_6098,N_1951,N_1375);
or U6099 (N_6099,N_2474,N_2673);
and U6100 (N_6100,N_4041,N_3527);
nand U6101 (N_6101,N_3773,N_1879);
or U6102 (N_6102,N_3826,N_659);
nor U6103 (N_6103,N_1889,N_3177);
or U6104 (N_6104,N_4734,N_1322);
or U6105 (N_6105,N_4684,N_3388);
nor U6106 (N_6106,N_1066,N_1369);
nor U6107 (N_6107,N_30,N_3318);
and U6108 (N_6108,N_3108,N_602);
or U6109 (N_6109,N_4312,N_654);
nand U6110 (N_6110,N_2148,N_1056);
nand U6111 (N_6111,N_3292,N_1849);
xor U6112 (N_6112,N_4452,N_3496);
xor U6113 (N_6113,N_1265,N_4259);
nand U6114 (N_6114,N_1507,N_1975);
and U6115 (N_6115,N_3706,N_1328);
and U6116 (N_6116,N_1666,N_2592);
and U6117 (N_6117,N_2495,N_223);
xor U6118 (N_6118,N_2801,N_4340);
and U6119 (N_6119,N_3314,N_3);
xor U6120 (N_6120,N_3213,N_3528);
xor U6121 (N_6121,N_750,N_3783);
nor U6122 (N_6122,N_1743,N_2819);
nand U6123 (N_6123,N_1301,N_2733);
nand U6124 (N_6124,N_1994,N_1793);
nor U6125 (N_6125,N_1912,N_412);
and U6126 (N_6126,N_623,N_4404);
or U6127 (N_6127,N_3547,N_3945);
or U6128 (N_6128,N_2565,N_4113);
xor U6129 (N_6129,N_1509,N_1919);
or U6130 (N_6130,N_411,N_1592);
nand U6131 (N_6131,N_3141,N_697);
or U6132 (N_6132,N_639,N_3931);
nor U6133 (N_6133,N_627,N_4911);
and U6134 (N_6134,N_1569,N_941);
nand U6135 (N_6135,N_1286,N_2044);
nand U6136 (N_6136,N_803,N_4667);
xnor U6137 (N_6137,N_73,N_72);
nand U6138 (N_6138,N_1011,N_1412);
xnor U6139 (N_6139,N_4190,N_1371);
and U6140 (N_6140,N_904,N_3142);
xor U6141 (N_6141,N_4068,N_495);
xnor U6142 (N_6142,N_4765,N_2085);
or U6143 (N_6143,N_817,N_314);
xnor U6144 (N_6144,N_354,N_3618);
xor U6145 (N_6145,N_1497,N_848);
and U6146 (N_6146,N_4134,N_1830);
and U6147 (N_6147,N_3705,N_499);
and U6148 (N_6148,N_2594,N_1442);
nor U6149 (N_6149,N_1443,N_1825);
or U6150 (N_6150,N_2433,N_2791);
nor U6151 (N_6151,N_4881,N_4251);
xnor U6152 (N_6152,N_3766,N_955);
or U6153 (N_6153,N_828,N_1922);
nor U6154 (N_6154,N_1973,N_2481);
nor U6155 (N_6155,N_1010,N_4690);
and U6156 (N_6156,N_1291,N_586);
xnor U6157 (N_6157,N_4368,N_963);
xor U6158 (N_6158,N_4591,N_2305);
xnor U6159 (N_6159,N_4960,N_2962);
nand U6160 (N_6160,N_2141,N_4854);
xor U6161 (N_6161,N_4829,N_1114);
xnor U6162 (N_6162,N_4981,N_1504);
or U6163 (N_6163,N_1843,N_744);
nand U6164 (N_6164,N_4003,N_1961);
nand U6165 (N_6165,N_1109,N_434);
and U6166 (N_6166,N_2630,N_4328);
nor U6167 (N_6167,N_255,N_787);
nor U6168 (N_6168,N_131,N_567);
nand U6169 (N_6169,N_38,N_513);
xor U6170 (N_6170,N_2751,N_870);
xnor U6171 (N_6171,N_3629,N_4602);
nand U6172 (N_6172,N_836,N_1123);
or U6173 (N_6173,N_4085,N_1122);
xnor U6174 (N_6174,N_87,N_1130);
nand U6175 (N_6175,N_1340,N_4235);
nand U6176 (N_6176,N_1172,N_1488);
nand U6177 (N_6177,N_4279,N_4577);
nand U6178 (N_6178,N_4094,N_3571);
and U6179 (N_6179,N_4946,N_3563);
nor U6180 (N_6180,N_2589,N_4154);
nand U6181 (N_6181,N_4902,N_2746);
xnor U6182 (N_6182,N_2470,N_1043);
or U6183 (N_6183,N_3034,N_281);
xnor U6184 (N_6184,N_2465,N_4800);
xnor U6185 (N_6185,N_507,N_3395);
or U6186 (N_6186,N_1885,N_1578);
and U6187 (N_6187,N_1542,N_3550);
nor U6188 (N_6188,N_4792,N_4506);
xnor U6189 (N_6189,N_221,N_2870);
xor U6190 (N_6190,N_3808,N_2256);
nor U6191 (N_6191,N_4121,N_1244);
xor U6192 (N_6192,N_2424,N_3048);
nand U6193 (N_6193,N_3277,N_4082);
or U6194 (N_6194,N_3003,N_3850);
nand U6195 (N_6195,N_4500,N_1544);
nand U6196 (N_6196,N_109,N_658);
or U6197 (N_6197,N_4347,N_547);
and U6198 (N_6198,N_2822,N_4853);
or U6199 (N_6199,N_1051,N_971);
xor U6200 (N_6200,N_2646,N_3620);
xnor U6201 (N_6201,N_2890,N_1247);
nand U6202 (N_6202,N_3418,N_3799);
and U6203 (N_6203,N_3074,N_389);
or U6204 (N_6204,N_2636,N_3487);
nor U6205 (N_6205,N_3237,N_1904);
nor U6206 (N_6206,N_886,N_4031);
nand U6207 (N_6207,N_2054,N_2234);
and U6208 (N_6208,N_2008,N_4176);
or U6209 (N_6209,N_399,N_2158);
nor U6210 (N_6210,N_3762,N_1714);
or U6211 (N_6211,N_2535,N_493);
nand U6212 (N_6212,N_4219,N_590);
nand U6213 (N_6213,N_4924,N_432);
or U6214 (N_6214,N_91,N_257);
and U6215 (N_6215,N_3968,N_3499);
nor U6216 (N_6216,N_260,N_1471);
nor U6217 (N_6217,N_4084,N_4999);
nand U6218 (N_6218,N_1129,N_2541);
or U6219 (N_6219,N_4930,N_2292);
and U6220 (N_6220,N_2823,N_1797);
nand U6221 (N_6221,N_4380,N_713);
nor U6222 (N_6222,N_18,N_1589);
xor U6223 (N_6223,N_1127,N_4434);
nand U6224 (N_6224,N_969,N_3903);
nand U6225 (N_6225,N_2201,N_2293);
nand U6226 (N_6226,N_4618,N_2430);
nor U6227 (N_6227,N_46,N_732);
or U6228 (N_6228,N_6,N_3061);
and U6229 (N_6229,N_696,N_2209);
nand U6230 (N_6230,N_1697,N_4348);
nand U6231 (N_6231,N_267,N_1117);
and U6232 (N_6232,N_3046,N_3262);
or U6233 (N_6233,N_2841,N_2753);
and U6234 (N_6234,N_1930,N_819);
nor U6235 (N_6235,N_4057,N_2859);
xnor U6236 (N_6236,N_3714,N_2872);
and U6237 (N_6237,N_4079,N_719);
or U6238 (N_6238,N_3950,N_3367);
nor U6239 (N_6239,N_288,N_801);
xor U6240 (N_6240,N_1426,N_1490);
xor U6241 (N_6241,N_635,N_2995);
or U6242 (N_6242,N_846,N_1180);
or U6243 (N_6243,N_1634,N_4326);
xor U6244 (N_6244,N_4136,N_4098);
xnor U6245 (N_6245,N_1953,N_543);
or U6246 (N_6246,N_3748,N_2132);
or U6247 (N_6247,N_3026,N_780);
nor U6248 (N_6248,N_3243,N_2249);
xnor U6249 (N_6249,N_2933,N_2032);
or U6250 (N_6250,N_931,N_3340);
and U6251 (N_6251,N_823,N_215);
and U6252 (N_6252,N_2779,N_3736);
nor U6253 (N_6253,N_4970,N_2306);
or U6254 (N_6254,N_1273,N_3255);
xnor U6255 (N_6255,N_2580,N_2621);
and U6256 (N_6256,N_946,N_3687);
nand U6257 (N_6257,N_3686,N_2356);
nor U6258 (N_6258,N_3995,N_3689);
or U6259 (N_6259,N_734,N_417);
xor U6260 (N_6260,N_2026,N_4020);
and U6261 (N_6261,N_4723,N_3373);
nand U6262 (N_6262,N_3818,N_1287);
xor U6263 (N_6263,N_875,N_4782);
nor U6264 (N_6264,N_3765,N_2310);
nand U6265 (N_6265,N_4438,N_3035);
nor U6266 (N_6266,N_1095,N_2518);
or U6267 (N_6267,N_42,N_580);
or U6268 (N_6268,N_1982,N_4471);
xor U6269 (N_6269,N_3428,N_1511);
xor U6270 (N_6270,N_4626,N_2406);
and U6271 (N_6271,N_2562,N_4373);
and U6272 (N_6272,N_4606,N_3371);
and U6273 (N_6273,N_2557,N_974);
or U6274 (N_6274,N_3892,N_4764);
nor U6275 (N_6275,N_4156,N_660);
nor U6276 (N_6276,N_3188,N_3135);
nor U6277 (N_6277,N_3856,N_3384);
nand U6278 (N_6278,N_4826,N_218);
xnor U6279 (N_6279,N_4425,N_2762);
nand U6280 (N_6280,N_975,N_1296);
xor U6281 (N_6281,N_1076,N_1720);
and U6282 (N_6282,N_3049,N_3375);
nand U6283 (N_6283,N_402,N_699);
xor U6284 (N_6284,N_2974,N_4406);
xnor U6285 (N_6285,N_1800,N_1263);
and U6286 (N_6286,N_4681,N_1600);
or U6287 (N_6287,N_3111,N_3448);
or U6288 (N_6288,N_4446,N_1350);
xor U6289 (N_6289,N_1993,N_4565);
nor U6290 (N_6290,N_1378,N_2689);
nor U6291 (N_6291,N_1220,N_3472);
xnor U6292 (N_6292,N_1246,N_2309);
and U6293 (N_6293,N_4002,N_1234);
nand U6294 (N_6294,N_103,N_1731);
xor U6295 (N_6295,N_1038,N_3829);
and U6296 (N_6296,N_2078,N_424);
xnor U6297 (N_6297,N_3657,N_4150);
nor U6298 (N_6298,N_4674,N_1481);
nand U6299 (N_6299,N_2684,N_2446);
or U6300 (N_6300,N_1568,N_2260);
and U6301 (N_6301,N_9,N_3253);
xnor U6302 (N_6302,N_4000,N_118);
and U6303 (N_6303,N_2023,N_3176);
nand U6304 (N_6304,N_4354,N_2377);
nand U6305 (N_6305,N_4991,N_2706);
or U6306 (N_6306,N_2975,N_4635);
nand U6307 (N_6307,N_2954,N_619);
xnor U6308 (N_6308,N_4821,N_2390);
nand U6309 (N_6309,N_915,N_4934);
or U6310 (N_6310,N_2196,N_3116);
or U6311 (N_6311,N_3643,N_1344);
or U6312 (N_6312,N_3182,N_4205);
xor U6313 (N_6313,N_484,N_325);
and U6314 (N_6314,N_175,N_888);
and U6315 (N_6315,N_4343,N_3912);
nand U6316 (N_6316,N_2624,N_35);
or U6317 (N_6317,N_4513,N_3479);
and U6318 (N_6318,N_1707,N_1617);
nor U6319 (N_6319,N_4653,N_3394);
or U6320 (N_6320,N_3150,N_3653);
or U6321 (N_6321,N_4108,N_1590);
xnor U6322 (N_6322,N_1200,N_3805);
nand U6323 (N_6323,N_4209,N_3181);
nor U6324 (N_6324,N_841,N_2443);
or U6325 (N_6325,N_958,N_4202);
xnor U6326 (N_6326,N_143,N_2198);
or U6327 (N_6327,N_1779,N_4547);
nand U6328 (N_6328,N_3052,N_2244);
or U6329 (N_6329,N_4575,N_1085);
xnor U6330 (N_6330,N_1166,N_4561);
and U6331 (N_6331,N_4297,N_3368);
and U6332 (N_6332,N_1610,N_2359);
or U6333 (N_6333,N_309,N_111);
nand U6334 (N_6334,N_962,N_2157);
xnor U6335 (N_6335,N_76,N_245);
and U6336 (N_6336,N_83,N_482);
nand U6337 (N_6337,N_1098,N_3769);
xor U6338 (N_6338,N_3480,N_2925);
nor U6339 (N_6339,N_2917,N_4240);
xnor U6340 (N_6340,N_2227,N_3708);
and U6341 (N_6341,N_1815,N_1534);
or U6342 (N_6342,N_3998,N_2364);
or U6343 (N_6343,N_723,N_1262);
and U6344 (N_6344,N_271,N_2615);
or U6345 (N_6345,N_2418,N_4724);
nand U6346 (N_6346,N_4,N_1221);
nor U6347 (N_6347,N_1763,N_2468);
xnor U6348 (N_6348,N_2001,N_1219);
and U6349 (N_6349,N_501,N_4879);
nand U6350 (N_6350,N_2591,N_2164);
and U6351 (N_6351,N_478,N_4388);
nand U6352 (N_6352,N_1280,N_2567);
or U6353 (N_6353,N_1002,N_900);
xnor U6354 (N_6354,N_1808,N_640);
xnor U6355 (N_6355,N_4607,N_3209);
nor U6356 (N_6356,N_4461,N_1577);
nor U6357 (N_6357,N_2548,N_3843);
or U6358 (N_6358,N_3275,N_4859);
and U6359 (N_6359,N_2834,N_239);
nand U6360 (N_6360,N_4707,N_292);
xor U6361 (N_6361,N_385,N_1268);
xnor U6362 (N_6362,N_3644,N_1866);
or U6363 (N_6363,N_157,N_4952);
nand U6364 (N_6364,N_3285,N_806);
nor U6365 (N_6365,N_1966,N_3498);
and U6366 (N_6366,N_1555,N_4941);
or U6367 (N_6367,N_2979,N_766);
nor U6368 (N_6368,N_934,N_3199);
and U6369 (N_6369,N_3989,N_3969);
xnor U6370 (N_6370,N_2540,N_4581);
nor U6371 (N_6371,N_1012,N_815);
or U6372 (N_6372,N_1,N_2921);
xnor U6373 (N_6373,N_1901,N_3349);
or U6374 (N_6374,N_2022,N_2693);
xnor U6375 (N_6375,N_1034,N_2509);
or U6376 (N_6376,N_2175,N_2024);
xor U6377 (N_6377,N_1736,N_2768);
and U6378 (N_6378,N_4882,N_3588);
and U6379 (N_6379,N_3273,N_4163);
or U6380 (N_6380,N_3101,N_4858);
xor U6381 (N_6381,N_2104,N_1447);
xor U6382 (N_6382,N_2911,N_901);
or U6383 (N_6383,N_3890,N_4586);
or U6384 (N_6384,N_4377,N_3771);
or U6385 (N_6385,N_2473,N_439);
or U6386 (N_6386,N_322,N_1498);
nor U6387 (N_6387,N_1661,N_3971);
xor U6388 (N_6388,N_638,N_2381);
nand U6389 (N_6389,N_1468,N_709);
nand U6390 (N_6390,N_1324,N_2447);
nor U6391 (N_6391,N_2714,N_3058);
or U6392 (N_6392,N_462,N_521);
nor U6393 (N_6393,N_4116,N_2804);
nor U6394 (N_6394,N_1929,N_760);
or U6395 (N_6395,N_4833,N_2810);
xor U6396 (N_6396,N_3239,N_1032);
nor U6397 (N_6397,N_3591,N_285);
and U6398 (N_6398,N_3567,N_408);
xor U6399 (N_6399,N_1539,N_274);
nor U6400 (N_6400,N_2076,N_1563);
xor U6401 (N_6401,N_3980,N_4660);
xor U6402 (N_6402,N_477,N_3500);
and U6403 (N_6403,N_1005,N_4819);
nor U6404 (N_6404,N_2189,N_1655);
nand U6405 (N_6405,N_1931,N_1659);
and U6406 (N_6406,N_2071,N_1362);
xnor U6407 (N_6407,N_387,N_4148);
xor U6408 (N_6408,N_725,N_3186);
nand U6409 (N_6409,N_1039,N_374);
or U6410 (N_6410,N_2561,N_795);
and U6411 (N_6411,N_816,N_1113);
nand U6412 (N_6412,N_4281,N_2212);
nor U6413 (N_6413,N_3408,N_868);
or U6414 (N_6414,N_3029,N_4741);
or U6415 (N_6415,N_1710,N_3389);
or U6416 (N_6416,N_2058,N_3126);
nand U6417 (N_6417,N_4105,N_220);
or U6418 (N_6418,N_1031,N_2028);
or U6419 (N_6419,N_4264,N_254);
or U6420 (N_6420,N_842,N_4253);
nand U6421 (N_6421,N_582,N_648);
and U6422 (N_6422,N_105,N_4709);
xor U6423 (N_6423,N_2388,N_3369);
or U6424 (N_6424,N_1693,N_1570);
nand U6425 (N_6425,N_3776,N_4067);
nand U6426 (N_6426,N_1390,N_4252);
nor U6427 (N_6427,N_3060,N_3796);
xnor U6428 (N_6428,N_2704,N_2010);
nand U6429 (N_6429,N_4541,N_3409);
or U6430 (N_6430,N_4016,N_1796);
and U6431 (N_6431,N_2575,N_4553);
nand U6432 (N_6432,N_3444,N_512);
and U6433 (N_6433,N_4387,N_2657);
xor U6434 (N_6434,N_4776,N_1745);
nand U6435 (N_6435,N_2101,N_1597);
nor U6436 (N_6436,N_651,N_4827);
nor U6437 (N_6437,N_3343,N_2515);
nor U6438 (N_6438,N_179,N_4769);
xnor U6439 (N_6439,N_3122,N_880);
nand U6440 (N_6440,N_490,N_2122);
xnor U6441 (N_6441,N_3344,N_2427);
and U6442 (N_6442,N_4390,N_811);
xor U6443 (N_6443,N_4015,N_455);
xor U6444 (N_6444,N_779,N_768);
nor U6445 (N_6445,N_4250,N_4429);
and U6446 (N_6446,N_2655,N_2990);
xnor U6447 (N_6447,N_4750,N_574);
xor U6448 (N_6448,N_2040,N_873);
or U6449 (N_6449,N_662,N_1658);
nor U6450 (N_6450,N_3304,N_4045);
nand U6451 (N_6451,N_463,N_3094);
or U6452 (N_6452,N_3354,N_2047);
xor U6453 (N_6453,N_19,N_555);
nand U6454 (N_6454,N_3646,N_4888);
or U6455 (N_6455,N_2303,N_2231);
nand U6456 (N_6456,N_1733,N_4316);
nor U6457 (N_6457,N_3422,N_40);
nor U6458 (N_6458,N_444,N_745);
nand U6459 (N_6459,N_3440,N_2682);
nand U6460 (N_6460,N_3293,N_4784);
and U6461 (N_6461,N_1809,N_2542);
nor U6462 (N_6462,N_2866,N_4043);
xor U6463 (N_6463,N_503,N_3648);
nor U6464 (N_6464,N_4682,N_2502);
xnor U6465 (N_6465,N_897,N_2412);
or U6466 (N_6466,N_3792,N_2331);
xor U6467 (N_6467,N_2988,N_1270);
or U6468 (N_6468,N_438,N_1300);
or U6469 (N_6469,N_644,N_2623);
xnor U6470 (N_6470,N_2874,N_961);
and U6471 (N_6471,N_155,N_2376);
and U6472 (N_6472,N_1283,N_2770);
or U6473 (N_6473,N_1586,N_4185);
nor U6474 (N_6474,N_4869,N_1088);
xnor U6475 (N_6475,N_532,N_1274);
nor U6476 (N_6476,N_3451,N_4756);
or U6477 (N_6477,N_2767,N_2813);
xor U6478 (N_6478,N_1352,N_2537);
and U6479 (N_6479,N_4313,N_4280);
nand U6480 (N_6480,N_3628,N_3966);
and U6481 (N_6481,N_3161,N_1189);
nand U6482 (N_6482,N_1374,N_1635);
xor U6483 (N_6483,N_3814,N_2649);
or U6484 (N_6484,N_110,N_2963);
nand U6485 (N_6485,N_2490,N_3599);
xnor U6486 (N_6486,N_1184,N_150);
and U6487 (N_6487,N_2358,N_3970);
nand U6488 (N_6488,N_3110,N_1142);
nor U6489 (N_6489,N_642,N_117);
or U6490 (N_6490,N_3231,N_465);
nand U6491 (N_6491,N_1035,N_3609);
nand U6492 (N_6492,N_1868,N_1409);
or U6493 (N_6493,N_522,N_58);
or U6494 (N_6494,N_4992,N_3173);
nand U6495 (N_6495,N_578,N_3568);
or U6496 (N_6496,N_3861,N_2280);
xnor U6497 (N_6497,N_2042,N_994);
xor U6498 (N_6498,N_1639,N_4323);
and U6499 (N_6499,N_2878,N_4990);
or U6500 (N_6500,N_2521,N_1238);
or U6501 (N_6501,N_845,N_871);
nand U6502 (N_6502,N_2005,N_2300);
xor U6503 (N_6503,N_4179,N_1876);
and U6504 (N_6504,N_4609,N_1431);
xor U6505 (N_6505,N_3732,N_4304);
xor U6506 (N_6506,N_2007,N_2037);
nand U6507 (N_6507,N_2740,N_740);
nand U6508 (N_6508,N_4168,N_1675);
nor U6509 (N_6509,N_4039,N_2551);
xor U6510 (N_6510,N_3427,N_3548);
nand U6511 (N_6511,N_2327,N_318);
nand U6512 (N_6512,N_4296,N_3611);
nand U6513 (N_6513,N_2829,N_3606);
and U6514 (N_6514,N_4767,N_2716);
and U6515 (N_6515,N_838,N_3625);
nor U6516 (N_6516,N_1314,N_3797);
xor U6517 (N_6517,N_666,N_2437);
xnor U6518 (N_6518,N_2508,N_4208);
and U6519 (N_6519,N_1628,N_884);
nand U6520 (N_6520,N_2564,N_1394);
nor U6521 (N_6521,N_2304,N_4948);
and U6522 (N_6522,N_2345,N_4019);
or U6523 (N_6523,N_2341,N_3317);
and U6524 (N_6524,N_1611,N_3542);
nor U6525 (N_6525,N_3767,N_4073);
xnor U6526 (N_6526,N_2969,N_2650);
nand U6527 (N_6527,N_3798,N_649);
nor U6528 (N_6528,N_2365,N_4661);
and U6529 (N_6529,N_2633,N_2251);
or U6530 (N_6530,N_3556,N_4181);
and U6531 (N_6531,N_4549,N_824);
nand U6532 (N_6532,N_4053,N_2238);
or U6533 (N_6533,N_1450,N_2073);
or U6534 (N_6534,N_63,N_4622);
nand U6535 (N_6535,N_3432,N_3331);
and U6536 (N_6536,N_2031,N_189);
xor U6537 (N_6537,N_1615,N_1385);
and U6538 (N_6538,N_2180,N_2402);
and U6539 (N_6539,N_4221,N_3063);
nor U6540 (N_6540,N_4324,N_4362);
nor U6541 (N_6541,N_2910,N_4178);
or U6542 (N_6542,N_226,N_154);
xor U6543 (N_6543,N_1936,N_1873);
nand U6544 (N_6544,N_213,N_813);
xnor U6545 (N_6545,N_2480,N_3162);
nand U6546 (N_6546,N_1356,N_4604);
and U6547 (N_6547,N_2096,N_2006);
nand U6548 (N_6548,N_3045,N_4732);
nand U6549 (N_6549,N_2207,N_2833);
nand U6550 (N_6550,N_973,N_1026);
xnor U6551 (N_6551,N_3376,N_1384);
or U6552 (N_6552,N_1407,N_4103);
and U6553 (N_6553,N_2348,N_2161);
or U6554 (N_6554,N_1152,N_2074);
xnor U6555 (N_6555,N_1689,N_3183);
nand U6556 (N_6556,N_1903,N_4417);
xnor U6557 (N_6557,N_749,N_1358);
and U6558 (N_6558,N_199,N_2836);
nor U6559 (N_6559,N_1651,N_55);
xor U6560 (N_6560,N_2725,N_3463);
xor U6561 (N_6561,N_3210,N_431);
xnor U6562 (N_6562,N_919,N_3037);
nand U6563 (N_6563,N_4111,N_3036);
xnor U6564 (N_6564,N_2929,N_2861);
nor U6565 (N_6565,N_1820,N_2940);
and U6566 (N_6566,N_2642,N_2426);
nand U6567 (N_6567,N_3923,N_2208);
or U6568 (N_6568,N_1752,N_3211);
xnor U6569 (N_6569,N_3225,N_2628);
nor U6570 (N_6570,N_3398,N_1252);
or U6571 (N_6571,N_2455,N_1377);
or U6572 (N_6572,N_2246,N_4936);
nor U6573 (N_6573,N_4868,N_1834);
xor U6574 (N_6574,N_4360,N_1874);
xnor U6575 (N_6575,N_2136,N_3323);
or U6576 (N_6576,N_97,N_390);
xnor U6577 (N_6577,N_2736,N_1255);
xor U6578 (N_6578,N_2448,N_2968);
nand U6579 (N_6579,N_4494,N_88);
or U6580 (N_6580,N_504,N_3617);
nand U6581 (N_6581,N_1249,N_4342);
and U6582 (N_6582,N_4558,N_4177);
and U6583 (N_6583,N_3385,N_943);
nand U6584 (N_6584,N_4937,N_2947);
or U6585 (N_6585,N_1613,N_784);
xor U6586 (N_6586,N_4804,N_3417);
xor U6587 (N_6587,N_1212,N_691);
nand U6588 (N_6588,N_4319,N_1472);
xnor U6589 (N_6589,N_1258,N_1171);
and U6590 (N_6590,N_4914,N_4490);
nand U6591 (N_6591,N_3217,N_4809);
and U6592 (N_6592,N_4907,N_1451);
nand U6593 (N_6593,N_1991,N_3857);
and U6594 (N_6594,N_3386,N_2734);
or U6595 (N_6595,N_1015,N_1440);
or U6596 (N_6596,N_3552,N_3893);
nor U6597 (N_6597,N_3577,N_1602);
nor U6598 (N_6598,N_4655,N_4773);
xor U6599 (N_6599,N_3130,N_3973);
xor U6600 (N_6600,N_183,N_3190);
and U6601 (N_6601,N_4917,N_4365);
and U6602 (N_6602,N_3120,N_4569);
or U6603 (N_6603,N_2965,N_4696);
nor U6604 (N_6604,N_3092,N_3929);
nor U6605 (N_6605,N_3873,N_2899);
nand U6606 (N_6606,N_3526,N_4225);
or U6607 (N_6607,N_1503,N_4248);
or U6608 (N_6608,N_777,N_2805);
or U6609 (N_6609,N_2117,N_1419);
xnor U6610 (N_6610,N_116,N_3447);
xnor U6611 (N_6611,N_2068,N_2808);
and U6612 (N_6612,N_4722,N_3612);
and U6613 (N_6613,N_4364,N_4583);
nand U6614 (N_6614,N_3131,N_4508);
or U6615 (N_6615,N_2320,N_1631);
or U6616 (N_6616,N_4473,N_3671);
and U6617 (N_6617,N_4736,N_953);
or U6618 (N_6618,N_414,N_3105);
nand U6619 (N_6619,N_4158,N_1923);
nor U6620 (N_6620,N_3238,N_728);
nand U6621 (N_6621,N_3436,N_1006);
or U6622 (N_6622,N_1014,N_1940);
nor U6623 (N_6623,N_2555,N_704);
nor U6624 (N_6624,N_2625,N_1566);
nand U6625 (N_6625,N_3975,N_1423);
xnor U6626 (N_6626,N_3532,N_4440);
nand U6627 (N_6627,N_60,N_187);
xnor U6628 (N_6628,N_3338,N_481);
nand U6629 (N_6629,N_2755,N_809);
nand U6630 (N_6630,N_4292,N_2419);
and U6631 (N_6631,N_2065,N_1422);
or U6632 (N_6632,N_2155,N_2891);
xor U6633 (N_6633,N_3441,N_4192);
nor U6634 (N_6634,N_1518,N_2440);
nand U6635 (N_6635,N_3602,N_4831);
xnor U6636 (N_6636,N_1652,N_185);
xor U6637 (N_6637,N_3192,N_4477);
xor U6638 (N_6638,N_3071,N_1864);
nand U6639 (N_6639,N_885,N_615);
and U6640 (N_6640,N_3791,N_1802);
or U6641 (N_6641,N_3282,N_3414);
xor U6642 (N_6642,N_3078,N_528);
xnor U6643 (N_6643,N_825,N_3403);
and U6644 (N_6644,N_2452,N_3641);
xnor U6645 (N_6645,N_1650,N_3031);
xnor U6646 (N_6646,N_3864,N_188);
nor U6647 (N_6647,N_1770,N_661);
xor U6648 (N_6648,N_4738,N_2677);
nand U6649 (N_6649,N_1718,N_2631);
and U6650 (N_6650,N_2092,N_3137);
xnor U6651 (N_6651,N_2366,N_1727);
nor U6652 (N_6652,N_4678,N_1527);
nor U6653 (N_6653,N_320,N_1494);
xnor U6654 (N_6654,N_1700,N_1696);
nand U6655 (N_6655,N_4962,N_3809);
xor U6656 (N_6656,N_3456,N_130);
xor U6657 (N_6657,N_589,N_4017);
or U6658 (N_6658,N_1486,N_3460);
and U6659 (N_6659,N_418,N_2513);
or U6660 (N_6660,N_3038,N_2647);
and U6661 (N_6661,N_3009,N_2241);
nand U6662 (N_6662,N_3658,N_1373);
nor U6663 (N_6663,N_2598,N_3693);
and U6664 (N_6664,N_3064,N_3608);
or U6665 (N_6665,N_351,N_4419);
nand U6666 (N_6666,N_4838,N_327);
nor U6667 (N_6667,N_4654,N_1687);
or U6668 (N_6668,N_123,N_4038);
and U6669 (N_6669,N_614,N_466);
nand U6670 (N_6670,N_177,N_4751);
or U6671 (N_6671,N_4184,N_3229);
nor U6672 (N_6672,N_3204,N_1000);
nand U6673 (N_6673,N_3374,N_2127);
and U6674 (N_6674,N_2577,N_3906);
and U6675 (N_6675,N_4906,N_3308);
nand U6676 (N_6676,N_371,N_2125);
or U6677 (N_6677,N_4802,N_13);
nand U6678 (N_6678,N_3206,N_487);
or U6679 (N_6679,N_3406,N_832);
or U6680 (N_6680,N_4011,N_3138);
xnor U6681 (N_6681,N_4710,N_2987);
or U6682 (N_6682,N_321,N_3566);
nand U6683 (N_6683,N_887,N_1822);
or U6684 (N_6684,N_715,N_4414);
and U6685 (N_6685,N_2944,N_4396);
xnor U6686 (N_6686,N_2912,N_2211);
nand U6687 (N_6687,N_1833,N_2868);
or U6688 (N_6688,N_2788,N_4822);
or U6689 (N_6689,N_241,N_2295);
nand U6690 (N_6690,N_3051,N_1310);
and U6691 (N_6691,N_2851,N_4303);
nor U6692 (N_6692,N_4109,N_1585);
xor U6693 (N_6693,N_4102,N_1159);
nand U6694 (N_6694,N_569,N_1144);
nor U6695 (N_6695,N_1646,N_746);
or U6696 (N_6696,N_1379,N_4632);
or U6697 (N_6697,N_1163,N_4231);
xnor U6698 (N_6698,N_1960,N_441);
nor U6699 (N_6699,N_2370,N_923);
or U6700 (N_6700,N_3442,N_219);
nand U6701 (N_6701,N_1530,N_2927);
nand U6702 (N_6702,N_3157,N_1591);
and U6703 (N_6703,N_2290,N_523);
and U6704 (N_6704,N_3446,N_980);
or U6705 (N_6705,N_2400,N_4044);
and U6706 (N_6706,N_3955,N_3477);
nor U6707 (N_6707,N_1368,N_2800);
or U6708 (N_6708,N_3889,N_4984);
nand U6709 (N_6709,N_443,N_2881);
nand U6710 (N_6710,N_2617,N_124);
and U6711 (N_6711,N_4908,N_2138);
xnor U6712 (N_6712,N_1094,N_1138);
and U6713 (N_6713,N_1535,N_2605);
xor U6714 (N_6714,N_4510,N_3258);
or U6715 (N_6715,N_2100,N_2826);
or U6716 (N_6716,N_508,N_505);
xnor U6717 (N_6717,N_682,N_4731);
nor U6718 (N_6718,N_4588,N_4433);
xnor U6719 (N_6719,N_258,N_3077);
nor U6720 (N_6720,N_304,N_2879);
and U6721 (N_6721,N_2318,N_2893);
and U6722 (N_6722,N_2326,N_4566);
xor U6723 (N_6723,N_1282,N_2750);
nand U6724 (N_6724,N_4649,N_4770);
nor U6725 (N_6725,N_1777,N_4877);
and U6726 (N_6726,N_3359,N_4080);
xor U6727 (N_6727,N_4289,N_2639);
nor U6728 (N_6728,N_4502,N_4207);
xnor U6729 (N_6729,N_3739,N_1721);
and U6730 (N_6730,N_4891,N_2214);
or U6731 (N_6731,N_4426,N_4825);
or U6732 (N_6732,N_368,N_2133);
or U6733 (N_6733,N_4813,N_4261);
and U6734 (N_6734,N_3325,N_1226);
nand U6735 (N_6735,N_61,N_3312);
nand U6736 (N_6736,N_4754,N_459);
and U6737 (N_6737,N_1376,N_3847);
and U6738 (N_6738,N_181,N_988);
xnor U6739 (N_6739,N_2109,N_4445);
xnor U6740 (N_6740,N_1963,N_3924);
nor U6741 (N_6741,N_275,N_1826);
nor U6742 (N_6742,N_3160,N_80);
nand U6743 (N_6743,N_4307,N_1583);
xor U6744 (N_6744,N_525,N_1979);
or U6745 (N_6745,N_4559,N_4743);
nor U6746 (N_6746,N_3166,N_4711);
nor U6747 (N_6747,N_4519,N_3303);
and U6748 (N_6748,N_3193,N_603);
xnor U6749 (N_6749,N_533,N_1435);
or U6750 (N_6750,N_370,N_4810);
and U6751 (N_6751,N_2278,N_208);
and U6752 (N_6752,N_3021,N_4410);
xor U6753 (N_6753,N_606,N_28);
and U6754 (N_6754,N_56,N_1893);
xor U6755 (N_6755,N_4556,N_3316);
and U6756 (N_6756,N_3284,N_1546);
nand U6757 (N_6757,N_996,N_2072);
or U6758 (N_6758,N_3665,N_1579);
or U6759 (N_6759,N_808,N_4349);
nand U6760 (N_6760,N_895,N_1131);
nor U6761 (N_6761,N_542,N_882);
or U6762 (N_6762,N_3327,N_2476);
nand U6763 (N_6763,N_4007,N_4735);
nand U6764 (N_6764,N_1227,N_1413);
and U6765 (N_6765,N_2838,N_4470);
nor U6766 (N_6766,N_3127,N_1934);
nor U6767 (N_6767,N_1971,N_939);
and U6768 (N_6768,N_4798,N_668);
nor U6769 (N_6769,N_178,N_4332);
nand U6770 (N_6770,N_336,N_1288);
and U6771 (N_6771,N_3565,N_4194);
xor U6772 (N_6772,N_752,N_705);
nand U6773 (N_6773,N_3434,N_25);
and U6774 (N_6774,N_565,N_991);
and U6775 (N_6775,N_464,N_3756);
nor U6776 (N_6776,N_3201,N_2635);
or U6777 (N_6777,N_3426,N_182);
or U6778 (N_6778,N_4409,N_3424);
nand U6779 (N_6779,N_4126,N_1232);
and U6780 (N_6780,N_3660,N_3070);
and U6781 (N_6781,N_1256,N_133);
nor U6782 (N_6782,N_976,N_3087);
nor U6783 (N_6783,N_4640,N_3507);
nor U6784 (N_6784,N_1909,N_3875);
nor U6785 (N_6785,N_4128,N_1609);
or U6786 (N_6786,N_820,N_5);
and U6787 (N_6787,N_2274,N_4969);
xnor U6788 (N_6788,N_1207,N_3810);
and U6789 (N_6789,N_3582,N_2273);
nand U6790 (N_6790,N_2730,N_4211);
nor U6791 (N_6791,N_2462,N_3015);
and U6792 (N_6792,N_2003,N_282);
nor U6793 (N_6793,N_3269,N_1317);
and U6794 (N_6794,N_396,N_2582);
nor U6795 (N_6795,N_3280,N_2057);
xnor U6796 (N_6796,N_1905,N_1787);
nor U6797 (N_6797,N_673,N_718);
nand U6798 (N_6798,N_134,N_1788);
or U6799 (N_6799,N_515,N_4605);
nand U6800 (N_6800,N_4491,N_3086);
nor U6801 (N_6801,N_2696,N_1186);
or U6802 (N_6802,N_4186,N_2784);
nor U6803 (N_6803,N_2475,N_3484);
and U6804 (N_6804,N_2583,N_4787);
and U6805 (N_6805,N_4314,N_2393);
or U6806 (N_6806,N_3650,N_2786);
nor U6807 (N_6807,N_599,N_1272);
nor U6808 (N_6808,N_3963,N_3294);
nor U6809 (N_6809,N_925,N_1134);
xnor U6810 (N_6810,N_148,N_388);
xor U6811 (N_6811,N_3777,N_3322);
xnor U6812 (N_6812,N_3900,N_775);
nor U6813 (N_6813,N_4294,N_3640);
and U6814 (N_6814,N_4531,N_3594);
nor U6815 (N_6815,N_4115,N_3133);
xor U6816 (N_6816,N_4835,N_2391);
nor U6817 (N_6817,N_2492,N_2875);
nor U6818 (N_6818,N_2529,N_4925);
nor U6819 (N_6819,N_2143,N_2156);
and U6820 (N_6820,N_2317,N_4584);
nor U6821 (N_6821,N_1524,N_739);
nand U6822 (N_6822,N_1565,N_1111);
or U6823 (N_6823,N_4580,N_1601);
xnor U6824 (N_6824,N_3579,N_1854);
xnor U6825 (N_6825,N_1119,N_2777);
and U6826 (N_6826,N_3751,N_4884);
xor U6827 (N_6827,N_280,N_2919);
and U6828 (N_6828,N_2747,N_1746);
and U6829 (N_6829,N_1185,N_2425);
nand U6830 (N_6830,N_2097,N_1416);
or U6831 (N_6831,N_2218,N_206);
and U6832 (N_6832,N_1987,N_724);
nor U6833 (N_6833,N_3466,N_2550);
and U6834 (N_6834,N_1983,N_583);
nor U6835 (N_6835,N_2226,N_4287);
nand U6836 (N_6836,N_3974,N_4611);
or U6837 (N_6837,N_2191,N_1495);
and U6838 (N_6838,N_675,N_2124);
xor U6839 (N_6839,N_3215,N_4544);
nand U6840 (N_6840,N_3543,N_3457);
xor U6841 (N_6841,N_2998,N_3822);
and U6842 (N_6842,N_2759,N_2279);
or U6843 (N_6843,N_3259,N_4894);
or U6844 (N_6844,N_2862,N_1045);
nor U6845 (N_6845,N_1470,N_1408);
xnor U6846 (N_6846,N_2959,N_1593);
nor U6847 (N_6847,N_500,N_1647);
and U6848 (N_6848,N_2086,N_192);
and U6849 (N_6849,N_3000,N_4469);
nand U6850 (N_6850,N_1789,N_2563);
and U6851 (N_6851,N_2600,N_3156);
nor U6852 (N_6852,N_3056,N_1190);
nand U6853 (N_6853,N_3904,N_3642);
or U6854 (N_6854,N_2276,N_2953);
xor U6855 (N_6855,N_653,N_2340);
or U6856 (N_6856,N_3041,N_4535);
nand U6857 (N_6857,N_4845,N_4101);
and U6858 (N_6858,N_4892,N_3613);
nor U6859 (N_6859,N_2483,N_1519);
or U6860 (N_6860,N_3604,N_3430);
nor U6861 (N_6861,N_4593,N_4107);
xnor U6862 (N_6862,N_1173,N_1126);
or U6863 (N_6863,N_2525,N_4890);
xor U6864 (N_6864,N_2742,N_277);
nand U6865 (N_6865,N_1548,N_2087);
and U6866 (N_6866,N_1778,N_1110);
nand U6867 (N_6867,N_2546,N_1935);
nor U6868 (N_6868,N_2916,N_1840);
nor U6869 (N_6869,N_2060,N_2609);
nor U6870 (N_6870,N_3987,N_4155);
or U6871 (N_6871,N_4641,N_3942);
or U6872 (N_6872,N_834,N_2960);
xor U6873 (N_6873,N_3458,N_2498);
xor U6874 (N_6874,N_2035,N_3469);
and U6875 (N_6875,N_1805,N_4487);
and U6876 (N_6876,N_3699,N_912);
nor U6877 (N_6877,N_2284,N_3978);
and U6878 (N_6878,N_1395,N_193);
xor U6879 (N_6879,N_4464,N_4138);
nand U6880 (N_6880,N_3140,N_1084);
nand U6881 (N_6881,N_2690,N_4985);
nor U6882 (N_6882,N_1501,N_4132);
xnor U6883 (N_6883,N_1115,N_4012);
or U6884 (N_6884,N_1522,N_2867);
and U6885 (N_6885,N_1070,N_2368);
and U6886 (N_6886,N_452,N_4857);
xor U6887 (N_6887,N_2107,N_1649);
and U6888 (N_6888,N_2250,N_968);
and U6889 (N_6889,N_4008,N_4634);
or U6890 (N_6890,N_2559,N_1086);
xnor U6891 (N_6891,N_4533,N_2371);
or U6892 (N_6892,N_1739,N_2272);
xor U6893 (N_6893,N_3806,N_2422);
and U6894 (N_6894,N_802,N_4402);
nand U6895 (N_6895,N_4229,N_2210);
or U6896 (N_6896,N_3601,N_1298);
nor U6897 (N_6897,N_2996,N_176);
or U6898 (N_6898,N_2217,N_655);
or U6899 (N_6899,N_3881,N_1847);
xor U6900 (N_6900,N_4817,N_829);
nand U6901 (N_6901,N_3683,N_2610);
xor U6902 (N_6902,N_1670,N_3267);
nor U6903 (N_6903,N_4983,N_2503);
nor U6904 (N_6904,N_3819,N_1846);
nor U6905 (N_6905,N_3926,N_156);
nand U6906 (N_6906,N_738,N_2053);
nor U6907 (N_6907,N_1678,N_224);
xor U6908 (N_6908,N_3450,N_741);
xor U6909 (N_6909,N_4537,N_2603);
xnor U6910 (N_6910,N_3710,N_4796);
xor U6911 (N_6911,N_3838,N_460);
xnor U6912 (N_6912,N_1239,N_3341);
nand U6913 (N_6913,N_2828,N_1584);
and U6914 (N_6914,N_1884,N_3198);
xnor U6915 (N_6915,N_4905,N_1387);
nor U6916 (N_6916,N_2749,N_3944);
or U6917 (N_6917,N_2507,N_2230);
xnor U6918 (N_6918,N_2662,N_2809);
nand U6919 (N_6919,N_2385,N_4430);
nand U6920 (N_6920,N_2436,N_3575);
nand U6921 (N_6921,N_2235,N_416);
and U6922 (N_6922,N_446,N_2653);
and U6923 (N_6923,N_2469,N_1943);
and U6924 (N_6924,N_721,N_2011);
and U6925 (N_6925,N_3964,N_2597);
nor U6926 (N_6926,N_1627,N_2173);
nor U6927 (N_6927,N_2342,N_617);
xor U6928 (N_6928,N_3937,N_3514);
and U6929 (N_6929,N_21,N_162);
nand U6930 (N_6930,N_3404,N_1538);
and U6931 (N_6931,N_2321,N_4554);
xnor U6932 (N_6932,N_48,N_1125);
nand U6933 (N_6933,N_1754,N_2233);
xor U6934 (N_6934,N_4717,N_1875);
and U6935 (N_6935,N_1968,N_3682);
nand U6936 (N_6936,N_337,N_2972);
nor U6937 (N_6937,N_310,N_494);
nand U6938 (N_6938,N_3770,N_3725);
xnor U6939 (N_6939,N_535,N_4733);
xnor U6940 (N_6940,N_2977,N_1827);
nor U6941 (N_6941,N_234,N_2369);
xor U6942 (N_6942,N_1531,N_3902);
xor U6943 (N_6943,N_3541,N_1406);
nor U6944 (N_6944,N_4573,N_1197);
and U6945 (N_6945,N_140,N_722);
nand U6946 (N_6946,N_4671,N_1918);
or U6947 (N_6947,N_4182,N_896);
nor U6948 (N_6948,N_129,N_3119);
and U6949 (N_6949,N_69,N_4482);
and U6950 (N_6950,N_4932,N_2643);
or U6951 (N_6951,N_2883,N_1571);
or U6952 (N_6952,N_4028,N_822);
or U6953 (N_6953,N_671,N_1618);
xnor U6954 (N_6954,N_3244,N_1913);
nor U6955 (N_6955,N_571,N_4701);
xnor U6956 (N_6956,N_94,N_4298);
and U6957 (N_6957,N_1619,N_3274);
or U6958 (N_6958,N_2045,N_4460);
nor U6959 (N_6959,N_2410,N_3290);
and U6960 (N_6960,N_492,N_3510);
nor U6961 (N_6961,N_1514,N_378);
or U6962 (N_6962,N_3415,N_754);
and U6963 (N_6963,N_1231,N_4197);
nor U6964 (N_6964,N_4385,N_313);
nor U6965 (N_6965,N_3845,N_2614);
xor U6966 (N_6966,N_1946,N_4598);
or U6967 (N_6967,N_3674,N_1626);
and U6968 (N_6968,N_4781,N_3656);
or U6969 (N_6969,N_3735,N_3786);
and U6970 (N_6970,N_3039,N_4995);
nand U6971 (N_6971,N_3750,N_940);
and U6972 (N_6972,N_305,N_4346);
xnor U6973 (N_6973,N_3581,N_4862);
nor U6974 (N_6974,N_2080,N_4214);
or U6975 (N_6975,N_1667,N_2678);
or U6976 (N_6976,N_4638,N_3803);
nand U6977 (N_6977,N_4762,N_3607);
nand U6978 (N_6978,N_4552,N_3832);
xnor U6979 (N_6979,N_2396,N_2775);
xnor U6980 (N_6980,N_4318,N_4075);
xnor U6981 (N_6981,N_4555,N_2420);
nand U6982 (N_6982,N_990,N_889);
or U6983 (N_6983,N_2831,N_121);
or U6984 (N_6984,N_2687,N_921);
or U6985 (N_6985,N_566,N_2444);
xnor U6986 (N_6986,N_3574,N_3834);
nand U6987 (N_6987,N_2607,N_570);
nand U6988 (N_6988,N_1236,N_2885);
xor U6989 (N_6989,N_3675,N_2027);
and U6990 (N_6990,N_4753,N_2825);
nor U6991 (N_6991,N_4454,N_4133);
nand U6992 (N_6992,N_4644,N_479);
or U6993 (N_6993,N_4366,N_2170);
nor U6994 (N_6994,N_4424,N_4315);
nor U6995 (N_6995,N_4840,N_2789);
and U6996 (N_6996,N_3028,N_2961);
xnor U6997 (N_6997,N_4860,N_3455);
nand U6998 (N_6998,N_1120,N_379);
nand U6999 (N_6999,N_2697,N_4885);
xor U7000 (N_7000,N_1099,N_1669);
and U7001 (N_7001,N_883,N_2694);
xor U7002 (N_7002,N_1679,N_2083);
or U7003 (N_7003,N_3464,N_629);
nand U7004 (N_7004,N_4824,N_1293);
or U7005 (N_7005,N_4563,N_605);
or U7006 (N_7006,N_1857,N_4876);
nand U7007 (N_7007,N_3825,N_1299);
xnor U7008 (N_7008,N_3232,N_1467);
nor U7009 (N_7009,N_4005,N_1735);
or U7010 (N_7010,N_145,N_3694);
and U7011 (N_7011,N_1654,N_2547);
nand U7012 (N_7012,N_302,N_3871);
and U7013 (N_7013,N_34,N_2852);
nor U7014 (N_7014,N_1001,N_3006);
nand U7015 (N_7015,N_1709,N_2266);
or U7016 (N_7016,N_126,N_4099);
nor U7017 (N_7017,N_1607,N_2691);
or U7018 (N_7018,N_3562,N_3545);
and U7019 (N_7019,N_2213,N_4401);
xor U7020 (N_7020,N_3896,N_2325);
nand U7021 (N_7021,N_4262,N_4988);
xnor U7022 (N_7022,N_4322,N_2763);
or U7023 (N_7023,N_4636,N_4254);
or U7024 (N_7024,N_4848,N_2807);
nand U7025 (N_7025,N_758,N_1277);
and U7026 (N_7026,N_4405,N_4714);
nand U7027 (N_7027,N_1192,N_2146);
nand U7028 (N_7028,N_1057,N_2679);
or U7029 (N_7029,N_27,N_1907);
xnor U7030 (N_7030,N_2999,N_2064);
or U7031 (N_7031,N_3898,N_947);
or U7032 (N_7032,N_202,N_2827);
or U7033 (N_7033,N_1575,N_2720);
or U7034 (N_7034,N_4359,N_4957);
nand U7035 (N_7035,N_4947,N_2020);
nor U7036 (N_7036,N_4972,N_4443);
and U7037 (N_7037,N_2177,N_2069);
nand U7038 (N_7038,N_393,N_3914);
xnor U7039 (N_7039,N_1942,N_4998);
and U7040 (N_7040,N_4672,N_2993);
xnor U7041 (N_7041,N_4130,N_2701);
nand U7042 (N_7042,N_4378,N_273);
nor U7043 (N_7043,N_422,N_4893);
nor U7044 (N_7044,N_847,N_1445);
or U7045 (N_7045,N_786,N_3200);
or U7046 (N_7046,N_1954,N_1381);
xor U7047 (N_7047,N_3570,N_2423);
and U7048 (N_7048,N_4968,N_3737);
or U7049 (N_7049,N_1101,N_1516);
and U7050 (N_7050,N_4866,N_2264);
nand U7051 (N_7051,N_1104,N_263);
nand U7052 (N_7052,N_3305,N_233);
xor U7053 (N_7053,N_4386,N_1992);
or U7054 (N_7054,N_1957,N_2780);
xor U7055 (N_7055,N_1108,N_1313);
or U7056 (N_7056,N_2270,N_2115);
or U7057 (N_7057,N_4070,N_107);
and U7058 (N_7058,N_4542,N_3827);
xor U7059 (N_7059,N_2267,N_4830);
nand U7060 (N_7060,N_4529,N_2328);
or U7061 (N_7061,N_2137,N_1520);
nor U7062 (N_7062,N_772,N_2036);
nor U7063 (N_7063,N_2590,N_1019);
nor U7064 (N_7064,N_3954,N_645);
nand U7065 (N_7065,N_372,N_2150);
nand U7066 (N_7066,N_32,N_3505);
nor U7067 (N_7067,N_3935,N_2848);
nand U7068 (N_7068,N_549,N_3245);
nor U7069 (N_7069,N_3927,N_3306);
nand U7070 (N_7070,N_3352,N_2500);
or U7071 (N_7071,N_4397,N_2254);
xnor U7072 (N_7072,N_4673,N_4528);
xor U7073 (N_7073,N_2699,N_4455);
nand U7074 (N_7074,N_3713,N_3264);
or U7075 (N_7075,N_4675,N_4904);
xnor U7076 (N_7076,N_4579,N_3911);
or U7077 (N_7077,N_3961,N_607);
xnor U7078 (N_7078,N_1449,N_1567);
nor U7079 (N_7079,N_2205,N_3268);
nand U7080 (N_7080,N_16,N_4943);
and U7081 (N_7081,N_4938,N_3621);
and U7082 (N_7082,N_2263,N_1257);
nand U7083 (N_7083,N_2277,N_1783);
xnor U7084 (N_7084,N_3057,N_3391);
nand U7085 (N_7085,N_373,N_3584);
nor U7086 (N_7086,N_3854,N_2110);
xor U7087 (N_7087,N_1078,N_3592);
or U7088 (N_7088,N_3148,N_1887);
nor U7089 (N_7089,N_323,N_1848);
and U7090 (N_7090,N_3517,N_1253);
nand U7091 (N_7091,N_899,N_4032);
nand U7092 (N_7092,N_4624,N_3257);
and U7093 (N_7093,N_138,N_810);
and U7094 (N_7094,N_1318,N_2528);
nand U7095 (N_7095,N_85,N_1928);
and U7096 (N_7096,N_1798,N_430);
nor U7097 (N_7097,N_3207,N_1926);
and U7098 (N_7098,N_3462,N_164);
xor U7099 (N_7099,N_222,N_1017);
and U7100 (N_7100,N_2311,N_4344);
nor U7101 (N_7101,N_3661,N_1740);
nand U7102 (N_7102,N_3248,N_3032);
nand U7103 (N_7103,N_948,N_4546);
nor U7104 (N_7104,N_4557,N_1053);
xor U7105 (N_7105,N_4797,N_2675);
and U7106 (N_7106,N_3128,N_2858);
or U7107 (N_7107,N_4524,N_2405);
xor U7108 (N_7108,N_3065,N_1897);
and U7109 (N_7109,N_2333,N_3720);
nor U7110 (N_7110,N_908,N_485);
or U7111 (N_7111,N_2139,N_1810);
nand U7112 (N_7112,N_3146,N_2458);
and U7113 (N_7113,N_685,N_1867);
nor U7114 (N_7114,N_3888,N_3651);
nor U7115 (N_7115,N_496,N_518);
nor U7116 (N_7116,N_3435,N_2135);
xnor U7117 (N_7117,N_488,N_4498);
and U7118 (N_7118,N_331,N_3153);
nor U7119 (N_7119,N_99,N_4030);
nand U7120 (N_7120,N_1477,N_100);
nor U7121 (N_7121,N_2754,N_2640);
or U7122 (N_7122,N_1359,N_714);
and U7123 (N_7123,N_626,N_355);
and U7124 (N_7124,N_4484,N_2142);
nor U7125 (N_7125,N_4457,N_2920);
and U7126 (N_7126,N_458,N_3718);
and U7127 (N_7127,N_349,N_3227);
and U7128 (N_7128,N_4367,N_1432);
and U7129 (N_7129,N_2471,N_1050);
nand U7130 (N_7130,N_3298,N_4072);
xor U7131 (N_7131,N_1425,N_1900);
xnor U7132 (N_7132,N_2394,N_2566);
or U7133 (N_7133,N_1097,N_1959);
nand U7134 (N_7134,N_4993,N_1603);
or U7135 (N_7135,N_4897,N_1023);
nand U7136 (N_7136,N_3627,N_90);
xnor U7137 (N_7137,N_3688,N_2692);
nand U7138 (N_7138,N_3531,N_3583);
or U7139 (N_7139,N_1165,N_4142);
and U7140 (N_7140,N_4463,N_1158);
xnor U7141 (N_7141,N_2644,N_2855);
nand U7142 (N_7142,N_3747,N_4119);
nand U7143 (N_7143,N_261,N_1505);
or U7144 (N_7144,N_3886,N_2952);
and U7145 (N_7145,N_881,N_2384);
or U7146 (N_7146,N_3997,N_4272);
nand U7147 (N_7147,N_1528,N_3632);
and U7148 (N_7148,N_2421,N_4895);
nor U7149 (N_7149,N_2744,N_1713);
nor U7150 (N_7150,N_2732,N_1167);
nor U7151 (N_7151,N_3145,N_3360);
nand U7152 (N_7152,N_3416,N_4227);
nor U7153 (N_7153,N_4258,N_914);
nor U7154 (N_7154,N_541,N_2338);
nand U7155 (N_7155,N_2956,N_986);
nor U7156 (N_7156,N_1366,N_1437);
and U7157 (N_7157,N_4685,N_3228);
nand U7158 (N_7158,N_3191,N_4980);
xnor U7159 (N_7159,N_198,N_2688);
nand U7160 (N_7160,N_894,N_3288);
nand U7161 (N_7161,N_2160,N_1878);
nor U7162 (N_7162,N_4499,N_4381);
nor U7163 (N_7163,N_3062,N_1181);
nor U7164 (N_7164,N_2611,N_2257);
or U7165 (N_7165,N_3922,N_2349);
and U7166 (N_7166,N_2985,N_1664);
and U7167 (N_7167,N_1329,N_2669);
and U7168 (N_7168,N_1690,N_4055);
or U7169 (N_7169,N_3236,N_3347);
and U7170 (N_7170,N_2055,N_1715);
or U7171 (N_7171,N_3986,N_4742);
xor U7172 (N_7172,N_2847,N_229);
nor U7173 (N_7173,N_1641,N_3824);
xnor U7174 (N_7174,N_445,N_45);
or U7175 (N_7175,N_4395,N_637);
nand U7176 (N_7176,N_531,N_3558);
or U7177 (N_7177,N_4599,N_4763);
nand U7178 (N_7178,N_1479,N_1164);
nand U7179 (N_7179,N_1228,N_3721);
nand U7180 (N_7180,N_1077,N_1260);
nand U7181 (N_7181,N_1028,N_4152);
or U7182 (N_7182,N_1676,N_765);
and U7183 (N_7183,N_1821,N_2472);
and U7184 (N_7184,N_4789,N_1824);
nand U7185 (N_7185,N_4066,N_1663);
or U7186 (N_7186,N_933,N_4056);
nor U7187 (N_7187,N_420,N_1537);
or U7188 (N_7188,N_1562,N_1660);
and U7189 (N_7189,N_2854,N_4740);
and U7190 (N_7190,N_3194,N_1480);
or U7191 (N_7191,N_2449,N_1630);
xnor U7192 (N_7192,N_2312,N_405);
or U7193 (N_7193,N_3745,N_4257);
nand U7194 (N_7194,N_872,N_4291);
or U7195 (N_7195,N_1016,N_3467);
nor U7196 (N_7196,N_4514,N_66);
and U7197 (N_7197,N_2889,N_3894);
nand U7198 (N_7198,N_4444,N_319);
and U7199 (N_7199,N_4256,N_4034);
and U7200 (N_7200,N_2089,N_4793);
xor U7201 (N_7201,N_1040,N_797);
or U7202 (N_7202,N_2324,N_1214);
nor U7203 (N_7203,N_1303,N_792);
and U7204 (N_7204,N_3454,N_2510);
and U7205 (N_7205,N_3351,N_3370);
or U7206 (N_7206,N_4949,N_863);
or U7207 (N_7207,N_3677,N_2253);
or U7208 (N_7208,N_3364,N_71);
or U7209 (N_7209,N_473,N_1243);
xor U7210 (N_7210,N_4987,N_978);
xnor U7211 (N_7211,N_3941,N_1240);
nor U7212 (N_7212,N_2360,N_3425);
nor U7213 (N_7213,N_1106,N_3758);
and U7214 (N_7214,N_2821,N_2221);
nand U7215 (N_7215,N_1691,N_1552);
xor U7216 (N_7216,N_4613,N_392);
nand U7217 (N_7217,N_3733,N_3610);
nand U7218 (N_7218,N_1037,N_1311);
or U7219 (N_7219,N_3321,N_36);
or U7220 (N_7220,N_3476,N_3155);
nand U7221 (N_7221,N_1853,N_1224);
nand U7222 (N_7222,N_3820,N_1361);
xnor U7223 (N_7223,N_4560,N_1845);
nor U7224 (N_7224,N_917,N_748);
or U7225 (N_7225,N_4512,N_2151);
xor U7226 (N_7226,N_82,N_300);
or U7227 (N_7227,N_52,N_3685);
or U7228 (N_7228,N_2228,N_3412);
nor U7229 (N_7229,N_4237,N_2815);
or U7230 (N_7230,N_558,N_2726);
and U7231 (N_7231,N_4160,N_3908);
nor U7232 (N_7232,N_4574,N_4216);
xor U7233 (N_7233,N_3019,N_1604);
or U7234 (N_7234,N_3187,N_2882);
xor U7235 (N_7235,N_2909,N_2012);
and U7236 (N_7236,N_4027,N_2840);
and U7237 (N_7237,N_4568,N_315);
or U7238 (N_7238,N_3930,N_4418);
or U7239 (N_7239,N_4306,N_3529);
xnor U7240 (N_7240,N_688,N_2014);
and U7241 (N_7241,N_246,N_1295);
or U7242 (N_7242,N_972,N_2401);
nand U7243 (N_7243,N_3332,N_4437);
xor U7244 (N_7244,N_2986,N_4435);
nand U7245 (N_7245,N_353,N_1747);
nand U7246 (N_7246,N_1305,N_4913);
nor U7247 (N_7247,N_1526,N_4187);
or U7248 (N_7248,N_1760,N_4912);
xnor U7249 (N_7249,N_2523,N_3569);
nor U7250 (N_7250,N_3473,N_3920);
xnor U7251 (N_7251,N_554,N_2181);
nor U7252 (N_7252,N_861,N_4059);
or U7253 (N_7253,N_995,N_3093);
or U7254 (N_7254,N_2432,N_677);
nand U7255 (N_7255,N_826,N_3667);
nand U7256 (N_7256,N_2526,N_2265);
nor U7257 (N_7257,N_268,N_4775);
nor U7258 (N_7258,N_4416,N_3158);
nor U7259 (N_7259,N_4900,N_4361);
xnor U7260 (N_7260,N_527,N_936);
and U7261 (N_7261,N_1018,N_360);
xor U7262 (N_7262,N_3534,N_3655);
or U7263 (N_7263,N_1517,N_3812);
nand U7264 (N_7264,N_4170,N_1061);
xor U7265 (N_7265,N_2897,N_86);
nand U7266 (N_7266,N_2344,N_4954);
xnor U7267 (N_7267,N_4394,N_1751);
nand U7268 (N_7268,N_1737,N_214);
nor U7269 (N_7269,N_1917,N_96);
nor U7270 (N_7270,N_1938,N_2585);
or U7271 (N_7271,N_4131,N_2797);
xor U7272 (N_7272,N_3726,N_4189);
xor U7273 (N_7273,N_2497,N_1640);
and U7274 (N_7274,N_1402,N_44);
nor U7275 (N_7275,N_3701,N_3795);
or U7276 (N_7276,N_3362,N_3421);
xor U7277 (N_7277,N_3938,N_2459);
or U7278 (N_7278,N_4725,N_1041);
nand U7279 (N_7279,N_1949,N_3411);
xor U7280 (N_7280,N_2417,N_4333);
nor U7281 (N_7281,N_2102,N_4545);
nand U7282 (N_7282,N_3494,N_3525);
nor U7283 (N_7283,N_293,N_3005);
or U7284 (N_7284,N_186,N_681);
and U7285 (N_7285,N_4760,N_2948);
nor U7286 (N_7286,N_4350,N_4033);
nor U7287 (N_7287,N_965,N_3296);
xor U7288 (N_7288,N_1267,N_1559);
nand U7289 (N_7289,N_1605,N_4637);
and U7290 (N_7290,N_1223,N_295);
nor U7291 (N_7291,N_2719,N_3121);
nor U7292 (N_7292,N_4166,N_3676);
and U7293 (N_7293,N_334,N_1872);
nor U7294 (N_7294,N_4608,N_913);
nand U7295 (N_7295,N_4823,N_4441);
nor U7296 (N_7296,N_4562,N_3080);
nor U7297 (N_7297,N_1549,N_342);
xnor U7298 (N_7298,N_1021,N_3749);
nand U7299 (N_7299,N_4887,N_3740);
or U7300 (N_7300,N_2431,N_1863);
xnor U7301 (N_7301,N_3947,N_1058);
or U7302 (N_7302,N_2332,N_634);
and U7303 (N_7303,N_4199,N_1160);
and U7304 (N_7304,N_2416,N_4518);
xor U7305 (N_7305,N_1828,N_979);
nor U7306 (N_7306,N_2531,N_1725);
nor U7307 (N_7307,N_1079,N_3174);
and U7308 (N_7308,N_4697,N_3772);
or U7309 (N_7309,N_1895,N_595);
nand U7310 (N_7310,N_3299,N_1860);
nand U7311 (N_7311,N_2695,N_2347);
xnor U7312 (N_7312,N_4712,N_4744);
xor U7313 (N_7313,N_3396,N_3018);
nand U7314 (N_7314,N_1653,N_4651);
xor U7315 (N_7315,N_4285,N_4918);
nor U7316 (N_7316,N_3184,N_4846);
xor U7317 (N_7317,N_1964,N_667);
xor U7318 (N_7318,N_4260,N_137);
or U7319 (N_7319,N_4159,N_4761);
nor U7320 (N_7320,N_4534,N_2352);
or U7321 (N_7321,N_3503,N_469);
xor U7322 (N_7322,N_3722,N_4210);
nand U7323 (N_7323,N_1748,N_4352);
nor U7324 (N_7324,N_3007,N_1100);
xnor U7325 (N_7325,N_4338,N_3339);
or U7326 (N_7326,N_236,N_4234);
xnor U7327 (N_7327,N_98,N_1989);
nand U7328 (N_7328,N_4594,N_4536);
xnor U7329 (N_7329,N_2079,N_3102);
nor U7330 (N_7330,N_2346,N_3560);
xnor U7331 (N_7331,N_2435,N_397);
or U7332 (N_7332,N_1343,N_1363);
or U7333 (N_7333,N_427,N_2658);
nand U7334 (N_7334,N_2178,N_3635);
and U7335 (N_7335,N_984,N_701);
or U7336 (N_7336,N_3636,N_2145);
nand U7337 (N_7337,N_4052,N_1062);
and U7338 (N_7338,N_2269,N_2323);
nand U7339 (N_7339,N_1762,N_2641);
and U7340 (N_7340,N_3129,N_3742);
nor U7341 (N_7341,N_3630,N_1454);
nand U7342 (N_7342,N_2991,N_1529);
xnor U7343 (N_7343,N_2316,N_4805);
nor U7344 (N_7344,N_2771,N_3724);
or U7345 (N_7345,N_3840,N_3081);
xnor U7346 (N_7346,N_1290,N_2404);
or U7347 (N_7347,N_4567,N_4766);
and U7348 (N_7348,N_2514,N_3493);
or U7349 (N_7349,N_4330,N_926);
xnor U7350 (N_7350,N_1711,N_514);
or U7351 (N_7351,N_4576,N_303);
nand U7352 (N_7352,N_2703,N_726);
nand U7353 (N_7353,N_1898,N_4679);
or U7354 (N_7354,N_665,N_1622);
or U7355 (N_7355,N_612,N_759);
nand U7356 (N_7356,N_2660,N_4864);
nand U7357 (N_7357,N_762,N_783);
and U7358 (N_7358,N_4861,N_3572);
and U7359 (N_7359,N_2670,N_2710);
nor U7360 (N_7360,N_1458,N_4125);
nor U7361 (N_7361,N_3216,N_4873);
nand U7362 (N_7362,N_2946,N_2319);
xnor U7363 (N_7363,N_1487,N_2530);
or U7364 (N_7364,N_2887,N_2877);
xor U7365 (N_7365,N_4247,N_814);
or U7366 (N_7366,N_4837,N_2197);
nand U7367 (N_7367,N_592,N_2793);
and U7368 (N_7368,N_2185,N_1396);
nor U7369 (N_7369,N_2464,N_1624);
xor U7370 (N_7370,N_3014,N_1154);
or U7371 (N_7371,N_4959,N_2372);
and U7372 (N_7372,N_3027,N_1758);
xnor U7373 (N_7373,N_1060,N_2683);
xor U7374 (N_7374,N_3622,N_4933);
or U7375 (N_7375,N_1841,N_1457);
and U7376 (N_7376,N_2259,N_1489);
or U7377 (N_7377,N_4811,N_4403);
nand U7378 (N_7378,N_2638,N_2860);
xor U7379 (N_7379,N_3781,N_641);
nand U7380 (N_7380,N_454,N_909);
nand U7381 (N_7381,N_4200,N_316);
or U7382 (N_7382,N_2034,N_2451);
and U7383 (N_7383,N_1974,N_2108);
nor U7384 (N_7384,N_587,N_2587);
nor U7385 (N_7385,N_1315,N_207);
nand U7386 (N_7386,N_727,N_4472);
and U7387 (N_7387,N_4521,N_1685);
and U7388 (N_7388,N_851,N_4757);
nand U7389 (N_7389,N_4407,N_2429);
nand U7390 (N_7390,N_1724,N_3996);
or U7391 (N_7391,N_3540,N_4867);
xnor U7392 (N_7392,N_2894,N_4686);
and U7393 (N_7393,N_2105,N_3934);
xor U7394 (N_7394,N_41,N_3821);
or U7395 (N_7395,N_1969,N_4620);
or U7396 (N_7396,N_1168,N_1316);
nand U7397 (N_7397,N_1145,N_596);
and U7398 (N_7398,N_4720,N_3691);
nand U7399 (N_7399,N_2203,N_1453);
nand U7400 (N_7400,N_1289,N_4703);
or U7401 (N_7401,N_613,N_1844);
xnor U7402 (N_7402,N_4841,N_1852);
nand U7403 (N_7403,N_999,N_1553);
nor U7404 (N_7404,N_3313,N_4171);
and U7405 (N_7405,N_856,N_180);
nand U7406 (N_7406,N_1582,N_4815);
nor U7407 (N_7407,N_1091,N_563);
nor U7408 (N_7408,N_1683,N_1997);
or U7409 (N_7409,N_4975,N_1049);
or U7410 (N_7410,N_2434,N_3143);
and U7411 (N_7411,N_1279,N_695);
or U7412 (N_7412,N_3868,N_369);
or U7413 (N_7413,N_616,N_3098);
xnor U7414 (N_7414,N_3703,N_1682);
xnor U7415 (N_7415,N_4283,N_2169);
and U7416 (N_7416,N_4302,N_1259);
xnor U7417 (N_7417,N_3301,N_2676);
or U7418 (N_7418,N_4137,N_2386);
xor U7419 (N_7419,N_4950,N_1421);
and U7420 (N_7420,N_3361,N_2994);
or U7421 (N_7421,N_160,N_2512);
or U7422 (N_7422,N_2938,N_1463);
xor U7423 (N_7423,N_15,N_364);
nor U7424 (N_7424,N_4293,N_2482);
and U7425 (N_7425,N_929,N_2399);
or U7426 (N_7426,N_2545,N_3286);
and U7427 (N_7427,N_29,N_4511);
xor U7428 (N_7428,N_4006,N_4021);
and U7429 (N_7429,N_2787,N_1784);
and U7430 (N_7430,N_2524,N_4719);
xnor U7431 (N_7431,N_4141,N_3595);
nor U7432 (N_7432,N_2123,N_3515);
nor U7433 (N_7433,N_4010,N_400);
nand U7434 (N_7434,N_1201,N_3043);
or U7435 (N_7435,N_1248,N_2397);
and U7436 (N_7436,N_891,N_3793);
nand U7437 (N_7437,N_3420,N_585);
nand U7438 (N_7438,N_877,N_3220);
xor U7439 (N_7439,N_2806,N_2121);
nor U7440 (N_7440,N_1523,N_4540);
xor U7441 (N_7441,N_1956,N_551);
nand U7442 (N_7442,N_1775,N_3511);
nor U7443 (N_7443,N_4692,N_1838);
and U7444 (N_7444,N_159,N_3879);
and U7445 (N_7445,N_2534,N_2602);
or U7446 (N_7446,N_3335,N_799);
or U7447 (N_7447,N_1712,N_1766);
xnor U7448 (N_7448,N_4994,N_163);
xnor U7449 (N_7449,N_1157,N_2286);
nor U7450 (N_7450,N_2802,N_546);
and U7451 (N_7451,N_1064,N_717);
nand U7452 (N_7452,N_3631,N_2206);
nor U7453 (N_7453,N_4439,N_560);
nand U7454 (N_7454,N_3419,N_855);
or U7455 (N_7455,N_981,N_4301);
xor U7456 (N_7456,N_1540,N_1309);
xnor U7457 (N_7457,N_1153,N_689);
xnor U7458 (N_7458,N_1178,N_2302);
and U7459 (N_7459,N_1475,N_3999);
nor U7460 (N_7460,N_4572,N_1036);
and U7461 (N_7461,N_1832,N_747);
xnor U7462 (N_7462,N_447,N_2075);
or U7463 (N_7463,N_530,N_2659);
or U7464 (N_7464,N_2748,N_510);
xor U7465 (N_7465,N_630,N_753);
nand U7466 (N_7466,N_4238,N_3250);
nand U7467 (N_7467,N_3637,N_4243);
and U7468 (N_7468,N_3668,N_1136);
and U7469 (N_7469,N_942,N_3993);
and U7470 (N_7470,N_3965,N_928);
or U7471 (N_7471,N_4706,N_960);
nand U7472 (N_7472,N_1105,N_4026);
xnor U7473 (N_7473,N_1430,N_4218);
xnor U7474 (N_7474,N_256,N_2030);
and U7475 (N_7475,N_4944,N_3587);
nand U7476 (N_7476,N_4064,N_2522);
xnor U7477 (N_7477,N_2757,N_3680);
xnor U7478 (N_7478,N_1836,N_544);
xnor U7479 (N_7479,N_332,N_3779);
xnor U7480 (N_7480,N_4311,N_3785);
and U7481 (N_7481,N_4974,N_57);
or U7482 (N_7482,N_2505,N_3271);
or U7483 (N_7483,N_4631,N_4415);
nor U7484 (N_7484,N_3580,N_1924);
nand U7485 (N_7485,N_572,N_1137);
and U7486 (N_7486,N_1806,N_1133);
and U7487 (N_7487,N_3342,N_3760);
xnor U7488 (N_7488,N_1183,N_1776);
nor U7489 (N_7489,N_3882,N_4239);
and U7490 (N_7490,N_2147,N_3149);
nand U7491 (N_7491,N_3952,N_1911);
nor U7492 (N_7492,N_1007,N_4603);
and U7493 (N_7493,N_289,N_2445);
nand U7494 (N_7494,N_161,N_2301);
or U7495 (N_7495,N_3985,N_1444);
or U7496 (N_7496,N_3084,N_3219);
xnor U7497 (N_7497,N_2973,N_2167);
nor U7498 (N_7498,N_141,N_4183);
and U7499 (N_7499,N_4139,N_4110);
and U7500 (N_7500,N_3427,N_2080);
xor U7501 (N_7501,N_3882,N_4475);
and U7502 (N_7502,N_1674,N_2887);
or U7503 (N_7503,N_4391,N_2752);
nor U7504 (N_7504,N_2786,N_3604);
nor U7505 (N_7505,N_4714,N_126);
nand U7506 (N_7506,N_3093,N_3110);
or U7507 (N_7507,N_2785,N_2493);
and U7508 (N_7508,N_4664,N_2897);
or U7509 (N_7509,N_4158,N_4951);
or U7510 (N_7510,N_1445,N_4202);
nand U7511 (N_7511,N_3177,N_3016);
nand U7512 (N_7512,N_631,N_444);
xor U7513 (N_7513,N_410,N_4258);
xnor U7514 (N_7514,N_2515,N_4976);
or U7515 (N_7515,N_4803,N_2198);
and U7516 (N_7516,N_2168,N_2667);
xnor U7517 (N_7517,N_2412,N_2204);
and U7518 (N_7518,N_1755,N_2373);
nor U7519 (N_7519,N_2037,N_781);
nand U7520 (N_7520,N_2367,N_1056);
nand U7521 (N_7521,N_2414,N_3485);
nor U7522 (N_7522,N_3224,N_4209);
nand U7523 (N_7523,N_348,N_2115);
or U7524 (N_7524,N_1393,N_792);
and U7525 (N_7525,N_222,N_326);
nor U7526 (N_7526,N_4670,N_897);
or U7527 (N_7527,N_1468,N_2790);
or U7528 (N_7528,N_2079,N_346);
nor U7529 (N_7529,N_707,N_3376);
or U7530 (N_7530,N_4874,N_3102);
nor U7531 (N_7531,N_3168,N_2691);
nand U7532 (N_7532,N_1431,N_2249);
or U7533 (N_7533,N_1277,N_550);
nand U7534 (N_7534,N_3789,N_147);
or U7535 (N_7535,N_147,N_1576);
nand U7536 (N_7536,N_4694,N_4592);
nor U7537 (N_7537,N_1258,N_2420);
nor U7538 (N_7538,N_2733,N_2621);
and U7539 (N_7539,N_3334,N_3012);
nor U7540 (N_7540,N_2673,N_2699);
and U7541 (N_7541,N_1055,N_4755);
and U7542 (N_7542,N_1843,N_3982);
nor U7543 (N_7543,N_4776,N_2134);
and U7544 (N_7544,N_508,N_3719);
nor U7545 (N_7545,N_1303,N_2032);
xor U7546 (N_7546,N_545,N_2250);
and U7547 (N_7547,N_283,N_1086);
xnor U7548 (N_7548,N_3633,N_2476);
and U7549 (N_7549,N_4446,N_4255);
nand U7550 (N_7550,N_1172,N_1684);
nand U7551 (N_7551,N_76,N_3791);
xnor U7552 (N_7552,N_2840,N_4794);
or U7553 (N_7553,N_3340,N_413);
or U7554 (N_7554,N_2537,N_4399);
xor U7555 (N_7555,N_2390,N_3714);
and U7556 (N_7556,N_2651,N_1861);
or U7557 (N_7557,N_2157,N_4136);
xnor U7558 (N_7558,N_4143,N_3445);
nor U7559 (N_7559,N_1685,N_4809);
xnor U7560 (N_7560,N_4821,N_3764);
nand U7561 (N_7561,N_4038,N_578);
and U7562 (N_7562,N_2554,N_3394);
or U7563 (N_7563,N_2042,N_14);
xor U7564 (N_7564,N_4191,N_2751);
xor U7565 (N_7565,N_4052,N_1969);
or U7566 (N_7566,N_3240,N_3348);
nor U7567 (N_7567,N_2514,N_4702);
and U7568 (N_7568,N_993,N_3890);
and U7569 (N_7569,N_4183,N_2948);
or U7570 (N_7570,N_2186,N_878);
xor U7571 (N_7571,N_1787,N_206);
and U7572 (N_7572,N_446,N_1272);
xnor U7573 (N_7573,N_2451,N_2109);
and U7574 (N_7574,N_3812,N_2340);
nor U7575 (N_7575,N_4067,N_683);
nand U7576 (N_7576,N_4533,N_703);
nand U7577 (N_7577,N_1912,N_4228);
and U7578 (N_7578,N_3884,N_2296);
xor U7579 (N_7579,N_2290,N_3374);
nor U7580 (N_7580,N_1583,N_3979);
or U7581 (N_7581,N_3591,N_4819);
nor U7582 (N_7582,N_4850,N_2086);
or U7583 (N_7583,N_1073,N_1134);
nor U7584 (N_7584,N_3054,N_3596);
nand U7585 (N_7585,N_857,N_3001);
nor U7586 (N_7586,N_766,N_3411);
or U7587 (N_7587,N_2475,N_4641);
xor U7588 (N_7588,N_2070,N_3081);
and U7589 (N_7589,N_671,N_2822);
nor U7590 (N_7590,N_4117,N_2471);
xnor U7591 (N_7591,N_2665,N_2733);
or U7592 (N_7592,N_3021,N_125);
nand U7593 (N_7593,N_2413,N_856);
nand U7594 (N_7594,N_4695,N_3913);
xnor U7595 (N_7595,N_3399,N_2048);
or U7596 (N_7596,N_2283,N_2424);
and U7597 (N_7597,N_2978,N_469);
nand U7598 (N_7598,N_3273,N_4113);
or U7599 (N_7599,N_437,N_4043);
or U7600 (N_7600,N_3514,N_154);
nand U7601 (N_7601,N_2837,N_583);
xnor U7602 (N_7602,N_944,N_2733);
nand U7603 (N_7603,N_787,N_4316);
nor U7604 (N_7604,N_4570,N_118);
xnor U7605 (N_7605,N_62,N_1635);
nor U7606 (N_7606,N_4886,N_2692);
nor U7607 (N_7607,N_2926,N_1839);
and U7608 (N_7608,N_1638,N_4946);
and U7609 (N_7609,N_3466,N_4331);
and U7610 (N_7610,N_1414,N_3110);
or U7611 (N_7611,N_4659,N_98);
xnor U7612 (N_7612,N_2626,N_508);
and U7613 (N_7613,N_1993,N_2941);
nor U7614 (N_7614,N_4487,N_715);
xnor U7615 (N_7615,N_3934,N_4705);
nand U7616 (N_7616,N_3436,N_3907);
xor U7617 (N_7617,N_2831,N_3289);
xnor U7618 (N_7618,N_1099,N_1823);
nand U7619 (N_7619,N_4690,N_512);
xor U7620 (N_7620,N_872,N_1573);
nand U7621 (N_7621,N_2760,N_1441);
xnor U7622 (N_7622,N_3366,N_3012);
nand U7623 (N_7623,N_3629,N_405);
nand U7624 (N_7624,N_3543,N_4753);
nand U7625 (N_7625,N_3246,N_2908);
and U7626 (N_7626,N_4548,N_4596);
or U7627 (N_7627,N_3336,N_243);
or U7628 (N_7628,N_4565,N_622);
nand U7629 (N_7629,N_67,N_4105);
nor U7630 (N_7630,N_2047,N_4763);
xor U7631 (N_7631,N_3740,N_1283);
and U7632 (N_7632,N_865,N_2192);
or U7633 (N_7633,N_137,N_1250);
or U7634 (N_7634,N_3475,N_2681);
xor U7635 (N_7635,N_3217,N_2799);
nor U7636 (N_7636,N_1871,N_336);
xor U7637 (N_7637,N_2636,N_3497);
xnor U7638 (N_7638,N_2769,N_2969);
nor U7639 (N_7639,N_1629,N_4152);
and U7640 (N_7640,N_1774,N_1090);
or U7641 (N_7641,N_670,N_3552);
xnor U7642 (N_7642,N_1206,N_1928);
nor U7643 (N_7643,N_2718,N_1991);
or U7644 (N_7644,N_2268,N_1209);
nor U7645 (N_7645,N_3202,N_1551);
nor U7646 (N_7646,N_4792,N_3823);
xor U7647 (N_7647,N_2212,N_3857);
xnor U7648 (N_7648,N_3575,N_92);
or U7649 (N_7649,N_1216,N_1786);
and U7650 (N_7650,N_3353,N_3620);
xor U7651 (N_7651,N_2104,N_1352);
or U7652 (N_7652,N_693,N_3062);
and U7653 (N_7653,N_1692,N_1815);
nand U7654 (N_7654,N_3083,N_4177);
or U7655 (N_7655,N_445,N_645);
xnor U7656 (N_7656,N_3459,N_750);
nand U7657 (N_7657,N_3984,N_3517);
nand U7658 (N_7658,N_3093,N_3510);
nand U7659 (N_7659,N_3019,N_2834);
or U7660 (N_7660,N_979,N_2328);
or U7661 (N_7661,N_1985,N_3361);
or U7662 (N_7662,N_3049,N_1806);
nand U7663 (N_7663,N_297,N_3111);
nand U7664 (N_7664,N_3751,N_3071);
and U7665 (N_7665,N_3483,N_800);
xor U7666 (N_7666,N_1093,N_2885);
and U7667 (N_7667,N_3956,N_2311);
xor U7668 (N_7668,N_4209,N_4956);
nand U7669 (N_7669,N_1300,N_3525);
nor U7670 (N_7670,N_1488,N_921);
nor U7671 (N_7671,N_3805,N_2318);
and U7672 (N_7672,N_870,N_3688);
nor U7673 (N_7673,N_3407,N_653);
xor U7674 (N_7674,N_1908,N_287);
xor U7675 (N_7675,N_982,N_2810);
or U7676 (N_7676,N_4946,N_2186);
or U7677 (N_7677,N_2442,N_3077);
xnor U7678 (N_7678,N_1503,N_2391);
or U7679 (N_7679,N_456,N_2353);
nor U7680 (N_7680,N_1626,N_3716);
nor U7681 (N_7681,N_2140,N_3481);
nand U7682 (N_7682,N_2711,N_1789);
nand U7683 (N_7683,N_4809,N_3241);
nor U7684 (N_7684,N_40,N_4742);
nor U7685 (N_7685,N_4466,N_4765);
and U7686 (N_7686,N_932,N_810);
or U7687 (N_7687,N_3774,N_2847);
nand U7688 (N_7688,N_2860,N_442);
xor U7689 (N_7689,N_2715,N_252);
xnor U7690 (N_7690,N_4704,N_1431);
xnor U7691 (N_7691,N_391,N_4309);
and U7692 (N_7692,N_3796,N_4665);
or U7693 (N_7693,N_4669,N_2937);
or U7694 (N_7694,N_3573,N_26);
nand U7695 (N_7695,N_3976,N_2641);
nor U7696 (N_7696,N_2576,N_212);
nand U7697 (N_7697,N_2298,N_4140);
xnor U7698 (N_7698,N_4651,N_3740);
xor U7699 (N_7699,N_302,N_992);
xnor U7700 (N_7700,N_3029,N_2184);
nand U7701 (N_7701,N_2746,N_1802);
and U7702 (N_7702,N_1,N_995);
nor U7703 (N_7703,N_1731,N_2089);
and U7704 (N_7704,N_4906,N_3525);
and U7705 (N_7705,N_3107,N_4061);
nor U7706 (N_7706,N_270,N_1546);
or U7707 (N_7707,N_2323,N_3978);
xor U7708 (N_7708,N_4441,N_3500);
or U7709 (N_7709,N_1392,N_2229);
nor U7710 (N_7710,N_344,N_4744);
nor U7711 (N_7711,N_3983,N_3372);
xor U7712 (N_7712,N_785,N_1028);
nor U7713 (N_7713,N_3142,N_4315);
nand U7714 (N_7714,N_2091,N_1266);
xor U7715 (N_7715,N_4882,N_2766);
or U7716 (N_7716,N_2809,N_214);
nor U7717 (N_7717,N_2078,N_2573);
xnor U7718 (N_7718,N_4527,N_2068);
xnor U7719 (N_7719,N_1972,N_1530);
nor U7720 (N_7720,N_4798,N_1744);
nor U7721 (N_7721,N_222,N_3473);
or U7722 (N_7722,N_455,N_70);
nand U7723 (N_7723,N_3415,N_3004);
or U7724 (N_7724,N_3474,N_2223);
or U7725 (N_7725,N_4860,N_1622);
xor U7726 (N_7726,N_4518,N_930);
nand U7727 (N_7727,N_949,N_2679);
nand U7728 (N_7728,N_4294,N_64);
and U7729 (N_7729,N_1283,N_3949);
xor U7730 (N_7730,N_4120,N_1201);
and U7731 (N_7731,N_4486,N_175);
or U7732 (N_7732,N_4793,N_4374);
xor U7733 (N_7733,N_1838,N_1977);
nand U7734 (N_7734,N_2630,N_4977);
nor U7735 (N_7735,N_4864,N_4210);
xnor U7736 (N_7736,N_2056,N_4290);
nor U7737 (N_7737,N_399,N_273);
xnor U7738 (N_7738,N_4456,N_889);
xor U7739 (N_7739,N_2382,N_4374);
nand U7740 (N_7740,N_3068,N_479);
nand U7741 (N_7741,N_1482,N_3186);
nand U7742 (N_7742,N_1311,N_3698);
nor U7743 (N_7743,N_1589,N_268);
nand U7744 (N_7744,N_3830,N_3833);
or U7745 (N_7745,N_2138,N_4710);
and U7746 (N_7746,N_4762,N_2343);
nand U7747 (N_7747,N_640,N_1597);
nor U7748 (N_7748,N_2288,N_51);
and U7749 (N_7749,N_1994,N_2421);
nor U7750 (N_7750,N_3978,N_3680);
nand U7751 (N_7751,N_1687,N_3853);
or U7752 (N_7752,N_4777,N_2307);
and U7753 (N_7753,N_4397,N_2491);
nor U7754 (N_7754,N_2416,N_3868);
nand U7755 (N_7755,N_278,N_129);
or U7756 (N_7756,N_2801,N_3271);
nor U7757 (N_7757,N_941,N_3626);
or U7758 (N_7758,N_279,N_3864);
nand U7759 (N_7759,N_3450,N_4618);
nand U7760 (N_7760,N_2125,N_3032);
xor U7761 (N_7761,N_4101,N_4067);
or U7762 (N_7762,N_2526,N_3744);
and U7763 (N_7763,N_4156,N_2257);
or U7764 (N_7764,N_1263,N_2005);
nor U7765 (N_7765,N_1981,N_2330);
nor U7766 (N_7766,N_2306,N_4791);
nor U7767 (N_7767,N_1292,N_3620);
and U7768 (N_7768,N_2867,N_1896);
xnor U7769 (N_7769,N_1295,N_1877);
and U7770 (N_7770,N_1252,N_4237);
nor U7771 (N_7771,N_2697,N_993);
xnor U7772 (N_7772,N_1590,N_1910);
xor U7773 (N_7773,N_485,N_4712);
nand U7774 (N_7774,N_3305,N_2880);
nor U7775 (N_7775,N_85,N_1355);
and U7776 (N_7776,N_3942,N_66);
nor U7777 (N_7777,N_2409,N_2899);
nor U7778 (N_7778,N_736,N_702);
xnor U7779 (N_7779,N_3841,N_4782);
nor U7780 (N_7780,N_1459,N_3907);
nand U7781 (N_7781,N_4589,N_2911);
and U7782 (N_7782,N_887,N_3062);
xor U7783 (N_7783,N_4468,N_1480);
nor U7784 (N_7784,N_3409,N_2938);
and U7785 (N_7785,N_3541,N_4464);
nand U7786 (N_7786,N_150,N_1034);
or U7787 (N_7787,N_2105,N_3623);
nor U7788 (N_7788,N_2828,N_4877);
and U7789 (N_7789,N_3748,N_4548);
xnor U7790 (N_7790,N_2828,N_2001);
nor U7791 (N_7791,N_2358,N_1249);
or U7792 (N_7792,N_2728,N_4495);
nand U7793 (N_7793,N_1723,N_2898);
nand U7794 (N_7794,N_2259,N_4801);
nor U7795 (N_7795,N_4909,N_245);
nand U7796 (N_7796,N_4774,N_2203);
nor U7797 (N_7797,N_4713,N_4463);
xnor U7798 (N_7798,N_1800,N_462);
nand U7799 (N_7799,N_4333,N_3447);
or U7800 (N_7800,N_1165,N_2415);
xor U7801 (N_7801,N_187,N_277);
xor U7802 (N_7802,N_821,N_181);
or U7803 (N_7803,N_770,N_4294);
or U7804 (N_7804,N_78,N_4064);
xnor U7805 (N_7805,N_645,N_17);
xor U7806 (N_7806,N_2854,N_1211);
and U7807 (N_7807,N_741,N_2204);
nor U7808 (N_7808,N_3947,N_558);
nand U7809 (N_7809,N_1702,N_3913);
or U7810 (N_7810,N_224,N_4680);
nand U7811 (N_7811,N_1706,N_3794);
xor U7812 (N_7812,N_3063,N_206);
or U7813 (N_7813,N_2681,N_1453);
or U7814 (N_7814,N_3763,N_3532);
nand U7815 (N_7815,N_913,N_3982);
and U7816 (N_7816,N_1464,N_1244);
nand U7817 (N_7817,N_3309,N_2103);
or U7818 (N_7818,N_2010,N_2365);
nand U7819 (N_7819,N_4666,N_4588);
xnor U7820 (N_7820,N_249,N_3450);
and U7821 (N_7821,N_1323,N_914);
or U7822 (N_7822,N_3072,N_3588);
nor U7823 (N_7823,N_2672,N_3322);
xor U7824 (N_7824,N_2341,N_4298);
or U7825 (N_7825,N_1590,N_807);
nor U7826 (N_7826,N_4055,N_1883);
and U7827 (N_7827,N_3515,N_1322);
xor U7828 (N_7828,N_3793,N_443);
xnor U7829 (N_7829,N_1625,N_2172);
xor U7830 (N_7830,N_3377,N_3821);
or U7831 (N_7831,N_640,N_242);
xor U7832 (N_7832,N_2009,N_2065);
and U7833 (N_7833,N_2742,N_454);
or U7834 (N_7834,N_1871,N_3514);
or U7835 (N_7835,N_3429,N_3978);
and U7836 (N_7836,N_1532,N_1633);
nor U7837 (N_7837,N_34,N_750);
xnor U7838 (N_7838,N_2598,N_597);
nor U7839 (N_7839,N_555,N_2884);
nand U7840 (N_7840,N_4317,N_4767);
nand U7841 (N_7841,N_1577,N_4046);
nor U7842 (N_7842,N_3381,N_2305);
xnor U7843 (N_7843,N_3933,N_2895);
nand U7844 (N_7844,N_1720,N_1719);
or U7845 (N_7845,N_3339,N_4538);
nor U7846 (N_7846,N_570,N_2573);
nand U7847 (N_7847,N_4664,N_3921);
nand U7848 (N_7848,N_1475,N_3331);
xor U7849 (N_7849,N_2150,N_2604);
and U7850 (N_7850,N_2161,N_860);
or U7851 (N_7851,N_3161,N_4879);
xnor U7852 (N_7852,N_59,N_1101);
nand U7853 (N_7853,N_3469,N_4239);
nand U7854 (N_7854,N_3755,N_2879);
nand U7855 (N_7855,N_3769,N_1170);
xor U7856 (N_7856,N_3505,N_3190);
xor U7857 (N_7857,N_3077,N_2360);
nand U7858 (N_7858,N_341,N_3582);
and U7859 (N_7859,N_2553,N_4188);
or U7860 (N_7860,N_1938,N_3938);
nor U7861 (N_7861,N_3347,N_4659);
nand U7862 (N_7862,N_4094,N_3108);
nor U7863 (N_7863,N_2658,N_4474);
nand U7864 (N_7864,N_751,N_1773);
nor U7865 (N_7865,N_231,N_3928);
nor U7866 (N_7866,N_1049,N_1526);
nor U7867 (N_7867,N_4304,N_3275);
nor U7868 (N_7868,N_4694,N_4570);
nor U7869 (N_7869,N_1322,N_771);
or U7870 (N_7870,N_3835,N_2355);
and U7871 (N_7871,N_2239,N_4919);
nand U7872 (N_7872,N_1474,N_2542);
nor U7873 (N_7873,N_1813,N_3949);
nand U7874 (N_7874,N_1781,N_4518);
nand U7875 (N_7875,N_342,N_23);
and U7876 (N_7876,N_3511,N_2224);
nand U7877 (N_7877,N_2553,N_1565);
nor U7878 (N_7878,N_4583,N_1241);
xor U7879 (N_7879,N_2288,N_910);
nand U7880 (N_7880,N_2483,N_4517);
or U7881 (N_7881,N_470,N_3177);
or U7882 (N_7882,N_2629,N_1891);
or U7883 (N_7883,N_789,N_4669);
nor U7884 (N_7884,N_2329,N_1284);
nor U7885 (N_7885,N_4215,N_2191);
xor U7886 (N_7886,N_412,N_4947);
or U7887 (N_7887,N_2289,N_2110);
and U7888 (N_7888,N_1709,N_1087);
nand U7889 (N_7889,N_1323,N_3252);
or U7890 (N_7890,N_3015,N_1200);
and U7891 (N_7891,N_2726,N_4716);
nor U7892 (N_7892,N_4393,N_3707);
and U7893 (N_7893,N_3665,N_673);
or U7894 (N_7894,N_3722,N_574);
or U7895 (N_7895,N_2477,N_1415);
and U7896 (N_7896,N_2323,N_717);
nand U7897 (N_7897,N_2475,N_1722);
xnor U7898 (N_7898,N_3594,N_4069);
nand U7899 (N_7899,N_2256,N_2106);
xnor U7900 (N_7900,N_1336,N_1296);
and U7901 (N_7901,N_3389,N_1357);
nor U7902 (N_7902,N_1231,N_3532);
and U7903 (N_7903,N_4882,N_1111);
or U7904 (N_7904,N_4828,N_2941);
xnor U7905 (N_7905,N_1220,N_1137);
xor U7906 (N_7906,N_613,N_2086);
nor U7907 (N_7907,N_3614,N_3032);
nor U7908 (N_7908,N_1149,N_1384);
or U7909 (N_7909,N_2480,N_3071);
nand U7910 (N_7910,N_2198,N_1112);
xnor U7911 (N_7911,N_3002,N_630);
or U7912 (N_7912,N_1206,N_1613);
nand U7913 (N_7913,N_3277,N_2570);
and U7914 (N_7914,N_2319,N_3204);
nand U7915 (N_7915,N_3294,N_618);
xnor U7916 (N_7916,N_1549,N_4285);
nor U7917 (N_7917,N_3829,N_4273);
and U7918 (N_7918,N_2186,N_3295);
and U7919 (N_7919,N_1049,N_3567);
nor U7920 (N_7920,N_1409,N_2411);
xnor U7921 (N_7921,N_1619,N_455);
or U7922 (N_7922,N_4754,N_1825);
or U7923 (N_7923,N_4194,N_541);
nand U7924 (N_7924,N_4371,N_2276);
nor U7925 (N_7925,N_4666,N_4583);
or U7926 (N_7926,N_290,N_252);
and U7927 (N_7927,N_290,N_15);
xnor U7928 (N_7928,N_1919,N_4113);
xnor U7929 (N_7929,N_4699,N_1137);
and U7930 (N_7930,N_1112,N_4328);
and U7931 (N_7931,N_2024,N_2621);
nor U7932 (N_7932,N_4312,N_2615);
nand U7933 (N_7933,N_1310,N_2456);
nor U7934 (N_7934,N_1434,N_3191);
nand U7935 (N_7935,N_2643,N_1477);
and U7936 (N_7936,N_2364,N_4193);
or U7937 (N_7937,N_4201,N_46);
xor U7938 (N_7938,N_1142,N_4937);
xor U7939 (N_7939,N_832,N_3460);
xor U7940 (N_7940,N_2439,N_3412);
nand U7941 (N_7941,N_2516,N_2009);
nor U7942 (N_7942,N_223,N_1879);
and U7943 (N_7943,N_4533,N_1351);
xnor U7944 (N_7944,N_2648,N_3093);
xnor U7945 (N_7945,N_11,N_396);
xnor U7946 (N_7946,N_851,N_4158);
xnor U7947 (N_7947,N_384,N_4134);
xor U7948 (N_7948,N_2272,N_3267);
nor U7949 (N_7949,N_221,N_3750);
nand U7950 (N_7950,N_2246,N_1474);
xor U7951 (N_7951,N_2594,N_1597);
xor U7952 (N_7952,N_208,N_3413);
nand U7953 (N_7953,N_4769,N_1521);
nor U7954 (N_7954,N_4594,N_2652);
nand U7955 (N_7955,N_1278,N_306);
or U7956 (N_7956,N_3936,N_988);
and U7957 (N_7957,N_4233,N_1074);
nand U7958 (N_7958,N_3861,N_1054);
nor U7959 (N_7959,N_4627,N_3729);
or U7960 (N_7960,N_2582,N_4139);
or U7961 (N_7961,N_4691,N_182);
nor U7962 (N_7962,N_4450,N_381);
nand U7963 (N_7963,N_4385,N_1336);
and U7964 (N_7964,N_4636,N_1928);
xor U7965 (N_7965,N_2358,N_402);
and U7966 (N_7966,N_1218,N_3837);
and U7967 (N_7967,N_2006,N_1324);
and U7968 (N_7968,N_1667,N_2062);
xor U7969 (N_7969,N_2914,N_1065);
nand U7970 (N_7970,N_829,N_1446);
nor U7971 (N_7971,N_4558,N_1330);
nand U7972 (N_7972,N_1612,N_1394);
nor U7973 (N_7973,N_3900,N_4437);
nor U7974 (N_7974,N_4833,N_2963);
or U7975 (N_7975,N_3393,N_1995);
xnor U7976 (N_7976,N_4228,N_1905);
or U7977 (N_7977,N_313,N_3765);
xnor U7978 (N_7978,N_3319,N_1981);
xnor U7979 (N_7979,N_4039,N_2579);
or U7980 (N_7980,N_4585,N_1352);
and U7981 (N_7981,N_3115,N_4651);
and U7982 (N_7982,N_3060,N_4115);
nand U7983 (N_7983,N_4177,N_411);
xnor U7984 (N_7984,N_3358,N_2528);
nand U7985 (N_7985,N_366,N_3433);
nor U7986 (N_7986,N_1796,N_2173);
and U7987 (N_7987,N_1638,N_2544);
and U7988 (N_7988,N_3886,N_2101);
nor U7989 (N_7989,N_3146,N_185);
nand U7990 (N_7990,N_2802,N_4073);
nand U7991 (N_7991,N_176,N_1548);
nor U7992 (N_7992,N_3355,N_4709);
nor U7993 (N_7993,N_2922,N_73);
and U7994 (N_7994,N_2317,N_2782);
nand U7995 (N_7995,N_3505,N_3175);
and U7996 (N_7996,N_3119,N_3478);
and U7997 (N_7997,N_2822,N_1110);
xor U7998 (N_7998,N_2564,N_651);
or U7999 (N_7999,N_4999,N_4205);
xnor U8000 (N_8000,N_1139,N_638);
xor U8001 (N_8001,N_4972,N_1047);
nor U8002 (N_8002,N_3522,N_709);
and U8003 (N_8003,N_4697,N_2109);
nor U8004 (N_8004,N_833,N_4419);
or U8005 (N_8005,N_2597,N_3988);
xor U8006 (N_8006,N_2422,N_2851);
xor U8007 (N_8007,N_3285,N_4989);
and U8008 (N_8008,N_3816,N_1085);
nor U8009 (N_8009,N_846,N_2469);
nor U8010 (N_8010,N_1375,N_2282);
or U8011 (N_8011,N_2716,N_4287);
nor U8012 (N_8012,N_2169,N_1984);
nor U8013 (N_8013,N_585,N_967);
xor U8014 (N_8014,N_3455,N_1162);
xnor U8015 (N_8015,N_3830,N_3025);
and U8016 (N_8016,N_732,N_3304);
xnor U8017 (N_8017,N_1369,N_4186);
or U8018 (N_8018,N_3756,N_1142);
nand U8019 (N_8019,N_764,N_1639);
xor U8020 (N_8020,N_593,N_3099);
nor U8021 (N_8021,N_237,N_4553);
nand U8022 (N_8022,N_4702,N_466);
nand U8023 (N_8023,N_735,N_3918);
and U8024 (N_8024,N_2677,N_1541);
nor U8025 (N_8025,N_4309,N_629);
nor U8026 (N_8026,N_3891,N_3149);
and U8027 (N_8027,N_2972,N_1137);
and U8028 (N_8028,N_168,N_911);
nand U8029 (N_8029,N_3878,N_507);
and U8030 (N_8030,N_863,N_2039);
and U8031 (N_8031,N_1724,N_4788);
or U8032 (N_8032,N_769,N_575);
nand U8033 (N_8033,N_3757,N_498);
nor U8034 (N_8034,N_4267,N_1117);
xor U8035 (N_8035,N_4730,N_3155);
nand U8036 (N_8036,N_1268,N_1019);
nor U8037 (N_8037,N_2485,N_1313);
nor U8038 (N_8038,N_4518,N_2438);
nor U8039 (N_8039,N_4792,N_2143);
nand U8040 (N_8040,N_3182,N_1991);
or U8041 (N_8041,N_4803,N_2923);
xor U8042 (N_8042,N_1260,N_4397);
or U8043 (N_8043,N_3816,N_53);
xor U8044 (N_8044,N_3393,N_3004);
xnor U8045 (N_8045,N_1456,N_2803);
nand U8046 (N_8046,N_2318,N_1587);
xor U8047 (N_8047,N_216,N_2297);
nand U8048 (N_8048,N_1035,N_369);
and U8049 (N_8049,N_1959,N_3520);
nand U8050 (N_8050,N_800,N_3744);
nand U8051 (N_8051,N_3805,N_4790);
nor U8052 (N_8052,N_2367,N_458);
nand U8053 (N_8053,N_2773,N_4563);
and U8054 (N_8054,N_3845,N_477);
nand U8055 (N_8055,N_770,N_3053);
nor U8056 (N_8056,N_2902,N_2014);
nor U8057 (N_8057,N_805,N_1175);
or U8058 (N_8058,N_480,N_855);
nor U8059 (N_8059,N_4137,N_3653);
or U8060 (N_8060,N_4418,N_3985);
xnor U8061 (N_8061,N_2581,N_4511);
or U8062 (N_8062,N_3510,N_288);
nor U8063 (N_8063,N_2929,N_1055);
or U8064 (N_8064,N_3119,N_4931);
nand U8065 (N_8065,N_3819,N_718);
nor U8066 (N_8066,N_2309,N_4798);
nand U8067 (N_8067,N_1591,N_709);
or U8068 (N_8068,N_2328,N_2477);
nor U8069 (N_8069,N_870,N_4618);
and U8070 (N_8070,N_1762,N_949);
xnor U8071 (N_8071,N_4898,N_4399);
and U8072 (N_8072,N_4802,N_1756);
and U8073 (N_8073,N_3294,N_2739);
nand U8074 (N_8074,N_1164,N_2615);
and U8075 (N_8075,N_3431,N_4674);
xnor U8076 (N_8076,N_2412,N_2755);
nor U8077 (N_8077,N_890,N_323);
and U8078 (N_8078,N_2794,N_3732);
and U8079 (N_8079,N_170,N_1673);
or U8080 (N_8080,N_4103,N_4246);
and U8081 (N_8081,N_4909,N_3346);
nand U8082 (N_8082,N_19,N_2203);
nor U8083 (N_8083,N_867,N_4556);
nor U8084 (N_8084,N_4976,N_1172);
or U8085 (N_8085,N_1001,N_1097);
or U8086 (N_8086,N_1955,N_3665);
nand U8087 (N_8087,N_3926,N_1946);
nor U8088 (N_8088,N_4870,N_275);
or U8089 (N_8089,N_4285,N_702);
xor U8090 (N_8090,N_4238,N_4287);
nand U8091 (N_8091,N_397,N_709);
xnor U8092 (N_8092,N_4169,N_1791);
and U8093 (N_8093,N_4624,N_1546);
xnor U8094 (N_8094,N_3788,N_2992);
nor U8095 (N_8095,N_870,N_3798);
nor U8096 (N_8096,N_1633,N_684);
nand U8097 (N_8097,N_334,N_2818);
or U8098 (N_8098,N_682,N_3330);
nor U8099 (N_8099,N_2758,N_1045);
or U8100 (N_8100,N_3673,N_2716);
nand U8101 (N_8101,N_4879,N_2705);
nand U8102 (N_8102,N_1792,N_1972);
xor U8103 (N_8103,N_2973,N_3662);
xnor U8104 (N_8104,N_4630,N_4845);
and U8105 (N_8105,N_3680,N_3202);
or U8106 (N_8106,N_1311,N_841);
and U8107 (N_8107,N_380,N_632);
nand U8108 (N_8108,N_85,N_803);
or U8109 (N_8109,N_4974,N_1080);
or U8110 (N_8110,N_4326,N_2041);
or U8111 (N_8111,N_3787,N_1999);
or U8112 (N_8112,N_2828,N_601);
xor U8113 (N_8113,N_2657,N_2842);
nand U8114 (N_8114,N_4407,N_481);
or U8115 (N_8115,N_3694,N_299);
and U8116 (N_8116,N_3117,N_3695);
nor U8117 (N_8117,N_402,N_3022);
xor U8118 (N_8118,N_189,N_329);
nand U8119 (N_8119,N_1980,N_3741);
nand U8120 (N_8120,N_4916,N_1154);
nor U8121 (N_8121,N_4257,N_3755);
xnor U8122 (N_8122,N_2798,N_1985);
or U8123 (N_8123,N_2839,N_200);
and U8124 (N_8124,N_1408,N_4071);
or U8125 (N_8125,N_2080,N_2827);
or U8126 (N_8126,N_2573,N_1898);
and U8127 (N_8127,N_2380,N_4117);
nor U8128 (N_8128,N_1563,N_40);
and U8129 (N_8129,N_2913,N_2031);
and U8130 (N_8130,N_4341,N_3017);
and U8131 (N_8131,N_1883,N_4229);
nand U8132 (N_8132,N_2017,N_1689);
and U8133 (N_8133,N_4423,N_3952);
nor U8134 (N_8134,N_3997,N_2584);
nand U8135 (N_8135,N_4117,N_2450);
or U8136 (N_8136,N_1379,N_157);
nor U8137 (N_8137,N_3963,N_2629);
xor U8138 (N_8138,N_4675,N_584);
nor U8139 (N_8139,N_1149,N_534);
or U8140 (N_8140,N_3433,N_3758);
xnor U8141 (N_8141,N_4177,N_1451);
nor U8142 (N_8142,N_3221,N_4138);
and U8143 (N_8143,N_2367,N_3683);
nor U8144 (N_8144,N_3630,N_1963);
nor U8145 (N_8145,N_3610,N_3872);
and U8146 (N_8146,N_3907,N_760);
xor U8147 (N_8147,N_2219,N_1835);
xnor U8148 (N_8148,N_994,N_3676);
xnor U8149 (N_8149,N_4996,N_4358);
and U8150 (N_8150,N_12,N_4117);
and U8151 (N_8151,N_3305,N_4788);
xor U8152 (N_8152,N_3916,N_3170);
nor U8153 (N_8153,N_1952,N_2285);
xnor U8154 (N_8154,N_792,N_863);
xor U8155 (N_8155,N_2858,N_20);
xnor U8156 (N_8156,N_3910,N_2968);
or U8157 (N_8157,N_4029,N_3279);
nand U8158 (N_8158,N_704,N_2740);
nor U8159 (N_8159,N_2877,N_93);
nor U8160 (N_8160,N_3566,N_85);
and U8161 (N_8161,N_4902,N_2934);
or U8162 (N_8162,N_294,N_3104);
nor U8163 (N_8163,N_1733,N_2320);
or U8164 (N_8164,N_1309,N_2289);
nand U8165 (N_8165,N_3529,N_2998);
nand U8166 (N_8166,N_3497,N_391);
nand U8167 (N_8167,N_521,N_4124);
nor U8168 (N_8168,N_3969,N_998);
nand U8169 (N_8169,N_59,N_722);
nor U8170 (N_8170,N_4914,N_1297);
and U8171 (N_8171,N_3534,N_922);
and U8172 (N_8172,N_2442,N_1273);
xnor U8173 (N_8173,N_3510,N_732);
nor U8174 (N_8174,N_4802,N_4859);
nor U8175 (N_8175,N_3311,N_4783);
and U8176 (N_8176,N_4590,N_2853);
or U8177 (N_8177,N_2819,N_3763);
or U8178 (N_8178,N_369,N_858);
or U8179 (N_8179,N_2653,N_1358);
and U8180 (N_8180,N_1010,N_1900);
nor U8181 (N_8181,N_953,N_3906);
and U8182 (N_8182,N_2844,N_173);
nor U8183 (N_8183,N_4756,N_2926);
xnor U8184 (N_8184,N_459,N_1792);
nor U8185 (N_8185,N_4999,N_3676);
nand U8186 (N_8186,N_3804,N_3056);
or U8187 (N_8187,N_4309,N_4784);
nand U8188 (N_8188,N_4476,N_2065);
and U8189 (N_8189,N_279,N_1852);
nor U8190 (N_8190,N_3182,N_4051);
nand U8191 (N_8191,N_1209,N_4834);
and U8192 (N_8192,N_4281,N_2585);
or U8193 (N_8193,N_2421,N_2937);
nor U8194 (N_8194,N_4752,N_4565);
nor U8195 (N_8195,N_3861,N_250);
xor U8196 (N_8196,N_3998,N_2349);
xor U8197 (N_8197,N_4686,N_4278);
or U8198 (N_8198,N_1473,N_3436);
or U8199 (N_8199,N_3913,N_3640);
and U8200 (N_8200,N_746,N_1199);
nor U8201 (N_8201,N_259,N_1654);
xor U8202 (N_8202,N_2348,N_1498);
nor U8203 (N_8203,N_359,N_1964);
nor U8204 (N_8204,N_4420,N_1415);
nor U8205 (N_8205,N_1370,N_4361);
nand U8206 (N_8206,N_4693,N_4313);
xnor U8207 (N_8207,N_4569,N_4008);
nand U8208 (N_8208,N_3422,N_1905);
xor U8209 (N_8209,N_4972,N_4371);
nor U8210 (N_8210,N_1272,N_2663);
nand U8211 (N_8211,N_3152,N_3433);
nor U8212 (N_8212,N_4818,N_50);
and U8213 (N_8213,N_1712,N_2926);
nand U8214 (N_8214,N_3607,N_2675);
nor U8215 (N_8215,N_1691,N_1010);
xnor U8216 (N_8216,N_2844,N_766);
or U8217 (N_8217,N_3698,N_3461);
and U8218 (N_8218,N_4662,N_2);
or U8219 (N_8219,N_254,N_2485);
nand U8220 (N_8220,N_3254,N_1452);
or U8221 (N_8221,N_4243,N_3044);
xor U8222 (N_8222,N_1201,N_3081);
and U8223 (N_8223,N_2292,N_2966);
nand U8224 (N_8224,N_3113,N_3133);
xnor U8225 (N_8225,N_2811,N_2135);
and U8226 (N_8226,N_4423,N_2712);
nand U8227 (N_8227,N_1738,N_2268);
or U8228 (N_8228,N_2846,N_3895);
and U8229 (N_8229,N_2760,N_1785);
and U8230 (N_8230,N_4213,N_4738);
or U8231 (N_8231,N_938,N_1084);
and U8232 (N_8232,N_3454,N_3721);
or U8233 (N_8233,N_1150,N_3220);
nor U8234 (N_8234,N_142,N_4862);
or U8235 (N_8235,N_1106,N_2959);
or U8236 (N_8236,N_1194,N_525);
nand U8237 (N_8237,N_4521,N_3994);
nand U8238 (N_8238,N_3352,N_1297);
nand U8239 (N_8239,N_2045,N_3803);
nor U8240 (N_8240,N_151,N_2002);
xor U8241 (N_8241,N_3454,N_3038);
or U8242 (N_8242,N_523,N_12);
xnor U8243 (N_8243,N_2218,N_584);
xnor U8244 (N_8244,N_2144,N_2150);
nand U8245 (N_8245,N_895,N_886);
nand U8246 (N_8246,N_4531,N_2280);
nor U8247 (N_8247,N_615,N_538);
nand U8248 (N_8248,N_2173,N_3420);
nor U8249 (N_8249,N_4378,N_380);
xnor U8250 (N_8250,N_3211,N_2906);
or U8251 (N_8251,N_3406,N_3438);
or U8252 (N_8252,N_3625,N_2467);
nand U8253 (N_8253,N_3177,N_1897);
nand U8254 (N_8254,N_2521,N_2992);
nand U8255 (N_8255,N_373,N_1897);
xnor U8256 (N_8256,N_2168,N_3161);
nand U8257 (N_8257,N_4717,N_3233);
and U8258 (N_8258,N_975,N_4004);
or U8259 (N_8259,N_4958,N_2290);
nor U8260 (N_8260,N_4465,N_3805);
nand U8261 (N_8261,N_3216,N_1638);
nor U8262 (N_8262,N_1895,N_2551);
and U8263 (N_8263,N_2082,N_1961);
or U8264 (N_8264,N_2112,N_4958);
or U8265 (N_8265,N_3722,N_3869);
xnor U8266 (N_8266,N_2710,N_4844);
nand U8267 (N_8267,N_799,N_4356);
nor U8268 (N_8268,N_4265,N_4586);
nand U8269 (N_8269,N_3733,N_81);
and U8270 (N_8270,N_318,N_3064);
nand U8271 (N_8271,N_4399,N_2189);
or U8272 (N_8272,N_3851,N_4523);
xor U8273 (N_8273,N_1028,N_1655);
nand U8274 (N_8274,N_4501,N_647);
or U8275 (N_8275,N_3002,N_565);
and U8276 (N_8276,N_867,N_395);
and U8277 (N_8277,N_4485,N_2018);
xnor U8278 (N_8278,N_4677,N_2214);
or U8279 (N_8279,N_2209,N_1055);
and U8280 (N_8280,N_918,N_1733);
xor U8281 (N_8281,N_2112,N_1211);
and U8282 (N_8282,N_1605,N_1034);
nand U8283 (N_8283,N_4410,N_4388);
or U8284 (N_8284,N_4916,N_2434);
nand U8285 (N_8285,N_4755,N_2647);
nor U8286 (N_8286,N_2555,N_30);
xor U8287 (N_8287,N_4560,N_2480);
xor U8288 (N_8288,N_214,N_1659);
xor U8289 (N_8289,N_4131,N_600);
and U8290 (N_8290,N_230,N_3569);
xnor U8291 (N_8291,N_4898,N_1419);
xor U8292 (N_8292,N_1844,N_3766);
xnor U8293 (N_8293,N_3774,N_2885);
xnor U8294 (N_8294,N_1481,N_4192);
nor U8295 (N_8295,N_2171,N_1763);
nor U8296 (N_8296,N_2325,N_2382);
nor U8297 (N_8297,N_1742,N_3230);
and U8298 (N_8298,N_3302,N_3700);
nand U8299 (N_8299,N_4606,N_1252);
xnor U8300 (N_8300,N_4841,N_3508);
xor U8301 (N_8301,N_976,N_663);
and U8302 (N_8302,N_4450,N_4863);
nand U8303 (N_8303,N_511,N_1694);
nor U8304 (N_8304,N_2981,N_3260);
nand U8305 (N_8305,N_4116,N_2194);
nand U8306 (N_8306,N_2232,N_1230);
nor U8307 (N_8307,N_3263,N_1264);
nand U8308 (N_8308,N_2279,N_2852);
nor U8309 (N_8309,N_2499,N_3587);
nand U8310 (N_8310,N_494,N_2279);
nor U8311 (N_8311,N_2224,N_949);
and U8312 (N_8312,N_1816,N_1373);
nand U8313 (N_8313,N_4530,N_3370);
xnor U8314 (N_8314,N_3775,N_2069);
or U8315 (N_8315,N_1993,N_4804);
xnor U8316 (N_8316,N_672,N_904);
and U8317 (N_8317,N_4651,N_3833);
nor U8318 (N_8318,N_3440,N_4994);
nor U8319 (N_8319,N_4046,N_2798);
nor U8320 (N_8320,N_2808,N_318);
nor U8321 (N_8321,N_1039,N_2244);
nand U8322 (N_8322,N_3203,N_405);
xor U8323 (N_8323,N_2009,N_4021);
nand U8324 (N_8324,N_4286,N_117);
xor U8325 (N_8325,N_3403,N_1849);
nor U8326 (N_8326,N_4106,N_3149);
or U8327 (N_8327,N_4081,N_3290);
and U8328 (N_8328,N_4138,N_1620);
nor U8329 (N_8329,N_3292,N_1259);
nor U8330 (N_8330,N_475,N_1442);
or U8331 (N_8331,N_3311,N_4316);
and U8332 (N_8332,N_1795,N_4486);
nand U8333 (N_8333,N_4659,N_2083);
xor U8334 (N_8334,N_320,N_1498);
nand U8335 (N_8335,N_3983,N_1948);
or U8336 (N_8336,N_1777,N_4416);
xor U8337 (N_8337,N_13,N_222);
nand U8338 (N_8338,N_2437,N_4907);
nor U8339 (N_8339,N_3751,N_2599);
nand U8340 (N_8340,N_3395,N_1508);
nor U8341 (N_8341,N_1429,N_3732);
xnor U8342 (N_8342,N_235,N_1287);
or U8343 (N_8343,N_2132,N_2450);
nand U8344 (N_8344,N_1799,N_401);
and U8345 (N_8345,N_1098,N_46);
nor U8346 (N_8346,N_2959,N_208);
xor U8347 (N_8347,N_901,N_4790);
xnor U8348 (N_8348,N_4078,N_1888);
nor U8349 (N_8349,N_347,N_1284);
nor U8350 (N_8350,N_1963,N_1161);
nor U8351 (N_8351,N_1082,N_4710);
and U8352 (N_8352,N_4508,N_3859);
xnor U8353 (N_8353,N_3054,N_37);
or U8354 (N_8354,N_2737,N_3043);
nand U8355 (N_8355,N_1571,N_540);
xor U8356 (N_8356,N_3567,N_4871);
xor U8357 (N_8357,N_2872,N_3853);
nor U8358 (N_8358,N_4412,N_2928);
or U8359 (N_8359,N_2311,N_3465);
nor U8360 (N_8360,N_1894,N_4143);
and U8361 (N_8361,N_3005,N_3058);
xor U8362 (N_8362,N_4465,N_1640);
xor U8363 (N_8363,N_1174,N_4289);
or U8364 (N_8364,N_2075,N_3044);
or U8365 (N_8365,N_664,N_1449);
nand U8366 (N_8366,N_4544,N_46);
nor U8367 (N_8367,N_3482,N_567);
nand U8368 (N_8368,N_4721,N_3276);
xnor U8369 (N_8369,N_1499,N_1066);
nor U8370 (N_8370,N_3205,N_175);
nor U8371 (N_8371,N_1788,N_1237);
nor U8372 (N_8372,N_38,N_1469);
or U8373 (N_8373,N_1955,N_884);
and U8374 (N_8374,N_1189,N_1939);
nand U8375 (N_8375,N_3281,N_1805);
or U8376 (N_8376,N_4055,N_1009);
xor U8377 (N_8377,N_2406,N_4790);
and U8378 (N_8378,N_2580,N_301);
or U8379 (N_8379,N_2091,N_141);
nand U8380 (N_8380,N_4205,N_2198);
nand U8381 (N_8381,N_2074,N_1346);
or U8382 (N_8382,N_2794,N_3028);
xnor U8383 (N_8383,N_451,N_2790);
and U8384 (N_8384,N_954,N_2512);
nand U8385 (N_8385,N_4261,N_2869);
or U8386 (N_8386,N_2030,N_1989);
or U8387 (N_8387,N_4546,N_4638);
and U8388 (N_8388,N_2500,N_1496);
or U8389 (N_8389,N_2424,N_545);
and U8390 (N_8390,N_3461,N_1633);
nor U8391 (N_8391,N_283,N_1398);
or U8392 (N_8392,N_2042,N_2237);
or U8393 (N_8393,N_1569,N_474);
nand U8394 (N_8394,N_3149,N_861);
nand U8395 (N_8395,N_3368,N_836);
nand U8396 (N_8396,N_587,N_3403);
nand U8397 (N_8397,N_3296,N_3017);
and U8398 (N_8398,N_4264,N_1118);
and U8399 (N_8399,N_4675,N_319);
nand U8400 (N_8400,N_3258,N_1873);
and U8401 (N_8401,N_1299,N_3283);
xnor U8402 (N_8402,N_4723,N_1241);
or U8403 (N_8403,N_1143,N_3874);
nand U8404 (N_8404,N_2750,N_2678);
xnor U8405 (N_8405,N_4248,N_3024);
nand U8406 (N_8406,N_4113,N_2850);
or U8407 (N_8407,N_4948,N_3971);
and U8408 (N_8408,N_1984,N_4339);
nand U8409 (N_8409,N_2265,N_3536);
nand U8410 (N_8410,N_2736,N_2874);
nor U8411 (N_8411,N_367,N_4250);
and U8412 (N_8412,N_2942,N_3180);
nand U8413 (N_8413,N_1277,N_3880);
or U8414 (N_8414,N_1986,N_4997);
and U8415 (N_8415,N_4924,N_465);
or U8416 (N_8416,N_2489,N_1669);
nand U8417 (N_8417,N_3096,N_2158);
nand U8418 (N_8418,N_2223,N_376);
nor U8419 (N_8419,N_2103,N_2718);
or U8420 (N_8420,N_27,N_3290);
xor U8421 (N_8421,N_512,N_1727);
and U8422 (N_8422,N_4583,N_3400);
xor U8423 (N_8423,N_2427,N_2824);
xnor U8424 (N_8424,N_4715,N_2389);
nand U8425 (N_8425,N_391,N_4497);
nand U8426 (N_8426,N_3376,N_2824);
nor U8427 (N_8427,N_1058,N_1316);
and U8428 (N_8428,N_884,N_2217);
nand U8429 (N_8429,N_3823,N_2126);
nor U8430 (N_8430,N_2837,N_192);
nand U8431 (N_8431,N_1854,N_2775);
or U8432 (N_8432,N_4961,N_1098);
xnor U8433 (N_8433,N_2463,N_4415);
and U8434 (N_8434,N_4222,N_4102);
or U8435 (N_8435,N_3334,N_53);
nand U8436 (N_8436,N_4788,N_4939);
nand U8437 (N_8437,N_4806,N_1217);
and U8438 (N_8438,N_4902,N_1526);
xor U8439 (N_8439,N_4497,N_275);
nand U8440 (N_8440,N_3841,N_3177);
or U8441 (N_8441,N_1681,N_4174);
or U8442 (N_8442,N_4051,N_1751);
and U8443 (N_8443,N_1353,N_620);
nor U8444 (N_8444,N_3316,N_2593);
or U8445 (N_8445,N_2883,N_3269);
nand U8446 (N_8446,N_2422,N_2930);
and U8447 (N_8447,N_1483,N_1732);
nand U8448 (N_8448,N_2908,N_3162);
and U8449 (N_8449,N_2502,N_2905);
or U8450 (N_8450,N_2120,N_4053);
nor U8451 (N_8451,N_4365,N_806);
xnor U8452 (N_8452,N_4112,N_1831);
nand U8453 (N_8453,N_3723,N_3016);
or U8454 (N_8454,N_189,N_4549);
or U8455 (N_8455,N_599,N_4804);
xnor U8456 (N_8456,N_4088,N_707);
xnor U8457 (N_8457,N_243,N_4498);
or U8458 (N_8458,N_2822,N_886);
and U8459 (N_8459,N_3493,N_3025);
and U8460 (N_8460,N_435,N_3468);
xor U8461 (N_8461,N_4049,N_549);
nor U8462 (N_8462,N_1217,N_1169);
xor U8463 (N_8463,N_3602,N_13);
and U8464 (N_8464,N_4888,N_2981);
and U8465 (N_8465,N_3990,N_1045);
xnor U8466 (N_8466,N_614,N_2161);
or U8467 (N_8467,N_3651,N_104);
nor U8468 (N_8468,N_4618,N_4646);
or U8469 (N_8469,N_2286,N_2774);
or U8470 (N_8470,N_3563,N_4396);
or U8471 (N_8471,N_2792,N_4782);
or U8472 (N_8472,N_1636,N_1001);
nand U8473 (N_8473,N_103,N_4999);
nand U8474 (N_8474,N_4604,N_402);
nor U8475 (N_8475,N_1639,N_2508);
and U8476 (N_8476,N_2441,N_1814);
xnor U8477 (N_8477,N_2454,N_481);
xnor U8478 (N_8478,N_1439,N_4299);
nand U8479 (N_8479,N_4790,N_2654);
and U8480 (N_8480,N_1543,N_1424);
and U8481 (N_8481,N_3737,N_1924);
nor U8482 (N_8482,N_4645,N_44);
nor U8483 (N_8483,N_3092,N_4319);
xor U8484 (N_8484,N_2623,N_1710);
and U8485 (N_8485,N_1119,N_2100);
or U8486 (N_8486,N_4371,N_4591);
xor U8487 (N_8487,N_250,N_1131);
nand U8488 (N_8488,N_806,N_2491);
nor U8489 (N_8489,N_3395,N_4561);
xnor U8490 (N_8490,N_3566,N_872);
and U8491 (N_8491,N_1965,N_3295);
or U8492 (N_8492,N_1868,N_2418);
or U8493 (N_8493,N_1532,N_3661);
or U8494 (N_8494,N_3346,N_310);
nor U8495 (N_8495,N_2706,N_4752);
xor U8496 (N_8496,N_1946,N_2940);
or U8497 (N_8497,N_835,N_4321);
nand U8498 (N_8498,N_3978,N_4396);
nor U8499 (N_8499,N_825,N_3332);
xor U8500 (N_8500,N_1032,N_4538);
xor U8501 (N_8501,N_4642,N_2016);
xnor U8502 (N_8502,N_3608,N_3258);
xor U8503 (N_8503,N_4189,N_4648);
nand U8504 (N_8504,N_4958,N_2674);
xor U8505 (N_8505,N_4599,N_3539);
nor U8506 (N_8506,N_4115,N_1962);
and U8507 (N_8507,N_1632,N_4701);
nor U8508 (N_8508,N_3679,N_3375);
and U8509 (N_8509,N_3130,N_4301);
xor U8510 (N_8510,N_782,N_2110);
nand U8511 (N_8511,N_1779,N_1758);
nand U8512 (N_8512,N_1348,N_935);
nand U8513 (N_8513,N_1789,N_2857);
or U8514 (N_8514,N_4244,N_3358);
and U8515 (N_8515,N_3331,N_12);
nand U8516 (N_8516,N_3782,N_426);
xor U8517 (N_8517,N_2682,N_473);
nor U8518 (N_8518,N_1452,N_1040);
or U8519 (N_8519,N_4589,N_3796);
or U8520 (N_8520,N_3510,N_2177);
nand U8521 (N_8521,N_4792,N_414);
nor U8522 (N_8522,N_1726,N_96);
nand U8523 (N_8523,N_2062,N_2743);
or U8524 (N_8524,N_4977,N_1691);
and U8525 (N_8525,N_1448,N_3306);
and U8526 (N_8526,N_1976,N_2172);
nor U8527 (N_8527,N_210,N_2144);
nand U8528 (N_8528,N_3617,N_4966);
nor U8529 (N_8529,N_2646,N_4311);
and U8530 (N_8530,N_1460,N_1305);
xor U8531 (N_8531,N_1334,N_3184);
and U8532 (N_8532,N_2613,N_3312);
nor U8533 (N_8533,N_627,N_4229);
nand U8534 (N_8534,N_1380,N_2971);
nor U8535 (N_8535,N_1298,N_4958);
xnor U8536 (N_8536,N_4858,N_3594);
xnor U8537 (N_8537,N_2221,N_1298);
nor U8538 (N_8538,N_1713,N_1715);
nand U8539 (N_8539,N_734,N_4338);
or U8540 (N_8540,N_2727,N_4461);
or U8541 (N_8541,N_3147,N_2713);
nand U8542 (N_8542,N_2708,N_2754);
and U8543 (N_8543,N_4918,N_2934);
nor U8544 (N_8544,N_3441,N_2992);
and U8545 (N_8545,N_437,N_2051);
or U8546 (N_8546,N_2114,N_1885);
and U8547 (N_8547,N_3812,N_1480);
xor U8548 (N_8548,N_2110,N_3573);
nor U8549 (N_8549,N_2197,N_1581);
or U8550 (N_8550,N_1695,N_1771);
and U8551 (N_8551,N_965,N_2958);
xor U8552 (N_8552,N_2987,N_3517);
nor U8553 (N_8553,N_1704,N_3720);
nand U8554 (N_8554,N_2976,N_3538);
and U8555 (N_8555,N_3011,N_1314);
or U8556 (N_8556,N_2453,N_717);
nand U8557 (N_8557,N_1491,N_2450);
nand U8558 (N_8558,N_2979,N_938);
nor U8559 (N_8559,N_3099,N_1943);
nor U8560 (N_8560,N_4775,N_3672);
nor U8561 (N_8561,N_4692,N_798);
nand U8562 (N_8562,N_3385,N_3309);
nor U8563 (N_8563,N_4243,N_2939);
nor U8564 (N_8564,N_970,N_2772);
and U8565 (N_8565,N_56,N_907);
and U8566 (N_8566,N_4467,N_1964);
and U8567 (N_8567,N_1255,N_4467);
and U8568 (N_8568,N_3104,N_4426);
nand U8569 (N_8569,N_1581,N_3105);
nand U8570 (N_8570,N_4452,N_3293);
or U8571 (N_8571,N_1452,N_68);
or U8572 (N_8572,N_397,N_752);
xor U8573 (N_8573,N_3202,N_4431);
nor U8574 (N_8574,N_90,N_104);
and U8575 (N_8575,N_642,N_2661);
or U8576 (N_8576,N_3950,N_3094);
and U8577 (N_8577,N_3079,N_2715);
nor U8578 (N_8578,N_93,N_2391);
or U8579 (N_8579,N_4635,N_2607);
xor U8580 (N_8580,N_3615,N_2376);
nor U8581 (N_8581,N_2646,N_268);
xor U8582 (N_8582,N_3846,N_4854);
nor U8583 (N_8583,N_2932,N_501);
and U8584 (N_8584,N_765,N_1487);
and U8585 (N_8585,N_4823,N_1015);
nor U8586 (N_8586,N_3560,N_2644);
or U8587 (N_8587,N_4842,N_3601);
or U8588 (N_8588,N_777,N_64);
or U8589 (N_8589,N_4995,N_684);
nor U8590 (N_8590,N_3548,N_4320);
nand U8591 (N_8591,N_3734,N_167);
xor U8592 (N_8592,N_1675,N_1094);
nor U8593 (N_8593,N_397,N_913);
xnor U8594 (N_8594,N_1550,N_3730);
nand U8595 (N_8595,N_3006,N_1603);
xnor U8596 (N_8596,N_1933,N_3593);
and U8597 (N_8597,N_353,N_3187);
nor U8598 (N_8598,N_3630,N_3645);
nor U8599 (N_8599,N_2759,N_1309);
nand U8600 (N_8600,N_3184,N_2898);
nand U8601 (N_8601,N_3562,N_4862);
and U8602 (N_8602,N_4015,N_2514);
xor U8603 (N_8603,N_4315,N_3330);
nor U8604 (N_8604,N_624,N_805);
nand U8605 (N_8605,N_1190,N_938);
and U8606 (N_8606,N_2343,N_3950);
xor U8607 (N_8607,N_427,N_2802);
or U8608 (N_8608,N_4390,N_4565);
nor U8609 (N_8609,N_1590,N_3933);
nand U8610 (N_8610,N_4039,N_4535);
nand U8611 (N_8611,N_2602,N_118);
or U8612 (N_8612,N_1232,N_3784);
nor U8613 (N_8613,N_3692,N_3704);
nand U8614 (N_8614,N_4587,N_2111);
xnor U8615 (N_8615,N_1677,N_3475);
xor U8616 (N_8616,N_3582,N_2282);
nand U8617 (N_8617,N_527,N_825);
or U8618 (N_8618,N_2039,N_4555);
or U8619 (N_8619,N_1020,N_439);
or U8620 (N_8620,N_1701,N_2748);
nand U8621 (N_8621,N_1059,N_4211);
and U8622 (N_8622,N_27,N_2818);
or U8623 (N_8623,N_2233,N_428);
or U8624 (N_8624,N_4971,N_4656);
nor U8625 (N_8625,N_2434,N_3710);
nor U8626 (N_8626,N_865,N_1896);
or U8627 (N_8627,N_3115,N_1507);
and U8628 (N_8628,N_2648,N_2895);
xnor U8629 (N_8629,N_2477,N_257);
nand U8630 (N_8630,N_1390,N_3329);
nor U8631 (N_8631,N_187,N_954);
xor U8632 (N_8632,N_950,N_4185);
or U8633 (N_8633,N_1278,N_84);
xnor U8634 (N_8634,N_2428,N_3241);
nand U8635 (N_8635,N_4393,N_864);
nor U8636 (N_8636,N_4399,N_2890);
nand U8637 (N_8637,N_2347,N_287);
nand U8638 (N_8638,N_2002,N_2808);
xnor U8639 (N_8639,N_3811,N_1603);
and U8640 (N_8640,N_168,N_56);
and U8641 (N_8641,N_3660,N_679);
nor U8642 (N_8642,N_407,N_3238);
nand U8643 (N_8643,N_2468,N_3);
or U8644 (N_8644,N_294,N_780);
xnor U8645 (N_8645,N_2692,N_4737);
and U8646 (N_8646,N_3305,N_637);
or U8647 (N_8647,N_403,N_877);
nand U8648 (N_8648,N_3821,N_3647);
or U8649 (N_8649,N_4362,N_3622);
nand U8650 (N_8650,N_3247,N_2614);
or U8651 (N_8651,N_3378,N_63);
and U8652 (N_8652,N_1073,N_2579);
nor U8653 (N_8653,N_3201,N_3688);
nor U8654 (N_8654,N_2762,N_1540);
and U8655 (N_8655,N_851,N_2862);
nor U8656 (N_8656,N_3641,N_4789);
and U8657 (N_8657,N_3372,N_2668);
and U8658 (N_8658,N_4421,N_4767);
xor U8659 (N_8659,N_4687,N_3095);
nor U8660 (N_8660,N_3416,N_4328);
or U8661 (N_8661,N_422,N_1905);
or U8662 (N_8662,N_1992,N_516);
and U8663 (N_8663,N_323,N_907);
or U8664 (N_8664,N_2980,N_2778);
nor U8665 (N_8665,N_2909,N_4417);
xnor U8666 (N_8666,N_4229,N_1447);
nor U8667 (N_8667,N_2267,N_2197);
and U8668 (N_8668,N_3277,N_1346);
nor U8669 (N_8669,N_1584,N_791);
and U8670 (N_8670,N_1792,N_259);
and U8671 (N_8671,N_3652,N_969);
xnor U8672 (N_8672,N_2910,N_3685);
and U8673 (N_8673,N_4111,N_2205);
xor U8674 (N_8674,N_574,N_4338);
or U8675 (N_8675,N_1619,N_3985);
and U8676 (N_8676,N_3620,N_1023);
or U8677 (N_8677,N_2534,N_1865);
or U8678 (N_8678,N_4049,N_3138);
xnor U8679 (N_8679,N_2170,N_1340);
and U8680 (N_8680,N_17,N_3469);
nand U8681 (N_8681,N_2341,N_2018);
and U8682 (N_8682,N_3368,N_4801);
xnor U8683 (N_8683,N_4130,N_249);
and U8684 (N_8684,N_1969,N_1671);
and U8685 (N_8685,N_769,N_975);
and U8686 (N_8686,N_1572,N_2126);
nor U8687 (N_8687,N_994,N_3412);
and U8688 (N_8688,N_4488,N_4506);
xnor U8689 (N_8689,N_1432,N_4764);
and U8690 (N_8690,N_265,N_559);
xnor U8691 (N_8691,N_4575,N_3162);
xor U8692 (N_8692,N_2267,N_3585);
and U8693 (N_8693,N_2807,N_3988);
nor U8694 (N_8694,N_3527,N_4750);
nand U8695 (N_8695,N_445,N_3526);
nor U8696 (N_8696,N_397,N_3184);
or U8697 (N_8697,N_125,N_4786);
and U8698 (N_8698,N_4824,N_720);
or U8699 (N_8699,N_3877,N_2530);
nor U8700 (N_8700,N_2916,N_1017);
and U8701 (N_8701,N_763,N_2465);
nor U8702 (N_8702,N_3877,N_4157);
nor U8703 (N_8703,N_4411,N_2979);
nand U8704 (N_8704,N_316,N_3913);
and U8705 (N_8705,N_912,N_4190);
and U8706 (N_8706,N_1559,N_1612);
or U8707 (N_8707,N_4201,N_1420);
nand U8708 (N_8708,N_2780,N_1789);
and U8709 (N_8709,N_3592,N_2606);
nor U8710 (N_8710,N_219,N_1449);
or U8711 (N_8711,N_2341,N_1646);
xnor U8712 (N_8712,N_114,N_3038);
and U8713 (N_8713,N_2342,N_2437);
or U8714 (N_8714,N_99,N_4605);
nor U8715 (N_8715,N_4097,N_4579);
xnor U8716 (N_8716,N_2090,N_1816);
or U8717 (N_8717,N_3340,N_4729);
nand U8718 (N_8718,N_113,N_2291);
nor U8719 (N_8719,N_4428,N_1174);
nand U8720 (N_8720,N_983,N_188);
xnor U8721 (N_8721,N_4406,N_1875);
or U8722 (N_8722,N_3439,N_1502);
xor U8723 (N_8723,N_3950,N_118);
or U8724 (N_8724,N_1739,N_3585);
xnor U8725 (N_8725,N_3212,N_3131);
nand U8726 (N_8726,N_4055,N_1457);
nor U8727 (N_8727,N_4063,N_1900);
nand U8728 (N_8728,N_277,N_82);
and U8729 (N_8729,N_866,N_2508);
nor U8730 (N_8730,N_208,N_1802);
and U8731 (N_8731,N_3757,N_372);
or U8732 (N_8732,N_4624,N_33);
nor U8733 (N_8733,N_1242,N_1314);
nand U8734 (N_8734,N_3630,N_3355);
nand U8735 (N_8735,N_576,N_2419);
and U8736 (N_8736,N_3809,N_4156);
xor U8737 (N_8737,N_1330,N_1961);
and U8738 (N_8738,N_1691,N_4196);
xnor U8739 (N_8739,N_4030,N_2094);
nand U8740 (N_8740,N_1685,N_3602);
or U8741 (N_8741,N_4353,N_4379);
nor U8742 (N_8742,N_4861,N_3085);
nand U8743 (N_8743,N_2950,N_2119);
nor U8744 (N_8744,N_3578,N_3098);
xor U8745 (N_8745,N_2754,N_745);
nor U8746 (N_8746,N_678,N_1900);
or U8747 (N_8747,N_3332,N_4988);
or U8748 (N_8748,N_3496,N_1244);
nand U8749 (N_8749,N_2551,N_865);
and U8750 (N_8750,N_830,N_4762);
and U8751 (N_8751,N_1277,N_3833);
xnor U8752 (N_8752,N_3566,N_1087);
nand U8753 (N_8753,N_2574,N_2677);
nor U8754 (N_8754,N_3639,N_4668);
nand U8755 (N_8755,N_1864,N_1887);
and U8756 (N_8756,N_4282,N_2594);
nand U8757 (N_8757,N_732,N_532);
and U8758 (N_8758,N_1860,N_2808);
or U8759 (N_8759,N_4448,N_4974);
or U8760 (N_8760,N_2923,N_304);
nand U8761 (N_8761,N_1995,N_2338);
or U8762 (N_8762,N_3399,N_4385);
nor U8763 (N_8763,N_2587,N_4465);
nand U8764 (N_8764,N_1040,N_225);
or U8765 (N_8765,N_1495,N_1331);
or U8766 (N_8766,N_1784,N_3271);
nor U8767 (N_8767,N_507,N_536);
xnor U8768 (N_8768,N_4124,N_507);
and U8769 (N_8769,N_2709,N_2801);
or U8770 (N_8770,N_1555,N_2685);
nand U8771 (N_8771,N_1477,N_4101);
or U8772 (N_8772,N_760,N_957);
and U8773 (N_8773,N_2668,N_2726);
or U8774 (N_8774,N_4832,N_1469);
and U8775 (N_8775,N_1628,N_4516);
nand U8776 (N_8776,N_939,N_577);
or U8777 (N_8777,N_4788,N_4318);
nand U8778 (N_8778,N_244,N_352);
xor U8779 (N_8779,N_102,N_4480);
nor U8780 (N_8780,N_3192,N_1635);
nor U8781 (N_8781,N_1037,N_3196);
xnor U8782 (N_8782,N_3087,N_709);
and U8783 (N_8783,N_2256,N_4920);
or U8784 (N_8784,N_2205,N_2577);
nand U8785 (N_8785,N_3608,N_3206);
nor U8786 (N_8786,N_347,N_1108);
nand U8787 (N_8787,N_2069,N_4417);
and U8788 (N_8788,N_3185,N_1990);
nor U8789 (N_8789,N_2945,N_3076);
nand U8790 (N_8790,N_3324,N_719);
or U8791 (N_8791,N_3138,N_2852);
nand U8792 (N_8792,N_930,N_1428);
or U8793 (N_8793,N_341,N_4372);
nor U8794 (N_8794,N_576,N_1020);
xor U8795 (N_8795,N_2361,N_4451);
nand U8796 (N_8796,N_3638,N_457);
nor U8797 (N_8797,N_899,N_634);
xor U8798 (N_8798,N_3848,N_4185);
and U8799 (N_8799,N_1029,N_2097);
or U8800 (N_8800,N_3941,N_2034);
xor U8801 (N_8801,N_4036,N_2122);
nor U8802 (N_8802,N_1329,N_4028);
nor U8803 (N_8803,N_2175,N_2591);
nand U8804 (N_8804,N_1924,N_799);
nor U8805 (N_8805,N_1187,N_2683);
nand U8806 (N_8806,N_4212,N_3271);
or U8807 (N_8807,N_3503,N_619);
or U8808 (N_8808,N_235,N_3466);
and U8809 (N_8809,N_612,N_3369);
and U8810 (N_8810,N_2163,N_4438);
and U8811 (N_8811,N_4945,N_215);
nor U8812 (N_8812,N_4361,N_1780);
or U8813 (N_8813,N_664,N_4842);
nor U8814 (N_8814,N_4092,N_4932);
or U8815 (N_8815,N_181,N_4536);
or U8816 (N_8816,N_1887,N_2796);
and U8817 (N_8817,N_526,N_387);
and U8818 (N_8818,N_1731,N_4898);
xnor U8819 (N_8819,N_4790,N_2429);
nor U8820 (N_8820,N_1419,N_286);
nor U8821 (N_8821,N_116,N_3337);
xnor U8822 (N_8822,N_4715,N_4198);
nor U8823 (N_8823,N_712,N_386);
and U8824 (N_8824,N_2600,N_4042);
nor U8825 (N_8825,N_3656,N_3874);
or U8826 (N_8826,N_2785,N_4810);
or U8827 (N_8827,N_2141,N_2371);
nand U8828 (N_8828,N_2451,N_1410);
xor U8829 (N_8829,N_991,N_4132);
and U8830 (N_8830,N_4591,N_4349);
and U8831 (N_8831,N_3225,N_2688);
and U8832 (N_8832,N_4392,N_4400);
and U8833 (N_8833,N_4913,N_3985);
nor U8834 (N_8834,N_4738,N_903);
or U8835 (N_8835,N_2680,N_209);
nand U8836 (N_8836,N_1961,N_409);
or U8837 (N_8837,N_957,N_1028);
and U8838 (N_8838,N_4570,N_3869);
nand U8839 (N_8839,N_1657,N_1430);
or U8840 (N_8840,N_1327,N_1915);
nand U8841 (N_8841,N_2121,N_945);
xor U8842 (N_8842,N_1283,N_456);
and U8843 (N_8843,N_1818,N_1490);
nor U8844 (N_8844,N_4537,N_1695);
xnor U8845 (N_8845,N_3701,N_2240);
nor U8846 (N_8846,N_1271,N_2062);
or U8847 (N_8847,N_4899,N_3708);
or U8848 (N_8848,N_3745,N_435);
nand U8849 (N_8849,N_4256,N_1534);
nand U8850 (N_8850,N_1656,N_69);
and U8851 (N_8851,N_4383,N_3078);
xor U8852 (N_8852,N_1112,N_4772);
xor U8853 (N_8853,N_3748,N_4792);
nor U8854 (N_8854,N_3093,N_4056);
xor U8855 (N_8855,N_2882,N_4411);
and U8856 (N_8856,N_3959,N_2675);
and U8857 (N_8857,N_4250,N_2006);
nand U8858 (N_8858,N_1883,N_4292);
nor U8859 (N_8859,N_3626,N_20);
xnor U8860 (N_8860,N_2783,N_4777);
xnor U8861 (N_8861,N_240,N_318);
xor U8862 (N_8862,N_2436,N_4832);
or U8863 (N_8863,N_224,N_1101);
and U8864 (N_8864,N_3531,N_1562);
and U8865 (N_8865,N_2850,N_2590);
xor U8866 (N_8866,N_1516,N_3636);
or U8867 (N_8867,N_3819,N_4901);
and U8868 (N_8868,N_1104,N_694);
xnor U8869 (N_8869,N_2034,N_1235);
nand U8870 (N_8870,N_1338,N_4542);
and U8871 (N_8871,N_4415,N_4899);
xor U8872 (N_8872,N_2556,N_1977);
nor U8873 (N_8873,N_806,N_3034);
or U8874 (N_8874,N_249,N_1511);
xnor U8875 (N_8875,N_2729,N_3389);
and U8876 (N_8876,N_4182,N_3537);
or U8877 (N_8877,N_11,N_2456);
nor U8878 (N_8878,N_2530,N_1523);
and U8879 (N_8879,N_4020,N_4301);
nor U8880 (N_8880,N_4266,N_4282);
nor U8881 (N_8881,N_1727,N_4152);
nor U8882 (N_8882,N_3110,N_1924);
or U8883 (N_8883,N_1228,N_4217);
or U8884 (N_8884,N_3764,N_3714);
or U8885 (N_8885,N_942,N_2956);
and U8886 (N_8886,N_856,N_4457);
or U8887 (N_8887,N_2721,N_142);
and U8888 (N_8888,N_3112,N_2110);
xnor U8889 (N_8889,N_3456,N_2771);
nand U8890 (N_8890,N_2948,N_1711);
nand U8891 (N_8891,N_1808,N_3218);
or U8892 (N_8892,N_3716,N_4399);
and U8893 (N_8893,N_4337,N_3281);
xor U8894 (N_8894,N_1387,N_1774);
or U8895 (N_8895,N_502,N_4791);
and U8896 (N_8896,N_2864,N_1738);
xor U8897 (N_8897,N_4065,N_4155);
xnor U8898 (N_8898,N_3028,N_209);
and U8899 (N_8899,N_3986,N_4886);
nand U8900 (N_8900,N_3300,N_245);
xor U8901 (N_8901,N_1068,N_3317);
or U8902 (N_8902,N_1229,N_807);
nor U8903 (N_8903,N_1780,N_184);
xnor U8904 (N_8904,N_4892,N_1870);
xor U8905 (N_8905,N_388,N_739);
xor U8906 (N_8906,N_583,N_3964);
and U8907 (N_8907,N_2678,N_2201);
xor U8908 (N_8908,N_3254,N_2072);
and U8909 (N_8909,N_1042,N_3191);
or U8910 (N_8910,N_1027,N_1992);
nor U8911 (N_8911,N_1157,N_3645);
nand U8912 (N_8912,N_3293,N_2694);
xnor U8913 (N_8913,N_687,N_4068);
nand U8914 (N_8914,N_1351,N_3047);
or U8915 (N_8915,N_1706,N_4540);
nand U8916 (N_8916,N_720,N_2436);
and U8917 (N_8917,N_3461,N_1987);
or U8918 (N_8918,N_472,N_3943);
xor U8919 (N_8919,N_2322,N_3056);
and U8920 (N_8920,N_3731,N_193);
and U8921 (N_8921,N_250,N_2414);
nand U8922 (N_8922,N_4235,N_4886);
nand U8923 (N_8923,N_2993,N_1849);
nand U8924 (N_8924,N_4852,N_3490);
or U8925 (N_8925,N_2389,N_1879);
nor U8926 (N_8926,N_4068,N_2573);
nand U8927 (N_8927,N_37,N_2904);
nor U8928 (N_8928,N_2256,N_2705);
nand U8929 (N_8929,N_1267,N_731);
xor U8930 (N_8930,N_4086,N_4934);
nor U8931 (N_8931,N_155,N_1886);
nor U8932 (N_8932,N_1408,N_2408);
nand U8933 (N_8933,N_530,N_3623);
and U8934 (N_8934,N_961,N_44);
nand U8935 (N_8935,N_2875,N_2260);
nand U8936 (N_8936,N_1077,N_2485);
xnor U8937 (N_8937,N_1700,N_783);
xnor U8938 (N_8938,N_2380,N_4637);
nand U8939 (N_8939,N_3689,N_2777);
or U8940 (N_8940,N_4783,N_4380);
nand U8941 (N_8941,N_2507,N_4706);
or U8942 (N_8942,N_993,N_1942);
xor U8943 (N_8943,N_2082,N_4961);
xnor U8944 (N_8944,N_3564,N_1597);
nor U8945 (N_8945,N_1942,N_4186);
or U8946 (N_8946,N_3066,N_4329);
nor U8947 (N_8947,N_3225,N_3692);
xor U8948 (N_8948,N_2781,N_3473);
or U8949 (N_8949,N_172,N_4853);
xor U8950 (N_8950,N_3626,N_4262);
xor U8951 (N_8951,N_3850,N_2022);
nand U8952 (N_8952,N_2696,N_2189);
nor U8953 (N_8953,N_3963,N_1208);
xor U8954 (N_8954,N_488,N_439);
nor U8955 (N_8955,N_585,N_1733);
and U8956 (N_8956,N_2466,N_528);
or U8957 (N_8957,N_3413,N_3663);
nand U8958 (N_8958,N_113,N_55);
and U8959 (N_8959,N_3710,N_4270);
or U8960 (N_8960,N_1630,N_313);
or U8961 (N_8961,N_2473,N_1681);
nand U8962 (N_8962,N_4935,N_4020);
or U8963 (N_8963,N_2492,N_416);
and U8964 (N_8964,N_3087,N_4591);
nand U8965 (N_8965,N_4597,N_4355);
xor U8966 (N_8966,N_3000,N_4726);
nor U8967 (N_8967,N_114,N_3543);
nor U8968 (N_8968,N_2149,N_4427);
or U8969 (N_8969,N_3443,N_936);
or U8970 (N_8970,N_3707,N_4864);
xor U8971 (N_8971,N_4596,N_3017);
nor U8972 (N_8972,N_4642,N_1087);
or U8973 (N_8973,N_4186,N_3770);
and U8974 (N_8974,N_3233,N_1523);
or U8975 (N_8975,N_2,N_1301);
xnor U8976 (N_8976,N_603,N_1996);
nand U8977 (N_8977,N_3615,N_865);
xnor U8978 (N_8978,N_1020,N_932);
or U8979 (N_8979,N_148,N_2988);
or U8980 (N_8980,N_1147,N_1252);
xor U8981 (N_8981,N_3910,N_4800);
nor U8982 (N_8982,N_2137,N_330);
xnor U8983 (N_8983,N_2546,N_4874);
and U8984 (N_8984,N_2356,N_4252);
nand U8985 (N_8985,N_3866,N_4116);
and U8986 (N_8986,N_3953,N_2897);
nor U8987 (N_8987,N_3928,N_3465);
xor U8988 (N_8988,N_3768,N_159);
nand U8989 (N_8989,N_3255,N_1338);
nor U8990 (N_8990,N_2877,N_3782);
or U8991 (N_8991,N_1996,N_4328);
nor U8992 (N_8992,N_4817,N_133);
xnor U8993 (N_8993,N_3079,N_4140);
nand U8994 (N_8994,N_783,N_4481);
nor U8995 (N_8995,N_2808,N_635);
nor U8996 (N_8996,N_2581,N_2644);
and U8997 (N_8997,N_4713,N_3975);
and U8998 (N_8998,N_1118,N_4478);
nor U8999 (N_8999,N_3045,N_2072);
nand U9000 (N_9000,N_140,N_1287);
or U9001 (N_9001,N_3345,N_497);
nand U9002 (N_9002,N_1823,N_1818);
and U9003 (N_9003,N_2777,N_297);
or U9004 (N_9004,N_471,N_2035);
or U9005 (N_9005,N_3124,N_4073);
and U9006 (N_9006,N_4890,N_3758);
nor U9007 (N_9007,N_2854,N_867);
nand U9008 (N_9008,N_2870,N_563);
or U9009 (N_9009,N_625,N_4546);
and U9010 (N_9010,N_10,N_1255);
nor U9011 (N_9011,N_125,N_2555);
xor U9012 (N_9012,N_2845,N_877);
xor U9013 (N_9013,N_2928,N_1813);
and U9014 (N_9014,N_4721,N_1624);
xor U9015 (N_9015,N_2060,N_4909);
or U9016 (N_9016,N_4207,N_902);
xor U9017 (N_9017,N_3914,N_277);
and U9018 (N_9018,N_1834,N_2013);
xor U9019 (N_9019,N_977,N_2733);
or U9020 (N_9020,N_4191,N_1026);
nor U9021 (N_9021,N_1468,N_902);
nor U9022 (N_9022,N_3848,N_2559);
nand U9023 (N_9023,N_2812,N_499);
or U9024 (N_9024,N_602,N_1578);
and U9025 (N_9025,N_4826,N_889);
nor U9026 (N_9026,N_4655,N_191);
nand U9027 (N_9027,N_3995,N_4969);
nand U9028 (N_9028,N_1000,N_2843);
xnor U9029 (N_9029,N_2741,N_3205);
and U9030 (N_9030,N_4678,N_1112);
nor U9031 (N_9031,N_1872,N_3063);
and U9032 (N_9032,N_1341,N_1310);
nand U9033 (N_9033,N_3021,N_1306);
nor U9034 (N_9034,N_905,N_912);
nand U9035 (N_9035,N_2156,N_4259);
nand U9036 (N_9036,N_4658,N_4815);
or U9037 (N_9037,N_4382,N_47);
or U9038 (N_9038,N_1705,N_3142);
and U9039 (N_9039,N_1642,N_4124);
xor U9040 (N_9040,N_3391,N_4462);
and U9041 (N_9041,N_2413,N_3742);
nand U9042 (N_9042,N_4858,N_4756);
or U9043 (N_9043,N_122,N_2403);
nand U9044 (N_9044,N_579,N_3124);
and U9045 (N_9045,N_2816,N_217);
nor U9046 (N_9046,N_2697,N_193);
nor U9047 (N_9047,N_4465,N_3961);
nand U9048 (N_9048,N_3749,N_3292);
xnor U9049 (N_9049,N_2439,N_2639);
nor U9050 (N_9050,N_617,N_3716);
or U9051 (N_9051,N_3086,N_4998);
nand U9052 (N_9052,N_1507,N_1189);
xnor U9053 (N_9053,N_2850,N_3549);
nand U9054 (N_9054,N_4455,N_2301);
nand U9055 (N_9055,N_127,N_2799);
nor U9056 (N_9056,N_2990,N_672);
xnor U9057 (N_9057,N_745,N_4809);
nand U9058 (N_9058,N_1446,N_2207);
nor U9059 (N_9059,N_2128,N_1483);
nor U9060 (N_9060,N_3489,N_2862);
and U9061 (N_9061,N_601,N_3404);
xnor U9062 (N_9062,N_4020,N_4923);
and U9063 (N_9063,N_4329,N_3450);
and U9064 (N_9064,N_1556,N_1997);
or U9065 (N_9065,N_514,N_3904);
and U9066 (N_9066,N_3631,N_1184);
or U9067 (N_9067,N_2704,N_501);
and U9068 (N_9068,N_497,N_2703);
or U9069 (N_9069,N_1615,N_4290);
nor U9070 (N_9070,N_3714,N_1294);
nand U9071 (N_9071,N_681,N_2053);
and U9072 (N_9072,N_1296,N_3433);
nor U9073 (N_9073,N_373,N_1742);
nand U9074 (N_9074,N_2241,N_3188);
or U9075 (N_9075,N_803,N_1386);
or U9076 (N_9076,N_2077,N_49);
and U9077 (N_9077,N_1043,N_1689);
nor U9078 (N_9078,N_1534,N_500);
or U9079 (N_9079,N_1759,N_1511);
and U9080 (N_9080,N_2045,N_3521);
nor U9081 (N_9081,N_2295,N_3913);
or U9082 (N_9082,N_1365,N_2193);
nand U9083 (N_9083,N_2449,N_2280);
nor U9084 (N_9084,N_2642,N_2573);
nor U9085 (N_9085,N_370,N_3152);
nand U9086 (N_9086,N_3843,N_4900);
and U9087 (N_9087,N_4415,N_3959);
nand U9088 (N_9088,N_409,N_3412);
or U9089 (N_9089,N_2714,N_422);
xor U9090 (N_9090,N_4000,N_4788);
xor U9091 (N_9091,N_3286,N_2948);
nor U9092 (N_9092,N_1517,N_4);
nor U9093 (N_9093,N_3411,N_4779);
nand U9094 (N_9094,N_501,N_3318);
or U9095 (N_9095,N_736,N_3456);
and U9096 (N_9096,N_2005,N_808);
nand U9097 (N_9097,N_3536,N_3111);
nand U9098 (N_9098,N_2376,N_3521);
and U9099 (N_9099,N_296,N_677);
or U9100 (N_9100,N_903,N_4096);
nand U9101 (N_9101,N_4886,N_2193);
nor U9102 (N_9102,N_1565,N_3594);
or U9103 (N_9103,N_2706,N_1722);
or U9104 (N_9104,N_44,N_128);
nor U9105 (N_9105,N_3116,N_4485);
nor U9106 (N_9106,N_3997,N_548);
xnor U9107 (N_9107,N_1676,N_3681);
xnor U9108 (N_9108,N_3216,N_313);
or U9109 (N_9109,N_171,N_1766);
or U9110 (N_9110,N_1807,N_2950);
and U9111 (N_9111,N_3532,N_3443);
and U9112 (N_9112,N_434,N_2666);
nor U9113 (N_9113,N_3777,N_4264);
xor U9114 (N_9114,N_2017,N_2859);
xor U9115 (N_9115,N_4073,N_491);
nand U9116 (N_9116,N_1443,N_4781);
and U9117 (N_9117,N_1296,N_1748);
or U9118 (N_9118,N_2201,N_4590);
nand U9119 (N_9119,N_245,N_2105);
xnor U9120 (N_9120,N_4108,N_1449);
or U9121 (N_9121,N_3908,N_2889);
and U9122 (N_9122,N_166,N_3987);
nand U9123 (N_9123,N_2109,N_2021);
and U9124 (N_9124,N_2964,N_742);
xor U9125 (N_9125,N_762,N_4766);
or U9126 (N_9126,N_2578,N_3063);
nor U9127 (N_9127,N_4619,N_4041);
xor U9128 (N_9128,N_4385,N_1367);
nor U9129 (N_9129,N_1179,N_1478);
nor U9130 (N_9130,N_4959,N_4883);
or U9131 (N_9131,N_4466,N_126);
nand U9132 (N_9132,N_1015,N_1624);
nand U9133 (N_9133,N_109,N_1232);
nand U9134 (N_9134,N_3176,N_2140);
nor U9135 (N_9135,N_1211,N_4408);
and U9136 (N_9136,N_3899,N_1649);
or U9137 (N_9137,N_1128,N_1722);
or U9138 (N_9138,N_4859,N_1976);
nor U9139 (N_9139,N_3680,N_4434);
or U9140 (N_9140,N_1894,N_3323);
or U9141 (N_9141,N_145,N_3873);
and U9142 (N_9142,N_4520,N_4323);
and U9143 (N_9143,N_3889,N_1259);
and U9144 (N_9144,N_832,N_4508);
nor U9145 (N_9145,N_3653,N_4062);
nand U9146 (N_9146,N_1207,N_3236);
nor U9147 (N_9147,N_1572,N_3445);
nor U9148 (N_9148,N_4616,N_4254);
and U9149 (N_9149,N_3536,N_374);
nand U9150 (N_9150,N_4962,N_2523);
and U9151 (N_9151,N_839,N_2219);
xor U9152 (N_9152,N_343,N_811);
nand U9153 (N_9153,N_3073,N_4067);
xor U9154 (N_9154,N_4831,N_899);
nor U9155 (N_9155,N_3269,N_4167);
nor U9156 (N_9156,N_1331,N_4905);
nand U9157 (N_9157,N_1969,N_1130);
xnor U9158 (N_9158,N_185,N_2869);
and U9159 (N_9159,N_3708,N_3636);
or U9160 (N_9160,N_2082,N_1103);
nand U9161 (N_9161,N_4222,N_3307);
xor U9162 (N_9162,N_2696,N_2455);
nor U9163 (N_9163,N_1934,N_1809);
xor U9164 (N_9164,N_1082,N_4322);
and U9165 (N_9165,N_422,N_1216);
and U9166 (N_9166,N_542,N_956);
nor U9167 (N_9167,N_1019,N_4943);
and U9168 (N_9168,N_3446,N_1390);
nor U9169 (N_9169,N_4811,N_3861);
and U9170 (N_9170,N_1604,N_2228);
and U9171 (N_9171,N_578,N_3481);
nor U9172 (N_9172,N_4939,N_3666);
nand U9173 (N_9173,N_1370,N_1581);
xor U9174 (N_9174,N_3372,N_3594);
and U9175 (N_9175,N_3895,N_3662);
nor U9176 (N_9176,N_4374,N_2961);
nor U9177 (N_9177,N_3044,N_1940);
or U9178 (N_9178,N_360,N_1982);
or U9179 (N_9179,N_3074,N_3301);
and U9180 (N_9180,N_4216,N_3035);
xnor U9181 (N_9181,N_4715,N_466);
and U9182 (N_9182,N_1347,N_3063);
nor U9183 (N_9183,N_3634,N_255);
nor U9184 (N_9184,N_655,N_2673);
nand U9185 (N_9185,N_1829,N_4673);
or U9186 (N_9186,N_4750,N_4715);
nor U9187 (N_9187,N_3012,N_1890);
or U9188 (N_9188,N_2612,N_2389);
nor U9189 (N_9189,N_4318,N_4333);
or U9190 (N_9190,N_2357,N_4092);
and U9191 (N_9191,N_2460,N_987);
xor U9192 (N_9192,N_4172,N_4821);
nor U9193 (N_9193,N_920,N_2392);
and U9194 (N_9194,N_3022,N_298);
nor U9195 (N_9195,N_4425,N_1582);
xnor U9196 (N_9196,N_139,N_1258);
or U9197 (N_9197,N_4572,N_4008);
nand U9198 (N_9198,N_1356,N_4203);
xor U9199 (N_9199,N_1239,N_1634);
xor U9200 (N_9200,N_233,N_69);
nand U9201 (N_9201,N_4463,N_1216);
nor U9202 (N_9202,N_238,N_1988);
nor U9203 (N_9203,N_1806,N_4395);
or U9204 (N_9204,N_3141,N_4583);
or U9205 (N_9205,N_250,N_1640);
nor U9206 (N_9206,N_2202,N_2032);
or U9207 (N_9207,N_1246,N_3233);
and U9208 (N_9208,N_1048,N_366);
or U9209 (N_9209,N_4186,N_1218);
nand U9210 (N_9210,N_153,N_392);
xor U9211 (N_9211,N_51,N_1720);
nor U9212 (N_9212,N_4544,N_1490);
or U9213 (N_9213,N_1135,N_1246);
nand U9214 (N_9214,N_549,N_1134);
or U9215 (N_9215,N_4107,N_1966);
xor U9216 (N_9216,N_143,N_2477);
nor U9217 (N_9217,N_3125,N_2256);
xnor U9218 (N_9218,N_2764,N_1832);
nand U9219 (N_9219,N_2315,N_2054);
or U9220 (N_9220,N_4801,N_4232);
nand U9221 (N_9221,N_3804,N_4803);
and U9222 (N_9222,N_1198,N_4650);
nand U9223 (N_9223,N_4081,N_3551);
nor U9224 (N_9224,N_1949,N_1708);
or U9225 (N_9225,N_3330,N_326);
nor U9226 (N_9226,N_1228,N_2035);
xnor U9227 (N_9227,N_3146,N_4198);
or U9228 (N_9228,N_103,N_1870);
nor U9229 (N_9229,N_3779,N_1930);
and U9230 (N_9230,N_334,N_4841);
and U9231 (N_9231,N_438,N_4852);
and U9232 (N_9232,N_1506,N_2503);
nor U9233 (N_9233,N_655,N_1334);
nand U9234 (N_9234,N_2810,N_3225);
xor U9235 (N_9235,N_594,N_3653);
or U9236 (N_9236,N_4665,N_2959);
nor U9237 (N_9237,N_2856,N_3624);
nor U9238 (N_9238,N_3639,N_1534);
and U9239 (N_9239,N_697,N_1155);
nor U9240 (N_9240,N_3230,N_2965);
xnor U9241 (N_9241,N_2182,N_307);
or U9242 (N_9242,N_748,N_4730);
and U9243 (N_9243,N_21,N_485);
nand U9244 (N_9244,N_4193,N_2270);
or U9245 (N_9245,N_2633,N_378);
nor U9246 (N_9246,N_1505,N_596);
nand U9247 (N_9247,N_1868,N_3635);
and U9248 (N_9248,N_2916,N_2277);
nor U9249 (N_9249,N_3,N_4646);
nor U9250 (N_9250,N_855,N_3816);
or U9251 (N_9251,N_4608,N_3962);
nor U9252 (N_9252,N_1997,N_2539);
nand U9253 (N_9253,N_2306,N_3639);
nand U9254 (N_9254,N_2249,N_1204);
nor U9255 (N_9255,N_1603,N_2862);
or U9256 (N_9256,N_2377,N_854);
nor U9257 (N_9257,N_4665,N_2628);
or U9258 (N_9258,N_1177,N_1468);
nor U9259 (N_9259,N_3156,N_971);
and U9260 (N_9260,N_1328,N_907);
and U9261 (N_9261,N_4361,N_4285);
or U9262 (N_9262,N_2084,N_1598);
or U9263 (N_9263,N_4818,N_3612);
xnor U9264 (N_9264,N_4118,N_2536);
or U9265 (N_9265,N_172,N_3389);
or U9266 (N_9266,N_1100,N_2768);
nor U9267 (N_9267,N_868,N_184);
nand U9268 (N_9268,N_1164,N_1555);
xnor U9269 (N_9269,N_205,N_4916);
and U9270 (N_9270,N_3156,N_2733);
nor U9271 (N_9271,N_2531,N_4309);
nand U9272 (N_9272,N_3172,N_582);
xor U9273 (N_9273,N_4866,N_408);
and U9274 (N_9274,N_4264,N_3765);
xor U9275 (N_9275,N_2492,N_2531);
xor U9276 (N_9276,N_4391,N_1923);
nand U9277 (N_9277,N_478,N_3927);
nor U9278 (N_9278,N_2897,N_4002);
and U9279 (N_9279,N_1515,N_674);
xor U9280 (N_9280,N_3612,N_4808);
xnor U9281 (N_9281,N_4998,N_511);
and U9282 (N_9282,N_3824,N_4669);
nor U9283 (N_9283,N_426,N_1438);
or U9284 (N_9284,N_2922,N_3483);
or U9285 (N_9285,N_1502,N_1166);
nor U9286 (N_9286,N_1725,N_926);
xnor U9287 (N_9287,N_1223,N_3851);
nor U9288 (N_9288,N_2479,N_3697);
nand U9289 (N_9289,N_3403,N_3301);
xnor U9290 (N_9290,N_49,N_1985);
nand U9291 (N_9291,N_2810,N_2076);
or U9292 (N_9292,N_3243,N_2733);
and U9293 (N_9293,N_2605,N_225);
xnor U9294 (N_9294,N_169,N_811);
nand U9295 (N_9295,N_1710,N_3442);
nor U9296 (N_9296,N_900,N_1362);
nand U9297 (N_9297,N_3235,N_484);
or U9298 (N_9298,N_4499,N_3721);
or U9299 (N_9299,N_4998,N_4445);
and U9300 (N_9300,N_1410,N_4516);
xnor U9301 (N_9301,N_2829,N_777);
or U9302 (N_9302,N_4476,N_3586);
and U9303 (N_9303,N_1565,N_1795);
or U9304 (N_9304,N_408,N_573);
nor U9305 (N_9305,N_3902,N_3384);
and U9306 (N_9306,N_2106,N_3187);
and U9307 (N_9307,N_1947,N_4907);
nand U9308 (N_9308,N_3045,N_619);
nor U9309 (N_9309,N_160,N_863);
or U9310 (N_9310,N_2476,N_3839);
xor U9311 (N_9311,N_3770,N_4442);
nor U9312 (N_9312,N_4726,N_4568);
or U9313 (N_9313,N_4535,N_214);
and U9314 (N_9314,N_1026,N_3095);
xnor U9315 (N_9315,N_2030,N_2147);
or U9316 (N_9316,N_1991,N_4308);
nor U9317 (N_9317,N_892,N_1415);
nand U9318 (N_9318,N_2102,N_1801);
xor U9319 (N_9319,N_3686,N_1798);
nand U9320 (N_9320,N_3066,N_4902);
nand U9321 (N_9321,N_4864,N_4135);
or U9322 (N_9322,N_2718,N_334);
xnor U9323 (N_9323,N_3624,N_927);
or U9324 (N_9324,N_4637,N_1389);
or U9325 (N_9325,N_2094,N_2341);
nand U9326 (N_9326,N_3869,N_2113);
nor U9327 (N_9327,N_1818,N_2556);
and U9328 (N_9328,N_436,N_2409);
and U9329 (N_9329,N_4570,N_3069);
and U9330 (N_9330,N_116,N_671);
nor U9331 (N_9331,N_991,N_2348);
nand U9332 (N_9332,N_1322,N_2309);
or U9333 (N_9333,N_3317,N_4718);
nor U9334 (N_9334,N_1439,N_301);
nand U9335 (N_9335,N_1243,N_4228);
nor U9336 (N_9336,N_1118,N_2945);
or U9337 (N_9337,N_1919,N_3965);
xor U9338 (N_9338,N_2875,N_3852);
or U9339 (N_9339,N_4842,N_4901);
and U9340 (N_9340,N_1859,N_2282);
or U9341 (N_9341,N_1200,N_83);
or U9342 (N_9342,N_1415,N_1735);
or U9343 (N_9343,N_1278,N_96);
nor U9344 (N_9344,N_244,N_4629);
xnor U9345 (N_9345,N_4471,N_4200);
nand U9346 (N_9346,N_1623,N_3909);
nand U9347 (N_9347,N_747,N_306);
nand U9348 (N_9348,N_2924,N_4486);
and U9349 (N_9349,N_2071,N_4521);
or U9350 (N_9350,N_1155,N_1731);
nor U9351 (N_9351,N_4906,N_1109);
xnor U9352 (N_9352,N_3854,N_1894);
nand U9353 (N_9353,N_873,N_2856);
and U9354 (N_9354,N_865,N_551);
nor U9355 (N_9355,N_3883,N_2701);
xnor U9356 (N_9356,N_470,N_18);
nand U9357 (N_9357,N_3313,N_1239);
nor U9358 (N_9358,N_1566,N_3900);
xor U9359 (N_9359,N_4891,N_3988);
xor U9360 (N_9360,N_4256,N_2682);
and U9361 (N_9361,N_4909,N_3909);
xnor U9362 (N_9362,N_1333,N_4402);
nand U9363 (N_9363,N_2625,N_2022);
or U9364 (N_9364,N_1635,N_3327);
nand U9365 (N_9365,N_4893,N_4725);
or U9366 (N_9366,N_4289,N_1610);
nor U9367 (N_9367,N_847,N_3041);
nor U9368 (N_9368,N_2539,N_2946);
xnor U9369 (N_9369,N_1322,N_4279);
and U9370 (N_9370,N_4554,N_2226);
xnor U9371 (N_9371,N_4758,N_2905);
nand U9372 (N_9372,N_2968,N_3244);
nor U9373 (N_9373,N_4191,N_3244);
nand U9374 (N_9374,N_3507,N_2061);
or U9375 (N_9375,N_3220,N_2453);
and U9376 (N_9376,N_3230,N_3340);
and U9377 (N_9377,N_447,N_4846);
xnor U9378 (N_9378,N_773,N_4121);
nand U9379 (N_9379,N_930,N_1394);
xor U9380 (N_9380,N_944,N_4783);
and U9381 (N_9381,N_4405,N_2962);
and U9382 (N_9382,N_3497,N_4522);
xor U9383 (N_9383,N_4637,N_3699);
nand U9384 (N_9384,N_1706,N_3156);
nor U9385 (N_9385,N_2875,N_1162);
and U9386 (N_9386,N_423,N_4609);
nor U9387 (N_9387,N_1121,N_4359);
nand U9388 (N_9388,N_1292,N_360);
xnor U9389 (N_9389,N_2911,N_3555);
xor U9390 (N_9390,N_4735,N_4945);
nor U9391 (N_9391,N_3622,N_483);
and U9392 (N_9392,N_746,N_1536);
nor U9393 (N_9393,N_2662,N_2980);
nor U9394 (N_9394,N_3230,N_2403);
and U9395 (N_9395,N_2537,N_3354);
and U9396 (N_9396,N_2888,N_968);
and U9397 (N_9397,N_2121,N_2797);
xor U9398 (N_9398,N_4152,N_2847);
nand U9399 (N_9399,N_3680,N_2610);
xor U9400 (N_9400,N_289,N_2602);
nor U9401 (N_9401,N_118,N_2192);
nand U9402 (N_9402,N_874,N_1126);
nor U9403 (N_9403,N_4604,N_2588);
and U9404 (N_9404,N_3260,N_494);
nand U9405 (N_9405,N_811,N_1597);
nand U9406 (N_9406,N_2801,N_1462);
and U9407 (N_9407,N_4242,N_937);
nor U9408 (N_9408,N_3443,N_242);
xnor U9409 (N_9409,N_1168,N_3318);
nor U9410 (N_9410,N_2635,N_12);
and U9411 (N_9411,N_4269,N_1392);
nor U9412 (N_9412,N_4289,N_1533);
and U9413 (N_9413,N_4910,N_1619);
and U9414 (N_9414,N_2902,N_3651);
xor U9415 (N_9415,N_1568,N_3729);
or U9416 (N_9416,N_2342,N_17);
xor U9417 (N_9417,N_4896,N_1100);
xor U9418 (N_9418,N_2709,N_1402);
and U9419 (N_9419,N_2059,N_4974);
nand U9420 (N_9420,N_3003,N_3793);
or U9421 (N_9421,N_2429,N_2427);
nor U9422 (N_9422,N_4652,N_2458);
nor U9423 (N_9423,N_3426,N_569);
and U9424 (N_9424,N_3837,N_4034);
nand U9425 (N_9425,N_1022,N_4340);
or U9426 (N_9426,N_3538,N_1683);
nand U9427 (N_9427,N_2440,N_2342);
or U9428 (N_9428,N_4920,N_2761);
nor U9429 (N_9429,N_1752,N_3414);
xor U9430 (N_9430,N_586,N_4025);
nand U9431 (N_9431,N_3716,N_4615);
and U9432 (N_9432,N_2288,N_2292);
nand U9433 (N_9433,N_3950,N_4879);
and U9434 (N_9434,N_2509,N_212);
nand U9435 (N_9435,N_1144,N_267);
or U9436 (N_9436,N_1485,N_1906);
xnor U9437 (N_9437,N_2502,N_794);
nand U9438 (N_9438,N_3252,N_3018);
xor U9439 (N_9439,N_548,N_1945);
xor U9440 (N_9440,N_3853,N_748);
xnor U9441 (N_9441,N_3087,N_3258);
nand U9442 (N_9442,N_3835,N_4322);
and U9443 (N_9443,N_3096,N_4916);
nand U9444 (N_9444,N_3236,N_3595);
nand U9445 (N_9445,N_3897,N_1980);
nor U9446 (N_9446,N_1914,N_2860);
nand U9447 (N_9447,N_4049,N_4792);
or U9448 (N_9448,N_1788,N_1657);
and U9449 (N_9449,N_3909,N_1627);
or U9450 (N_9450,N_2858,N_305);
nor U9451 (N_9451,N_1115,N_3777);
nand U9452 (N_9452,N_2613,N_3767);
and U9453 (N_9453,N_3511,N_2390);
or U9454 (N_9454,N_1143,N_4795);
nor U9455 (N_9455,N_4884,N_4614);
nand U9456 (N_9456,N_1770,N_3737);
and U9457 (N_9457,N_1009,N_1239);
nor U9458 (N_9458,N_139,N_2285);
and U9459 (N_9459,N_2540,N_2423);
nor U9460 (N_9460,N_2501,N_4930);
xor U9461 (N_9461,N_979,N_2081);
or U9462 (N_9462,N_3536,N_2453);
or U9463 (N_9463,N_3805,N_948);
nand U9464 (N_9464,N_2779,N_902);
xor U9465 (N_9465,N_2958,N_3521);
nand U9466 (N_9466,N_4043,N_2643);
xnor U9467 (N_9467,N_4781,N_282);
nor U9468 (N_9468,N_3993,N_359);
or U9469 (N_9469,N_4332,N_580);
or U9470 (N_9470,N_1339,N_2869);
xnor U9471 (N_9471,N_4164,N_3777);
nor U9472 (N_9472,N_3729,N_1766);
xor U9473 (N_9473,N_3604,N_1656);
nor U9474 (N_9474,N_3937,N_137);
xor U9475 (N_9475,N_4147,N_2540);
and U9476 (N_9476,N_822,N_774);
nor U9477 (N_9477,N_2376,N_3421);
or U9478 (N_9478,N_1979,N_4227);
and U9479 (N_9479,N_1757,N_1232);
nand U9480 (N_9480,N_4865,N_141);
nor U9481 (N_9481,N_2271,N_158);
nor U9482 (N_9482,N_3495,N_99);
nand U9483 (N_9483,N_2070,N_77);
and U9484 (N_9484,N_2942,N_3781);
nand U9485 (N_9485,N_4572,N_2423);
nand U9486 (N_9486,N_81,N_218);
xor U9487 (N_9487,N_709,N_2165);
xor U9488 (N_9488,N_4988,N_390);
xor U9489 (N_9489,N_341,N_3843);
or U9490 (N_9490,N_131,N_2419);
or U9491 (N_9491,N_2724,N_2254);
or U9492 (N_9492,N_831,N_4766);
xor U9493 (N_9493,N_1486,N_3840);
xor U9494 (N_9494,N_2837,N_4014);
nor U9495 (N_9495,N_1092,N_2704);
and U9496 (N_9496,N_4557,N_3038);
xnor U9497 (N_9497,N_3912,N_863);
xor U9498 (N_9498,N_4371,N_4314);
nor U9499 (N_9499,N_4185,N_2224);
nand U9500 (N_9500,N_1719,N_454);
or U9501 (N_9501,N_3524,N_2616);
nor U9502 (N_9502,N_4088,N_1412);
and U9503 (N_9503,N_720,N_3268);
nand U9504 (N_9504,N_3130,N_4235);
xor U9505 (N_9505,N_3783,N_1128);
nor U9506 (N_9506,N_761,N_1285);
and U9507 (N_9507,N_4855,N_37);
and U9508 (N_9508,N_4455,N_850);
nand U9509 (N_9509,N_4091,N_3663);
and U9510 (N_9510,N_2292,N_589);
nor U9511 (N_9511,N_737,N_2891);
nand U9512 (N_9512,N_1127,N_1478);
xnor U9513 (N_9513,N_2245,N_2253);
and U9514 (N_9514,N_4366,N_2752);
nor U9515 (N_9515,N_4644,N_1244);
xor U9516 (N_9516,N_3353,N_653);
nand U9517 (N_9517,N_2569,N_3430);
nand U9518 (N_9518,N_2710,N_3515);
nor U9519 (N_9519,N_1761,N_4804);
nor U9520 (N_9520,N_567,N_2613);
nand U9521 (N_9521,N_3602,N_4700);
nor U9522 (N_9522,N_939,N_3242);
or U9523 (N_9523,N_3730,N_4687);
xnor U9524 (N_9524,N_4729,N_1782);
and U9525 (N_9525,N_709,N_1113);
and U9526 (N_9526,N_2677,N_1197);
nand U9527 (N_9527,N_2953,N_1233);
nor U9528 (N_9528,N_579,N_1064);
and U9529 (N_9529,N_2206,N_2602);
nand U9530 (N_9530,N_2011,N_1307);
nand U9531 (N_9531,N_2385,N_791);
or U9532 (N_9532,N_3986,N_3700);
nand U9533 (N_9533,N_3200,N_3639);
xnor U9534 (N_9534,N_2510,N_4479);
nand U9535 (N_9535,N_1372,N_1482);
xor U9536 (N_9536,N_4237,N_3661);
nor U9537 (N_9537,N_4689,N_2375);
xor U9538 (N_9538,N_2868,N_2355);
or U9539 (N_9539,N_4606,N_4592);
xor U9540 (N_9540,N_3949,N_3599);
nor U9541 (N_9541,N_239,N_4302);
nor U9542 (N_9542,N_1601,N_4581);
and U9543 (N_9543,N_4740,N_1111);
or U9544 (N_9544,N_4446,N_3117);
xnor U9545 (N_9545,N_1889,N_2527);
and U9546 (N_9546,N_2022,N_662);
nor U9547 (N_9547,N_1493,N_890);
nand U9548 (N_9548,N_4154,N_4473);
and U9549 (N_9549,N_4398,N_2043);
nor U9550 (N_9550,N_4034,N_3761);
nor U9551 (N_9551,N_1438,N_893);
or U9552 (N_9552,N_4888,N_1783);
and U9553 (N_9553,N_3359,N_200);
nand U9554 (N_9554,N_2166,N_3353);
xnor U9555 (N_9555,N_839,N_4590);
or U9556 (N_9556,N_3512,N_3761);
nand U9557 (N_9557,N_2459,N_2328);
or U9558 (N_9558,N_2304,N_907);
nor U9559 (N_9559,N_2083,N_1471);
or U9560 (N_9560,N_4795,N_783);
xnor U9561 (N_9561,N_4849,N_734);
nor U9562 (N_9562,N_4971,N_3688);
nand U9563 (N_9563,N_4094,N_1024);
nand U9564 (N_9564,N_1838,N_1485);
or U9565 (N_9565,N_3464,N_1056);
or U9566 (N_9566,N_3333,N_3794);
nand U9567 (N_9567,N_3005,N_4899);
xor U9568 (N_9568,N_1858,N_1405);
nor U9569 (N_9569,N_4016,N_284);
or U9570 (N_9570,N_137,N_359);
nor U9571 (N_9571,N_394,N_829);
or U9572 (N_9572,N_2333,N_4737);
nor U9573 (N_9573,N_1323,N_2784);
and U9574 (N_9574,N_44,N_406);
xnor U9575 (N_9575,N_1230,N_4076);
or U9576 (N_9576,N_4764,N_4821);
nor U9577 (N_9577,N_4211,N_4351);
xor U9578 (N_9578,N_2261,N_2702);
and U9579 (N_9579,N_4018,N_947);
and U9580 (N_9580,N_2488,N_683);
nor U9581 (N_9581,N_4546,N_2199);
and U9582 (N_9582,N_3230,N_4581);
or U9583 (N_9583,N_438,N_2092);
or U9584 (N_9584,N_2263,N_1043);
nand U9585 (N_9585,N_3635,N_2758);
xor U9586 (N_9586,N_423,N_1875);
and U9587 (N_9587,N_2990,N_3433);
xnor U9588 (N_9588,N_2349,N_1925);
nor U9589 (N_9589,N_2363,N_565);
nor U9590 (N_9590,N_2064,N_3352);
xor U9591 (N_9591,N_3668,N_1692);
xnor U9592 (N_9592,N_1172,N_3084);
or U9593 (N_9593,N_1704,N_3905);
or U9594 (N_9594,N_1714,N_1394);
nor U9595 (N_9595,N_832,N_3601);
xnor U9596 (N_9596,N_4916,N_156);
nand U9597 (N_9597,N_996,N_2190);
xnor U9598 (N_9598,N_3605,N_1051);
nand U9599 (N_9599,N_3222,N_2661);
nor U9600 (N_9600,N_4693,N_1977);
or U9601 (N_9601,N_1323,N_2109);
and U9602 (N_9602,N_612,N_4048);
nor U9603 (N_9603,N_2393,N_4094);
xor U9604 (N_9604,N_3656,N_575);
xnor U9605 (N_9605,N_426,N_484);
and U9606 (N_9606,N_4384,N_4729);
xnor U9607 (N_9607,N_4613,N_2727);
or U9608 (N_9608,N_1412,N_4830);
nor U9609 (N_9609,N_2868,N_1718);
or U9610 (N_9610,N_238,N_176);
nor U9611 (N_9611,N_4698,N_1949);
or U9612 (N_9612,N_3676,N_4661);
and U9613 (N_9613,N_3136,N_4230);
xor U9614 (N_9614,N_3844,N_1468);
xor U9615 (N_9615,N_104,N_823);
nor U9616 (N_9616,N_565,N_416);
nor U9617 (N_9617,N_4323,N_3874);
or U9618 (N_9618,N_2300,N_296);
and U9619 (N_9619,N_1132,N_1487);
xor U9620 (N_9620,N_1426,N_2174);
or U9621 (N_9621,N_242,N_426);
nand U9622 (N_9622,N_2899,N_4701);
nor U9623 (N_9623,N_4304,N_3637);
or U9624 (N_9624,N_3901,N_2971);
or U9625 (N_9625,N_3959,N_4570);
xor U9626 (N_9626,N_931,N_849);
and U9627 (N_9627,N_1754,N_2306);
nor U9628 (N_9628,N_1715,N_1672);
xnor U9629 (N_9629,N_3053,N_4588);
nand U9630 (N_9630,N_3072,N_428);
and U9631 (N_9631,N_1547,N_2277);
nand U9632 (N_9632,N_1167,N_4913);
and U9633 (N_9633,N_4873,N_843);
and U9634 (N_9634,N_4277,N_4628);
or U9635 (N_9635,N_2523,N_850);
nor U9636 (N_9636,N_3367,N_2602);
or U9637 (N_9637,N_4256,N_2952);
xnor U9638 (N_9638,N_1685,N_2589);
xnor U9639 (N_9639,N_377,N_4812);
nor U9640 (N_9640,N_1780,N_3631);
and U9641 (N_9641,N_2940,N_1952);
xnor U9642 (N_9642,N_1257,N_1764);
nor U9643 (N_9643,N_4829,N_3602);
or U9644 (N_9644,N_4596,N_2522);
or U9645 (N_9645,N_3378,N_1277);
or U9646 (N_9646,N_4596,N_701);
or U9647 (N_9647,N_3445,N_350);
xor U9648 (N_9648,N_3079,N_1901);
and U9649 (N_9649,N_4553,N_3099);
nor U9650 (N_9650,N_806,N_730);
and U9651 (N_9651,N_2882,N_4169);
nor U9652 (N_9652,N_736,N_4232);
nor U9653 (N_9653,N_2688,N_2695);
xor U9654 (N_9654,N_4293,N_3123);
or U9655 (N_9655,N_606,N_4722);
or U9656 (N_9656,N_821,N_1998);
nor U9657 (N_9657,N_2768,N_224);
nor U9658 (N_9658,N_3521,N_1547);
nor U9659 (N_9659,N_3092,N_4611);
and U9660 (N_9660,N_1504,N_746);
nand U9661 (N_9661,N_3298,N_4464);
nor U9662 (N_9662,N_4576,N_4890);
or U9663 (N_9663,N_1611,N_3793);
and U9664 (N_9664,N_2641,N_677);
and U9665 (N_9665,N_4597,N_4933);
nand U9666 (N_9666,N_1059,N_3064);
nor U9667 (N_9667,N_2225,N_2667);
xor U9668 (N_9668,N_4682,N_4001);
and U9669 (N_9669,N_4924,N_4799);
nor U9670 (N_9670,N_3082,N_1246);
and U9671 (N_9671,N_193,N_1200);
xor U9672 (N_9672,N_354,N_795);
nand U9673 (N_9673,N_4197,N_2334);
nor U9674 (N_9674,N_3347,N_4622);
nand U9675 (N_9675,N_3407,N_1491);
or U9676 (N_9676,N_50,N_2775);
nand U9677 (N_9677,N_3184,N_4819);
and U9678 (N_9678,N_750,N_3520);
nor U9679 (N_9679,N_958,N_4820);
nor U9680 (N_9680,N_4100,N_3881);
or U9681 (N_9681,N_2728,N_4776);
nor U9682 (N_9682,N_4114,N_1287);
nor U9683 (N_9683,N_403,N_1903);
xor U9684 (N_9684,N_3800,N_1496);
nand U9685 (N_9685,N_3254,N_3484);
xnor U9686 (N_9686,N_1720,N_223);
xnor U9687 (N_9687,N_351,N_2798);
nand U9688 (N_9688,N_457,N_43);
or U9689 (N_9689,N_3959,N_2138);
nor U9690 (N_9690,N_2491,N_3384);
nand U9691 (N_9691,N_3559,N_3684);
xor U9692 (N_9692,N_3478,N_4531);
or U9693 (N_9693,N_1934,N_3617);
nor U9694 (N_9694,N_3186,N_4907);
or U9695 (N_9695,N_2736,N_3169);
nor U9696 (N_9696,N_1061,N_4987);
nor U9697 (N_9697,N_1822,N_3570);
nand U9698 (N_9698,N_2608,N_729);
and U9699 (N_9699,N_1446,N_4857);
nor U9700 (N_9700,N_1992,N_905);
or U9701 (N_9701,N_1983,N_851);
nand U9702 (N_9702,N_3085,N_1304);
xnor U9703 (N_9703,N_2649,N_850);
nor U9704 (N_9704,N_18,N_3137);
xnor U9705 (N_9705,N_4168,N_229);
nand U9706 (N_9706,N_4977,N_4609);
or U9707 (N_9707,N_172,N_1315);
and U9708 (N_9708,N_640,N_2996);
and U9709 (N_9709,N_486,N_3703);
xor U9710 (N_9710,N_4100,N_958);
and U9711 (N_9711,N_3830,N_4216);
and U9712 (N_9712,N_2921,N_695);
xor U9713 (N_9713,N_3780,N_87);
nand U9714 (N_9714,N_4343,N_4883);
nor U9715 (N_9715,N_3994,N_727);
nor U9716 (N_9716,N_1431,N_4456);
nand U9717 (N_9717,N_4681,N_4480);
and U9718 (N_9718,N_4028,N_1831);
xnor U9719 (N_9719,N_700,N_4244);
nand U9720 (N_9720,N_534,N_2986);
nand U9721 (N_9721,N_4579,N_1160);
nand U9722 (N_9722,N_1957,N_3077);
nor U9723 (N_9723,N_412,N_1173);
and U9724 (N_9724,N_2828,N_1193);
nand U9725 (N_9725,N_3117,N_1367);
xnor U9726 (N_9726,N_3143,N_2027);
or U9727 (N_9727,N_4769,N_1910);
xnor U9728 (N_9728,N_2151,N_1299);
and U9729 (N_9729,N_3542,N_1899);
or U9730 (N_9730,N_1851,N_3611);
nor U9731 (N_9731,N_3813,N_2524);
xnor U9732 (N_9732,N_2354,N_4639);
xor U9733 (N_9733,N_1520,N_4574);
and U9734 (N_9734,N_4976,N_2920);
nor U9735 (N_9735,N_1579,N_1188);
and U9736 (N_9736,N_849,N_954);
nand U9737 (N_9737,N_3125,N_4598);
or U9738 (N_9738,N_2008,N_4580);
nand U9739 (N_9739,N_1844,N_4122);
or U9740 (N_9740,N_509,N_1966);
or U9741 (N_9741,N_2941,N_4810);
or U9742 (N_9742,N_3006,N_329);
or U9743 (N_9743,N_2385,N_3237);
or U9744 (N_9744,N_3405,N_958);
and U9745 (N_9745,N_3378,N_859);
or U9746 (N_9746,N_84,N_3302);
xor U9747 (N_9747,N_2643,N_1730);
nor U9748 (N_9748,N_4073,N_1421);
or U9749 (N_9749,N_3182,N_2029);
and U9750 (N_9750,N_563,N_3447);
or U9751 (N_9751,N_1873,N_135);
or U9752 (N_9752,N_2739,N_2853);
and U9753 (N_9753,N_3187,N_3243);
and U9754 (N_9754,N_2286,N_4996);
nor U9755 (N_9755,N_798,N_4728);
nand U9756 (N_9756,N_4638,N_3511);
nand U9757 (N_9757,N_3355,N_3175);
and U9758 (N_9758,N_1074,N_4931);
and U9759 (N_9759,N_2262,N_3925);
xnor U9760 (N_9760,N_2505,N_1789);
xor U9761 (N_9761,N_2039,N_4819);
and U9762 (N_9762,N_3718,N_4582);
or U9763 (N_9763,N_3754,N_1901);
or U9764 (N_9764,N_2138,N_2229);
nand U9765 (N_9765,N_3872,N_4884);
and U9766 (N_9766,N_2045,N_1244);
or U9767 (N_9767,N_545,N_2457);
nor U9768 (N_9768,N_2334,N_1183);
and U9769 (N_9769,N_289,N_3871);
xor U9770 (N_9770,N_1748,N_3126);
nor U9771 (N_9771,N_3583,N_1258);
and U9772 (N_9772,N_1637,N_1642);
nand U9773 (N_9773,N_2536,N_2898);
and U9774 (N_9774,N_2889,N_486);
xnor U9775 (N_9775,N_610,N_612);
xnor U9776 (N_9776,N_1134,N_1425);
nand U9777 (N_9777,N_487,N_4611);
nand U9778 (N_9778,N_1160,N_2912);
and U9779 (N_9779,N_1742,N_4582);
nand U9780 (N_9780,N_4551,N_3369);
or U9781 (N_9781,N_2104,N_3668);
or U9782 (N_9782,N_2952,N_3730);
xnor U9783 (N_9783,N_1295,N_4143);
or U9784 (N_9784,N_2201,N_1839);
and U9785 (N_9785,N_1866,N_3984);
and U9786 (N_9786,N_3405,N_427);
and U9787 (N_9787,N_2157,N_4650);
and U9788 (N_9788,N_3814,N_1007);
or U9789 (N_9789,N_1913,N_1573);
nand U9790 (N_9790,N_4346,N_4012);
and U9791 (N_9791,N_4385,N_3210);
xnor U9792 (N_9792,N_2093,N_4785);
nand U9793 (N_9793,N_11,N_2180);
nand U9794 (N_9794,N_549,N_4248);
or U9795 (N_9795,N_2728,N_224);
and U9796 (N_9796,N_1142,N_3551);
nand U9797 (N_9797,N_1133,N_4905);
nor U9798 (N_9798,N_2737,N_3853);
and U9799 (N_9799,N_3583,N_2342);
xnor U9800 (N_9800,N_1534,N_2080);
or U9801 (N_9801,N_141,N_4357);
nor U9802 (N_9802,N_211,N_3784);
or U9803 (N_9803,N_4415,N_2482);
or U9804 (N_9804,N_2416,N_3832);
nand U9805 (N_9805,N_2525,N_4508);
nand U9806 (N_9806,N_1322,N_1094);
or U9807 (N_9807,N_1505,N_4006);
xnor U9808 (N_9808,N_4544,N_4874);
or U9809 (N_9809,N_2363,N_2250);
xnor U9810 (N_9810,N_285,N_40);
or U9811 (N_9811,N_1108,N_690);
nand U9812 (N_9812,N_1778,N_2380);
nand U9813 (N_9813,N_3264,N_1192);
or U9814 (N_9814,N_3860,N_2954);
xnor U9815 (N_9815,N_3367,N_2597);
nor U9816 (N_9816,N_3075,N_1667);
xnor U9817 (N_9817,N_1273,N_4286);
nor U9818 (N_9818,N_1114,N_4536);
xor U9819 (N_9819,N_523,N_3849);
and U9820 (N_9820,N_4556,N_4439);
nor U9821 (N_9821,N_569,N_3264);
or U9822 (N_9822,N_3874,N_2416);
xnor U9823 (N_9823,N_2681,N_3817);
nand U9824 (N_9824,N_474,N_186);
and U9825 (N_9825,N_1548,N_1536);
nor U9826 (N_9826,N_1450,N_4856);
or U9827 (N_9827,N_1544,N_2271);
nand U9828 (N_9828,N_4473,N_1884);
or U9829 (N_9829,N_7,N_161);
and U9830 (N_9830,N_699,N_1784);
xor U9831 (N_9831,N_3032,N_3402);
nand U9832 (N_9832,N_1511,N_262);
or U9833 (N_9833,N_2805,N_4747);
and U9834 (N_9834,N_3245,N_4892);
or U9835 (N_9835,N_4194,N_3375);
and U9836 (N_9836,N_2649,N_4185);
xnor U9837 (N_9837,N_1094,N_3435);
xnor U9838 (N_9838,N_1710,N_3284);
xor U9839 (N_9839,N_1283,N_1745);
nand U9840 (N_9840,N_3779,N_4815);
nand U9841 (N_9841,N_1343,N_391);
or U9842 (N_9842,N_63,N_2841);
and U9843 (N_9843,N_4611,N_1648);
xnor U9844 (N_9844,N_425,N_217);
or U9845 (N_9845,N_3153,N_502);
nand U9846 (N_9846,N_4206,N_2694);
or U9847 (N_9847,N_3264,N_38);
or U9848 (N_9848,N_1558,N_788);
nor U9849 (N_9849,N_2208,N_1804);
xor U9850 (N_9850,N_3439,N_2585);
and U9851 (N_9851,N_2072,N_4520);
xor U9852 (N_9852,N_3053,N_3940);
nand U9853 (N_9853,N_989,N_1575);
nand U9854 (N_9854,N_2693,N_2252);
and U9855 (N_9855,N_2557,N_1940);
and U9856 (N_9856,N_1228,N_4978);
xor U9857 (N_9857,N_4524,N_768);
xnor U9858 (N_9858,N_177,N_4100);
and U9859 (N_9859,N_3600,N_675);
nor U9860 (N_9860,N_3692,N_2758);
and U9861 (N_9861,N_2744,N_419);
and U9862 (N_9862,N_2998,N_1645);
nand U9863 (N_9863,N_4680,N_680);
and U9864 (N_9864,N_4884,N_1020);
nand U9865 (N_9865,N_1788,N_40);
and U9866 (N_9866,N_1568,N_3404);
and U9867 (N_9867,N_4618,N_2265);
or U9868 (N_9868,N_1550,N_1877);
nand U9869 (N_9869,N_4321,N_2438);
or U9870 (N_9870,N_4134,N_2990);
nor U9871 (N_9871,N_3052,N_4743);
or U9872 (N_9872,N_796,N_3368);
and U9873 (N_9873,N_2626,N_3776);
and U9874 (N_9874,N_882,N_4767);
nor U9875 (N_9875,N_3489,N_3411);
and U9876 (N_9876,N_2379,N_3569);
and U9877 (N_9877,N_3587,N_1228);
and U9878 (N_9878,N_4674,N_531);
nand U9879 (N_9879,N_1833,N_2942);
nor U9880 (N_9880,N_3980,N_574);
nand U9881 (N_9881,N_4775,N_715);
and U9882 (N_9882,N_514,N_3701);
nand U9883 (N_9883,N_2260,N_4615);
or U9884 (N_9884,N_2139,N_2907);
xnor U9885 (N_9885,N_442,N_1039);
nor U9886 (N_9886,N_2863,N_4475);
or U9887 (N_9887,N_2241,N_3929);
nand U9888 (N_9888,N_3634,N_3259);
nor U9889 (N_9889,N_4458,N_2420);
nand U9890 (N_9890,N_2003,N_509);
nand U9891 (N_9891,N_3323,N_2636);
nor U9892 (N_9892,N_3613,N_1865);
nor U9893 (N_9893,N_837,N_1960);
nor U9894 (N_9894,N_1021,N_1348);
and U9895 (N_9895,N_3601,N_4800);
and U9896 (N_9896,N_918,N_703);
nand U9897 (N_9897,N_1788,N_4600);
or U9898 (N_9898,N_1950,N_2849);
or U9899 (N_9899,N_80,N_3396);
and U9900 (N_9900,N_1477,N_3527);
nand U9901 (N_9901,N_3392,N_444);
and U9902 (N_9902,N_4321,N_4874);
or U9903 (N_9903,N_2915,N_1898);
and U9904 (N_9904,N_704,N_4263);
nand U9905 (N_9905,N_2339,N_4013);
and U9906 (N_9906,N_3595,N_2716);
and U9907 (N_9907,N_4538,N_4070);
and U9908 (N_9908,N_326,N_2764);
xor U9909 (N_9909,N_486,N_4154);
or U9910 (N_9910,N_797,N_4665);
or U9911 (N_9911,N_2370,N_4096);
nand U9912 (N_9912,N_932,N_3810);
or U9913 (N_9913,N_1575,N_3692);
nor U9914 (N_9914,N_4,N_3373);
nor U9915 (N_9915,N_3125,N_4525);
nand U9916 (N_9916,N_4664,N_4946);
or U9917 (N_9917,N_1902,N_1230);
nand U9918 (N_9918,N_1795,N_3986);
and U9919 (N_9919,N_4902,N_1310);
and U9920 (N_9920,N_3191,N_4623);
xor U9921 (N_9921,N_1136,N_4764);
nand U9922 (N_9922,N_4960,N_2999);
nand U9923 (N_9923,N_4550,N_1435);
or U9924 (N_9924,N_3729,N_1010);
nor U9925 (N_9925,N_1576,N_3916);
nor U9926 (N_9926,N_3585,N_1415);
and U9927 (N_9927,N_453,N_452);
and U9928 (N_9928,N_2317,N_3364);
xor U9929 (N_9929,N_1904,N_402);
or U9930 (N_9930,N_4593,N_1218);
or U9931 (N_9931,N_272,N_4850);
nand U9932 (N_9932,N_2174,N_512);
or U9933 (N_9933,N_1708,N_2055);
xor U9934 (N_9934,N_678,N_2488);
nor U9935 (N_9935,N_4794,N_1164);
nand U9936 (N_9936,N_4719,N_297);
xor U9937 (N_9937,N_1315,N_4997);
or U9938 (N_9938,N_4954,N_4493);
nor U9939 (N_9939,N_1717,N_1079);
and U9940 (N_9940,N_2076,N_189);
nor U9941 (N_9941,N_4518,N_2404);
xor U9942 (N_9942,N_978,N_3231);
and U9943 (N_9943,N_4259,N_3186);
nand U9944 (N_9944,N_2539,N_4537);
xnor U9945 (N_9945,N_1553,N_1061);
xnor U9946 (N_9946,N_4935,N_1082);
nor U9947 (N_9947,N_1314,N_4376);
nor U9948 (N_9948,N_3699,N_2494);
or U9949 (N_9949,N_4380,N_1667);
or U9950 (N_9950,N_1183,N_360);
xor U9951 (N_9951,N_162,N_4897);
xor U9952 (N_9952,N_4427,N_4130);
or U9953 (N_9953,N_877,N_3334);
and U9954 (N_9954,N_451,N_4056);
xor U9955 (N_9955,N_4471,N_1763);
or U9956 (N_9956,N_605,N_3685);
nor U9957 (N_9957,N_3116,N_4658);
xnor U9958 (N_9958,N_4887,N_2447);
and U9959 (N_9959,N_4113,N_3956);
xnor U9960 (N_9960,N_4939,N_2085);
nor U9961 (N_9961,N_119,N_2702);
xnor U9962 (N_9962,N_4235,N_2976);
and U9963 (N_9963,N_1263,N_957);
nor U9964 (N_9964,N_1887,N_3152);
or U9965 (N_9965,N_402,N_221);
nor U9966 (N_9966,N_4286,N_2906);
or U9967 (N_9967,N_3443,N_312);
or U9968 (N_9968,N_561,N_3927);
nand U9969 (N_9969,N_3391,N_769);
nand U9970 (N_9970,N_138,N_2489);
and U9971 (N_9971,N_4173,N_88);
or U9972 (N_9972,N_2843,N_2474);
nand U9973 (N_9973,N_1937,N_3381);
nand U9974 (N_9974,N_3847,N_3357);
and U9975 (N_9975,N_4391,N_242);
and U9976 (N_9976,N_1061,N_2035);
and U9977 (N_9977,N_827,N_265);
or U9978 (N_9978,N_2539,N_3916);
nand U9979 (N_9979,N_935,N_82);
nor U9980 (N_9980,N_103,N_1477);
and U9981 (N_9981,N_639,N_513);
and U9982 (N_9982,N_1566,N_1275);
nand U9983 (N_9983,N_2043,N_4016);
nand U9984 (N_9984,N_4833,N_3463);
nor U9985 (N_9985,N_2964,N_4766);
nand U9986 (N_9986,N_141,N_4414);
or U9987 (N_9987,N_1790,N_4287);
or U9988 (N_9988,N_1219,N_3580);
xnor U9989 (N_9989,N_3630,N_1019);
nor U9990 (N_9990,N_3526,N_1247);
and U9991 (N_9991,N_4664,N_1103);
nand U9992 (N_9992,N_947,N_909);
and U9993 (N_9993,N_3650,N_4589);
xnor U9994 (N_9994,N_603,N_1100);
and U9995 (N_9995,N_2303,N_4114);
nand U9996 (N_9996,N_763,N_4064);
nand U9997 (N_9997,N_1056,N_81);
and U9998 (N_9998,N_4107,N_2108);
nor U9999 (N_9999,N_4843,N_3781);
and UO_0 (O_0,N_7491,N_5822);
or UO_1 (O_1,N_5377,N_8822);
nand UO_2 (O_2,N_6660,N_9165);
nand UO_3 (O_3,N_7404,N_7100);
nor UO_4 (O_4,N_6458,N_5080);
nand UO_5 (O_5,N_8340,N_5921);
and UO_6 (O_6,N_6986,N_9238);
nand UO_7 (O_7,N_7048,N_7354);
and UO_8 (O_8,N_8211,N_9770);
xnor UO_9 (O_9,N_8953,N_8331);
xor UO_10 (O_10,N_9331,N_9949);
nor UO_11 (O_11,N_8086,N_6368);
xor UO_12 (O_12,N_6580,N_9071);
nor UO_13 (O_13,N_9609,N_8716);
or UO_14 (O_14,N_6569,N_9135);
and UO_15 (O_15,N_8568,N_7023);
xor UO_16 (O_16,N_7992,N_5067);
or UO_17 (O_17,N_6880,N_7334);
or UO_18 (O_18,N_8948,N_7996);
nand UO_19 (O_19,N_5324,N_7041);
nor UO_20 (O_20,N_9481,N_7359);
xor UO_21 (O_21,N_8563,N_8096);
xnor UO_22 (O_22,N_6198,N_5084);
xor UO_23 (O_23,N_6129,N_7378);
or UO_24 (O_24,N_5985,N_8532);
or UO_25 (O_25,N_7074,N_9838);
and UO_26 (O_26,N_9439,N_7292);
xnor UO_27 (O_27,N_7667,N_6445);
nand UO_28 (O_28,N_9551,N_5969);
or UO_29 (O_29,N_8961,N_7436);
and UO_30 (O_30,N_6517,N_5480);
xor UO_31 (O_31,N_7202,N_7165);
and UO_32 (O_32,N_8482,N_9700);
nand UO_33 (O_33,N_5479,N_5538);
and UO_34 (O_34,N_8681,N_6246);
or UO_35 (O_35,N_7123,N_6339);
or UO_36 (O_36,N_5651,N_6111);
nor UO_37 (O_37,N_8296,N_8533);
xnor UO_38 (O_38,N_8425,N_9529);
nand UO_39 (O_39,N_9448,N_6364);
or UO_40 (O_40,N_5580,N_5163);
and UO_41 (O_41,N_6542,N_8869);
nand UO_42 (O_42,N_6902,N_8417);
xor UO_43 (O_43,N_5903,N_7556);
xor UO_44 (O_44,N_8105,N_6725);
xor UO_45 (O_45,N_8255,N_9455);
and UO_46 (O_46,N_5059,N_6108);
and UO_47 (O_47,N_9421,N_6679);
and UO_48 (O_48,N_8945,N_7775);
or UO_49 (O_49,N_5607,N_6860);
or UO_50 (O_50,N_6003,N_9900);
nor UO_51 (O_51,N_7628,N_9022);
nand UO_52 (O_52,N_8384,N_8597);
and UO_53 (O_53,N_8079,N_6876);
xor UO_54 (O_54,N_5265,N_5924);
nand UO_55 (O_55,N_5487,N_6021);
xor UO_56 (O_56,N_7283,N_9161);
nor UO_57 (O_57,N_5795,N_9323);
nand UO_58 (O_58,N_5861,N_8808);
or UO_59 (O_59,N_6649,N_7559);
xnor UO_60 (O_60,N_6510,N_8844);
and UO_61 (O_61,N_9304,N_8438);
and UO_62 (O_62,N_5096,N_8672);
and UO_63 (O_63,N_6826,N_8906);
or UO_64 (O_64,N_6352,N_6016);
nand UO_65 (O_65,N_9756,N_8832);
or UO_66 (O_66,N_9419,N_6276);
or UO_67 (O_67,N_6544,N_8594);
or UO_68 (O_68,N_9681,N_8726);
xor UO_69 (O_69,N_5052,N_9658);
and UO_70 (O_70,N_6837,N_6599);
and UO_71 (O_71,N_6944,N_6162);
xnor UO_72 (O_72,N_8210,N_6655);
and UO_73 (O_73,N_9961,N_7546);
and UO_74 (O_74,N_5185,N_8101);
nand UO_75 (O_75,N_6567,N_5405);
nand UO_76 (O_76,N_6565,N_8898);
nor UO_77 (O_77,N_9833,N_7357);
nor UO_78 (O_78,N_9485,N_7510);
nor UO_79 (O_79,N_8846,N_6716);
nor UO_80 (O_80,N_7180,N_6728);
nand UO_81 (O_81,N_6365,N_5657);
and UO_82 (O_82,N_6997,N_9340);
nor UO_83 (O_83,N_7243,N_5991);
nand UO_84 (O_84,N_8629,N_6305);
and UO_85 (O_85,N_6832,N_8671);
xnor UO_86 (O_86,N_7710,N_9416);
and UO_87 (O_87,N_7274,N_7657);
nand UO_88 (O_88,N_7066,N_6605);
or UO_89 (O_89,N_5249,N_7050);
xnor UO_90 (O_90,N_5177,N_5264);
xnor UO_91 (O_91,N_7690,N_7679);
or UO_92 (O_92,N_7248,N_6233);
and UO_93 (O_93,N_9823,N_9082);
or UO_94 (O_94,N_6402,N_5213);
and UO_95 (O_95,N_8003,N_7881);
xnor UO_96 (O_96,N_9830,N_8700);
or UO_97 (O_97,N_5642,N_6110);
nand UO_98 (O_98,N_5430,N_5963);
nor UO_99 (O_99,N_9192,N_9289);
or UO_100 (O_100,N_6887,N_9489);
or UO_101 (O_101,N_5227,N_6069);
nor UO_102 (O_102,N_6275,N_9755);
or UO_103 (O_103,N_6284,N_8656);
and UO_104 (O_104,N_6273,N_5415);
nand UO_105 (O_105,N_6055,N_8024);
xor UO_106 (O_106,N_7371,N_8029);
or UO_107 (O_107,N_7153,N_6718);
xnor UO_108 (O_108,N_5128,N_8374);
nand UO_109 (O_109,N_7383,N_8649);
nand UO_110 (O_110,N_6283,N_5863);
and UO_111 (O_111,N_8395,N_9167);
nand UO_112 (O_112,N_9213,N_7007);
or UO_113 (O_113,N_6504,N_9404);
nor UO_114 (O_114,N_9166,N_9328);
xnor UO_115 (O_115,N_7680,N_8880);
nor UO_116 (O_116,N_5803,N_9454);
nand UO_117 (O_117,N_6680,N_7964);
nor UO_118 (O_118,N_5228,N_5178);
and UO_119 (O_119,N_6636,N_6988);
nand UO_120 (O_120,N_5211,N_7024);
xor UO_121 (O_121,N_7316,N_6508);
nand UO_122 (O_122,N_5899,N_6023);
and UO_123 (O_123,N_5563,N_9270);
nor UO_124 (O_124,N_6318,N_8390);
xnor UO_125 (O_125,N_5073,N_6614);
nand UO_126 (O_126,N_5477,N_6755);
or UO_127 (O_127,N_9889,N_6644);
xnor UO_128 (O_128,N_8803,N_5910);
and UO_129 (O_129,N_8021,N_8461);
and UO_130 (O_130,N_6325,N_5194);
and UO_131 (O_131,N_8531,N_8062);
or UO_132 (O_132,N_8962,N_7224);
nand UO_133 (O_133,N_8475,N_6366);
and UO_134 (O_134,N_8058,N_9875);
xor UO_135 (O_135,N_9663,N_6072);
xor UO_136 (O_136,N_7476,N_7718);
nand UO_137 (O_137,N_9980,N_9730);
nor UO_138 (O_138,N_7837,N_6581);
nand UO_139 (O_139,N_6123,N_6376);
and UO_140 (O_140,N_8811,N_8717);
nand UO_141 (O_141,N_9133,N_5797);
xnor UO_142 (O_142,N_9036,N_5849);
nand UO_143 (O_143,N_5804,N_5455);
xor UO_144 (O_144,N_6439,N_9278);
nand UO_145 (O_145,N_9390,N_8366);
nand UO_146 (O_146,N_6178,N_8769);
nor UO_147 (O_147,N_8185,N_5782);
and UO_148 (O_148,N_6908,N_8462);
xnor UO_149 (O_149,N_5351,N_8666);
xor UO_150 (O_150,N_9447,N_5190);
and UO_151 (O_151,N_8715,N_9470);
nor UO_152 (O_152,N_6646,N_9850);
and UO_153 (O_153,N_5749,N_7502);
nor UO_154 (O_154,N_5644,N_9595);
or UO_155 (O_155,N_5353,N_7276);
nand UO_156 (O_156,N_7769,N_7126);
xor UO_157 (O_157,N_7926,N_8378);
or UO_158 (O_158,N_5337,N_5575);
or UO_159 (O_159,N_8827,N_9179);
or UO_160 (O_160,N_9468,N_5608);
xnor UO_161 (O_161,N_6747,N_9648);
and UO_162 (O_162,N_9661,N_7373);
or UO_163 (O_163,N_8966,N_7249);
nor UO_164 (O_164,N_5315,N_8860);
nor UO_165 (O_165,N_8895,N_5394);
or UO_166 (O_166,N_5775,N_6555);
xnor UO_167 (O_167,N_6289,N_9726);
and UO_168 (O_168,N_8712,N_7551);
nand UO_169 (O_169,N_5446,N_7712);
xor UO_170 (O_170,N_9637,N_8027);
xor UO_171 (O_171,N_8166,N_9533);
xnor UO_172 (O_172,N_5335,N_5202);
nor UO_173 (O_173,N_8491,N_9585);
or UO_174 (O_174,N_6813,N_6962);
xnor UO_175 (O_175,N_6589,N_7326);
nor UO_176 (O_176,N_8134,N_5103);
and UO_177 (O_177,N_7159,N_7227);
nand UO_178 (O_178,N_8249,N_8601);
xnor UO_179 (O_179,N_7372,N_7433);
and UO_180 (O_180,N_7856,N_8925);
nor UO_181 (O_181,N_7825,N_6480);
xor UO_182 (O_182,N_7445,N_6076);
nor UO_183 (O_183,N_5182,N_9043);
nand UO_184 (O_184,N_7393,N_8234);
nor UO_185 (O_185,N_5242,N_7259);
nor UO_186 (O_186,N_5902,N_6877);
nand UO_187 (O_187,N_9001,N_5197);
or UO_188 (O_188,N_5271,N_7079);
nor UO_189 (O_189,N_7238,N_5937);
xor UO_190 (O_190,N_8921,N_9079);
xnor UO_191 (O_191,N_9784,N_6241);
or UO_192 (O_192,N_6004,N_5340);
and UO_193 (O_193,N_7113,N_5938);
or UO_194 (O_194,N_9591,N_8085);
and UO_195 (O_195,N_7056,N_5320);
nand UO_196 (O_196,N_5133,N_9651);
xor UO_197 (O_197,N_5681,N_9189);
and UO_198 (O_198,N_9397,N_9400);
xnor UO_199 (O_199,N_9907,N_6541);
and UO_200 (O_200,N_6929,N_6691);
nand UO_201 (O_201,N_7797,N_6203);
or UO_202 (O_202,N_8509,N_7446);
nand UO_203 (O_203,N_9157,N_7658);
nor UO_204 (O_204,N_6562,N_7924);
nand UO_205 (O_205,N_6503,N_5138);
nor UO_206 (O_206,N_9228,N_9575);
or UO_207 (O_207,N_6613,N_8406);
nand UO_208 (O_208,N_7405,N_5208);
or UO_209 (O_209,N_5541,N_6191);
and UO_210 (O_210,N_7652,N_8454);
xor UO_211 (O_211,N_7970,N_7443);
xnor UO_212 (O_212,N_7432,N_8675);
nor UO_213 (O_213,N_8753,N_6668);
xnor UO_214 (O_214,N_5166,N_9062);
nand UO_215 (O_215,N_7668,N_7196);
nand UO_216 (O_216,N_5892,N_8773);
nand UO_217 (O_217,N_7342,N_8534);
xor UO_218 (O_218,N_6999,N_6166);
and UO_219 (O_219,N_7329,N_5475);
and UO_220 (O_220,N_6782,N_9955);
xnor UO_221 (O_221,N_5702,N_5582);
or UO_222 (O_222,N_8289,N_6073);
and UO_223 (O_223,N_7175,N_7246);
nand UO_224 (O_224,N_5734,N_5019);
nor UO_225 (O_225,N_8645,N_7469);
nand UO_226 (O_226,N_6847,N_9703);
or UO_227 (O_227,N_9232,N_5342);
xnor UO_228 (O_228,N_5186,N_9993);
and UO_229 (O_229,N_8152,N_6874);
nor UO_230 (O_230,N_8548,N_7385);
xnor UO_231 (O_231,N_9796,N_9965);
nand UO_232 (O_232,N_6026,N_5508);
nor UO_233 (O_233,N_5445,N_9910);
nor UO_234 (O_234,N_8008,N_7218);
xnor UO_235 (O_235,N_7633,N_8588);
and UO_236 (O_236,N_6735,N_8908);
or UO_237 (O_237,N_5896,N_9716);
and UO_238 (O_238,N_8522,N_5788);
and UO_239 (O_239,N_5281,N_9386);
nand UO_240 (O_240,N_6617,N_7968);
or UO_241 (O_241,N_6978,N_6309);
nor UO_242 (O_242,N_7273,N_8269);
nor UO_243 (O_243,N_6709,N_5267);
or UO_244 (O_244,N_9361,N_5998);
xnor UO_245 (O_245,N_5539,N_7823);
xnor UO_246 (O_246,N_7872,N_6615);
xnor UO_247 (O_247,N_5677,N_5365);
nand UO_248 (O_248,N_9476,N_9208);
nand UO_249 (O_249,N_8922,N_9747);
and UO_250 (O_250,N_5021,N_5470);
nor UO_251 (O_251,N_7632,N_8212);
or UO_252 (O_252,N_5511,N_9868);
nor UO_253 (O_253,N_7197,N_6047);
xor UO_254 (O_254,N_7922,N_5906);
and UO_255 (O_255,N_7596,N_8812);
nand UO_256 (O_256,N_5278,N_9858);
nand UO_257 (O_257,N_6359,N_5319);
nand UO_258 (O_258,N_7729,N_8957);
or UO_259 (O_259,N_6363,N_5196);
and UO_260 (O_260,N_5483,N_9911);
nand UO_261 (O_261,N_5950,N_7104);
or UO_262 (O_262,N_8574,N_6682);
and UO_263 (O_263,N_5215,N_6206);
nand UO_264 (O_264,N_8361,N_7960);
nand UO_265 (O_265,N_6556,N_7937);
and UO_266 (O_266,N_5341,N_8333);
xor UO_267 (O_267,N_9798,N_7470);
nand UO_268 (O_268,N_6585,N_8539);
nand UO_269 (O_269,N_7128,N_9725);
and UO_270 (O_270,N_8490,N_6103);
and UO_271 (O_271,N_9244,N_9906);
nand UO_272 (O_272,N_5557,N_7941);
xnor UO_273 (O_273,N_9358,N_7642);
nand UO_274 (O_274,N_5529,N_9441);
or UO_275 (O_275,N_6518,N_9553);
and UO_276 (O_276,N_5567,N_5785);
nand UO_277 (O_277,N_5500,N_8841);
nand UO_278 (O_278,N_9745,N_9574);
or UO_279 (O_279,N_8848,N_8026);
nor UO_280 (O_280,N_5834,N_8173);
and UO_281 (O_281,N_8694,N_7913);
nor UO_282 (O_282,N_8485,N_8776);
nand UO_283 (O_283,N_6548,N_5041);
and UO_284 (O_284,N_5743,N_9638);
and UO_285 (O_285,N_8541,N_7473);
and UO_286 (O_286,N_5363,N_7528);
nor UO_287 (O_287,N_7265,N_8550);
nand UO_288 (O_288,N_5591,N_6296);
and UO_289 (O_289,N_8604,N_8767);
nand UO_290 (O_290,N_6189,N_9538);
nor UO_291 (O_291,N_7363,N_5720);
xnor UO_292 (O_292,N_6736,N_8742);
xnor UO_293 (O_293,N_9191,N_8151);
nor UO_294 (O_294,N_9256,N_7200);
or UO_295 (O_295,N_5326,N_7808);
or UO_296 (O_296,N_5206,N_9002);
and UO_297 (O_297,N_6209,N_5030);
and UO_298 (O_298,N_6657,N_7855);
xnor UO_299 (O_299,N_6340,N_8248);
nor UO_300 (O_300,N_6200,N_8505);
xnor UO_301 (O_301,N_9921,N_6373);
xnor UO_302 (O_302,N_5544,N_7489);
or UO_303 (O_303,N_7150,N_9998);
nor UO_304 (O_304,N_6750,N_8992);
and UO_305 (O_305,N_5710,N_5643);
xnor UO_306 (O_306,N_7814,N_5514);
or UO_307 (O_307,N_9445,N_7799);
and UO_308 (O_308,N_5993,N_6319);
nand UO_309 (O_309,N_6637,N_5649);
or UO_310 (O_310,N_6345,N_7314);
and UO_311 (O_311,N_7131,N_9307);
nor UO_312 (O_312,N_9004,N_9557);
or UO_313 (O_313,N_5787,N_9500);
or UO_314 (O_314,N_6979,N_8022);
or UO_315 (O_315,N_6194,N_5684);
nand UO_316 (O_316,N_8787,N_7903);
nor UO_317 (O_317,N_9241,N_6868);
nand UO_318 (O_318,N_7776,N_8068);
or UO_319 (O_319,N_9336,N_6520);
and UO_320 (O_320,N_5081,N_5612);
nand UO_321 (O_321,N_6041,N_9916);
and UO_322 (O_322,N_7984,N_7089);
nor UO_323 (O_323,N_5095,N_5489);
and UO_324 (O_324,N_8687,N_5069);
xor UO_325 (O_325,N_6465,N_6120);
xnor UO_326 (O_326,N_9430,N_8695);
nor UO_327 (O_327,N_6809,N_6576);
xnor UO_328 (O_328,N_5505,N_6824);
nand UO_329 (O_329,N_9413,N_7802);
or UO_330 (O_330,N_5844,N_9261);
nand UO_331 (O_331,N_9114,N_8701);
or UO_332 (O_332,N_8758,N_7655);
nand UO_333 (O_333,N_5247,N_8737);
and UO_334 (O_334,N_6022,N_6941);
nand UO_335 (O_335,N_6591,N_8518);
or UO_336 (O_336,N_9621,N_8217);
nor UO_337 (O_337,N_9527,N_9060);
nand UO_338 (O_338,N_5396,N_5655);
and UO_339 (O_339,N_5379,N_6949);
xor UO_340 (O_340,N_8087,N_6081);
nor UO_341 (O_341,N_8614,N_7784);
or UO_342 (O_342,N_6767,N_6590);
xnor UO_343 (O_343,N_8332,N_5023);
nor UO_344 (O_344,N_7804,N_7882);
xnor UO_345 (O_345,N_6303,N_6171);
or UO_346 (O_346,N_7261,N_5244);
nor UO_347 (O_347,N_9660,N_7121);
and UO_348 (O_348,N_6766,N_8162);
nand UO_349 (O_349,N_9344,N_8891);
nor UO_350 (O_350,N_9675,N_9878);
or UO_351 (O_351,N_6870,N_5527);
and UO_352 (O_352,N_7832,N_9223);
xor UO_353 (O_353,N_5158,N_6659);
nand UO_354 (O_354,N_5916,N_5685);
nand UO_355 (O_355,N_6444,N_9733);
xnor UO_356 (O_356,N_7086,N_6956);
xnor UO_357 (O_357,N_5725,N_6742);
xor UO_358 (O_358,N_9507,N_8426);
and UO_359 (O_359,N_9573,N_8202);
or UO_360 (O_360,N_8581,N_7969);
and UO_361 (O_361,N_8423,N_8394);
nor UO_362 (O_362,N_7627,N_8724);
or UO_363 (O_363,N_7174,N_5980);
or UO_364 (O_364,N_7390,N_7387);
nor UO_365 (O_365,N_7599,N_8281);
nand UO_366 (O_366,N_8250,N_7186);
and UO_367 (O_367,N_8368,N_7009);
nand UO_368 (O_368,N_9409,N_7073);
or UO_369 (O_369,N_8463,N_9535);
nand UO_370 (O_370,N_8639,N_9801);
nor UO_371 (O_371,N_7058,N_9836);
xor UO_372 (O_372,N_7835,N_5668);
nor UO_373 (O_373,N_6223,N_5046);
xnor UO_374 (O_374,N_5613,N_7439);
and UO_375 (O_375,N_7555,N_7212);
nand UO_376 (O_376,N_6952,N_5490);
nor UO_377 (O_377,N_5156,N_7717);
and UO_378 (O_378,N_5172,N_8868);
and UO_379 (O_379,N_9946,N_8819);
xor UO_380 (O_380,N_9092,N_8225);
xnor UO_381 (O_381,N_5589,N_6674);
xnor UO_382 (O_382,N_7571,N_8515);
and UO_383 (O_383,N_8823,N_5088);
or UO_384 (O_384,N_7967,N_5548);
nor UO_385 (O_385,N_6056,N_6843);
nor UO_386 (O_386,N_7025,N_7010);
or UO_387 (O_387,N_5359,N_7155);
xor UO_388 (O_388,N_5473,N_9377);
xor UO_389 (O_389,N_5276,N_5165);
xnor UO_390 (O_390,N_5303,N_6360);
or UO_391 (O_391,N_6446,N_5389);
xor UO_392 (O_392,N_5779,N_7144);
and UO_393 (O_393,N_8057,N_5332);
nor UO_394 (O_394,N_5735,N_7262);
or UO_395 (O_395,N_8488,N_7195);
xor UO_396 (O_396,N_6842,N_5707);
nor UO_397 (O_397,N_5530,N_5586);
and UO_398 (O_398,N_5058,N_7026);
nand UO_399 (O_399,N_5524,N_5123);
xor UO_400 (O_400,N_8793,N_8916);
nor UO_401 (O_401,N_6831,N_5703);
nor UO_402 (O_402,N_6921,N_9615);
and UO_403 (O_403,N_5828,N_5953);
nor UO_404 (O_404,N_7241,N_6307);
nor UO_405 (O_405,N_6292,N_6764);
or UO_406 (O_406,N_5181,N_5983);
xor UO_407 (O_407,N_9284,N_5061);
and UO_408 (O_408,N_5056,N_8081);
nor UO_409 (O_409,N_7997,N_9146);
nand UO_410 (O_410,N_6253,N_9486);
or UO_411 (O_411,N_6799,N_8006);
nor UO_412 (O_412,N_9147,N_9987);
nor UO_413 (O_413,N_9087,N_6934);
nand UO_414 (O_414,N_9922,N_6492);
xor UO_415 (O_415,N_7253,N_7598);
nor UO_416 (O_416,N_7971,N_7019);
nand UO_417 (O_417,N_9851,N_7461);
nand UO_418 (O_418,N_6916,N_5131);
xnor UO_419 (O_419,N_5770,N_7785);
nor UO_420 (O_420,N_6851,N_7403);
or UO_421 (O_421,N_7409,N_9140);
xor UO_422 (O_422,N_9547,N_7688);
and UO_423 (O_423,N_9629,N_9866);
and UO_424 (O_424,N_9246,N_9075);
nand UO_425 (O_425,N_8558,N_7410);
xnor UO_426 (O_426,N_6579,N_5831);
nand UO_427 (O_427,N_7157,N_6564);
nor UO_428 (O_428,N_7464,N_5578);
xnor UO_429 (O_429,N_7929,N_6463);
nor UO_430 (O_430,N_5907,N_6172);
or UO_431 (O_431,N_5339,N_7766);
and UO_432 (O_432,N_7302,N_9522);
nand UO_433 (O_433,N_9953,N_8591);
xnor UO_434 (O_434,N_8038,N_5029);
or UO_435 (O_435,N_5225,N_9294);
and UO_436 (O_436,N_6037,N_9064);
nor UO_437 (O_437,N_8888,N_6149);
nand UO_438 (O_438,N_9190,N_7819);
nand UO_439 (O_439,N_7391,N_7810);
and UO_440 (O_440,N_5328,N_9711);
and UO_441 (O_441,N_5357,N_5696);
nor UO_442 (O_442,N_9348,N_8839);
xnor UO_443 (O_443,N_8207,N_6400);
and UO_444 (O_444,N_5101,N_9540);
and UO_445 (O_445,N_9329,N_5176);
nand UO_446 (O_446,N_9584,N_5015);
nand UO_447 (O_447,N_8586,N_8497);
nand UO_448 (O_448,N_7234,N_7156);
and UO_449 (O_449,N_5425,N_9963);
nand UO_450 (O_450,N_5155,N_8195);
xor UO_451 (O_451,N_5409,N_6386);
and UO_452 (O_452,N_5219,N_9118);
nand UO_453 (O_453,N_6210,N_5767);
nor UO_454 (O_454,N_9872,N_5625);
and UO_455 (O_455,N_8399,N_5708);
and UO_456 (O_456,N_5967,N_6048);
nand UO_457 (O_457,N_9084,N_9917);
nor UO_458 (O_458,N_5118,N_9990);
nor UO_459 (O_459,N_8163,N_9059);
or UO_460 (O_460,N_7597,N_6036);
or UO_461 (O_461,N_6749,N_8242);
and UO_462 (O_462,N_9536,N_7656);
xnor UO_463 (O_463,N_8039,N_7952);
nand UO_464 (O_464,N_8348,N_6337);
nand UO_465 (O_465,N_5089,N_8609);
nand UO_466 (O_466,N_7643,N_8633);
nand UO_467 (O_467,N_5535,N_5074);
nand UO_468 (O_468,N_9628,N_8713);
nor UO_469 (O_469,N_5298,N_9510);
xor UO_470 (O_470,N_6794,N_8718);
and UO_471 (O_471,N_6028,N_6090);
or UO_472 (O_472,N_7242,N_9727);
nand UO_473 (O_473,N_7358,N_5540);
and UO_474 (O_474,N_6177,N_6554);
and UO_475 (O_475,N_6966,N_7504);
and UO_476 (O_476,N_5635,N_6814);
nor UO_477 (O_477,N_5521,N_9426);
and UO_478 (O_478,N_5929,N_6093);
xnor UO_479 (O_479,N_8752,N_5671);
nand UO_480 (O_480,N_9456,N_5952);
nand UO_481 (O_481,N_7361,N_6892);
xnor UO_482 (O_482,N_6746,N_9694);
xor UO_483 (O_483,N_5436,N_7211);
nand UO_484 (O_484,N_8141,N_6933);
or UO_485 (O_485,N_6633,N_5465);
nand UO_486 (O_486,N_5371,N_6597);
and UO_487 (O_487,N_6230,N_9717);
and UO_488 (O_488,N_6840,N_8053);
nand UO_489 (O_489,N_6791,N_8342);
or UO_490 (O_490,N_9279,N_5758);
or UO_491 (O_491,N_9052,N_7552);
and UO_492 (O_492,N_8354,N_9349);
and UO_493 (O_493,N_7068,N_9475);
nand UO_494 (O_494,N_6031,N_5988);
nor UO_495 (O_495,N_5414,N_8440);
xnor UO_496 (O_496,N_5756,N_8472);
xor UO_497 (O_497,N_9106,N_8865);
xor UO_498 (O_498,N_9549,N_9433);
xor UO_499 (O_499,N_8924,N_8199);
nor UO_500 (O_500,N_8389,N_7032);
and UO_501 (O_501,N_8034,N_9030);
and UO_502 (O_502,N_9412,N_5372);
nor UO_503 (O_503,N_5615,N_9995);
nand UO_504 (O_504,N_7985,N_7001);
xor UO_505 (O_505,N_6375,N_6486);
and UO_506 (O_506,N_9296,N_7807);
xor UO_507 (O_507,N_8449,N_7138);
nor UO_508 (O_508,N_7748,N_5981);
nor UO_509 (O_509,N_5390,N_7338);
nand UO_510 (O_510,N_5486,N_6552);
xnor UO_511 (O_511,N_9517,N_7389);
or UO_512 (O_512,N_8535,N_5746);
and UO_513 (O_513,N_6664,N_7549);
nand UO_514 (O_514,N_7475,N_8862);
xnor UO_515 (O_515,N_9085,N_6001);
and UO_516 (O_516,N_5000,N_5587);
nand UO_517 (O_517,N_5574,N_8257);
nor UO_518 (O_518,N_9245,N_8587);
nand UO_519 (O_519,N_8504,N_8772);
and UO_520 (O_520,N_8387,N_6798);
xnor UO_521 (O_521,N_6134,N_7083);
nor UO_522 (O_522,N_6060,N_8284);
and UO_523 (O_523,N_5510,N_6416);
nand UO_524 (O_524,N_5007,N_8165);
and UO_525 (O_525,N_8683,N_7989);
or UO_526 (O_526,N_9218,N_7311);
nor UO_527 (O_527,N_8741,N_9642);
nand UO_528 (O_528,N_6351,N_9369);
nand UO_529 (O_529,N_5609,N_8734);
nor UO_530 (O_530,N_8460,N_9652);
and UO_531 (O_531,N_9318,N_7654);
nand UO_532 (O_532,N_5960,N_6724);
nor UO_533 (O_533,N_6050,N_7568);
or UO_534 (O_534,N_6354,N_6068);
nand UO_535 (O_535,N_5542,N_6385);
nand UO_536 (O_536,N_8524,N_6411);
and UO_537 (O_537,N_8892,N_6040);
and UO_538 (O_538,N_6396,N_9446);
nand UO_539 (O_539,N_8089,N_7723);
nor UO_540 (O_540,N_9291,N_5078);
or UO_541 (O_541,N_8635,N_5545);
and UO_542 (O_542,N_5853,N_6648);
nor UO_543 (O_543,N_8178,N_8730);
or UO_544 (O_544,N_6574,N_6417);
xnor UO_545 (O_545,N_8690,N_8648);
and UO_546 (O_546,N_5060,N_5485);
nor UO_547 (O_547,N_6271,N_6784);
nand UO_548 (O_548,N_9011,N_8873);
nand UO_549 (O_549,N_5502,N_8598);
and UO_550 (O_550,N_8209,N_7313);
xnor UO_551 (O_551,N_5816,N_6312);
xor UO_552 (O_552,N_8866,N_7310);
and UO_553 (O_553,N_9634,N_7308);
xnor UO_554 (O_554,N_9089,N_8124);
nand UO_555 (O_555,N_5454,N_8551);
nor UO_556 (O_556,N_6490,N_8420);
or UO_557 (O_557,N_9217,N_5117);
nand UO_558 (O_558,N_7811,N_9699);
or UO_559 (O_559,N_6815,N_8343);
or UO_560 (O_560,N_9069,N_7282);
nor UO_561 (O_561,N_6509,N_9359);
xnor UO_562 (O_562,N_9765,N_5238);
nand UO_563 (O_563,N_6881,N_8744);
or UO_564 (O_564,N_9346,N_7909);
xor UO_565 (O_565,N_6521,N_6095);
nor UO_566 (O_566,N_6044,N_7696);
or UO_567 (O_567,N_6607,N_6109);
xor UO_568 (O_568,N_6852,N_8964);
nand UO_569 (O_569,N_9160,N_6690);
or UO_570 (O_570,N_8381,N_5552);
or UO_571 (O_571,N_5498,N_6977);
nand UO_572 (O_572,N_6694,N_8201);
xnor UO_573 (O_573,N_5879,N_6954);
or UO_574 (O_574,N_7382,N_5360);
nand UO_575 (O_575,N_7479,N_8806);
nor UO_576 (O_576,N_9149,N_5013);
or UO_577 (O_577,N_9898,N_5579);
nor UO_578 (O_578,N_8627,N_5291);
nand UO_579 (O_579,N_9313,N_6092);
nand UO_580 (O_580,N_9364,N_7983);
nand UO_581 (O_581,N_9602,N_9554);
nor UO_582 (O_582,N_6789,N_9193);
nor UO_583 (O_583,N_6361,N_9094);
or UO_584 (O_584,N_8042,N_6228);
nor UO_585 (O_585,N_8043,N_9463);
nor UO_586 (O_586,N_9119,N_6260);
or UO_587 (O_587,N_9504,N_5385);
or UO_588 (O_588,N_7897,N_9372);
or UO_589 (O_589,N_9178,N_9671);
nor UO_590 (O_590,N_8608,N_5382);
nand UO_591 (O_591,N_5576,N_9761);
xor UO_592 (O_592,N_7565,N_6115);
and UO_593 (O_593,N_6519,N_6827);
xor UO_594 (O_594,N_9180,N_7269);
or UO_595 (O_595,N_7143,N_9783);
or UO_596 (O_596,N_9376,N_7573);
and UO_597 (O_597,N_9128,N_7545);
nand UO_598 (O_598,N_6464,N_5808);
or UO_599 (O_599,N_8590,N_7072);
and UO_600 (O_600,N_7773,N_5909);
nand UO_601 (O_601,N_5772,N_6692);
nor UO_602 (O_602,N_7392,N_7675);
nand UO_603 (O_603,N_6392,N_5755);
xnor UO_604 (O_604,N_9210,N_7994);
and UO_605 (O_605,N_5979,N_6256);
nor UO_606 (O_606,N_8362,N_7965);
nor UO_607 (O_607,N_5588,N_7017);
xnor UO_608 (O_608,N_6467,N_6147);
and UO_609 (O_609,N_9186,N_7621);
or UO_610 (O_610,N_5151,N_5971);
or UO_611 (O_611,N_8929,N_8765);
nand UO_612 (O_612,N_9368,N_8377);
xor UO_613 (O_613,N_9854,N_9937);
xnor UO_614 (O_614,N_5105,N_8792);
xnor UO_615 (O_615,N_7531,N_6713);
and UO_616 (O_616,N_7541,N_5594);
and UO_617 (O_617,N_9235,N_5221);
and UO_618 (O_618,N_7695,N_6971);
or UO_619 (O_619,N_8364,N_5986);
nand UO_620 (O_620,N_7430,N_7672);
nand UO_621 (O_621,N_7051,N_7284);
nor UO_622 (O_622,N_8188,N_9646);
xnor UO_623 (O_623,N_7305,N_8047);
or UO_624 (O_624,N_9352,N_6672);
and UO_625 (O_625,N_6154,N_7986);
nor UO_626 (O_626,N_8932,N_5035);
and UO_627 (O_627,N_5934,N_9687);
nand UO_628 (O_628,N_9102,N_7517);
nor UO_629 (O_629,N_5120,N_6522);
or UO_630 (O_630,N_5241,N_6610);
xor UO_631 (O_631,N_9017,N_7147);
nor UO_632 (O_632,N_6981,N_9176);
xor UO_633 (O_633,N_9045,N_7917);
nand UO_634 (O_634,N_6453,N_6907);
or UO_635 (O_635,N_6408,N_8685);
xnor UO_636 (O_636,N_6141,N_5596);
xor UO_637 (O_637,N_9325,N_6170);
nor UO_638 (O_638,N_6891,N_6557);
nand UO_639 (O_639,N_8153,N_9027);
nand UO_640 (O_640,N_9918,N_6277);
xor UO_641 (O_641,N_7615,N_5330);
nor UO_642 (O_642,N_5287,N_5883);
and UO_643 (O_643,N_9467,N_7481);
nand UO_644 (O_644,N_6744,N_8527);
or UO_645 (O_645,N_7008,N_6410);
nor UO_646 (O_646,N_6096,N_5433);
or UO_647 (O_647,N_8191,N_7004);
or UO_648 (O_648,N_7312,N_9579);
xnor UO_649 (O_649,N_6098,N_7171);
xor UO_650 (O_650,N_7813,N_5153);
or UO_651 (O_651,N_7677,N_6059);
and UO_652 (O_652,N_5139,N_9490);
nor UO_653 (O_653,N_6409,N_9127);
nand UO_654 (O_654,N_7827,N_8684);
nor UO_655 (O_655,N_6653,N_9626);
and UO_656 (O_656,N_9099,N_6358);
or UO_657 (O_657,N_7786,N_9145);
nor UO_658 (O_658,N_8689,N_8126);
nand UO_659 (O_659,N_6732,N_7257);
nor UO_660 (O_660,N_8893,N_8142);
and UO_661 (O_661,N_8877,N_7523);
xor UO_662 (O_662,N_8442,N_5248);
nand UO_663 (O_663,N_7140,N_8098);
and UO_664 (O_664,N_5106,N_5189);
or UO_665 (O_665,N_5650,N_9183);
nand UO_666 (O_666,N_6926,N_6261);
and UO_667 (O_667,N_6451,N_7562);
or UO_668 (O_668,N_5269,N_8147);
nor UO_669 (O_669,N_7044,N_6602);
and UO_670 (O_670,N_9880,N_9198);
nor UO_671 (O_671,N_9752,N_9012);
and UO_672 (O_672,N_5482,N_8206);
or UO_673 (O_673,N_6466,N_7137);
nor UO_674 (O_674,N_6295,N_8761);
xor UO_675 (O_675,N_5600,N_5125);
nand UO_676 (O_676,N_7374,N_9105);
and UO_677 (O_677,N_5819,N_7664);
and UO_678 (O_678,N_5786,N_5661);
nand UO_679 (O_679,N_6017,N_7570);
and UO_680 (O_680,N_9627,N_8405);
nand UO_681 (O_681,N_9684,N_7154);
xor UO_682 (O_682,N_7830,N_9498);
xor UO_683 (O_683,N_9542,N_6404);
or UO_684 (O_684,N_6395,N_9046);
and UO_685 (O_685,N_7423,N_5146);
xor UO_686 (O_686,N_6174,N_8556);
or UO_687 (O_687,N_7898,N_5690);
and UO_688 (O_688,N_9205,N_9616);
nand UO_689 (O_689,N_9355,N_9954);
xor UO_690 (O_690,N_9534,N_9605);
and UO_691 (O_691,N_9237,N_5009);
nor UO_692 (O_692,N_8971,N_8371);
nand UO_693 (O_693,N_6300,N_9919);
nand UO_694 (O_694,N_9138,N_5025);
nor UO_695 (O_695,N_5395,N_9255);
nor UO_696 (O_696,N_8602,N_6299);
and UO_697 (O_697,N_8816,N_9158);
and UO_698 (O_698,N_7822,N_8216);
and UO_699 (O_699,N_5705,N_7637);
xnor UO_700 (O_700,N_6627,N_6769);
nor UO_701 (O_701,N_7759,N_9015);
xnor UO_702 (O_702,N_5272,N_5001);
nor UO_703 (O_703,N_6856,N_7649);
nor UO_704 (O_704,N_6058,N_6454);
nor UO_705 (O_705,N_8080,N_7975);
xnor UO_706 (O_706,N_8227,N_5142);
and UO_707 (O_707,N_8259,N_6432);
xnor UO_708 (O_708,N_6274,N_6267);
xor UO_709 (O_709,N_8018,N_7425);
and UO_710 (O_710,N_8224,N_8538);
nor UO_711 (O_711,N_5412,N_5744);
nor UO_712 (O_712,N_7330,N_5590);
nand UO_713 (O_713,N_5918,N_9940);
and UO_714 (O_714,N_6461,N_6878);
or UO_715 (O_715,N_8421,N_9668);
and UO_716 (O_716,N_7756,N_7355);
or UO_717 (O_717,N_7442,N_6297);
xor UO_718 (O_718,N_7458,N_8624);
nand UO_719 (O_719,N_8930,N_5229);
nand UO_720 (O_720,N_6362,N_9974);
nor UO_721 (O_721,N_6370,N_7400);
and UO_722 (O_722,N_6201,N_5391);
and UO_723 (O_723,N_6057,N_6357);
nand UO_724 (O_724,N_6083,N_5961);
nor UO_725 (O_725,N_8118,N_6217);
xnor UO_726 (O_726,N_8498,N_5312);
nor UO_727 (O_727,N_6775,N_7901);
nor UO_728 (O_728,N_5322,N_8247);
xnor UO_729 (O_729,N_7750,N_9014);
xor UO_730 (O_730,N_6899,N_7752);
or UO_731 (O_731,N_7315,N_9287);
and UO_732 (O_732,N_8400,N_7685);
or UO_733 (O_733,N_5718,N_9824);
nor UO_734 (O_734,N_9797,N_6214);
xnor UO_735 (O_735,N_9530,N_9406);
nor UO_736 (O_736,N_9113,N_8200);
nand UO_737 (O_737,N_5411,N_8386);
or UO_738 (O_738,N_7204,N_6401);
xnor UO_739 (O_739,N_5876,N_5410);
xnor UO_740 (O_740,N_6583,N_7593);
and UO_741 (O_741,N_9883,N_7868);
nor UO_742 (O_742,N_9257,N_5491);
and UO_743 (O_743,N_9174,N_9981);
and UO_744 (O_744,N_8130,N_9405);
xnor UO_745 (O_745,N_9748,N_5719);
and UO_746 (O_746,N_9403,N_6528);
nor UO_747 (O_747,N_9090,N_9964);
xor UO_748 (O_748,N_9659,N_5716);
and UO_749 (O_749,N_8218,N_8998);
nand UO_750 (O_750,N_5006,N_8445);
nor UO_751 (O_751,N_7040,N_8478);
nor UO_752 (O_752,N_7250,N_6777);
nand UO_753 (O_753,N_6006,N_5184);
or UO_754 (O_754,N_6866,N_7709);
xnor UO_755 (O_755,N_6960,N_9923);
and UO_756 (O_756,N_6850,N_5968);
nor UO_757 (O_757,N_7947,N_9086);
nor UO_758 (O_758,N_6169,N_5317);
nand UO_759 (O_759,N_9239,N_6712);
nand UO_760 (O_760,N_7659,N_7177);
or UO_761 (O_761,N_8621,N_6711);
nand UO_762 (O_762,N_8369,N_9499);
xnor UO_763 (O_763,N_9131,N_7506);
and UO_764 (O_764,N_6243,N_5783);
nor UO_765 (O_765,N_7018,N_5122);
and UO_766 (O_766,N_6857,N_9704);
nor UO_767 (O_767,N_8545,N_6810);
nand UO_768 (O_768,N_6460,N_6656);
nor UO_769 (O_769,N_8974,N_6051);
and UO_770 (O_770,N_7999,N_9632);
nor UO_771 (O_771,N_9673,N_6421);
xor UO_772 (O_772,N_9996,N_8337);
or UO_773 (O_773,N_5691,N_6684);
and UO_774 (O_774,N_8879,N_7500);
xor UO_775 (O_775,N_9357,N_8870);
and UO_776 (O_776,N_8290,N_9713);
nand UO_777 (O_777,N_9861,N_9926);
xor UO_778 (O_778,N_7539,N_6595);
nand UO_779 (O_779,N_6094,N_9674);
or UO_780 (O_780,N_9379,N_9513);
and UO_781 (O_781,N_6500,N_6195);
nor UO_782 (O_782,N_7203,N_7182);
nand UO_783 (O_783,N_9061,N_8644);
or UO_784 (O_784,N_7603,N_8074);
nand UO_785 (O_785,N_5043,N_5466);
xor UO_786 (O_786,N_6053,N_9818);
nor UO_787 (O_787,N_7959,N_9077);
nand UO_788 (O_788,N_7336,N_9019);
nand UO_789 (O_789,N_9164,N_5914);
nor UO_790 (O_790,N_5966,N_7701);
nand UO_791 (O_791,N_5068,N_7581);
xor UO_792 (O_792,N_7127,N_6516);
xor UO_793 (O_793,N_5799,N_7589);
nand UO_794 (O_794,N_8000,N_6776);
nor UO_795 (O_795,N_9594,N_9526);
xor UO_796 (O_796,N_5205,N_7891);
or UO_797 (O_797,N_5620,N_8232);
or UO_798 (O_798,N_8418,N_6127);
nor UO_799 (O_799,N_9480,N_5806);
or UO_800 (O_800,N_7244,N_9231);
nand UO_801 (O_801,N_9908,N_5399);
xor UO_802 (O_802,N_8969,N_9427);
nor UO_803 (O_803,N_5289,N_9250);
xor UO_804 (O_804,N_7857,N_8778);
nand UO_805 (O_805,N_8537,N_7438);
xor UO_806 (O_806,N_8064,N_7053);
nand UO_807 (O_807,N_6598,N_8301);
nand UO_808 (O_808,N_6043,N_9610);
nand UO_809 (O_809,N_5859,N_9775);
nand UO_810 (O_810,N_5936,N_9787);
nor UO_811 (O_811,N_8923,N_8519);
nand UO_812 (O_812,N_8770,N_6049);
xor UO_813 (O_813,N_5077,N_6687);
or UO_814 (O_814,N_6806,N_6306);
xor UO_815 (O_815,N_9947,N_8297);
nor UO_816 (O_816,N_7918,N_7402);
or UO_817 (O_817,N_6512,N_6790);
or UO_818 (O_818,N_5300,N_9265);
nor UO_819 (O_819,N_6608,N_8311);
xor UO_820 (O_820,N_5543,N_6754);
or UO_821 (O_821,N_7399,N_6144);
nor UO_822 (O_822,N_8536,N_5602);
or UO_823 (O_823,N_5972,N_7585);
or UO_824 (O_824,N_8810,N_9525);
nand UO_825 (O_825,N_6157,N_9010);
nor UO_826 (O_826,N_5086,N_5672);
or UO_827 (O_827,N_6222,N_7514);
or UO_828 (O_828,N_5314,N_9185);
nor UO_829 (O_829,N_7493,N_6291);
nor UO_830 (O_830,N_6118,N_9395);
nor UO_831 (O_831,N_7979,N_7303);
nand UO_832 (O_832,N_9508,N_8465);
xor UO_833 (O_833,N_7020,N_9227);
and UO_834 (O_834,N_7420,N_8205);
nand UO_835 (O_835,N_9472,N_5424);
xnor UO_836 (O_836,N_8376,N_8951);
nor UO_837 (O_837,N_8315,N_6524);
nand UO_838 (O_838,N_5619,N_6990);
xnor UO_839 (O_839,N_5935,N_8170);
nor UO_840 (O_840,N_7287,N_6367);
nor UO_841 (O_841,N_5878,N_6443);
nand UO_842 (O_842,N_9096,N_5995);
and UO_843 (O_843,N_7448,N_6859);
or UO_844 (O_844,N_5132,N_5053);
xor UO_845 (O_845,N_8180,N_9882);
and UO_846 (O_846,N_9865,N_8258);
nor UO_847 (O_847,N_7604,N_7741);
xnor UO_848 (O_848,N_9399,N_9273);
nand UO_849 (O_849,N_6785,N_7240);
or UO_850 (O_850,N_9672,N_8268);
nand UO_851 (O_851,N_7594,N_5065);
nand UO_852 (O_852,N_9976,N_8313);
nand UO_853 (O_853,N_6846,N_7839);
and UO_854 (O_854,N_7467,N_9766);
nor UO_855 (O_855,N_8031,N_7012);
xor UO_856 (O_856,N_8104,N_7721);
xor UO_857 (O_857,N_5519,N_7638);
xor UO_858 (O_858,N_8020,N_9840);
and UO_859 (O_859,N_6739,N_8009);
nand UO_860 (O_860,N_7116,N_5114);
nand UO_861 (O_861,N_7337,N_7818);
xnor UO_862 (O_862,N_8896,N_9654);
xor UO_863 (O_863,N_6202,N_5085);
nor UO_864 (O_864,N_6168,N_5261);
nand UO_865 (O_865,N_8464,N_5008);
nor UO_866 (O_866,N_8424,N_5222);
nand UO_867 (O_867,N_8030,N_9308);
and UO_868 (O_868,N_9853,N_8867);
nand UO_869 (O_869,N_7081,N_9655);
or UO_870 (O_870,N_8956,N_8190);
xnor UO_871 (O_871,N_5994,N_9018);
nand UO_872 (O_872,N_9502,N_9989);
or UO_873 (O_873,N_8011,N_5932);
xor UO_874 (O_874,N_7109,N_9614);
xnor UO_875 (O_875,N_6343,N_5833);
or UO_876 (O_876,N_5022,N_5904);
nand UO_877 (O_877,N_5848,N_6349);
xnor UO_878 (O_878,N_8573,N_8041);
nand UO_879 (O_879,N_5945,N_6717);
nand UO_880 (O_880,N_5860,N_6531);
nand UO_881 (O_881,N_8499,N_8357);
nand UO_882 (O_882,N_9962,N_6561);
nand UO_883 (O_883,N_8655,N_7762);
or UO_884 (O_884,N_6264,N_9000);
or UO_885 (O_885,N_9539,N_8899);
nor UO_886 (O_886,N_5641,N_5152);
nand UO_887 (O_887,N_8582,N_6864);
nand UO_888 (O_888,N_7437,N_6126);
xnor UO_889 (O_889,N_8857,N_9442);
and UO_890 (O_890,N_8999,N_5495);
nand UO_891 (O_891,N_5239,N_7779);
nand UO_892 (O_892,N_9590,N_5667);
or UO_893 (O_893,N_7746,N_8061);
xor UO_894 (O_894,N_6654,N_8557);
and UO_895 (O_895,N_8106,N_5183);
xor UO_896 (O_896,N_8063,N_8322);
nand UO_897 (O_897,N_9982,N_5275);
xor UO_898 (O_898,N_9519,N_5044);
and UO_899 (O_899,N_5422,N_6932);
or UO_900 (O_900,N_7449,N_7101);
and UO_901 (O_901,N_9263,N_5234);
and UO_902 (O_902,N_5062,N_9870);
or UO_903 (O_903,N_9449,N_7170);
or UO_904 (O_904,N_5871,N_9887);
or UO_905 (O_905,N_5599,N_8559);
xor UO_906 (O_906,N_9777,N_8336);
and UO_907 (O_907,N_6281,N_6231);
nand UO_908 (O_908,N_8078,N_5393);
nor UO_909 (O_909,N_5135,N_9471);
xnor UO_910 (O_910,N_5627,N_5572);
nand UO_911 (O_911,N_8670,N_9735);
nand UO_912 (O_912,N_7459,N_6248);
nor UO_913 (O_913,N_7322,N_9458);
xnor UO_914 (O_914,N_7052,N_8012);
xor UO_915 (O_915,N_6896,N_9473);
or UO_916 (O_916,N_8155,N_6704);
xnor UO_917 (O_917,N_6671,N_9664);
nand UO_918 (O_918,N_7030,N_5124);
or UO_919 (O_919,N_5614,N_6252);
xnor UO_920 (O_920,N_7133,N_5481);
and UO_921 (O_921,N_7877,N_8145);
or UO_922 (O_922,N_5811,N_7801);
xor UO_923 (O_923,N_6477,N_9267);
and UO_924 (O_924,N_7745,N_9088);
nand UO_925 (O_925,N_6020,N_9242);
xor UO_926 (O_926,N_6425,N_6763);
nor UO_927 (O_927,N_5948,N_7927);
xnor UO_928 (O_928,N_9562,N_6835);
or UO_929 (O_929,N_5835,N_8264);
or UO_930 (O_930,N_6729,N_7817);
nor UO_931 (O_931,N_8707,N_6313);
and UO_932 (O_932,N_7843,N_5143);
and UO_933 (O_933,N_9063,N_6805);
nor UO_934 (O_934,N_7694,N_6188);
or UO_935 (O_935,N_7998,N_9129);
xnor UO_936 (O_936,N_6871,N_5869);
or UO_937 (O_937,N_8976,N_7576);
nor UO_938 (O_938,N_6216,N_8763);
xor UO_939 (O_939,N_7455,N_9091);
and UO_940 (O_940,N_6922,N_9083);
nor UO_941 (O_941,N_5306,N_5888);
nor UO_942 (O_942,N_8585,N_8859);
and UO_943 (O_943,N_5191,N_6288);
or UO_944 (O_944,N_8853,N_9184);
xor UO_945 (O_945,N_6244,N_5180);
xnor UO_946 (O_946,N_8466,N_6000);
or UO_947 (O_947,N_5516,N_5235);
and UO_948 (O_948,N_8845,N_9842);
xnor UO_949 (O_949,N_6667,N_6844);
or UO_950 (O_950,N_9742,N_8220);
and UO_951 (O_951,N_8698,N_7457);
or UO_952 (O_952,N_5843,N_9815);
and UO_953 (O_953,N_5622,N_9657);
and UO_954 (O_954,N_8825,N_5024);
xnor UO_955 (O_955,N_9835,N_6976);
and UO_956 (O_956,N_8091,N_5361);
and UO_957 (O_957,N_8618,N_8595);
nor UO_958 (O_958,N_8046,N_8033);
and UO_959 (O_959,N_9862,N_9316);
nor UO_960 (O_960,N_7345,N_9807);
xor UO_961 (O_961,N_9792,N_6418);
or UO_962 (O_962,N_8221,N_8448);
or UO_963 (O_963,N_5683,N_8959);
and UO_964 (O_964,N_6029,N_5977);
nor UO_965 (O_965,N_6738,N_5435);
xor UO_966 (O_966,N_8795,N_5413);
and UO_967 (O_967,N_8628,N_9169);
and UO_968 (O_968,N_5729,N_6335);
and UO_969 (O_969,N_8937,N_9806);
nor UO_970 (O_970,N_9207,N_9588);
nor UO_971 (O_971,N_9689,N_9056);
or UO_972 (O_972,N_9805,N_6483);
and UO_973 (O_973,N_9641,N_8764);
nor UO_974 (O_974,N_6091,N_7348);
and UO_975 (O_975,N_8760,N_8302);
nor UO_976 (O_976,N_6472,N_7478);
and UO_977 (O_977,N_9774,N_5447);
or UO_978 (O_978,N_9493,N_5174);
nor UO_979 (O_979,N_7554,N_8025);
and UO_980 (O_980,N_6038,N_8659);
nor UO_981 (O_981,N_7692,N_6326);
nand UO_982 (O_982,N_7720,N_8642);
or UO_983 (O_983,N_8528,N_8745);
or UO_984 (O_984,N_5846,N_6991);
or UO_985 (O_985,N_6885,N_5714);
and UO_986 (O_986,N_8731,N_5216);
xor UO_987 (O_987,N_7375,N_5870);
nand UO_988 (O_988,N_9679,N_6423);
nor UO_989 (O_989,N_8107,N_8843);
or UO_990 (O_990,N_5984,N_7125);
or UO_991 (O_991,N_7064,N_9702);
nor UO_992 (O_992,N_7974,N_8972);
nand UO_993 (O_993,N_8875,N_9782);
xnor UO_994 (O_994,N_7906,N_5531);
nor UO_995 (O_995,N_6139,N_5604);
xnor UO_996 (O_996,N_8372,N_7873);
nor UO_997 (O_997,N_8349,N_5711);
xnor UO_998 (O_998,N_5329,N_9967);
and UO_999 (O_999,N_9763,N_7787);
and UO_1000 (O_1000,N_9956,N_8254);
nand UO_1001 (O_1001,N_9141,N_5751);
and UO_1002 (O_1002,N_5978,N_9452);
nor UO_1003 (O_1003,N_7487,N_5823);
or UO_1004 (O_1004,N_5263,N_6219);
xnor UO_1005 (O_1005,N_7039,N_7700);
nor UO_1006 (O_1006,N_8392,N_8913);
or UO_1007 (O_1007,N_7496,N_8780);
xor UO_1008 (O_1008,N_9435,N_9220);
and UO_1009 (O_1009,N_5533,N_7118);
xor UO_1010 (O_1010,N_8692,N_5780);
xor UO_1011 (O_1011,N_7092,N_5581);
nand UO_1012 (O_1012,N_7115,N_9813);
nor UO_1013 (O_1013,N_8229,N_9034);
nand UO_1014 (O_1014,N_8230,N_6701);
or UO_1015 (O_1015,N_6193,N_5992);
nand UO_1016 (O_1016,N_8260,N_7160);
nand UO_1017 (O_1017,N_7714,N_8066);
nand UO_1018 (O_1018,N_6459,N_6331);
or UO_1019 (O_1019,N_8316,N_8833);
xnor UO_1020 (O_1020,N_6533,N_7865);
nand UO_1021 (O_1021,N_8968,N_5201);
xnor UO_1022 (O_1022,N_5805,N_7728);
nor UO_1023 (O_1023,N_6128,N_9764);
xor UO_1024 (O_1024,N_9678,N_6689);
or UO_1025 (O_1025,N_6184,N_8599);
nand UO_1026 (O_1026,N_5274,N_9281);
or UO_1027 (O_1027,N_8314,N_7796);
and UO_1028 (O_1028,N_8097,N_6619);
nor UO_1029 (O_1029,N_8223,N_8511);
nand UO_1030 (O_1030,N_6993,N_6164);
nor UO_1031 (O_1031,N_9951,N_5384);
or UO_1032 (O_1032,N_9760,N_8164);
or UO_1033 (O_1033,N_9721,N_7201);
nand UO_1034 (O_1034,N_8820,N_8732);
nor UO_1035 (O_1035,N_9363,N_8775);
nor UO_1036 (O_1036,N_9960,N_6811);
nand UO_1037 (O_1037,N_7260,N_7669);
nand UO_1038 (O_1038,N_6247,N_7911);
xnor UO_1039 (O_1039,N_5923,N_5397);
nand UO_1040 (O_1040,N_5673,N_7290);
nand UO_1041 (O_1041,N_9986,N_9686);
xnor UO_1042 (O_1042,N_6974,N_7406);
nand UO_1043 (O_1043,N_5378,N_8495);
xnor UO_1044 (O_1044,N_8016,N_9367);
xnor UO_1045 (O_1045,N_9293,N_5097);
nand UO_1046 (O_1046,N_7703,N_8049);
nand UO_1047 (O_1047,N_7281,N_9819);
xor UO_1048 (O_1048,N_5374,N_9903);
nor UO_1049 (O_1049,N_7447,N_9886);
or UO_1050 (O_1050,N_5733,N_7760);
nand UO_1051 (O_1051,N_9708,N_9125);
nand UO_1052 (O_1052,N_9685,N_8710);
or UO_1053 (O_1053,N_9778,N_9020);
xnor UO_1054 (O_1054,N_7846,N_6584);
xnor UO_1055 (O_1055,N_6014,N_9751);
or UO_1056 (O_1056,N_8275,N_9572);
xnor UO_1057 (O_1057,N_8800,N_8887);
nand UO_1058 (O_1058,N_8514,N_8198);
or UO_1059 (O_1059,N_6975,N_8496);
nand UO_1060 (O_1060,N_7548,N_5036);
xnor UO_1061 (O_1061,N_5631,N_6573);
or UO_1062 (O_1062,N_9877,N_6086);
nand UO_1063 (O_1063,N_8804,N_8327);
or UO_1064 (O_1064,N_7702,N_7600);
xnor UO_1065 (O_1065,N_9859,N_7607);
nor UO_1066 (O_1066,N_8443,N_8263);
nor UO_1067 (O_1067,N_8037,N_6931);
nand UO_1068 (O_1068,N_6484,N_8244);
nor UO_1069 (O_1069,N_8756,N_9767);
and UO_1070 (O_1070,N_5829,N_5145);
and UO_1071 (O_1071,N_9326,N_7230);
or UO_1072 (O_1072,N_6208,N_7958);
and UO_1073 (O_1073,N_5866,N_7080);
nand UO_1074 (O_1074,N_8186,N_6983);
xnor UO_1075 (O_1075,N_6624,N_6726);
or UO_1076 (O_1076,N_9123,N_7161);
nor UO_1077 (O_1077,N_7309,N_6105);
nand UO_1078 (O_1078,N_8874,N_6015);
nand UO_1079 (O_1079,N_7853,N_7626);
or UO_1080 (O_1080,N_8856,N_8453);
and UO_1081 (O_1081,N_6125,N_9172);
xor UO_1082 (O_1082,N_8430,N_7172);
nor UO_1083 (O_1083,N_5741,N_8204);
nand UO_1084 (O_1084,N_7090,N_7384);
nor UO_1085 (O_1085,N_5373,N_6628);
and UO_1086 (O_1086,N_9863,N_6647);
or UO_1087 (O_1087,N_7914,N_8542);
and UO_1088 (O_1088,N_8852,N_8697);
nand UO_1089 (O_1089,N_5911,N_8459);
nand UO_1090 (O_1090,N_9639,N_8214);
xor UO_1091 (O_1091,N_8251,N_8751);
and UO_1092 (O_1092,N_9896,N_6570);
and UO_1093 (O_1093,N_9389,N_5905);
nor UO_1094 (O_1094,N_5054,N_7609);
and UO_1095 (O_1095,N_8876,N_5082);
or UO_1096 (O_1096,N_6630,N_7844);
nand UO_1097 (O_1097,N_8653,N_8993);
xnor UO_1098 (O_1098,N_5845,N_7821);
nand UO_1099 (O_1099,N_5908,N_8015);
xnor UO_1100 (O_1100,N_8991,N_6435);
and UO_1101 (O_1101,N_8138,N_5776);
nand UO_1102 (O_1102,N_9633,N_6786);
nand UO_1103 (O_1103,N_7772,N_9879);
or UO_1104 (O_1104,N_7091,N_5944);
nor UO_1105 (O_1105,N_6911,N_5223);
and UO_1106 (O_1106,N_7869,N_6502);
and UO_1107 (O_1107,N_7468,N_6221);
nor UO_1108 (O_1108,N_9600,N_6848);
and UO_1109 (O_1109,N_9617,N_9768);
and UO_1110 (O_1110,N_6770,N_9249);
or UO_1111 (O_1111,N_6783,N_6237);
xor UO_1112 (O_1112,N_5618,N_5406);
nand UO_1113 (O_1113,N_8253,N_5638);
nor UO_1114 (O_1114,N_9757,N_6529);
nand UO_1115 (O_1115,N_6820,N_8934);
xor UO_1116 (O_1116,N_8375,N_7751);
nor UO_1117 (O_1117,N_9827,N_5940);
and UO_1118 (O_1118,N_5679,N_9800);
or UO_1119 (O_1119,N_7108,N_5258);
nand UO_1120 (O_1120,N_6612,N_5458);
xnor UO_1121 (O_1121,N_7737,N_7219);
nor UO_1122 (O_1122,N_8910,N_7508);
and UO_1123 (O_1123,N_9154,N_7483);
and UO_1124 (O_1124,N_9491,N_5997);
nand UO_1125 (O_1125,N_9469,N_6913);
nor UO_1126 (O_1126,N_6234,N_6587);
and UO_1127 (O_1127,N_5352,N_9997);
or UO_1128 (O_1128,N_7272,N_7255);
nand UO_1129 (O_1129,N_5345,N_9593);
or UO_1130 (O_1130,N_5562,N_8279);
nand UO_1131 (O_1131,N_7905,N_5640);
and UO_1132 (O_1132,N_8855,N_8660);
nor UO_1133 (O_1133,N_5532,N_8413);
and UO_1134 (O_1134,N_9970,N_7263);
nor UO_1135 (O_1135,N_8347,N_7353);
and UO_1136 (O_1136,N_6005,N_6969);
nand UO_1137 (O_1137,N_6918,N_8002);
nand UO_1138 (O_1138,N_9566,N_7953);
nand UO_1139 (O_1139,N_8678,N_8477);
and UO_1140 (O_1140,N_9163,N_7907);
nand UO_1141 (O_1141,N_5407,N_9984);
or UO_1142 (O_1142,N_7031,N_8437);
and UO_1143 (O_1143,N_6515,N_9816);
or UO_1144 (O_1144,N_5606,N_9843);
or UO_1145 (O_1145,N_5419,N_9795);
nand UO_1146 (O_1146,N_5686,N_6800);
or UO_1147 (O_1147,N_5577,N_6635);
nand UO_1148 (O_1148,N_5310,N_6886);
nand UO_1149 (O_1149,N_6663,N_6027);
or UO_1150 (O_1150,N_6829,N_7601);
xor UO_1151 (O_1151,N_9958,N_8076);
xnor UO_1152 (O_1152,N_9266,N_6116);
or UO_1153 (O_1153,N_6838,N_9669);
and UO_1154 (O_1154,N_5654,N_9315);
nand UO_1155 (O_1155,N_8788,N_6287);
or UO_1156 (O_1156,N_7574,N_6302);
nand UO_1157 (O_1157,N_8641,N_8391);
nand UO_1158 (O_1158,N_7826,N_7884);
nor UO_1159 (O_1159,N_8955,N_8093);
nor UO_1160 (O_1160,N_8849,N_5777);
nand UO_1161 (O_1161,N_9607,N_5838);
nand UO_1162 (O_1162,N_7507,N_8168);
nand UO_1163 (O_1163,N_7164,N_5592);
nand UO_1164 (O_1164,N_5877,N_9939);
nand UO_1165 (O_1165,N_5955,N_7484);
or UO_1166 (O_1166,N_7715,N_7828);
nor UO_1167 (O_1167,N_5136,N_5949);
xnor UO_1168 (O_1168,N_7043,N_8243);
or UO_1169 (O_1169,N_6158,N_8189);
xnor UO_1170 (O_1170,N_9565,N_7613);
nand UO_1171 (O_1171,N_7644,N_7299);
nand UO_1172 (O_1172,N_6320,N_8977);
and UO_1173 (O_1173,N_8851,N_9860);
xnor UO_1174 (O_1174,N_6316,N_8779);
nor UO_1175 (O_1175,N_8578,N_8620);
nand UO_1176 (O_1176,N_7511,N_9881);
nand UO_1177 (O_1177,N_5217,N_5566);
or UO_1178 (O_1178,N_6371,N_5040);
and UO_1179 (O_1179,N_7727,N_8663);
nor UO_1180 (O_1180,N_6441,N_5639);
nand UO_1181 (O_1181,N_6390,N_7676);
and UO_1182 (O_1182,N_8786,N_5209);
xor UO_1183 (O_1183,N_9959,N_6009);
and UO_1184 (O_1184,N_6821,N_9341);
and UO_1185 (O_1185,N_7747,N_7572);
or UO_1186 (O_1186,N_8565,N_5658);
or UO_1187 (O_1187,N_6626,N_7226);
or UO_1188 (O_1188,N_8940,N_7946);
and UO_1189 (O_1189,N_9428,N_7793);
nand UO_1190 (O_1190,N_6161,N_8654);
xnor UO_1191 (O_1191,N_7078,N_5154);
nand UO_1192 (O_1192,N_7167,N_5555);
and UO_1193 (O_1193,N_9108,N_7771);
and UO_1194 (O_1194,N_5110,N_8291);
and UO_1195 (O_1195,N_7838,N_8324);
nand UO_1196 (O_1196,N_7792,N_8917);
or UO_1197 (O_1197,N_8351,N_5355);
or UO_1198 (O_1198,N_5347,N_7707);
and UO_1199 (O_1199,N_9321,N_9338);
xnor UO_1200 (O_1200,N_7189,N_7660);
nor UO_1201 (O_1201,N_6731,N_8231);
and UO_1202 (O_1202,N_6699,N_6265);
xnor UO_1203 (O_1203,N_7237,N_6804);
xnor UO_1204 (O_1204,N_8987,N_5771);
or UO_1205 (O_1205,N_6963,N_5366);
and UO_1206 (O_1206,N_6951,N_9107);
or UO_1207 (O_1207,N_6982,N_8723);
xnor UO_1208 (O_1208,N_6493,N_5647);
nand UO_1209 (O_1209,N_8323,N_5109);
nor UO_1210 (O_1210,N_5441,N_7434);
xor UO_1211 (O_1211,N_9116,N_5063);
and UO_1212 (O_1212,N_5796,N_9366);
xnor UO_1213 (O_1213,N_7398,N_7158);
or UO_1214 (O_1214,N_8181,N_8261);
nor UO_1215 (O_1215,N_9758,N_7097);
xnor UO_1216 (O_1216,N_9224,N_7791);
nor UO_1217 (O_1217,N_5825,N_8809);
nor UO_1218 (O_1218,N_8664,N_6251);
xnor UO_1219 (O_1219,N_7534,N_6315);
xor UO_1220 (O_1220,N_6393,N_5957);
and UO_1221 (O_1221,N_6269,N_8794);
xnor UO_1222 (O_1222,N_8240,N_6412);
nand UO_1223 (O_1223,N_8900,N_7795);
nor UO_1224 (O_1224,N_7421,N_7770);
nor UO_1225 (O_1225,N_7289,N_6571);
xnor UO_1226 (O_1226,N_6153,N_9631);
nand UO_1227 (O_1227,N_7013,N_9691);
or UO_1228 (O_1228,N_9832,N_6761);
and UO_1229 (O_1229,N_5864,N_5768);
and UO_1230 (O_1230,N_5724,N_6002);
xnor UO_1231 (O_1231,N_8838,N_8815);
nand UO_1232 (O_1232,N_9779,N_8319);
or UO_1233 (O_1233,N_8306,N_5827);
or UO_1234 (O_1234,N_8150,N_6119);
xnor UO_1235 (O_1235,N_6327,N_6479);
nand UO_1236 (O_1236,N_8520,N_9936);
nand UO_1237 (O_1237,N_8722,N_6629);
or UO_1238 (O_1238,N_9032,N_6839);
and UO_1239 (O_1239,N_8566,N_9211);
xor UO_1240 (O_1240,N_9852,N_5951);
or UO_1241 (O_1241,N_9643,N_8543);
xor UO_1242 (O_1242,N_5450,N_5309);
and UO_1243 (O_1243,N_9236,N_7093);
nand UO_1244 (O_1244,N_9794,N_5930);
and UO_1245 (O_1245,N_8182,N_5503);
xnor UO_1246 (O_1246,N_8280,N_8433);
and UO_1247 (O_1247,N_6150,N_5461);
xnor UO_1248 (O_1248,N_5973,N_5499);
xnor UO_1249 (O_1249,N_9829,N_8045);
nor UO_1250 (O_1250,N_5731,N_6700);
xnor UO_1251 (O_1251,N_7887,N_5049);
nor UO_1252 (O_1252,N_6547,N_7317);
or UO_1253 (O_1253,N_9202,N_9247);
nor UO_1254 (O_1254,N_6272,N_8277);
xor UO_1255 (O_1255,N_9929,N_8222);
or UO_1256 (O_1256,N_6526,N_5912);
nor UO_1257 (O_1257,N_9994,N_5534);
xnor UO_1258 (O_1258,N_6324,N_9168);
nor UO_1259 (O_1259,N_7370,N_7509);
xor UO_1260 (O_1260,N_7112,N_8890);
nor UO_1261 (O_1261,N_6197,N_8881);
and UO_1262 (O_1262,N_6780,N_6447);
or UO_1263 (O_1263,N_9968,N_7662);
nand UO_1264 (O_1264,N_7103,N_8864);
xor UO_1265 (O_1265,N_8335,N_8826);
and UO_1266 (O_1266,N_8419,N_8167);
and UO_1267 (O_1267,N_7681,N_5296);
nand UO_1268 (O_1268,N_6973,N_5840);
nand UO_1269 (O_1269,N_8650,N_6879);
and UO_1270 (O_1270,N_6082,N_9892);
or UO_1271 (O_1271,N_9724,N_5874);
nand UO_1272 (O_1272,N_9812,N_5598);
nand UO_1273 (O_1273,N_9979,N_6873);
nand UO_1274 (O_1274,N_6910,N_9057);
or UO_1275 (O_1275,N_6218,N_5872);
nor UO_1276 (O_1276,N_7169,N_6278);
xnor UO_1277 (O_1277,N_8884,N_7592);
nor UO_1278 (O_1278,N_9450,N_9924);
nand UO_1279 (O_1279,N_8549,N_9143);
nand UO_1280 (O_1280,N_7647,N_8032);
and UO_1281 (O_1281,N_8305,N_5715);
nand UO_1282 (O_1282,N_6498,N_7217);
and UO_1283 (O_1283,N_7047,N_7663);
xnor UO_1284 (O_1284,N_9196,N_7774);
or UO_1285 (O_1285,N_7324,N_9142);
or UO_1286 (O_1286,N_5387,N_9544);
or UO_1287 (O_1287,N_5965,N_6560);
nor UO_1288 (O_1288,N_7622,N_7297);
nor UO_1289 (O_1289,N_5926,N_9311);
nand UO_1290 (O_1290,N_7129,N_7278);
or UO_1291 (O_1291,N_9104,N_8122);
or UO_1292 (O_1292,N_9564,N_7735);
nor UO_1293 (O_1293,N_6482,N_5826);
or UO_1294 (O_1294,N_8561,N_6262);
or UO_1295 (O_1295,N_5996,N_7896);
and UO_1296 (O_1296,N_6807,N_7102);
or UO_1297 (O_1297,N_9201,N_5802);
nand UO_1298 (O_1298,N_5583,N_7650);
or UO_1299 (O_1299,N_9076,N_9740);
and UO_1300 (O_1300,N_7347,N_6391);
or UO_1301 (O_1301,N_9869,N_5233);
and UO_1302 (O_1302,N_6117,N_8136);
and UO_1303 (O_1303,N_6753,N_6097);
xnor UO_1304 (O_1304,N_9891,N_9457);
nand UO_1305 (O_1305,N_7397,N_5457);
nor UO_1306 (O_1306,N_7344,N_7215);
nor UO_1307 (O_1307,N_5325,N_9398);
xnor UO_1308 (O_1308,N_5467,N_5438);
or UO_1309 (O_1309,N_9277,N_5119);
nand UO_1310 (O_1310,N_6996,N_6032);
or UO_1311 (O_1311,N_7286,N_8446);
nand UO_1312 (O_1312,N_9408,N_6836);
and UO_1313 (O_1313,N_9382,N_5652);
xor UO_1314 (O_1314,N_8798,N_9120);
nand UO_1315 (O_1315,N_5501,N_9411);
nand UO_1316 (O_1316,N_6199,N_8219);
nand UO_1317 (O_1317,N_7577,N_7666);
or UO_1318 (O_1318,N_8128,N_6436);
or UO_1319 (O_1319,N_6350,N_6972);
nand UO_1320 (O_1320,N_8861,N_5416);
nor UO_1321 (O_1321,N_7412,N_5236);
nand UO_1322 (O_1322,N_7059,N_5260);
nand UO_1323 (O_1323,N_9952,N_9276);
xnor UO_1324 (O_1324,N_5472,N_9285);
nor UO_1325 (O_1325,N_5898,N_6757);
xor UO_1326 (O_1326,N_5653,N_6948);
or UO_1327 (O_1327,N_6752,N_5693);
xnor UO_1328 (O_1328,N_6114,N_7699);
nor UO_1329 (O_1329,N_8077,N_8802);
nand UO_1330 (O_1330,N_6901,N_9581);
nor UO_1331 (O_1331,N_9942,N_8630);
and UO_1332 (O_1332,N_9596,N_9656);
nand UO_1333 (O_1333,N_8579,N_5913);
nor UO_1334 (O_1334,N_8293,N_9546);
xor UO_1335 (O_1335,N_8233,N_7122);
nand UO_1336 (O_1336,N_9601,N_7132);
nand UO_1337 (O_1337,N_7492,N_7407);
nand UO_1338 (O_1338,N_8355,N_5559);
or UO_1339 (O_1339,N_5839,N_5569);
nand UO_1340 (O_1340,N_8799,N_6758);
nor UO_1341 (O_1341,N_9410,N_6322);
or UO_1342 (O_1342,N_6087,N_6180);
or UO_1343 (O_1343,N_7307,N_5368);
nor UO_1344 (O_1344,N_9381,N_8102);
or UO_1345 (O_1345,N_5349,N_6818);
nand UO_1346 (O_1346,N_9440,N_6955);
and UO_1347 (O_1347,N_9303,N_6787);
xnor UO_1348 (O_1348,N_5231,N_5894);
nor UO_1349 (O_1349,N_7199,N_9005);
nor UO_1350 (O_1350,N_5307,N_7046);
or UO_1351 (O_1351,N_7049,N_8784);
nand UO_1352 (O_1352,N_5891,N_8938);
xor UO_1353 (O_1353,N_6077,N_5931);
nand UO_1354 (O_1354,N_8317,N_6212);
xor UO_1355 (O_1355,N_7364,N_5694);
and UO_1356 (O_1356,N_9676,N_8949);
nand UO_1357 (O_1357,N_5739,N_5546);
xor UO_1358 (O_1358,N_8014,N_6293);
or UO_1359 (O_1359,N_6532,N_9252);
nor UO_1360 (O_1360,N_9461,N_6033);
and UO_1361 (O_1361,N_5295,N_9153);
nand UO_1362 (O_1362,N_9384,N_5753);
nand UO_1363 (O_1363,N_5885,N_6010);
or UO_1364 (O_1364,N_8738,N_7815);
xnor UO_1365 (O_1365,N_8646,N_9556);
and UO_1366 (O_1366,N_7452,N_9033);
and UO_1367 (O_1367,N_9156,N_9230);
and UO_1368 (O_1368,N_5942,N_7945);
and UO_1369 (O_1369,N_6998,N_5726);
nor UO_1370 (O_1370,N_9744,N_5515);
and UO_1371 (O_1371,N_9492,N_9081);
xnor UO_1372 (O_1372,N_5875,N_5016);
and UO_1373 (O_1373,N_7726,N_5517);
or UO_1374 (O_1374,N_6342,N_7529);
nand UO_1375 (O_1375,N_7879,N_5224);
nand UO_1376 (O_1376,N_9187,N_8050);
nor UO_1377 (O_1377,N_5273,N_9194);
xnor UO_1378 (O_1378,N_8235,N_7367);
nand UO_1379 (O_1379,N_9680,N_8169);
and UO_1380 (O_1380,N_6917,N_5747);
nor UO_1381 (O_1381,N_6693,N_5187);
nand UO_1382 (O_1382,N_5327,N_7851);
nand UO_1383 (O_1383,N_5220,N_9054);
nor UO_1384 (O_1384,N_6514,N_5230);
xor UO_1385 (O_1385,N_8408,N_7028);
or UO_1386 (O_1386,N_5832,N_8404);
and UO_1387 (O_1387,N_5199,N_7288);
nand UO_1388 (O_1388,N_5417,N_6406);
or UO_1389 (O_1389,N_5915,N_7954);
and UO_1390 (O_1390,N_7943,N_5442);
and UO_1391 (O_1391,N_5426,N_8902);
nor UO_1392 (O_1392,N_9322,N_5865);
or UO_1393 (O_1393,N_6182,N_9009);
or UO_1394 (O_1394,N_7413,N_7862);
and UO_1395 (O_1395,N_7185,N_6298);
or UO_1396 (O_1396,N_6965,N_8728);
xnor UO_1397 (O_1397,N_7542,N_9286);
or UO_1398 (O_1398,N_8552,N_8402);
and UO_1399 (O_1399,N_8474,N_9503);
or UO_1400 (O_1400,N_9791,N_6867);
or UO_1401 (O_1401,N_8975,N_5293);
or UO_1402 (O_1402,N_9620,N_9066);
nand UO_1403 (O_1403,N_8226,N_9319);
nor UO_1404 (O_1404,N_8978,N_6642);
nand UO_1405 (O_1405,N_7494,N_6145);
and UO_1406 (O_1406,N_8177,N_9608);
nand UO_1407 (O_1407,N_9375,N_6347);
nand UO_1408 (O_1408,N_6468,N_6167);
xnor UO_1409 (O_1409,N_8990,N_8457);
and UO_1410 (O_1410,N_9552,N_9931);
or UO_1411 (O_1411,N_8640,N_6507);
and UO_1412 (O_1412,N_6388,N_7346);
xnor UO_1413 (O_1413,N_6906,N_6136);
or UO_1414 (O_1414,N_5161,N_9649);
nand UO_1415 (O_1415,N_9324,N_5429);
and UO_1416 (O_1416,N_8546,N_6751);
nor UO_1417 (O_1417,N_9705,N_8278);
and UO_1418 (O_1418,N_7561,N_7820);
nand UO_1419 (O_1419,N_7266,N_6304);
nor UO_1420 (O_1420,N_9333,N_5282);
nand UO_1421 (O_1421,N_9973,N_8652);
or UO_1422 (O_1422,N_6121,N_6394);
or UO_1423 (O_1423,N_8662,N_9888);
nor UO_1424 (O_1424,N_9762,N_7567);
nor UO_1425 (O_1425,N_5943,N_9712);
xnor UO_1426 (O_1426,N_8526,N_8393);
and UO_1427 (O_1427,N_8338,N_9932);
and UO_1428 (O_1428,N_5670,N_7380);
nor UO_1429 (O_1429,N_8797,N_5492);
or UO_1430 (O_1430,N_7148,N_7641);
xnor UO_1431 (O_1431,N_9203,N_7184);
and UO_1432 (O_1432,N_6355,N_8572);
nand UO_1433 (O_1433,N_6737,N_6430);
or UO_1434 (O_1434,N_9569,N_5551);
nand UO_1435 (O_1435,N_7719,N_7408);
and UO_1436 (O_1436,N_5769,N_9347);
or UO_1437 (O_1437,N_5821,N_8282);
nand UO_1438 (O_1438,N_6414,N_9934);
xor UO_1439 (O_1439,N_9589,N_9373);
xor UO_1440 (O_1440,N_9305,N_8193);
nor UO_1441 (O_1441,N_8237,N_7119);
or UO_1442 (O_1442,N_6328,N_8651);
or UO_1443 (O_1443,N_8740,N_9139);
nand UO_1444 (O_1444,N_6112,N_7841);
nand UO_1445 (O_1445,N_6356,N_8367);
nand UO_1446 (O_1446,N_9814,N_6861);
xor UO_1447 (O_1447,N_9563,N_8783);
nor UO_1448 (O_1448,N_9938,N_5164);
xor UO_1449 (O_1449,N_6229,N_8241);
or UO_1450 (O_1450,N_9876,N_8939);
nand UO_1451 (O_1451,N_9234,N_5810);
nand UO_1452 (O_1452,N_6792,N_9548);
xnor UO_1453 (O_1453,N_5757,N_8699);
nand UO_1454 (O_1454,N_6448,N_5676);
nor UO_1455 (O_1455,N_6165,N_7065);
and UO_1456 (O_1456,N_9845,N_6543);
nor UO_1457 (O_1457,N_7993,N_6148);
or UO_1458 (O_1458,N_7029,N_7803);
and UO_1459 (O_1459,N_5401,N_9999);
and UO_1460 (O_1460,N_5790,N_8560);
and UO_1461 (O_1461,N_5440,N_7733);
and UO_1462 (O_1462,N_8441,N_7267);
and UO_1463 (O_1463,N_5842,N_8796);
xor UO_1464 (O_1464,N_5836,N_7360);
nand UO_1465 (O_1465,N_6677,N_6883);
nand UO_1466 (O_1466,N_7094,N_8894);
nand UO_1467 (O_1467,N_5203,N_8246);
xor UO_1468 (O_1468,N_6823,N_8885);
xor UO_1469 (O_1469,N_8157,N_9512);
nor UO_1470 (O_1470,N_5112,N_6816);
nand UO_1471 (O_1471,N_6474,N_7925);
nor UO_1472 (O_1472,N_5459,N_9109);
nor UO_1473 (O_1473,N_6723,N_7225);
nor UO_1474 (O_1474,N_9541,N_7332);
nor UO_1475 (O_1475,N_9356,N_8435);
and UO_1476 (O_1476,N_9501,N_9514);
nor UO_1477 (O_1477,N_6334,N_6549);
xor UO_1478 (O_1478,N_5283,N_5506);
nand UO_1479 (O_1479,N_8606,N_9342);
or UO_1480 (O_1480,N_6173,N_6707);
nor UO_1481 (O_1481,N_7340,N_8208);
nand UO_1482 (O_1482,N_6681,N_5884);
and UO_1483 (O_1483,N_6936,N_6487);
nor UO_1484 (O_1484,N_9635,N_8149);
xnor UO_1485 (O_1485,N_5381,N_8774);
nand UO_1486 (O_1486,N_7145,N_8084);
nand UO_1487 (O_1487,N_8749,N_9524);
nand UO_1488 (O_1488,N_7863,N_5987);
xnor UO_1489 (O_1489,N_9478,N_6506);
or UO_1490 (O_1490,N_5646,N_6898);
nor UO_1491 (O_1491,N_9698,N_5752);
or UO_1492 (O_1492,N_9810,N_7369);
or UO_1493 (O_1493,N_5255,N_7236);
nand UO_1494 (O_1494,N_8516,N_8048);
and UO_1495 (O_1495,N_5079,N_6476);
nand UO_1496 (O_1496,N_8135,N_9173);
and UO_1497 (O_1497,N_5798,N_8397);
or UO_1498 (O_1498,N_5193,N_8941);
nor UO_1499 (O_1499,N_7636,N_6497);
endmodule