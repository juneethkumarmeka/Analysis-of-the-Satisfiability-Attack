module basic_1500_15000_2000_10_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_34,In_1381);
nand U1 (N_1,In_1322,In_1435);
and U2 (N_2,In_242,In_713);
nor U3 (N_3,In_1144,In_93);
nor U4 (N_4,In_871,In_380);
nand U5 (N_5,In_237,In_284);
nor U6 (N_6,In_903,In_1237);
xor U7 (N_7,In_644,In_383);
nand U8 (N_8,In_712,In_689);
or U9 (N_9,In_862,In_577);
nand U10 (N_10,In_549,In_57);
nor U11 (N_11,In_1443,In_1226);
and U12 (N_12,In_97,In_290);
nand U13 (N_13,In_1192,In_39);
and U14 (N_14,In_904,In_304);
nand U15 (N_15,In_1429,In_357);
nor U16 (N_16,In_1148,In_1297);
and U17 (N_17,In_951,In_771);
or U18 (N_18,In_981,In_1196);
and U19 (N_19,In_857,In_556);
and U20 (N_20,In_341,In_1191);
nor U21 (N_21,In_1127,In_491);
nor U22 (N_22,In_465,In_757);
or U23 (N_23,In_338,In_752);
and U24 (N_24,In_10,In_1221);
nor U25 (N_25,In_589,In_1092);
and U26 (N_26,In_730,In_222);
and U27 (N_27,In_1211,In_1366);
and U28 (N_28,In_68,In_675);
nand U29 (N_29,In_1491,In_1270);
nor U30 (N_30,In_459,In_762);
nand U31 (N_31,In_368,In_160);
or U32 (N_32,In_1496,In_287);
nand U33 (N_33,In_444,In_88);
nand U34 (N_34,In_568,In_1255);
xor U35 (N_35,In_1202,In_821);
nor U36 (N_36,In_317,In_1485);
or U37 (N_37,In_79,In_761);
nand U38 (N_38,In_480,In_831);
nor U39 (N_39,In_662,In_633);
nand U40 (N_40,In_63,In_519);
and U41 (N_41,In_132,In_126);
and U42 (N_42,In_728,In_807);
or U43 (N_43,In_106,In_103);
nand U44 (N_44,In_345,In_1220);
nand U45 (N_45,In_766,In_472);
and U46 (N_46,In_427,In_1200);
nor U47 (N_47,In_471,In_81);
nor U48 (N_48,In_939,In_1389);
nand U49 (N_49,In_1415,In_926);
nor U50 (N_50,In_124,In_748);
or U51 (N_51,In_369,In_227);
nand U52 (N_52,In_782,In_925);
or U53 (N_53,In_1019,In_1261);
nand U54 (N_54,In_300,In_1124);
nor U55 (N_55,In_964,In_1121);
nand U56 (N_56,In_869,In_687);
or U57 (N_57,In_94,In_113);
or U58 (N_58,In_1136,In_592);
nand U59 (N_59,In_924,In_350);
nand U60 (N_60,In_143,In_492);
and U61 (N_61,In_1084,In_234);
nor U62 (N_62,In_250,In_572);
and U63 (N_63,In_282,In_681);
or U64 (N_64,In_815,In_880);
nor U65 (N_65,In_796,In_1336);
nor U66 (N_66,In_54,In_179);
and U67 (N_67,In_1348,In_1341);
nand U68 (N_68,In_1360,In_927);
nor U69 (N_69,In_99,In_198);
or U70 (N_70,In_355,In_733);
nand U71 (N_71,In_354,In_1331);
or U72 (N_72,In_166,In_396);
nand U73 (N_73,In_1292,In_630);
or U74 (N_74,In_732,In_117);
and U75 (N_75,In_1117,In_348);
or U76 (N_76,In_213,In_1024);
nor U77 (N_77,In_1342,In_1377);
nor U78 (N_78,In_1390,In_588);
nor U79 (N_79,In_1154,In_1449);
and U80 (N_80,In_886,In_1495);
or U81 (N_81,In_878,In_703);
or U82 (N_82,In_605,In_1394);
nor U83 (N_83,In_55,In_858);
nor U84 (N_84,In_1278,In_1434);
and U85 (N_85,In_935,In_1268);
nor U86 (N_86,In_1418,In_521);
or U87 (N_87,In_1284,In_1146);
or U88 (N_88,In_940,In_1368);
nor U89 (N_89,In_1420,In_210);
nand U90 (N_90,In_990,In_1151);
or U91 (N_91,In_1033,In_629);
nand U92 (N_92,In_1138,In_1424);
nand U93 (N_93,In_252,In_42);
or U94 (N_94,In_911,In_421);
or U95 (N_95,In_1344,In_1359);
or U96 (N_96,In_508,In_150);
or U97 (N_97,In_646,In_1437);
nor U98 (N_98,In_810,In_848);
or U99 (N_99,In_1119,In_86);
nor U100 (N_100,In_76,In_1286);
and U101 (N_101,In_1419,In_929);
and U102 (N_102,In_1379,In_1014);
nor U103 (N_103,In_373,In_907);
and U104 (N_104,In_297,In_961);
and U105 (N_105,In_534,In_984);
nor U106 (N_106,In_1209,In_817);
or U107 (N_107,In_11,In_1294);
nand U108 (N_108,In_835,In_1256);
and U109 (N_109,In_1214,In_726);
nand U110 (N_110,In_777,In_1216);
or U111 (N_111,In_1006,In_507);
and U112 (N_112,In_46,In_310);
nor U113 (N_113,In_454,In_923);
nor U114 (N_114,In_545,In_1452);
or U115 (N_115,In_799,In_1269);
or U116 (N_116,In_488,In_1493);
or U117 (N_117,In_944,In_696);
nand U118 (N_118,In_468,In_403);
nor U119 (N_119,In_1364,In_275);
nand U120 (N_120,In_331,In_95);
and U121 (N_121,In_1012,In_1349);
xnor U122 (N_122,In_1258,In_288);
or U123 (N_123,In_390,In_426);
nand U124 (N_124,In_420,In_978);
nor U125 (N_125,In_82,In_147);
nand U126 (N_126,In_1334,In_970);
and U127 (N_127,In_746,In_567);
and U128 (N_128,In_755,In_191);
and U129 (N_129,In_187,In_538);
or U130 (N_130,In_1126,In_385);
nand U131 (N_131,In_679,In_1345);
nor U132 (N_132,In_1451,In_793);
or U133 (N_133,In_725,In_361);
nor U134 (N_134,In_1131,In_729);
nand U135 (N_135,In_1271,In_1038);
and U136 (N_136,In_772,In_405);
or U137 (N_137,In_685,In_74);
nand U138 (N_138,In_1018,In_408);
and U139 (N_139,In_335,In_6);
or U140 (N_140,In_44,In_531);
nand U141 (N_141,In_1480,In_631);
and U142 (N_142,In_812,In_255);
and U143 (N_143,In_1458,In_1078);
or U144 (N_144,In_975,In_1099);
nor U145 (N_145,In_25,In_482);
nor U146 (N_146,In_319,In_21);
or U147 (N_147,In_122,In_425);
nor U148 (N_148,In_316,In_625);
nand U149 (N_149,In_1369,In_749);
or U150 (N_150,In_3,In_906);
or U151 (N_151,In_1115,In_1179);
nand U152 (N_152,In_291,In_1027);
nor U153 (N_153,In_214,In_352);
nor U154 (N_154,In_220,In_334);
nand U155 (N_155,In_9,In_804);
nor U156 (N_156,In_389,In_1158);
or U157 (N_157,In_968,In_497);
and U158 (N_158,In_314,In_1464);
nand U159 (N_159,In_879,In_516);
or U160 (N_160,In_1071,In_228);
nor U161 (N_161,In_722,In_1408);
nor U162 (N_162,In_1484,In_170);
or U163 (N_163,In_461,In_194);
or U164 (N_164,In_1110,In_905);
or U165 (N_165,In_1152,In_1048);
or U166 (N_166,In_1059,In_641);
or U167 (N_167,In_834,In_30);
or U168 (N_168,In_1143,In_1350);
or U169 (N_169,In_1276,In_1194);
nand U170 (N_170,In_829,In_1353);
or U171 (N_171,In_18,In_43);
nand U172 (N_172,In_1260,In_5);
nand U173 (N_173,In_229,In_131);
and U174 (N_174,In_1135,In_359);
nand U175 (N_175,In_945,In_820);
or U176 (N_176,In_253,In_700);
nor U177 (N_177,In_1186,In_402);
or U178 (N_178,In_1188,In_384);
nor U179 (N_179,In_138,In_1282);
or U180 (N_180,In_684,In_230);
or U181 (N_181,In_649,In_261);
nor U182 (N_182,In_1210,In_1250);
and U183 (N_183,In_394,In_381);
nand U184 (N_184,In_558,In_1106);
nor U185 (N_185,In_1306,In_1430);
and U186 (N_186,In_717,In_1487);
or U187 (N_187,In_583,In_1241);
and U188 (N_188,In_702,In_153);
nor U189 (N_189,In_667,In_1102);
and U190 (N_190,In_109,In_443);
nor U191 (N_191,In_1346,In_1497);
and U192 (N_192,In_1343,In_524);
and U193 (N_193,In_526,In_315);
xnor U194 (N_194,In_1373,In_233);
nor U195 (N_195,In_745,In_1053);
nor U196 (N_196,In_349,In_24);
nand U197 (N_197,In_1446,In_175);
and U198 (N_198,In_606,In_1118);
or U199 (N_199,In_1242,In_72);
nor U200 (N_200,In_1448,In_655);
xor U201 (N_201,In_1397,In_1040);
nand U202 (N_202,In_870,In_636);
or U203 (N_203,In_1213,In_1317);
and U204 (N_204,In_794,In_654);
nand U205 (N_205,In_1468,In_1032);
nor U206 (N_206,In_1052,In_706);
or U207 (N_207,In_1382,In_1441);
nor U208 (N_208,In_37,In_1174);
xor U209 (N_209,In_270,In_1266);
or U210 (N_210,In_596,In_1312);
nor U211 (N_211,In_1181,In_223);
or U212 (N_212,In_118,In_785);
nand U213 (N_213,In_330,In_550);
and U214 (N_214,In_579,In_540);
and U215 (N_215,In_650,In_841);
or U216 (N_216,In_1080,In_578);
nand U217 (N_217,In_477,In_133);
nor U218 (N_218,In_1469,In_1083);
and U219 (N_219,In_140,In_98);
nand U220 (N_220,In_298,In_1045);
nor U221 (N_221,In_813,In_429);
nor U222 (N_222,In_165,In_487);
nor U223 (N_223,In_744,In_693);
and U224 (N_224,In_1228,In_895);
or U225 (N_225,In_274,In_1204);
nor U226 (N_226,In_888,In_863);
or U227 (N_227,In_678,In_1488);
nand U228 (N_228,In_983,In_914);
nor U229 (N_229,In_249,In_205);
and U230 (N_230,In_435,In_876);
nand U231 (N_231,In_245,In_321);
nor U232 (N_232,In_900,In_783);
and U233 (N_233,In_406,In_1470);
nor U234 (N_234,In_816,In_707);
nor U235 (N_235,In_1462,In_199);
and U236 (N_236,In_1310,In_466);
nor U237 (N_237,In_62,In_273);
and U238 (N_238,In_1130,In_172);
and U239 (N_239,In_1238,In_1016);
or U240 (N_240,In_1251,In_340);
and U241 (N_241,In_423,In_1476);
nand U242 (N_242,In_660,In_20);
nor U243 (N_243,In_1277,In_854);
nand U244 (N_244,In_741,In_195);
nand U245 (N_245,In_756,In_514);
and U246 (N_246,In_1316,In_1330);
nand U247 (N_247,In_149,In_963);
and U248 (N_248,In_1161,In_960);
nand U249 (N_249,In_1232,In_773);
nor U250 (N_250,In_343,In_1299);
and U251 (N_251,In_714,In_1421);
or U252 (N_252,In_1447,In_77);
nand U253 (N_253,In_720,In_825);
nor U254 (N_254,In_1372,In_1090);
nand U255 (N_255,In_544,In_155);
or U256 (N_256,In_1002,In_1122);
nor U257 (N_257,In_1004,In_1219);
or U258 (N_258,In_38,In_114);
or U259 (N_259,In_285,In_177);
nor U260 (N_260,In_1304,In_1086);
and U261 (N_261,In_1329,In_916);
nand U262 (N_262,In_872,In_1159);
and U263 (N_263,In_144,In_603);
or U264 (N_264,In_246,In_467);
nor U265 (N_265,In_202,In_1326);
and U266 (N_266,In_392,In_792);
xor U267 (N_267,In_683,In_27);
nor U268 (N_268,In_758,In_1378);
or U269 (N_269,In_1172,In_808);
or U270 (N_270,In_36,In_966);
and U271 (N_271,In_1054,In_1463);
nor U272 (N_272,In_1386,In_850);
nor U273 (N_273,In_174,In_329);
nand U274 (N_274,In_16,In_840);
and U275 (N_275,In_494,In_943);
nand U276 (N_276,In_613,In_1020);
nor U277 (N_277,In_499,In_948);
or U278 (N_278,In_1094,In_1363);
nor U279 (N_279,In_674,In_58);
nor U280 (N_280,In_176,In_1474);
or U281 (N_281,In_987,In_128);
and U282 (N_282,In_653,In_1058);
nand U283 (N_283,In_1478,In_374);
and U284 (N_284,In_115,In_1489);
nor U285 (N_285,In_740,In_784);
xor U286 (N_286,In_192,In_1340);
nor U287 (N_287,In_163,In_867);
and U288 (N_288,In_610,In_955);
nor U289 (N_289,In_826,In_1383);
or U290 (N_290,In_1233,In_565);
or U291 (N_291,In_1205,In_0);
nor U292 (N_292,In_1290,In_953);
and U293 (N_293,In_885,In_293);
nor U294 (N_294,In_372,In_1281);
nor U295 (N_295,In_1140,In_982);
nand U296 (N_296,In_600,In_735);
nand U297 (N_297,In_224,In_937);
or U298 (N_298,In_1400,In_1);
nand U299 (N_299,In_1347,In_1267);
and U300 (N_300,In_35,In_506);
nor U301 (N_301,In_621,In_204);
and U302 (N_302,In_1401,In_988);
xnor U303 (N_303,In_1178,In_690);
xor U304 (N_304,In_894,In_457);
or U305 (N_305,In_881,In_377);
and U306 (N_306,In_1450,In_364);
nand U307 (N_307,In_1185,In_1472);
and U308 (N_308,In_1007,In_186);
nand U309 (N_309,In_669,In_1407);
or U310 (N_310,In_611,In_809);
or U311 (N_311,In_645,In_1298);
or U312 (N_312,In_1236,In_292);
or U313 (N_313,In_1166,In_1065);
and U314 (N_314,In_1145,In_1153);
nor U315 (N_315,In_324,In_1272);
or U316 (N_316,In_1457,In_569);
nand U317 (N_317,In_837,In_1384);
nand U318 (N_318,In_325,In_620);
and U319 (N_319,In_573,In_1142);
nor U320 (N_320,In_861,In_1259);
and U321 (N_321,In_439,In_864);
nand U322 (N_322,In_1338,In_433);
and U323 (N_323,In_500,In_502);
or U324 (N_324,In_1376,In_1300);
nor U325 (N_325,In_989,In_560);
nand U326 (N_326,In_1055,In_1413);
nand U327 (N_327,In_995,In_263);
and U328 (N_328,In_597,In_1093);
nor U329 (N_329,In_278,In_56);
and U330 (N_330,In_208,In_201);
and U331 (N_331,In_416,In_281);
nor U332 (N_332,In_264,In_607);
or U333 (N_333,In_437,In_1223);
and U334 (N_334,In_962,In_440);
nand U335 (N_335,In_485,In_226);
or U336 (N_336,In_469,In_299);
or U337 (N_337,In_434,In_1165);
nand U338 (N_338,In_48,In_1050);
or U339 (N_339,In_604,In_686);
nand U340 (N_340,In_590,In_1182);
nand U341 (N_341,In_709,In_1440);
or U342 (N_342,In_901,In_1125);
and U343 (N_343,In_1461,In_279);
and U344 (N_344,In_193,In_481);
nand U345 (N_345,In_618,In_307);
nor U346 (N_346,In_1275,In_136);
nand U347 (N_347,In_798,In_1081);
nand U348 (N_348,In_883,In_407);
or U349 (N_349,In_814,In_1380);
nor U350 (N_350,In_770,In_1067);
and U351 (N_351,In_371,In_619);
nand U352 (N_352,In_1410,In_1147);
or U353 (N_353,In_543,In_1393);
or U354 (N_354,In_1392,In_708);
nand U355 (N_355,In_1481,In_146);
and U356 (N_356,In_120,In_346);
nand U357 (N_357,In_452,In_1456);
or U358 (N_358,In_1001,In_490);
and U359 (N_359,In_517,In_1077);
nand U360 (N_360,In_1325,In_1471);
nor U361 (N_361,In_173,In_13);
nand U362 (N_362,In_1168,In_1302);
nor U363 (N_363,In_1402,In_1351);
and U364 (N_364,In_890,In_1075);
nand U365 (N_365,In_609,In_1163);
nand U366 (N_366,In_1149,In_855);
nand U367 (N_367,In_1167,In_464);
nand U368 (N_368,In_476,In_387);
xnor U369 (N_369,In_1107,In_161);
xor U370 (N_370,In_542,In_1431);
nand U371 (N_371,In_313,In_1328);
nand U372 (N_372,In_723,In_1483);
nor U373 (N_373,In_1466,In_1439);
and U374 (N_374,In_257,In_156);
nor U375 (N_375,In_366,In_789);
nor U376 (N_376,In_1010,In_1318);
nor U377 (N_377,In_775,In_677);
nor U378 (N_378,In_1103,In_788);
and U379 (N_379,In_759,In_397);
nand U380 (N_380,In_1070,In_33);
or U381 (N_381,In_1460,In_1246);
nor U382 (N_382,In_1104,In_887);
nand U383 (N_383,In_130,In_638);
nand U384 (N_384,In_698,In_742);
nand U385 (N_385,In_1465,In_455);
or U386 (N_386,In_266,In_305);
nor U387 (N_387,In_811,In_721);
nand U388 (N_388,In_333,In_206);
and U389 (N_389,In_69,In_1253);
and U390 (N_390,In_1422,In_828);
and U391 (N_391,In_286,In_236);
nor U392 (N_392,In_1028,In_694);
and U393 (N_393,In_157,In_853);
and U394 (N_394,In_1433,In_1482);
nor U395 (N_395,In_1164,In_1370);
and U396 (N_396,In_376,In_110);
nor U397 (N_397,In_941,In_412);
and U398 (N_398,In_501,In_1137);
or U399 (N_399,In_134,In_167);
nor U400 (N_400,In_1051,In_436);
and U401 (N_401,In_111,In_294);
nor U402 (N_402,In_268,In_1222);
nand U403 (N_403,In_66,In_456);
nand U404 (N_404,In_142,In_493);
nand U405 (N_405,In_447,In_1239);
or U406 (N_406,In_453,In_1490);
and U407 (N_407,In_805,In_145);
nor U408 (N_408,In_216,In_979);
nor U409 (N_409,In_189,In_1287);
nor U410 (N_410,In_267,In_637);
or U411 (N_411,In_395,In_451);
nand U412 (N_412,In_1247,In_496);
nand U413 (N_413,In_965,In_976);
nand U414 (N_414,In_422,In_239);
and U415 (N_415,In_1293,In_84);
or U416 (N_416,In_673,In_1332);
and U417 (N_417,In_51,In_1034);
nand U418 (N_418,In_1438,In_530);
and U419 (N_419,In_415,In_428);
nor U420 (N_420,In_1358,In_116);
and U421 (N_421,In_779,In_78);
nand U422 (N_422,In_652,In_769);
nor U423 (N_423,In_936,In_541);
xnor U424 (N_424,In_238,In_28);
and U425 (N_425,In_1396,In_564);
or U426 (N_426,In_893,In_362);
nand U427 (N_427,In_67,In_1009);
nor U428 (N_428,In_289,In_1230);
or U429 (N_429,In_1475,In_363);
nor U430 (N_430,In_185,In_296);
or U431 (N_431,In_938,In_1013);
nor U432 (N_432,In_739,In_101);
nor U433 (N_433,In_1057,In_909);
nand U434 (N_434,In_998,In_986);
nand U435 (N_435,In_595,In_399);
and U436 (N_436,In_247,In_1215);
nand U437 (N_437,In_441,In_1008);
and U438 (N_438,In_29,In_1409);
nand U439 (N_439,In_866,In_581);
or U440 (N_440,In_884,In_1073);
nand U441 (N_441,In_1017,In_1187);
nor U442 (N_442,In_1025,In_1324);
or U443 (N_443,In_1229,In_642);
nand U444 (N_444,In_522,In_917);
and U445 (N_445,In_308,In_1085);
or U446 (N_446,In_235,In_119);
nor U447 (N_447,In_1217,In_505);
nor U448 (N_448,In_657,In_539);
nand U449 (N_449,In_999,In_715);
or U450 (N_450,In_697,In_1074);
or U451 (N_451,In_393,In_985);
nor U452 (N_452,In_462,In_932);
and U453 (N_453,In_1206,In_1335);
nand U454 (N_454,In_865,In_535);
and U455 (N_455,In_92,In_753);
nor U456 (N_456,In_2,In_1425);
nor U457 (N_457,In_1030,In_190);
nand U458 (N_458,In_328,In_580);
nor U459 (N_459,In_1207,In_896);
and U460 (N_460,In_692,In_1101);
nor U461 (N_461,In_949,In_875);
nand U462 (N_462,In_971,In_891);
nand U463 (N_463,In_908,In_1162);
nand U464 (N_464,In_410,In_431);
nand U465 (N_465,In_232,In_1072);
nand U466 (N_466,In_1399,In_1395);
and U467 (N_467,In_1371,In_1498);
or U468 (N_468,In_31,In_913);
nand U469 (N_469,In_337,In_209);
and U470 (N_470,In_358,In_1218);
nand U471 (N_471,In_1307,In_533);
nand U472 (N_472,In_910,In_921);
and U473 (N_473,In_557,In_1313);
and U474 (N_474,In_96,In_849);
nor U475 (N_475,In_1279,In_1288);
nand U476 (N_476,In_1337,In_1291);
nor U477 (N_477,In_169,In_575);
or U478 (N_478,In_659,In_561);
or U479 (N_479,In_776,In_152);
nand U480 (N_480,In_523,In_859);
or U481 (N_481,In_75,In_135);
and U482 (N_482,In_85,In_1355);
or U483 (N_483,In_323,In_1467);
nor U484 (N_484,In_892,In_15);
or U485 (N_485,In_1432,In_902);
and U486 (N_486,In_1046,In_790);
and U487 (N_487,In_129,In_634);
and U488 (N_488,In_52,In_486);
nor U489 (N_489,In_551,In_1169);
or U490 (N_490,In_845,In_718);
or U491 (N_491,In_53,In_622);
nor U492 (N_492,In_1225,In_993);
nor U493 (N_493,In_1327,In_400);
and U494 (N_494,In_1160,In_1303);
and U495 (N_495,In_515,In_882);
and U496 (N_496,In_992,In_1333);
or U497 (N_497,In_448,In_125);
and U498 (N_498,In_178,In_484);
nor U499 (N_499,In_599,In_764);
and U500 (N_500,In_168,In_382);
nand U501 (N_501,In_417,In_1082);
and U502 (N_502,In_158,In_419);
or U503 (N_503,In_1319,In_80);
nor U504 (N_504,In_1039,In_302);
nor U505 (N_505,In_474,In_1029);
nand U506 (N_506,In_360,In_272);
and U507 (N_507,In_1398,In_1494);
nor U508 (N_508,In_475,In_928);
nor U509 (N_509,In_1455,In_671);
nand U510 (N_510,In_1442,In_1454);
and U511 (N_511,In_1109,In_470);
nand U512 (N_512,In_954,In_1320);
nand U513 (N_513,In_1087,In_73);
nand U514 (N_514,In_873,In_391);
nand U515 (N_515,In_432,In_184);
nand U516 (N_516,In_1063,In_743);
and U517 (N_517,In_260,In_1044);
or U518 (N_518,In_547,In_1037);
or U519 (N_519,In_1245,In_154);
and U520 (N_520,In_1023,In_1295);
nand U521 (N_521,In_1375,In_503);
and U522 (N_522,In_219,In_1352);
or U523 (N_523,In_70,In_180);
or U524 (N_524,In_1416,In_483);
and U525 (N_525,In_727,In_1388);
or U526 (N_526,In_4,In_1309);
nand U527 (N_527,In_1096,In_1129);
and U528 (N_528,In_525,In_1305);
nor U529 (N_529,In_663,In_919);
nor U530 (N_530,In_958,In_563);
and U531 (N_531,In_1227,In_244);
or U532 (N_532,In_552,In_100);
nand U533 (N_533,In_912,In_1428);
nor U534 (N_534,In_258,In_585);
or U535 (N_535,In_90,In_701);
nor U536 (N_536,In_303,In_112);
nor U537 (N_537,In_856,In_370);
nand U538 (N_538,In_1041,In_1445);
nor U539 (N_539,In_635,In_868);
nand U540 (N_540,In_378,In_240);
nand U541 (N_541,In_554,In_123);
nand U542 (N_542,In_196,In_1254);
nand U543 (N_543,In_1022,In_22);
nor U544 (N_544,In_1095,In_1183);
nor U545 (N_545,In_774,In_778);
nor U546 (N_546,In_833,In_254);
nor U547 (N_547,In_584,In_1354);
nor U548 (N_548,In_915,In_1444);
xnor U549 (N_549,In_768,In_1120);
and U550 (N_550,In_137,In_277);
or U551 (N_551,In_724,In_780);
nor U552 (N_552,In_7,In_26);
and U553 (N_553,In_498,In_942);
and U554 (N_554,In_972,In_842);
nor U555 (N_555,In_736,In_947);
nand U556 (N_556,In_760,In_819);
or U557 (N_557,In_1231,In_1274);
nand U558 (N_558,In_711,In_1499);
nor U559 (N_559,In_218,In_473);
and U560 (N_560,In_791,In_509);
and U561 (N_561,In_61,In_19);
nor U562 (N_562,In_1426,In_665);
nand U563 (N_563,In_1177,In_401);
nand U564 (N_564,In_301,In_795);
nand U565 (N_565,In_1365,In_930);
or U566 (N_566,In_1189,In_1190);
nand U567 (N_567,In_716,In_1003);
nand U568 (N_568,In_1301,In_1112);
and U569 (N_569,In_40,In_217);
or U570 (N_570,In_594,In_1088);
nor U571 (N_571,In_151,In_1000);
nor U572 (N_572,In_632,In_832);
nand U573 (N_573,In_91,In_1035);
and U574 (N_574,In_64,In_747);
nor U575 (N_575,In_695,In_734);
and U576 (N_576,In_1098,In_351);
and U577 (N_577,In_513,In_1321);
nor U578 (N_578,In_553,In_957);
or U579 (N_579,In_676,In_87);
and U580 (N_580,In_148,In_1252);
nand U581 (N_581,In_946,In_386);
nand U582 (N_582,In_1141,In_801);
nand U583 (N_583,In_576,In_1404);
nor U584 (N_584,In_1011,In_1062);
and U585 (N_585,In_107,In_449);
or U586 (N_586,In_977,In_1170);
and U587 (N_587,In_311,In_1289);
xor U588 (N_588,In_105,In_510);
or U589 (N_589,In_1235,In_839);
or U590 (N_590,In_666,In_897);
nor U591 (N_591,In_787,In_108);
nor U592 (N_592,In_877,In_478);
or U593 (N_593,In_181,In_922);
or U594 (N_594,In_566,In_1243);
nand U595 (N_595,In_899,In_1273);
or U596 (N_596,In_1339,In_719);
and U597 (N_597,In_280,In_846);
nor U598 (N_598,In_1116,In_283);
or U599 (N_599,In_750,In_591);
or U600 (N_600,In_624,In_889);
nor U601 (N_601,In_537,In_860);
and U602 (N_602,In_1296,In_643);
nand U603 (N_603,In_200,In_991);
and U604 (N_604,In_822,In_45);
nand U605 (N_605,In_8,In_1234);
or U606 (N_606,In_626,In_570);
nand U607 (N_607,In_326,In_1385);
xor U608 (N_608,In_1417,In_1257);
and U609 (N_609,In_847,In_994);
and U610 (N_610,In_1105,In_183);
nor U611 (N_611,In_1201,In_32);
and U612 (N_612,In_141,In_738);
and U613 (N_613,In_339,In_1049);
nor U614 (N_614,In_710,In_571);
and U615 (N_615,In_1477,In_824);
or U616 (N_616,In_797,In_1031);
nor U617 (N_617,In_959,In_353);
nand U618 (N_618,In_1133,In_1405);
nand U619 (N_619,In_388,In_1056);
and U620 (N_620,In_670,In_1362);
or U621 (N_621,In_164,In_664);
and U622 (N_622,In_852,In_737);
nand U623 (N_623,In_559,In_1356);
nor U624 (N_624,In_1367,In_418);
or U625 (N_625,In_682,In_1026);
nand U626 (N_626,In_1157,In_705);
nand U627 (N_627,In_1411,In_271);
nand U628 (N_628,In_1180,In_104);
and U629 (N_629,In_511,In_956);
nand U630 (N_630,In_1021,In_1043);
and U631 (N_631,In_1171,In_159);
nor U632 (N_632,In_269,In_1114);
nand U633 (N_633,In_446,In_1212);
nor U634 (N_634,In_1280,In_512);
nor U635 (N_635,In_997,In_731);
and U636 (N_636,In_967,In_639);
or U637 (N_637,In_379,In_398);
nand U638 (N_638,In_139,In_479);
and U639 (N_639,In_404,In_898);
nor U640 (N_640,In_786,In_1374);
or U641 (N_641,In_680,In_127);
nor U642 (N_642,In_598,In_615);
and U643 (N_643,In_952,In_1492);
and U644 (N_644,In_950,In_1453);
nor U645 (N_645,In_691,In_640);
nand U646 (N_646,In_256,In_648);
or U647 (N_647,In_874,In_241);
or U648 (N_648,In_49,In_207);
and U649 (N_649,In_555,In_23);
nor U650 (N_650,In_309,In_1089);
nand U651 (N_651,In_215,In_934);
xnor U652 (N_652,In_844,In_1097);
nand U653 (N_653,In_1015,In_342);
nand U654 (N_654,In_1066,In_562);
nand U655 (N_655,In_375,In_413);
and U656 (N_656,In_1208,In_751);
nand U657 (N_657,In_212,In_1199);
nor U658 (N_658,In_50,In_688);
nor U659 (N_659,In_1262,In_102);
nor U660 (N_660,In_617,In_1091);
nor U661 (N_661,In_1047,In_781);
and U662 (N_662,In_409,In_532);
nand U663 (N_663,In_1387,In_243);
nor U664 (N_664,In_322,In_1005);
and U665 (N_665,In_647,In_356);
nor U666 (N_666,In_344,In_65);
nor U667 (N_667,In_1357,In_445);
and U668 (N_668,In_1197,In_1060);
nor U669 (N_669,In_614,In_836);
and U670 (N_670,In_489,In_248);
and U671 (N_671,In_1193,In_838);
or U672 (N_672,In_616,In_1132);
and U673 (N_673,In_587,In_1283);
nand U674 (N_674,In_231,In_1473);
nand U675 (N_675,In_1176,In_754);
nand U676 (N_676,In_320,In_528);
nand U677 (N_677,In_450,In_704);
nor U678 (N_678,In_1264,In_295);
or U679 (N_679,In_1113,In_536);
or U680 (N_680,In_593,In_851);
nand U681 (N_681,In_262,In_546);
and U682 (N_682,In_211,In_627);
and U683 (N_683,In_1108,In_1061);
nor U684 (N_684,In_1195,In_1079);
nand U685 (N_685,In_933,In_520);
nor U686 (N_686,In_203,In_1249);
and U687 (N_687,In_623,In_612);
nand U688 (N_688,In_527,In_162);
nor U689 (N_689,In_424,In_1184);
xor U690 (N_690,In_121,In_800);
and U691 (N_691,In_1175,In_306);
nor U692 (N_692,In_969,In_504);
or U693 (N_693,In_974,In_518);
nand U694 (N_694,In_438,In_365);
nand U695 (N_695,In_803,In_818);
and U696 (N_696,In_89,In_197);
and U697 (N_697,In_586,In_765);
nor U698 (N_698,In_1414,In_1459);
and U699 (N_699,In_318,In_602);
or U700 (N_700,In_1064,In_1224);
or U701 (N_701,In_495,In_1315);
or U702 (N_702,In_1412,In_656);
nand U703 (N_703,In_601,In_1263);
or U704 (N_704,In_574,In_83);
and U705 (N_705,In_14,In_1100);
or U706 (N_706,In_529,In_763);
and U707 (N_707,In_582,In_608);
nor U708 (N_708,In_996,In_668);
nor U709 (N_709,In_60,In_843);
nor U710 (N_710,In_1486,In_1198);
and U711 (N_711,In_463,In_1128);
and U712 (N_712,In_276,In_188);
nor U713 (N_713,In_336,In_12);
and U714 (N_714,In_1156,In_41);
nor U715 (N_715,In_259,In_347);
nor U716 (N_716,In_548,In_658);
nor U717 (N_717,In_628,In_1139);
nand U718 (N_718,In_171,In_931);
nor U719 (N_719,In_1323,In_327);
and U720 (N_720,In_1076,In_1036);
or U721 (N_721,In_920,In_332);
nand U722 (N_722,In_1134,In_47);
or U723 (N_723,In_460,In_1427);
nor U724 (N_724,In_1314,In_1406);
and U725 (N_725,In_823,In_71);
or U726 (N_726,In_1203,In_1308);
nand U727 (N_727,In_1042,In_802);
nand U728 (N_728,In_1155,In_367);
or U729 (N_729,In_827,In_1123);
nand U730 (N_730,In_830,In_1285);
and U731 (N_731,In_1479,In_1068);
or U732 (N_732,In_1391,In_1311);
and U733 (N_733,In_265,In_225);
and U734 (N_734,In_1248,In_1069);
nand U735 (N_735,In_1173,In_221);
nor U736 (N_736,In_806,In_699);
nand U737 (N_737,In_1244,In_251);
nor U738 (N_738,In_973,In_651);
nor U739 (N_739,In_17,In_59);
nor U740 (N_740,In_1403,In_1361);
and U741 (N_741,In_1111,In_414);
nand U742 (N_742,In_442,In_767);
nor U743 (N_743,In_1265,In_1150);
or U744 (N_744,In_312,In_182);
nand U745 (N_745,In_672,In_411);
nand U746 (N_746,In_980,In_430);
and U747 (N_747,In_661,In_1240);
or U748 (N_748,In_458,In_1436);
nand U749 (N_749,In_918,In_1423);
and U750 (N_750,In_1002,In_1092);
or U751 (N_751,In_1360,In_863);
nand U752 (N_752,In_307,In_1335);
and U753 (N_753,In_395,In_312);
nor U754 (N_754,In_838,In_656);
or U755 (N_755,In_1366,In_1068);
nor U756 (N_756,In_585,In_699);
nor U757 (N_757,In_1056,In_378);
and U758 (N_758,In_809,In_354);
or U759 (N_759,In_547,In_992);
nor U760 (N_760,In_1059,In_247);
nor U761 (N_761,In_270,In_122);
and U762 (N_762,In_1472,In_562);
nand U763 (N_763,In_574,In_563);
or U764 (N_764,In_991,In_1268);
nor U765 (N_765,In_232,In_22);
or U766 (N_766,In_263,In_740);
or U767 (N_767,In_1341,In_1157);
or U768 (N_768,In_1396,In_248);
nor U769 (N_769,In_985,In_627);
nor U770 (N_770,In_1446,In_491);
or U771 (N_771,In_609,In_1167);
nand U772 (N_772,In_258,In_1229);
nor U773 (N_773,In_1241,In_753);
nor U774 (N_774,In_394,In_626);
or U775 (N_775,In_744,In_728);
or U776 (N_776,In_819,In_622);
nor U777 (N_777,In_427,In_1416);
nor U778 (N_778,In_845,In_879);
nor U779 (N_779,In_446,In_288);
nand U780 (N_780,In_82,In_381);
or U781 (N_781,In_13,In_208);
nor U782 (N_782,In_631,In_506);
or U783 (N_783,In_567,In_1117);
and U784 (N_784,In_1110,In_101);
nor U785 (N_785,In_1232,In_1005);
nand U786 (N_786,In_170,In_59);
or U787 (N_787,In_302,In_484);
nand U788 (N_788,In_263,In_1387);
nand U789 (N_789,In_852,In_960);
nor U790 (N_790,In_1482,In_451);
and U791 (N_791,In_1211,In_608);
or U792 (N_792,In_641,In_931);
xnor U793 (N_793,In_174,In_1229);
nor U794 (N_794,In_1092,In_890);
and U795 (N_795,In_1494,In_93);
and U796 (N_796,In_1175,In_999);
or U797 (N_797,In_1133,In_170);
nor U798 (N_798,In_164,In_104);
nor U799 (N_799,In_421,In_1497);
xor U800 (N_800,In_356,In_86);
nor U801 (N_801,In_1114,In_378);
and U802 (N_802,In_359,In_1107);
nor U803 (N_803,In_322,In_1227);
nand U804 (N_804,In_715,In_730);
or U805 (N_805,In_303,In_239);
nand U806 (N_806,In_85,In_209);
nor U807 (N_807,In_305,In_1429);
or U808 (N_808,In_926,In_909);
nand U809 (N_809,In_481,In_765);
and U810 (N_810,In_382,In_1051);
nand U811 (N_811,In_822,In_292);
and U812 (N_812,In_826,In_387);
and U813 (N_813,In_243,In_229);
nor U814 (N_814,In_360,In_1280);
nor U815 (N_815,In_511,In_299);
and U816 (N_816,In_1430,In_551);
nor U817 (N_817,In_977,In_1039);
and U818 (N_818,In_718,In_294);
or U819 (N_819,In_179,In_542);
nand U820 (N_820,In_1353,In_812);
or U821 (N_821,In_1391,In_1150);
nor U822 (N_822,In_1422,In_160);
and U823 (N_823,In_667,In_139);
or U824 (N_824,In_782,In_1107);
nor U825 (N_825,In_982,In_1076);
nand U826 (N_826,In_260,In_801);
and U827 (N_827,In_546,In_1133);
and U828 (N_828,In_411,In_562);
nor U829 (N_829,In_1202,In_470);
and U830 (N_830,In_1039,In_140);
or U831 (N_831,In_287,In_1287);
nand U832 (N_832,In_715,In_713);
or U833 (N_833,In_455,In_410);
nand U834 (N_834,In_907,In_1058);
and U835 (N_835,In_837,In_678);
or U836 (N_836,In_886,In_642);
or U837 (N_837,In_1313,In_148);
or U838 (N_838,In_1301,In_205);
or U839 (N_839,In_1159,In_921);
and U840 (N_840,In_477,In_182);
and U841 (N_841,In_1337,In_533);
and U842 (N_842,In_1166,In_1089);
nor U843 (N_843,In_462,In_283);
nor U844 (N_844,In_337,In_324);
nor U845 (N_845,In_1140,In_1137);
and U846 (N_846,In_584,In_547);
nand U847 (N_847,In_1430,In_747);
nand U848 (N_848,In_188,In_893);
nor U849 (N_849,In_725,In_147);
or U850 (N_850,In_292,In_172);
and U851 (N_851,In_869,In_405);
or U852 (N_852,In_303,In_592);
and U853 (N_853,In_354,In_413);
nor U854 (N_854,In_713,In_1276);
nor U855 (N_855,In_208,In_657);
nand U856 (N_856,In_190,In_323);
nor U857 (N_857,In_472,In_823);
or U858 (N_858,In_191,In_809);
and U859 (N_859,In_1102,In_255);
and U860 (N_860,In_212,In_836);
and U861 (N_861,In_957,In_1084);
nor U862 (N_862,In_1372,In_1289);
and U863 (N_863,In_1285,In_1005);
and U864 (N_864,In_843,In_1022);
nor U865 (N_865,In_524,In_227);
and U866 (N_866,In_181,In_601);
nor U867 (N_867,In_955,In_17);
nand U868 (N_868,In_865,In_474);
or U869 (N_869,In_1425,In_820);
nor U870 (N_870,In_634,In_966);
nor U871 (N_871,In_522,In_1089);
and U872 (N_872,In_1486,In_72);
and U873 (N_873,In_369,In_360);
nor U874 (N_874,In_294,In_670);
and U875 (N_875,In_1024,In_902);
nor U876 (N_876,In_610,In_1394);
nand U877 (N_877,In_503,In_1352);
nand U878 (N_878,In_910,In_80);
or U879 (N_879,In_1220,In_276);
and U880 (N_880,In_570,In_256);
or U881 (N_881,In_1402,In_1154);
nand U882 (N_882,In_1495,In_819);
and U883 (N_883,In_940,In_1231);
and U884 (N_884,In_772,In_205);
nand U885 (N_885,In_1330,In_1190);
nor U886 (N_886,In_1022,In_981);
nand U887 (N_887,In_1088,In_40);
or U888 (N_888,In_1451,In_1249);
nand U889 (N_889,In_198,In_18);
and U890 (N_890,In_159,In_55);
or U891 (N_891,In_1232,In_641);
nand U892 (N_892,In_739,In_1048);
or U893 (N_893,In_803,In_977);
or U894 (N_894,In_893,In_903);
and U895 (N_895,In_735,In_896);
nor U896 (N_896,In_297,In_1310);
and U897 (N_897,In_469,In_722);
nor U898 (N_898,In_278,In_935);
nor U899 (N_899,In_934,In_578);
and U900 (N_900,In_619,In_361);
nor U901 (N_901,In_776,In_961);
and U902 (N_902,In_1433,In_1457);
and U903 (N_903,In_1019,In_484);
and U904 (N_904,In_976,In_1123);
or U905 (N_905,In_155,In_415);
nor U906 (N_906,In_975,In_360);
nand U907 (N_907,In_1071,In_674);
nor U908 (N_908,In_615,In_967);
nor U909 (N_909,In_424,In_1009);
or U910 (N_910,In_166,In_668);
or U911 (N_911,In_666,In_372);
nor U912 (N_912,In_1068,In_1416);
nand U913 (N_913,In_478,In_126);
and U914 (N_914,In_1289,In_805);
xnor U915 (N_915,In_491,In_484);
and U916 (N_916,In_432,In_1249);
nand U917 (N_917,In_204,In_6);
or U918 (N_918,In_861,In_185);
and U919 (N_919,In_368,In_1440);
or U920 (N_920,In_566,In_1007);
nor U921 (N_921,In_1340,In_435);
nor U922 (N_922,In_935,In_1441);
nand U923 (N_923,In_375,In_836);
xor U924 (N_924,In_443,In_124);
nand U925 (N_925,In_280,In_1318);
nand U926 (N_926,In_751,In_274);
or U927 (N_927,In_912,In_904);
nor U928 (N_928,In_433,In_629);
or U929 (N_929,In_890,In_1390);
nand U930 (N_930,In_1165,In_1252);
nor U931 (N_931,In_845,In_1392);
or U932 (N_932,In_438,In_828);
and U933 (N_933,In_1420,In_608);
and U934 (N_934,In_454,In_729);
and U935 (N_935,In_457,In_649);
nor U936 (N_936,In_929,In_1260);
nand U937 (N_937,In_776,In_1455);
or U938 (N_938,In_41,In_1236);
nor U939 (N_939,In_1034,In_1448);
nor U940 (N_940,In_1127,In_838);
or U941 (N_941,In_1271,In_1154);
nor U942 (N_942,In_359,In_484);
and U943 (N_943,In_124,In_921);
or U944 (N_944,In_133,In_1071);
and U945 (N_945,In_565,In_1399);
nor U946 (N_946,In_694,In_133);
nor U947 (N_947,In_1214,In_27);
nand U948 (N_948,In_1475,In_547);
or U949 (N_949,In_1324,In_428);
nand U950 (N_950,In_1359,In_844);
or U951 (N_951,In_514,In_1257);
or U952 (N_952,In_651,In_1027);
or U953 (N_953,In_329,In_387);
nand U954 (N_954,In_1071,In_961);
nand U955 (N_955,In_1301,In_1388);
and U956 (N_956,In_89,In_1448);
nand U957 (N_957,In_1385,In_522);
nor U958 (N_958,In_638,In_1124);
or U959 (N_959,In_989,In_109);
nand U960 (N_960,In_1266,In_1267);
nor U961 (N_961,In_1473,In_693);
nor U962 (N_962,In_1412,In_1426);
nand U963 (N_963,In_577,In_1223);
nand U964 (N_964,In_876,In_1061);
or U965 (N_965,In_1178,In_922);
xnor U966 (N_966,In_1169,In_1068);
nor U967 (N_967,In_480,In_1425);
nand U968 (N_968,In_1017,In_996);
or U969 (N_969,In_841,In_912);
or U970 (N_970,In_663,In_509);
or U971 (N_971,In_892,In_81);
and U972 (N_972,In_187,In_557);
nor U973 (N_973,In_889,In_1397);
and U974 (N_974,In_1099,In_1127);
or U975 (N_975,In_609,In_870);
nand U976 (N_976,In_260,In_526);
and U977 (N_977,In_618,In_1071);
and U978 (N_978,In_1470,In_1448);
and U979 (N_979,In_1424,In_909);
nand U980 (N_980,In_1324,In_681);
or U981 (N_981,In_131,In_684);
nor U982 (N_982,In_1440,In_473);
and U983 (N_983,In_190,In_1369);
or U984 (N_984,In_187,In_243);
nor U985 (N_985,In_793,In_1100);
nor U986 (N_986,In_1001,In_328);
nand U987 (N_987,In_540,In_1265);
nand U988 (N_988,In_419,In_710);
nor U989 (N_989,In_1202,In_760);
or U990 (N_990,In_24,In_1151);
nand U991 (N_991,In_1079,In_181);
nand U992 (N_992,In_1497,In_500);
or U993 (N_993,In_590,In_850);
nand U994 (N_994,In_641,In_106);
nand U995 (N_995,In_1245,In_884);
or U996 (N_996,In_524,In_951);
or U997 (N_997,In_1483,In_101);
nand U998 (N_998,In_1499,In_896);
and U999 (N_999,In_587,In_237);
and U1000 (N_1000,In_60,In_315);
or U1001 (N_1001,In_500,In_162);
or U1002 (N_1002,In_250,In_1409);
and U1003 (N_1003,In_497,In_635);
nand U1004 (N_1004,In_537,In_438);
or U1005 (N_1005,In_651,In_489);
nand U1006 (N_1006,In_1204,In_86);
or U1007 (N_1007,In_1449,In_281);
or U1008 (N_1008,In_557,In_730);
and U1009 (N_1009,In_1244,In_1146);
nand U1010 (N_1010,In_1028,In_1308);
and U1011 (N_1011,In_1058,In_844);
and U1012 (N_1012,In_936,In_62);
nand U1013 (N_1013,In_81,In_868);
nand U1014 (N_1014,In_658,In_1426);
nor U1015 (N_1015,In_468,In_425);
nand U1016 (N_1016,In_813,In_180);
nor U1017 (N_1017,In_1417,In_1125);
and U1018 (N_1018,In_812,In_734);
or U1019 (N_1019,In_461,In_959);
nand U1020 (N_1020,In_455,In_1109);
or U1021 (N_1021,In_62,In_1434);
and U1022 (N_1022,In_669,In_847);
or U1023 (N_1023,In_283,In_841);
nor U1024 (N_1024,In_1314,In_1014);
nand U1025 (N_1025,In_165,In_258);
nor U1026 (N_1026,In_1436,In_1292);
or U1027 (N_1027,In_1089,In_838);
nor U1028 (N_1028,In_381,In_319);
nand U1029 (N_1029,In_1242,In_1366);
or U1030 (N_1030,In_1460,In_989);
or U1031 (N_1031,In_60,In_214);
nand U1032 (N_1032,In_1047,In_1285);
or U1033 (N_1033,In_1477,In_352);
nand U1034 (N_1034,In_428,In_1303);
and U1035 (N_1035,In_1471,In_38);
nor U1036 (N_1036,In_171,In_307);
nand U1037 (N_1037,In_1313,In_337);
or U1038 (N_1038,In_1181,In_478);
nor U1039 (N_1039,In_1114,In_423);
nor U1040 (N_1040,In_1217,In_1167);
and U1041 (N_1041,In_418,In_1255);
or U1042 (N_1042,In_437,In_769);
and U1043 (N_1043,In_584,In_237);
nor U1044 (N_1044,In_1286,In_227);
nor U1045 (N_1045,In_49,In_744);
and U1046 (N_1046,In_907,In_1110);
or U1047 (N_1047,In_960,In_1083);
or U1048 (N_1048,In_314,In_631);
nor U1049 (N_1049,In_1415,In_384);
nand U1050 (N_1050,In_668,In_1106);
or U1051 (N_1051,In_10,In_1247);
nand U1052 (N_1052,In_677,In_801);
nand U1053 (N_1053,In_557,In_1494);
or U1054 (N_1054,In_338,In_148);
and U1055 (N_1055,In_251,In_1167);
and U1056 (N_1056,In_323,In_233);
and U1057 (N_1057,In_191,In_1338);
nor U1058 (N_1058,In_713,In_433);
nand U1059 (N_1059,In_270,In_1166);
or U1060 (N_1060,In_1291,In_285);
or U1061 (N_1061,In_102,In_1118);
and U1062 (N_1062,In_860,In_1409);
nand U1063 (N_1063,In_1373,In_1246);
nor U1064 (N_1064,In_866,In_1296);
nor U1065 (N_1065,In_839,In_1319);
or U1066 (N_1066,In_1113,In_330);
nand U1067 (N_1067,In_1041,In_228);
nor U1068 (N_1068,In_611,In_157);
or U1069 (N_1069,In_228,In_293);
nor U1070 (N_1070,In_115,In_756);
or U1071 (N_1071,In_863,In_964);
or U1072 (N_1072,In_1301,In_426);
and U1073 (N_1073,In_272,In_1280);
nand U1074 (N_1074,In_65,In_129);
nand U1075 (N_1075,In_298,In_652);
and U1076 (N_1076,In_1201,In_769);
or U1077 (N_1077,In_187,In_297);
and U1078 (N_1078,In_1272,In_25);
and U1079 (N_1079,In_1244,In_1079);
and U1080 (N_1080,In_1308,In_540);
nand U1081 (N_1081,In_1041,In_1025);
or U1082 (N_1082,In_444,In_1389);
nor U1083 (N_1083,In_1163,In_868);
or U1084 (N_1084,In_1390,In_651);
nor U1085 (N_1085,In_711,In_196);
nand U1086 (N_1086,In_968,In_589);
and U1087 (N_1087,In_626,In_251);
nor U1088 (N_1088,In_1017,In_387);
nor U1089 (N_1089,In_6,In_844);
nand U1090 (N_1090,In_887,In_531);
nor U1091 (N_1091,In_1210,In_323);
nand U1092 (N_1092,In_1021,In_273);
nor U1093 (N_1093,In_442,In_506);
nor U1094 (N_1094,In_802,In_690);
nand U1095 (N_1095,In_71,In_614);
or U1096 (N_1096,In_1298,In_821);
nand U1097 (N_1097,In_1316,In_195);
or U1098 (N_1098,In_393,In_684);
or U1099 (N_1099,In_1146,In_6);
nand U1100 (N_1100,In_26,In_932);
nor U1101 (N_1101,In_1216,In_759);
nand U1102 (N_1102,In_316,In_123);
nand U1103 (N_1103,In_914,In_958);
and U1104 (N_1104,In_599,In_1383);
nor U1105 (N_1105,In_498,In_51);
and U1106 (N_1106,In_1165,In_110);
nor U1107 (N_1107,In_812,In_162);
and U1108 (N_1108,In_14,In_1478);
nor U1109 (N_1109,In_253,In_1162);
and U1110 (N_1110,In_1378,In_925);
nand U1111 (N_1111,In_936,In_15);
nor U1112 (N_1112,In_816,In_1265);
and U1113 (N_1113,In_1290,In_955);
nor U1114 (N_1114,In_450,In_609);
and U1115 (N_1115,In_756,In_1043);
nand U1116 (N_1116,In_326,In_359);
and U1117 (N_1117,In_556,In_1066);
nor U1118 (N_1118,In_305,In_1312);
nor U1119 (N_1119,In_831,In_694);
and U1120 (N_1120,In_1238,In_1350);
nand U1121 (N_1121,In_605,In_1085);
nor U1122 (N_1122,In_1279,In_517);
nand U1123 (N_1123,In_895,In_585);
nor U1124 (N_1124,In_882,In_969);
nor U1125 (N_1125,In_70,In_1102);
and U1126 (N_1126,In_1049,In_810);
nor U1127 (N_1127,In_1357,In_297);
nand U1128 (N_1128,In_1304,In_936);
and U1129 (N_1129,In_569,In_787);
or U1130 (N_1130,In_20,In_577);
or U1131 (N_1131,In_101,In_573);
or U1132 (N_1132,In_376,In_240);
nor U1133 (N_1133,In_1202,In_466);
or U1134 (N_1134,In_1296,In_299);
or U1135 (N_1135,In_617,In_530);
nor U1136 (N_1136,In_446,In_799);
nor U1137 (N_1137,In_1333,In_1417);
nor U1138 (N_1138,In_60,In_1436);
nand U1139 (N_1139,In_659,In_819);
and U1140 (N_1140,In_772,In_1203);
and U1141 (N_1141,In_1356,In_1431);
nor U1142 (N_1142,In_1432,In_1433);
nor U1143 (N_1143,In_733,In_174);
and U1144 (N_1144,In_53,In_525);
or U1145 (N_1145,In_69,In_999);
nand U1146 (N_1146,In_772,In_951);
and U1147 (N_1147,In_1013,In_771);
and U1148 (N_1148,In_92,In_486);
nand U1149 (N_1149,In_676,In_321);
nor U1150 (N_1150,In_1246,In_1345);
nor U1151 (N_1151,In_869,In_520);
nand U1152 (N_1152,In_979,In_1412);
and U1153 (N_1153,In_1041,In_784);
or U1154 (N_1154,In_677,In_675);
nand U1155 (N_1155,In_1481,In_1240);
nor U1156 (N_1156,In_1425,In_585);
nor U1157 (N_1157,In_1378,In_1034);
nand U1158 (N_1158,In_1141,In_602);
or U1159 (N_1159,In_410,In_300);
nor U1160 (N_1160,In_1037,In_767);
or U1161 (N_1161,In_423,In_1105);
and U1162 (N_1162,In_1165,In_451);
or U1163 (N_1163,In_835,In_710);
or U1164 (N_1164,In_536,In_1272);
nand U1165 (N_1165,In_325,In_806);
or U1166 (N_1166,In_682,In_204);
and U1167 (N_1167,In_853,In_19);
or U1168 (N_1168,In_472,In_47);
nand U1169 (N_1169,In_1284,In_120);
or U1170 (N_1170,In_515,In_568);
and U1171 (N_1171,In_1114,In_247);
nand U1172 (N_1172,In_1371,In_700);
and U1173 (N_1173,In_906,In_410);
nand U1174 (N_1174,In_868,In_75);
nand U1175 (N_1175,In_1435,In_494);
or U1176 (N_1176,In_107,In_1242);
nand U1177 (N_1177,In_1435,In_1243);
or U1178 (N_1178,In_305,In_824);
and U1179 (N_1179,In_325,In_1472);
or U1180 (N_1180,In_691,In_243);
or U1181 (N_1181,In_1416,In_1324);
nor U1182 (N_1182,In_631,In_44);
or U1183 (N_1183,In_940,In_1393);
nand U1184 (N_1184,In_1497,In_1079);
nor U1185 (N_1185,In_223,In_481);
and U1186 (N_1186,In_255,In_1366);
nand U1187 (N_1187,In_569,In_262);
nand U1188 (N_1188,In_1294,In_666);
nand U1189 (N_1189,In_838,In_551);
or U1190 (N_1190,In_1087,In_229);
or U1191 (N_1191,In_1206,In_212);
nand U1192 (N_1192,In_264,In_33);
nand U1193 (N_1193,In_166,In_1433);
or U1194 (N_1194,In_959,In_76);
nor U1195 (N_1195,In_368,In_329);
nand U1196 (N_1196,In_1196,In_40);
and U1197 (N_1197,In_1175,In_360);
nand U1198 (N_1198,In_704,In_325);
nand U1199 (N_1199,In_99,In_203);
nand U1200 (N_1200,In_34,In_1240);
and U1201 (N_1201,In_558,In_341);
or U1202 (N_1202,In_422,In_398);
nand U1203 (N_1203,In_1041,In_1276);
nor U1204 (N_1204,In_95,In_701);
nand U1205 (N_1205,In_1299,In_1204);
nor U1206 (N_1206,In_555,In_790);
and U1207 (N_1207,In_140,In_533);
nand U1208 (N_1208,In_807,In_1332);
nand U1209 (N_1209,In_878,In_302);
nor U1210 (N_1210,In_414,In_517);
or U1211 (N_1211,In_774,In_243);
nand U1212 (N_1212,In_805,In_643);
or U1213 (N_1213,In_545,In_1291);
nor U1214 (N_1214,In_749,In_701);
or U1215 (N_1215,In_83,In_693);
or U1216 (N_1216,In_977,In_1116);
and U1217 (N_1217,In_883,In_1464);
and U1218 (N_1218,In_844,In_201);
nor U1219 (N_1219,In_334,In_1429);
nand U1220 (N_1220,In_988,In_526);
nand U1221 (N_1221,In_1290,In_1221);
and U1222 (N_1222,In_30,In_1486);
or U1223 (N_1223,In_753,In_5);
and U1224 (N_1224,In_1029,In_1024);
nand U1225 (N_1225,In_14,In_666);
nor U1226 (N_1226,In_1342,In_530);
nand U1227 (N_1227,In_922,In_943);
or U1228 (N_1228,In_3,In_1311);
and U1229 (N_1229,In_56,In_1006);
nand U1230 (N_1230,In_1013,In_342);
and U1231 (N_1231,In_1409,In_407);
or U1232 (N_1232,In_644,In_1241);
or U1233 (N_1233,In_1378,In_1202);
nand U1234 (N_1234,In_1097,In_364);
or U1235 (N_1235,In_718,In_758);
nor U1236 (N_1236,In_1229,In_979);
or U1237 (N_1237,In_1336,In_638);
or U1238 (N_1238,In_691,In_848);
nand U1239 (N_1239,In_471,In_1057);
nor U1240 (N_1240,In_1364,In_1086);
or U1241 (N_1241,In_1196,In_518);
nor U1242 (N_1242,In_82,In_506);
nand U1243 (N_1243,In_61,In_1446);
nor U1244 (N_1244,In_717,In_872);
xnor U1245 (N_1245,In_372,In_837);
and U1246 (N_1246,In_157,In_326);
and U1247 (N_1247,In_1465,In_324);
and U1248 (N_1248,In_1014,In_592);
or U1249 (N_1249,In_227,In_1085);
or U1250 (N_1250,In_1216,In_869);
nor U1251 (N_1251,In_105,In_207);
nand U1252 (N_1252,In_116,In_922);
or U1253 (N_1253,In_1255,In_518);
nand U1254 (N_1254,In_75,In_356);
or U1255 (N_1255,In_174,In_487);
or U1256 (N_1256,In_273,In_635);
nor U1257 (N_1257,In_646,In_49);
nand U1258 (N_1258,In_948,In_1494);
nand U1259 (N_1259,In_325,In_417);
nor U1260 (N_1260,In_812,In_275);
nor U1261 (N_1261,In_1062,In_1489);
or U1262 (N_1262,In_846,In_897);
nor U1263 (N_1263,In_1082,In_662);
and U1264 (N_1264,In_968,In_1194);
nor U1265 (N_1265,In_192,In_951);
nor U1266 (N_1266,In_672,In_1417);
nand U1267 (N_1267,In_16,In_1025);
nor U1268 (N_1268,In_1167,In_625);
nand U1269 (N_1269,In_1195,In_500);
nor U1270 (N_1270,In_27,In_1424);
and U1271 (N_1271,In_57,In_266);
and U1272 (N_1272,In_1210,In_690);
and U1273 (N_1273,In_956,In_18);
or U1274 (N_1274,In_722,In_976);
nor U1275 (N_1275,In_1213,In_1358);
nand U1276 (N_1276,In_1217,In_1136);
or U1277 (N_1277,In_189,In_485);
or U1278 (N_1278,In_561,In_9);
or U1279 (N_1279,In_1076,In_333);
or U1280 (N_1280,In_905,In_506);
nor U1281 (N_1281,In_75,In_436);
nor U1282 (N_1282,In_1226,In_1120);
nand U1283 (N_1283,In_352,In_1392);
nand U1284 (N_1284,In_848,In_177);
nand U1285 (N_1285,In_493,In_863);
nand U1286 (N_1286,In_1473,In_819);
nand U1287 (N_1287,In_999,In_24);
nand U1288 (N_1288,In_272,In_411);
and U1289 (N_1289,In_486,In_1086);
or U1290 (N_1290,In_654,In_1189);
nor U1291 (N_1291,In_1293,In_1248);
or U1292 (N_1292,In_927,In_16);
or U1293 (N_1293,In_945,In_587);
and U1294 (N_1294,In_393,In_914);
nor U1295 (N_1295,In_1246,In_686);
nand U1296 (N_1296,In_576,In_1469);
nor U1297 (N_1297,In_887,In_1457);
or U1298 (N_1298,In_1249,In_1321);
or U1299 (N_1299,In_1482,In_1496);
and U1300 (N_1300,In_157,In_20);
or U1301 (N_1301,In_1040,In_1073);
nor U1302 (N_1302,In_1257,In_727);
nand U1303 (N_1303,In_341,In_531);
and U1304 (N_1304,In_1099,In_1263);
nand U1305 (N_1305,In_122,In_488);
nand U1306 (N_1306,In_901,In_1294);
nand U1307 (N_1307,In_1089,In_530);
nor U1308 (N_1308,In_1163,In_849);
nor U1309 (N_1309,In_890,In_435);
nand U1310 (N_1310,In_187,In_921);
nand U1311 (N_1311,In_133,In_1367);
or U1312 (N_1312,In_29,In_173);
and U1313 (N_1313,In_1211,In_564);
or U1314 (N_1314,In_1159,In_129);
or U1315 (N_1315,In_200,In_1319);
nand U1316 (N_1316,In_18,In_1209);
nand U1317 (N_1317,In_30,In_511);
nand U1318 (N_1318,In_64,In_423);
and U1319 (N_1319,In_605,In_648);
nor U1320 (N_1320,In_991,In_431);
or U1321 (N_1321,In_995,In_580);
and U1322 (N_1322,In_1199,In_297);
nand U1323 (N_1323,In_29,In_1336);
nor U1324 (N_1324,In_395,In_1184);
nor U1325 (N_1325,In_758,In_588);
nor U1326 (N_1326,In_501,In_602);
nand U1327 (N_1327,In_1215,In_151);
nand U1328 (N_1328,In_608,In_122);
and U1329 (N_1329,In_1432,In_1379);
or U1330 (N_1330,In_791,In_41);
nor U1331 (N_1331,In_605,In_694);
and U1332 (N_1332,In_755,In_797);
and U1333 (N_1333,In_762,In_348);
or U1334 (N_1334,In_12,In_212);
nor U1335 (N_1335,In_4,In_766);
nor U1336 (N_1336,In_202,In_776);
nor U1337 (N_1337,In_1412,In_587);
nand U1338 (N_1338,In_1353,In_349);
nand U1339 (N_1339,In_83,In_1183);
or U1340 (N_1340,In_350,In_1457);
or U1341 (N_1341,In_950,In_925);
or U1342 (N_1342,In_230,In_1448);
nor U1343 (N_1343,In_526,In_636);
nand U1344 (N_1344,In_922,In_132);
nand U1345 (N_1345,In_312,In_749);
nand U1346 (N_1346,In_798,In_200);
or U1347 (N_1347,In_199,In_173);
nor U1348 (N_1348,In_803,In_710);
nor U1349 (N_1349,In_790,In_832);
and U1350 (N_1350,In_1103,In_972);
and U1351 (N_1351,In_794,In_1038);
nand U1352 (N_1352,In_1336,In_273);
and U1353 (N_1353,In_48,In_785);
nor U1354 (N_1354,In_1372,In_462);
nand U1355 (N_1355,In_522,In_1186);
nand U1356 (N_1356,In_907,In_496);
or U1357 (N_1357,In_307,In_416);
nand U1358 (N_1358,In_546,In_473);
or U1359 (N_1359,In_1228,In_825);
nand U1360 (N_1360,In_489,In_1);
or U1361 (N_1361,In_570,In_21);
nor U1362 (N_1362,In_1411,In_331);
and U1363 (N_1363,In_1415,In_1437);
and U1364 (N_1364,In_85,In_79);
nor U1365 (N_1365,In_394,In_1493);
nor U1366 (N_1366,In_1097,In_229);
and U1367 (N_1367,In_414,In_876);
or U1368 (N_1368,In_403,In_1278);
nand U1369 (N_1369,In_1462,In_1376);
or U1370 (N_1370,In_1021,In_223);
or U1371 (N_1371,In_753,In_1046);
or U1372 (N_1372,In_834,In_1280);
and U1373 (N_1373,In_106,In_1385);
and U1374 (N_1374,In_945,In_1347);
nand U1375 (N_1375,In_855,In_209);
nand U1376 (N_1376,In_740,In_1313);
nor U1377 (N_1377,In_304,In_827);
nor U1378 (N_1378,In_709,In_917);
nand U1379 (N_1379,In_1340,In_1338);
or U1380 (N_1380,In_193,In_1170);
nand U1381 (N_1381,In_13,In_788);
and U1382 (N_1382,In_456,In_1165);
nor U1383 (N_1383,In_647,In_209);
and U1384 (N_1384,In_462,In_875);
or U1385 (N_1385,In_1014,In_826);
xnor U1386 (N_1386,In_194,In_47);
nor U1387 (N_1387,In_68,In_93);
nand U1388 (N_1388,In_1436,In_701);
or U1389 (N_1389,In_868,In_379);
and U1390 (N_1390,In_613,In_1026);
or U1391 (N_1391,In_1337,In_23);
or U1392 (N_1392,In_609,In_1022);
xnor U1393 (N_1393,In_650,In_480);
nand U1394 (N_1394,In_1335,In_1315);
nand U1395 (N_1395,In_1166,In_139);
nor U1396 (N_1396,In_855,In_1295);
nand U1397 (N_1397,In_1077,In_262);
nor U1398 (N_1398,In_1226,In_427);
nand U1399 (N_1399,In_1146,In_187);
and U1400 (N_1400,In_1175,In_555);
and U1401 (N_1401,In_1438,In_260);
nor U1402 (N_1402,In_1376,In_448);
or U1403 (N_1403,In_1192,In_455);
and U1404 (N_1404,In_949,In_901);
nor U1405 (N_1405,In_1450,In_269);
nor U1406 (N_1406,In_881,In_592);
and U1407 (N_1407,In_588,In_519);
or U1408 (N_1408,In_1199,In_65);
nor U1409 (N_1409,In_593,In_805);
nand U1410 (N_1410,In_1048,In_759);
and U1411 (N_1411,In_1045,In_774);
nor U1412 (N_1412,In_393,In_977);
nor U1413 (N_1413,In_1077,In_1495);
nand U1414 (N_1414,In_582,In_40);
nor U1415 (N_1415,In_1442,In_1118);
and U1416 (N_1416,In_675,In_592);
or U1417 (N_1417,In_1467,In_1368);
nor U1418 (N_1418,In_1018,In_830);
and U1419 (N_1419,In_1320,In_245);
and U1420 (N_1420,In_611,In_36);
and U1421 (N_1421,In_200,In_1239);
or U1422 (N_1422,In_1411,In_967);
nand U1423 (N_1423,In_714,In_1177);
nand U1424 (N_1424,In_485,In_1255);
xnor U1425 (N_1425,In_1457,In_417);
nand U1426 (N_1426,In_279,In_168);
and U1427 (N_1427,In_1087,In_289);
and U1428 (N_1428,In_564,In_1274);
and U1429 (N_1429,In_1000,In_1030);
and U1430 (N_1430,In_831,In_1445);
nand U1431 (N_1431,In_696,In_407);
nor U1432 (N_1432,In_1485,In_1115);
nand U1433 (N_1433,In_603,In_635);
or U1434 (N_1434,In_1252,In_410);
or U1435 (N_1435,In_603,In_507);
nand U1436 (N_1436,In_7,In_891);
nand U1437 (N_1437,In_653,In_338);
nand U1438 (N_1438,In_651,In_1286);
nor U1439 (N_1439,In_626,In_657);
nand U1440 (N_1440,In_646,In_1281);
and U1441 (N_1441,In_1469,In_1306);
nor U1442 (N_1442,In_1310,In_1301);
or U1443 (N_1443,In_415,In_655);
nor U1444 (N_1444,In_677,In_346);
nand U1445 (N_1445,In_361,In_1406);
nand U1446 (N_1446,In_1446,In_815);
nand U1447 (N_1447,In_1083,In_728);
and U1448 (N_1448,In_627,In_602);
nand U1449 (N_1449,In_570,In_3);
nor U1450 (N_1450,In_418,In_933);
or U1451 (N_1451,In_793,In_1452);
nor U1452 (N_1452,In_848,In_463);
or U1453 (N_1453,In_496,In_1171);
or U1454 (N_1454,In_1068,In_976);
nor U1455 (N_1455,In_476,In_558);
or U1456 (N_1456,In_342,In_1299);
and U1457 (N_1457,In_641,In_1244);
nor U1458 (N_1458,In_589,In_1368);
or U1459 (N_1459,In_1144,In_759);
nor U1460 (N_1460,In_307,In_717);
nand U1461 (N_1461,In_571,In_851);
nand U1462 (N_1462,In_244,In_699);
nor U1463 (N_1463,In_895,In_237);
nand U1464 (N_1464,In_339,In_864);
nand U1465 (N_1465,In_1384,In_1107);
nor U1466 (N_1466,In_1365,In_506);
or U1467 (N_1467,In_188,In_1430);
and U1468 (N_1468,In_1478,In_3);
and U1469 (N_1469,In_726,In_655);
and U1470 (N_1470,In_585,In_1400);
and U1471 (N_1471,In_1379,In_321);
and U1472 (N_1472,In_550,In_995);
nor U1473 (N_1473,In_602,In_936);
or U1474 (N_1474,In_1201,In_619);
nor U1475 (N_1475,In_396,In_1172);
and U1476 (N_1476,In_333,In_798);
nor U1477 (N_1477,In_281,In_254);
and U1478 (N_1478,In_214,In_1210);
or U1479 (N_1479,In_741,In_403);
nand U1480 (N_1480,In_26,In_1300);
nand U1481 (N_1481,In_1136,In_63);
and U1482 (N_1482,In_501,In_1249);
nand U1483 (N_1483,In_618,In_840);
nor U1484 (N_1484,In_894,In_975);
nor U1485 (N_1485,In_535,In_970);
nand U1486 (N_1486,In_1054,In_1068);
or U1487 (N_1487,In_489,In_690);
nand U1488 (N_1488,In_601,In_1108);
or U1489 (N_1489,In_646,In_379);
or U1490 (N_1490,In_870,In_778);
nand U1491 (N_1491,In_46,In_1037);
nor U1492 (N_1492,In_1052,In_1307);
nand U1493 (N_1493,In_420,In_1198);
nor U1494 (N_1494,In_217,In_364);
and U1495 (N_1495,In_797,In_758);
nor U1496 (N_1496,In_518,In_1061);
and U1497 (N_1497,In_940,In_830);
or U1498 (N_1498,In_396,In_325);
or U1499 (N_1499,In_1414,In_50);
and U1500 (N_1500,N_1245,N_80);
and U1501 (N_1501,N_679,N_945);
or U1502 (N_1502,N_1164,N_1086);
or U1503 (N_1503,N_6,N_135);
and U1504 (N_1504,N_215,N_1088);
nor U1505 (N_1505,N_783,N_587);
or U1506 (N_1506,N_568,N_1497);
and U1507 (N_1507,N_136,N_529);
and U1508 (N_1508,N_506,N_1243);
and U1509 (N_1509,N_315,N_362);
or U1510 (N_1510,N_249,N_320);
nand U1511 (N_1511,N_865,N_387);
and U1512 (N_1512,N_1343,N_752);
and U1513 (N_1513,N_98,N_173);
and U1514 (N_1514,N_629,N_475);
nand U1515 (N_1515,N_1479,N_318);
nand U1516 (N_1516,N_672,N_862);
or U1517 (N_1517,N_429,N_1242);
and U1518 (N_1518,N_470,N_533);
nand U1519 (N_1519,N_992,N_145);
and U1520 (N_1520,N_1252,N_877);
or U1521 (N_1521,N_1004,N_831);
or U1522 (N_1522,N_159,N_511);
or U1523 (N_1523,N_1454,N_282);
and U1524 (N_1524,N_122,N_123);
nor U1525 (N_1525,N_1420,N_1030);
nand U1526 (N_1526,N_1101,N_346);
and U1527 (N_1527,N_644,N_896);
and U1528 (N_1528,N_422,N_1283);
or U1529 (N_1529,N_182,N_171);
and U1530 (N_1530,N_786,N_332);
nor U1531 (N_1531,N_289,N_1264);
nor U1532 (N_1532,N_1147,N_298);
nand U1533 (N_1533,N_1150,N_925);
nor U1534 (N_1534,N_1351,N_868);
or U1535 (N_1535,N_348,N_360);
nor U1536 (N_1536,N_307,N_707);
or U1537 (N_1537,N_26,N_1319);
nand U1538 (N_1538,N_915,N_1160);
nand U1539 (N_1539,N_1445,N_833);
nand U1540 (N_1540,N_499,N_764);
nor U1541 (N_1541,N_1492,N_151);
and U1542 (N_1542,N_848,N_652);
and U1543 (N_1543,N_1300,N_1165);
nand U1544 (N_1544,N_258,N_818);
nor U1545 (N_1545,N_325,N_857);
nand U1546 (N_1546,N_690,N_932);
or U1547 (N_1547,N_460,N_542);
or U1548 (N_1548,N_1034,N_402);
nand U1549 (N_1549,N_948,N_727);
nand U1550 (N_1550,N_699,N_1281);
nand U1551 (N_1551,N_166,N_1026);
and U1552 (N_1552,N_381,N_793);
nand U1553 (N_1553,N_850,N_1382);
or U1554 (N_1554,N_1306,N_751);
nor U1555 (N_1555,N_3,N_711);
nor U1556 (N_1556,N_639,N_1294);
or U1557 (N_1557,N_0,N_1403);
or U1558 (N_1558,N_227,N_1220);
and U1559 (N_1559,N_95,N_409);
nand U1560 (N_1560,N_1096,N_1366);
nand U1561 (N_1561,N_1452,N_937);
nor U1562 (N_1562,N_1289,N_1200);
nand U1563 (N_1563,N_1464,N_445);
nand U1564 (N_1564,N_1129,N_594);
and U1565 (N_1565,N_243,N_397);
and U1566 (N_1566,N_1120,N_344);
and U1567 (N_1567,N_263,N_434);
and U1568 (N_1568,N_61,N_373);
nor U1569 (N_1569,N_1008,N_112);
or U1570 (N_1570,N_37,N_914);
nor U1571 (N_1571,N_955,N_374);
or U1572 (N_1572,N_438,N_338);
nand U1573 (N_1573,N_247,N_188);
nand U1574 (N_1574,N_428,N_701);
nor U1575 (N_1575,N_1333,N_1203);
and U1576 (N_1576,N_512,N_1254);
nand U1577 (N_1577,N_846,N_461);
or U1578 (N_1578,N_980,N_815);
nor U1579 (N_1579,N_1286,N_1077);
nand U1580 (N_1580,N_59,N_546);
nand U1581 (N_1581,N_109,N_1495);
nand U1582 (N_1582,N_192,N_1483);
nor U1583 (N_1583,N_496,N_847);
or U1584 (N_1584,N_279,N_1419);
nor U1585 (N_1585,N_423,N_83);
nand U1586 (N_1586,N_1353,N_1292);
and U1587 (N_1587,N_820,N_371);
nor U1588 (N_1588,N_216,N_5);
nor U1589 (N_1589,N_114,N_1107);
nor U1590 (N_1590,N_1211,N_294);
nor U1591 (N_1591,N_1131,N_1484);
nand U1592 (N_1592,N_1177,N_432);
nand U1593 (N_1593,N_1100,N_609);
nor U1594 (N_1594,N_796,N_927);
nand U1595 (N_1595,N_899,N_1237);
and U1596 (N_1596,N_745,N_1308);
xor U1597 (N_1597,N_1023,N_177);
and U1598 (N_1598,N_40,N_947);
or U1599 (N_1599,N_991,N_1079);
nand U1600 (N_1600,N_1095,N_798);
nand U1601 (N_1601,N_1036,N_933);
nor U1602 (N_1602,N_1324,N_897);
and U1603 (N_1603,N_558,N_446);
and U1604 (N_1604,N_1146,N_36);
nor U1605 (N_1605,N_984,N_242);
nand U1606 (N_1606,N_1271,N_230);
or U1607 (N_1607,N_465,N_238);
nor U1608 (N_1608,N_363,N_606);
or U1609 (N_1609,N_1209,N_1408);
and U1610 (N_1610,N_839,N_1463);
or U1611 (N_1611,N_125,N_1132);
or U1612 (N_1612,N_1084,N_907);
or U1613 (N_1613,N_27,N_585);
or U1614 (N_1614,N_29,N_401);
nand U1615 (N_1615,N_375,N_1002);
and U1616 (N_1616,N_99,N_1453);
and U1617 (N_1617,N_730,N_368);
or U1618 (N_1618,N_1087,N_1193);
nand U1619 (N_1619,N_1470,N_290);
or U1620 (N_1620,N_142,N_658);
and U1621 (N_1621,N_710,N_882);
and U1622 (N_1622,N_211,N_1066);
or U1623 (N_1623,N_597,N_938);
nand U1624 (N_1624,N_632,N_1094);
nand U1625 (N_1625,N_2,N_525);
and U1626 (N_1626,N_1080,N_874);
and U1627 (N_1627,N_723,N_653);
or U1628 (N_1628,N_1431,N_873);
nor U1629 (N_1629,N_28,N_190);
and U1630 (N_1630,N_769,N_1438);
nand U1631 (N_1631,N_153,N_510);
nand U1632 (N_1632,N_1293,N_1202);
nand U1633 (N_1633,N_271,N_954);
or U1634 (N_1634,N_1191,N_1327);
nand U1635 (N_1635,N_56,N_167);
nor U1636 (N_1636,N_601,N_757);
nor U1637 (N_1637,N_1065,N_256);
or U1638 (N_1638,N_861,N_418);
or U1639 (N_1639,N_508,N_1170);
and U1640 (N_1640,N_891,N_220);
or U1641 (N_1641,N_1093,N_58);
nand U1642 (N_1642,N_305,N_1444);
or U1643 (N_1643,N_715,N_518);
or U1644 (N_1644,N_901,N_185);
or U1645 (N_1645,N_1090,N_931);
nor U1646 (N_1646,N_16,N_453);
and U1647 (N_1647,N_442,N_93);
or U1648 (N_1648,N_19,N_1284);
nand U1649 (N_1649,N_675,N_8);
nor U1650 (N_1650,N_110,N_1450);
or U1651 (N_1651,N_959,N_260);
or U1652 (N_1652,N_547,N_414);
nor U1653 (N_1653,N_49,N_791);
and U1654 (N_1654,N_1236,N_1429);
nor U1655 (N_1655,N_566,N_1447);
nor U1656 (N_1656,N_550,N_553);
nand U1657 (N_1657,N_458,N_281);
and U1658 (N_1658,N_316,N_531);
nand U1659 (N_1659,N_649,N_1285);
and U1660 (N_1660,N_299,N_394);
and U1661 (N_1661,N_398,N_604);
or U1662 (N_1662,N_1223,N_217);
or U1663 (N_1663,N_1109,N_127);
or U1664 (N_1664,N_1265,N_163);
nand U1665 (N_1665,N_1457,N_82);
nor U1666 (N_1666,N_538,N_1486);
or U1667 (N_1667,N_1471,N_1054);
nor U1668 (N_1668,N_656,N_255);
nand U1669 (N_1669,N_666,N_384);
or U1670 (N_1670,N_253,N_1040);
nand U1671 (N_1671,N_48,N_170);
nand U1672 (N_1672,N_1155,N_1375);
and U1673 (N_1673,N_1339,N_1121);
or U1674 (N_1674,N_102,N_700);
or U1675 (N_1675,N_749,N_840);
and U1676 (N_1676,N_1378,N_1033);
nand U1677 (N_1677,N_435,N_495);
or U1678 (N_1678,N_990,N_1348);
or U1679 (N_1679,N_1051,N_1298);
nor U1680 (N_1680,N_1190,N_1325);
nor U1681 (N_1681,N_501,N_822);
nand U1682 (N_1682,N_717,N_214);
nand U1683 (N_1683,N_426,N_702);
or U1684 (N_1684,N_1296,N_934);
and U1685 (N_1685,N_433,N_1031);
nor U1686 (N_1686,N_708,N_459);
nor U1687 (N_1687,N_150,N_1244);
xor U1688 (N_1688,N_235,N_718);
and U1689 (N_1689,N_772,N_244);
nand U1690 (N_1690,N_369,N_199);
nor U1691 (N_1691,N_842,N_548);
or U1692 (N_1692,N_334,N_1276);
nand U1693 (N_1693,N_494,N_1250);
and U1694 (N_1694,N_773,N_448);
and U1695 (N_1695,N_664,N_623);
or U1696 (N_1696,N_1380,N_1393);
or U1697 (N_1697,N_1230,N_541);
or U1698 (N_1698,N_724,N_964);
nand U1699 (N_1699,N_1417,N_330);
nor U1700 (N_1700,N_104,N_1466);
nand U1701 (N_1701,N_1000,N_880);
and U1702 (N_1702,N_1186,N_1239);
nor U1703 (N_1703,N_1421,N_812);
or U1704 (N_1704,N_339,N_795);
nand U1705 (N_1705,N_340,N_578);
or U1706 (N_1706,N_272,N_1459);
or U1707 (N_1707,N_46,N_1003);
nand U1708 (N_1708,N_1161,N_257);
nor U1709 (N_1709,N_1316,N_69);
or U1710 (N_1710,N_1020,N_570);
nand U1711 (N_1711,N_187,N_999);
nand U1712 (N_1712,N_828,N_1398);
nand U1713 (N_1713,N_1210,N_703);
nand U1714 (N_1714,N_799,N_826);
nor U1715 (N_1715,N_302,N_686);
nor U1716 (N_1716,N_1303,N_476);
nand U1717 (N_1717,N_457,N_1422);
or U1718 (N_1718,N_872,N_728);
nor U1719 (N_1719,N_143,N_890);
and U1720 (N_1720,N_1208,N_391);
nand U1721 (N_1721,N_68,N_780);
nor U1722 (N_1722,N_24,N_1342);
nor U1723 (N_1723,N_884,N_583);
or U1724 (N_1724,N_1414,N_1487);
and U1725 (N_1725,N_1169,N_204);
or U1726 (N_1726,N_892,N_906);
nor U1727 (N_1727,N_408,N_107);
nand U1728 (N_1728,N_157,N_160);
and U1729 (N_1729,N_407,N_73);
or U1730 (N_1730,N_1180,N_1355);
nand U1731 (N_1731,N_851,N_678);
and U1732 (N_1732,N_1269,N_1105);
and U1733 (N_1733,N_960,N_837);
nor U1734 (N_1734,N_345,N_834);
xor U1735 (N_1735,N_519,N_579);
nor U1736 (N_1736,N_1061,N_57);
nand U1737 (N_1737,N_1374,N_572);
nor U1738 (N_1738,N_1405,N_1340);
and U1739 (N_1739,N_186,N_1410);
nand U1740 (N_1740,N_50,N_349);
nor U1741 (N_1741,N_264,N_1081);
and U1742 (N_1742,N_403,N_836);
or U1743 (N_1743,N_957,N_844);
nor U1744 (N_1744,N_661,N_673);
or U1745 (N_1745,N_189,N_905);
or U1746 (N_1746,N_638,N_224);
and U1747 (N_1747,N_406,N_329);
or U1748 (N_1748,N_12,N_805);
nor U1749 (N_1749,N_1295,N_813);
or U1750 (N_1750,N_1110,N_592);
nand U1751 (N_1751,N_1145,N_580);
nand U1752 (N_1752,N_477,N_497);
or U1753 (N_1753,N_869,N_76);
or U1754 (N_1754,N_712,N_1038);
nand U1755 (N_1755,N_84,N_1423);
nand U1756 (N_1756,N_787,N_1233);
nand U1757 (N_1757,N_498,N_956);
nand U1758 (N_1758,N_209,N_737);
nand U1759 (N_1759,N_1262,N_935);
nor U1760 (N_1760,N_845,N_981);
nor U1761 (N_1761,N_936,N_1307);
nand U1762 (N_1762,N_1205,N_286);
and U1763 (N_1763,N_74,N_1485);
nor U1764 (N_1764,N_168,N_790);
and U1765 (N_1765,N_1221,N_326);
nand U1766 (N_1766,N_1021,N_1402);
nand U1767 (N_1767,N_467,N_1217);
nand U1768 (N_1768,N_1187,N_9);
or U1769 (N_1769,N_509,N_1213);
or U1770 (N_1770,N_612,N_1028);
and U1771 (N_1771,N_941,N_968);
nor U1772 (N_1772,N_1392,N_917);
and U1773 (N_1773,N_118,N_978);
and U1774 (N_1774,N_450,N_66);
and U1775 (N_1775,N_988,N_1474);
and U1776 (N_1776,N_1019,N_474);
nand U1777 (N_1777,N_288,N_1331);
nor U1778 (N_1778,N_361,N_1256);
or U1779 (N_1779,N_856,N_1416);
and U1780 (N_1780,N_989,N_1199);
or U1781 (N_1781,N_1025,N_676);
and U1782 (N_1782,N_1473,N_1071);
or U1783 (N_1783,N_169,N_888);
nor U1784 (N_1784,N_627,N_91);
or U1785 (N_1785,N_296,N_536);
nand U1786 (N_1786,N_1151,N_79);
or U1787 (N_1787,N_908,N_1427);
nor U1788 (N_1788,N_804,N_1032);
nor U1789 (N_1789,N_1194,N_356);
and U1790 (N_1790,N_327,N_228);
nand U1791 (N_1791,N_1435,N_1389);
or U1792 (N_1792,N_889,N_514);
or U1793 (N_1793,N_101,N_1229);
nand U1794 (N_1794,N_337,N_165);
nor U1795 (N_1795,N_176,N_549);
and U1796 (N_1796,N_400,N_1103);
nand U1797 (N_1797,N_172,N_500);
or U1798 (N_1798,N_1192,N_688);
and U1799 (N_1799,N_376,N_1360);
and U1800 (N_1800,N_1232,N_921);
or U1801 (N_1801,N_1078,N_1070);
or U1802 (N_1802,N_1044,N_912);
and U1803 (N_1803,N_534,N_1171);
and U1804 (N_1804,N_291,N_1130);
and U1805 (N_1805,N_266,N_174);
or U1806 (N_1806,N_424,N_218);
xor U1807 (N_1807,N_270,N_222);
or U1808 (N_1808,N_1060,N_1411);
xnor U1809 (N_1809,N_1490,N_1162);
or U1810 (N_1810,N_939,N_994);
nand U1811 (N_1811,N_567,N_952);
or U1812 (N_1812,N_1489,N_561);
nor U1813 (N_1813,N_1240,N_201);
nor U1814 (N_1814,N_962,N_492);
nor U1815 (N_1815,N_1255,N_807);
nor U1816 (N_1816,N_23,N_1368);
nor U1817 (N_1817,N_1415,N_1461);
or U1818 (N_1818,N_1052,N_1446);
nor U1819 (N_1819,N_382,N_685);
and U1820 (N_1820,N_1041,N_1059);
and U1821 (N_1821,N_449,N_479);
nor U1822 (N_1822,N_823,N_1361);
or U1823 (N_1823,N_1238,N_1207);
and U1824 (N_1824,N_687,N_358);
and U1825 (N_1825,N_949,N_134);
or U1826 (N_1826,N_1451,N_1126);
nor U1827 (N_1827,N_483,N_670);
nand U1828 (N_1828,N_353,N_859);
or U1829 (N_1829,N_1055,N_1072);
nor U1830 (N_1830,N_1228,N_1182);
or U1831 (N_1831,N_54,N_207);
nand U1832 (N_1832,N_589,N_116);
and U1833 (N_1833,N_887,N_559);
and U1834 (N_1834,N_532,N_1321);
or U1835 (N_1835,N_808,N_265);
and U1836 (N_1836,N_343,N_540);
nand U1837 (N_1837,N_146,N_1115);
or U1838 (N_1838,N_1311,N_1323);
and U1839 (N_1839,N_254,N_226);
and U1840 (N_1840,N_181,N_1278);
or U1841 (N_1841,N_65,N_716);
nand U1842 (N_1842,N_208,N_415);
and U1843 (N_1843,N_904,N_827);
nand U1844 (N_1844,N_1179,N_53);
or U1845 (N_1845,N_1369,N_390);
nand U1846 (N_1846,N_1215,N_386);
nand U1847 (N_1847,N_1291,N_755);
and U1848 (N_1848,N_96,N_493);
nand U1849 (N_1849,N_1112,N_1432);
and U1850 (N_1850,N_333,N_997);
or U1851 (N_1851,N_328,N_771);
or U1852 (N_1852,N_1288,N_618);
and U1853 (N_1853,N_669,N_1472);
and U1854 (N_1854,N_1365,N_640);
nand U1855 (N_1855,N_898,N_761);
nand U1856 (N_1856,N_1400,N_473);
nand U1857 (N_1857,N_696,N_814);
or U1858 (N_1858,N_439,N_1035);
nand U1859 (N_1859,N_1124,N_444);
nand U1860 (N_1860,N_645,N_776);
and U1861 (N_1861,N_725,N_1045);
nor U1862 (N_1862,N_193,N_1082);
and U1863 (N_1863,N_194,N_113);
and U1864 (N_1864,N_1449,N_735);
or U1865 (N_1865,N_779,N_748);
or U1866 (N_1866,N_746,N_1477);
nor U1867 (N_1867,N_895,N_87);
and U1868 (N_1868,N_1196,N_359);
or U1869 (N_1869,N_21,N_1394);
nand U1870 (N_1870,N_641,N_1185);
xnor U1871 (N_1871,N_683,N_705);
nor U1872 (N_1872,N_86,N_775);
or U1873 (N_1873,N_636,N_1128);
nand U1874 (N_1874,N_71,N_1277);
nand U1875 (N_1875,N_85,N_1430);
or U1876 (N_1876,N_789,N_240);
nor U1877 (N_1877,N_1274,N_619);
nor U1878 (N_1878,N_1058,N_614);
nor U1879 (N_1879,N_753,N_1290);
nand U1880 (N_1880,N_393,N_692);
nor U1881 (N_1881,N_689,N_367);
and U1882 (N_1882,N_1063,N_33);
and U1883 (N_1883,N_1253,N_794);
nand U1884 (N_1884,N_1068,N_1337);
nor U1885 (N_1885,N_197,N_694);
or U1886 (N_1886,N_385,N_132);
nor U1887 (N_1887,N_293,N_1313);
and U1888 (N_1888,N_1304,N_1143);
and U1889 (N_1889,N_1258,N_563);
nor U1890 (N_1890,N_396,N_262);
and U1891 (N_1891,N_517,N_431);
nor U1892 (N_1892,N_900,N_1388);
xor U1893 (N_1893,N_809,N_1386);
or U1894 (N_1894,N_824,N_156);
nor U1895 (N_1895,N_1302,N_974);
nor U1896 (N_1896,N_383,N_1166);
or U1897 (N_1897,N_1158,N_714);
nor U1898 (N_1898,N_1201,N_45);
and U1899 (N_1899,N_451,N_88);
or U1900 (N_1900,N_1263,N_631);
nand U1901 (N_1901,N_203,N_395);
and U1902 (N_1902,N_950,N_1029);
nand U1903 (N_1903,N_484,N_321);
nand U1904 (N_1904,N_292,N_1279);
nand U1905 (N_1905,N_961,N_357);
nor U1906 (N_1906,N_1106,N_137);
nand U1907 (N_1907,N_565,N_468);
or U1908 (N_1908,N_1475,N_1345);
or U1909 (N_1909,N_10,N_885);
nand U1910 (N_1910,N_1156,N_1049);
nand U1911 (N_1911,N_963,N_1280);
and U1912 (N_1912,N_1122,N_421);
xnor U1913 (N_1913,N_1259,N_743);
or U1914 (N_1914,N_64,N_909);
and U1915 (N_1915,N_1442,N_1048);
nor U1916 (N_1916,N_392,N_51);
nand U1917 (N_1917,N_562,N_1005);
and U1918 (N_1918,N_1257,N_1373);
or U1919 (N_1919,N_624,N_1136);
and U1920 (N_1920,N_237,N_1039);
nand U1921 (N_1921,N_622,N_1440);
and U1922 (N_1922,N_754,N_854);
or U1923 (N_1923,N_1305,N_1225);
and U1924 (N_1924,N_616,N_1141);
nand U1925 (N_1925,N_1067,N_1367);
xnor U1926 (N_1926,N_1317,N_350);
nor U1927 (N_1927,N_34,N_1249);
or U1928 (N_1928,N_1108,N_1);
and U1929 (N_1929,N_605,N_489);
or U1930 (N_1930,N_1496,N_278);
or U1931 (N_1931,N_817,N_1183);
nand U1932 (N_1932,N_259,N_513);
nor U1933 (N_1933,N_505,N_1015);
and U1934 (N_1934,N_1138,N_399);
and U1935 (N_1935,N_731,N_996);
nor U1936 (N_1936,N_31,N_128);
nor U1937 (N_1937,N_317,N_721);
or U1938 (N_1938,N_158,N_552);
and U1939 (N_1939,N_1314,N_1270);
and U1940 (N_1940,N_634,N_835);
or U1941 (N_1941,N_741,N_577);
and U1942 (N_1942,N_760,N_821);
and U1943 (N_1943,N_411,N_767);
or U1944 (N_1944,N_527,N_1123);
nand U1945 (N_1945,N_918,N_1482);
and U1946 (N_1946,N_602,N_681);
nor U1947 (N_1947,N_1214,N_147);
and U1948 (N_1948,N_586,N_312);
or U1949 (N_1949,N_115,N_1175);
nand U1950 (N_1950,N_1409,N_946);
or U1951 (N_1951,N_539,N_1198);
or U1952 (N_1952,N_1467,N_229);
nand U1953 (N_1953,N_706,N_191);
and U1954 (N_1954,N_953,N_599);
nor U1955 (N_1955,N_364,N_1001);
nor U1956 (N_1956,N_858,N_180);
nor U1957 (N_1957,N_929,N_277);
nand U1958 (N_1958,N_1381,N_800);
nor U1959 (N_1959,N_855,N_152);
and U1960 (N_1960,N_853,N_693);
nand U1961 (N_1961,N_677,N_452);
nor U1962 (N_1962,N_1330,N_52);
nand U1963 (N_1963,N_516,N_63);
and U1964 (N_1964,N_736,N_124);
and U1965 (N_1965,N_867,N_1212);
nor U1966 (N_1966,N_674,N_910);
nand U1967 (N_1967,N_979,N_485);
or U1968 (N_1968,N_811,N_1009);
and U1969 (N_1969,N_922,N_1139);
nand U1970 (N_1970,N_309,N_55);
xor U1971 (N_1971,N_301,N_695);
and U1972 (N_1972,N_621,N_1069);
and U1973 (N_1973,N_633,N_1352);
or U1974 (N_1974,N_419,N_902);
nor U1975 (N_1975,N_1178,N_911);
or U1976 (N_1976,N_223,N_117);
or U1977 (N_1977,N_471,N_1493);
or U1978 (N_1978,N_1137,N_967);
or U1979 (N_1979,N_1462,N_744);
and U1980 (N_1980,N_883,N_626);
and U1981 (N_1981,N_1116,N_1406);
nor U1982 (N_1982,N_697,N_43);
nor U1983 (N_1983,N_1251,N_521);
nand U1984 (N_1984,N_841,N_970);
and U1985 (N_1985,N_766,N_1465);
and U1986 (N_1986,N_405,N_860);
and U1987 (N_1987,N_1234,N_491);
nor U1988 (N_1988,N_284,N_1336);
nand U1989 (N_1989,N_179,N_94);
and U1990 (N_1990,N_919,N_261);
nor U1991 (N_1991,N_667,N_441);
and U1992 (N_1992,N_557,N_1455);
nor U1993 (N_1993,N_591,N_1379);
and U1994 (N_1994,N_863,N_665);
nor U1995 (N_1995,N_610,N_221);
nor U1996 (N_1996,N_1387,N_232);
or U1997 (N_1997,N_1359,N_722);
and U1998 (N_1998,N_704,N_1390);
nor U1999 (N_1999,N_588,N_881);
and U2000 (N_2000,N_1152,N_129);
or U2001 (N_2001,N_838,N_89);
nor U2002 (N_2002,N_273,N_141);
and U2003 (N_2003,N_280,N_607);
or U2004 (N_2004,N_1476,N_893);
or U2005 (N_2005,N_269,N_1439);
nand U2006 (N_2006,N_388,N_1142);
nor U2007 (N_2007,N_455,N_782);
or U2008 (N_2008,N_611,N_944);
nand U2009 (N_2009,N_544,N_1266);
and U2010 (N_2010,N_1433,N_1011);
nor U2011 (N_2011,N_600,N_584);
and U2012 (N_2012,N_1231,N_648);
or U2013 (N_2013,N_380,N_574);
and U2014 (N_2014,N_1341,N_200);
nor U2015 (N_2015,N_545,N_322);
or U2016 (N_2016,N_42,N_1469);
nand U2017 (N_2017,N_336,N_971);
or U2018 (N_2018,N_1407,N_870);
or U2019 (N_2019,N_1188,N_758);
nand U2020 (N_2020,N_77,N_225);
nor U2021 (N_2021,N_575,N_903);
or U2022 (N_2022,N_252,N_178);
nor U2023 (N_2023,N_130,N_1372);
or U2024 (N_2024,N_233,N_1356);
nand U2025 (N_2025,N_1260,N_11);
or U2026 (N_2026,N_871,N_515);
nand U2027 (N_2027,N_977,N_788);
and U2028 (N_2028,N_354,N_1006);
nor U2029 (N_2029,N_1144,N_245);
nand U2030 (N_2030,N_430,N_440);
or U2031 (N_2031,N_478,N_1318);
and U2032 (N_2032,N_762,N_90);
nor U2033 (N_2033,N_416,N_982);
nand U2034 (N_2034,N_1272,N_1322);
or U2035 (N_2035,N_366,N_620);
nand U2036 (N_2036,N_487,N_617);
and U2037 (N_2037,N_998,N_377);
and U2038 (N_2038,N_378,N_684);
and U2039 (N_2039,N_105,N_1172);
or U2040 (N_2040,N_7,N_436);
and U2041 (N_2041,N_41,N_643);
and U2042 (N_2042,N_67,N_747);
or U2043 (N_2043,N_1224,N_319);
nand U2044 (N_2044,N_1468,N_139);
nand U2045 (N_2045,N_1099,N_149);
nor U2046 (N_2046,N_819,N_1089);
or U2047 (N_2047,N_195,N_379);
and U2048 (N_2048,N_1309,N_323);
nor U2049 (N_2049,N_1418,N_530);
nor U2050 (N_2050,N_1184,N_781);
nor U2051 (N_2051,N_507,N_1267);
nand U2052 (N_2052,N_965,N_1426);
and U2053 (N_2053,N_32,N_916);
nand U2054 (N_2054,N_966,N_590);
nand U2055 (N_2055,N_729,N_1349);
nor U2056 (N_2056,N_72,N_1007);
or U2057 (N_2057,N_464,N_1370);
nor U2058 (N_2058,N_210,N_1118);
or U2059 (N_2059,N_303,N_285);
nor U2060 (N_2060,N_986,N_973);
or U2061 (N_2061,N_206,N_806);
and U2062 (N_2062,N_1494,N_1085);
and U2063 (N_2063,N_987,N_1062);
and U2064 (N_2064,N_732,N_275);
and U2065 (N_2065,N_1364,N_1301);
and U2066 (N_2066,N_1013,N_22);
and U2067 (N_2067,N_1226,N_1273);
nand U2068 (N_2068,N_1114,N_926);
and U2069 (N_2069,N_1346,N_763);
nand U2070 (N_2070,N_1127,N_35);
and U2071 (N_2071,N_810,N_1261);
and U2072 (N_2072,N_866,N_1074);
or U2073 (N_2073,N_1241,N_1326);
nand U2074 (N_2074,N_1014,N_100);
and U2075 (N_2075,N_1219,N_680);
nor U2076 (N_2076,N_1376,N_138);
nor U2077 (N_2077,N_1363,N_928);
nor U2078 (N_2078,N_297,N_615);
nand U2079 (N_2079,N_1395,N_734);
or U2080 (N_2080,N_886,N_1246);
nor U2081 (N_2081,N_942,N_598);
nand U2082 (N_2082,N_1443,N_843);
and U2083 (N_2083,N_482,N_14);
nand U2084 (N_2084,N_1282,N_196);
nor U2085 (N_2085,N_650,N_162);
or U2086 (N_2086,N_502,N_581);
nor U2087 (N_2087,N_236,N_287);
nor U2088 (N_2088,N_62,N_164);
nand U2089 (N_2089,N_713,N_668);
or U2090 (N_2090,N_4,N_1216);
nand U2091 (N_2091,N_13,N_792);
nor U2092 (N_2092,N_1154,N_556);
nor U2093 (N_2093,N_198,N_573);
nand U2094 (N_2094,N_930,N_662);
nand U2095 (N_2095,N_924,N_1159);
and U2096 (N_2096,N_310,N_1377);
nor U2097 (N_2097,N_276,N_1227);
nor U2098 (N_2098,N_691,N_248);
and U2099 (N_2099,N_231,N_389);
and U2100 (N_2100,N_1498,N_1491);
or U2101 (N_2101,N_1022,N_522);
or U2102 (N_2102,N_646,N_1218);
and U2103 (N_2103,N_103,N_797);
nand U2104 (N_2104,N_1056,N_133);
or U2105 (N_2105,N_1458,N_1133);
or U2106 (N_2106,N_1168,N_698);
nand U2107 (N_2107,N_347,N_1010);
nor U2108 (N_2108,N_1053,N_1396);
nor U2109 (N_2109,N_596,N_535);
and U2110 (N_2110,N_1268,N_503);
nand U2111 (N_2111,N_1092,N_184);
or U2112 (N_2112,N_463,N_1206);
or U2113 (N_2113,N_306,N_410);
nand U2114 (N_2114,N_267,N_106);
nor U2115 (N_2115,N_1204,N_20);
and U2116 (N_2116,N_1017,N_951);
nand U2117 (N_2117,N_969,N_1488);
or U2118 (N_2118,N_995,N_785);
and U2119 (N_2119,N_576,N_148);
nor U2120 (N_2120,N_894,N_1287);
and U2121 (N_2121,N_663,N_1350);
nand U2122 (N_2122,N_1012,N_630);
nand U2123 (N_2123,N_1397,N_1113);
and U2124 (N_2124,N_239,N_1434);
nand U2125 (N_2125,N_308,N_1098);
or U2126 (N_2126,N_720,N_1335);
nor U2127 (N_2127,N_1385,N_923);
or U2128 (N_2128,N_420,N_274);
and U2129 (N_2129,N_1358,N_1425);
nor U2130 (N_2130,N_472,N_342);
nor U2131 (N_2131,N_47,N_603);
and U2132 (N_2132,N_1299,N_1073);
nand U2133 (N_2133,N_1117,N_1413);
or U2134 (N_2134,N_1176,N_830);
and U2135 (N_2135,N_1167,N_311);
or U2136 (N_2136,N_613,N_560);
and U2137 (N_2137,N_976,N_1140);
nand U2138 (N_2138,N_1437,N_756);
or U2139 (N_2139,N_372,N_1027);
nor U2140 (N_2140,N_1157,N_1235);
nor U2141 (N_2141,N_654,N_250);
nand U2142 (N_2142,N_175,N_739);
or U2143 (N_2143,N_647,N_38);
nor U2144 (N_2144,N_111,N_335);
xnor U2145 (N_2145,N_81,N_268);
or U2146 (N_2146,N_15,N_504);
and U2147 (N_2147,N_412,N_1354);
and U2148 (N_2148,N_331,N_1310);
or U2149 (N_2149,N_940,N_1197);
nand U2150 (N_2150,N_456,N_875);
or U2151 (N_2151,N_571,N_1480);
xor U2152 (N_2152,N_30,N_324);
nor U2153 (N_2153,N_300,N_759);
nand U2154 (N_2154,N_341,N_682);
or U2155 (N_2155,N_1499,N_719);
or U2156 (N_2156,N_490,N_219);
nand U2157 (N_2157,N_879,N_1448);
nor U2158 (N_2158,N_803,N_355);
nor U2159 (N_2159,N_593,N_770);
nor U2160 (N_2160,N_283,N_537);
nand U2161 (N_2161,N_120,N_816);
nor U2162 (N_2162,N_778,N_832);
nand U2163 (N_2163,N_543,N_126);
and U2164 (N_2164,N_1371,N_801);
and U2165 (N_2165,N_709,N_1441);
or U2166 (N_2166,N_70,N_60);
and U2167 (N_2167,N_1119,N_205);
nand U2168 (N_2168,N_1057,N_1362);
and U2169 (N_2169,N_183,N_1134);
nor U2170 (N_2170,N_404,N_1018);
nand U2171 (N_2171,N_768,N_314);
and U2172 (N_2172,N_1174,N_993);
or U2173 (N_2173,N_1104,N_628);
or U2174 (N_2174,N_144,N_295);
or U2175 (N_2175,N_983,N_246);
or U2176 (N_2176,N_1338,N_1401);
and U2177 (N_2177,N_738,N_1047);
nor U2178 (N_2178,N_528,N_802);
or U2179 (N_2179,N_523,N_17);
and U2180 (N_2180,N_480,N_608);
nand U2181 (N_2181,N_1163,N_1328);
nand U2182 (N_2182,N_551,N_1412);
or U2183 (N_2183,N_1478,N_1195);
nor U2184 (N_2184,N_659,N_469);
nand U2185 (N_2185,N_1297,N_774);
nor U2186 (N_2186,N_1076,N_765);
and U2187 (N_2187,N_852,N_1111);
or U2188 (N_2188,N_671,N_1247);
nor U2189 (N_2189,N_161,N_75);
nor U2190 (N_2190,N_108,N_1248);
nor U2191 (N_2191,N_78,N_1148);
or U2192 (N_2192,N_1275,N_1383);
or U2193 (N_2193,N_1428,N_425);
or U2194 (N_2194,N_140,N_1091);
nand U2195 (N_2195,N_1149,N_564);
nand U2196 (N_2196,N_876,N_121);
nand U2197 (N_2197,N_1347,N_443);
or U2198 (N_2198,N_975,N_466);
nand U2199 (N_2199,N_1102,N_1456);
or U2200 (N_2200,N_972,N_1075);
and U2201 (N_2201,N_417,N_18);
or U2202 (N_2202,N_554,N_733);
or U2203 (N_2203,N_829,N_750);
nand U2204 (N_2204,N_943,N_1334);
nor U2205 (N_2205,N_1312,N_825);
nor U2206 (N_2206,N_1042,N_251);
and U2207 (N_2207,N_365,N_454);
nor U2208 (N_2208,N_1357,N_1320);
nor U2209 (N_2209,N_726,N_447);
and U2210 (N_2210,N_582,N_241);
nor U2211 (N_2211,N_119,N_1436);
nor U2212 (N_2212,N_520,N_1315);
nand U2213 (N_2213,N_437,N_657);
or U2214 (N_2214,N_524,N_635);
nor U2215 (N_2215,N_742,N_595);
nor U2216 (N_2216,N_1222,N_486);
nor U2217 (N_2217,N_555,N_25);
or U2218 (N_2218,N_212,N_1391);
nor U2219 (N_2219,N_39,N_1125);
nor U2220 (N_2220,N_351,N_155);
nor U2221 (N_2221,N_202,N_1083);
or U2222 (N_2222,N_1050,N_958);
or U2223 (N_2223,N_1135,N_920);
nor U2224 (N_2224,N_660,N_625);
nor U2225 (N_2225,N_526,N_413);
nand U2226 (N_2226,N_1399,N_985);
nor U2227 (N_2227,N_1064,N_864);
and U2228 (N_2228,N_1173,N_427);
nand U2229 (N_2229,N_1024,N_213);
nor U2230 (N_2230,N_1181,N_1424);
nand U2231 (N_2231,N_849,N_488);
or U2232 (N_2232,N_784,N_154);
and U2233 (N_2233,N_1344,N_92);
and U2234 (N_2234,N_878,N_304);
nand U2235 (N_2235,N_1046,N_97);
nor U2236 (N_2236,N_234,N_777);
or U2237 (N_2237,N_1384,N_1016);
nand U2238 (N_2238,N_462,N_651);
xor U2239 (N_2239,N_352,N_740);
or U2240 (N_2240,N_569,N_1481);
nor U2241 (N_2241,N_313,N_481);
nor U2242 (N_2242,N_44,N_913);
nand U2243 (N_2243,N_1460,N_642);
nand U2244 (N_2244,N_1332,N_637);
and U2245 (N_2245,N_1329,N_1404);
or U2246 (N_2246,N_1037,N_131);
and U2247 (N_2247,N_1153,N_370);
nor U2248 (N_2248,N_1189,N_1097);
nand U2249 (N_2249,N_1043,N_655);
or U2250 (N_2250,N_15,N_1186);
and U2251 (N_2251,N_783,N_937);
nor U2252 (N_2252,N_1243,N_665);
or U2253 (N_2253,N_53,N_947);
nand U2254 (N_2254,N_719,N_435);
nor U2255 (N_2255,N_525,N_890);
and U2256 (N_2256,N_1411,N_1266);
and U2257 (N_2257,N_18,N_1396);
nor U2258 (N_2258,N_553,N_1015);
nand U2259 (N_2259,N_1415,N_956);
nor U2260 (N_2260,N_234,N_669);
or U2261 (N_2261,N_544,N_877);
and U2262 (N_2262,N_776,N_591);
or U2263 (N_2263,N_1145,N_1247);
nand U2264 (N_2264,N_841,N_103);
nor U2265 (N_2265,N_585,N_653);
nor U2266 (N_2266,N_416,N_57);
or U2267 (N_2267,N_854,N_1120);
nor U2268 (N_2268,N_999,N_238);
nand U2269 (N_2269,N_1319,N_895);
or U2270 (N_2270,N_259,N_523);
and U2271 (N_2271,N_1190,N_11);
and U2272 (N_2272,N_79,N_742);
or U2273 (N_2273,N_224,N_715);
nand U2274 (N_2274,N_69,N_781);
and U2275 (N_2275,N_270,N_991);
nor U2276 (N_2276,N_1044,N_245);
nand U2277 (N_2277,N_941,N_889);
or U2278 (N_2278,N_693,N_1481);
nand U2279 (N_2279,N_657,N_537);
nor U2280 (N_2280,N_378,N_745);
nand U2281 (N_2281,N_976,N_1441);
nor U2282 (N_2282,N_537,N_1396);
or U2283 (N_2283,N_250,N_1390);
nor U2284 (N_2284,N_92,N_1089);
and U2285 (N_2285,N_113,N_396);
and U2286 (N_2286,N_1104,N_1066);
and U2287 (N_2287,N_1492,N_257);
nand U2288 (N_2288,N_563,N_1279);
nand U2289 (N_2289,N_1196,N_791);
and U2290 (N_2290,N_43,N_814);
nand U2291 (N_2291,N_552,N_1108);
and U2292 (N_2292,N_1212,N_908);
and U2293 (N_2293,N_858,N_857);
nor U2294 (N_2294,N_1117,N_976);
nor U2295 (N_2295,N_792,N_958);
or U2296 (N_2296,N_388,N_286);
nand U2297 (N_2297,N_178,N_1396);
or U2298 (N_2298,N_286,N_326);
and U2299 (N_2299,N_870,N_1401);
nand U2300 (N_2300,N_1468,N_1454);
nand U2301 (N_2301,N_790,N_958);
and U2302 (N_2302,N_930,N_679);
nand U2303 (N_2303,N_23,N_351);
nor U2304 (N_2304,N_1312,N_47);
nor U2305 (N_2305,N_450,N_814);
nand U2306 (N_2306,N_1194,N_1176);
or U2307 (N_2307,N_1070,N_1364);
or U2308 (N_2308,N_844,N_1110);
and U2309 (N_2309,N_249,N_1462);
nand U2310 (N_2310,N_467,N_1463);
nor U2311 (N_2311,N_1262,N_1198);
or U2312 (N_2312,N_186,N_1171);
nand U2313 (N_2313,N_670,N_410);
and U2314 (N_2314,N_589,N_439);
nand U2315 (N_2315,N_1057,N_306);
and U2316 (N_2316,N_811,N_125);
nand U2317 (N_2317,N_178,N_368);
and U2318 (N_2318,N_619,N_1461);
or U2319 (N_2319,N_966,N_818);
nand U2320 (N_2320,N_244,N_1064);
and U2321 (N_2321,N_608,N_996);
nor U2322 (N_2322,N_1355,N_715);
and U2323 (N_2323,N_1210,N_172);
nor U2324 (N_2324,N_105,N_1068);
and U2325 (N_2325,N_1221,N_917);
and U2326 (N_2326,N_1386,N_1147);
or U2327 (N_2327,N_1125,N_11);
nand U2328 (N_2328,N_379,N_1412);
nor U2329 (N_2329,N_242,N_864);
nor U2330 (N_2330,N_920,N_1264);
or U2331 (N_2331,N_736,N_1034);
nand U2332 (N_2332,N_1310,N_1420);
nor U2333 (N_2333,N_1038,N_877);
or U2334 (N_2334,N_1470,N_379);
nand U2335 (N_2335,N_391,N_1303);
nor U2336 (N_2336,N_1299,N_1243);
and U2337 (N_2337,N_193,N_666);
nand U2338 (N_2338,N_1254,N_1068);
or U2339 (N_2339,N_1045,N_1248);
and U2340 (N_2340,N_612,N_406);
or U2341 (N_2341,N_132,N_1333);
nand U2342 (N_2342,N_1239,N_349);
nor U2343 (N_2343,N_581,N_1069);
nand U2344 (N_2344,N_940,N_222);
or U2345 (N_2345,N_289,N_536);
or U2346 (N_2346,N_1366,N_427);
nor U2347 (N_2347,N_1405,N_1008);
and U2348 (N_2348,N_260,N_1317);
and U2349 (N_2349,N_604,N_339);
and U2350 (N_2350,N_1374,N_1465);
or U2351 (N_2351,N_211,N_1108);
nor U2352 (N_2352,N_262,N_1199);
nor U2353 (N_2353,N_563,N_781);
or U2354 (N_2354,N_824,N_24);
and U2355 (N_2355,N_874,N_401);
or U2356 (N_2356,N_1061,N_1393);
or U2357 (N_2357,N_1464,N_549);
and U2358 (N_2358,N_298,N_253);
nand U2359 (N_2359,N_684,N_1323);
or U2360 (N_2360,N_301,N_114);
nor U2361 (N_2361,N_117,N_514);
or U2362 (N_2362,N_933,N_1103);
and U2363 (N_2363,N_692,N_998);
or U2364 (N_2364,N_1208,N_84);
and U2365 (N_2365,N_1426,N_7);
nand U2366 (N_2366,N_404,N_759);
or U2367 (N_2367,N_327,N_1438);
nand U2368 (N_2368,N_891,N_1298);
nand U2369 (N_2369,N_1333,N_1167);
xor U2370 (N_2370,N_1330,N_937);
nor U2371 (N_2371,N_467,N_308);
and U2372 (N_2372,N_441,N_792);
nand U2373 (N_2373,N_476,N_288);
or U2374 (N_2374,N_613,N_1000);
or U2375 (N_2375,N_503,N_551);
and U2376 (N_2376,N_985,N_1278);
or U2377 (N_2377,N_297,N_237);
or U2378 (N_2378,N_1093,N_786);
nand U2379 (N_2379,N_511,N_1308);
nor U2380 (N_2380,N_1297,N_972);
or U2381 (N_2381,N_747,N_194);
nor U2382 (N_2382,N_1185,N_1127);
or U2383 (N_2383,N_656,N_1137);
xnor U2384 (N_2384,N_1404,N_560);
nand U2385 (N_2385,N_1339,N_478);
nand U2386 (N_2386,N_1079,N_1006);
nand U2387 (N_2387,N_206,N_731);
nor U2388 (N_2388,N_521,N_763);
nand U2389 (N_2389,N_326,N_644);
or U2390 (N_2390,N_659,N_144);
nand U2391 (N_2391,N_490,N_1152);
nor U2392 (N_2392,N_83,N_1456);
nand U2393 (N_2393,N_619,N_1232);
and U2394 (N_2394,N_457,N_218);
and U2395 (N_2395,N_1141,N_98);
nand U2396 (N_2396,N_811,N_333);
nor U2397 (N_2397,N_445,N_872);
nand U2398 (N_2398,N_898,N_249);
or U2399 (N_2399,N_1433,N_725);
and U2400 (N_2400,N_1083,N_966);
and U2401 (N_2401,N_828,N_1101);
nand U2402 (N_2402,N_430,N_972);
and U2403 (N_2403,N_1359,N_1435);
and U2404 (N_2404,N_492,N_1218);
or U2405 (N_2405,N_784,N_1255);
nor U2406 (N_2406,N_585,N_451);
nand U2407 (N_2407,N_812,N_623);
and U2408 (N_2408,N_905,N_398);
or U2409 (N_2409,N_49,N_819);
nand U2410 (N_2410,N_789,N_1161);
nor U2411 (N_2411,N_875,N_802);
or U2412 (N_2412,N_606,N_834);
or U2413 (N_2413,N_184,N_1488);
or U2414 (N_2414,N_249,N_548);
or U2415 (N_2415,N_623,N_540);
and U2416 (N_2416,N_1305,N_520);
nand U2417 (N_2417,N_56,N_1309);
nor U2418 (N_2418,N_968,N_1208);
or U2419 (N_2419,N_1328,N_1430);
nand U2420 (N_2420,N_1261,N_453);
nor U2421 (N_2421,N_978,N_703);
nor U2422 (N_2422,N_932,N_698);
nor U2423 (N_2423,N_472,N_605);
or U2424 (N_2424,N_290,N_247);
or U2425 (N_2425,N_436,N_1176);
or U2426 (N_2426,N_366,N_630);
nor U2427 (N_2427,N_517,N_225);
and U2428 (N_2428,N_111,N_516);
and U2429 (N_2429,N_899,N_926);
or U2430 (N_2430,N_386,N_414);
and U2431 (N_2431,N_803,N_216);
nor U2432 (N_2432,N_66,N_524);
nor U2433 (N_2433,N_804,N_787);
and U2434 (N_2434,N_1217,N_1215);
nand U2435 (N_2435,N_1264,N_1000);
nor U2436 (N_2436,N_1098,N_405);
nor U2437 (N_2437,N_1241,N_728);
and U2438 (N_2438,N_1053,N_1285);
or U2439 (N_2439,N_868,N_782);
nor U2440 (N_2440,N_698,N_36);
or U2441 (N_2441,N_1365,N_1372);
and U2442 (N_2442,N_276,N_1012);
or U2443 (N_2443,N_1384,N_1485);
and U2444 (N_2444,N_1267,N_128);
nand U2445 (N_2445,N_310,N_322);
nor U2446 (N_2446,N_683,N_460);
nand U2447 (N_2447,N_581,N_1238);
nand U2448 (N_2448,N_1051,N_1147);
nand U2449 (N_2449,N_820,N_794);
nand U2450 (N_2450,N_1230,N_294);
or U2451 (N_2451,N_1219,N_628);
and U2452 (N_2452,N_669,N_1388);
nand U2453 (N_2453,N_743,N_171);
and U2454 (N_2454,N_681,N_1199);
or U2455 (N_2455,N_1423,N_1015);
nand U2456 (N_2456,N_166,N_1324);
nand U2457 (N_2457,N_1268,N_551);
and U2458 (N_2458,N_1283,N_297);
nand U2459 (N_2459,N_1057,N_962);
nor U2460 (N_2460,N_950,N_254);
and U2461 (N_2461,N_544,N_228);
and U2462 (N_2462,N_643,N_1112);
nor U2463 (N_2463,N_614,N_123);
nand U2464 (N_2464,N_480,N_1242);
nand U2465 (N_2465,N_1204,N_164);
nor U2466 (N_2466,N_185,N_271);
xnor U2467 (N_2467,N_909,N_929);
and U2468 (N_2468,N_438,N_894);
nor U2469 (N_2469,N_1468,N_1372);
nand U2470 (N_2470,N_497,N_128);
nand U2471 (N_2471,N_280,N_1348);
nor U2472 (N_2472,N_933,N_1113);
or U2473 (N_2473,N_1018,N_1318);
nor U2474 (N_2474,N_1105,N_1453);
nand U2475 (N_2475,N_118,N_612);
or U2476 (N_2476,N_649,N_1484);
nor U2477 (N_2477,N_667,N_805);
and U2478 (N_2478,N_534,N_876);
nor U2479 (N_2479,N_1426,N_725);
nand U2480 (N_2480,N_1197,N_723);
and U2481 (N_2481,N_164,N_1035);
nor U2482 (N_2482,N_1174,N_557);
and U2483 (N_2483,N_960,N_331);
or U2484 (N_2484,N_917,N_1287);
and U2485 (N_2485,N_988,N_269);
nand U2486 (N_2486,N_1456,N_1175);
or U2487 (N_2487,N_683,N_545);
and U2488 (N_2488,N_373,N_30);
and U2489 (N_2489,N_206,N_1339);
nor U2490 (N_2490,N_668,N_633);
and U2491 (N_2491,N_685,N_1229);
nor U2492 (N_2492,N_1420,N_139);
nand U2493 (N_2493,N_859,N_506);
or U2494 (N_2494,N_1190,N_752);
or U2495 (N_2495,N_175,N_1017);
nor U2496 (N_2496,N_291,N_852);
and U2497 (N_2497,N_112,N_1322);
nand U2498 (N_2498,N_858,N_697);
nand U2499 (N_2499,N_671,N_916);
nand U2500 (N_2500,N_291,N_968);
or U2501 (N_2501,N_174,N_409);
nand U2502 (N_2502,N_280,N_721);
or U2503 (N_2503,N_892,N_327);
or U2504 (N_2504,N_252,N_352);
nor U2505 (N_2505,N_577,N_1219);
nor U2506 (N_2506,N_1221,N_704);
nor U2507 (N_2507,N_69,N_406);
nor U2508 (N_2508,N_891,N_629);
nand U2509 (N_2509,N_919,N_351);
or U2510 (N_2510,N_70,N_170);
nor U2511 (N_2511,N_525,N_9);
or U2512 (N_2512,N_324,N_375);
nor U2513 (N_2513,N_909,N_808);
or U2514 (N_2514,N_288,N_10);
nand U2515 (N_2515,N_1300,N_686);
or U2516 (N_2516,N_383,N_212);
or U2517 (N_2517,N_49,N_1083);
xnor U2518 (N_2518,N_544,N_515);
or U2519 (N_2519,N_436,N_878);
or U2520 (N_2520,N_1232,N_1061);
nand U2521 (N_2521,N_884,N_35);
or U2522 (N_2522,N_71,N_728);
and U2523 (N_2523,N_56,N_660);
and U2524 (N_2524,N_846,N_375);
and U2525 (N_2525,N_835,N_1474);
nand U2526 (N_2526,N_1197,N_1255);
and U2527 (N_2527,N_1003,N_1254);
and U2528 (N_2528,N_1130,N_417);
nor U2529 (N_2529,N_1165,N_691);
nand U2530 (N_2530,N_1305,N_797);
or U2531 (N_2531,N_148,N_1120);
or U2532 (N_2532,N_816,N_50);
and U2533 (N_2533,N_51,N_448);
and U2534 (N_2534,N_3,N_1260);
nand U2535 (N_2535,N_876,N_197);
nand U2536 (N_2536,N_1304,N_1322);
nor U2537 (N_2537,N_34,N_193);
nand U2538 (N_2538,N_1168,N_704);
or U2539 (N_2539,N_995,N_13);
or U2540 (N_2540,N_907,N_1120);
nand U2541 (N_2541,N_337,N_1417);
and U2542 (N_2542,N_601,N_1372);
nor U2543 (N_2543,N_150,N_257);
nand U2544 (N_2544,N_249,N_316);
nand U2545 (N_2545,N_1129,N_498);
or U2546 (N_2546,N_1253,N_1406);
nor U2547 (N_2547,N_759,N_83);
and U2548 (N_2548,N_166,N_996);
nand U2549 (N_2549,N_675,N_1232);
and U2550 (N_2550,N_579,N_769);
nor U2551 (N_2551,N_761,N_335);
or U2552 (N_2552,N_600,N_1354);
nor U2553 (N_2553,N_697,N_548);
or U2554 (N_2554,N_292,N_12);
and U2555 (N_2555,N_610,N_573);
nor U2556 (N_2556,N_178,N_1014);
nand U2557 (N_2557,N_361,N_1469);
nand U2558 (N_2558,N_1499,N_757);
nor U2559 (N_2559,N_109,N_586);
or U2560 (N_2560,N_1391,N_578);
or U2561 (N_2561,N_729,N_18);
nor U2562 (N_2562,N_1260,N_720);
or U2563 (N_2563,N_795,N_1229);
nor U2564 (N_2564,N_951,N_109);
or U2565 (N_2565,N_274,N_622);
nor U2566 (N_2566,N_716,N_1178);
or U2567 (N_2567,N_394,N_393);
nor U2568 (N_2568,N_535,N_572);
and U2569 (N_2569,N_174,N_1362);
nand U2570 (N_2570,N_979,N_166);
and U2571 (N_2571,N_322,N_739);
and U2572 (N_2572,N_9,N_1459);
and U2573 (N_2573,N_698,N_1095);
or U2574 (N_2574,N_1101,N_1388);
and U2575 (N_2575,N_1456,N_1157);
nand U2576 (N_2576,N_199,N_553);
nand U2577 (N_2577,N_1399,N_1195);
nor U2578 (N_2578,N_552,N_715);
or U2579 (N_2579,N_1339,N_1480);
and U2580 (N_2580,N_939,N_1420);
nor U2581 (N_2581,N_974,N_155);
nand U2582 (N_2582,N_1165,N_1062);
or U2583 (N_2583,N_369,N_1227);
or U2584 (N_2584,N_418,N_1266);
nand U2585 (N_2585,N_390,N_529);
and U2586 (N_2586,N_266,N_133);
nor U2587 (N_2587,N_820,N_188);
or U2588 (N_2588,N_1432,N_497);
nor U2589 (N_2589,N_593,N_219);
nand U2590 (N_2590,N_560,N_574);
or U2591 (N_2591,N_1397,N_733);
and U2592 (N_2592,N_1458,N_564);
and U2593 (N_2593,N_1193,N_485);
or U2594 (N_2594,N_1001,N_723);
or U2595 (N_2595,N_1274,N_841);
or U2596 (N_2596,N_912,N_5);
and U2597 (N_2597,N_538,N_1045);
and U2598 (N_2598,N_666,N_436);
nor U2599 (N_2599,N_1267,N_159);
or U2600 (N_2600,N_1246,N_382);
nor U2601 (N_2601,N_355,N_1096);
and U2602 (N_2602,N_371,N_457);
nand U2603 (N_2603,N_1224,N_1297);
nor U2604 (N_2604,N_855,N_987);
or U2605 (N_2605,N_1042,N_770);
nand U2606 (N_2606,N_339,N_1199);
and U2607 (N_2607,N_210,N_1358);
or U2608 (N_2608,N_86,N_9);
nand U2609 (N_2609,N_873,N_1035);
and U2610 (N_2610,N_548,N_387);
nand U2611 (N_2611,N_99,N_1192);
or U2612 (N_2612,N_298,N_621);
nand U2613 (N_2613,N_1205,N_1068);
and U2614 (N_2614,N_838,N_995);
nor U2615 (N_2615,N_151,N_1482);
or U2616 (N_2616,N_623,N_1040);
nand U2617 (N_2617,N_1395,N_1497);
and U2618 (N_2618,N_1413,N_792);
nor U2619 (N_2619,N_1434,N_34);
nor U2620 (N_2620,N_1260,N_94);
or U2621 (N_2621,N_1496,N_285);
nand U2622 (N_2622,N_1460,N_271);
or U2623 (N_2623,N_240,N_95);
nor U2624 (N_2624,N_768,N_371);
nand U2625 (N_2625,N_10,N_63);
nand U2626 (N_2626,N_1424,N_547);
and U2627 (N_2627,N_218,N_1294);
nor U2628 (N_2628,N_739,N_711);
or U2629 (N_2629,N_1330,N_497);
nor U2630 (N_2630,N_986,N_1234);
nand U2631 (N_2631,N_1363,N_1462);
or U2632 (N_2632,N_142,N_715);
or U2633 (N_2633,N_1120,N_1420);
nand U2634 (N_2634,N_248,N_343);
nor U2635 (N_2635,N_103,N_325);
xnor U2636 (N_2636,N_962,N_498);
or U2637 (N_2637,N_1442,N_256);
and U2638 (N_2638,N_1071,N_287);
nor U2639 (N_2639,N_1448,N_1061);
and U2640 (N_2640,N_330,N_296);
or U2641 (N_2641,N_111,N_1061);
or U2642 (N_2642,N_690,N_185);
and U2643 (N_2643,N_422,N_1449);
or U2644 (N_2644,N_1337,N_1314);
and U2645 (N_2645,N_1078,N_30);
nor U2646 (N_2646,N_168,N_1221);
or U2647 (N_2647,N_846,N_81);
nor U2648 (N_2648,N_1484,N_193);
nand U2649 (N_2649,N_404,N_70);
nor U2650 (N_2650,N_1220,N_68);
or U2651 (N_2651,N_582,N_711);
nand U2652 (N_2652,N_794,N_997);
or U2653 (N_2653,N_475,N_117);
nor U2654 (N_2654,N_1282,N_641);
and U2655 (N_2655,N_995,N_540);
nand U2656 (N_2656,N_472,N_1475);
and U2657 (N_2657,N_1323,N_992);
or U2658 (N_2658,N_903,N_1407);
and U2659 (N_2659,N_102,N_377);
and U2660 (N_2660,N_252,N_359);
nand U2661 (N_2661,N_1475,N_24);
nor U2662 (N_2662,N_1113,N_1215);
nand U2663 (N_2663,N_582,N_636);
or U2664 (N_2664,N_50,N_623);
or U2665 (N_2665,N_474,N_319);
or U2666 (N_2666,N_499,N_941);
nand U2667 (N_2667,N_1313,N_1027);
nor U2668 (N_2668,N_715,N_493);
or U2669 (N_2669,N_919,N_1158);
and U2670 (N_2670,N_328,N_1482);
nand U2671 (N_2671,N_307,N_305);
nor U2672 (N_2672,N_1493,N_310);
and U2673 (N_2673,N_1347,N_607);
and U2674 (N_2674,N_213,N_850);
or U2675 (N_2675,N_880,N_752);
nor U2676 (N_2676,N_748,N_780);
nand U2677 (N_2677,N_549,N_45);
nor U2678 (N_2678,N_1143,N_953);
nand U2679 (N_2679,N_909,N_1400);
or U2680 (N_2680,N_959,N_1435);
or U2681 (N_2681,N_856,N_776);
nor U2682 (N_2682,N_963,N_1350);
or U2683 (N_2683,N_278,N_265);
xnor U2684 (N_2684,N_130,N_1317);
nand U2685 (N_2685,N_541,N_1310);
or U2686 (N_2686,N_1250,N_934);
nand U2687 (N_2687,N_1256,N_1063);
nor U2688 (N_2688,N_1250,N_99);
nand U2689 (N_2689,N_1424,N_1047);
and U2690 (N_2690,N_242,N_918);
nand U2691 (N_2691,N_1415,N_602);
and U2692 (N_2692,N_987,N_1230);
nand U2693 (N_2693,N_870,N_274);
nand U2694 (N_2694,N_686,N_520);
or U2695 (N_2695,N_295,N_1304);
nand U2696 (N_2696,N_1404,N_1034);
and U2697 (N_2697,N_413,N_768);
nand U2698 (N_2698,N_693,N_159);
or U2699 (N_2699,N_642,N_622);
or U2700 (N_2700,N_1180,N_1424);
and U2701 (N_2701,N_963,N_1475);
and U2702 (N_2702,N_1216,N_1049);
and U2703 (N_2703,N_796,N_1294);
and U2704 (N_2704,N_902,N_137);
nand U2705 (N_2705,N_1072,N_667);
or U2706 (N_2706,N_494,N_677);
nand U2707 (N_2707,N_1206,N_1031);
or U2708 (N_2708,N_1491,N_642);
nor U2709 (N_2709,N_491,N_896);
or U2710 (N_2710,N_1414,N_1097);
or U2711 (N_2711,N_1121,N_203);
nand U2712 (N_2712,N_722,N_884);
nor U2713 (N_2713,N_88,N_46);
or U2714 (N_2714,N_616,N_1092);
or U2715 (N_2715,N_1176,N_1436);
nand U2716 (N_2716,N_568,N_1309);
nor U2717 (N_2717,N_419,N_842);
nand U2718 (N_2718,N_629,N_575);
nor U2719 (N_2719,N_223,N_941);
or U2720 (N_2720,N_308,N_838);
or U2721 (N_2721,N_1394,N_709);
nor U2722 (N_2722,N_1170,N_46);
nor U2723 (N_2723,N_1207,N_1494);
and U2724 (N_2724,N_542,N_318);
nor U2725 (N_2725,N_1045,N_674);
nor U2726 (N_2726,N_644,N_362);
or U2727 (N_2727,N_828,N_28);
nor U2728 (N_2728,N_652,N_94);
or U2729 (N_2729,N_679,N_1352);
and U2730 (N_2730,N_1191,N_30);
and U2731 (N_2731,N_1209,N_309);
and U2732 (N_2732,N_892,N_614);
nor U2733 (N_2733,N_209,N_467);
nand U2734 (N_2734,N_429,N_414);
and U2735 (N_2735,N_1307,N_1107);
nand U2736 (N_2736,N_1438,N_861);
and U2737 (N_2737,N_793,N_59);
nand U2738 (N_2738,N_1150,N_812);
or U2739 (N_2739,N_38,N_1344);
and U2740 (N_2740,N_1229,N_1189);
nand U2741 (N_2741,N_719,N_24);
or U2742 (N_2742,N_25,N_518);
nand U2743 (N_2743,N_1044,N_235);
and U2744 (N_2744,N_674,N_707);
or U2745 (N_2745,N_1250,N_935);
nand U2746 (N_2746,N_250,N_134);
or U2747 (N_2747,N_161,N_1460);
nand U2748 (N_2748,N_1039,N_1223);
and U2749 (N_2749,N_396,N_231);
nand U2750 (N_2750,N_44,N_481);
and U2751 (N_2751,N_708,N_1415);
nor U2752 (N_2752,N_228,N_787);
and U2753 (N_2753,N_1215,N_1233);
or U2754 (N_2754,N_676,N_1373);
nor U2755 (N_2755,N_1060,N_272);
nor U2756 (N_2756,N_1370,N_834);
nand U2757 (N_2757,N_1054,N_203);
nor U2758 (N_2758,N_575,N_295);
or U2759 (N_2759,N_108,N_1275);
xnor U2760 (N_2760,N_552,N_794);
nor U2761 (N_2761,N_482,N_620);
nand U2762 (N_2762,N_1058,N_128);
nand U2763 (N_2763,N_465,N_192);
and U2764 (N_2764,N_327,N_1194);
nand U2765 (N_2765,N_944,N_1322);
and U2766 (N_2766,N_429,N_274);
nor U2767 (N_2767,N_227,N_73);
and U2768 (N_2768,N_761,N_1243);
xor U2769 (N_2769,N_663,N_449);
or U2770 (N_2770,N_107,N_212);
or U2771 (N_2771,N_724,N_928);
nor U2772 (N_2772,N_1100,N_765);
nand U2773 (N_2773,N_1023,N_1474);
and U2774 (N_2774,N_805,N_511);
nand U2775 (N_2775,N_577,N_48);
nor U2776 (N_2776,N_583,N_266);
nand U2777 (N_2777,N_661,N_1039);
or U2778 (N_2778,N_934,N_944);
and U2779 (N_2779,N_1493,N_809);
and U2780 (N_2780,N_385,N_1458);
and U2781 (N_2781,N_48,N_775);
nand U2782 (N_2782,N_494,N_1211);
and U2783 (N_2783,N_1311,N_809);
xnor U2784 (N_2784,N_231,N_879);
nor U2785 (N_2785,N_1351,N_841);
and U2786 (N_2786,N_947,N_488);
xor U2787 (N_2787,N_1357,N_1363);
nand U2788 (N_2788,N_445,N_805);
nand U2789 (N_2789,N_1448,N_923);
and U2790 (N_2790,N_714,N_55);
or U2791 (N_2791,N_828,N_1238);
and U2792 (N_2792,N_445,N_1473);
or U2793 (N_2793,N_782,N_1418);
nand U2794 (N_2794,N_558,N_159);
nor U2795 (N_2795,N_739,N_1250);
nand U2796 (N_2796,N_36,N_854);
nand U2797 (N_2797,N_1216,N_666);
nand U2798 (N_2798,N_917,N_790);
nand U2799 (N_2799,N_449,N_1280);
nor U2800 (N_2800,N_570,N_1293);
xnor U2801 (N_2801,N_1398,N_1194);
and U2802 (N_2802,N_429,N_1306);
or U2803 (N_2803,N_1499,N_1348);
and U2804 (N_2804,N_1230,N_23);
and U2805 (N_2805,N_501,N_92);
or U2806 (N_2806,N_1282,N_442);
nand U2807 (N_2807,N_14,N_223);
or U2808 (N_2808,N_176,N_1073);
nand U2809 (N_2809,N_223,N_135);
nor U2810 (N_2810,N_1392,N_634);
nor U2811 (N_2811,N_1479,N_664);
nand U2812 (N_2812,N_695,N_191);
or U2813 (N_2813,N_1250,N_304);
and U2814 (N_2814,N_763,N_1387);
and U2815 (N_2815,N_1412,N_13);
nor U2816 (N_2816,N_268,N_443);
nand U2817 (N_2817,N_257,N_1263);
and U2818 (N_2818,N_125,N_799);
nor U2819 (N_2819,N_207,N_1234);
nor U2820 (N_2820,N_146,N_983);
nand U2821 (N_2821,N_844,N_1173);
and U2822 (N_2822,N_477,N_1212);
or U2823 (N_2823,N_808,N_1465);
or U2824 (N_2824,N_1068,N_1404);
or U2825 (N_2825,N_1305,N_618);
or U2826 (N_2826,N_82,N_1378);
or U2827 (N_2827,N_560,N_1265);
and U2828 (N_2828,N_717,N_1217);
or U2829 (N_2829,N_691,N_391);
or U2830 (N_2830,N_1111,N_1429);
nor U2831 (N_2831,N_548,N_307);
nand U2832 (N_2832,N_1085,N_1372);
and U2833 (N_2833,N_1027,N_340);
nand U2834 (N_2834,N_374,N_312);
and U2835 (N_2835,N_828,N_967);
nor U2836 (N_2836,N_1340,N_31);
and U2837 (N_2837,N_683,N_493);
or U2838 (N_2838,N_1400,N_426);
and U2839 (N_2839,N_724,N_1150);
or U2840 (N_2840,N_1346,N_1048);
nand U2841 (N_2841,N_1380,N_1059);
and U2842 (N_2842,N_1162,N_992);
or U2843 (N_2843,N_547,N_1073);
and U2844 (N_2844,N_933,N_510);
nor U2845 (N_2845,N_636,N_567);
nor U2846 (N_2846,N_853,N_756);
nand U2847 (N_2847,N_234,N_915);
nor U2848 (N_2848,N_624,N_1197);
nand U2849 (N_2849,N_1499,N_9);
or U2850 (N_2850,N_489,N_1479);
or U2851 (N_2851,N_1362,N_1167);
or U2852 (N_2852,N_37,N_512);
and U2853 (N_2853,N_77,N_1170);
and U2854 (N_2854,N_307,N_75);
nor U2855 (N_2855,N_135,N_1443);
or U2856 (N_2856,N_933,N_320);
or U2857 (N_2857,N_689,N_143);
nand U2858 (N_2858,N_1372,N_26);
nand U2859 (N_2859,N_614,N_1013);
and U2860 (N_2860,N_835,N_1304);
nor U2861 (N_2861,N_658,N_716);
and U2862 (N_2862,N_1108,N_924);
nor U2863 (N_2863,N_475,N_1000);
and U2864 (N_2864,N_695,N_1123);
or U2865 (N_2865,N_507,N_150);
or U2866 (N_2866,N_1400,N_885);
xnor U2867 (N_2867,N_44,N_1260);
nor U2868 (N_2868,N_453,N_1430);
and U2869 (N_2869,N_1087,N_458);
and U2870 (N_2870,N_1416,N_1051);
nand U2871 (N_2871,N_29,N_715);
or U2872 (N_2872,N_703,N_1460);
nor U2873 (N_2873,N_1122,N_1105);
nor U2874 (N_2874,N_958,N_170);
nand U2875 (N_2875,N_41,N_801);
nor U2876 (N_2876,N_1419,N_958);
nor U2877 (N_2877,N_328,N_670);
nor U2878 (N_2878,N_1323,N_793);
nor U2879 (N_2879,N_1286,N_101);
or U2880 (N_2880,N_513,N_35);
nor U2881 (N_2881,N_311,N_150);
or U2882 (N_2882,N_1434,N_1216);
or U2883 (N_2883,N_657,N_404);
nor U2884 (N_2884,N_561,N_537);
or U2885 (N_2885,N_686,N_442);
nand U2886 (N_2886,N_1301,N_249);
or U2887 (N_2887,N_172,N_448);
nand U2888 (N_2888,N_576,N_996);
nand U2889 (N_2889,N_1035,N_471);
and U2890 (N_2890,N_916,N_1011);
and U2891 (N_2891,N_8,N_1233);
nand U2892 (N_2892,N_646,N_1026);
or U2893 (N_2893,N_1459,N_426);
or U2894 (N_2894,N_306,N_803);
nor U2895 (N_2895,N_29,N_1291);
nand U2896 (N_2896,N_1183,N_675);
and U2897 (N_2897,N_945,N_1393);
and U2898 (N_2898,N_1274,N_848);
and U2899 (N_2899,N_1409,N_1091);
nor U2900 (N_2900,N_798,N_789);
and U2901 (N_2901,N_792,N_1104);
and U2902 (N_2902,N_149,N_628);
nand U2903 (N_2903,N_1499,N_422);
nor U2904 (N_2904,N_487,N_671);
or U2905 (N_2905,N_59,N_1272);
or U2906 (N_2906,N_576,N_1460);
or U2907 (N_2907,N_450,N_339);
nand U2908 (N_2908,N_956,N_598);
and U2909 (N_2909,N_447,N_1266);
or U2910 (N_2910,N_585,N_1264);
and U2911 (N_2911,N_437,N_498);
or U2912 (N_2912,N_437,N_722);
and U2913 (N_2913,N_1182,N_1261);
nor U2914 (N_2914,N_607,N_1158);
xor U2915 (N_2915,N_897,N_1308);
nand U2916 (N_2916,N_1275,N_854);
nand U2917 (N_2917,N_650,N_454);
nor U2918 (N_2918,N_1088,N_359);
and U2919 (N_2919,N_444,N_154);
nor U2920 (N_2920,N_1449,N_519);
nand U2921 (N_2921,N_1434,N_222);
nor U2922 (N_2922,N_741,N_396);
and U2923 (N_2923,N_921,N_1422);
or U2924 (N_2924,N_1181,N_1081);
and U2925 (N_2925,N_773,N_1111);
and U2926 (N_2926,N_16,N_797);
nor U2927 (N_2927,N_1160,N_94);
nor U2928 (N_2928,N_822,N_770);
or U2929 (N_2929,N_1153,N_436);
and U2930 (N_2930,N_898,N_9);
and U2931 (N_2931,N_1293,N_457);
nand U2932 (N_2932,N_1308,N_40);
nand U2933 (N_2933,N_1152,N_568);
and U2934 (N_2934,N_323,N_771);
nor U2935 (N_2935,N_471,N_777);
nand U2936 (N_2936,N_1288,N_321);
or U2937 (N_2937,N_627,N_631);
and U2938 (N_2938,N_155,N_54);
nand U2939 (N_2939,N_811,N_1279);
and U2940 (N_2940,N_439,N_86);
nor U2941 (N_2941,N_522,N_1106);
or U2942 (N_2942,N_1498,N_778);
nor U2943 (N_2943,N_1005,N_935);
and U2944 (N_2944,N_314,N_1227);
nand U2945 (N_2945,N_1457,N_1479);
or U2946 (N_2946,N_154,N_294);
and U2947 (N_2947,N_756,N_718);
nor U2948 (N_2948,N_788,N_939);
or U2949 (N_2949,N_1155,N_1087);
nor U2950 (N_2950,N_1363,N_1045);
nor U2951 (N_2951,N_221,N_1225);
nor U2952 (N_2952,N_819,N_296);
nand U2953 (N_2953,N_897,N_348);
or U2954 (N_2954,N_975,N_163);
and U2955 (N_2955,N_688,N_740);
nor U2956 (N_2956,N_543,N_1054);
nand U2957 (N_2957,N_528,N_286);
nand U2958 (N_2958,N_25,N_888);
or U2959 (N_2959,N_812,N_62);
or U2960 (N_2960,N_1440,N_1451);
nand U2961 (N_2961,N_1445,N_988);
nand U2962 (N_2962,N_980,N_782);
and U2963 (N_2963,N_357,N_184);
or U2964 (N_2964,N_1214,N_905);
nand U2965 (N_2965,N_216,N_313);
nand U2966 (N_2966,N_969,N_653);
nand U2967 (N_2967,N_193,N_878);
and U2968 (N_2968,N_761,N_57);
or U2969 (N_2969,N_725,N_1107);
or U2970 (N_2970,N_1451,N_410);
nor U2971 (N_2971,N_1257,N_1496);
and U2972 (N_2972,N_952,N_905);
nor U2973 (N_2973,N_446,N_1032);
or U2974 (N_2974,N_519,N_1368);
nor U2975 (N_2975,N_800,N_248);
nor U2976 (N_2976,N_1245,N_365);
or U2977 (N_2977,N_1171,N_939);
nor U2978 (N_2978,N_1262,N_617);
and U2979 (N_2979,N_417,N_149);
and U2980 (N_2980,N_72,N_1363);
and U2981 (N_2981,N_294,N_599);
or U2982 (N_2982,N_789,N_214);
and U2983 (N_2983,N_395,N_1248);
nor U2984 (N_2984,N_427,N_1045);
and U2985 (N_2985,N_211,N_474);
and U2986 (N_2986,N_307,N_991);
and U2987 (N_2987,N_1176,N_1421);
nand U2988 (N_2988,N_524,N_309);
nor U2989 (N_2989,N_950,N_1224);
nor U2990 (N_2990,N_479,N_1173);
or U2991 (N_2991,N_703,N_1008);
nor U2992 (N_2992,N_410,N_1295);
nand U2993 (N_2993,N_813,N_186);
or U2994 (N_2994,N_228,N_746);
nand U2995 (N_2995,N_633,N_847);
nor U2996 (N_2996,N_1005,N_211);
nor U2997 (N_2997,N_53,N_1040);
and U2998 (N_2998,N_477,N_1002);
and U2999 (N_2999,N_224,N_1123);
nor U3000 (N_3000,N_2169,N_1618);
nand U3001 (N_3001,N_2965,N_2488);
and U3002 (N_3002,N_1676,N_2691);
nor U3003 (N_3003,N_2650,N_2144);
nor U3004 (N_3004,N_2321,N_2643);
nand U3005 (N_3005,N_1641,N_2452);
nor U3006 (N_3006,N_2656,N_2323);
or U3007 (N_3007,N_2127,N_2133);
nand U3008 (N_3008,N_2463,N_2353);
or U3009 (N_3009,N_2423,N_2581);
nand U3010 (N_3010,N_2897,N_2399);
nand U3011 (N_3011,N_2411,N_2555);
and U3012 (N_3012,N_2922,N_1867);
nand U3013 (N_3013,N_2003,N_2453);
or U3014 (N_3014,N_2436,N_1740);
or U3015 (N_3015,N_1525,N_1855);
nand U3016 (N_3016,N_2087,N_2468);
or U3017 (N_3017,N_1577,N_2341);
nand U3018 (N_3018,N_2621,N_2472);
nor U3019 (N_3019,N_1610,N_2794);
nor U3020 (N_3020,N_2545,N_1904);
nor U3021 (N_3021,N_2798,N_1848);
and U3022 (N_3022,N_2601,N_2908);
nand U3023 (N_3023,N_2486,N_1596);
xnor U3024 (N_3024,N_2749,N_2303);
nand U3025 (N_3025,N_2067,N_2597);
or U3026 (N_3026,N_2574,N_1960);
and U3027 (N_3027,N_1861,N_1520);
and U3028 (N_3028,N_2460,N_2276);
nor U3029 (N_3029,N_2782,N_2646);
or U3030 (N_3030,N_1844,N_2311);
or U3031 (N_3031,N_2812,N_2924);
nor U3032 (N_3032,N_1615,N_2790);
nand U3033 (N_3033,N_2520,N_2449);
or U3034 (N_3034,N_2529,N_1812);
nand U3035 (N_3035,N_1672,N_2803);
or U3036 (N_3036,N_1707,N_2700);
and U3037 (N_3037,N_2192,N_2751);
nor U3038 (N_3038,N_1967,N_2204);
nand U3039 (N_3039,N_2179,N_2573);
nor U3040 (N_3040,N_1652,N_1912);
or U3041 (N_3041,N_2333,N_2247);
and U3042 (N_3042,N_1993,N_2838);
and U3043 (N_3043,N_1661,N_2910);
nor U3044 (N_3044,N_2006,N_1738);
nand U3045 (N_3045,N_2930,N_2065);
or U3046 (N_3046,N_2830,N_1764);
or U3047 (N_3047,N_2027,N_2739);
nand U3048 (N_3048,N_2864,N_1626);
nor U3049 (N_3049,N_2148,N_2562);
or U3050 (N_3050,N_2177,N_1851);
and U3051 (N_3051,N_2015,N_2622);
and U3052 (N_3052,N_2318,N_2605);
nor U3053 (N_3053,N_2263,N_1801);
and U3054 (N_3054,N_2270,N_2326);
and U3055 (N_3055,N_1959,N_1826);
or U3056 (N_3056,N_2892,N_2888);
nand U3057 (N_3057,N_2037,N_2957);
and U3058 (N_3058,N_2315,N_1731);
nand U3059 (N_3059,N_1601,N_2858);
nor U3060 (N_3060,N_2603,N_2365);
and U3061 (N_3061,N_1978,N_2776);
nor U3062 (N_3062,N_1905,N_2666);
and U3063 (N_3063,N_2469,N_1706);
and U3064 (N_3064,N_2216,N_2822);
or U3065 (N_3065,N_1581,N_2625);
nand U3066 (N_3066,N_2199,N_2079);
and U3067 (N_3067,N_1933,N_1782);
or U3068 (N_3068,N_1723,N_2450);
and U3069 (N_3069,N_2781,N_2843);
or U3070 (N_3070,N_2648,N_2617);
nor U3071 (N_3071,N_1825,N_2714);
or U3072 (N_3072,N_2939,N_2388);
nor U3073 (N_3073,N_2357,N_2075);
nor U3074 (N_3074,N_2633,N_2147);
and U3075 (N_3075,N_2701,N_1957);
nor U3076 (N_3076,N_2162,N_2498);
nor U3077 (N_3077,N_2461,N_1939);
nor U3078 (N_3078,N_2972,N_1598);
or U3079 (N_3079,N_1646,N_2827);
and U3080 (N_3080,N_1711,N_2733);
nand U3081 (N_3081,N_2506,N_2408);
and U3082 (N_3082,N_2278,N_2538);
nor U3083 (N_3083,N_2268,N_2402);
or U3084 (N_3084,N_1755,N_2122);
and U3085 (N_3085,N_2811,N_2525);
nor U3086 (N_3086,N_2364,N_1657);
nand U3087 (N_3087,N_2481,N_2870);
and U3088 (N_3088,N_2391,N_2308);
nor U3089 (N_3089,N_2835,N_2663);
and U3090 (N_3090,N_1749,N_1669);
and U3091 (N_3091,N_2259,N_2706);
nor U3092 (N_3092,N_2502,N_2026);
nand U3093 (N_3093,N_1504,N_2293);
and U3094 (N_3094,N_2234,N_2890);
nand U3095 (N_3095,N_1971,N_1881);
nand U3096 (N_3096,N_2396,N_2580);
or U3097 (N_3097,N_2630,N_2089);
nor U3098 (N_3098,N_2425,N_1607);
nor U3099 (N_3099,N_2667,N_2119);
nor U3100 (N_3100,N_2334,N_2592);
xor U3101 (N_3101,N_2445,N_1695);
nor U3102 (N_3102,N_1846,N_2677);
or U3103 (N_3103,N_2832,N_2768);
and U3104 (N_3104,N_2310,N_2921);
and U3105 (N_3105,N_2490,N_2915);
nand U3106 (N_3106,N_2505,N_1856);
and U3107 (N_3107,N_2049,N_2418);
and U3108 (N_3108,N_2415,N_1770);
nor U3109 (N_3109,N_2424,N_2126);
and U3110 (N_3110,N_2242,N_1974);
or U3111 (N_3111,N_1759,N_1666);
nor U3112 (N_3112,N_2947,N_1629);
or U3113 (N_3113,N_2245,N_2745);
and U3114 (N_3114,N_2374,N_2657);
nor U3115 (N_3115,N_1945,N_1627);
and U3116 (N_3116,N_2236,N_2211);
nand U3117 (N_3117,N_1976,N_2740);
or U3118 (N_3118,N_1820,N_2807);
and U3119 (N_3119,N_2684,N_2362);
nand U3120 (N_3120,N_2732,N_2635);
and U3121 (N_3121,N_2721,N_2936);
and U3122 (N_3122,N_1886,N_2028);
nand U3123 (N_3123,N_1754,N_2896);
nor U3124 (N_3124,N_1547,N_1563);
and U3125 (N_3125,N_2431,N_1728);
or U3126 (N_3126,N_2419,N_2363);
nor U3127 (N_3127,N_1732,N_1823);
nor U3128 (N_3128,N_1690,N_1704);
and U3129 (N_3129,N_1613,N_1771);
and U3130 (N_3130,N_2379,N_2531);
nand U3131 (N_3131,N_2039,N_2076);
and U3132 (N_3132,N_2096,N_2130);
xnor U3133 (N_3133,N_2381,N_1756);
nand U3134 (N_3134,N_1748,N_2097);
and U3135 (N_3135,N_2715,N_1857);
or U3136 (N_3136,N_1570,N_2029);
and U3137 (N_3137,N_1545,N_2971);
or U3138 (N_3138,N_1818,N_2871);
or U3139 (N_3139,N_2564,N_1784);
and U3140 (N_3140,N_1722,N_2937);
and U3141 (N_3141,N_2779,N_2378);
and U3142 (N_3142,N_1788,N_1936);
or U3143 (N_3143,N_2271,N_2124);
and U3144 (N_3144,N_2865,N_2591);
nor U3145 (N_3145,N_2702,N_2285);
and U3146 (N_3146,N_2705,N_2552);
and U3147 (N_3147,N_2136,N_2101);
nand U3148 (N_3148,N_2874,N_1662);
or U3149 (N_3149,N_1579,N_1860);
or U3150 (N_3150,N_2788,N_1573);
nor U3151 (N_3151,N_2501,N_2058);
xor U3152 (N_3152,N_2135,N_2766);
or U3153 (N_3153,N_2084,N_2833);
nand U3154 (N_3154,N_1864,N_2772);
nand U3155 (N_3155,N_2856,N_1888);
nor U3156 (N_3156,N_1816,N_1724);
and U3157 (N_3157,N_1914,N_1941);
or U3158 (N_3158,N_2291,N_1981);
xor U3159 (N_3159,N_2823,N_2683);
nand U3160 (N_3160,N_2183,N_2482);
nor U3161 (N_3161,N_2241,N_2267);
or U3162 (N_3162,N_1530,N_2227);
xor U3163 (N_3163,N_2763,N_2685);
nor U3164 (N_3164,N_1875,N_1542);
and U3165 (N_3165,N_2462,N_1561);
nor U3166 (N_3166,N_1878,N_1595);
or U3167 (N_3167,N_2283,N_2406);
and U3168 (N_3168,N_2497,N_2593);
nand U3169 (N_3169,N_1638,N_2298);
nand U3170 (N_3170,N_2831,N_2269);
or U3171 (N_3171,N_2180,N_2330);
or U3172 (N_3172,N_2828,N_1997);
nor U3173 (N_3173,N_2933,N_1528);
or U3174 (N_3174,N_2528,N_2273);
nand U3175 (N_3175,N_2149,N_2240);
or U3176 (N_3176,N_2371,N_1813);
and U3177 (N_3177,N_2989,N_2422);
nand U3178 (N_3178,N_2613,N_2035);
nand U3179 (N_3179,N_2111,N_1958);
nor U3180 (N_3180,N_2712,N_2639);
and U3181 (N_3181,N_2343,N_1849);
nor U3182 (N_3182,N_1983,N_1757);
and U3183 (N_3183,N_1510,N_2878);
nor U3184 (N_3184,N_2629,N_1776);
nand U3185 (N_3185,N_2166,N_2647);
nand U3186 (N_3186,N_2530,N_1966);
nand U3187 (N_3187,N_2840,N_2687);
nand U3188 (N_3188,N_1989,N_1691);
and U3189 (N_3189,N_2264,N_2138);
or U3190 (N_3190,N_2140,N_1650);
or U3191 (N_3191,N_2671,N_2641);
nor U3192 (N_3192,N_2404,N_2352);
and U3193 (N_3193,N_1946,N_1558);
nand U3194 (N_3194,N_1847,N_2286);
nand U3195 (N_3195,N_1681,N_2430);
or U3196 (N_3196,N_2172,N_2297);
nor U3197 (N_3197,N_1932,N_1962);
or U3198 (N_3198,N_2756,N_2295);
or U3199 (N_3199,N_1677,N_2351);
or U3200 (N_3200,N_2025,N_1827);
and U3201 (N_3201,N_2917,N_1747);
or U3202 (N_3202,N_2458,N_1972);
and U3203 (N_3203,N_2775,N_2694);
nor U3204 (N_3204,N_2072,N_2350);
nand U3205 (N_3205,N_2061,N_2883);
and U3206 (N_3206,N_2438,N_2727);
and U3207 (N_3207,N_2519,N_2932);
or U3208 (N_3208,N_1639,N_1511);
and U3209 (N_3209,N_2679,N_2281);
or U3210 (N_3210,N_2993,N_2369);
nand U3211 (N_3211,N_2532,N_2880);
or U3212 (N_3212,N_2125,N_1877);
or U3213 (N_3213,N_1645,N_2572);
and U3214 (N_3214,N_2723,N_2959);
or U3215 (N_3215,N_1990,N_1992);
nor U3216 (N_3216,N_1979,N_2439);
nor U3217 (N_3217,N_2158,N_2332);
or U3218 (N_3218,N_2695,N_1947);
and U3219 (N_3219,N_2335,N_2561);
and U3220 (N_3220,N_1567,N_2596);
and U3221 (N_3221,N_2770,N_2475);
nor U3222 (N_3222,N_2217,N_1995);
and U3223 (N_3223,N_2654,N_2595);
and U3224 (N_3224,N_1798,N_1987);
nor U3225 (N_3225,N_2797,N_2673);
nor U3226 (N_3226,N_2214,N_1557);
or U3227 (N_3227,N_2255,N_2219);
and U3228 (N_3228,N_2464,N_1965);
or U3229 (N_3229,N_2307,N_1822);
and U3230 (N_3230,N_2556,N_1665);
nor U3231 (N_3231,N_2547,N_1506);
and U3232 (N_3232,N_2994,N_2952);
nor U3233 (N_3233,N_2022,N_2342);
and U3234 (N_3234,N_2891,N_2550);
or U3235 (N_3235,N_1840,N_2612);
nand U3236 (N_3236,N_2316,N_2886);
nand U3237 (N_3237,N_2692,N_2320);
or U3238 (N_3238,N_2304,N_2730);
or U3239 (N_3239,N_2563,N_2070);
nand U3240 (N_3240,N_2467,N_2394);
nor U3241 (N_3241,N_1741,N_1745);
or U3242 (N_3242,N_2116,N_1929);
nor U3243 (N_3243,N_1658,N_1546);
and U3244 (N_3244,N_1514,N_1744);
or U3245 (N_3245,N_2786,N_2471);
or U3246 (N_3246,N_1964,N_2534);
and U3247 (N_3247,N_2082,N_2287);
or U3248 (N_3248,N_2875,N_2009);
or U3249 (N_3249,N_2748,N_1729);
and U3250 (N_3250,N_2551,N_1642);
nor U3251 (N_3251,N_1508,N_2808);
nand U3252 (N_3252,N_2017,N_2569);
nand U3253 (N_3253,N_2277,N_2454);
or U3254 (N_3254,N_2491,N_1562);
nand U3255 (N_3255,N_1739,N_2544);
nor U3256 (N_3256,N_1513,N_2068);
or U3257 (N_3257,N_2385,N_2305);
nor U3258 (N_3258,N_2750,N_2681);
nand U3259 (N_3259,N_1869,N_2873);
nor U3260 (N_3260,N_2031,N_1519);
or U3261 (N_3261,N_2707,N_1634);
nand U3262 (N_3262,N_2253,N_2095);
nor U3263 (N_3263,N_2642,N_1931);
or U3264 (N_3264,N_1512,N_2852);
nand U3265 (N_3265,N_2905,N_2901);
nand U3266 (N_3266,N_1950,N_2818);
nand U3267 (N_3267,N_2451,N_2187);
or U3268 (N_3268,N_2086,N_2110);
nor U3269 (N_3269,N_1906,N_2688);
nand U3270 (N_3270,N_2405,N_1709);
nand U3271 (N_3271,N_2328,N_2474);
or U3272 (N_3272,N_2115,N_1951);
and U3273 (N_3273,N_2724,N_1783);
nor U3274 (N_3274,N_1921,N_1673);
and U3275 (N_3275,N_2774,N_2817);
and U3276 (N_3276,N_2954,N_2403);
xor U3277 (N_3277,N_2628,N_2173);
and U3278 (N_3278,N_2146,N_2778);
or U3279 (N_3279,N_2210,N_1616);
nor U3280 (N_3280,N_1687,N_2568);
and U3281 (N_3281,N_1725,N_1791);
or U3282 (N_3282,N_2160,N_2213);
or U3283 (N_3283,N_2949,N_1894);
and U3284 (N_3284,N_2645,N_2558);
and U3285 (N_3285,N_2296,N_2393);
nand U3286 (N_3286,N_2982,N_2324);
nor U3287 (N_3287,N_2537,N_2785);
nor U3288 (N_3288,N_1876,N_1643);
nor U3289 (N_3289,N_2670,N_2690);
nor U3290 (N_3290,N_2717,N_2951);
or U3291 (N_3291,N_1780,N_2627);
and U3292 (N_3292,N_1803,N_2644);
nand U3293 (N_3293,N_2893,N_2810);
nand U3294 (N_3294,N_2016,N_2784);
nor U3295 (N_3295,N_2623,N_1517);
nor U3296 (N_3296,N_2984,N_1600);
and U3297 (N_3297,N_2383,N_1539);
nor U3298 (N_3298,N_2361,N_2309);
nor U3299 (N_3299,N_1996,N_1922);
nand U3300 (N_3300,N_1899,N_2877);
or U3301 (N_3301,N_1674,N_2854);
nor U3302 (N_3302,N_2000,N_2791);
nor U3303 (N_3303,N_2163,N_2448);
and U3304 (N_3304,N_1796,N_2652);
and U3305 (N_3305,N_2659,N_1841);
nand U3306 (N_3306,N_1765,N_1663);
and U3307 (N_3307,N_1790,N_2367);
nor U3308 (N_3308,N_2289,N_1719);
nand U3309 (N_3309,N_2985,N_2664);
nor U3310 (N_3310,N_1915,N_2728);
nor U3311 (N_3311,N_1986,N_1938);
nor U3312 (N_3312,N_2539,N_1647);
nand U3313 (N_3313,N_2262,N_2799);
or U3314 (N_3314,N_2631,N_2196);
and U3315 (N_3315,N_2407,N_2608);
or U3316 (N_3316,N_2209,N_1631);
nand U3317 (N_3317,N_2389,N_2510);
nand U3318 (N_3318,N_2226,N_1838);
nand U3319 (N_3319,N_2741,N_2239);
nand U3320 (N_3320,N_2319,N_2536);
or U3321 (N_3321,N_2024,N_2599);
nand U3322 (N_3322,N_1679,N_2237);
nand U3323 (N_3323,N_2703,N_2021);
or U3324 (N_3324,N_2836,N_2429);
and U3325 (N_3325,N_1799,N_2548);
nand U3326 (N_3326,N_2434,N_2384);
nor U3327 (N_3327,N_1735,N_2863);
and U3328 (N_3328,N_2764,N_1830);
or U3329 (N_3329,N_1806,N_2524);
nor U3330 (N_3330,N_1715,N_2566);
or U3331 (N_3331,N_1516,N_2041);
or U3332 (N_3332,N_2988,N_2432);
or U3333 (N_3333,N_2649,N_1943);
nand U3334 (N_3334,N_2198,N_2494);
nand U3335 (N_3335,N_1970,N_1828);
or U3336 (N_3336,N_2946,N_2571);
and U3337 (N_3337,N_1649,N_2195);
and U3338 (N_3338,N_1544,N_2129);
or U3339 (N_3339,N_2256,N_2855);
and U3340 (N_3340,N_2614,N_2996);
nor U3341 (N_3341,N_2800,N_2261);
nand U3342 (N_3342,N_2682,N_2489);
or U3343 (N_3343,N_1608,N_2669);
nand U3344 (N_3344,N_1689,N_1815);
and U3345 (N_3345,N_1742,N_2420);
nand U3346 (N_3346,N_1630,N_2752);
and U3347 (N_3347,N_2493,N_1602);
nand U3348 (N_3348,N_1637,N_2167);
nor U3349 (N_3349,N_2059,N_1696);
nand U3350 (N_3350,N_2911,N_1872);
and U3351 (N_3351,N_1717,N_2934);
or U3352 (N_3352,N_2105,N_2322);
or U3353 (N_3353,N_1761,N_2841);
nor U3354 (N_3354,N_2976,N_2992);
or U3355 (N_3355,N_2746,N_1760);
and U3356 (N_3356,N_2698,N_2624);
nor U3357 (N_3357,N_2182,N_1835);
and U3358 (N_3358,N_1683,N_1590);
or U3359 (N_3359,N_2968,N_1623);
or U3360 (N_3360,N_2912,N_2260);
and U3361 (N_3361,N_2722,N_2280);
nor U3362 (N_3362,N_1895,N_2540);
nand U3363 (N_3363,N_2437,N_2662);
nor U3364 (N_3364,N_1575,N_2963);
and U3365 (N_3365,N_2272,N_2619);
or U3366 (N_3366,N_2773,N_2980);
nand U3367 (N_3367,N_1944,N_2104);
nand U3368 (N_3368,N_2676,N_2373);
and U3369 (N_3369,N_1998,N_1862);
and U3370 (N_3370,N_2206,N_2473);
or U3371 (N_3371,N_1786,N_2184);
and U3372 (N_3372,N_2109,N_2123);
or U3373 (N_3373,N_1656,N_2857);
or U3374 (N_3374,N_1538,N_1699);
and U3375 (N_3375,N_1734,N_2066);
or U3376 (N_3376,N_2274,N_2620);
and U3377 (N_3377,N_2360,N_2386);
nand U3378 (N_3378,N_2761,N_1721);
nor U3379 (N_3379,N_2435,N_2523);
and U3380 (N_3380,N_2159,N_2598);
nand U3381 (N_3381,N_1720,N_1829);
and U3382 (N_3382,N_2584,N_2178);
nor U3383 (N_3383,N_1503,N_2979);
nor U3384 (N_3384,N_1540,N_1926);
nand U3385 (N_3385,N_2056,N_2653);
nand U3386 (N_3386,N_2767,N_1902);
nand U3387 (N_3387,N_1651,N_1660);
or U3388 (N_3388,N_2943,N_1664);
and U3389 (N_3389,N_2758,N_1781);
or U3390 (N_3390,N_2132,N_1777);
and U3391 (N_3391,N_1908,N_2604);
and U3392 (N_3392,N_2114,N_2466);
or U3393 (N_3393,N_1953,N_2678);
nor U3394 (N_3394,N_2983,N_2103);
nor U3395 (N_3395,N_2340,N_2380);
nand U3396 (N_3396,N_2421,N_1807);
nand U3397 (N_3397,N_2668,N_2238);
or U3398 (N_3398,N_2050,N_1527);
and U3399 (N_3399,N_2935,N_2007);
nor U3400 (N_3400,N_2348,N_2073);
and U3401 (N_3401,N_2010,N_1582);
nor U3402 (N_3402,N_2139,N_2977);
nor U3403 (N_3403,N_2969,N_1587);
or U3404 (N_3404,N_2508,N_2141);
nor U3405 (N_3405,N_2521,N_2579);
nand U3406 (N_3406,N_2554,N_2106);
or U3407 (N_3407,N_1963,N_1751);
and U3408 (N_3408,N_2484,N_1583);
or U3409 (N_3409,N_1569,N_2747);
and U3410 (N_3410,N_1554,N_1940);
and U3411 (N_3411,N_1800,N_2013);
and U3412 (N_3412,N_2244,N_1534);
and U3413 (N_3413,N_1773,N_2477);
nor U3414 (N_3414,N_1716,N_2543);
or U3415 (N_3415,N_1622,N_2894);
xor U3416 (N_3416,N_1948,N_1633);
xor U3417 (N_3417,N_2457,N_1743);
nand U3418 (N_3418,N_2314,N_2953);
nor U3419 (N_3419,N_2884,N_2713);
or U3420 (N_3420,N_1833,N_2938);
or U3421 (N_3421,N_1680,N_1507);
nor U3422 (N_3422,N_1584,N_2809);
nor U3423 (N_3423,N_2686,N_1909);
or U3424 (N_3424,N_1712,N_2377);
and U3425 (N_3425,N_2966,N_2522);
nand U3426 (N_3426,N_2233,N_1994);
nor U3427 (N_3427,N_2222,N_1737);
or U3428 (N_3428,N_2459,N_2931);
and U3429 (N_3429,N_2414,N_2736);
and U3430 (N_3430,N_1655,N_1531);
and U3431 (N_3431,N_2825,N_1973);
nand U3432 (N_3432,N_2997,N_1697);
or U3433 (N_3433,N_1714,N_2338);
nand U3434 (N_3434,N_2004,N_2533);
nand U3435 (N_3435,N_2171,N_2063);
or U3436 (N_3436,N_1819,N_2899);
nand U3437 (N_3437,N_2517,N_1795);
and U3438 (N_3438,N_2428,N_2860);
nor U3439 (N_3439,N_2387,N_2588);
nor U3440 (N_3440,N_2229,N_2928);
and U3441 (N_3441,N_1693,N_2476);
or U3442 (N_3442,N_2306,N_2567);
nor U3443 (N_3443,N_2134,N_2853);
and U3444 (N_3444,N_2585,N_2651);
or U3445 (N_3445,N_1576,N_2987);
nand U3446 (N_3446,N_1975,N_2783);
or U3447 (N_3447,N_1518,N_2615);
and U3448 (N_3448,N_2704,N_1515);
and U3449 (N_3449,N_2051,N_2680);
nand U3450 (N_3450,N_2275,N_2602);
nand U3451 (N_3451,N_1809,N_2535);
or U3452 (N_3452,N_1614,N_2046);
nand U3453 (N_3453,N_2478,N_2586);
nand U3454 (N_3454,N_2197,N_2012);
and U3455 (N_3455,N_2176,N_1949);
nand U3456 (N_3456,N_2885,N_1956);
nand U3457 (N_3457,N_2672,N_2327);
and U3458 (N_3458,N_2055,N_1532);
nor U3459 (N_3459,N_1736,N_2409);
nor U3460 (N_3460,N_2057,N_1802);
and U3461 (N_3461,N_2033,N_1644);
and U3462 (N_3462,N_2765,N_2804);
and U3463 (N_3463,N_2030,N_2975);
nand U3464 (N_3464,N_1805,N_2292);
nand U3465 (N_3465,N_2290,N_2094);
xor U3466 (N_3466,N_2720,N_2868);
nand U3467 (N_3467,N_1556,N_2043);
nand U3468 (N_3468,N_2416,N_1678);
nand U3469 (N_3469,N_2401,N_2675);
nand U3470 (N_3470,N_2060,N_2862);
nand U3471 (N_3471,N_1927,N_1866);
and U3472 (N_3472,N_1670,N_1549);
nor U3473 (N_3473,N_1535,N_1935);
and U3474 (N_3474,N_2040,N_1885);
nand U3475 (N_3475,N_2413,N_2882);
nand U3476 (N_3476,N_1636,N_2848);
or U3477 (N_3477,N_2526,N_2844);
nand U3478 (N_3478,N_2689,N_2755);
and U3479 (N_3479,N_2900,N_2907);
and U3480 (N_3480,N_1892,N_2881);
and U3481 (N_3481,N_2153,N_2117);
or U3482 (N_3482,N_2250,N_1701);
nand U3483 (N_3483,N_2231,N_1694);
and U3484 (N_3484,N_2507,N_2802);
nor U3485 (N_3485,N_2045,N_1865);
and U3486 (N_3486,N_1814,N_2339);
and U3487 (N_3487,N_1592,N_2092);
xor U3488 (N_3488,N_2816,N_1811);
or U3489 (N_3489,N_1852,N_2926);
nand U3490 (N_3490,N_2441,N_2560);
or U3491 (N_3491,N_2824,N_2801);
or U3492 (N_3492,N_2071,N_2313);
nand U3493 (N_3493,N_2102,N_1859);
nor U3494 (N_3494,N_1821,N_1917);
xor U3495 (N_3495,N_2834,N_1850);
or U3496 (N_3496,N_1620,N_1889);
or U3497 (N_3497,N_2956,N_2610);
or U3498 (N_3498,N_1836,N_2034);
or U3499 (N_3499,N_2826,N_2193);
or U3500 (N_3500,N_1952,N_2638);
nor U3501 (N_3501,N_2577,N_1916);
nand U3502 (N_3502,N_1928,N_2990);
or U3503 (N_3503,N_2795,N_2837);
nor U3504 (N_3504,N_2819,N_2455);
or U3505 (N_3505,N_1883,N_1873);
nor U3506 (N_3506,N_1937,N_1565);
or U3507 (N_3507,N_1843,N_2175);
nand U3508 (N_3508,N_2375,N_1871);
nor U3509 (N_3509,N_2978,N_2575);
nand U3510 (N_3510,N_2872,N_1900);
or U3511 (N_3511,N_2249,N_2866);
nand U3512 (N_3512,N_2511,N_1934);
or U3513 (N_3513,N_2944,N_2410);
and U3514 (N_3514,N_2549,N_2091);
nor U3515 (N_3515,N_1591,N_1619);
or U3516 (N_3516,N_2587,N_2048);
nor U3517 (N_3517,N_2470,N_1903);
and U3518 (N_3518,N_1523,N_2190);
or U3519 (N_3519,N_1999,N_2496);
nand U3520 (N_3520,N_2083,N_2796);
nand U3521 (N_3521,N_2640,N_1635);
and U3522 (N_3522,N_2142,N_1685);
nor U3523 (N_3523,N_2266,N_2780);
nand U3524 (N_3524,N_2107,N_1555);
nor U3525 (N_3525,N_2074,N_2230);
or U3526 (N_3526,N_1564,N_2443);
or U3527 (N_3527,N_1919,N_1609);
or U3528 (N_3528,N_2557,N_2062);
and U3529 (N_3529,N_1560,N_1671);
and U3530 (N_3530,N_2867,N_2174);
and U3531 (N_3531,N_2235,N_2546);
and U3532 (N_3532,N_2618,N_2787);
and U3533 (N_3533,N_2697,N_1718);
or U3534 (N_3534,N_2194,N_2916);
or U3535 (N_3535,N_1692,N_2927);
nand U3536 (N_3536,N_2081,N_2128);
nor U3537 (N_3537,N_2696,N_2078);
or U3538 (N_3538,N_2516,N_2359);
nor U3539 (N_3539,N_2080,N_1837);
nand U3540 (N_3540,N_2923,N_2077);
or U3541 (N_3541,N_2165,N_2914);
or U3542 (N_3542,N_2356,N_1597);
nor U3543 (N_3543,N_2509,N_2920);
or U3544 (N_3544,N_1611,N_2945);
nor U3545 (N_3545,N_1961,N_1980);
or U3546 (N_3546,N_1891,N_1984);
and U3547 (N_3547,N_1500,N_1551);
nor U3548 (N_3548,N_2246,N_2895);
nor U3549 (N_3549,N_2582,N_1775);
or U3550 (N_3550,N_1785,N_2054);
or U3551 (N_3551,N_2583,N_2941);
nor U3552 (N_3552,N_1804,N_1988);
nand U3553 (N_3553,N_1896,N_2759);
nor U3554 (N_3554,N_1752,N_1529);
nor U3555 (N_3555,N_2479,N_2088);
nand U3556 (N_3556,N_1659,N_2918);
nor U3557 (N_3557,N_2589,N_2312);
and U3558 (N_3558,N_1955,N_1746);
and U3559 (N_3559,N_2215,N_2368);
or U3560 (N_3560,N_1559,N_2252);
nor U3561 (N_3561,N_2186,N_1778);
or U3562 (N_3562,N_1880,N_1668);
nand U3563 (N_3563,N_2734,N_2729);
or U3564 (N_3564,N_2207,N_2578);
nor U3565 (N_3565,N_2738,N_1521);
nor U3566 (N_3566,N_2632,N_2850);
or U3567 (N_3567,N_2805,N_2559);
or U3568 (N_3568,N_2331,N_1787);
and U3569 (N_3569,N_1907,N_1705);
nand U3570 (N_3570,N_1632,N_2861);
or U3571 (N_3571,N_1920,N_1910);
and U3572 (N_3572,N_2150,N_2876);
nand U3573 (N_3573,N_2018,N_1968);
nor U3574 (N_3574,N_2829,N_2869);
nand U3575 (N_3575,N_2433,N_2069);
nand U3576 (N_3576,N_2145,N_2337);
or U3577 (N_3577,N_2299,N_1688);
and U3578 (N_3578,N_2064,N_2036);
nand U3579 (N_3579,N_2121,N_2440);
and U3580 (N_3580,N_1792,N_2336);
nor U3581 (N_3581,N_2228,N_2655);
and U3582 (N_3582,N_1789,N_2973);
and U3583 (N_3583,N_1628,N_2325);
or U3584 (N_3584,N_2929,N_2346);
and U3585 (N_3585,N_1870,N_1654);
and U3586 (N_3586,N_1686,N_1753);
and U3587 (N_3587,N_1586,N_2693);
and U3588 (N_3588,N_2372,N_1923);
nor U3589 (N_3589,N_1969,N_2904);
or U3590 (N_3590,N_1911,N_2634);
nand U3591 (N_3591,N_1703,N_2725);
nand U3592 (N_3592,N_2397,N_2212);
nor U3593 (N_3593,N_2637,N_2913);
and U3594 (N_3594,N_2446,N_2813);
nor U3595 (N_3595,N_2302,N_2020);
and U3596 (N_3596,N_2847,N_2225);
or U3597 (N_3597,N_2376,N_2014);
nand U3598 (N_3598,N_2181,N_1772);
and U3599 (N_3599,N_2300,N_1653);
and U3600 (N_3600,N_2726,N_1794);
and U3601 (N_3601,N_1552,N_1726);
nor U3602 (N_3602,N_2842,N_2754);
and U3603 (N_3603,N_2485,N_1713);
nand U3604 (N_3604,N_2345,N_2925);
nand U3605 (N_3605,N_1991,N_2008);
nand U3606 (N_3606,N_1684,N_2909);
nand U3607 (N_3607,N_2156,N_1750);
or U3608 (N_3608,N_1874,N_2719);
or U3609 (N_3609,N_2108,N_2626);
nand U3610 (N_3610,N_2232,N_1566);
xor U3611 (N_3611,N_1954,N_1700);
nor U3612 (N_3612,N_2185,N_1580);
nand U3613 (N_3613,N_1817,N_2366);
xor U3614 (N_3614,N_2845,N_2518);
or U3615 (N_3615,N_1522,N_1767);
and U3616 (N_3616,N_1768,N_1730);
nand U3617 (N_3617,N_2355,N_1882);
or U3618 (N_3618,N_1733,N_2282);
and U3619 (N_3619,N_2170,N_2742);
or U3620 (N_3620,N_1509,N_1762);
xnor U3621 (N_3621,N_1548,N_1808);
and U3622 (N_3622,N_2998,N_1502);
nor U3623 (N_3623,N_1863,N_2711);
and U3624 (N_3624,N_2962,N_1890);
or U3625 (N_3625,N_2942,N_2958);
nand U3626 (N_3626,N_2201,N_1779);
nor U3627 (N_3627,N_2395,N_2955);
nor U3628 (N_3628,N_2038,N_1572);
nand U3629 (N_3629,N_2168,N_2248);
nor U3630 (N_3630,N_2191,N_2301);
nand U3631 (N_3631,N_2220,N_2223);
nor U3632 (N_3632,N_2793,N_1536);
nand U3633 (N_3633,N_2161,N_1553);
nor U3634 (N_3634,N_2019,N_2757);
or U3635 (N_3635,N_2120,N_2118);
or U3636 (N_3636,N_2771,N_1537);
and U3637 (N_3637,N_2480,N_2131);
or U3638 (N_3638,N_2203,N_2221);
nand U3639 (N_3639,N_2155,N_2042);
and U3640 (N_3640,N_2288,N_2284);
and U3641 (N_3641,N_1588,N_2205);
nor U3642 (N_3642,N_2565,N_1842);
or U3643 (N_3643,N_1612,N_1918);
and U3644 (N_3644,N_2098,N_2344);
and U3645 (N_3645,N_2594,N_2044);
and U3646 (N_3646,N_2789,N_1603);
or U3647 (N_3647,N_2514,N_1571);
nor U3648 (N_3648,N_2504,N_2906);
or U3649 (N_3649,N_1605,N_1593);
nand U3650 (N_3650,N_2814,N_1625);
nor U3651 (N_3651,N_2961,N_2661);
nor U3652 (N_3652,N_1708,N_2390);
or U3653 (N_3653,N_2699,N_1925);
nand U3654 (N_3654,N_2815,N_2735);
and U3655 (N_3655,N_1793,N_2032);
and U3656 (N_3656,N_2294,N_2011);
nand U3657 (N_3657,N_1702,N_2100);
and U3658 (N_3658,N_1698,N_1845);
and U3659 (N_3659,N_1810,N_1854);
and U3660 (N_3660,N_2317,N_1505);
nor U3661 (N_3661,N_2606,N_1853);
and U3662 (N_3662,N_1824,N_2991);
or U3663 (N_3663,N_1648,N_2708);
nor U3664 (N_3664,N_2329,N_2254);
nand U3665 (N_3665,N_2718,N_2887);
or U3666 (N_3666,N_2903,N_2053);
or U3667 (N_3667,N_2821,N_2164);
nor U3668 (N_3668,N_2093,N_1578);
nor U3669 (N_3669,N_1524,N_2553);
nand U3670 (N_3670,N_2113,N_2851);
nor U3671 (N_3671,N_2940,N_2487);
and U3672 (N_3672,N_2417,N_1893);
nand U3673 (N_3673,N_2731,N_2716);
nor U3674 (N_3674,N_2442,N_2005);
nand U3675 (N_3675,N_2354,N_2964);
or U3676 (N_3676,N_1897,N_2710);
or U3677 (N_3677,N_2806,N_2279);
nand U3678 (N_3678,N_1727,N_2099);
and U3679 (N_3679,N_2265,N_1606);
and U3680 (N_3680,N_2218,N_1640);
or U3681 (N_3681,N_1839,N_2743);
nor U3682 (N_3682,N_2513,N_2709);
and U3683 (N_3683,N_1879,N_2570);
nor U3684 (N_3684,N_1913,N_1682);
and U3685 (N_3685,N_2607,N_2085);
nand U3686 (N_3686,N_2889,N_2981);
or U3687 (N_3687,N_2349,N_2737);
nor U3688 (N_3688,N_1501,N_1832);
or U3689 (N_3689,N_2660,N_2849);
nor U3690 (N_3690,N_2358,N_2137);
and U3691 (N_3691,N_2444,N_2967);
and U3692 (N_3692,N_2658,N_2465);
and U3693 (N_3693,N_2541,N_2258);
xor U3694 (N_3694,N_1930,N_2143);
and U3695 (N_3695,N_1550,N_1982);
nand U3696 (N_3696,N_2202,N_2902);
and U3697 (N_3697,N_2152,N_2492);
nand U3698 (N_3698,N_2753,N_2047);
nor U3699 (N_3699,N_2974,N_2839);
or U3700 (N_3700,N_1533,N_1898);
xor U3701 (N_3701,N_2576,N_2769);
nor U3702 (N_3702,N_2636,N_2999);
nor U3703 (N_3703,N_2898,N_2762);
nand U3704 (N_3704,N_2224,N_1769);
nor U3705 (N_3705,N_2590,N_2948);
or U3706 (N_3706,N_2500,N_2512);
nand U3707 (N_3707,N_1667,N_2483);
nand U3708 (N_3708,N_2495,N_2398);
or U3709 (N_3709,N_2447,N_1585);
nand U3710 (N_3710,N_1621,N_2188);
nor U3711 (N_3711,N_1526,N_2200);
nor U3712 (N_3712,N_2002,N_2515);
or U3713 (N_3713,N_2792,N_1884);
and U3714 (N_3714,N_2090,N_2542);
nor U3715 (N_3715,N_1831,N_1599);
or U3716 (N_3716,N_2347,N_2744);
nand U3717 (N_3717,N_1774,N_2257);
and U3718 (N_3718,N_2382,N_1541);
or U3719 (N_3719,N_2616,N_2052);
or U3720 (N_3720,N_1901,N_2665);
or U3721 (N_3721,N_2970,N_2527);
nor U3722 (N_3722,N_2499,N_1675);
nor U3723 (N_3723,N_1924,N_2001);
or U3724 (N_3724,N_2400,N_2950);
nand U3725 (N_3725,N_2251,N_2846);
or U3726 (N_3726,N_2427,N_2426);
nand U3727 (N_3727,N_1985,N_1568);
nor U3728 (N_3728,N_2370,N_1887);
nand U3729 (N_3729,N_2919,N_2392);
or U3730 (N_3730,N_1594,N_2112);
or U3731 (N_3731,N_2154,N_2820);
nor U3732 (N_3732,N_2600,N_1763);
nor U3733 (N_3733,N_2503,N_1589);
and U3734 (N_3734,N_2859,N_2157);
nand U3735 (N_3735,N_2151,N_1604);
nor U3736 (N_3736,N_2879,N_1617);
nand U3737 (N_3737,N_2674,N_1543);
xnor U3738 (N_3738,N_2609,N_2760);
nor U3739 (N_3739,N_2611,N_1858);
nor U3740 (N_3740,N_1710,N_1834);
and U3741 (N_3741,N_2189,N_2243);
xnor U3742 (N_3742,N_1574,N_1797);
or U3743 (N_3743,N_1624,N_2995);
and U3744 (N_3744,N_2023,N_2412);
nor U3745 (N_3745,N_1766,N_2960);
nand U3746 (N_3746,N_1942,N_1868);
and U3747 (N_3747,N_2456,N_2777);
or U3748 (N_3748,N_2208,N_2986);
nor U3749 (N_3749,N_1977,N_1758);
nand U3750 (N_3750,N_2625,N_2611);
or U3751 (N_3751,N_2925,N_2334);
nand U3752 (N_3752,N_2496,N_2837);
or U3753 (N_3753,N_2719,N_2163);
nor U3754 (N_3754,N_2858,N_2013);
or U3755 (N_3755,N_2137,N_1653);
nor U3756 (N_3756,N_1649,N_2356);
nand U3757 (N_3757,N_1540,N_2702);
nand U3758 (N_3758,N_2034,N_2503);
xor U3759 (N_3759,N_2999,N_2425);
nand U3760 (N_3760,N_1984,N_1739);
nand U3761 (N_3761,N_2083,N_2637);
nor U3762 (N_3762,N_1566,N_1698);
and U3763 (N_3763,N_2664,N_1744);
nor U3764 (N_3764,N_2758,N_2448);
nor U3765 (N_3765,N_2228,N_2944);
and U3766 (N_3766,N_1994,N_1998);
nor U3767 (N_3767,N_1583,N_2004);
nand U3768 (N_3768,N_2147,N_2635);
or U3769 (N_3769,N_1820,N_2363);
nor U3770 (N_3770,N_2099,N_1596);
nor U3771 (N_3771,N_2954,N_2944);
nor U3772 (N_3772,N_2289,N_2715);
or U3773 (N_3773,N_2105,N_1729);
or U3774 (N_3774,N_1793,N_2968);
or U3775 (N_3775,N_2501,N_1736);
nor U3776 (N_3776,N_2173,N_1830);
or U3777 (N_3777,N_2124,N_1553);
nor U3778 (N_3778,N_1779,N_2476);
and U3779 (N_3779,N_1910,N_1887);
nor U3780 (N_3780,N_2551,N_2871);
nand U3781 (N_3781,N_2602,N_2106);
and U3782 (N_3782,N_2871,N_2672);
or U3783 (N_3783,N_2480,N_2624);
or U3784 (N_3784,N_2171,N_2364);
or U3785 (N_3785,N_2128,N_2114);
or U3786 (N_3786,N_2086,N_2736);
and U3787 (N_3787,N_1841,N_2218);
nor U3788 (N_3788,N_2577,N_1897);
nand U3789 (N_3789,N_1878,N_2892);
nand U3790 (N_3790,N_1754,N_1917);
nor U3791 (N_3791,N_2829,N_1547);
and U3792 (N_3792,N_2953,N_2415);
nor U3793 (N_3793,N_2042,N_2684);
and U3794 (N_3794,N_2429,N_2550);
nand U3795 (N_3795,N_1570,N_1609);
xnor U3796 (N_3796,N_2429,N_1568);
nor U3797 (N_3797,N_1975,N_2807);
or U3798 (N_3798,N_2414,N_2627);
and U3799 (N_3799,N_2602,N_2963);
or U3800 (N_3800,N_1775,N_2780);
or U3801 (N_3801,N_2283,N_2009);
or U3802 (N_3802,N_2819,N_1768);
or U3803 (N_3803,N_1906,N_1736);
and U3804 (N_3804,N_1758,N_2593);
nor U3805 (N_3805,N_1502,N_2068);
nor U3806 (N_3806,N_2251,N_2511);
nand U3807 (N_3807,N_2446,N_2757);
nand U3808 (N_3808,N_2956,N_2198);
nor U3809 (N_3809,N_1919,N_2044);
nor U3810 (N_3810,N_2135,N_1850);
nor U3811 (N_3811,N_1910,N_2497);
nand U3812 (N_3812,N_2221,N_2097);
and U3813 (N_3813,N_2380,N_2721);
nand U3814 (N_3814,N_2450,N_2389);
or U3815 (N_3815,N_1915,N_1838);
nor U3816 (N_3816,N_1908,N_1921);
nand U3817 (N_3817,N_2360,N_2371);
or U3818 (N_3818,N_2791,N_1636);
xor U3819 (N_3819,N_1531,N_1863);
or U3820 (N_3820,N_2581,N_2796);
and U3821 (N_3821,N_2611,N_1520);
nand U3822 (N_3822,N_1626,N_1948);
or U3823 (N_3823,N_2025,N_1853);
or U3824 (N_3824,N_1926,N_2675);
or U3825 (N_3825,N_2780,N_2282);
or U3826 (N_3826,N_1809,N_1769);
and U3827 (N_3827,N_1586,N_2518);
or U3828 (N_3828,N_2046,N_2162);
nand U3829 (N_3829,N_2902,N_2523);
and U3830 (N_3830,N_1732,N_2311);
nor U3831 (N_3831,N_2634,N_1892);
nor U3832 (N_3832,N_2686,N_1683);
nor U3833 (N_3833,N_2856,N_1628);
nand U3834 (N_3834,N_1920,N_1885);
nor U3835 (N_3835,N_2866,N_2507);
or U3836 (N_3836,N_1959,N_2575);
or U3837 (N_3837,N_2511,N_1824);
and U3838 (N_3838,N_2436,N_1853);
and U3839 (N_3839,N_2177,N_2113);
and U3840 (N_3840,N_2936,N_2396);
nand U3841 (N_3841,N_2174,N_2368);
nor U3842 (N_3842,N_2308,N_2546);
or U3843 (N_3843,N_2564,N_2031);
nand U3844 (N_3844,N_1920,N_2544);
and U3845 (N_3845,N_2970,N_2447);
and U3846 (N_3846,N_2967,N_2074);
nor U3847 (N_3847,N_2903,N_2996);
nor U3848 (N_3848,N_2287,N_2195);
or U3849 (N_3849,N_2876,N_2410);
or U3850 (N_3850,N_1749,N_1526);
nor U3851 (N_3851,N_2077,N_1646);
and U3852 (N_3852,N_2921,N_2910);
or U3853 (N_3853,N_2203,N_2673);
nor U3854 (N_3854,N_2218,N_2863);
or U3855 (N_3855,N_2992,N_1802);
and U3856 (N_3856,N_2513,N_2125);
or U3857 (N_3857,N_2037,N_2086);
or U3858 (N_3858,N_2036,N_1972);
and U3859 (N_3859,N_1512,N_2473);
and U3860 (N_3860,N_2402,N_1543);
or U3861 (N_3861,N_2667,N_2211);
nor U3862 (N_3862,N_2232,N_2931);
nor U3863 (N_3863,N_2211,N_1730);
xor U3864 (N_3864,N_2200,N_2124);
nand U3865 (N_3865,N_2065,N_2448);
nor U3866 (N_3866,N_2788,N_2424);
or U3867 (N_3867,N_2102,N_1715);
nor U3868 (N_3868,N_2690,N_1789);
nand U3869 (N_3869,N_2171,N_2028);
and U3870 (N_3870,N_2482,N_2490);
and U3871 (N_3871,N_2099,N_2419);
nor U3872 (N_3872,N_2367,N_2986);
and U3873 (N_3873,N_2637,N_2538);
nand U3874 (N_3874,N_2202,N_2473);
nand U3875 (N_3875,N_2687,N_2076);
nor U3876 (N_3876,N_2946,N_2910);
nand U3877 (N_3877,N_2022,N_2635);
nor U3878 (N_3878,N_2615,N_2499);
nand U3879 (N_3879,N_2331,N_1877);
nand U3880 (N_3880,N_2275,N_2003);
nor U3881 (N_3881,N_2121,N_1620);
nand U3882 (N_3882,N_2282,N_2506);
nor U3883 (N_3883,N_2720,N_2311);
or U3884 (N_3884,N_2844,N_1618);
nor U3885 (N_3885,N_2180,N_2011);
and U3886 (N_3886,N_2976,N_2216);
nand U3887 (N_3887,N_1662,N_2440);
or U3888 (N_3888,N_1774,N_1865);
or U3889 (N_3889,N_2533,N_2670);
and U3890 (N_3890,N_2063,N_2775);
nand U3891 (N_3891,N_2282,N_1690);
or U3892 (N_3892,N_2068,N_1659);
and U3893 (N_3893,N_2327,N_2587);
or U3894 (N_3894,N_1600,N_1820);
or U3895 (N_3895,N_1740,N_1933);
nor U3896 (N_3896,N_2955,N_2174);
nand U3897 (N_3897,N_2546,N_1904);
nand U3898 (N_3898,N_2925,N_1548);
nand U3899 (N_3899,N_2676,N_1503);
nand U3900 (N_3900,N_1818,N_2454);
or U3901 (N_3901,N_2176,N_2556);
and U3902 (N_3902,N_1934,N_2369);
or U3903 (N_3903,N_1522,N_2136);
nor U3904 (N_3904,N_2449,N_2688);
nor U3905 (N_3905,N_2121,N_2397);
and U3906 (N_3906,N_2285,N_2157);
nand U3907 (N_3907,N_2487,N_1804);
nor U3908 (N_3908,N_1770,N_1768);
and U3909 (N_3909,N_2354,N_1592);
and U3910 (N_3910,N_1769,N_2331);
nand U3911 (N_3911,N_2479,N_2363);
nor U3912 (N_3912,N_2675,N_1539);
and U3913 (N_3913,N_2462,N_2560);
nor U3914 (N_3914,N_2828,N_2258);
nor U3915 (N_3915,N_2337,N_2747);
nand U3916 (N_3916,N_2913,N_1953);
or U3917 (N_3917,N_2087,N_1852);
and U3918 (N_3918,N_1772,N_1987);
nand U3919 (N_3919,N_2527,N_2549);
and U3920 (N_3920,N_2393,N_1628);
and U3921 (N_3921,N_2610,N_2285);
nand U3922 (N_3922,N_1621,N_2879);
nand U3923 (N_3923,N_1997,N_2826);
nor U3924 (N_3924,N_1672,N_1628);
xnor U3925 (N_3925,N_2891,N_2562);
or U3926 (N_3926,N_2527,N_2691);
nand U3927 (N_3927,N_2616,N_2239);
nand U3928 (N_3928,N_2802,N_2472);
or U3929 (N_3929,N_2608,N_2980);
or U3930 (N_3930,N_2219,N_2949);
and U3931 (N_3931,N_2890,N_2716);
nand U3932 (N_3932,N_2485,N_1973);
nor U3933 (N_3933,N_2371,N_2713);
nand U3934 (N_3934,N_2348,N_2748);
and U3935 (N_3935,N_1831,N_1753);
nand U3936 (N_3936,N_1550,N_2585);
or U3937 (N_3937,N_2279,N_2506);
and U3938 (N_3938,N_1767,N_2720);
nand U3939 (N_3939,N_1910,N_2792);
or U3940 (N_3940,N_1642,N_1538);
nand U3941 (N_3941,N_1771,N_2127);
nand U3942 (N_3942,N_1716,N_1993);
or U3943 (N_3943,N_2894,N_1997);
nand U3944 (N_3944,N_2293,N_1847);
nand U3945 (N_3945,N_1784,N_1668);
and U3946 (N_3946,N_2777,N_1583);
nor U3947 (N_3947,N_2908,N_1725);
and U3948 (N_3948,N_1617,N_2374);
nand U3949 (N_3949,N_2672,N_1878);
or U3950 (N_3950,N_2213,N_1850);
or U3951 (N_3951,N_2799,N_2394);
or U3952 (N_3952,N_1914,N_2209);
nor U3953 (N_3953,N_2161,N_2031);
nor U3954 (N_3954,N_2311,N_1903);
nor U3955 (N_3955,N_1808,N_2945);
and U3956 (N_3956,N_2982,N_2235);
or U3957 (N_3957,N_1982,N_1930);
nand U3958 (N_3958,N_2325,N_2202);
or U3959 (N_3959,N_1975,N_2759);
nand U3960 (N_3960,N_1966,N_2905);
and U3961 (N_3961,N_2134,N_2991);
nand U3962 (N_3962,N_2188,N_2485);
nand U3963 (N_3963,N_2452,N_2753);
or U3964 (N_3964,N_2893,N_2080);
and U3965 (N_3965,N_1726,N_2631);
nand U3966 (N_3966,N_2935,N_2559);
or U3967 (N_3967,N_1880,N_2715);
xor U3968 (N_3968,N_2388,N_1915);
nor U3969 (N_3969,N_2688,N_2762);
and U3970 (N_3970,N_2123,N_2503);
or U3971 (N_3971,N_1631,N_2855);
and U3972 (N_3972,N_1803,N_2203);
nor U3973 (N_3973,N_1897,N_1751);
or U3974 (N_3974,N_1719,N_2521);
and U3975 (N_3975,N_2972,N_2343);
and U3976 (N_3976,N_2153,N_2873);
nand U3977 (N_3977,N_1834,N_2105);
nand U3978 (N_3978,N_2311,N_1714);
and U3979 (N_3979,N_1837,N_2617);
nand U3980 (N_3980,N_2559,N_2550);
or U3981 (N_3981,N_1610,N_2345);
nor U3982 (N_3982,N_1786,N_2208);
or U3983 (N_3983,N_1715,N_2558);
and U3984 (N_3984,N_2058,N_1647);
or U3985 (N_3985,N_1684,N_1548);
or U3986 (N_3986,N_2142,N_2902);
nand U3987 (N_3987,N_1974,N_2319);
and U3988 (N_3988,N_1677,N_1606);
nor U3989 (N_3989,N_1842,N_2516);
nand U3990 (N_3990,N_1817,N_1987);
nand U3991 (N_3991,N_2090,N_2627);
and U3992 (N_3992,N_1854,N_1671);
or U3993 (N_3993,N_1568,N_2690);
nand U3994 (N_3994,N_2292,N_1685);
nor U3995 (N_3995,N_2396,N_2524);
or U3996 (N_3996,N_1595,N_1540);
and U3997 (N_3997,N_2268,N_2841);
nor U3998 (N_3998,N_2946,N_1825);
and U3999 (N_3999,N_2649,N_2701);
nand U4000 (N_4000,N_2532,N_2330);
or U4001 (N_4001,N_2818,N_1756);
or U4002 (N_4002,N_2367,N_2903);
or U4003 (N_4003,N_2671,N_2352);
nor U4004 (N_4004,N_2148,N_1674);
nor U4005 (N_4005,N_1857,N_2923);
nand U4006 (N_4006,N_2102,N_2830);
nor U4007 (N_4007,N_2721,N_2868);
or U4008 (N_4008,N_2652,N_2889);
nor U4009 (N_4009,N_2235,N_1525);
nor U4010 (N_4010,N_2611,N_2556);
nand U4011 (N_4011,N_2492,N_1844);
and U4012 (N_4012,N_2858,N_2170);
nand U4013 (N_4013,N_2390,N_2288);
or U4014 (N_4014,N_1620,N_2487);
and U4015 (N_4015,N_2125,N_2866);
nand U4016 (N_4016,N_2302,N_2164);
or U4017 (N_4017,N_1674,N_2532);
nor U4018 (N_4018,N_2985,N_2924);
nor U4019 (N_4019,N_2475,N_2381);
nor U4020 (N_4020,N_2335,N_2685);
nand U4021 (N_4021,N_2687,N_2662);
nor U4022 (N_4022,N_2248,N_2060);
nand U4023 (N_4023,N_2430,N_1875);
nor U4024 (N_4024,N_1633,N_2690);
and U4025 (N_4025,N_2871,N_1577);
and U4026 (N_4026,N_2710,N_1611);
nor U4027 (N_4027,N_2620,N_1569);
nor U4028 (N_4028,N_2682,N_2834);
and U4029 (N_4029,N_1662,N_2590);
and U4030 (N_4030,N_2706,N_1952);
nor U4031 (N_4031,N_1876,N_2505);
or U4032 (N_4032,N_1534,N_2670);
nor U4033 (N_4033,N_2108,N_1616);
nor U4034 (N_4034,N_2175,N_2900);
nor U4035 (N_4035,N_1922,N_1661);
nor U4036 (N_4036,N_1583,N_2478);
nor U4037 (N_4037,N_2693,N_2724);
nand U4038 (N_4038,N_2699,N_2644);
and U4039 (N_4039,N_1939,N_1980);
nand U4040 (N_4040,N_1802,N_2631);
or U4041 (N_4041,N_2187,N_2455);
and U4042 (N_4042,N_2684,N_2675);
or U4043 (N_4043,N_2009,N_2941);
nor U4044 (N_4044,N_2852,N_2128);
nand U4045 (N_4045,N_2073,N_2632);
nor U4046 (N_4046,N_1871,N_2493);
and U4047 (N_4047,N_2473,N_2094);
and U4048 (N_4048,N_2075,N_1502);
nor U4049 (N_4049,N_2344,N_1542);
or U4050 (N_4050,N_2883,N_2961);
and U4051 (N_4051,N_2637,N_2464);
or U4052 (N_4052,N_2841,N_2941);
and U4053 (N_4053,N_2620,N_2464);
nand U4054 (N_4054,N_2246,N_2760);
nand U4055 (N_4055,N_1599,N_2901);
or U4056 (N_4056,N_2435,N_2293);
nor U4057 (N_4057,N_2956,N_2180);
nor U4058 (N_4058,N_2603,N_2311);
nor U4059 (N_4059,N_1586,N_1739);
nor U4060 (N_4060,N_2335,N_2126);
nand U4061 (N_4061,N_2167,N_1718);
and U4062 (N_4062,N_2433,N_2532);
nor U4063 (N_4063,N_2851,N_1963);
and U4064 (N_4064,N_2954,N_2782);
or U4065 (N_4065,N_2360,N_2163);
and U4066 (N_4066,N_1785,N_2821);
xor U4067 (N_4067,N_1875,N_2582);
nor U4068 (N_4068,N_1986,N_2111);
nand U4069 (N_4069,N_1913,N_1765);
nand U4070 (N_4070,N_2954,N_1988);
and U4071 (N_4071,N_1659,N_2007);
and U4072 (N_4072,N_2436,N_1554);
nor U4073 (N_4073,N_1654,N_2224);
and U4074 (N_4074,N_2693,N_1550);
nand U4075 (N_4075,N_1612,N_1552);
or U4076 (N_4076,N_1750,N_2573);
and U4077 (N_4077,N_2708,N_2758);
and U4078 (N_4078,N_2835,N_1812);
or U4079 (N_4079,N_2974,N_1515);
and U4080 (N_4080,N_2256,N_2740);
nand U4081 (N_4081,N_1711,N_2245);
nor U4082 (N_4082,N_2741,N_2563);
nor U4083 (N_4083,N_2700,N_2443);
nand U4084 (N_4084,N_1516,N_2976);
nor U4085 (N_4085,N_1590,N_2947);
nor U4086 (N_4086,N_1759,N_2357);
or U4087 (N_4087,N_2787,N_1921);
nor U4088 (N_4088,N_2054,N_1895);
nand U4089 (N_4089,N_1942,N_1682);
or U4090 (N_4090,N_1642,N_2826);
nor U4091 (N_4091,N_2055,N_1805);
or U4092 (N_4092,N_2424,N_2681);
and U4093 (N_4093,N_2875,N_2515);
or U4094 (N_4094,N_1989,N_2397);
or U4095 (N_4095,N_2678,N_2971);
and U4096 (N_4096,N_2438,N_2894);
nand U4097 (N_4097,N_2582,N_2374);
nand U4098 (N_4098,N_1714,N_2630);
and U4099 (N_4099,N_1882,N_1726);
nor U4100 (N_4100,N_2958,N_2029);
or U4101 (N_4101,N_1962,N_2557);
and U4102 (N_4102,N_1827,N_2598);
and U4103 (N_4103,N_2986,N_2338);
or U4104 (N_4104,N_2572,N_2557);
nor U4105 (N_4105,N_1946,N_1878);
nand U4106 (N_4106,N_2068,N_2604);
and U4107 (N_4107,N_2994,N_2495);
nor U4108 (N_4108,N_1874,N_2340);
nand U4109 (N_4109,N_1751,N_2482);
and U4110 (N_4110,N_2958,N_1582);
nand U4111 (N_4111,N_2463,N_1538);
or U4112 (N_4112,N_1812,N_1515);
and U4113 (N_4113,N_2393,N_1663);
or U4114 (N_4114,N_2148,N_2409);
nand U4115 (N_4115,N_1646,N_2069);
nor U4116 (N_4116,N_2637,N_2049);
and U4117 (N_4117,N_1580,N_2026);
and U4118 (N_4118,N_2343,N_2845);
nor U4119 (N_4119,N_2478,N_1830);
and U4120 (N_4120,N_2916,N_2139);
nand U4121 (N_4121,N_1860,N_2131);
and U4122 (N_4122,N_2093,N_1972);
nand U4123 (N_4123,N_2725,N_2017);
or U4124 (N_4124,N_2620,N_1809);
or U4125 (N_4125,N_1598,N_2079);
and U4126 (N_4126,N_2067,N_2606);
and U4127 (N_4127,N_2775,N_2824);
or U4128 (N_4128,N_2857,N_2954);
nor U4129 (N_4129,N_2449,N_2017);
nor U4130 (N_4130,N_1800,N_1786);
nand U4131 (N_4131,N_2973,N_2929);
or U4132 (N_4132,N_1964,N_2975);
nand U4133 (N_4133,N_2786,N_2229);
and U4134 (N_4134,N_2197,N_2676);
or U4135 (N_4135,N_2450,N_2177);
and U4136 (N_4136,N_2472,N_2018);
and U4137 (N_4137,N_2527,N_2847);
nand U4138 (N_4138,N_2877,N_1981);
nor U4139 (N_4139,N_2772,N_2814);
nand U4140 (N_4140,N_1956,N_2754);
or U4141 (N_4141,N_1730,N_1704);
or U4142 (N_4142,N_2471,N_1820);
nor U4143 (N_4143,N_2131,N_2726);
and U4144 (N_4144,N_2960,N_1969);
and U4145 (N_4145,N_1793,N_2137);
or U4146 (N_4146,N_2562,N_1629);
nor U4147 (N_4147,N_2261,N_2860);
or U4148 (N_4148,N_2661,N_1686);
and U4149 (N_4149,N_2614,N_1970);
nand U4150 (N_4150,N_2658,N_2160);
and U4151 (N_4151,N_2799,N_1933);
and U4152 (N_4152,N_1599,N_1619);
nor U4153 (N_4153,N_1779,N_2870);
nor U4154 (N_4154,N_2415,N_2500);
and U4155 (N_4155,N_1912,N_1634);
nand U4156 (N_4156,N_2250,N_2147);
and U4157 (N_4157,N_2948,N_1633);
or U4158 (N_4158,N_2285,N_1939);
nor U4159 (N_4159,N_2595,N_2990);
or U4160 (N_4160,N_2938,N_2832);
or U4161 (N_4161,N_2103,N_2909);
nand U4162 (N_4162,N_2804,N_2755);
and U4163 (N_4163,N_2873,N_2679);
and U4164 (N_4164,N_2086,N_1569);
nor U4165 (N_4165,N_2331,N_2248);
nor U4166 (N_4166,N_2199,N_2266);
or U4167 (N_4167,N_2266,N_1816);
and U4168 (N_4168,N_2331,N_2049);
or U4169 (N_4169,N_2215,N_2627);
nor U4170 (N_4170,N_1969,N_1813);
nor U4171 (N_4171,N_2439,N_1747);
and U4172 (N_4172,N_2997,N_2585);
and U4173 (N_4173,N_2451,N_2496);
nor U4174 (N_4174,N_1503,N_2358);
nor U4175 (N_4175,N_1732,N_1803);
and U4176 (N_4176,N_2360,N_1919);
and U4177 (N_4177,N_2392,N_1648);
or U4178 (N_4178,N_1641,N_2751);
or U4179 (N_4179,N_1716,N_2137);
nor U4180 (N_4180,N_2940,N_2290);
and U4181 (N_4181,N_2775,N_2294);
nor U4182 (N_4182,N_1537,N_1757);
or U4183 (N_4183,N_2650,N_2822);
or U4184 (N_4184,N_2653,N_2501);
and U4185 (N_4185,N_2468,N_1993);
nand U4186 (N_4186,N_2623,N_2953);
or U4187 (N_4187,N_1615,N_1706);
nor U4188 (N_4188,N_2789,N_2003);
nor U4189 (N_4189,N_2965,N_2297);
or U4190 (N_4190,N_2429,N_2455);
nor U4191 (N_4191,N_1934,N_1849);
and U4192 (N_4192,N_1803,N_2968);
and U4193 (N_4193,N_2810,N_2158);
nand U4194 (N_4194,N_1847,N_2459);
nor U4195 (N_4195,N_1699,N_1959);
nand U4196 (N_4196,N_1517,N_1946);
nand U4197 (N_4197,N_2204,N_2284);
nor U4198 (N_4198,N_2930,N_2537);
nor U4199 (N_4199,N_1898,N_2343);
nor U4200 (N_4200,N_2451,N_1720);
nor U4201 (N_4201,N_1536,N_1608);
nand U4202 (N_4202,N_2442,N_2016);
nand U4203 (N_4203,N_2699,N_1543);
and U4204 (N_4204,N_1785,N_2555);
nor U4205 (N_4205,N_2635,N_1601);
and U4206 (N_4206,N_2666,N_2651);
nor U4207 (N_4207,N_2426,N_2431);
nand U4208 (N_4208,N_1929,N_2958);
or U4209 (N_4209,N_1988,N_2948);
or U4210 (N_4210,N_1716,N_1889);
nor U4211 (N_4211,N_1653,N_2797);
and U4212 (N_4212,N_2739,N_1820);
nor U4213 (N_4213,N_1598,N_1558);
and U4214 (N_4214,N_2531,N_2951);
nand U4215 (N_4215,N_2675,N_2284);
and U4216 (N_4216,N_1687,N_2403);
nor U4217 (N_4217,N_2247,N_2387);
and U4218 (N_4218,N_2480,N_1973);
and U4219 (N_4219,N_1858,N_2221);
or U4220 (N_4220,N_2064,N_1970);
and U4221 (N_4221,N_2285,N_1749);
or U4222 (N_4222,N_2486,N_2644);
nor U4223 (N_4223,N_2473,N_2006);
and U4224 (N_4224,N_2193,N_2656);
or U4225 (N_4225,N_1987,N_2532);
nor U4226 (N_4226,N_2900,N_2308);
nand U4227 (N_4227,N_1841,N_2768);
nand U4228 (N_4228,N_2100,N_2956);
and U4229 (N_4229,N_2486,N_2214);
nor U4230 (N_4230,N_2866,N_1995);
or U4231 (N_4231,N_2996,N_2311);
nand U4232 (N_4232,N_2300,N_2457);
nor U4233 (N_4233,N_1577,N_2987);
and U4234 (N_4234,N_2127,N_2308);
and U4235 (N_4235,N_2125,N_2337);
or U4236 (N_4236,N_2712,N_1934);
nor U4237 (N_4237,N_2757,N_2169);
and U4238 (N_4238,N_2076,N_1748);
and U4239 (N_4239,N_1863,N_2526);
and U4240 (N_4240,N_2089,N_2731);
and U4241 (N_4241,N_2912,N_2613);
or U4242 (N_4242,N_2829,N_2762);
nand U4243 (N_4243,N_2174,N_2334);
and U4244 (N_4244,N_1557,N_2762);
or U4245 (N_4245,N_2666,N_1842);
or U4246 (N_4246,N_1538,N_2058);
or U4247 (N_4247,N_2195,N_1756);
or U4248 (N_4248,N_2143,N_1565);
nand U4249 (N_4249,N_2327,N_2841);
or U4250 (N_4250,N_1914,N_2039);
nand U4251 (N_4251,N_2039,N_1614);
nand U4252 (N_4252,N_2114,N_1697);
nand U4253 (N_4253,N_2320,N_1545);
nand U4254 (N_4254,N_2501,N_2385);
nor U4255 (N_4255,N_1811,N_2188);
and U4256 (N_4256,N_1547,N_2756);
and U4257 (N_4257,N_2044,N_2138);
or U4258 (N_4258,N_1969,N_1721);
and U4259 (N_4259,N_2324,N_2774);
and U4260 (N_4260,N_2998,N_2944);
nor U4261 (N_4261,N_2212,N_2580);
or U4262 (N_4262,N_2028,N_2644);
nand U4263 (N_4263,N_1937,N_2953);
or U4264 (N_4264,N_2181,N_2646);
and U4265 (N_4265,N_2936,N_2358);
and U4266 (N_4266,N_1910,N_2514);
nand U4267 (N_4267,N_2986,N_2083);
nor U4268 (N_4268,N_2460,N_1925);
nand U4269 (N_4269,N_2665,N_2105);
nand U4270 (N_4270,N_2624,N_1907);
or U4271 (N_4271,N_1961,N_2793);
nand U4272 (N_4272,N_1538,N_2739);
nand U4273 (N_4273,N_1764,N_1811);
nand U4274 (N_4274,N_2487,N_2277);
nor U4275 (N_4275,N_2788,N_1724);
xnor U4276 (N_4276,N_2364,N_2334);
or U4277 (N_4277,N_1993,N_2407);
and U4278 (N_4278,N_2904,N_1858);
nor U4279 (N_4279,N_1509,N_1606);
nor U4280 (N_4280,N_2514,N_2434);
and U4281 (N_4281,N_2126,N_2557);
or U4282 (N_4282,N_2721,N_1819);
nor U4283 (N_4283,N_1842,N_2621);
nor U4284 (N_4284,N_2287,N_2813);
or U4285 (N_4285,N_2958,N_1705);
nand U4286 (N_4286,N_1604,N_1549);
and U4287 (N_4287,N_2869,N_2978);
or U4288 (N_4288,N_2383,N_1762);
nand U4289 (N_4289,N_1904,N_1926);
nand U4290 (N_4290,N_2100,N_2880);
nand U4291 (N_4291,N_2821,N_2437);
nand U4292 (N_4292,N_2999,N_2246);
and U4293 (N_4293,N_2643,N_2416);
and U4294 (N_4294,N_2114,N_1648);
or U4295 (N_4295,N_2573,N_2495);
nand U4296 (N_4296,N_2782,N_2308);
nor U4297 (N_4297,N_2178,N_1921);
or U4298 (N_4298,N_2578,N_2140);
nor U4299 (N_4299,N_2003,N_2826);
nor U4300 (N_4300,N_2925,N_1537);
or U4301 (N_4301,N_2175,N_2405);
nand U4302 (N_4302,N_1706,N_2964);
nand U4303 (N_4303,N_1769,N_2420);
nand U4304 (N_4304,N_2421,N_2468);
nor U4305 (N_4305,N_1712,N_2582);
and U4306 (N_4306,N_2451,N_1676);
or U4307 (N_4307,N_1773,N_2339);
and U4308 (N_4308,N_1968,N_2321);
and U4309 (N_4309,N_2479,N_2819);
nor U4310 (N_4310,N_2496,N_2840);
and U4311 (N_4311,N_2852,N_1657);
or U4312 (N_4312,N_2536,N_2449);
nand U4313 (N_4313,N_2125,N_1978);
nand U4314 (N_4314,N_2445,N_1958);
and U4315 (N_4315,N_2967,N_1921);
nor U4316 (N_4316,N_1778,N_2845);
and U4317 (N_4317,N_2259,N_2701);
and U4318 (N_4318,N_2435,N_2563);
and U4319 (N_4319,N_2705,N_2317);
and U4320 (N_4320,N_2714,N_1745);
and U4321 (N_4321,N_2388,N_2212);
and U4322 (N_4322,N_2506,N_2109);
or U4323 (N_4323,N_2180,N_2097);
and U4324 (N_4324,N_2638,N_1818);
xnor U4325 (N_4325,N_2682,N_1618);
nor U4326 (N_4326,N_2911,N_2527);
nand U4327 (N_4327,N_1653,N_2648);
or U4328 (N_4328,N_2101,N_2872);
or U4329 (N_4329,N_2472,N_1882);
nand U4330 (N_4330,N_2534,N_2793);
nor U4331 (N_4331,N_2776,N_1671);
or U4332 (N_4332,N_2398,N_2020);
and U4333 (N_4333,N_2327,N_2833);
nor U4334 (N_4334,N_2981,N_2096);
or U4335 (N_4335,N_1714,N_1667);
nor U4336 (N_4336,N_2750,N_2810);
or U4337 (N_4337,N_2831,N_2226);
nor U4338 (N_4338,N_2897,N_2413);
or U4339 (N_4339,N_1575,N_2895);
nand U4340 (N_4340,N_2180,N_2713);
nand U4341 (N_4341,N_2273,N_2979);
or U4342 (N_4342,N_2154,N_2030);
or U4343 (N_4343,N_2854,N_2232);
nand U4344 (N_4344,N_2726,N_2846);
and U4345 (N_4345,N_2300,N_1945);
or U4346 (N_4346,N_1524,N_2993);
and U4347 (N_4347,N_2317,N_1837);
nand U4348 (N_4348,N_2531,N_2661);
nand U4349 (N_4349,N_2407,N_2749);
and U4350 (N_4350,N_2207,N_2569);
nor U4351 (N_4351,N_2588,N_1519);
nor U4352 (N_4352,N_1768,N_1544);
and U4353 (N_4353,N_2190,N_1856);
or U4354 (N_4354,N_2824,N_2317);
nand U4355 (N_4355,N_2599,N_2120);
and U4356 (N_4356,N_2578,N_2216);
or U4357 (N_4357,N_2887,N_2977);
and U4358 (N_4358,N_1696,N_2203);
and U4359 (N_4359,N_2520,N_2085);
or U4360 (N_4360,N_1649,N_2212);
or U4361 (N_4361,N_1914,N_2717);
nand U4362 (N_4362,N_1560,N_2458);
and U4363 (N_4363,N_2106,N_2885);
or U4364 (N_4364,N_1808,N_1966);
nor U4365 (N_4365,N_1924,N_1547);
and U4366 (N_4366,N_2115,N_2182);
nor U4367 (N_4367,N_1733,N_1932);
or U4368 (N_4368,N_2624,N_1554);
nand U4369 (N_4369,N_1939,N_2719);
or U4370 (N_4370,N_1653,N_2198);
and U4371 (N_4371,N_2570,N_2685);
nand U4372 (N_4372,N_2294,N_2314);
and U4373 (N_4373,N_1850,N_1523);
and U4374 (N_4374,N_2155,N_2660);
and U4375 (N_4375,N_2607,N_2109);
nor U4376 (N_4376,N_1912,N_2986);
nor U4377 (N_4377,N_2577,N_2905);
nor U4378 (N_4378,N_2791,N_2786);
and U4379 (N_4379,N_2196,N_2324);
nor U4380 (N_4380,N_1711,N_2036);
nor U4381 (N_4381,N_2933,N_2567);
or U4382 (N_4382,N_2946,N_1589);
nor U4383 (N_4383,N_2727,N_2068);
or U4384 (N_4384,N_1785,N_2419);
nand U4385 (N_4385,N_2669,N_2169);
nand U4386 (N_4386,N_2474,N_2939);
nor U4387 (N_4387,N_1842,N_1715);
nor U4388 (N_4388,N_2453,N_2580);
nand U4389 (N_4389,N_1997,N_1829);
or U4390 (N_4390,N_1896,N_2282);
nor U4391 (N_4391,N_2853,N_2141);
nand U4392 (N_4392,N_1909,N_1974);
and U4393 (N_4393,N_1548,N_1617);
nor U4394 (N_4394,N_2751,N_1695);
nor U4395 (N_4395,N_2320,N_1521);
nor U4396 (N_4396,N_1769,N_1839);
and U4397 (N_4397,N_2617,N_1653);
and U4398 (N_4398,N_1982,N_2719);
nor U4399 (N_4399,N_2758,N_2960);
or U4400 (N_4400,N_2225,N_2198);
or U4401 (N_4401,N_1984,N_1805);
and U4402 (N_4402,N_1973,N_2066);
or U4403 (N_4403,N_2098,N_1985);
nand U4404 (N_4404,N_2836,N_2747);
nand U4405 (N_4405,N_2013,N_1971);
and U4406 (N_4406,N_2299,N_2210);
and U4407 (N_4407,N_2455,N_1966);
nor U4408 (N_4408,N_1794,N_2116);
and U4409 (N_4409,N_2779,N_2419);
nand U4410 (N_4410,N_2750,N_2764);
nand U4411 (N_4411,N_2227,N_1842);
and U4412 (N_4412,N_2580,N_1580);
nand U4413 (N_4413,N_1501,N_1992);
or U4414 (N_4414,N_1670,N_2106);
or U4415 (N_4415,N_2270,N_2201);
nor U4416 (N_4416,N_2486,N_2728);
and U4417 (N_4417,N_2527,N_1897);
nor U4418 (N_4418,N_2130,N_2742);
and U4419 (N_4419,N_1944,N_1517);
and U4420 (N_4420,N_2684,N_2942);
nand U4421 (N_4421,N_2551,N_2411);
or U4422 (N_4422,N_2331,N_2987);
or U4423 (N_4423,N_2381,N_1696);
and U4424 (N_4424,N_2006,N_2345);
nor U4425 (N_4425,N_2817,N_1974);
or U4426 (N_4426,N_1568,N_1685);
nand U4427 (N_4427,N_2875,N_2653);
nand U4428 (N_4428,N_1717,N_2635);
nand U4429 (N_4429,N_2143,N_2405);
nor U4430 (N_4430,N_1860,N_2764);
xor U4431 (N_4431,N_2383,N_2989);
or U4432 (N_4432,N_2613,N_1626);
nor U4433 (N_4433,N_2964,N_2116);
nand U4434 (N_4434,N_1509,N_2273);
and U4435 (N_4435,N_2428,N_1760);
or U4436 (N_4436,N_2470,N_1839);
or U4437 (N_4437,N_1707,N_2293);
nand U4438 (N_4438,N_1596,N_1748);
nor U4439 (N_4439,N_2841,N_2209);
nor U4440 (N_4440,N_2898,N_1616);
and U4441 (N_4441,N_2686,N_1694);
and U4442 (N_4442,N_1690,N_2093);
and U4443 (N_4443,N_2779,N_2584);
and U4444 (N_4444,N_1608,N_2345);
and U4445 (N_4445,N_1851,N_2644);
xor U4446 (N_4446,N_2066,N_2883);
nand U4447 (N_4447,N_2267,N_2429);
or U4448 (N_4448,N_2186,N_2884);
nor U4449 (N_4449,N_2303,N_2993);
and U4450 (N_4450,N_2340,N_1784);
or U4451 (N_4451,N_1721,N_1806);
nand U4452 (N_4452,N_2136,N_1934);
and U4453 (N_4453,N_2095,N_2137);
nor U4454 (N_4454,N_2263,N_2608);
nor U4455 (N_4455,N_2560,N_2535);
nor U4456 (N_4456,N_2432,N_1520);
nor U4457 (N_4457,N_1909,N_2030);
or U4458 (N_4458,N_1934,N_1575);
nand U4459 (N_4459,N_2146,N_2918);
nor U4460 (N_4460,N_2685,N_2520);
and U4461 (N_4461,N_1814,N_2299);
and U4462 (N_4462,N_2676,N_2609);
and U4463 (N_4463,N_2798,N_2903);
nor U4464 (N_4464,N_2507,N_2549);
nor U4465 (N_4465,N_1926,N_2695);
nor U4466 (N_4466,N_2382,N_2873);
or U4467 (N_4467,N_1612,N_2369);
nor U4468 (N_4468,N_2849,N_1933);
and U4469 (N_4469,N_2244,N_1742);
and U4470 (N_4470,N_1994,N_1699);
nor U4471 (N_4471,N_2029,N_1552);
nor U4472 (N_4472,N_1953,N_1521);
and U4473 (N_4473,N_2085,N_2946);
nor U4474 (N_4474,N_2533,N_2078);
or U4475 (N_4475,N_2929,N_2424);
or U4476 (N_4476,N_2915,N_1975);
nor U4477 (N_4477,N_1897,N_2852);
nor U4478 (N_4478,N_2987,N_2060);
nand U4479 (N_4479,N_2504,N_1876);
nor U4480 (N_4480,N_2455,N_2116);
nand U4481 (N_4481,N_1750,N_2362);
nor U4482 (N_4482,N_2983,N_2404);
nand U4483 (N_4483,N_2830,N_1864);
nand U4484 (N_4484,N_2978,N_2540);
and U4485 (N_4485,N_2804,N_2494);
and U4486 (N_4486,N_2578,N_2468);
or U4487 (N_4487,N_1964,N_2759);
or U4488 (N_4488,N_2675,N_1924);
or U4489 (N_4489,N_1931,N_1729);
nor U4490 (N_4490,N_2072,N_2399);
nor U4491 (N_4491,N_2382,N_2425);
or U4492 (N_4492,N_1604,N_2030);
and U4493 (N_4493,N_1783,N_2523);
nand U4494 (N_4494,N_2083,N_1509);
or U4495 (N_4495,N_1506,N_1983);
or U4496 (N_4496,N_2684,N_1706);
nand U4497 (N_4497,N_2595,N_2407);
or U4498 (N_4498,N_2398,N_1809);
nor U4499 (N_4499,N_1586,N_2173);
or U4500 (N_4500,N_4285,N_3443);
or U4501 (N_4501,N_3296,N_3458);
or U4502 (N_4502,N_4154,N_3416);
and U4503 (N_4503,N_4082,N_4200);
nand U4504 (N_4504,N_3011,N_3943);
nor U4505 (N_4505,N_4129,N_4034);
or U4506 (N_4506,N_4273,N_3204);
nand U4507 (N_4507,N_3932,N_4127);
or U4508 (N_4508,N_3609,N_3560);
xnor U4509 (N_4509,N_4225,N_3836);
nand U4510 (N_4510,N_4404,N_3916);
and U4511 (N_4511,N_4165,N_3874);
nor U4512 (N_4512,N_4291,N_4201);
nand U4513 (N_4513,N_3522,N_4118);
or U4514 (N_4514,N_4195,N_3155);
nand U4515 (N_4515,N_3133,N_3840);
and U4516 (N_4516,N_3956,N_4356);
or U4517 (N_4517,N_4022,N_4375);
xnor U4518 (N_4518,N_3175,N_4333);
or U4519 (N_4519,N_4467,N_3909);
or U4520 (N_4520,N_3855,N_3048);
or U4521 (N_4521,N_4015,N_3374);
and U4522 (N_4522,N_4402,N_3156);
and U4523 (N_4523,N_3883,N_3819);
nor U4524 (N_4524,N_3983,N_3553);
nand U4525 (N_4525,N_3832,N_3814);
or U4526 (N_4526,N_4303,N_3165);
and U4527 (N_4527,N_3394,N_4458);
nand U4528 (N_4528,N_3525,N_4236);
nand U4529 (N_4529,N_3232,N_3886);
nor U4530 (N_4530,N_4270,N_4120);
nor U4531 (N_4531,N_3988,N_3263);
and U4532 (N_4532,N_4013,N_4395);
or U4533 (N_4533,N_3278,N_4049);
xor U4534 (N_4534,N_3537,N_3391);
nand U4535 (N_4535,N_4144,N_3171);
nand U4536 (N_4536,N_3892,N_3856);
or U4537 (N_4537,N_3474,N_4256);
and U4538 (N_4538,N_4260,N_3835);
and U4539 (N_4539,N_3024,N_3573);
nand U4540 (N_4540,N_4253,N_4481);
nand U4541 (N_4541,N_3066,N_4194);
and U4542 (N_4542,N_4489,N_4114);
xnor U4543 (N_4543,N_4204,N_4104);
nor U4544 (N_4544,N_4282,N_3585);
nand U4545 (N_4545,N_3216,N_4327);
nor U4546 (N_4546,N_4183,N_3080);
or U4547 (N_4547,N_3332,N_3422);
nand U4548 (N_4548,N_4143,N_4418);
and U4549 (N_4549,N_3392,N_3464);
and U4550 (N_4550,N_4370,N_4242);
or U4551 (N_4551,N_3183,N_4365);
nor U4552 (N_4552,N_4400,N_3690);
nand U4553 (N_4553,N_3272,N_3775);
and U4554 (N_4554,N_3334,N_3100);
or U4555 (N_4555,N_3815,N_3423);
or U4556 (N_4556,N_3357,N_3505);
or U4557 (N_4557,N_3549,N_3297);
or U4558 (N_4558,N_3169,N_4492);
nor U4559 (N_4559,N_3681,N_4245);
nand U4560 (N_4560,N_4284,N_4459);
and U4561 (N_4561,N_3338,N_3099);
nor U4562 (N_4562,N_4463,N_3212);
and U4563 (N_4563,N_4248,N_4440);
or U4564 (N_4564,N_3208,N_3828);
and U4565 (N_4565,N_4086,N_3259);
and U4566 (N_4566,N_3222,N_3527);
and U4567 (N_4567,N_4430,N_3049);
or U4568 (N_4568,N_4336,N_3791);
nand U4569 (N_4569,N_3950,N_4071);
nor U4570 (N_4570,N_3979,N_3999);
or U4571 (N_4571,N_3426,N_4151);
nand U4572 (N_4572,N_3646,N_3345);
nor U4573 (N_4573,N_4385,N_4388);
and U4574 (N_4574,N_3327,N_4098);
nor U4575 (N_4575,N_3403,N_4043);
nor U4576 (N_4576,N_3056,N_3306);
or U4577 (N_4577,N_3853,N_3982);
or U4578 (N_4578,N_3589,N_3055);
or U4579 (N_4579,N_3352,N_3355);
nor U4580 (N_4580,N_3105,N_4277);
or U4581 (N_4581,N_3301,N_3157);
nor U4582 (N_4582,N_4217,N_4229);
or U4583 (N_4583,N_3688,N_3287);
nor U4584 (N_4584,N_4206,N_3533);
and U4585 (N_4585,N_4093,N_3177);
nor U4586 (N_4586,N_3405,N_3419);
or U4587 (N_4587,N_3262,N_3981);
and U4588 (N_4588,N_4132,N_3510);
and U4589 (N_4589,N_3975,N_3907);
and U4590 (N_4590,N_3502,N_3662);
and U4591 (N_4591,N_3253,N_3842);
and U4592 (N_4592,N_3800,N_4171);
or U4593 (N_4593,N_3472,N_3057);
nand U4594 (N_4594,N_3752,N_4239);
and U4595 (N_4595,N_4450,N_4212);
and U4596 (N_4596,N_4462,N_4480);
nor U4597 (N_4597,N_4329,N_4044);
and U4598 (N_4598,N_3670,N_4424);
and U4599 (N_4599,N_4369,N_3843);
or U4600 (N_4600,N_4042,N_3616);
nand U4601 (N_4601,N_3768,N_4081);
and U4602 (N_4602,N_3424,N_3729);
and U4603 (N_4603,N_3315,N_4235);
and U4604 (N_4604,N_3656,N_3031);
nor U4605 (N_4605,N_3487,N_3314);
and U4606 (N_4606,N_4393,N_3132);
nand U4607 (N_4607,N_4172,N_4208);
or U4608 (N_4608,N_3453,N_3028);
and U4609 (N_4609,N_4167,N_3034);
nor U4610 (N_4610,N_4448,N_3205);
nand U4611 (N_4611,N_3337,N_3331);
and U4612 (N_4612,N_4032,N_4255);
nand U4613 (N_4613,N_3279,N_3083);
nor U4614 (N_4614,N_3620,N_3737);
nor U4615 (N_4615,N_3808,N_3861);
or U4616 (N_4616,N_4061,N_3063);
nand U4617 (N_4617,N_3087,N_4301);
nor U4618 (N_4618,N_3606,N_3241);
nand U4619 (N_4619,N_3528,N_3753);
or U4620 (N_4620,N_3077,N_3199);
and U4621 (N_4621,N_3123,N_3020);
nand U4622 (N_4622,N_3784,N_4487);
and U4623 (N_4623,N_3265,N_3353);
or U4624 (N_4624,N_3696,N_3811);
or U4625 (N_4625,N_3967,N_3161);
and U4626 (N_4626,N_3546,N_3460);
nand U4627 (N_4627,N_3079,N_4115);
nor U4628 (N_4628,N_4296,N_4037);
and U4629 (N_4629,N_3266,N_3891);
or U4630 (N_4630,N_3703,N_3863);
nand U4631 (N_4631,N_3035,N_3303);
and U4632 (N_4632,N_4415,N_3381);
nor U4633 (N_4633,N_3299,N_3320);
and U4634 (N_4634,N_3640,N_4221);
and U4635 (N_4635,N_3793,N_3897);
or U4636 (N_4636,N_4444,N_3516);
and U4637 (N_4637,N_3629,N_4233);
nor U4638 (N_4638,N_3110,N_3172);
nand U4639 (N_4639,N_4435,N_3860);
and U4640 (N_4640,N_3326,N_3007);
or U4641 (N_4641,N_3715,N_3408);
or U4642 (N_4642,N_3582,N_3642);
nand U4643 (N_4643,N_4371,N_3657);
nor U4644 (N_4644,N_3548,N_3968);
and U4645 (N_4645,N_3624,N_4353);
or U4646 (N_4646,N_3196,N_3709);
or U4647 (N_4647,N_3672,N_4361);
nand U4648 (N_4648,N_3052,N_3722);
nand U4649 (N_4649,N_3558,N_3978);
and U4650 (N_4650,N_3429,N_3275);
and U4651 (N_4651,N_4470,N_4137);
nand U4652 (N_4652,N_3188,N_3952);
nor U4653 (N_4653,N_4139,N_3494);
nand U4654 (N_4654,N_4320,N_4328);
nand U4655 (N_4655,N_4192,N_3865);
or U4656 (N_4656,N_3653,N_3484);
and U4657 (N_4657,N_3803,N_3668);
nand U4658 (N_4658,N_3714,N_4142);
nor U4659 (N_4659,N_3910,N_4173);
or U4660 (N_4660,N_4457,N_4306);
and U4661 (N_4661,N_3894,N_3748);
nand U4662 (N_4662,N_4307,N_3389);
or U4663 (N_4663,N_3089,N_3902);
and U4664 (N_4664,N_3849,N_3112);
nor U4665 (N_4665,N_3936,N_3039);
nand U4666 (N_4666,N_3141,N_3837);
and U4667 (N_4667,N_3746,N_3185);
nor U4668 (N_4668,N_4378,N_4461);
or U4669 (N_4669,N_4437,N_4138);
nor U4670 (N_4670,N_3248,N_4247);
nand U4671 (N_4671,N_3693,N_3711);
nand U4672 (N_4672,N_3673,N_3858);
or U4673 (N_4673,N_3520,N_3747);
nand U4674 (N_4674,N_4368,N_3705);
nor U4675 (N_4675,N_3015,N_3201);
nand U4676 (N_4676,N_3158,N_3261);
nand U4677 (N_4677,N_3434,N_3237);
and U4678 (N_4678,N_3953,N_3147);
nand U4679 (N_4679,N_4429,N_4309);
and U4680 (N_4680,N_3862,N_4485);
nand U4681 (N_4681,N_3876,N_4259);
nand U4682 (N_4682,N_3300,N_3985);
and U4683 (N_4683,N_3859,N_4454);
nand U4684 (N_4684,N_4413,N_3984);
or U4685 (N_4685,N_3065,N_4325);
nand U4686 (N_4686,N_3554,N_3682);
nand U4687 (N_4687,N_3749,N_3578);
or U4688 (N_4688,N_3648,N_3519);
nand U4689 (N_4689,N_3704,N_4261);
and U4690 (N_4690,N_4055,N_3721);
nor U4691 (N_4691,N_3428,N_3281);
nand U4692 (N_4692,N_4384,N_3053);
nor U4693 (N_4693,N_4460,N_4408);
or U4694 (N_4694,N_4023,N_3799);
nor U4695 (N_4695,N_3193,N_3166);
nor U4696 (N_4696,N_3625,N_3944);
and U4697 (N_4697,N_3603,N_4308);
nor U4698 (N_4698,N_3634,N_3942);
or U4699 (N_4699,N_3732,N_4092);
nor U4700 (N_4700,N_4477,N_3102);
and U4701 (N_4701,N_4178,N_3313);
and U4702 (N_4702,N_3929,N_3698);
nor U4703 (N_4703,N_3765,N_3900);
xnor U4704 (N_4704,N_4390,N_3276);
nor U4705 (N_4705,N_4283,N_3664);
or U4706 (N_4706,N_3068,N_3257);
nand U4707 (N_4707,N_3202,N_4106);
and U4708 (N_4708,N_3798,N_4153);
nor U4709 (N_4709,N_3750,N_3319);
nor U4710 (N_4710,N_3927,N_3540);
nand U4711 (N_4711,N_3187,N_3933);
or U4712 (N_4712,N_3008,N_4258);
nand U4713 (N_4713,N_3877,N_3127);
nor U4714 (N_4714,N_3960,N_3884);
or U4715 (N_4715,N_3866,N_3779);
nand U4716 (N_4716,N_3150,N_4059);
nand U4717 (N_4717,N_3587,N_4315);
nor U4718 (N_4718,N_3027,N_4088);
or U4719 (N_4719,N_3255,N_3564);
or U4720 (N_4720,N_3251,N_4170);
nor U4721 (N_4721,N_4311,N_3783);
nand U4722 (N_4722,N_3919,N_3115);
nand U4723 (N_4723,N_3777,N_3120);
and U4724 (N_4724,N_4210,N_3621);
nand U4725 (N_4725,N_4338,N_3989);
nand U4726 (N_4726,N_4422,N_3545);
or U4727 (N_4727,N_4169,N_3937);
nor U4728 (N_4728,N_3240,N_3782);
nor U4729 (N_4729,N_3179,N_4264);
nor U4730 (N_4730,N_3647,N_3486);
nand U4731 (N_4731,N_3764,N_3277);
nor U4732 (N_4732,N_3140,N_3666);
nand U4733 (N_4733,N_3191,N_4111);
and U4734 (N_4734,N_3758,N_4438);
or U4735 (N_4735,N_3513,N_3043);
nand U4736 (N_4736,N_4441,N_3743);
and U4737 (N_4737,N_3234,N_3440);
nor U4738 (N_4738,N_4380,N_3005);
and U4739 (N_4739,N_4045,N_3563);
nor U4740 (N_4740,N_3605,N_3162);
nor U4741 (N_4741,N_3993,N_3991);
or U4742 (N_4742,N_4004,N_3821);
and U4743 (N_4743,N_4156,N_3214);
nor U4744 (N_4744,N_3718,N_3333);
nand U4745 (N_4745,N_3471,N_3113);
nand U4746 (N_4746,N_3371,N_4240);
and U4747 (N_4747,N_3467,N_4340);
or U4748 (N_4748,N_4050,N_3622);
or U4749 (N_4749,N_3612,N_4318);
nand U4750 (N_4750,N_3741,N_3774);
nor U4751 (N_4751,N_3555,N_3385);
and U4752 (N_4752,N_3360,N_3069);
xnor U4753 (N_4753,N_4381,N_4272);
or U4754 (N_4754,N_4160,N_3760);
nor U4755 (N_4755,N_4068,N_3367);
or U4756 (N_4756,N_4271,N_4374);
and U4757 (N_4757,N_3448,N_3482);
nand U4758 (N_4758,N_3675,N_3192);
or U4759 (N_4759,N_4376,N_4432);
and U4760 (N_4760,N_3496,N_3759);
nor U4761 (N_4761,N_3805,N_3432);
nor U4762 (N_4762,N_3081,N_3042);
and U4763 (N_4763,N_3233,N_3570);
and U4764 (N_4764,N_3086,N_3380);
and U4765 (N_4765,N_4084,N_3059);
nand U4766 (N_4766,N_3700,N_4399);
and U4767 (N_4767,N_3896,N_4300);
or U4768 (N_4768,N_4348,N_3219);
or U4769 (N_4769,N_3845,N_3957);
nor U4770 (N_4770,N_3444,N_4005);
nor U4771 (N_4771,N_3073,N_4266);
nand U4772 (N_4772,N_4124,N_3885);
or U4773 (N_4773,N_3996,N_4476);
nand U4774 (N_4774,N_4234,N_3571);
or U4775 (N_4775,N_3071,N_3200);
nand U4776 (N_4776,N_4162,N_4286);
and U4777 (N_4777,N_3365,N_3308);
nand U4778 (N_4778,N_4038,N_3173);
and U4779 (N_4779,N_3637,N_3454);
and U4780 (N_4780,N_3145,N_4145);
or U4781 (N_4781,N_3004,N_3022);
or U4782 (N_4782,N_4067,N_3480);
and U4783 (N_4783,N_3931,N_4449);
or U4784 (N_4784,N_3713,N_3117);
nor U4785 (N_4785,N_3364,N_4113);
nand U4786 (N_4786,N_3131,N_3441);
nand U4787 (N_4787,N_4150,N_4297);
nor U4788 (N_4788,N_3506,N_4222);
or U4789 (N_4789,N_4317,N_4464);
nand U4790 (N_4790,N_4265,N_3271);
and U4791 (N_4791,N_4251,N_3001);
and U4792 (N_4792,N_4499,N_4105);
nor U4793 (N_4793,N_3209,N_3317);
nor U4794 (N_4794,N_4313,N_3321);
nand U4795 (N_4795,N_3706,N_3676);
and U4796 (N_4796,N_4227,N_3854);
or U4797 (N_4797,N_3868,N_3913);
and U4798 (N_4798,N_4349,N_3610);
nor U4799 (N_4799,N_3146,N_3654);
nor U4800 (N_4800,N_3766,N_3139);
nor U4801 (N_4801,N_3725,N_4080);
or U4802 (N_4802,N_3776,N_3207);
nor U4803 (N_4803,N_3189,N_4198);
and U4804 (N_4804,N_4493,N_3598);
or U4805 (N_4805,N_4215,N_3457);
nand U4806 (N_4806,N_4189,N_3125);
nor U4807 (N_4807,N_3658,N_3134);
and U4808 (N_4808,N_4213,N_3745);
nor U4809 (N_4809,N_3959,N_4063);
and U4810 (N_4810,N_3816,N_3070);
or U4811 (N_4811,N_3669,N_3010);
or U4812 (N_4812,N_3905,N_3017);
nand U4813 (N_4813,N_3093,N_4252);
nand U4814 (N_4814,N_4275,N_3149);
or U4815 (N_4815,N_4020,N_3411);
or U4816 (N_4816,N_3002,N_3971);
nand U4817 (N_4817,N_3839,N_3559);
nand U4818 (N_4818,N_4048,N_3243);
and U4819 (N_4819,N_3304,N_3930);
and U4820 (N_4820,N_4214,N_4434);
or U4821 (N_4821,N_3286,N_3674);
nand U4822 (N_4822,N_4382,N_3270);
nand U4823 (N_4823,N_3438,N_3607);
nand U4824 (N_4824,N_3763,N_4030);
nand U4825 (N_4825,N_4394,N_4482);
nor U4826 (N_4826,N_4047,N_3997);
and U4827 (N_4827,N_3879,N_3918);
or U4828 (N_4828,N_3901,N_3249);
nor U4829 (N_4829,N_3801,N_4339);
nand U4830 (N_4830,N_3402,N_3807);
xor U4831 (N_4831,N_3492,N_4119);
nand U4832 (N_4832,N_3493,N_4312);
and U4833 (N_4833,N_4359,N_3386);
nor U4834 (N_4834,N_4290,N_4396);
nor U4835 (N_4835,N_4383,N_3906);
and U4836 (N_4836,N_4330,N_4117);
or U4837 (N_4837,N_3325,N_3641);
and U4838 (N_4838,N_4428,N_4324);
or U4839 (N_4839,N_3632,N_3795);
and U4840 (N_4840,N_4414,N_3142);
and U4841 (N_4841,N_4116,N_3437);
or U4842 (N_4842,N_3462,N_3794);
nand U4843 (N_4843,N_4219,N_3660);
or U4844 (N_4844,N_3498,N_3124);
nand U4845 (N_4845,N_4474,N_3054);
nand U4846 (N_4846,N_3692,N_4326);
or U4847 (N_4847,N_3116,N_3267);
nand U4848 (N_4848,N_3822,N_3871);
nor U4849 (N_4849,N_3994,N_3128);
or U4850 (N_4850,N_3912,N_3524);
nor U4851 (N_4851,N_4427,N_3834);
nand U4852 (N_4852,N_3890,N_3459);
xor U4853 (N_4853,N_3618,N_3590);
or U4854 (N_4854,N_3501,N_3178);
nand U4855 (N_4855,N_4083,N_4392);
nand U4856 (N_4856,N_4070,N_3414);
nor U4857 (N_4857,N_4310,N_3407);
nor U4858 (N_4858,N_3870,N_3818);
or U4859 (N_4859,N_3736,N_3707);
nand U4860 (N_4860,N_4164,N_3898);
and U4861 (N_4861,N_3723,N_3060);
nor U4862 (N_4862,N_3726,N_3136);
xnor U4863 (N_4863,N_3449,N_3580);
or U4864 (N_4864,N_3154,N_4455);
nand U4865 (N_4865,N_3823,N_4405);
and U4866 (N_4866,N_3121,N_4280);
or U4867 (N_4867,N_3223,N_4419);
or U4868 (N_4868,N_3804,N_3290);
nor U4869 (N_4869,N_4094,N_3771);
or U4870 (N_4870,N_3881,N_4026);
nor U4871 (N_4871,N_4299,N_3298);
nand U4872 (N_4872,N_3351,N_3170);
nand U4873 (N_4873,N_3581,N_3029);
and U4874 (N_4874,N_4387,N_3370);
nand U4875 (N_4875,N_3934,N_4146);
nand U4876 (N_4876,N_4095,N_4135);
or U4877 (N_4877,N_3252,N_3097);
and U4878 (N_4878,N_4334,N_3787);
nand U4879 (N_4879,N_3159,N_4193);
nor U4880 (N_4880,N_3288,N_4377);
and U4881 (N_4881,N_4011,N_3095);
nor U4882 (N_4882,N_3577,N_3476);
nand U4883 (N_4883,N_3305,N_3036);
nand U4884 (N_4884,N_4295,N_3965);
and U4885 (N_4885,N_3283,N_4269);
or U4886 (N_4886,N_3312,N_4244);
nand U4887 (N_4887,N_4343,N_3176);
nand U4888 (N_4888,N_3401,N_4168);
nor U4889 (N_4889,N_3733,N_4029);
nand U4890 (N_4890,N_4197,N_3358);
and U4891 (N_4891,N_4465,N_3938);
nand U4892 (N_4892,N_3349,N_4421);
nor U4893 (N_4893,N_4230,N_3311);
nand U4894 (N_4894,N_3523,N_3211);
or U4895 (N_4895,N_4495,N_4278);
nand U4896 (N_4896,N_3652,N_3363);
nor U4897 (N_4897,N_3148,N_3848);
nor U4898 (N_4898,N_3122,N_4466);
or U4899 (N_4899,N_3023,N_3514);
nand U4900 (N_4900,N_4108,N_3686);
nor U4901 (N_4901,N_3377,N_4121);
and U4902 (N_4902,N_3427,N_4177);
nand U4903 (N_4903,N_3037,N_4000);
nor U4904 (N_4904,N_3562,N_3235);
and U4905 (N_4905,N_3517,N_3948);
and U4906 (N_4906,N_3130,N_3250);
nand U4907 (N_4907,N_3220,N_4077);
and U4908 (N_4908,N_4122,N_3796);
or U4909 (N_4909,N_4207,N_4398);
nor U4910 (N_4910,N_3539,N_3995);
xor U4911 (N_4911,N_3406,N_3384);
nor U4912 (N_4912,N_3344,N_3160);
nand U4913 (N_4913,N_4134,N_4347);
and U4914 (N_4914,N_3404,N_3309);
nand U4915 (N_4915,N_3339,N_3786);
nand U4916 (N_4916,N_3468,N_4436);
nor U4917 (N_4917,N_3511,N_3274);
or U4918 (N_4918,N_4141,N_3033);
or U4919 (N_4919,N_3908,N_3850);
and U4920 (N_4920,N_3247,N_4102);
nand U4921 (N_4921,N_4469,N_3683);
nor U4922 (N_4922,N_4451,N_3186);
nand U4923 (N_4923,N_3797,N_4498);
nand U4924 (N_4924,N_3108,N_3551);
xor U4925 (N_4925,N_3119,N_4025);
or U4926 (N_4926,N_3926,N_3827);
nor U4927 (N_4927,N_3593,N_3181);
or U4928 (N_4928,N_3972,N_3829);
and U4929 (N_4929,N_3280,N_3973);
and U4930 (N_4930,N_3844,N_3198);
and U4931 (N_4931,N_3684,N_4079);
nor U4932 (N_4932,N_4069,N_3882);
nand U4933 (N_4933,N_3728,N_3591);
or U4934 (N_4934,N_3710,N_4223);
or U4935 (N_4935,N_4445,N_3639);
nand U4936 (N_4936,N_4496,N_3477);
nor U4937 (N_4937,N_3481,N_3756);
nand U4938 (N_4938,N_4323,N_3268);
or U4939 (N_4939,N_4335,N_3712);
or U4940 (N_4940,N_3221,N_4267);
nor U4941 (N_4941,N_4226,N_3630);
and U4942 (N_4942,N_4497,N_3359);
or U4943 (N_4943,N_3534,N_3966);
and U4944 (N_4944,N_4019,N_3269);
or U4945 (N_4945,N_4345,N_3461);
and U4946 (N_4946,N_3663,N_4231);
and U4947 (N_4947,N_4257,N_3413);
or U4948 (N_4948,N_3810,N_4130);
nor U4949 (N_4949,N_3644,N_3026);
and U4950 (N_4950,N_3659,N_3078);
or U4951 (N_4951,N_4220,N_3767);
nor U4952 (N_4952,N_4012,N_3399);
or U4953 (N_4953,N_3203,N_3792);
nand U4954 (N_4954,N_4243,N_4484);
nor U4955 (N_4955,N_3447,N_3388);
and U4956 (N_4956,N_3163,N_4010);
nor U4957 (N_4957,N_4006,N_3627);
nor U4958 (N_4958,N_3594,N_3601);
nand U4959 (N_4959,N_3708,N_3336);
or U4960 (N_4960,N_3076,N_4288);
nand U4961 (N_4961,N_4040,N_4052);
nand U4962 (N_4962,N_4289,N_4494);
or U4963 (N_4963,N_3439,N_4447);
and U4964 (N_4964,N_4468,N_3701);
nor U4965 (N_4965,N_3425,N_4107);
nor U4966 (N_4966,N_4155,N_4076);
and U4967 (N_4967,N_4411,N_3228);
and U4968 (N_4968,N_3695,N_3769);
nor U4969 (N_4969,N_4147,N_3226);
nand U4970 (N_4970,N_4109,N_3949);
or U4971 (N_4971,N_3103,N_3574);
nand U4972 (N_4972,N_3961,N_3813);
or U4973 (N_4973,N_3045,N_4100);
nand U4974 (N_4974,N_4016,N_3636);
or U4975 (N_4975,N_3258,N_3293);
nand U4976 (N_4976,N_4075,N_3939);
nand U4977 (N_4977,N_3809,N_3397);
and U4978 (N_4978,N_3928,N_3963);
nand U4979 (N_4979,N_3626,N_3899);
or U4980 (N_4980,N_3025,N_4054);
and U4981 (N_4981,N_3922,N_4191);
and U4982 (N_4982,N_3180,N_4174);
nand U4983 (N_4983,N_3526,N_3084);
nand U4984 (N_4984,N_3608,N_3781);
nor U4985 (N_4985,N_4148,N_4416);
or U4986 (N_4986,N_3174,N_3151);
nand U4987 (N_4987,N_3872,N_3244);
or U4988 (N_4988,N_3535,N_3550);
nor U4989 (N_4989,N_4302,N_3378);
or U4990 (N_4990,N_3393,N_3830);
nor U4991 (N_4991,N_4407,N_3041);
and U4992 (N_4992,N_3831,N_3218);
nand U4993 (N_4993,N_3046,N_3980);
and U4994 (N_4994,N_3542,N_3164);
and U4995 (N_4995,N_4003,N_3780);
nor U4996 (N_4996,N_3802,N_3479);
nand U4997 (N_4997,N_3512,N_3770);
or U4998 (N_4998,N_3569,N_3435);
nand U4999 (N_4999,N_3238,N_4331);
nor U5000 (N_5000,N_3082,N_4238);
nand U5001 (N_5001,N_3739,N_3575);
nand U5002 (N_5002,N_4062,N_3806);
or U5003 (N_5003,N_3168,N_3592);
and U5004 (N_5004,N_3679,N_3323);
nand U5005 (N_5005,N_3295,N_4035);
nor U5006 (N_5006,N_3184,N_4166);
nand U5007 (N_5007,N_4366,N_4136);
nand U5008 (N_5008,N_4412,N_4473);
nand U5009 (N_5009,N_4058,N_3597);
nand U5010 (N_5010,N_4483,N_3012);
nand U5011 (N_5011,N_3284,N_3294);
or U5012 (N_5012,N_4332,N_3348);
or U5013 (N_5013,N_3264,N_3072);
and U5014 (N_5014,N_3873,N_4279);
nand U5015 (N_5015,N_4099,N_3356);
xnor U5016 (N_5016,N_3665,N_3310);
or U5017 (N_5017,N_4180,N_3092);
nor U5018 (N_5018,N_4018,N_3455);
nand U5019 (N_5019,N_3469,N_4033);
nor U5020 (N_5020,N_3206,N_4292);
nand U5021 (N_5021,N_4237,N_3547);
and U5022 (N_5022,N_3941,N_4446);
or U5023 (N_5023,N_4294,N_3418);
nor U5024 (N_5024,N_3602,N_3347);
and U5025 (N_5025,N_4149,N_4216);
or U5026 (N_5026,N_4001,N_4479);
or U5027 (N_5027,N_3572,N_4008);
nand U5028 (N_5028,N_3515,N_3047);
nand U5029 (N_5029,N_3478,N_4046);
nor U5030 (N_5030,N_3285,N_3490);
and U5031 (N_5031,N_3445,N_3561);
nand U5032 (N_5032,N_3757,N_3436);
nor U5033 (N_5033,N_3864,N_4028);
nand U5034 (N_5034,N_4490,N_4228);
nor U5035 (N_5035,N_3410,N_3489);
or U5036 (N_5036,N_3667,N_4041);
nor U5037 (N_5037,N_4126,N_4128);
nand U5038 (N_5038,N_3613,N_4262);
nor U5039 (N_5039,N_4187,N_3246);
or U5040 (N_5040,N_4182,N_3631);
or U5041 (N_5041,N_3838,N_3000);
and U5042 (N_5042,N_3346,N_3735);
and U5043 (N_5043,N_3003,N_4097);
nand U5044 (N_5044,N_3504,N_3935);
or U5045 (N_5045,N_4472,N_4249);
nor U5046 (N_5046,N_4158,N_3521);
or U5047 (N_5047,N_4274,N_3111);
nand U5048 (N_5048,N_3372,N_3499);
nor U5049 (N_5049,N_3040,N_3488);
nand U5050 (N_5050,N_3064,N_3431);
or U5051 (N_5051,N_4420,N_3552);
or U5052 (N_5052,N_3109,N_4456);
and U5053 (N_5053,N_3740,N_3878);
and U5054 (N_5054,N_3376,N_3887);
nor U5055 (N_5055,N_4321,N_3847);
nor U5056 (N_5056,N_3213,N_3006);
nand U5057 (N_5057,N_3236,N_4232);
and U5058 (N_5058,N_3051,N_3964);
xor U5059 (N_5059,N_4352,N_3731);
nand U5060 (N_5060,N_3677,N_3584);
xnor U5061 (N_5061,N_3651,N_3421);
nand U5062 (N_5062,N_3307,N_4031);
nand U5063 (N_5063,N_4185,N_4110);
or U5064 (N_5064,N_3595,N_4205);
nand U5065 (N_5065,N_4342,N_3529);
nand U5066 (N_5066,N_3789,N_3417);
nand U5067 (N_5067,N_3826,N_4403);
nor U5068 (N_5068,N_3452,N_4196);
or U5069 (N_5069,N_4159,N_3014);
nor U5070 (N_5070,N_4157,N_3538);
nand U5071 (N_5071,N_3369,N_3224);
and U5072 (N_5072,N_3604,N_4268);
or U5073 (N_5073,N_3229,N_3152);
nor U5074 (N_5074,N_3361,N_3869);
nand U5075 (N_5075,N_3329,N_3450);
or U5076 (N_5076,N_3409,N_3566);
nor U5077 (N_5077,N_3075,N_3106);
nand U5078 (N_5078,N_4066,N_3857);
nor U5079 (N_5079,N_3340,N_3144);
and U5080 (N_5080,N_4057,N_3643);
or U5081 (N_5081,N_3466,N_3727);
nor U5082 (N_5082,N_3330,N_4475);
and U5083 (N_5083,N_4344,N_4009);
or U5084 (N_5084,N_4372,N_3716);
or U5085 (N_5085,N_3947,N_4188);
nand U5086 (N_5086,N_3483,N_3567);
nand U5087 (N_5087,N_4017,N_3530);
nand U5088 (N_5088,N_4246,N_4360);
nor U5089 (N_5089,N_3456,N_3091);
and U5090 (N_5090,N_3889,N_3565);
nor U5091 (N_5091,N_3851,N_3254);
nor U5092 (N_5092,N_3825,N_3430);
and U5093 (N_5093,N_4391,N_3904);
nand U5094 (N_5094,N_3962,N_4305);
and U5095 (N_5095,N_3375,N_3992);
and U5096 (N_5096,N_3242,N_4007);
nor U5097 (N_5097,N_3446,N_3846);
or U5098 (N_5098,N_3062,N_4367);
and U5099 (N_5099,N_4452,N_4224);
and U5100 (N_5100,N_4354,N_4373);
nand U5101 (N_5101,N_3536,N_4417);
and U5102 (N_5102,N_3273,N_3761);
nand U5103 (N_5103,N_3951,N_4478);
and U5104 (N_5104,N_3691,N_3009);
and U5105 (N_5105,N_4241,N_3543);
xnor U5106 (N_5106,N_4211,N_4409);
nand U5107 (N_5107,N_3720,N_3788);
or U5108 (N_5108,N_3812,N_3400);
nand U5109 (N_5109,N_3485,N_4397);
nor U5110 (N_5110,N_4074,N_4103);
nand U5111 (N_5111,N_3342,N_3291);
nand U5112 (N_5112,N_3599,N_4389);
or U5113 (N_5113,N_3210,N_3596);
nand U5114 (N_5114,N_3335,N_4064);
nand U5115 (N_5115,N_3302,N_3541);
nand U5116 (N_5116,N_3579,N_4152);
and U5117 (N_5117,N_3778,N_3619);
or U5118 (N_5118,N_4176,N_3194);
nand U5119 (N_5119,N_3104,N_3649);
or U5120 (N_5120,N_4298,N_3465);
nand U5121 (N_5121,N_3114,N_3678);
or U5122 (N_5122,N_4021,N_3544);
nor U5123 (N_5123,N_3955,N_4471);
and U5124 (N_5124,N_3583,N_3373);
nand U5125 (N_5125,N_4039,N_3239);
nor U5126 (N_5126,N_3379,N_3067);
or U5127 (N_5127,N_3350,N_3638);
nand U5128 (N_5128,N_4014,N_3030);
or U5129 (N_5129,N_4488,N_4087);
nor U5130 (N_5130,N_4431,N_3227);
and U5131 (N_5131,N_4036,N_3888);
or U5132 (N_5132,N_3197,N_3058);
or U5133 (N_5133,N_3893,N_4090);
nand U5134 (N_5134,N_3911,N_3925);
nand U5135 (N_5135,N_4089,N_4175);
nand U5136 (N_5136,N_3382,N_4202);
nor U5137 (N_5137,N_3328,N_3050);
or U5138 (N_5138,N_3702,N_3717);
or U5139 (N_5139,N_4491,N_3532);
nand U5140 (N_5140,N_4181,N_3762);
nor U5141 (N_5141,N_4024,N_3463);
nand U5142 (N_5142,N_4423,N_3420);
nand U5143 (N_5143,N_3442,N_3038);
or U5144 (N_5144,N_4002,N_3615);
or U5145 (N_5145,N_3772,N_4254);
and U5146 (N_5146,N_3699,N_3671);
or U5147 (N_5147,N_3685,N_3032);
nand U5148 (N_5148,N_4351,N_4053);
or U5149 (N_5149,N_4101,N_3895);
and U5150 (N_5150,N_4078,N_3867);
and U5151 (N_5151,N_4358,N_3491);
nand U5152 (N_5152,N_4341,N_3354);
nor U5153 (N_5153,N_3260,N_3924);
or U5154 (N_5154,N_3633,N_3387);
and U5155 (N_5155,N_4433,N_4131);
nor U5156 (N_5156,N_3085,N_3946);
nand U5157 (N_5157,N_3990,N_4364);
or U5158 (N_5158,N_3969,N_3974);
nor U5159 (N_5159,N_3013,N_3628);
and U5160 (N_5160,N_3341,N_4486);
or U5161 (N_5161,N_4314,N_3917);
or U5162 (N_5162,N_4442,N_3508);
nor U5163 (N_5163,N_3680,N_3215);
nor U5164 (N_5164,N_3195,N_3182);
or U5165 (N_5165,N_3383,N_3153);
or U5166 (N_5166,N_4184,N_3088);
or U5167 (N_5167,N_3126,N_4091);
and U5168 (N_5168,N_3324,N_3509);
or U5169 (N_5169,N_3987,N_3433);
nand U5170 (N_5170,N_3366,N_4263);
nand U5171 (N_5171,N_3824,N_4218);
or U5172 (N_5172,N_4406,N_4161);
nand U5173 (N_5173,N_3129,N_3833);
and U5174 (N_5174,N_3958,N_3137);
or U5175 (N_5175,N_3841,N_3470);
nand U5176 (N_5176,N_3650,N_3096);
nor U5177 (N_5177,N_3094,N_3245);
or U5178 (N_5178,N_3940,N_3880);
nand U5179 (N_5179,N_4426,N_3923);
and U5180 (N_5180,N_3820,N_4293);
or U5181 (N_5181,N_3817,N_3473);
nor U5182 (N_5182,N_4319,N_3167);
and U5183 (N_5183,N_4276,N_3507);
nor U5184 (N_5184,N_3118,N_4401);
and U5185 (N_5185,N_3576,N_3368);
or U5186 (N_5186,N_3738,N_3362);
nand U5187 (N_5187,N_3256,N_4056);
nor U5188 (N_5188,N_3316,N_3395);
xnor U5189 (N_5189,N_4250,N_4281);
nor U5190 (N_5190,N_3586,N_3945);
and U5191 (N_5191,N_3986,N_3903);
or U5192 (N_5192,N_4363,N_3343);
nand U5193 (N_5193,N_3661,N_3531);
and U5194 (N_5194,N_3623,N_4027);
nor U5195 (N_5195,N_4060,N_3322);
nor U5196 (N_5196,N_3568,N_3230);
nand U5197 (N_5197,N_3915,N_4209);
or U5198 (N_5198,N_4316,N_3914);
nor U5199 (N_5199,N_4386,N_3282);
nor U5200 (N_5200,N_4112,N_3518);
nor U5201 (N_5201,N_4072,N_3021);
and U5202 (N_5202,N_3977,N_3694);
nor U5203 (N_5203,N_4085,N_3225);
and U5204 (N_5204,N_3687,N_3645);
nor U5205 (N_5205,N_4346,N_3920);
nand U5206 (N_5206,N_3090,N_4350);
nor U5207 (N_5207,N_3190,N_3143);
xnor U5208 (N_5208,N_3588,N_3289);
nand U5209 (N_5209,N_3390,N_3734);
or U5210 (N_5210,N_4096,N_3135);
nand U5211 (N_5211,N_3852,N_3557);
nor U5212 (N_5212,N_3475,N_3451);
or U5213 (N_5213,N_3396,N_3138);
nand U5214 (N_5214,N_3724,N_4125);
nor U5215 (N_5215,N_3755,N_4133);
nand U5216 (N_5216,N_4190,N_4357);
nor U5217 (N_5217,N_4179,N_3719);
nand U5218 (N_5218,N_3074,N_3231);
xor U5219 (N_5219,N_3016,N_3556);
nor U5220 (N_5220,N_4362,N_3614);
and U5221 (N_5221,N_3217,N_3318);
or U5222 (N_5222,N_3998,N_4355);
and U5223 (N_5223,N_3635,N_3398);
nand U5224 (N_5224,N_3503,N_4379);
nand U5225 (N_5225,N_4140,N_3921);
nand U5226 (N_5226,N_3018,N_3611);
nand U5227 (N_5227,N_4287,N_4425);
or U5228 (N_5228,N_3773,N_3742);
or U5229 (N_5229,N_4322,N_3655);
nand U5230 (N_5230,N_4051,N_3415);
or U5231 (N_5231,N_3754,N_4439);
and U5232 (N_5232,N_3600,N_4163);
and U5233 (N_5233,N_3292,N_4443);
and U5234 (N_5234,N_3689,N_3617);
nor U5235 (N_5235,N_3495,N_3101);
or U5236 (N_5236,N_4186,N_3744);
nand U5237 (N_5237,N_4203,N_3730);
nor U5238 (N_5238,N_4337,N_4453);
nand U5239 (N_5239,N_3098,N_3970);
nor U5240 (N_5240,N_3061,N_4123);
or U5241 (N_5241,N_3954,N_3044);
nand U5242 (N_5242,N_3019,N_3107);
nor U5243 (N_5243,N_3697,N_3497);
and U5244 (N_5244,N_4065,N_3500);
nor U5245 (N_5245,N_4410,N_4199);
and U5246 (N_5246,N_4304,N_3875);
nand U5247 (N_5247,N_3790,N_4073);
and U5248 (N_5248,N_3751,N_3976);
and U5249 (N_5249,N_3412,N_3785);
nor U5250 (N_5250,N_3976,N_3178);
and U5251 (N_5251,N_4383,N_3326);
and U5252 (N_5252,N_3073,N_3928);
nor U5253 (N_5253,N_4020,N_4317);
or U5254 (N_5254,N_3336,N_4029);
nor U5255 (N_5255,N_4083,N_3378);
and U5256 (N_5256,N_4460,N_3865);
or U5257 (N_5257,N_4308,N_3910);
and U5258 (N_5258,N_3832,N_3654);
or U5259 (N_5259,N_3673,N_4086);
and U5260 (N_5260,N_3724,N_4197);
and U5261 (N_5261,N_3597,N_3736);
or U5262 (N_5262,N_4376,N_3947);
nor U5263 (N_5263,N_3535,N_3590);
and U5264 (N_5264,N_3992,N_3011);
or U5265 (N_5265,N_3255,N_3930);
xnor U5266 (N_5266,N_3074,N_4033);
xor U5267 (N_5267,N_3045,N_3624);
or U5268 (N_5268,N_4338,N_4266);
or U5269 (N_5269,N_3390,N_4094);
or U5270 (N_5270,N_4488,N_3414);
nand U5271 (N_5271,N_3826,N_4185);
nand U5272 (N_5272,N_3667,N_3872);
or U5273 (N_5273,N_3577,N_4073);
and U5274 (N_5274,N_4259,N_4444);
and U5275 (N_5275,N_3341,N_3650);
or U5276 (N_5276,N_3858,N_3914);
and U5277 (N_5277,N_3026,N_3462);
or U5278 (N_5278,N_4164,N_3010);
and U5279 (N_5279,N_4116,N_3027);
and U5280 (N_5280,N_4301,N_3926);
xor U5281 (N_5281,N_4062,N_4195);
nand U5282 (N_5282,N_3340,N_3934);
and U5283 (N_5283,N_4018,N_3555);
nor U5284 (N_5284,N_3264,N_3010);
or U5285 (N_5285,N_4154,N_3267);
or U5286 (N_5286,N_4269,N_3704);
nand U5287 (N_5287,N_4426,N_3594);
or U5288 (N_5288,N_3935,N_3093);
nor U5289 (N_5289,N_3875,N_3712);
and U5290 (N_5290,N_3715,N_4480);
nor U5291 (N_5291,N_3806,N_3684);
nand U5292 (N_5292,N_4321,N_4269);
and U5293 (N_5293,N_3443,N_4404);
or U5294 (N_5294,N_3519,N_3625);
or U5295 (N_5295,N_3888,N_3499);
or U5296 (N_5296,N_3766,N_3606);
or U5297 (N_5297,N_4497,N_3294);
and U5298 (N_5298,N_3357,N_4433);
nand U5299 (N_5299,N_3932,N_4063);
and U5300 (N_5300,N_4316,N_3664);
or U5301 (N_5301,N_3181,N_3962);
nand U5302 (N_5302,N_4033,N_3966);
and U5303 (N_5303,N_3424,N_3394);
and U5304 (N_5304,N_4026,N_4052);
and U5305 (N_5305,N_3655,N_3355);
or U5306 (N_5306,N_3035,N_4226);
nand U5307 (N_5307,N_4025,N_3186);
or U5308 (N_5308,N_3828,N_3226);
nor U5309 (N_5309,N_3102,N_4109);
nand U5310 (N_5310,N_4192,N_4228);
nor U5311 (N_5311,N_4493,N_4290);
or U5312 (N_5312,N_4005,N_4070);
nor U5313 (N_5313,N_3182,N_3978);
nand U5314 (N_5314,N_3571,N_3959);
and U5315 (N_5315,N_3047,N_4225);
or U5316 (N_5316,N_4257,N_4024);
and U5317 (N_5317,N_3302,N_3735);
or U5318 (N_5318,N_4084,N_3413);
nor U5319 (N_5319,N_3702,N_4297);
nand U5320 (N_5320,N_4329,N_3934);
or U5321 (N_5321,N_3306,N_4317);
nand U5322 (N_5322,N_3709,N_3885);
and U5323 (N_5323,N_4437,N_3548);
and U5324 (N_5324,N_3092,N_3969);
or U5325 (N_5325,N_3446,N_4495);
or U5326 (N_5326,N_3122,N_3660);
or U5327 (N_5327,N_3803,N_3873);
or U5328 (N_5328,N_3369,N_3452);
nor U5329 (N_5329,N_3283,N_3023);
and U5330 (N_5330,N_4339,N_4020);
and U5331 (N_5331,N_3562,N_4390);
nor U5332 (N_5332,N_3300,N_3848);
and U5333 (N_5333,N_3736,N_3532);
nand U5334 (N_5334,N_4440,N_3759);
or U5335 (N_5335,N_3238,N_3699);
and U5336 (N_5336,N_3920,N_4000);
or U5337 (N_5337,N_3896,N_3557);
nand U5338 (N_5338,N_3205,N_4231);
nand U5339 (N_5339,N_3746,N_3854);
nor U5340 (N_5340,N_3753,N_4142);
and U5341 (N_5341,N_3307,N_3837);
nand U5342 (N_5342,N_3589,N_3330);
and U5343 (N_5343,N_3276,N_3318);
nand U5344 (N_5344,N_3380,N_3544);
and U5345 (N_5345,N_3353,N_3929);
and U5346 (N_5346,N_4240,N_4115);
nor U5347 (N_5347,N_4290,N_4402);
nand U5348 (N_5348,N_3715,N_3636);
or U5349 (N_5349,N_4063,N_3282);
and U5350 (N_5350,N_3899,N_4049);
and U5351 (N_5351,N_3012,N_3557);
or U5352 (N_5352,N_3191,N_3254);
nor U5353 (N_5353,N_3915,N_3014);
nor U5354 (N_5354,N_3807,N_4444);
and U5355 (N_5355,N_3144,N_4358);
nor U5356 (N_5356,N_4100,N_4058);
nand U5357 (N_5357,N_3751,N_3980);
and U5358 (N_5358,N_3944,N_3868);
and U5359 (N_5359,N_3397,N_3723);
or U5360 (N_5360,N_3047,N_3060);
or U5361 (N_5361,N_4410,N_3933);
nor U5362 (N_5362,N_4348,N_3993);
nand U5363 (N_5363,N_3176,N_3346);
and U5364 (N_5364,N_3456,N_3287);
nand U5365 (N_5365,N_4132,N_3362);
xnor U5366 (N_5366,N_3345,N_4082);
or U5367 (N_5367,N_4436,N_4434);
and U5368 (N_5368,N_4412,N_4489);
and U5369 (N_5369,N_4042,N_3327);
nand U5370 (N_5370,N_3304,N_3992);
nor U5371 (N_5371,N_3277,N_3290);
nor U5372 (N_5372,N_3637,N_4146);
nor U5373 (N_5373,N_3311,N_3737);
and U5374 (N_5374,N_3332,N_3287);
nand U5375 (N_5375,N_3837,N_3271);
or U5376 (N_5376,N_3108,N_3151);
or U5377 (N_5377,N_3539,N_3433);
or U5378 (N_5378,N_3373,N_4141);
or U5379 (N_5379,N_4243,N_4246);
or U5380 (N_5380,N_3308,N_4203);
and U5381 (N_5381,N_3444,N_3774);
or U5382 (N_5382,N_4333,N_3795);
nand U5383 (N_5383,N_4218,N_4065);
or U5384 (N_5384,N_3921,N_3125);
and U5385 (N_5385,N_3791,N_3865);
nand U5386 (N_5386,N_3813,N_4009);
nand U5387 (N_5387,N_3491,N_3578);
and U5388 (N_5388,N_3650,N_4409);
nand U5389 (N_5389,N_4456,N_3038);
nor U5390 (N_5390,N_3076,N_3409);
or U5391 (N_5391,N_3777,N_3234);
and U5392 (N_5392,N_3109,N_3725);
and U5393 (N_5393,N_4166,N_4167);
nor U5394 (N_5394,N_3966,N_4156);
and U5395 (N_5395,N_3061,N_3153);
nand U5396 (N_5396,N_4496,N_3076);
and U5397 (N_5397,N_3962,N_4145);
and U5398 (N_5398,N_3001,N_3614);
nor U5399 (N_5399,N_4035,N_3119);
or U5400 (N_5400,N_3265,N_4496);
nand U5401 (N_5401,N_3399,N_4137);
nor U5402 (N_5402,N_3810,N_3225);
and U5403 (N_5403,N_3800,N_4162);
nor U5404 (N_5404,N_3197,N_4076);
nand U5405 (N_5405,N_4330,N_4124);
or U5406 (N_5406,N_3914,N_4279);
or U5407 (N_5407,N_3687,N_3400);
and U5408 (N_5408,N_3260,N_3000);
nand U5409 (N_5409,N_4357,N_4318);
and U5410 (N_5410,N_4189,N_4482);
nand U5411 (N_5411,N_3154,N_4360);
and U5412 (N_5412,N_3682,N_4128);
and U5413 (N_5413,N_3501,N_3224);
and U5414 (N_5414,N_4134,N_3411);
nor U5415 (N_5415,N_3246,N_3467);
nand U5416 (N_5416,N_3988,N_3716);
and U5417 (N_5417,N_3474,N_3273);
nand U5418 (N_5418,N_3931,N_4451);
nand U5419 (N_5419,N_3410,N_3942);
and U5420 (N_5420,N_3595,N_3253);
nand U5421 (N_5421,N_4321,N_3516);
or U5422 (N_5422,N_3506,N_3938);
nand U5423 (N_5423,N_3517,N_3577);
nor U5424 (N_5424,N_3116,N_3925);
and U5425 (N_5425,N_3255,N_4351);
nand U5426 (N_5426,N_3035,N_3343);
nand U5427 (N_5427,N_3607,N_4280);
nor U5428 (N_5428,N_4094,N_3412);
nor U5429 (N_5429,N_3958,N_3412);
and U5430 (N_5430,N_3497,N_3317);
or U5431 (N_5431,N_3390,N_4028);
or U5432 (N_5432,N_4438,N_3745);
nand U5433 (N_5433,N_4403,N_3101);
nand U5434 (N_5434,N_3148,N_4129);
or U5435 (N_5435,N_4492,N_3685);
nor U5436 (N_5436,N_4323,N_3187);
nand U5437 (N_5437,N_3284,N_3155);
nand U5438 (N_5438,N_3999,N_3009);
nor U5439 (N_5439,N_3421,N_4461);
nor U5440 (N_5440,N_4288,N_3718);
nand U5441 (N_5441,N_4165,N_4086);
nor U5442 (N_5442,N_3297,N_3666);
and U5443 (N_5443,N_3027,N_4149);
nor U5444 (N_5444,N_3985,N_4462);
nand U5445 (N_5445,N_4112,N_3260);
or U5446 (N_5446,N_3369,N_3843);
nor U5447 (N_5447,N_3787,N_3070);
or U5448 (N_5448,N_4200,N_3270);
xnor U5449 (N_5449,N_3986,N_3202);
and U5450 (N_5450,N_4042,N_3134);
nand U5451 (N_5451,N_4190,N_4230);
nand U5452 (N_5452,N_4035,N_3042);
nor U5453 (N_5453,N_3206,N_3161);
and U5454 (N_5454,N_3392,N_3033);
nand U5455 (N_5455,N_4263,N_3653);
and U5456 (N_5456,N_4299,N_4444);
nor U5457 (N_5457,N_4406,N_3472);
or U5458 (N_5458,N_4445,N_4320);
nor U5459 (N_5459,N_4304,N_4216);
and U5460 (N_5460,N_3557,N_3789);
or U5461 (N_5461,N_3177,N_3708);
and U5462 (N_5462,N_4344,N_3319);
nand U5463 (N_5463,N_3674,N_3438);
nor U5464 (N_5464,N_3260,N_4231);
or U5465 (N_5465,N_3514,N_3204);
xor U5466 (N_5466,N_4367,N_4373);
and U5467 (N_5467,N_3773,N_3792);
nor U5468 (N_5468,N_3545,N_4103);
or U5469 (N_5469,N_3153,N_3215);
nor U5470 (N_5470,N_3589,N_3615);
and U5471 (N_5471,N_3501,N_3899);
nor U5472 (N_5472,N_4400,N_4059);
or U5473 (N_5473,N_3962,N_3718);
and U5474 (N_5474,N_3961,N_3537);
nor U5475 (N_5475,N_3511,N_3046);
nor U5476 (N_5476,N_4426,N_4344);
nand U5477 (N_5477,N_4104,N_3674);
nand U5478 (N_5478,N_3799,N_3747);
nor U5479 (N_5479,N_3805,N_3907);
or U5480 (N_5480,N_4466,N_4332);
or U5481 (N_5481,N_3975,N_3581);
or U5482 (N_5482,N_3846,N_4305);
nor U5483 (N_5483,N_4356,N_3042);
nor U5484 (N_5484,N_4053,N_4346);
and U5485 (N_5485,N_3819,N_3182);
or U5486 (N_5486,N_4317,N_3346);
nor U5487 (N_5487,N_3653,N_4443);
nor U5488 (N_5488,N_4101,N_3751);
xor U5489 (N_5489,N_3098,N_3648);
nand U5490 (N_5490,N_4432,N_3240);
nor U5491 (N_5491,N_4295,N_4110);
nand U5492 (N_5492,N_3790,N_3093);
nor U5493 (N_5493,N_4451,N_3661);
nand U5494 (N_5494,N_4069,N_4418);
or U5495 (N_5495,N_4402,N_4179);
nor U5496 (N_5496,N_4388,N_3882);
or U5497 (N_5497,N_3302,N_3758);
or U5498 (N_5498,N_4281,N_3667);
nand U5499 (N_5499,N_4067,N_3243);
nor U5500 (N_5500,N_4100,N_4172);
nand U5501 (N_5501,N_3630,N_3664);
nand U5502 (N_5502,N_4405,N_3682);
and U5503 (N_5503,N_3920,N_3805);
or U5504 (N_5504,N_3247,N_3113);
nand U5505 (N_5505,N_4058,N_3933);
nand U5506 (N_5506,N_4032,N_4195);
or U5507 (N_5507,N_3805,N_3733);
nand U5508 (N_5508,N_3488,N_3121);
or U5509 (N_5509,N_4310,N_4374);
nand U5510 (N_5510,N_3755,N_3347);
nand U5511 (N_5511,N_4240,N_3759);
nor U5512 (N_5512,N_3879,N_3673);
nor U5513 (N_5513,N_3639,N_4416);
and U5514 (N_5514,N_4263,N_3854);
nor U5515 (N_5515,N_3117,N_4201);
or U5516 (N_5516,N_3244,N_4226);
and U5517 (N_5517,N_4408,N_3444);
nand U5518 (N_5518,N_3053,N_4121);
or U5519 (N_5519,N_3615,N_3441);
and U5520 (N_5520,N_3747,N_3145);
or U5521 (N_5521,N_4079,N_3068);
nand U5522 (N_5522,N_4182,N_3534);
nand U5523 (N_5523,N_3606,N_3430);
and U5524 (N_5524,N_4431,N_3586);
nand U5525 (N_5525,N_3529,N_4471);
nand U5526 (N_5526,N_3419,N_3044);
nor U5527 (N_5527,N_3502,N_3332);
or U5528 (N_5528,N_3536,N_4393);
and U5529 (N_5529,N_4265,N_3653);
xor U5530 (N_5530,N_4340,N_3708);
and U5531 (N_5531,N_3413,N_3989);
or U5532 (N_5532,N_3162,N_4381);
and U5533 (N_5533,N_4419,N_3866);
nor U5534 (N_5534,N_4303,N_3063);
or U5535 (N_5535,N_3640,N_3550);
and U5536 (N_5536,N_3095,N_4191);
or U5537 (N_5537,N_3211,N_3426);
xor U5538 (N_5538,N_3500,N_3122);
nand U5539 (N_5539,N_4129,N_3221);
and U5540 (N_5540,N_3577,N_3750);
nand U5541 (N_5541,N_4318,N_3647);
nand U5542 (N_5542,N_4378,N_3459);
nor U5543 (N_5543,N_4470,N_3883);
nor U5544 (N_5544,N_3477,N_4428);
nand U5545 (N_5545,N_4251,N_3493);
and U5546 (N_5546,N_4083,N_4478);
nand U5547 (N_5547,N_3255,N_3099);
nand U5548 (N_5548,N_3830,N_3897);
or U5549 (N_5549,N_4243,N_4302);
or U5550 (N_5550,N_4387,N_3044);
or U5551 (N_5551,N_3936,N_3799);
nand U5552 (N_5552,N_3308,N_3823);
nor U5553 (N_5553,N_4223,N_4136);
nand U5554 (N_5554,N_4457,N_3772);
and U5555 (N_5555,N_4419,N_3129);
or U5556 (N_5556,N_3191,N_4232);
nand U5557 (N_5557,N_3325,N_3095);
and U5558 (N_5558,N_3788,N_3264);
nor U5559 (N_5559,N_3074,N_4210);
and U5560 (N_5560,N_3372,N_3646);
nand U5561 (N_5561,N_4416,N_4307);
nor U5562 (N_5562,N_3519,N_4073);
nor U5563 (N_5563,N_3660,N_4230);
nand U5564 (N_5564,N_3951,N_4337);
nand U5565 (N_5565,N_3498,N_3996);
and U5566 (N_5566,N_4264,N_3002);
nor U5567 (N_5567,N_4197,N_3560);
nor U5568 (N_5568,N_4093,N_4393);
and U5569 (N_5569,N_3112,N_3205);
nor U5570 (N_5570,N_3148,N_3654);
or U5571 (N_5571,N_3690,N_3022);
nand U5572 (N_5572,N_4292,N_4137);
or U5573 (N_5573,N_3187,N_3769);
nand U5574 (N_5574,N_4335,N_3073);
or U5575 (N_5575,N_3747,N_3243);
or U5576 (N_5576,N_3437,N_3060);
nand U5577 (N_5577,N_4427,N_4377);
or U5578 (N_5578,N_3940,N_3689);
and U5579 (N_5579,N_3458,N_4478);
or U5580 (N_5580,N_3855,N_4124);
nor U5581 (N_5581,N_3831,N_3718);
or U5582 (N_5582,N_3259,N_4328);
nor U5583 (N_5583,N_4317,N_4052);
nor U5584 (N_5584,N_4389,N_4023);
nand U5585 (N_5585,N_3891,N_3616);
or U5586 (N_5586,N_3475,N_4379);
nor U5587 (N_5587,N_3151,N_4042);
or U5588 (N_5588,N_4411,N_3393);
nand U5589 (N_5589,N_3296,N_4075);
nand U5590 (N_5590,N_4023,N_3537);
nand U5591 (N_5591,N_3806,N_4145);
nor U5592 (N_5592,N_3915,N_3601);
nor U5593 (N_5593,N_4449,N_3635);
and U5594 (N_5594,N_3221,N_4495);
or U5595 (N_5595,N_4470,N_3646);
or U5596 (N_5596,N_4372,N_3173);
nand U5597 (N_5597,N_3675,N_3391);
nor U5598 (N_5598,N_3059,N_3648);
nor U5599 (N_5599,N_3732,N_3008);
or U5600 (N_5600,N_3281,N_3398);
nor U5601 (N_5601,N_3618,N_3370);
or U5602 (N_5602,N_3214,N_4438);
nor U5603 (N_5603,N_3539,N_4454);
nor U5604 (N_5604,N_3772,N_4272);
or U5605 (N_5605,N_3662,N_4079);
or U5606 (N_5606,N_4107,N_4142);
nand U5607 (N_5607,N_3020,N_4390);
nor U5608 (N_5608,N_3265,N_3143);
or U5609 (N_5609,N_3524,N_4110);
nand U5610 (N_5610,N_3600,N_4381);
nor U5611 (N_5611,N_4062,N_3876);
and U5612 (N_5612,N_3611,N_3115);
and U5613 (N_5613,N_3253,N_3594);
nor U5614 (N_5614,N_3043,N_4481);
and U5615 (N_5615,N_3014,N_3971);
and U5616 (N_5616,N_3120,N_3307);
nand U5617 (N_5617,N_3683,N_3068);
or U5618 (N_5618,N_3885,N_4482);
and U5619 (N_5619,N_3736,N_3720);
xor U5620 (N_5620,N_4208,N_3412);
nor U5621 (N_5621,N_3829,N_3126);
and U5622 (N_5622,N_3562,N_3186);
xor U5623 (N_5623,N_3772,N_4329);
or U5624 (N_5624,N_3889,N_4239);
and U5625 (N_5625,N_3108,N_4330);
and U5626 (N_5626,N_3029,N_3573);
or U5627 (N_5627,N_4012,N_4309);
nor U5628 (N_5628,N_3950,N_4145);
and U5629 (N_5629,N_4358,N_3133);
and U5630 (N_5630,N_4050,N_4269);
or U5631 (N_5631,N_3233,N_3415);
and U5632 (N_5632,N_3285,N_3210);
and U5633 (N_5633,N_3886,N_4022);
and U5634 (N_5634,N_3997,N_4161);
nand U5635 (N_5635,N_3218,N_3784);
nand U5636 (N_5636,N_3713,N_3402);
and U5637 (N_5637,N_3329,N_3314);
nor U5638 (N_5638,N_3263,N_4172);
nor U5639 (N_5639,N_3182,N_4033);
and U5640 (N_5640,N_4114,N_3486);
nand U5641 (N_5641,N_3242,N_4419);
and U5642 (N_5642,N_4058,N_4380);
or U5643 (N_5643,N_4322,N_3159);
nand U5644 (N_5644,N_3793,N_3650);
nor U5645 (N_5645,N_3686,N_4084);
nand U5646 (N_5646,N_4375,N_3099);
and U5647 (N_5647,N_4342,N_3953);
nand U5648 (N_5648,N_3325,N_4457);
and U5649 (N_5649,N_4456,N_3662);
or U5650 (N_5650,N_3651,N_4030);
and U5651 (N_5651,N_3216,N_3255);
and U5652 (N_5652,N_3952,N_3754);
or U5653 (N_5653,N_3196,N_3248);
or U5654 (N_5654,N_4202,N_3357);
and U5655 (N_5655,N_3906,N_4227);
and U5656 (N_5656,N_3549,N_3894);
and U5657 (N_5657,N_4174,N_3072);
nand U5658 (N_5658,N_3811,N_3436);
and U5659 (N_5659,N_4102,N_3342);
nand U5660 (N_5660,N_3631,N_4342);
or U5661 (N_5661,N_3601,N_3497);
or U5662 (N_5662,N_3082,N_3437);
nand U5663 (N_5663,N_3557,N_3906);
or U5664 (N_5664,N_3353,N_4412);
xnor U5665 (N_5665,N_4398,N_3464);
nor U5666 (N_5666,N_4384,N_4377);
nand U5667 (N_5667,N_4380,N_3830);
nand U5668 (N_5668,N_3036,N_3861);
nand U5669 (N_5669,N_3353,N_3548);
and U5670 (N_5670,N_4017,N_3075);
nor U5671 (N_5671,N_4432,N_4399);
and U5672 (N_5672,N_3719,N_4285);
nand U5673 (N_5673,N_4028,N_4264);
xnor U5674 (N_5674,N_4114,N_4142);
or U5675 (N_5675,N_3154,N_3106);
and U5676 (N_5676,N_4329,N_4233);
nor U5677 (N_5677,N_4205,N_4199);
nor U5678 (N_5678,N_3375,N_3161);
or U5679 (N_5679,N_4338,N_3619);
nand U5680 (N_5680,N_3148,N_3053);
or U5681 (N_5681,N_3094,N_4472);
nand U5682 (N_5682,N_3056,N_4491);
and U5683 (N_5683,N_4176,N_3741);
and U5684 (N_5684,N_4365,N_4092);
nand U5685 (N_5685,N_3132,N_4388);
nand U5686 (N_5686,N_3144,N_3624);
nand U5687 (N_5687,N_3034,N_3126);
and U5688 (N_5688,N_3555,N_4404);
or U5689 (N_5689,N_4170,N_4123);
or U5690 (N_5690,N_4250,N_4186);
or U5691 (N_5691,N_3701,N_4329);
nand U5692 (N_5692,N_3695,N_3059);
or U5693 (N_5693,N_3410,N_4413);
nand U5694 (N_5694,N_3274,N_4274);
nor U5695 (N_5695,N_3800,N_3278);
and U5696 (N_5696,N_4140,N_3897);
nor U5697 (N_5697,N_4409,N_3855);
nand U5698 (N_5698,N_3750,N_3340);
or U5699 (N_5699,N_4314,N_3313);
nor U5700 (N_5700,N_3607,N_3170);
or U5701 (N_5701,N_3449,N_3008);
and U5702 (N_5702,N_3325,N_4222);
nand U5703 (N_5703,N_4359,N_3382);
nand U5704 (N_5704,N_3792,N_3551);
nor U5705 (N_5705,N_4062,N_3598);
and U5706 (N_5706,N_3168,N_4457);
xnor U5707 (N_5707,N_4479,N_3356);
nand U5708 (N_5708,N_3305,N_4012);
or U5709 (N_5709,N_4327,N_3729);
and U5710 (N_5710,N_3309,N_3568);
nor U5711 (N_5711,N_3609,N_3055);
or U5712 (N_5712,N_4350,N_3689);
and U5713 (N_5713,N_3431,N_3380);
nor U5714 (N_5714,N_3049,N_3750);
nand U5715 (N_5715,N_3068,N_3163);
nand U5716 (N_5716,N_3349,N_3384);
nand U5717 (N_5717,N_3744,N_4276);
or U5718 (N_5718,N_3863,N_3190);
and U5719 (N_5719,N_4468,N_3171);
or U5720 (N_5720,N_3046,N_4107);
nor U5721 (N_5721,N_3478,N_3055);
nand U5722 (N_5722,N_3629,N_3405);
or U5723 (N_5723,N_4163,N_4003);
nand U5724 (N_5724,N_4091,N_3147);
or U5725 (N_5725,N_4476,N_4185);
nor U5726 (N_5726,N_3919,N_3829);
nand U5727 (N_5727,N_3300,N_3115);
or U5728 (N_5728,N_3146,N_4176);
or U5729 (N_5729,N_3835,N_4195);
or U5730 (N_5730,N_4371,N_4101);
or U5731 (N_5731,N_4445,N_3575);
nand U5732 (N_5732,N_4418,N_4268);
and U5733 (N_5733,N_3240,N_3055);
nand U5734 (N_5734,N_3426,N_3296);
nand U5735 (N_5735,N_4112,N_4310);
nor U5736 (N_5736,N_4281,N_3900);
nand U5737 (N_5737,N_4290,N_3903);
and U5738 (N_5738,N_4156,N_3525);
and U5739 (N_5739,N_4393,N_4308);
or U5740 (N_5740,N_3990,N_3996);
and U5741 (N_5741,N_4093,N_4100);
nor U5742 (N_5742,N_4091,N_4266);
and U5743 (N_5743,N_3437,N_3911);
nor U5744 (N_5744,N_3523,N_4025);
or U5745 (N_5745,N_4001,N_3444);
or U5746 (N_5746,N_3550,N_3211);
nand U5747 (N_5747,N_3900,N_3857);
and U5748 (N_5748,N_3414,N_3404);
or U5749 (N_5749,N_3463,N_4259);
or U5750 (N_5750,N_3186,N_3451);
or U5751 (N_5751,N_3474,N_4457);
or U5752 (N_5752,N_3280,N_3804);
nor U5753 (N_5753,N_3882,N_3152);
nand U5754 (N_5754,N_4235,N_3194);
or U5755 (N_5755,N_4161,N_4209);
and U5756 (N_5756,N_4231,N_4453);
nor U5757 (N_5757,N_3034,N_3594);
or U5758 (N_5758,N_3768,N_3631);
and U5759 (N_5759,N_3785,N_3934);
nand U5760 (N_5760,N_3074,N_4364);
and U5761 (N_5761,N_3622,N_4209);
nor U5762 (N_5762,N_4301,N_3360);
and U5763 (N_5763,N_3487,N_3012);
or U5764 (N_5764,N_4171,N_3193);
or U5765 (N_5765,N_4333,N_3121);
or U5766 (N_5766,N_3629,N_3239);
nor U5767 (N_5767,N_3013,N_3814);
nand U5768 (N_5768,N_3146,N_3277);
and U5769 (N_5769,N_3296,N_4041);
and U5770 (N_5770,N_3034,N_3592);
or U5771 (N_5771,N_3454,N_3763);
nand U5772 (N_5772,N_3149,N_4137);
and U5773 (N_5773,N_3874,N_3458);
and U5774 (N_5774,N_3682,N_3451);
nor U5775 (N_5775,N_3751,N_3343);
and U5776 (N_5776,N_4183,N_4063);
nand U5777 (N_5777,N_3752,N_3780);
and U5778 (N_5778,N_3343,N_3211);
or U5779 (N_5779,N_4164,N_3634);
and U5780 (N_5780,N_4374,N_3425);
nand U5781 (N_5781,N_3854,N_3861);
and U5782 (N_5782,N_3016,N_4189);
and U5783 (N_5783,N_3184,N_4312);
or U5784 (N_5784,N_4479,N_4222);
and U5785 (N_5785,N_4432,N_3816);
nand U5786 (N_5786,N_4385,N_3189);
or U5787 (N_5787,N_4372,N_3126);
and U5788 (N_5788,N_3342,N_4138);
nor U5789 (N_5789,N_3779,N_4428);
nor U5790 (N_5790,N_3843,N_4117);
nand U5791 (N_5791,N_4216,N_4116);
nor U5792 (N_5792,N_3454,N_3213);
and U5793 (N_5793,N_3879,N_4259);
and U5794 (N_5794,N_3619,N_4160);
nand U5795 (N_5795,N_3851,N_4284);
nand U5796 (N_5796,N_3717,N_3272);
nor U5797 (N_5797,N_3658,N_3411);
and U5798 (N_5798,N_4268,N_3210);
or U5799 (N_5799,N_4321,N_3434);
nand U5800 (N_5800,N_3184,N_3352);
or U5801 (N_5801,N_3158,N_4360);
nand U5802 (N_5802,N_3427,N_3776);
and U5803 (N_5803,N_4176,N_3746);
nand U5804 (N_5804,N_3507,N_3765);
nand U5805 (N_5805,N_3419,N_3168);
nand U5806 (N_5806,N_3392,N_4205);
and U5807 (N_5807,N_4040,N_3927);
or U5808 (N_5808,N_3409,N_3963);
or U5809 (N_5809,N_4371,N_3462);
nor U5810 (N_5810,N_4283,N_3037);
nor U5811 (N_5811,N_3303,N_3700);
nand U5812 (N_5812,N_4205,N_3380);
xnor U5813 (N_5813,N_4426,N_4474);
nand U5814 (N_5814,N_4247,N_3500);
nand U5815 (N_5815,N_3856,N_3383);
and U5816 (N_5816,N_4283,N_3347);
or U5817 (N_5817,N_4074,N_3438);
and U5818 (N_5818,N_4020,N_4296);
and U5819 (N_5819,N_4371,N_4031);
or U5820 (N_5820,N_3199,N_4289);
and U5821 (N_5821,N_3716,N_3471);
nand U5822 (N_5822,N_4051,N_3820);
nor U5823 (N_5823,N_4225,N_3034);
nor U5824 (N_5824,N_3300,N_4469);
nand U5825 (N_5825,N_3761,N_4042);
nand U5826 (N_5826,N_4078,N_3167);
nand U5827 (N_5827,N_3093,N_3038);
or U5828 (N_5828,N_4391,N_3616);
and U5829 (N_5829,N_3158,N_3724);
or U5830 (N_5830,N_4009,N_4154);
nor U5831 (N_5831,N_3690,N_3805);
and U5832 (N_5832,N_3709,N_3932);
or U5833 (N_5833,N_4273,N_3503);
nor U5834 (N_5834,N_4214,N_3238);
nand U5835 (N_5835,N_4316,N_3550);
nor U5836 (N_5836,N_3951,N_3932);
and U5837 (N_5837,N_3146,N_3586);
and U5838 (N_5838,N_3093,N_3456);
or U5839 (N_5839,N_3694,N_3608);
nand U5840 (N_5840,N_4485,N_4400);
nand U5841 (N_5841,N_3229,N_3349);
nor U5842 (N_5842,N_3433,N_4495);
or U5843 (N_5843,N_3660,N_3651);
or U5844 (N_5844,N_3746,N_4388);
and U5845 (N_5845,N_3717,N_3397);
nor U5846 (N_5846,N_3991,N_3826);
or U5847 (N_5847,N_4259,N_3618);
and U5848 (N_5848,N_3861,N_3148);
or U5849 (N_5849,N_4346,N_3389);
nand U5850 (N_5850,N_3276,N_3356);
nand U5851 (N_5851,N_4399,N_3932);
and U5852 (N_5852,N_3199,N_3883);
nor U5853 (N_5853,N_4236,N_3595);
and U5854 (N_5854,N_3586,N_3565);
nand U5855 (N_5855,N_4317,N_3738);
and U5856 (N_5856,N_4349,N_4482);
nor U5857 (N_5857,N_4405,N_4359);
or U5858 (N_5858,N_4280,N_3189);
and U5859 (N_5859,N_4131,N_4377);
nand U5860 (N_5860,N_3962,N_4118);
and U5861 (N_5861,N_3958,N_3066);
nand U5862 (N_5862,N_4125,N_3458);
nor U5863 (N_5863,N_3825,N_4330);
nand U5864 (N_5864,N_4025,N_3500);
nor U5865 (N_5865,N_3601,N_3593);
and U5866 (N_5866,N_3549,N_4326);
nand U5867 (N_5867,N_3929,N_3760);
nand U5868 (N_5868,N_3344,N_4333);
nand U5869 (N_5869,N_3956,N_3682);
nand U5870 (N_5870,N_3278,N_4433);
or U5871 (N_5871,N_4282,N_3244);
nand U5872 (N_5872,N_3825,N_3100);
or U5873 (N_5873,N_3331,N_4275);
nor U5874 (N_5874,N_3428,N_3218);
nand U5875 (N_5875,N_3964,N_3713);
nor U5876 (N_5876,N_3786,N_4312);
nor U5877 (N_5877,N_4485,N_4160);
or U5878 (N_5878,N_3659,N_3991);
nor U5879 (N_5879,N_4329,N_4478);
and U5880 (N_5880,N_3239,N_3015);
nand U5881 (N_5881,N_3865,N_3986);
nor U5882 (N_5882,N_3160,N_3861);
and U5883 (N_5883,N_3865,N_3217);
nand U5884 (N_5884,N_3792,N_3994);
nor U5885 (N_5885,N_3379,N_3978);
or U5886 (N_5886,N_3836,N_4018);
nand U5887 (N_5887,N_4411,N_3278);
nor U5888 (N_5888,N_3372,N_4190);
nand U5889 (N_5889,N_4231,N_3309);
and U5890 (N_5890,N_3187,N_3688);
nor U5891 (N_5891,N_4113,N_3275);
or U5892 (N_5892,N_3605,N_4380);
nor U5893 (N_5893,N_3733,N_3538);
nor U5894 (N_5894,N_3737,N_3673);
nor U5895 (N_5895,N_4017,N_4189);
or U5896 (N_5896,N_4490,N_4073);
nor U5897 (N_5897,N_3935,N_4341);
nor U5898 (N_5898,N_4402,N_4309);
nor U5899 (N_5899,N_3843,N_4346);
and U5900 (N_5900,N_3305,N_3851);
nor U5901 (N_5901,N_3914,N_3131);
nand U5902 (N_5902,N_4014,N_3614);
xor U5903 (N_5903,N_3461,N_4385);
nand U5904 (N_5904,N_4386,N_3958);
nand U5905 (N_5905,N_3784,N_3976);
and U5906 (N_5906,N_4131,N_3388);
xnor U5907 (N_5907,N_3191,N_3828);
or U5908 (N_5908,N_3493,N_3647);
nor U5909 (N_5909,N_3385,N_4083);
nor U5910 (N_5910,N_3728,N_4034);
and U5911 (N_5911,N_3848,N_4204);
nand U5912 (N_5912,N_3659,N_3458);
or U5913 (N_5913,N_4291,N_3436);
nor U5914 (N_5914,N_3342,N_3428);
or U5915 (N_5915,N_3673,N_3600);
nor U5916 (N_5916,N_3746,N_4298);
nand U5917 (N_5917,N_4394,N_4113);
nand U5918 (N_5918,N_4399,N_4147);
and U5919 (N_5919,N_4367,N_3939);
nor U5920 (N_5920,N_3745,N_3576);
nand U5921 (N_5921,N_4247,N_4414);
nand U5922 (N_5922,N_4449,N_3891);
nor U5923 (N_5923,N_4374,N_4026);
and U5924 (N_5924,N_3161,N_4490);
and U5925 (N_5925,N_4399,N_3583);
and U5926 (N_5926,N_3750,N_4451);
nand U5927 (N_5927,N_4484,N_3818);
and U5928 (N_5928,N_3030,N_3486);
nand U5929 (N_5929,N_4237,N_4437);
nand U5930 (N_5930,N_3553,N_3068);
or U5931 (N_5931,N_4246,N_4280);
nand U5932 (N_5932,N_3834,N_3370);
or U5933 (N_5933,N_4373,N_4384);
nand U5934 (N_5934,N_3722,N_3888);
nor U5935 (N_5935,N_3746,N_4425);
nor U5936 (N_5936,N_3466,N_3598);
and U5937 (N_5937,N_3319,N_4364);
nand U5938 (N_5938,N_3211,N_3094);
and U5939 (N_5939,N_4461,N_4271);
and U5940 (N_5940,N_3077,N_4401);
nand U5941 (N_5941,N_3251,N_4294);
and U5942 (N_5942,N_4047,N_3988);
nand U5943 (N_5943,N_3262,N_3649);
nor U5944 (N_5944,N_4011,N_3891);
xnor U5945 (N_5945,N_3103,N_4378);
or U5946 (N_5946,N_4498,N_4117);
or U5947 (N_5947,N_4126,N_4426);
nand U5948 (N_5948,N_3475,N_3943);
nand U5949 (N_5949,N_3653,N_3677);
or U5950 (N_5950,N_4173,N_3944);
and U5951 (N_5951,N_3565,N_3216);
and U5952 (N_5952,N_3083,N_4026);
and U5953 (N_5953,N_3301,N_3554);
nand U5954 (N_5954,N_4385,N_4404);
and U5955 (N_5955,N_4319,N_3275);
nand U5956 (N_5956,N_3201,N_3318);
nand U5957 (N_5957,N_4121,N_3481);
or U5958 (N_5958,N_3223,N_3522);
and U5959 (N_5959,N_3458,N_4275);
and U5960 (N_5960,N_3530,N_3169);
nor U5961 (N_5961,N_4245,N_3158);
or U5962 (N_5962,N_3427,N_4482);
and U5963 (N_5963,N_3383,N_4126);
or U5964 (N_5964,N_4317,N_3956);
or U5965 (N_5965,N_4317,N_4443);
nand U5966 (N_5966,N_4495,N_4356);
or U5967 (N_5967,N_3063,N_4089);
nand U5968 (N_5968,N_3853,N_3104);
nand U5969 (N_5969,N_4093,N_3766);
or U5970 (N_5970,N_3288,N_3019);
nand U5971 (N_5971,N_4099,N_3822);
nor U5972 (N_5972,N_3674,N_3320);
nor U5973 (N_5973,N_4494,N_3417);
nor U5974 (N_5974,N_3326,N_4422);
nor U5975 (N_5975,N_4306,N_3711);
nor U5976 (N_5976,N_3369,N_3050);
or U5977 (N_5977,N_3778,N_4320);
nand U5978 (N_5978,N_4135,N_3399);
nand U5979 (N_5979,N_3601,N_4365);
or U5980 (N_5980,N_3574,N_3515);
nor U5981 (N_5981,N_3713,N_3715);
nor U5982 (N_5982,N_3588,N_4295);
or U5983 (N_5983,N_4229,N_3479);
and U5984 (N_5984,N_4390,N_3494);
and U5985 (N_5985,N_3186,N_4426);
or U5986 (N_5986,N_4368,N_3467);
nor U5987 (N_5987,N_3577,N_3915);
nor U5988 (N_5988,N_4041,N_4228);
nor U5989 (N_5989,N_4025,N_4091);
and U5990 (N_5990,N_3398,N_3881);
and U5991 (N_5991,N_3477,N_4010);
nand U5992 (N_5992,N_3075,N_3870);
nor U5993 (N_5993,N_4443,N_4074);
and U5994 (N_5994,N_3881,N_3778);
or U5995 (N_5995,N_3310,N_3425);
or U5996 (N_5996,N_3262,N_3985);
nand U5997 (N_5997,N_3400,N_3965);
nor U5998 (N_5998,N_3902,N_4150);
and U5999 (N_5999,N_3992,N_3402);
nand U6000 (N_6000,N_5241,N_5287);
nor U6001 (N_6001,N_5879,N_5814);
nor U6002 (N_6002,N_5930,N_5871);
or U6003 (N_6003,N_4506,N_4617);
nand U6004 (N_6004,N_4794,N_4786);
or U6005 (N_6005,N_4827,N_5670);
nand U6006 (N_6006,N_5615,N_5932);
or U6007 (N_6007,N_4881,N_4503);
or U6008 (N_6008,N_4672,N_4998);
and U6009 (N_6009,N_4890,N_5053);
nand U6010 (N_6010,N_5583,N_5321);
and U6011 (N_6011,N_5128,N_5412);
or U6012 (N_6012,N_4835,N_4846);
or U6013 (N_6013,N_5338,N_5268);
nor U6014 (N_6014,N_4746,N_4787);
or U6015 (N_6015,N_4957,N_5774);
nand U6016 (N_6016,N_5194,N_5870);
or U6017 (N_6017,N_5980,N_4984);
nand U6018 (N_6018,N_5675,N_5815);
and U6019 (N_6019,N_5666,N_4988);
nor U6020 (N_6020,N_5999,N_5979);
or U6021 (N_6021,N_4513,N_4934);
nor U6022 (N_6022,N_5405,N_5007);
nor U6023 (N_6023,N_5488,N_5586);
or U6024 (N_6024,N_4959,N_4833);
nor U6025 (N_6025,N_4917,N_5643);
and U6026 (N_6026,N_5107,N_5334);
and U6027 (N_6027,N_5428,N_4812);
nand U6028 (N_6028,N_5411,N_4990);
nand U6029 (N_6029,N_5136,N_4622);
nor U6030 (N_6030,N_4640,N_5937);
and U6031 (N_6031,N_4875,N_5591);
or U6032 (N_6032,N_4508,N_4913);
nor U6033 (N_6033,N_5475,N_5792);
or U6034 (N_6034,N_4755,N_4578);
or U6035 (N_6035,N_5968,N_5523);
or U6036 (N_6036,N_5348,N_5333);
or U6037 (N_6037,N_5209,N_5202);
and U6038 (N_6038,N_4981,N_5876);
nand U6039 (N_6039,N_4546,N_5365);
or U6040 (N_6040,N_5878,N_5469);
or U6041 (N_6041,N_4790,N_5441);
and U6042 (N_6042,N_5808,N_4541);
nor U6043 (N_6043,N_4977,N_4710);
nand U6044 (N_6044,N_5032,N_5204);
nor U6045 (N_6045,N_4500,N_5948);
nor U6046 (N_6046,N_5433,N_5279);
nor U6047 (N_6047,N_5703,N_5788);
or U6048 (N_6048,N_5942,N_5851);
xnor U6049 (N_6049,N_5250,N_5843);
and U6050 (N_6050,N_5350,N_4894);
nor U6051 (N_6051,N_5579,N_4570);
nor U6052 (N_6052,N_4825,N_4861);
and U6053 (N_6053,N_4597,N_5751);
and U6054 (N_6054,N_5067,N_4751);
nor U6055 (N_6055,N_4901,N_5787);
nand U6056 (N_6056,N_5259,N_5595);
or U6057 (N_6057,N_5311,N_5035);
or U6058 (N_6058,N_5904,N_4590);
or U6059 (N_6059,N_5885,N_4902);
nor U6060 (N_6060,N_5533,N_4769);
nand U6061 (N_6061,N_4759,N_5526);
nand U6062 (N_6062,N_5477,N_5087);
and U6063 (N_6063,N_5802,N_5747);
or U6064 (N_6064,N_4719,N_5654);
or U6065 (N_6065,N_5228,N_5418);
nand U6066 (N_6066,N_5356,N_5465);
nand U6067 (N_6067,N_5599,N_5807);
and U6068 (N_6068,N_5688,N_5380);
or U6069 (N_6069,N_5436,N_5375);
or U6070 (N_6070,N_5247,N_4528);
nand U6071 (N_6071,N_5264,N_4594);
nand U6072 (N_6072,N_5818,N_5946);
nor U6073 (N_6073,N_5208,N_5978);
nand U6074 (N_6074,N_5507,N_5112);
and U6075 (N_6075,N_4591,N_5759);
and U6076 (N_6076,N_4515,N_5221);
nor U6077 (N_6077,N_5455,N_5622);
nor U6078 (N_6078,N_5327,N_5297);
and U6079 (N_6079,N_5163,N_5237);
nand U6080 (N_6080,N_5608,N_5026);
or U6081 (N_6081,N_5600,N_4615);
or U6082 (N_6082,N_4932,N_5200);
or U6083 (N_6083,N_5379,N_5960);
nand U6084 (N_6084,N_5116,N_5423);
or U6085 (N_6085,N_5308,N_4763);
or U6086 (N_6086,N_5407,N_4952);
nor U6087 (N_6087,N_5076,N_4983);
or U6088 (N_6088,N_5520,N_5033);
or U6089 (N_6089,N_4668,N_4664);
nor U6090 (N_6090,N_5636,N_4946);
nor U6091 (N_6091,N_5660,N_4726);
nor U6092 (N_6092,N_5577,N_5668);
and U6093 (N_6093,N_4967,N_5013);
and U6094 (N_6094,N_5552,N_5069);
nor U6095 (N_6095,N_4539,N_4625);
and U6096 (N_6096,N_5425,N_5664);
nand U6097 (N_6097,N_5752,N_5830);
and U6098 (N_6098,N_4855,N_5746);
nand U6099 (N_6099,N_5711,N_5722);
and U6100 (N_6100,N_5037,N_5039);
and U6101 (N_6101,N_5716,N_4750);
and U6102 (N_6102,N_5219,N_5998);
nand U6103 (N_6103,N_4580,N_5663);
and U6104 (N_6104,N_5971,N_5385);
nor U6105 (N_6105,N_5789,N_5314);
nand U6106 (N_6106,N_5610,N_5189);
or U6107 (N_6107,N_5854,N_5175);
nand U6108 (N_6108,N_5148,N_5881);
nor U6109 (N_6109,N_5681,N_5972);
nor U6110 (N_6110,N_5938,N_5933);
nand U6111 (N_6111,N_5756,N_5392);
nand U6112 (N_6112,N_5563,N_5238);
nand U6113 (N_6113,N_5042,N_5626);
or U6114 (N_6114,N_5757,N_5578);
nor U6115 (N_6115,N_5531,N_5955);
nand U6116 (N_6116,N_4607,N_5398);
and U6117 (N_6117,N_5060,N_5165);
or U6118 (N_6118,N_4814,N_5918);
and U6119 (N_6119,N_4791,N_4912);
nor U6120 (N_6120,N_5289,N_4840);
and U6121 (N_6121,N_5750,N_5827);
or U6122 (N_6122,N_5656,N_5288);
or U6123 (N_6123,N_5482,N_4837);
or U6124 (N_6124,N_4898,N_5653);
and U6125 (N_6125,N_4511,N_5928);
nand U6126 (N_6126,N_5139,N_4799);
or U6127 (N_6127,N_4976,N_5905);
or U6128 (N_6128,N_5995,N_5466);
nand U6129 (N_6129,N_5419,N_5280);
and U6130 (N_6130,N_4699,N_4757);
or U6131 (N_6131,N_4658,N_5718);
nor U6132 (N_6132,N_5501,N_5158);
nor U6133 (N_6133,N_5129,N_5066);
and U6134 (N_6134,N_5431,N_5273);
nand U6135 (N_6135,N_5853,N_5902);
nand U6136 (N_6136,N_5147,N_5882);
nor U6137 (N_6137,N_5731,N_5335);
or U6138 (N_6138,N_4659,N_5456);
nand U6139 (N_6139,N_4850,N_5068);
or U6140 (N_6140,N_5406,N_5554);
and U6141 (N_6141,N_5893,N_5263);
or U6142 (N_6142,N_5645,N_5628);
nand U6143 (N_6143,N_4953,N_4880);
and U6144 (N_6144,N_5100,N_5230);
xnor U6145 (N_6145,N_4639,N_5201);
nand U6146 (N_6146,N_4765,N_5498);
or U6147 (N_6147,N_5266,N_5292);
nor U6148 (N_6148,N_5071,N_5006);
and U6149 (N_6149,N_4738,N_5721);
or U6150 (N_6150,N_5867,N_4691);
nand U6151 (N_6151,N_5420,N_5040);
nand U6152 (N_6152,N_4651,N_5801);
or U6153 (N_6153,N_5001,N_4903);
and U6154 (N_6154,N_5614,N_5530);
or U6155 (N_6155,N_4978,N_4773);
or U6156 (N_6156,N_4793,N_5872);
nand U6157 (N_6157,N_5640,N_5063);
nand U6158 (N_6158,N_5239,N_5075);
and U6159 (N_6159,N_5157,N_4713);
or U6160 (N_6160,N_5778,N_4676);
nor U6161 (N_6161,N_5355,N_4925);
or U6162 (N_6162,N_4756,N_5144);
and U6163 (N_6163,N_5499,N_4845);
nand U6164 (N_6164,N_4944,N_5088);
and U6165 (N_6165,N_5771,N_5492);
or U6166 (N_6166,N_4857,N_4636);
nand U6167 (N_6167,N_5700,N_5537);
and U6168 (N_6168,N_5191,N_4975);
nand U6169 (N_6169,N_5549,N_4531);
or U6170 (N_6170,N_5319,N_5059);
and U6171 (N_6171,N_5278,N_5984);
nor U6172 (N_6172,N_4721,N_4993);
nand U6173 (N_6173,N_5835,N_5803);
or U6174 (N_6174,N_5956,N_4911);
nand U6175 (N_6175,N_5233,N_5326);
or U6176 (N_6176,N_5532,N_5570);
nand U6177 (N_6177,N_5251,N_4781);
nand U6178 (N_6178,N_4551,N_5495);
nand U6179 (N_6179,N_5305,N_5766);
nor U6180 (N_6180,N_5647,N_5582);
and U6181 (N_6181,N_5565,N_5220);
nand U6182 (N_6182,N_4667,N_4961);
nor U6183 (N_6183,N_5486,N_4542);
and U6184 (N_6184,N_4574,N_4628);
and U6185 (N_6185,N_5849,N_5895);
and U6186 (N_6186,N_5439,N_5396);
or U6187 (N_6187,N_4821,N_5702);
and U6188 (N_6188,N_5360,N_4777);
nand U6189 (N_6189,N_5672,N_5038);
nand U6190 (N_6190,N_5864,N_4882);
and U6191 (N_6191,N_5625,N_5502);
nor U6192 (N_6192,N_5755,N_4657);
nor U6193 (N_6193,N_4697,N_5254);
or U6194 (N_6194,N_5354,N_5836);
nor U6195 (N_6195,N_5317,N_4963);
and U6196 (N_6196,N_4991,N_5080);
or U6197 (N_6197,N_4899,N_4836);
or U6198 (N_6198,N_5353,N_5991);
nor U6199 (N_6199,N_4569,N_4938);
or U6200 (N_6200,N_5503,N_5667);
nand U6201 (N_6201,N_4908,N_5318);
nand U6202 (N_6202,N_5468,N_5917);
or U6203 (N_6203,N_4631,N_5840);
nand U6204 (N_6204,N_5581,N_5519);
and U6205 (N_6205,N_4645,N_4516);
and U6206 (N_6206,N_5105,N_4728);
and U6207 (N_6207,N_5696,N_4604);
and U6208 (N_6208,N_5467,N_5249);
and U6209 (N_6209,N_4867,N_5648);
and U6210 (N_6210,N_5546,N_5868);
or U6211 (N_6211,N_4758,N_5939);
nor U6212 (N_6212,N_5886,N_5203);
nor U6213 (N_6213,N_5393,N_5715);
or U6214 (N_6214,N_5291,N_5437);
and U6215 (N_6215,N_5720,N_5739);
or U6216 (N_6216,N_4620,N_5275);
nor U6217 (N_6217,N_5394,N_5661);
nand U6218 (N_6218,N_5847,N_4919);
nand U6219 (N_6219,N_4895,N_5142);
nor U6220 (N_6220,N_4596,N_4807);
nand U6221 (N_6221,N_5497,N_4655);
nand U6222 (N_6222,N_5265,N_4583);
or U6223 (N_6223,N_5812,N_4588);
or U6224 (N_6224,N_5769,N_4599);
or U6225 (N_6225,N_5440,N_5103);
nand U6226 (N_6226,N_4815,N_5281);
or U6227 (N_6227,N_5062,N_5257);
or U6228 (N_6228,N_5235,N_5434);
or U6229 (N_6229,N_4892,N_5206);
nand U6230 (N_6230,N_5816,N_5464);
nor U6231 (N_6231,N_5368,N_5585);
nor U6232 (N_6232,N_5382,N_4740);
nand U6233 (N_6233,N_5186,N_5953);
nor U6234 (N_6234,N_4562,N_4711);
or U6235 (N_6235,N_5635,N_5331);
and U6236 (N_6236,N_5262,N_5791);
or U6237 (N_6237,N_5470,N_5008);
and U6238 (N_6238,N_5480,N_5458);
nand U6239 (N_6239,N_4709,N_5992);
or U6240 (N_6240,N_4571,N_5985);
or U6241 (N_6241,N_5555,N_4810);
and U6242 (N_6242,N_5810,N_4708);
or U6243 (N_6243,N_4884,N_4730);
nor U6244 (N_6244,N_5556,N_5424);
nor U6245 (N_6245,N_5034,N_4842);
nor U6246 (N_6246,N_5115,N_5146);
or U6247 (N_6247,N_5574,N_5962);
nor U6248 (N_6248,N_5179,N_5003);
nor U6249 (N_6249,N_5779,N_4572);
nand U6250 (N_6250,N_4962,N_4669);
nand U6251 (N_6251,N_5121,N_5841);
and U6252 (N_6252,N_5374,N_5481);
nor U6253 (N_6253,N_5054,N_4703);
nor U6254 (N_6254,N_4598,N_5977);
nand U6255 (N_6255,N_4933,N_5196);
nand U6256 (N_6256,N_5997,N_5631);
nand U6257 (N_6257,N_5564,N_5457);
or U6258 (N_6258,N_5929,N_5414);
or U6259 (N_6259,N_5020,N_5234);
nor U6260 (N_6260,N_4512,N_4869);
nor U6261 (N_6261,N_5540,N_5861);
and U6262 (N_6262,N_5276,N_4841);
nand U6263 (N_6263,N_4966,N_5744);
or U6264 (N_6264,N_5347,N_5261);
and U6265 (N_6265,N_5964,N_4678);
nor U6266 (N_6266,N_5487,N_5214);
or U6267 (N_6267,N_5123,N_5073);
nand U6268 (N_6268,N_5567,N_5909);
nor U6269 (N_6269,N_5633,N_5652);
nor U6270 (N_6270,N_5361,N_5730);
nand U6271 (N_6271,N_5258,N_5912);
or U6272 (N_6272,N_4564,N_5126);
nor U6273 (N_6273,N_5114,N_5606);
nor U6274 (N_6274,N_4929,N_5785);
and U6275 (N_6275,N_5620,N_4679);
and U6276 (N_6276,N_5745,N_5869);
or U6277 (N_6277,N_5800,N_5517);
nand U6278 (N_6278,N_5012,N_4577);
and U6279 (N_6279,N_4712,N_5834);
and U6280 (N_6280,N_5435,N_4951);
and U6281 (N_6281,N_4600,N_5761);
nor U6282 (N_6282,N_5072,N_5575);
or U6283 (N_6283,N_4886,N_5920);
and U6284 (N_6284,N_4502,N_4715);
nor U6285 (N_6285,N_5557,N_5632);
nand U6286 (N_6286,N_5850,N_4762);
nand U6287 (N_6287,N_4656,N_5969);
nand U6288 (N_6288,N_5124,N_4538);
and U6289 (N_6289,N_5337,N_4930);
and U6290 (N_6290,N_5764,N_4973);
and U6291 (N_6291,N_5944,N_5504);
or U6292 (N_6292,N_5083,N_5132);
nor U6293 (N_6293,N_4947,N_5539);
nor U6294 (N_6294,N_4641,N_4960);
or U6295 (N_6295,N_5272,N_5438);
nand U6296 (N_6296,N_4563,N_5691);
or U6297 (N_6297,N_5036,N_5838);
or U6298 (N_6298,N_5547,N_4918);
or U6299 (N_6299,N_5400,N_4737);
nand U6300 (N_6300,N_5819,N_4839);
nor U6301 (N_6301,N_4732,N_5111);
nor U6302 (N_6302,N_5728,N_4870);
nor U6303 (N_6303,N_5174,N_5192);
and U6304 (N_6304,N_4540,N_5195);
or U6305 (N_6305,N_5223,N_5644);
or U6306 (N_6306,N_5940,N_5754);
or U6307 (N_6307,N_5908,N_4816);
and U6308 (N_6308,N_4614,N_5941);
and U6309 (N_6309,N_5889,N_5478);
nor U6310 (N_6310,N_5094,N_5358);
and U6311 (N_6311,N_4566,N_4956);
and U6312 (N_6312,N_4789,N_4921);
nor U6313 (N_6313,N_5176,N_4505);
nand U6314 (N_6314,N_5796,N_4865);
or U6315 (N_6315,N_5536,N_5710);
nor U6316 (N_6316,N_5910,N_5683);
nand U6317 (N_6317,N_4771,N_5029);
nor U6318 (N_6318,N_5322,N_5846);
or U6319 (N_6319,N_5044,N_4525);
or U6320 (N_6320,N_5863,N_4684);
xor U6321 (N_6321,N_5782,N_5994);
or U6322 (N_6322,N_4811,N_4647);
nor U6323 (N_6323,N_5155,N_5500);
or U6324 (N_6324,N_4927,N_5887);
nor U6325 (N_6325,N_4736,N_5270);
or U6326 (N_6326,N_5274,N_5429);
or U6327 (N_6327,N_4904,N_4748);
or U6328 (N_6328,N_5544,N_5023);
nand U6329 (N_6329,N_4584,N_4928);
and U6330 (N_6330,N_5762,N_5336);
and U6331 (N_6331,N_5826,N_4958);
nand U6332 (N_6332,N_4702,N_5133);
nor U6333 (N_6333,N_5805,N_5389);
and U6334 (N_6334,N_5187,N_5970);
nor U6335 (N_6335,N_4926,N_5216);
and U6336 (N_6336,N_5143,N_5590);
nor U6337 (N_6337,N_5852,N_5047);
nand U6338 (N_6338,N_5639,N_5104);
nor U6339 (N_6339,N_5516,N_5786);
and U6340 (N_6340,N_5089,N_4660);
or U6341 (N_6341,N_5253,N_5749);
nor U6342 (N_6342,N_4548,N_5024);
nor U6343 (N_6343,N_4831,N_5988);
nor U6344 (N_6344,N_4705,N_5588);
and U6345 (N_6345,N_5890,N_5943);
nand U6346 (N_6346,N_5106,N_5027);
or U6347 (N_6347,N_5426,N_5444);
or U6348 (N_6348,N_4948,N_5416);
nor U6349 (N_6349,N_5461,N_5198);
nor U6350 (N_6350,N_5213,N_5102);
nor U6351 (N_6351,N_5101,N_5952);
and U6352 (N_6352,N_4752,N_5476);
nand U6353 (N_6353,N_5733,N_4969);
nor U6354 (N_6354,N_5587,N_4729);
nor U6355 (N_6355,N_4545,N_4792);
or U6356 (N_6356,N_4767,N_5673);
nand U6357 (N_6357,N_5343,N_5282);
and U6358 (N_6358,N_5776,N_5513);
nand U6359 (N_6359,N_4685,N_4858);
nand U6360 (N_6360,N_4768,N_5430);
and U6361 (N_6361,N_4554,N_5099);
xnor U6362 (N_6362,N_5496,N_4995);
or U6363 (N_6363,N_4876,N_5596);
and U6364 (N_6364,N_5093,N_5646);
nand U6365 (N_6365,N_5432,N_5891);
or U6366 (N_6366,N_5658,N_4537);
nor U6367 (N_6367,N_4618,N_5659);
and U6368 (N_6368,N_5052,N_5491);
nand U6369 (N_6369,N_5451,N_5218);
nor U6370 (N_6370,N_5562,N_5580);
nor U6371 (N_6371,N_5357,N_5485);
and U6372 (N_6372,N_5914,N_4907);
or U6373 (N_6373,N_5415,N_5510);
and U6374 (N_6374,N_5760,N_5877);
nand U6375 (N_6375,N_5712,N_4783);
and U6376 (N_6376,N_5346,N_5010);
nand U6377 (N_6377,N_5168,N_4509);
or U6378 (N_6378,N_4828,N_5775);
nand U6379 (N_6379,N_5859,N_5684);
nand U6380 (N_6380,N_4897,N_4761);
nand U6381 (N_6381,N_5695,N_5138);
or U6382 (N_6382,N_5307,N_5309);
or U6383 (N_6383,N_5302,N_5922);
nand U6384 (N_6384,N_4695,N_5572);
nand U6385 (N_6385,N_5804,N_5641);
nor U6386 (N_6386,N_5450,N_4700);
or U6387 (N_6387,N_4868,N_4714);
and U6388 (N_6388,N_5260,N_5207);
nand U6389 (N_6389,N_4687,N_4813);
or U6390 (N_6390,N_4587,N_4915);
nor U6391 (N_6391,N_4605,N_4682);
and U6392 (N_6392,N_5915,N_5092);
or U6393 (N_6393,N_5898,N_5742);
nand U6394 (N_6394,N_5957,N_4873);
and U6395 (N_6395,N_5183,N_4671);
nor U6396 (N_6396,N_5848,N_5351);
xor U6397 (N_6397,N_4706,N_4611);
nor U6398 (N_6398,N_5427,N_4922);
or U6399 (N_6399,N_4996,N_5484);
and U6400 (N_6400,N_4782,N_5058);
nand U6401 (N_6401,N_4533,N_5171);
nand U6402 (N_6402,N_4725,N_5662);
and U6403 (N_6403,N_4866,N_4519);
and U6404 (N_6404,N_5773,N_4802);
nand U6405 (N_6405,N_4891,N_4940);
or U6406 (N_6406,N_5949,N_4510);
nor U6407 (N_6407,N_5387,N_5973);
nor U6408 (N_6408,N_5244,N_5874);
nand U6409 (N_6409,N_5597,N_5701);
or U6410 (N_6410,N_4637,N_4733);
or U6411 (N_6411,N_4801,N_5799);
nor U6412 (N_6412,N_4523,N_5443);
nand U6413 (N_6413,N_4749,N_5086);
nand U6414 (N_6414,N_5299,N_5125);
nand U6415 (N_6415,N_5657,N_4501);
nor U6416 (N_6416,N_5763,N_5592);
or U6417 (N_6417,N_5152,N_5185);
or U6418 (N_6418,N_5772,N_5388);
xor U6419 (N_6419,N_4621,N_5794);
and U6420 (N_6420,N_5137,N_5951);
or U6421 (N_6421,N_5873,N_5397);
nand U6422 (N_6422,N_5224,N_4734);
and U6423 (N_6423,N_5031,N_5018);
and U6424 (N_6424,N_4955,N_5151);
and U6425 (N_6425,N_4602,N_4559);
and U6426 (N_6426,N_5550,N_5091);
nor U6427 (N_6427,N_5506,N_5674);
or U6428 (N_6428,N_5736,N_4595);
nand U6429 (N_6429,N_5911,N_5097);
nand U6430 (N_6430,N_4673,N_5377);
or U6431 (N_6431,N_5950,N_4690);
and U6432 (N_6432,N_5623,N_4731);
nor U6433 (N_6433,N_5584,N_5896);
or U6434 (N_6434,N_5081,N_5837);
nor U6435 (N_6435,N_5806,N_5824);
or U6436 (N_6436,N_5271,N_4834);
nand U6437 (N_6437,N_5986,N_5817);
and U6438 (N_6438,N_5095,N_4661);
nor U6439 (N_6439,N_4633,N_5341);
nor U6440 (N_6440,N_5990,N_5593);
or U6441 (N_6441,N_5833,N_4601);
or U6442 (N_6442,N_5916,N_4754);
nand U6443 (N_6443,N_4923,N_4796);
or U6444 (N_6444,N_5931,N_5845);
or U6445 (N_6445,N_5677,N_5372);
and U6446 (N_6446,N_4644,N_5390);
and U6447 (N_6447,N_5611,N_5967);
nor U6448 (N_6448,N_5212,N_5051);
nor U6449 (N_6449,N_5795,N_5686);
nor U6450 (N_6450,N_5413,N_5935);
and U6451 (N_6451,N_5320,N_5541);
nand U6452 (N_6452,N_5605,N_4526);
nor U6453 (N_6453,N_5529,N_5188);
and U6454 (N_6454,N_4585,N_4819);
and U6455 (N_6455,N_5079,N_5924);
nor U6456 (N_6456,N_5630,N_5310);
or U6457 (N_6457,N_5777,N_5894);
or U6458 (N_6458,N_5906,N_5245);
nor U6459 (N_6459,N_4696,N_4677);
or U6460 (N_6460,N_5897,N_4507);
nor U6461 (N_6461,N_5511,N_4883);
nand U6462 (N_6462,N_5892,N_4534);
or U6463 (N_6463,N_5002,N_5162);
or U6464 (N_6464,N_4924,N_5923);
and U6465 (N_6465,N_5958,N_5522);
and U6466 (N_6466,N_4809,N_4608);
nand U6467 (N_6467,N_5243,N_4980);
or U6468 (N_6468,N_5449,N_4698);
and U6469 (N_6469,N_5726,N_4643);
or U6470 (N_6470,N_5323,N_4909);
and U6471 (N_6471,N_4735,N_4649);
nand U6472 (N_6472,N_4517,N_4889);
nand U6473 (N_6473,N_4775,N_4972);
nand U6474 (N_6474,N_4727,N_5154);
and U6475 (N_6475,N_5781,N_4527);
and U6476 (N_6476,N_5240,N_4674);
nand U6477 (N_6477,N_5493,N_4530);
and U6478 (N_6478,N_5021,N_5352);
nor U6479 (N_6479,N_4544,N_5727);
and U6480 (N_6480,N_5284,N_4560);
nor U6481 (N_6481,N_5370,N_5172);
or U6482 (N_6482,N_4558,N_4522);
and U6483 (N_6483,N_5134,N_5028);
nor U6484 (N_6484,N_4844,N_5118);
nor U6485 (N_6485,N_4985,N_5514);
and U6486 (N_6486,N_4627,N_5061);
nor U6487 (N_6487,N_4823,N_5373);
and U6488 (N_6488,N_4910,N_5056);
nor U6489 (N_6489,N_5490,N_5617);
and U6490 (N_6490,N_5559,N_4974);
nand U6491 (N_6491,N_5383,N_4616);
or U6492 (N_6492,N_5669,N_5880);
and U6493 (N_6493,N_5651,N_4798);
nor U6494 (N_6494,N_5576,N_5828);
and U6495 (N_6495,N_5793,N_5974);
nor U6496 (N_6496,N_4720,N_5452);
nor U6497 (N_6497,N_4680,N_5976);
nand U6498 (N_6498,N_5215,N_5011);
nand U6499 (N_6499,N_5145,N_4686);
and U6500 (N_6500,N_5131,N_4610);
nand U6501 (N_6501,N_4764,N_5589);
nand U6502 (N_6502,N_4612,N_5820);
nand U6503 (N_6503,N_5604,N_5164);
nor U6504 (N_6504,N_5098,N_4805);
nor U6505 (N_6505,N_5169,N_4654);
nand U6506 (N_6506,N_4994,N_4888);
nor U6507 (N_6507,N_4770,N_5831);
nor U6508 (N_6508,N_5705,N_5524);
and U6509 (N_6509,N_5734,N_5222);
nor U6510 (N_6510,N_5085,N_4854);
or U6511 (N_6511,N_4856,N_4646);
nor U6512 (N_6512,N_4688,N_5558);
nor U6513 (N_6513,N_4650,N_5921);
nor U6514 (N_6514,N_4986,N_5332);
or U6515 (N_6515,N_4532,N_5634);
or U6516 (N_6516,N_4634,N_4997);
or U6517 (N_6517,N_5982,N_5694);
nand U6518 (N_6518,N_4670,N_5638);
nor U6519 (N_6519,N_4666,N_5913);
nand U6520 (N_6520,N_5989,N_5573);
nand U6521 (N_6521,N_5560,N_5117);
or U6522 (N_6522,N_4935,N_4609);
and U6523 (N_6523,N_5603,N_5369);
nand U6524 (N_6524,N_4822,N_5494);
nor U6525 (N_6525,N_5410,N_5242);
nand U6526 (N_6526,N_5717,N_5016);
and U6527 (N_6527,N_5509,N_5609);
xnor U6528 (N_6528,N_5875,N_4629);
nand U6529 (N_6529,N_4520,N_4843);
nor U6530 (N_6530,N_4987,N_4518);
nand U6531 (N_6531,N_5790,N_5050);
nor U6532 (N_6532,N_4693,N_4784);
or U6533 (N_6533,N_5167,N_5678);
nor U6534 (N_6534,N_5655,N_5693);
nor U6535 (N_6535,N_4945,N_4536);
nand U6536 (N_6536,N_5697,N_4968);
nor U6537 (N_6537,N_5569,N_5065);
nor U6538 (N_6538,N_5542,N_5166);
or U6539 (N_6539,N_4852,N_4941);
nand U6540 (N_6540,N_4859,N_4999);
nand U6541 (N_6541,N_5304,N_5594);
nor U6542 (N_6542,N_4626,N_5566);
nand U6543 (N_6543,N_4896,N_5161);
nand U6544 (N_6544,N_5724,N_4905);
and U6545 (N_6545,N_5286,N_5000);
nor U6546 (N_6546,N_5190,N_5883);
and U6547 (N_6547,N_4879,N_5043);
nor U6548 (N_6548,N_5947,N_5709);
and U6549 (N_6549,N_4779,N_5489);
and U6550 (N_6550,N_5900,N_5090);
or U6551 (N_6551,N_4553,N_5809);
or U6552 (N_6552,N_5345,N_5707);
and U6553 (N_6553,N_4785,N_5865);
nor U6554 (N_6554,N_5505,N_5181);
xnor U6555 (N_6555,N_5538,N_5698);
nand U6556 (N_6556,N_4603,N_5135);
or U6557 (N_6557,N_5607,N_4795);
and U6558 (N_6558,N_5708,N_5723);
nor U6559 (N_6559,N_5740,N_5463);
nor U6560 (N_6560,N_4832,N_5535);
nor U6561 (N_6561,N_4623,N_5300);
and U6562 (N_6562,N_5231,N_5682);
nand U6563 (N_6563,N_5981,N_5680);
or U6564 (N_6564,N_5445,N_5621);
nor U6565 (N_6565,N_5363,N_4982);
or U6566 (N_6566,N_4906,N_5474);
or U6567 (N_6567,N_4878,N_5743);
or U6568 (N_6568,N_5844,N_4916);
nor U6569 (N_6569,N_5009,N_4653);
and U6570 (N_6570,N_5246,N_5899);
nor U6571 (N_6571,N_5184,N_4665);
nor U6572 (N_6572,N_5512,N_4683);
and U6573 (N_6573,N_4849,N_4630);
nand U6574 (N_6574,N_5294,N_5017);
nand U6575 (N_6575,N_5312,N_5177);
and U6576 (N_6576,N_4797,N_5765);
nor U6577 (N_6577,N_5741,N_4556);
nor U6578 (N_6578,N_5160,N_5619);
or U6579 (N_6579,N_4937,N_5401);
or U6580 (N_6580,N_5462,N_4642);
nor U6581 (N_6581,N_5903,N_5330);
and U6582 (N_6582,N_5735,N_4524);
nor U6583 (N_6583,N_5267,N_4561);
nor U6584 (N_6584,N_5127,N_5324);
nor U6585 (N_6585,N_5005,N_5855);
or U6586 (N_6586,N_5293,N_5315);
nand U6587 (N_6587,N_4826,N_5395);
nor U6588 (N_6588,N_4803,N_5367);
nor U6589 (N_6589,N_4514,N_5046);
nand U6590 (N_6590,N_5109,N_5901);
nand U6591 (N_6591,N_4549,N_4724);
nor U6592 (N_6592,N_5699,N_4900);
and U6593 (N_6593,N_5528,N_5856);
nand U6594 (N_6594,N_5961,N_4838);
and U6595 (N_6595,N_4589,N_5719);
and U6596 (N_6596,N_5409,N_4694);
and U6597 (N_6597,N_4971,N_5340);
and U6598 (N_6598,N_4864,N_5296);
nor U6599 (N_6599,N_5996,N_4954);
nor U6600 (N_6600,N_5758,N_4851);
and U6601 (N_6601,N_5022,N_5153);
nand U6602 (N_6602,N_5290,N_5983);
nand U6603 (N_6603,N_5770,N_5140);
nor U6604 (N_6604,N_5829,N_5534);
and U6605 (N_6605,N_5447,N_4776);
nand U6606 (N_6606,N_5704,N_5676);
nor U6607 (N_6607,N_5084,N_5601);
nand U6608 (N_6608,N_5687,N_5548);
or U6609 (N_6609,N_4943,N_4613);
or U6610 (N_6610,N_4808,N_5252);
and U6611 (N_6611,N_5078,N_5783);
or U6612 (N_6612,N_5422,N_5649);
and U6613 (N_6613,N_4565,N_5232);
or U6614 (N_6614,N_5460,N_5386);
or U6615 (N_6615,N_4745,N_5637);
nand U6616 (N_6616,N_5255,N_5738);
nor U6617 (N_6617,N_5515,N_4887);
nor U6618 (N_6618,N_5277,N_5193);
nand U6619 (N_6619,N_4872,N_4817);
nand U6620 (N_6620,N_5384,N_5842);
nand U6621 (N_6621,N_5884,N_4624);
nand U6622 (N_6622,N_5141,N_5295);
nand U6623 (N_6623,N_5074,N_5064);
nor U6624 (N_6624,N_5568,N_5963);
nand U6625 (N_6625,N_5329,N_4989);
nand U6626 (N_6626,N_5473,N_4753);
nand U6627 (N_6627,N_4555,N_5442);
and U6628 (N_6628,N_5987,N_5823);
nor U6629 (N_6629,N_5096,N_5627);
or U6630 (N_6630,N_4939,N_5399);
nor U6631 (N_6631,N_5170,N_5402);
or U6632 (N_6632,N_5954,N_5014);
nand U6633 (N_6633,N_4920,N_5376);
nand U6634 (N_6634,N_4521,N_4579);
or U6635 (N_6635,N_5325,N_5199);
or U6636 (N_6636,N_5182,N_4723);
nand U6637 (N_6637,N_4829,N_4979);
nand U6638 (N_6638,N_5618,N_5349);
nor U6639 (N_6639,N_5713,N_5725);
or U6640 (N_6640,N_4567,N_5448);
and U6641 (N_6641,N_5811,N_5553);
or U6642 (N_6642,N_5813,N_5689);
or U6643 (N_6643,N_5561,N_4965);
or U6644 (N_6644,N_4722,N_5381);
and U6645 (N_6645,N_4931,N_4582);
or U6646 (N_6646,N_5359,N_5342);
or U6647 (N_6647,N_4552,N_4778);
and U6648 (N_6648,N_4704,N_5934);
or U6649 (N_6649,N_5965,N_4593);
nand U6650 (N_6650,N_4830,N_4675);
nor U6651 (N_6651,N_5966,N_4744);
and U6652 (N_6652,N_5768,N_4635);
or U6653 (N_6653,N_5180,N_5454);
nand U6654 (N_6654,N_5403,N_5404);
and U6655 (N_6655,N_4914,N_5225);
or U6656 (N_6656,N_5945,N_4550);
or U6657 (N_6657,N_4586,N_5665);
or U6658 (N_6658,N_5748,N_5256);
nand U6659 (N_6659,N_5472,N_5690);
nand U6660 (N_6660,N_5925,N_4619);
or U6661 (N_6661,N_4741,N_4743);
nor U6662 (N_6662,N_5479,N_5518);
nand U6663 (N_6663,N_5119,N_4557);
or U6664 (N_6664,N_5366,N_5391);
and U6665 (N_6665,N_5825,N_5780);
nand U6666 (N_6666,N_5149,N_5571);
nand U6667 (N_6667,N_5862,N_5753);
and U6668 (N_6668,N_5459,N_5408);
or U6669 (N_6669,N_5993,N_4950);
nor U6670 (N_6670,N_4862,N_4681);
and U6671 (N_6671,N_5650,N_4529);
nor U6672 (N_6672,N_5298,N_4581);
or U6673 (N_6673,N_5371,N_5927);
nand U6674 (N_6674,N_5082,N_5729);
nand U6675 (N_6675,N_5839,N_4747);
nor U6676 (N_6676,N_4663,N_5858);
nand U6677 (N_6677,N_5421,N_5784);
and U6678 (N_6678,N_5378,N_5888);
nor U6679 (N_6679,N_5236,N_4717);
nor U6680 (N_6680,N_4874,N_4638);
nand U6681 (N_6681,N_5822,N_5303);
or U6682 (N_6682,N_4800,N_5269);
nand U6683 (N_6683,N_4718,N_4760);
nor U6684 (N_6684,N_5602,N_4632);
nand U6685 (N_6685,N_5598,N_5197);
nand U6686 (N_6686,N_4893,N_4606);
or U6687 (N_6687,N_5798,N_5210);
nor U6688 (N_6688,N_5364,N_5642);
or U6689 (N_6689,N_5316,N_5113);
nand U6690 (N_6690,N_5797,N_5205);
and U6691 (N_6691,N_5616,N_5313);
and U6692 (N_6692,N_5737,N_5866);
nand U6693 (N_6693,N_5679,N_5227);
or U6694 (N_6694,N_4780,N_4568);
nor U6695 (N_6695,N_4949,N_4774);
or U6696 (N_6696,N_4847,N_5907);
or U6697 (N_6697,N_5453,N_4824);
nor U6698 (N_6698,N_4739,N_5173);
or U6699 (N_6699,N_4772,N_5483);
and U6700 (N_6700,N_5417,N_5521);
nand U6701 (N_6701,N_5692,N_5077);
and U6702 (N_6702,N_4964,N_5229);
nor U6703 (N_6703,N_5545,N_5025);
nand U6704 (N_6704,N_4692,N_4871);
and U6705 (N_6705,N_5714,N_5049);
nor U6706 (N_6706,N_5821,N_5339);
nor U6707 (N_6707,N_4970,N_5612);
nor U6708 (N_6708,N_4860,N_4504);
and U6709 (N_6709,N_4820,N_4689);
or U6710 (N_6710,N_4575,N_4806);
xor U6711 (N_6711,N_5108,N_4701);
nand U6712 (N_6712,N_5527,N_4707);
nor U6713 (N_6713,N_5767,N_5045);
nor U6714 (N_6714,N_5362,N_4662);
and U6715 (N_6715,N_5159,N_5156);
or U6716 (N_6716,N_5732,N_5344);
and U6717 (N_6717,N_5015,N_4652);
nor U6718 (N_6718,N_4804,N_5936);
nand U6719 (N_6719,N_5226,N_4885);
and U6720 (N_6720,N_5122,N_4942);
and U6721 (N_6721,N_5030,N_5629);
and U6722 (N_6722,N_5328,N_5178);
and U6723 (N_6723,N_5471,N_5055);
or U6724 (N_6724,N_5624,N_5004);
nor U6725 (N_6725,N_5525,N_5211);
nand U6726 (N_6726,N_5706,N_5130);
xnor U6727 (N_6727,N_5508,N_5150);
and U6728 (N_6728,N_4716,N_4853);
nor U6729 (N_6729,N_5919,N_4543);
and U6730 (N_6730,N_5110,N_4547);
nand U6731 (N_6731,N_5019,N_4576);
nor U6732 (N_6732,N_4592,N_4535);
nand U6733 (N_6733,N_5832,N_4818);
or U6734 (N_6734,N_4863,N_5285);
nand U6735 (N_6735,N_5306,N_5048);
nor U6736 (N_6736,N_5857,N_5283);
or U6737 (N_6737,N_5551,N_4848);
or U6738 (N_6738,N_5301,N_5685);
nor U6739 (N_6739,N_5959,N_5120);
nor U6740 (N_6740,N_4788,N_4766);
or U6741 (N_6741,N_4992,N_5543);
or U6742 (N_6742,N_4936,N_5860);
xor U6743 (N_6743,N_4742,N_5070);
and U6744 (N_6744,N_5217,N_5926);
and U6745 (N_6745,N_5446,N_5613);
or U6746 (N_6746,N_5248,N_5041);
nor U6747 (N_6747,N_4648,N_5671);
and U6748 (N_6748,N_5975,N_5057);
and U6749 (N_6749,N_4573,N_4877);
and U6750 (N_6750,N_5669,N_4599);
or U6751 (N_6751,N_4711,N_4643);
nand U6752 (N_6752,N_4549,N_5363);
nand U6753 (N_6753,N_5486,N_4960);
and U6754 (N_6754,N_5685,N_5701);
and U6755 (N_6755,N_4537,N_5050);
and U6756 (N_6756,N_5732,N_5812);
or U6757 (N_6757,N_5258,N_5399);
or U6758 (N_6758,N_5406,N_4557);
or U6759 (N_6759,N_5841,N_5356);
and U6760 (N_6760,N_4717,N_5552);
nand U6761 (N_6761,N_4577,N_5258);
or U6762 (N_6762,N_5431,N_4953);
or U6763 (N_6763,N_4818,N_4770);
and U6764 (N_6764,N_4638,N_4850);
nand U6765 (N_6765,N_5997,N_5661);
nor U6766 (N_6766,N_5632,N_4961);
or U6767 (N_6767,N_5072,N_5396);
or U6768 (N_6768,N_5054,N_4718);
nor U6769 (N_6769,N_4596,N_5430);
nor U6770 (N_6770,N_5377,N_5117);
nor U6771 (N_6771,N_5079,N_5773);
and U6772 (N_6772,N_4596,N_5775);
nand U6773 (N_6773,N_5463,N_5328);
or U6774 (N_6774,N_5473,N_4625);
and U6775 (N_6775,N_4655,N_5978);
nand U6776 (N_6776,N_4913,N_5935);
or U6777 (N_6777,N_5304,N_4558);
or U6778 (N_6778,N_5374,N_4680);
nor U6779 (N_6779,N_5140,N_4694);
nor U6780 (N_6780,N_5505,N_5846);
nand U6781 (N_6781,N_5418,N_5617);
and U6782 (N_6782,N_5439,N_4820);
or U6783 (N_6783,N_4951,N_4833);
nand U6784 (N_6784,N_5276,N_5832);
nor U6785 (N_6785,N_5285,N_4626);
nand U6786 (N_6786,N_5500,N_4888);
nand U6787 (N_6787,N_5804,N_4547);
nand U6788 (N_6788,N_5285,N_5526);
nor U6789 (N_6789,N_5538,N_4901);
and U6790 (N_6790,N_4963,N_5136);
or U6791 (N_6791,N_4783,N_5723);
or U6792 (N_6792,N_4520,N_5478);
or U6793 (N_6793,N_5185,N_5846);
and U6794 (N_6794,N_5786,N_5662);
nor U6795 (N_6795,N_5700,N_4807);
or U6796 (N_6796,N_5505,N_5501);
or U6797 (N_6797,N_5350,N_5124);
nand U6798 (N_6798,N_5106,N_5264);
and U6799 (N_6799,N_5715,N_4879);
and U6800 (N_6800,N_5662,N_5265);
and U6801 (N_6801,N_5334,N_5295);
or U6802 (N_6802,N_5832,N_5579);
nor U6803 (N_6803,N_5504,N_5990);
and U6804 (N_6804,N_5051,N_5180);
or U6805 (N_6805,N_5364,N_5614);
nand U6806 (N_6806,N_4502,N_5351);
and U6807 (N_6807,N_5249,N_5029);
or U6808 (N_6808,N_5244,N_4724);
nand U6809 (N_6809,N_4958,N_5272);
or U6810 (N_6810,N_5993,N_5279);
or U6811 (N_6811,N_5641,N_4546);
nor U6812 (N_6812,N_5040,N_5264);
nor U6813 (N_6813,N_4939,N_5944);
nand U6814 (N_6814,N_5950,N_5311);
xor U6815 (N_6815,N_5200,N_5234);
nand U6816 (N_6816,N_4695,N_4935);
nor U6817 (N_6817,N_5687,N_5635);
or U6818 (N_6818,N_4678,N_4849);
nand U6819 (N_6819,N_5621,N_5118);
and U6820 (N_6820,N_5342,N_5203);
nand U6821 (N_6821,N_5874,N_5724);
or U6822 (N_6822,N_4722,N_5123);
and U6823 (N_6823,N_4581,N_4749);
nor U6824 (N_6824,N_5437,N_5705);
and U6825 (N_6825,N_5056,N_5070);
and U6826 (N_6826,N_5370,N_5025);
nand U6827 (N_6827,N_5281,N_5173);
nand U6828 (N_6828,N_5607,N_5191);
and U6829 (N_6829,N_5747,N_5230);
or U6830 (N_6830,N_5203,N_5713);
or U6831 (N_6831,N_4775,N_5268);
and U6832 (N_6832,N_4832,N_5021);
nor U6833 (N_6833,N_5387,N_4638);
nand U6834 (N_6834,N_5871,N_5380);
nor U6835 (N_6835,N_4721,N_5097);
nor U6836 (N_6836,N_5597,N_4761);
and U6837 (N_6837,N_5916,N_5290);
nor U6838 (N_6838,N_4598,N_5379);
and U6839 (N_6839,N_5108,N_4671);
xor U6840 (N_6840,N_5661,N_5738);
nand U6841 (N_6841,N_5296,N_5996);
and U6842 (N_6842,N_5114,N_4989);
nand U6843 (N_6843,N_5297,N_5159);
nor U6844 (N_6844,N_4700,N_5340);
or U6845 (N_6845,N_5680,N_5600);
and U6846 (N_6846,N_5591,N_5822);
nand U6847 (N_6847,N_4768,N_5175);
nand U6848 (N_6848,N_5777,N_5068);
nand U6849 (N_6849,N_4653,N_4913);
and U6850 (N_6850,N_5484,N_5386);
nand U6851 (N_6851,N_5171,N_5814);
and U6852 (N_6852,N_5525,N_5500);
nor U6853 (N_6853,N_5030,N_5690);
and U6854 (N_6854,N_5039,N_5558);
nor U6855 (N_6855,N_5315,N_5146);
nor U6856 (N_6856,N_5005,N_5726);
nor U6857 (N_6857,N_4921,N_5055);
and U6858 (N_6858,N_5537,N_4862);
and U6859 (N_6859,N_4989,N_5150);
nand U6860 (N_6860,N_5942,N_5482);
or U6861 (N_6861,N_5520,N_4674);
or U6862 (N_6862,N_5170,N_4854);
and U6863 (N_6863,N_5961,N_5507);
nor U6864 (N_6864,N_4895,N_4957);
and U6865 (N_6865,N_5945,N_4769);
nand U6866 (N_6866,N_5235,N_5779);
nor U6867 (N_6867,N_4727,N_5633);
and U6868 (N_6868,N_5068,N_4838);
or U6869 (N_6869,N_5096,N_4947);
nand U6870 (N_6870,N_5416,N_5910);
nor U6871 (N_6871,N_5405,N_4718);
and U6872 (N_6872,N_5717,N_5959);
or U6873 (N_6873,N_5324,N_5694);
nor U6874 (N_6874,N_5054,N_5953);
or U6875 (N_6875,N_5116,N_5731);
nand U6876 (N_6876,N_5285,N_5977);
nor U6877 (N_6877,N_5376,N_4829);
nor U6878 (N_6878,N_5328,N_5714);
or U6879 (N_6879,N_5240,N_5650);
and U6880 (N_6880,N_4821,N_5573);
nand U6881 (N_6881,N_5295,N_5692);
or U6882 (N_6882,N_4661,N_4743);
and U6883 (N_6883,N_5862,N_5607);
nor U6884 (N_6884,N_5763,N_5227);
or U6885 (N_6885,N_5071,N_5078);
and U6886 (N_6886,N_5411,N_5187);
nor U6887 (N_6887,N_5846,N_5762);
and U6888 (N_6888,N_4791,N_4582);
or U6889 (N_6889,N_4825,N_5858);
nand U6890 (N_6890,N_4734,N_4766);
or U6891 (N_6891,N_4642,N_5076);
or U6892 (N_6892,N_5955,N_4542);
and U6893 (N_6893,N_5083,N_5002);
and U6894 (N_6894,N_4864,N_5229);
nor U6895 (N_6895,N_5823,N_5732);
nand U6896 (N_6896,N_5296,N_4701);
or U6897 (N_6897,N_5946,N_5140);
nand U6898 (N_6898,N_4700,N_5043);
nor U6899 (N_6899,N_5488,N_4987);
and U6900 (N_6900,N_5053,N_5002);
nand U6901 (N_6901,N_4822,N_5627);
and U6902 (N_6902,N_5577,N_5782);
nand U6903 (N_6903,N_4729,N_5707);
nor U6904 (N_6904,N_5464,N_5161);
xnor U6905 (N_6905,N_5367,N_4721);
or U6906 (N_6906,N_4720,N_5697);
and U6907 (N_6907,N_5731,N_4507);
or U6908 (N_6908,N_5924,N_5959);
nand U6909 (N_6909,N_5717,N_5800);
and U6910 (N_6910,N_5286,N_4608);
nor U6911 (N_6911,N_5633,N_4896);
nand U6912 (N_6912,N_4672,N_4730);
nand U6913 (N_6913,N_5812,N_4771);
nor U6914 (N_6914,N_5334,N_5218);
or U6915 (N_6915,N_4781,N_5055);
nand U6916 (N_6916,N_4520,N_4699);
and U6917 (N_6917,N_5083,N_5055);
and U6918 (N_6918,N_5847,N_5474);
and U6919 (N_6919,N_5991,N_4658);
and U6920 (N_6920,N_4666,N_5987);
nor U6921 (N_6921,N_4544,N_5915);
nor U6922 (N_6922,N_4718,N_5519);
nor U6923 (N_6923,N_5851,N_5986);
or U6924 (N_6924,N_5885,N_4862);
nor U6925 (N_6925,N_4867,N_5872);
nor U6926 (N_6926,N_5699,N_5698);
nor U6927 (N_6927,N_5312,N_5948);
nor U6928 (N_6928,N_5700,N_4935);
nor U6929 (N_6929,N_4607,N_4714);
nor U6930 (N_6930,N_4895,N_4873);
nand U6931 (N_6931,N_4574,N_5632);
and U6932 (N_6932,N_4729,N_5540);
nor U6933 (N_6933,N_5621,N_4748);
or U6934 (N_6934,N_5294,N_5061);
nor U6935 (N_6935,N_5408,N_4586);
or U6936 (N_6936,N_5479,N_5317);
nand U6937 (N_6937,N_5346,N_4683);
or U6938 (N_6938,N_4790,N_5705);
and U6939 (N_6939,N_4801,N_4822);
or U6940 (N_6940,N_4509,N_4905);
and U6941 (N_6941,N_4614,N_5089);
nor U6942 (N_6942,N_5182,N_5846);
or U6943 (N_6943,N_5967,N_5489);
xor U6944 (N_6944,N_4795,N_4721);
nor U6945 (N_6945,N_5104,N_4889);
or U6946 (N_6946,N_5668,N_5638);
or U6947 (N_6947,N_4717,N_4838);
and U6948 (N_6948,N_5230,N_4881);
nor U6949 (N_6949,N_5073,N_5995);
or U6950 (N_6950,N_4910,N_4736);
and U6951 (N_6951,N_4710,N_4533);
or U6952 (N_6952,N_4850,N_5036);
and U6953 (N_6953,N_4985,N_4931);
and U6954 (N_6954,N_5668,N_5136);
or U6955 (N_6955,N_5945,N_5940);
and U6956 (N_6956,N_4545,N_5381);
nand U6957 (N_6957,N_5013,N_5407);
and U6958 (N_6958,N_5260,N_5100);
nand U6959 (N_6959,N_4545,N_5041);
nor U6960 (N_6960,N_5685,N_4544);
and U6961 (N_6961,N_5714,N_5651);
or U6962 (N_6962,N_5604,N_5388);
nand U6963 (N_6963,N_5375,N_4582);
nor U6964 (N_6964,N_5858,N_5431);
nor U6965 (N_6965,N_4857,N_4980);
nor U6966 (N_6966,N_4539,N_4765);
and U6967 (N_6967,N_5433,N_4562);
and U6968 (N_6968,N_5296,N_5465);
nor U6969 (N_6969,N_5364,N_5879);
nor U6970 (N_6970,N_5747,N_5099);
nand U6971 (N_6971,N_4508,N_5329);
nor U6972 (N_6972,N_5747,N_5214);
or U6973 (N_6973,N_5981,N_4932);
nand U6974 (N_6974,N_5318,N_5781);
nand U6975 (N_6975,N_5990,N_4700);
and U6976 (N_6976,N_4640,N_4678);
and U6977 (N_6977,N_4902,N_4648);
and U6978 (N_6978,N_5912,N_5109);
nand U6979 (N_6979,N_5722,N_4715);
and U6980 (N_6980,N_5592,N_5294);
nand U6981 (N_6981,N_5253,N_5747);
and U6982 (N_6982,N_5626,N_4924);
nand U6983 (N_6983,N_5846,N_4808);
nand U6984 (N_6984,N_4973,N_4953);
or U6985 (N_6985,N_5607,N_4906);
nor U6986 (N_6986,N_5444,N_4667);
or U6987 (N_6987,N_5995,N_5392);
or U6988 (N_6988,N_4990,N_5809);
nor U6989 (N_6989,N_4501,N_4624);
or U6990 (N_6990,N_5239,N_4850);
and U6991 (N_6991,N_5794,N_4996);
and U6992 (N_6992,N_5396,N_5966);
or U6993 (N_6993,N_4830,N_4572);
nand U6994 (N_6994,N_5264,N_5819);
nand U6995 (N_6995,N_4956,N_4707);
and U6996 (N_6996,N_5924,N_5509);
nor U6997 (N_6997,N_5494,N_5901);
or U6998 (N_6998,N_4716,N_5659);
or U6999 (N_6999,N_5128,N_5847);
nand U7000 (N_7000,N_5215,N_5697);
or U7001 (N_7001,N_4566,N_4506);
and U7002 (N_7002,N_5279,N_5250);
nand U7003 (N_7003,N_5737,N_4813);
or U7004 (N_7004,N_5754,N_4956);
nor U7005 (N_7005,N_5469,N_5504);
or U7006 (N_7006,N_5404,N_5275);
nor U7007 (N_7007,N_5688,N_5996);
and U7008 (N_7008,N_5701,N_5653);
or U7009 (N_7009,N_5335,N_5619);
nor U7010 (N_7010,N_5550,N_5460);
and U7011 (N_7011,N_5722,N_4858);
or U7012 (N_7012,N_5269,N_4828);
nor U7013 (N_7013,N_5476,N_5908);
nor U7014 (N_7014,N_5971,N_5679);
nand U7015 (N_7015,N_5929,N_5430);
or U7016 (N_7016,N_5736,N_5476);
or U7017 (N_7017,N_5087,N_4641);
nand U7018 (N_7018,N_5457,N_4793);
or U7019 (N_7019,N_5647,N_5548);
and U7020 (N_7020,N_4743,N_5552);
and U7021 (N_7021,N_5600,N_4620);
or U7022 (N_7022,N_5784,N_4511);
or U7023 (N_7023,N_4962,N_5410);
nor U7024 (N_7024,N_5627,N_5503);
nand U7025 (N_7025,N_4733,N_5902);
or U7026 (N_7026,N_4740,N_4985);
or U7027 (N_7027,N_4559,N_5963);
nand U7028 (N_7028,N_4877,N_5425);
and U7029 (N_7029,N_4617,N_5381);
nand U7030 (N_7030,N_5783,N_4772);
or U7031 (N_7031,N_5233,N_4837);
or U7032 (N_7032,N_4980,N_5291);
nor U7033 (N_7033,N_4865,N_4540);
or U7034 (N_7034,N_5742,N_5493);
or U7035 (N_7035,N_4748,N_4510);
or U7036 (N_7036,N_4600,N_5071);
and U7037 (N_7037,N_5631,N_5954);
nand U7038 (N_7038,N_4510,N_4667);
and U7039 (N_7039,N_5283,N_4608);
nand U7040 (N_7040,N_5454,N_4524);
nand U7041 (N_7041,N_5485,N_4693);
or U7042 (N_7042,N_5969,N_4643);
and U7043 (N_7043,N_5556,N_5591);
and U7044 (N_7044,N_5723,N_5797);
nand U7045 (N_7045,N_4783,N_4877);
nor U7046 (N_7046,N_5435,N_5932);
nand U7047 (N_7047,N_5690,N_5268);
nand U7048 (N_7048,N_5563,N_5253);
or U7049 (N_7049,N_4772,N_5253);
nor U7050 (N_7050,N_4523,N_4812);
and U7051 (N_7051,N_4953,N_5724);
or U7052 (N_7052,N_5545,N_4981);
or U7053 (N_7053,N_5217,N_5753);
and U7054 (N_7054,N_5239,N_5985);
nand U7055 (N_7055,N_5331,N_4556);
or U7056 (N_7056,N_5630,N_5062);
xor U7057 (N_7057,N_5207,N_4575);
xnor U7058 (N_7058,N_5398,N_4501);
or U7059 (N_7059,N_4679,N_5939);
nand U7060 (N_7060,N_5348,N_5890);
nand U7061 (N_7061,N_4645,N_5206);
nor U7062 (N_7062,N_5864,N_4615);
or U7063 (N_7063,N_5087,N_4825);
or U7064 (N_7064,N_5210,N_4979);
and U7065 (N_7065,N_4560,N_5807);
nand U7066 (N_7066,N_5316,N_4886);
nor U7067 (N_7067,N_5484,N_5409);
nand U7068 (N_7068,N_5412,N_5791);
nor U7069 (N_7069,N_5701,N_4943);
nand U7070 (N_7070,N_5383,N_5090);
or U7071 (N_7071,N_5807,N_4941);
nor U7072 (N_7072,N_5756,N_4897);
and U7073 (N_7073,N_5327,N_4869);
nand U7074 (N_7074,N_5377,N_4565);
and U7075 (N_7075,N_5947,N_4695);
or U7076 (N_7076,N_5583,N_5661);
or U7077 (N_7077,N_5422,N_5931);
or U7078 (N_7078,N_5451,N_5034);
or U7079 (N_7079,N_5164,N_4811);
nor U7080 (N_7080,N_5224,N_5327);
nand U7081 (N_7081,N_5301,N_5471);
nand U7082 (N_7082,N_5047,N_5984);
or U7083 (N_7083,N_4830,N_5996);
nand U7084 (N_7084,N_5596,N_5311);
or U7085 (N_7085,N_5725,N_5614);
and U7086 (N_7086,N_5450,N_4740);
nand U7087 (N_7087,N_5593,N_5311);
or U7088 (N_7088,N_4824,N_4649);
nor U7089 (N_7089,N_5677,N_4569);
nor U7090 (N_7090,N_5026,N_5538);
and U7091 (N_7091,N_5300,N_5765);
nand U7092 (N_7092,N_4596,N_4576);
nand U7093 (N_7093,N_5032,N_4513);
or U7094 (N_7094,N_4720,N_4938);
and U7095 (N_7095,N_5935,N_5151);
nor U7096 (N_7096,N_5773,N_5266);
nand U7097 (N_7097,N_4949,N_4722);
or U7098 (N_7098,N_5606,N_5746);
nor U7099 (N_7099,N_5069,N_5725);
and U7100 (N_7100,N_5092,N_5601);
nand U7101 (N_7101,N_5075,N_5356);
or U7102 (N_7102,N_4998,N_4721);
and U7103 (N_7103,N_5296,N_5212);
and U7104 (N_7104,N_5259,N_4579);
nor U7105 (N_7105,N_5928,N_4932);
or U7106 (N_7106,N_5987,N_4861);
nand U7107 (N_7107,N_5781,N_5286);
nand U7108 (N_7108,N_4994,N_5082);
nor U7109 (N_7109,N_5180,N_4974);
nor U7110 (N_7110,N_5313,N_5253);
nor U7111 (N_7111,N_4805,N_4631);
and U7112 (N_7112,N_5892,N_5901);
or U7113 (N_7113,N_5666,N_4698);
nand U7114 (N_7114,N_4968,N_4753);
nor U7115 (N_7115,N_5392,N_4836);
and U7116 (N_7116,N_5343,N_4576);
nor U7117 (N_7117,N_5775,N_4577);
or U7118 (N_7118,N_4886,N_5752);
nor U7119 (N_7119,N_4811,N_5839);
or U7120 (N_7120,N_4985,N_5289);
or U7121 (N_7121,N_4757,N_5893);
nand U7122 (N_7122,N_5025,N_5857);
or U7123 (N_7123,N_4891,N_5928);
and U7124 (N_7124,N_5704,N_5005);
nor U7125 (N_7125,N_4738,N_4537);
nand U7126 (N_7126,N_5029,N_5859);
and U7127 (N_7127,N_5939,N_5091);
or U7128 (N_7128,N_5344,N_4531);
xnor U7129 (N_7129,N_4639,N_4892);
and U7130 (N_7130,N_5564,N_4811);
or U7131 (N_7131,N_5017,N_4923);
or U7132 (N_7132,N_5032,N_4996);
and U7133 (N_7133,N_5946,N_4503);
nand U7134 (N_7134,N_5211,N_4704);
nor U7135 (N_7135,N_4718,N_4635);
or U7136 (N_7136,N_5759,N_5669);
and U7137 (N_7137,N_4932,N_5908);
or U7138 (N_7138,N_5507,N_5900);
nor U7139 (N_7139,N_4842,N_5084);
nor U7140 (N_7140,N_4583,N_5033);
or U7141 (N_7141,N_5110,N_4761);
and U7142 (N_7142,N_5164,N_5131);
and U7143 (N_7143,N_5213,N_4776);
or U7144 (N_7144,N_5287,N_4742);
or U7145 (N_7145,N_5585,N_5916);
or U7146 (N_7146,N_5613,N_5502);
nor U7147 (N_7147,N_5041,N_5028);
nor U7148 (N_7148,N_5502,N_5164);
and U7149 (N_7149,N_5179,N_5593);
nand U7150 (N_7150,N_5481,N_4532);
or U7151 (N_7151,N_4514,N_5657);
and U7152 (N_7152,N_5301,N_4666);
or U7153 (N_7153,N_4529,N_5169);
and U7154 (N_7154,N_4582,N_5728);
and U7155 (N_7155,N_4827,N_4996);
or U7156 (N_7156,N_4694,N_5808);
or U7157 (N_7157,N_4710,N_5779);
nand U7158 (N_7158,N_5533,N_4630);
nor U7159 (N_7159,N_5653,N_5707);
nand U7160 (N_7160,N_5785,N_4532);
or U7161 (N_7161,N_5719,N_5670);
nor U7162 (N_7162,N_5716,N_4564);
and U7163 (N_7163,N_5455,N_5777);
or U7164 (N_7164,N_5026,N_5994);
nand U7165 (N_7165,N_5107,N_5965);
or U7166 (N_7166,N_5762,N_5283);
and U7167 (N_7167,N_5312,N_5586);
or U7168 (N_7168,N_4620,N_5582);
or U7169 (N_7169,N_5949,N_5569);
nand U7170 (N_7170,N_5497,N_4828);
nor U7171 (N_7171,N_5187,N_4985);
or U7172 (N_7172,N_5338,N_5665);
nor U7173 (N_7173,N_4899,N_5331);
nor U7174 (N_7174,N_4816,N_5112);
xor U7175 (N_7175,N_5954,N_5822);
nor U7176 (N_7176,N_5963,N_4858);
nor U7177 (N_7177,N_4931,N_5047);
nand U7178 (N_7178,N_4854,N_5973);
xor U7179 (N_7179,N_5047,N_4755);
nor U7180 (N_7180,N_5768,N_5838);
or U7181 (N_7181,N_4844,N_5671);
or U7182 (N_7182,N_5910,N_4584);
and U7183 (N_7183,N_5102,N_5462);
nand U7184 (N_7184,N_5238,N_5134);
nand U7185 (N_7185,N_5640,N_4836);
nor U7186 (N_7186,N_5969,N_5385);
and U7187 (N_7187,N_5007,N_5305);
or U7188 (N_7188,N_5139,N_5552);
nand U7189 (N_7189,N_4599,N_4845);
and U7190 (N_7190,N_5802,N_5697);
nand U7191 (N_7191,N_4947,N_4622);
or U7192 (N_7192,N_4836,N_4968);
or U7193 (N_7193,N_5974,N_5339);
nand U7194 (N_7194,N_5791,N_5691);
or U7195 (N_7195,N_4693,N_5189);
nand U7196 (N_7196,N_4928,N_5699);
and U7197 (N_7197,N_5383,N_5095);
and U7198 (N_7198,N_5448,N_5207);
or U7199 (N_7199,N_4502,N_5827);
or U7200 (N_7200,N_5609,N_4953);
or U7201 (N_7201,N_5195,N_4888);
nand U7202 (N_7202,N_4601,N_5002);
and U7203 (N_7203,N_4502,N_5465);
and U7204 (N_7204,N_5376,N_4746);
and U7205 (N_7205,N_5935,N_5248);
and U7206 (N_7206,N_4876,N_4546);
nand U7207 (N_7207,N_5537,N_4636);
nor U7208 (N_7208,N_5989,N_5104);
nor U7209 (N_7209,N_4648,N_5391);
or U7210 (N_7210,N_5415,N_5907);
nor U7211 (N_7211,N_4898,N_5191);
or U7212 (N_7212,N_5287,N_4812);
nor U7213 (N_7213,N_5958,N_5252);
or U7214 (N_7214,N_5149,N_5577);
nand U7215 (N_7215,N_4620,N_4933);
nor U7216 (N_7216,N_5822,N_5950);
or U7217 (N_7217,N_5318,N_5843);
and U7218 (N_7218,N_5991,N_5072);
or U7219 (N_7219,N_5821,N_4812);
and U7220 (N_7220,N_5237,N_5731);
nand U7221 (N_7221,N_5617,N_4826);
nand U7222 (N_7222,N_5358,N_5023);
nor U7223 (N_7223,N_5282,N_4793);
nor U7224 (N_7224,N_5751,N_4920);
and U7225 (N_7225,N_4513,N_4967);
nand U7226 (N_7226,N_5877,N_4606);
or U7227 (N_7227,N_5803,N_4849);
and U7228 (N_7228,N_5704,N_4870);
or U7229 (N_7229,N_4799,N_5400);
nor U7230 (N_7230,N_5696,N_4584);
nand U7231 (N_7231,N_4664,N_4765);
nand U7232 (N_7232,N_4608,N_4849);
and U7233 (N_7233,N_4720,N_4768);
and U7234 (N_7234,N_5674,N_5159);
or U7235 (N_7235,N_5859,N_4777);
nand U7236 (N_7236,N_5685,N_5528);
nand U7237 (N_7237,N_5780,N_5849);
nor U7238 (N_7238,N_5099,N_5307);
nor U7239 (N_7239,N_5677,N_5433);
and U7240 (N_7240,N_4583,N_4762);
nand U7241 (N_7241,N_5272,N_5153);
nor U7242 (N_7242,N_4531,N_4879);
nand U7243 (N_7243,N_4584,N_4587);
nor U7244 (N_7244,N_5255,N_4739);
and U7245 (N_7245,N_5394,N_5353);
nor U7246 (N_7246,N_4664,N_5364);
nand U7247 (N_7247,N_5543,N_5295);
and U7248 (N_7248,N_5712,N_5867);
and U7249 (N_7249,N_5515,N_5313);
and U7250 (N_7250,N_4697,N_5738);
nand U7251 (N_7251,N_5671,N_5707);
nor U7252 (N_7252,N_4501,N_5114);
and U7253 (N_7253,N_5204,N_5914);
or U7254 (N_7254,N_5255,N_5692);
or U7255 (N_7255,N_4804,N_5913);
and U7256 (N_7256,N_5438,N_5946);
and U7257 (N_7257,N_4781,N_5068);
nor U7258 (N_7258,N_4603,N_5722);
and U7259 (N_7259,N_5131,N_4919);
nand U7260 (N_7260,N_4918,N_5827);
nor U7261 (N_7261,N_5339,N_5448);
and U7262 (N_7262,N_5428,N_4701);
nand U7263 (N_7263,N_5431,N_5213);
or U7264 (N_7264,N_4957,N_5457);
nand U7265 (N_7265,N_5553,N_5386);
nand U7266 (N_7266,N_5667,N_4830);
nand U7267 (N_7267,N_4734,N_5836);
nor U7268 (N_7268,N_5790,N_4866);
nor U7269 (N_7269,N_5462,N_5040);
nand U7270 (N_7270,N_4670,N_5135);
and U7271 (N_7271,N_4948,N_5950);
and U7272 (N_7272,N_4568,N_5865);
and U7273 (N_7273,N_4898,N_5667);
nand U7274 (N_7274,N_4577,N_5704);
nand U7275 (N_7275,N_4773,N_4501);
or U7276 (N_7276,N_4751,N_5451);
or U7277 (N_7277,N_4918,N_4938);
and U7278 (N_7278,N_4555,N_5039);
or U7279 (N_7279,N_5723,N_5435);
xnor U7280 (N_7280,N_4622,N_5906);
or U7281 (N_7281,N_4687,N_4718);
or U7282 (N_7282,N_4926,N_5992);
nor U7283 (N_7283,N_5723,N_5841);
nand U7284 (N_7284,N_5631,N_5447);
or U7285 (N_7285,N_5730,N_4861);
nand U7286 (N_7286,N_4570,N_5990);
and U7287 (N_7287,N_5597,N_5536);
nand U7288 (N_7288,N_5683,N_5647);
nand U7289 (N_7289,N_5356,N_5050);
nand U7290 (N_7290,N_4657,N_5024);
nor U7291 (N_7291,N_5304,N_5517);
nand U7292 (N_7292,N_4988,N_5942);
nor U7293 (N_7293,N_5253,N_4798);
and U7294 (N_7294,N_5450,N_5896);
or U7295 (N_7295,N_5547,N_5463);
and U7296 (N_7296,N_4786,N_5196);
nand U7297 (N_7297,N_4605,N_5104);
nor U7298 (N_7298,N_5766,N_5656);
nand U7299 (N_7299,N_5957,N_5646);
and U7300 (N_7300,N_5855,N_5258);
nand U7301 (N_7301,N_5280,N_5796);
nand U7302 (N_7302,N_4798,N_5855);
and U7303 (N_7303,N_5977,N_5508);
nand U7304 (N_7304,N_5908,N_5996);
or U7305 (N_7305,N_5607,N_4954);
and U7306 (N_7306,N_4810,N_4614);
or U7307 (N_7307,N_5859,N_5176);
nand U7308 (N_7308,N_5065,N_5205);
nor U7309 (N_7309,N_5192,N_4852);
nor U7310 (N_7310,N_5474,N_5389);
or U7311 (N_7311,N_5367,N_5206);
or U7312 (N_7312,N_5953,N_4616);
or U7313 (N_7313,N_4732,N_5380);
nor U7314 (N_7314,N_5837,N_4969);
nand U7315 (N_7315,N_5846,N_5868);
nand U7316 (N_7316,N_4976,N_5568);
and U7317 (N_7317,N_5777,N_5930);
nand U7318 (N_7318,N_5472,N_5464);
nand U7319 (N_7319,N_5194,N_4717);
nand U7320 (N_7320,N_5020,N_5805);
or U7321 (N_7321,N_4580,N_4597);
nand U7322 (N_7322,N_5716,N_5336);
and U7323 (N_7323,N_5947,N_5662);
or U7324 (N_7324,N_5428,N_5450);
and U7325 (N_7325,N_4806,N_4945);
nand U7326 (N_7326,N_4991,N_5300);
or U7327 (N_7327,N_5385,N_5104);
and U7328 (N_7328,N_5396,N_5711);
xnor U7329 (N_7329,N_4821,N_5633);
nand U7330 (N_7330,N_5097,N_5155);
or U7331 (N_7331,N_4744,N_4623);
xor U7332 (N_7332,N_5532,N_5976);
nand U7333 (N_7333,N_5531,N_5951);
and U7334 (N_7334,N_5627,N_5072);
and U7335 (N_7335,N_5537,N_5348);
and U7336 (N_7336,N_5221,N_4537);
nand U7337 (N_7337,N_5012,N_5551);
and U7338 (N_7338,N_5907,N_5617);
nor U7339 (N_7339,N_4910,N_5454);
nand U7340 (N_7340,N_5549,N_5234);
or U7341 (N_7341,N_5858,N_5220);
nand U7342 (N_7342,N_5456,N_5117);
nor U7343 (N_7343,N_5264,N_5467);
and U7344 (N_7344,N_4676,N_4991);
or U7345 (N_7345,N_4998,N_5549);
and U7346 (N_7346,N_5301,N_4968);
or U7347 (N_7347,N_5536,N_4882);
nand U7348 (N_7348,N_4972,N_5426);
and U7349 (N_7349,N_5632,N_5971);
nor U7350 (N_7350,N_5503,N_5931);
or U7351 (N_7351,N_4782,N_4837);
nor U7352 (N_7352,N_4837,N_5533);
and U7353 (N_7353,N_4745,N_5275);
nor U7354 (N_7354,N_5061,N_4734);
and U7355 (N_7355,N_5194,N_5213);
nor U7356 (N_7356,N_5823,N_5081);
and U7357 (N_7357,N_5423,N_5408);
or U7358 (N_7358,N_5042,N_5027);
and U7359 (N_7359,N_5512,N_4960);
or U7360 (N_7360,N_5304,N_4653);
and U7361 (N_7361,N_4943,N_5939);
nand U7362 (N_7362,N_4744,N_5123);
nand U7363 (N_7363,N_4629,N_5142);
nor U7364 (N_7364,N_5286,N_5738);
nor U7365 (N_7365,N_5586,N_4739);
nor U7366 (N_7366,N_5496,N_4765);
or U7367 (N_7367,N_5559,N_5548);
or U7368 (N_7368,N_4926,N_5372);
or U7369 (N_7369,N_4745,N_5900);
nand U7370 (N_7370,N_5740,N_5783);
nand U7371 (N_7371,N_5181,N_5250);
nor U7372 (N_7372,N_5088,N_5200);
and U7373 (N_7373,N_4852,N_5643);
nand U7374 (N_7374,N_4844,N_4865);
nand U7375 (N_7375,N_5843,N_5448);
nand U7376 (N_7376,N_5823,N_5411);
xnor U7377 (N_7377,N_5338,N_5983);
nor U7378 (N_7378,N_5381,N_5345);
nand U7379 (N_7379,N_5123,N_5927);
nor U7380 (N_7380,N_5019,N_4735);
and U7381 (N_7381,N_5785,N_5787);
and U7382 (N_7382,N_5646,N_4854);
nor U7383 (N_7383,N_4763,N_4520);
and U7384 (N_7384,N_5640,N_5511);
nor U7385 (N_7385,N_4894,N_5870);
nor U7386 (N_7386,N_5469,N_5064);
nor U7387 (N_7387,N_5757,N_5195);
nand U7388 (N_7388,N_4658,N_4562);
nand U7389 (N_7389,N_4881,N_4873);
and U7390 (N_7390,N_4745,N_4513);
and U7391 (N_7391,N_5238,N_5213);
or U7392 (N_7392,N_5499,N_5358);
nand U7393 (N_7393,N_5143,N_4965);
xor U7394 (N_7394,N_5338,N_4834);
nor U7395 (N_7395,N_4551,N_4541);
and U7396 (N_7396,N_4576,N_5835);
nor U7397 (N_7397,N_4556,N_4562);
or U7398 (N_7398,N_4546,N_5654);
nand U7399 (N_7399,N_5236,N_4965);
nor U7400 (N_7400,N_5849,N_5152);
and U7401 (N_7401,N_4727,N_5073);
nand U7402 (N_7402,N_5838,N_5484);
nand U7403 (N_7403,N_5362,N_4883);
and U7404 (N_7404,N_5046,N_5251);
and U7405 (N_7405,N_5189,N_5521);
nand U7406 (N_7406,N_5400,N_5707);
nor U7407 (N_7407,N_5589,N_4595);
nand U7408 (N_7408,N_4652,N_4858);
and U7409 (N_7409,N_5628,N_5650);
and U7410 (N_7410,N_5138,N_4774);
or U7411 (N_7411,N_5134,N_5027);
nand U7412 (N_7412,N_4703,N_5684);
nor U7413 (N_7413,N_4790,N_5105);
or U7414 (N_7414,N_5617,N_4797);
and U7415 (N_7415,N_5314,N_4671);
nand U7416 (N_7416,N_5041,N_4534);
nor U7417 (N_7417,N_4562,N_4542);
or U7418 (N_7418,N_4780,N_4785);
and U7419 (N_7419,N_4539,N_5147);
and U7420 (N_7420,N_5696,N_5318);
nor U7421 (N_7421,N_5176,N_5689);
nor U7422 (N_7422,N_5661,N_5072);
or U7423 (N_7423,N_4749,N_5486);
nand U7424 (N_7424,N_5569,N_4770);
or U7425 (N_7425,N_5431,N_5785);
or U7426 (N_7426,N_5135,N_5854);
nand U7427 (N_7427,N_4544,N_4549);
and U7428 (N_7428,N_5486,N_4849);
nand U7429 (N_7429,N_5628,N_4958);
and U7430 (N_7430,N_4570,N_5950);
nor U7431 (N_7431,N_5436,N_5870);
or U7432 (N_7432,N_4729,N_5053);
or U7433 (N_7433,N_4954,N_4661);
or U7434 (N_7434,N_5109,N_4578);
and U7435 (N_7435,N_5093,N_5974);
nor U7436 (N_7436,N_5547,N_5998);
and U7437 (N_7437,N_5527,N_5117);
nor U7438 (N_7438,N_5541,N_5602);
nor U7439 (N_7439,N_4611,N_5492);
nand U7440 (N_7440,N_4553,N_4528);
nor U7441 (N_7441,N_5574,N_5588);
and U7442 (N_7442,N_5091,N_4549);
nor U7443 (N_7443,N_4667,N_5469);
and U7444 (N_7444,N_4975,N_5265);
nor U7445 (N_7445,N_5027,N_5715);
nand U7446 (N_7446,N_5721,N_5574);
or U7447 (N_7447,N_5098,N_4848);
and U7448 (N_7448,N_5659,N_4517);
and U7449 (N_7449,N_5800,N_5473);
nand U7450 (N_7450,N_5024,N_5689);
nor U7451 (N_7451,N_5973,N_4605);
or U7452 (N_7452,N_5092,N_4503);
and U7453 (N_7453,N_5596,N_5838);
or U7454 (N_7454,N_5840,N_5429);
and U7455 (N_7455,N_5270,N_5708);
or U7456 (N_7456,N_5369,N_4722);
nand U7457 (N_7457,N_4919,N_5142);
or U7458 (N_7458,N_5259,N_4539);
and U7459 (N_7459,N_5777,N_4640);
nand U7460 (N_7460,N_5720,N_5318);
and U7461 (N_7461,N_5061,N_4755);
nand U7462 (N_7462,N_4855,N_4768);
nand U7463 (N_7463,N_5642,N_5465);
or U7464 (N_7464,N_5931,N_4639);
nor U7465 (N_7465,N_5947,N_5723);
and U7466 (N_7466,N_4734,N_5876);
or U7467 (N_7467,N_5842,N_4997);
nor U7468 (N_7468,N_5649,N_4924);
or U7469 (N_7469,N_4704,N_4502);
or U7470 (N_7470,N_5910,N_4765);
and U7471 (N_7471,N_4652,N_5512);
nand U7472 (N_7472,N_4844,N_4714);
or U7473 (N_7473,N_5511,N_5469);
or U7474 (N_7474,N_4809,N_4693);
and U7475 (N_7475,N_5864,N_5941);
nand U7476 (N_7476,N_4605,N_5514);
nor U7477 (N_7477,N_5852,N_5551);
and U7478 (N_7478,N_4782,N_4517);
nand U7479 (N_7479,N_4797,N_4666);
or U7480 (N_7480,N_5782,N_5870);
and U7481 (N_7481,N_5563,N_5949);
nor U7482 (N_7482,N_4798,N_4748);
and U7483 (N_7483,N_4785,N_5420);
nor U7484 (N_7484,N_4969,N_5129);
nand U7485 (N_7485,N_5768,N_4840);
nand U7486 (N_7486,N_4685,N_5608);
nor U7487 (N_7487,N_5379,N_4626);
nand U7488 (N_7488,N_4930,N_4837);
and U7489 (N_7489,N_5693,N_4587);
and U7490 (N_7490,N_5756,N_4712);
or U7491 (N_7491,N_5943,N_5313);
or U7492 (N_7492,N_5511,N_5785);
nor U7493 (N_7493,N_4618,N_5065);
nand U7494 (N_7494,N_5212,N_5356);
nand U7495 (N_7495,N_5354,N_4744);
nand U7496 (N_7496,N_4976,N_4941);
nand U7497 (N_7497,N_5778,N_5143);
or U7498 (N_7498,N_4620,N_5479);
and U7499 (N_7499,N_5748,N_4979);
and U7500 (N_7500,N_7429,N_7305);
and U7501 (N_7501,N_6479,N_6812);
nand U7502 (N_7502,N_6393,N_7184);
and U7503 (N_7503,N_6966,N_7078);
nand U7504 (N_7504,N_6662,N_7232);
nor U7505 (N_7505,N_6496,N_6001);
nor U7506 (N_7506,N_6108,N_6971);
or U7507 (N_7507,N_7027,N_6984);
nor U7508 (N_7508,N_6699,N_7371);
nand U7509 (N_7509,N_7032,N_6989);
and U7510 (N_7510,N_7056,N_6463);
nand U7511 (N_7511,N_6953,N_7460);
nand U7512 (N_7512,N_6171,N_6593);
nor U7513 (N_7513,N_6738,N_6180);
or U7514 (N_7514,N_6586,N_7143);
nand U7515 (N_7515,N_7196,N_6655);
and U7516 (N_7516,N_6865,N_6977);
and U7517 (N_7517,N_6383,N_7492);
nand U7518 (N_7518,N_6147,N_6248);
nand U7519 (N_7519,N_6945,N_6684);
nor U7520 (N_7520,N_6567,N_6535);
and U7521 (N_7521,N_6735,N_6657);
nor U7522 (N_7522,N_6163,N_7077);
and U7523 (N_7523,N_6194,N_7281);
nand U7524 (N_7524,N_6722,N_7046);
nor U7525 (N_7525,N_6247,N_6770);
and U7526 (N_7526,N_7261,N_7259);
nand U7527 (N_7527,N_7158,N_6161);
nand U7528 (N_7528,N_6861,N_6588);
nand U7529 (N_7529,N_6183,N_6753);
nor U7530 (N_7530,N_6355,N_6771);
or U7531 (N_7531,N_7308,N_7242);
nand U7532 (N_7532,N_7166,N_7226);
nor U7533 (N_7533,N_6538,N_6294);
and U7534 (N_7534,N_6307,N_6358);
nor U7535 (N_7535,N_6271,N_6300);
and U7536 (N_7536,N_6200,N_7432);
or U7537 (N_7537,N_6202,N_6299);
or U7538 (N_7538,N_7381,N_7187);
nor U7539 (N_7539,N_7017,N_6086);
nand U7540 (N_7540,N_6042,N_6846);
nor U7541 (N_7541,N_6095,N_7491);
nand U7542 (N_7542,N_6745,N_6159);
and U7543 (N_7543,N_6851,N_7446);
or U7544 (N_7544,N_6497,N_7055);
nand U7545 (N_7545,N_7193,N_7401);
xor U7546 (N_7546,N_6533,N_7263);
and U7547 (N_7547,N_6033,N_6808);
or U7548 (N_7548,N_7434,N_6581);
and U7549 (N_7549,N_7202,N_6352);
nand U7550 (N_7550,N_6346,N_6616);
nor U7551 (N_7551,N_6956,N_7477);
or U7552 (N_7552,N_6893,N_6103);
nand U7553 (N_7553,N_6158,N_7102);
and U7554 (N_7554,N_7262,N_7181);
nor U7555 (N_7555,N_7011,N_7339);
nor U7556 (N_7556,N_6118,N_6900);
nand U7557 (N_7557,N_7264,N_6908);
nand U7558 (N_7558,N_6372,N_6857);
nand U7559 (N_7559,N_6020,N_6281);
nor U7560 (N_7560,N_6913,N_6709);
xor U7561 (N_7561,N_6316,N_6816);
and U7562 (N_7562,N_6916,N_7209);
nand U7563 (N_7563,N_6006,N_6119);
and U7564 (N_7564,N_6007,N_7274);
or U7565 (N_7565,N_6345,N_6363);
nor U7566 (N_7566,N_7229,N_7285);
nor U7567 (N_7567,N_7349,N_6492);
or U7568 (N_7568,N_6727,N_6650);
or U7569 (N_7569,N_6637,N_7178);
nand U7570 (N_7570,N_7185,N_7215);
nor U7571 (N_7571,N_6458,N_6004);
nor U7572 (N_7572,N_6031,N_6870);
nand U7573 (N_7573,N_7214,N_7223);
and U7574 (N_7574,N_7266,N_6721);
or U7575 (N_7575,N_6211,N_6029);
or U7576 (N_7576,N_6388,N_7064);
nor U7577 (N_7577,N_7130,N_7124);
nor U7578 (N_7578,N_6573,N_7085);
and U7579 (N_7579,N_6380,N_6368);
nor U7580 (N_7580,N_6754,N_6992);
and U7581 (N_7581,N_6157,N_7246);
or U7582 (N_7582,N_6401,N_6071);
xnor U7583 (N_7583,N_7065,N_7071);
nand U7584 (N_7584,N_6451,N_6400);
nor U7585 (N_7585,N_6545,N_6057);
nor U7586 (N_7586,N_6547,N_6472);
nand U7587 (N_7587,N_6235,N_7438);
nand U7588 (N_7588,N_7272,N_6610);
or U7589 (N_7589,N_6072,N_7174);
nand U7590 (N_7590,N_6841,N_7092);
nor U7591 (N_7591,N_6192,N_6566);
nand U7592 (N_7592,N_7475,N_7292);
and U7593 (N_7593,N_7177,N_7362);
nor U7594 (N_7594,N_7467,N_6671);
nand U7595 (N_7595,N_6903,N_6416);
and U7596 (N_7596,N_6540,N_7322);
nor U7597 (N_7597,N_6392,N_6452);
nor U7598 (N_7598,N_7424,N_6078);
and U7599 (N_7599,N_6634,N_6667);
or U7600 (N_7600,N_7353,N_7219);
and U7601 (N_7601,N_6933,N_6359);
nand U7602 (N_7602,N_7313,N_6606);
nor U7603 (N_7603,N_6411,N_6869);
and U7604 (N_7604,N_7099,N_6319);
nand U7605 (N_7605,N_6246,N_7470);
or U7606 (N_7606,N_6322,N_6844);
and U7607 (N_7607,N_7109,N_7089);
nand U7608 (N_7608,N_6925,N_7142);
and U7609 (N_7609,N_6189,N_7410);
nand U7610 (N_7610,N_6850,N_6543);
or U7611 (N_7611,N_6744,N_6982);
nand U7612 (N_7612,N_7128,N_7405);
and U7613 (N_7613,N_6466,N_7194);
and U7614 (N_7614,N_7041,N_6898);
nand U7615 (N_7615,N_6418,N_6026);
xnor U7616 (N_7616,N_6414,N_7180);
and U7617 (N_7617,N_6115,N_6750);
and U7618 (N_7618,N_6424,N_7135);
nand U7619 (N_7619,N_6387,N_7016);
nand U7620 (N_7620,N_6509,N_7358);
nor U7621 (N_7621,N_6384,N_6758);
nor U7622 (N_7622,N_7039,N_6914);
or U7623 (N_7623,N_6652,N_6876);
and U7624 (N_7624,N_6120,N_6341);
and U7625 (N_7625,N_7478,N_7307);
and U7626 (N_7626,N_6325,N_7275);
nor U7627 (N_7627,N_7412,N_7076);
and U7628 (N_7628,N_6499,N_6902);
or U7629 (N_7629,N_7472,N_6223);
and U7630 (N_7630,N_7463,N_6923);
or U7631 (N_7631,N_6921,N_6131);
and U7632 (N_7632,N_7002,N_7427);
nor U7633 (N_7633,N_7101,N_7119);
nor U7634 (N_7634,N_6886,N_6105);
nand U7635 (N_7635,N_6045,N_7456);
or U7636 (N_7636,N_6934,N_7356);
nand U7637 (N_7637,N_6556,N_6153);
nand U7638 (N_7638,N_6531,N_6706);
nand U7639 (N_7639,N_7377,N_7132);
nor U7640 (N_7640,N_6892,N_6884);
or U7641 (N_7641,N_7160,N_6952);
and U7642 (N_7642,N_7114,N_7311);
nor U7643 (N_7643,N_6824,N_7058);
nor U7644 (N_7644,N_7480,N_6685);
or U7645 (N_7645,N_6469,N_7398);
or U7646 (N_7646,N_6944,N_6516);
nor U7647 (N_7647,N_6257,N_7100);
nor U7648 (N_7648,N_7172,N_6594);
nor U7649 (N_7649,N_6752,N_6957);
and U7650 (N_7650,N_6795,N_7498);
or U7651 (N_7651,N_6802,N_6085);
or U7652 (N_7652,N_6951,N_6522);
or U7653 (N_7653,N_7222,N_7473);
or U7654 (N_7654,N_6204,N_7073);
and U7655 (N_7655,N_7332,N_6833);
nand U7656 (N_7656,N_7331,N_7328);
nor U7657 (N_7657,N_7413,N_6421);
nand U7658 (N_7658,N_6048,N_6948);
nor U7659 (N_7659,N_6149,N_6700);
and U7660 (N_7660,N_6324,N_6236);
or U7661 (N_7661,N_7437,N_7125);
and U7662 (N_7662,N_7448,N_7452);
or U7663 (N_7663,N_6590,N_6631);
nand U7664 (N_7664,N_6651,N_6602);
nor U7665 (N_7665,N_6162,N_7117);
and U7666 (N_7666,N_6170,N_7228);
and U7667 (N_7667,N_6221,N_6151);
and U7668 (N_7668,N_7428,N_7403);
nor U7669 (N_7669,N_7159,N_6726);
nand U7670 (N_7670,N_6612,N_6690);
or U7671 (N_7671,N_6768,N_6036);
nand U7672 (N_7672,N_6224,N_6417);
or U7673 (N_7673,N_6014,N_6798);
and U7674 (N_7674,N_6676,N_6043);
nand U7675 (N_7675,N_7249,N_6765);
nand U7676 (N_7676,N_6058,N_6051);
nor U7677 (N_7677,N_7097,N_7203);
or U7678 (N_7678,N_6222,N_6284);
nand U7679 (N_7679,N_6068,N_6260);
nor U7680 (N_7680,N_6361,N_7454);
or U7681 (N_7681,N_6818,N_7256);
or U7682 (N_7682,N_6308,N_6412);
nor U7683 (N_7683,N_6261,N_7208);
nand U7684 (N_7684,N_6932,N_6691);
or U7685 (N_7685,N_6664,N_7442);
nor U7686 (N_7686,N_6199,N_6196);
or U7687 (N_7687,N_6054,N_6137);
or U7688 (N_7688,N_6461,N_6258);
and U7689 (N_7689,N_6680,N_7450);
and U7690 (N_7690,N_6350,N_6519);
nand U7691 (N_7691,N_7451,N_6521);
nand U7692 (N_7692,N_7207,N_6460);
and U7693 (N_7693,N_6832,N_6658);
nor U7694 (N_7694,N_7306,N_7050);
nor U7695 (N_7695,N_7350,N_6367);
and U7696 (N_7696,N_6471,N_7329);
or U7697 (N_7697,N_6836,N_6369);
nor U7698 (N_7698,N_6339,N_7360);
nor U7699 (N_7699,N_6641,N_7149);
nor U7700 (N_7700,N_6974,N_6599);
or U7701 (N_7701,N_6114,N_7230);
nand U7702 (N_7702,N_7344,N_6696);
nand U7703 (N_7703,N_6090,N_7170);
or U7704 (N_7704,N_6807,N_6840);
and U7705 (N_7705,N_6872,N_6629);
nor U7706 (N_7706,N_7265,N_7171);
nand U7707 (N_7707,N_6182,N_7009);
nor U7708 (N_7708,N_6973,N_7310);
or U7709 (N_7709,N_6077,N_7147);
nor U7710 (N_7710,N_6897,N_7420);
or U7711 (N_7711,N_6267,N_6589);
and U7712 (N_7712,N_6666,N_6734);
nand U7713 (N_7713,N_7024,N_6644);
nor U7714 (N_7714,N_7019,N_7186);
and U7715 (N_7715,N_7459,N_7043);
or U7716 (N_7716,N_6191,N_7048);
or U7717 (N_7717,N_6718,N_6785);
nand U7718 (N_7718,N_6856,N_6373);
nand U7719 (N_7719,N_7270,N_6291);
or U7720 (N_7720,N_6433,N_6164);
nand U7721 (N_7721,N_6990,N_6927);
and U7722 (N_7722,N_7237,N_6817);
nand U7723 (N_7723,N_6789,N_6849);
and U7724 (N_7724,N_7443,N_7179);
nor U7725 (N_7725,N_6842,N_7378);
nand U7726 (N_7726,N_7372,N_6292);
nor U7727 (N_7727,N_7040,N_6148);
nand U7728 (N_7728,N_6866,N_6782);
nand U7729 (N_7729,N_6862,N_6140);
nor U7730 (N_7730,N_6428,N_7200);
nand U7731 (N_7731,N_7031,N_6225);
and U7732 (N_7732,N_7425,N_7444);
nand U7733 (N_7733,N_7391,N_6883);
nand U7734 (N_7734,N_7131,N_7284);
nor U7735 (N_7735,N_6498,N_7494);
and U7736 (N_7736,N_6524,N_6129);
nand U7737 (N_7737,N_6265,N_6595);
nor U7738 (N_7738,N_7008,N_7062);
nor U7739 (N_7739,N_7038,N_6623);
nor U7740 (N_7740,N_7144,N_7188);
or U7741 (N_7741,N_6582,N_7318);
or U7742 (N_7742,N_6541,N_7216);
or U7743 (N_7743,N_6490,N_6038);
xor U7744 (N_7744,N_6126,N_6829);
or U7745 (N_7745,N_7258,N_6733);
and U7746 (N_7746,N_6512,N_6141);
and U7747 (N_7747,N_6441,N_6574);
nand U7748 (N_7748,N_6993,N_7396);
or U7749 (N_7749,N_7383,N_7288);
and U7750 (N_7750,N_6008,N_6987);
nand U7751 (N_7751,N_7397,N_6674);
nand U7752 (N_7752,N_6740,N_6776);
nand U7753 (N_7753,N_6122,N_7123);
nor U7754 (N_7754,N_6028,N_7118);
nand U7755 (N_7755,N_6178,N_7220);
nand U7756 (N_7756,N_6935,N_7049);
nor U7757 (N_7757,N_6213,N_6330);
nand U7758 (N_7758,N_7471,N_7212);
and U7759 (N_7759,N_6675,N_6943);
nand U7760 (N_7760,N_7431,N_6081);
or U7761 (N_7761,N_6475,N_6198);
nand U7762 (N_7762,N_6348,N_7022);
nand U7763 (N_7763,N_6124,N_6059);
and U7764 (N_7764,N_7485,N_7345);
and U7765 (N_7765,N_7000,N_6918);
and U7766 (N_7766,N_7340,N_6797);
nor U7767 (N_7767,N_6578,N_6473);
nand U7768 (N_7768,N_6751,N_6814);
nand U7769 (N_7769,N_7139,N_7302);
nand U7770 (N_7770,N_7441,N_7495);
and U7771 (N_7771,N_6985,N_6321);
or U7772 (N_7772,N_6929,N_6881);
nor U7773 (N_7773,N_7342,N_7445);
or U7774 (N_7774,N_6939,N_7369);
nand U7775 (N_7775,N_6130,N_6713);
nor U7776 (N_7776,N_6378,N_6167);
nor U7777 (N_7777,N_7301,N_7368);
and U7778 (N_7778,N_6701,N_6517);
nor U7779 (N_7779,N_6431,N_6591);
and U7780 (N_7780,N_6875,N_6649);
or U7781 (N_7781,N_6732,N_6229);
and U7782 (N_7782,N_6470,N_6710);
nand U7783 (N_7783,N_7376,N_6825);
and U7784 (N_7784,N_7324,N_6518);
and U7785 (N_7785,N_7387,N_7169);
or U7786 (N_7786,N_6160,N_6584);
nor U7787 (N_7787,N_6279,N_6988);
nor U7788 (N_7788,N_6962,N_6216);
nor U7789 (N_7789,N_6268,N_7030);
or U7790 (N_7790,N_7276,N_7476);
and U7791 (N_7791,N_6201,N_6207);
and U7792 (N_7792,N_7115,N_6653);
nand U7793 (N_7793,N_6370,N_7218);
or U7794 (N_7794,N_7148,N_6154);
nor U7795 (N_7795,N_7252,N_7462);
nand U7796 (N_7796,N_7210,N_6835);
nand U7797 (N_7797,N_6636,N_6080);
and U7798 (N_7798,N_6301,N_6603);
nand U7799 (N_7799,N_6000,N_6780);
nor U7800 (N_7800,N_6228,N_6289);
or U7801 (N_7801,N_7354,N_7379);
nor U7802 (N_7802,N_6572,N_7296);
or U7803 (N_7803,N_6293,N_6609);
or U7804 (N_7804,N_6273,N_6642);
nor U7805 (N_7805,N_6999,N_7217);
and U7806 (N_7806,N_6009,N_6082);
or U7807 (N_7807,N_6600,N_6430);
or U7808 (N_7808,N_7290,N_6374);
and U7809 (N_7809,N_6663,N_7298);
nor U7810 (N_7810,N_6190,N_6793);
nand U7811 (N_7811,N_6672,N_6855);
nand U7812 (N_7812,N_6834,N_6654);
nand U7813 (N_7813,N_7028,N_7074);
nor U7814 (N_7814,N_7173,N_6169);
xor U7815 (N_7815,N_7026,N_7493);
nand U7816 (N_7816,N_6117,N_6731);
nor U7817 (N_7817,N_7343,N_7094);
and U7818 (N_7818,N_6774,N_6544);
xor U7819 (N_7819,N_6262,N_6564);
or U7820 (N_7820,N_7294,N_7414);
or U7821 (N_7821,N_6027,N_6375);
nor U7822 (N_7822,N_6830,N_6422);
and U7823 (N_7823,N_7066,N_6963);
nor U7824 (N_7824,N_6483,N_6063);
or U7825 (N_7825,N_7394,N_6232);
or U7826 (N_7826,N_7162,N_6208);
and U7827 (N_7827,N_6764,N_6894);
nor U7828 (N_7828,N_6910,N_7183);
nor U7829 (N_7829,N_7090,N_6116);
or U7830 (N_7830,N_6739,N_6134);
nor U7831 (N_7831,N_6254,N_6579);
nor U7832 (N_7832,N_6349,N_6060);
nand U7833 (N_7833,N_6845,N_6410);
nand U7834 (N_7834,N_6156,N_6478);
nor U7835 (N_7835,N_7151,N_6702);
or U7836 (N_7836,N_6215,N_6557);
nand U7837 (N_7837,N_7426,N_6371);
or U7838 (N_7838,N_6280,N_6565);
or U7839 (N_7839,N_6917,N_7087);
or U7840 (N_7840,N_7481,N_6759);
nand U7841 (N_7841,N_6069,N_6404);
and U7842 (N_7842,N_6486,N_6094);
and U7843 (N_7843,N_7325,N_6976);
and U7844 (N_7844,N_6711,N_7205);
and U7845 (N_7845,N_7435,N_7269);
nand U7846 (N_7846,N_6109,N_6692);
and U7847 (N_7847,N_6212,N_7007);
and U7848 (N_7848,N_6139,N_6704);
and U7849 (N_7849,N_6455,N_6708);
and U7850 (N_7850,N_7464,N_7057);
and U7851 (N_7851,N_6724,N_6551);
and U7852 (N_7852,N_7436,N_6174);
nand U7853 (N_7853,N_7374,N_6340);
and U7854 (N_7854,N_7164,N_6890);
nor U7855 (N_7855,N_6364,N_7384);
nor U7856 (N_7856,N_7213,N_7053);
or U7857 (N_7857,N_6907,N_6438);
or U7858 (N_7858,N_6332,N_6442);
or U7859 (N_7859,N_7399,N_6563);
nand U7860 (N_7860,N_6243,N_6259);
and U7861 (N_7861,N_6050,N_6019);
nand U7862 (N_7862,N_7300,N_6044);
and U7863 (N_7863,N_6767,N_7075);
and U7864 (N_7864,N_6459,N_6747);
nor U7865 (N_7865,N_6885,N_7061);
nor U7866 (N_7866,N_7201,N_6687);
and U7867 (N_7867,N_7150,N_6270);
nor U7868 (N_7868,N_6320,N_7081);
and U7869 (N_7869,N_6310,N_6937);
nor U7870 (N_7870,N_6756,N_7453);
nand U7871 (N_7871,N_6569,N_6436);
nand U7872 (N_7872,N_6608,N_6357);
and U7873 (N_7873,N_7333,N_6177);
nand U7874 (N_7874,N_6282,N_6089);
nor U7875 (N_7875,N_6462,N_6398);
or U7876 (N_7876,N_6439,N_6295);
nand U7877 (N_7877,N_7244,N_6523);
nor U7878 (N_7878,N_7382,N_6853);
nor U7879 (N_7879,N_6495,N_6012);
or U7880 (N_7880,N_7108,N_7156);
nor U7881 (N_7881,N_6444,N_6858);
and U7882 (N_7882,N_6227,N_6707);
or U7883 (N_7883,N_6097,N_6576);
nor U7884 (N_7884,N_6511,N_6079);
and U7885 (N_7885,N_6016,N_7280);
and U7886 (N_7886,N_6803,N_7006);
or U7887 (N_7887,N_7140,N_6389);
nor U7888 (N_7888,N_6661,N_6693);
nand U7889 (N_7889,N_7120,N_7366);
and U7890 (N_7890,N_6810,N_6450);
or U7891 (N_7891,N_6112,N_6408);
nand U7892 (N_7892,N_7239,N_6627);
nand U7893 (N_7893,N_7336,N_6668);
nand U7894 (N_7894,N_6904,N_7357);
nor U7895 (N_7895,N_7326,N_7012);
or U7896 (N_7896,N_7337,N_6464);
nand U7897 (N_7897,N_7465,N_6510);
nand U7898 (N_7898,N_7104,N_6413);
or U7899 (N_7899,N_6723,N_7279);
nand U7900 (N_7900,N_7330,N_7407);
and U7901 (N_7901,N_7385,N_6193);
nor U7902 (N_7902,N_6166,N_7316);
nor U7903 (N_7903,N_6536,N_6587);
nor U7904 (N_7904,N_6597,N_7153);
or U7905 (N_7905,N_6763,N_7315);
and U7906 (N_7906,N_7025,N_6781);
and U7907 (N_7907,N_6277,N_7241);
or U7908 (N_7908,N_6741,N_7327);
or U7909 (N_7909,N_7402,N_6195);
and U7910 (N_7910,N_6240,N_6087);
nor U7911 (N_7911,N_6394,N_6091);
nand U7912 (N_7912,N_6306,N_6947);
or U7913 (N_7913,N_6622,N_6125);
and U7914 (N_7914,N_6928,N_6678);
nand U7915 (N_7915,N_6084,N_6405);
or U7916 (N_7916,N_6978,N_6773);
or U7917 (N_7917,N_7386,N_6783);
nand U7918 (N_7918,N_7406,N_6342);
or U7919 (N_7919,N_6874,N_6083);
nand U7920 (N_7920,N_6467,N_6715);
nor U7921 (N_7921,N_7367,N_6525);
and U7922 (N_7922,N_6023,N_6991);
or U7923 (N_7923,N_6092,N_6312);
nor U7924 (N_7924,N_6214,N_7321);
xnor U7925 (N_7925,N_6245,N_6986);
nor U7926 (N_7926,N_6304,N_7157);
nand U7927 (N_7927,N_7251,N_7496);
nand U7928 (N_7928,N_7036,N_6757);
and U7929 (N_7929,N_6983,N_6099);
nor U7930 (N_7930,N_6491,N_7091);
or U7931 (N_7931,N_6677,N_7499);
and U7932 (N_7932,N_7192,N_6296);
and U7933 (N_7933,N_6217,N_7334);
nor U7934 (N_7934,N_6784,N_6186);
or U7935 (N_7935,N_6298,N_6453);
and U7936 (N_7936,N_6168,N_6560);
nor U7937 (N_7937,N_6647,N_6867);
and U7938 (N_7938,N_6843,N_6303);
nor U7939 (N_7939,N_7278,N_6456);
xnor U7940 (N_7940,N_6882,N_7419);
nand U7941 (N_7941,N_6263,N_6796);
and U7942 (N_7942,N_6396,N_6336);
xnor U7943 (N_7943,N_6755,N_6055);
nand U7944 (N_7944,N_7415,N_7234);
or U7945 (N_7945,N_6682,N_6936);
or U7946 (N_7946,N_6011,N_7001);
nor U7947 (N_7947,N_6972,N_6437);
nor U7948 (N_7948,N_7355,N_6219);
and U7949 (N_7949,N_6924,N_7195);
and U7950 (N_7950,N_7121,N_6203);
or U7951 (N_7951,N_6482,N_6274);
nand U7952 (N_7952,N_7020,N_6127);
or U7953 (N_7953,N_6537,N_7154);
or U7954 (N_7954,N_6283,N_7457);
and U7955 (N_7955,N_6896,N_6252);
or U7956 (N_7956,N_6746,N_6505);
nand U7957 (N_7957,N_6804,N_6242);
or U7958 (N_7958,N_7422,N_6965);
nand U7959 (N_7959,N_6239,N_6575);
nand U7960 (N_7960,N_6061,N_7189);
and U7961 (N_7961,N_7260,N_6448);
nand U7962 (N_7962,N_7167,N_7421);
or U7963 (N_7963,N_6930,N_6487);
and U7964 (N_7964,N_7411,N_6749);
or U7965 (N_7965,N_6555,N_6493);
nand U7966 (N_7966,N_6362,N_6730);
nor U7967 (N_7967,N_6021,N_6381);
nor U7968 (N_7968,N_6873,N_6297);
and U7969 (N_7969,N_6397,N_7314);
or U7970 (N_7970,N_6290,N_6425);
nor U7971 (N_7971,N_6305,N_6500);
and U7972 (N_7972,N_6419,N_6905);
or U7973 (N_7973,N_6040,N_7127);
and U7974 (N_7974,N_7072,N_6800);
or U7975 (N_7975,N_6328,N_7003);
nor U7976 (N_7976,N_6527,N_7069);
or U7977 (N_7977,N_6220,N_6766);
nand U7978 (N_7978,N_6942,N_7286);
and U7979 (N_7979,N_6039,N_6546);
nor U7980 (N_7980,N_7088,N_6403);
or U7981 (N_7981,N_6507,N_7034);
nor U7982 (N_7982,N_6679,N_7045);
nor U7983 (N_7983,N_6792,N_7293);
and U7984 (N_7984,N_6970,N_6353);
nor U7985 (N_7985,N_7093,N_7359);
nor U7986 (N_7986,N_6915,N_6703);
nand U7987 (N_7987,N_7341,N_6474);
nor U7988 (N_7988,N_6377,N_6695);
nor U7989 (N_7989,N_6101,N_7067);
nand U7990 (N_7990,N_7137,N_6185);
nor U7991 (N_7991,N_6619,N_7113);
or U7992 (N_7992,N_7303,N_6088);
or U7993 (N_7993,N_6777,N_6694);
and U7994 (N_7994,N_6107,N_7176);
and U7995 (N_7995,N_7488,N_6035);
nand U7996 (N_7996,N_7133,N_6683);
and U7997 (N_7997,N_7317,N_7486);
nor U7998 (N_7998,N_6601,N_6996);
or U7999 (N_7999,N_7042,N_6104);
nand U8000 (N_8000,N_6820,N_7106);
nor U8001 (N_8001,N_6981,N_6697);
nand U8002 (N_8002,N_6964,N_6617);
and U8003 (N_8003,N_6457,N_6852);
or U8004 (N_8004,N_6822,N_6052);
or U8005 (N_8005,N_6628,N_6465);
and U8006 (N_8006,N_6630,N_7271);
or U8007 (N_8007,N_7487,N_6554);
nand U8008 (N_8008,N_6686,N_6176);
or U8009 (N_8009,N_6761,N_6669);
and U8010 (N_8010,N_7105,N_6003);
nand U8011 (N_8011,N_7400,N_6504);
or U8012 (N_8012,N_6705,N_7235);
or U8013 (N_8013,N_6689,N_6356);
nand U8014 (N_8014,N_6188,N_6877);
nor U8015 (N_8015,N_7323,N_7250);
nand U8016 (N_8016,N_7455,N_6323);
nor U8017 (N_8017,N_6717,N_6256);
or U8018 (N_8018,N_7309,N_6347);
nor U8019 (N_8019,N_6041,N_6468);
or U8020 (N_8020,N_6351,N_6429);
nand U8021 (N_8021,N_6794,N_6549);
and U8022 (N_8022,N_6906,N_6698);
and U8023 (N_8023,N_6476,N_6454);
or U8024 (N_8024,N_6909,N_7490);
nand U8025 (N_8025,N_7389,N_6670);
and U8026 (N_8026,N_6278,N_7243);
nor U8027 (N_8027,N_6447,N_6681);
nor U8028 (N_8028,N_6879,N_6821);
nor U8029 (N_8029,N_6234,N_6010);
nand U8030 (N_8030,N_6656,N_6379);
nor U8031 (N_8031,N_7483,N_7163);
and U8032 (N_8032,N_7458,N_6539);
and U8033 (N_8033,N_6074,N_6813);
nor U8034 (N_8034,N_6266,N_6571);
nor U8035 (N_8035,N_7297,N_6809);
or U8036 (N_8036,N_6331,N_6955);
nand U8037 (N_8037,N_7393,N_7257);
nor U8038 (N_8038,N_6864,N_6831);
and U8039 (N_8039,N_6618,N_6249);
nor U8040 (N_8040,N_6534,N_7238);
and U8041 (N_8041,N_6714,N_7392);
nor U8042 (N_8042,N_6365,N_7267);
or U8043 (N_8043,N_6210,N_6998);
nor U8044 (N_8044,N_6206,N_6197);
nor U8045 (N_8045,N_7489,N_7283);
nand U8046 (N_8046,N_7060,N_7165);
nor U8047 (N_8047,N_6434,N_6760);
nand U8048 (N_8048,N_6772,N_6570);
nor U8049 (N_8049,N_6311,N_6994);
or U8050 (N_8050,N_7033,N_6067);
and U8051 (N_8051,N_6502,N_6343);
nor U8052 (N_8052,N_6244,N_6360);
and U8053 (N_8053,N_6805,N_7111);
nor U8054 (N_8054,N_6920,N_7245);
nand U8055 (N_8055,N_6209,N_7136);
nand U8056 (N_8056,N_6728,N_6123);
nand U8057 (N_8057,N_6172,N_6911);
and U8058 (N_8058,N_6013,N_6859);
nand U8059 (N_8059,N_6583,N_7497);
nor U8060 (N_8060,N_7004,N_7199);
or U8061 (N_8061,N_6940,N_6113);
nor U8062 (N_8062,N_6390,N_6995);
and U8063 (N_8063,N_6526,N_6880);
and U8064 (N_8064,N_6848,N_7380);
nor U8065 (N_8065,N_6309,N_7395);
and U8066 (N_8066,N_6187,N_7107);
nor U8067 (N_8067,N_6409,N_7375);
or U8068 (N_8068,N_6145,N_7051);
nor U8069 (N_8069,N_6287,N_6643);
and U8070 (N_8070,N_6110,N_7231);
nand U8071 (N_8071,N_7474,N_7273);
and U8072 (N_8072,N_6338,N_7338);
and U8073 (N_8073,N_7138,N_6959);
nand U8074 (N_8074,N_7433,N_7079);
or U8075 (N_8075,N_6899,N_6329);
or U8076 (N_8076,N_6056,N_7206);
nand U8077 (N_8077,N_6819,N_6286);
and U8078 (N_8078,N_6264,N_6326);
and U8079 (N_8079,N_7198,N_6585);
and U8080 (N_8080,N_7005,N_6762);
and U8081 (N_8081,N_6826,N_6335);
nand U8082 (N_8082,N_7319,N_6032);
or U8083 (N_8083,N_7095,N_6786);
nand U8084 (N_8084,N_6288,N_6950);
nor U8085 (N_8085,N_7335,N_6138);
and U8086 (N_8086,N_6231,N_6313);
nor U8087 (N_8087,N_7352,N_6787);
or U8088 (N_8088,N_6508,N_7084);
and U8089 (N_8089,N_6888,N_7035);
nand U8090 (N_8090,N_7346,N_6165);
or U8091 (N_8091,N_6725,N_7240);
nand U8092 (N_8092,N_6719,N_7122);
or U8093 (N_8093,N_7018,N_6395);
or U8094 (N_8094,N_7096,N_6066);
or U8095 (N_8095,N_7146,N_7225);
or U8096 (N_8096,N_6423,N_6596);
and U8097 (N_8097,N_7254,N_7417);
and U8098 (N_8098,N_6484,N_7347);
nand U8099 (N_8099,N_6960,N_6427);
nand U8100 (N_8100,N_7190,N_6748);
xnor U8101 (N_8101,N_6237,N_6251);
nand U8102 (N_8102,N_6135,N_6173);
nor U8103 (N_8103,N_6432,N_6337);
nand U8104 (N_8104,N_6002,N_6559);
or U8105 (N_8105,N_7145,N_6065);
nor U8106 (N_8106,N_6230,N_6382);
and U8107 (N_8107,N_6302,N_6577);
nor U8108 (N_8108,N_6376,N_6047);
or U8109 (N_8109,N_7015,N_7068);
and U8110 (N_8110,N_6954,N_6961);
nand U8111 (N_8111,N_6878,N_6548);
or U8112 (N_8112,N_7126,N_6407);
or U8113 (N_8113,N_6152,N_7010);
nor U8114 (N_8114,N_7277,N_7365);
nor U8115 (N_8115,N_7233,N_6635);
nor U8116 (N_8116,N_6901,N_6184);
nor U8117 (N_8117,N_6979,N_6111);
and U8118 (N_8118,N_6515,N_6736);
nand U8119 (N_8119,N_6098,N_6318);
or U8120 (N_8120,N_6737,N_6530);
nand U8121 (N_8121,N_6868,N_6070);
and U8122 (N_8122,N_6506,N_6646);
or U8123 (N_8123,N_6621,N_6863);
and U8124 (N_8124,N_6645,N_6806);
nand U8125 (N_8125,N_6481,N_6179);
and U8126 (N_8126,N_7221,N_6558);
and U8127 (N_8127,N_7282,N_6155);
and U8128 (N_8128,N_7320,N_6561);
and U8129 (N_8129,N_6605,N_6391);
and U8130 (N_8130,N_6399,N_7440);
or U8131 (N_8131,N_7110,N_7052);
or U8132 (N_8132,N_7255,N_6344);
nor U8133 (N_8133,N_6847,N_6811);
or U8134 (N_8134,N_6967,N_7461);
or U8135 (N_8135,N_6030,N_6034);
nor U8136 (N_8136,N_6485,N_7482);
or U8137 (N_8137,N_6017,N_6542);
or U8138 (N_8138,N_6386,N_6790);
and U8139 (N_8139,N_7348,N_6778);
and U8140 (N_8140,N_7227,N_6823);
nand U8141 (N_8141,N_6489,N_6175);
nand U8142 (N_8142,N_6659,N_6688);
nand U8143 (N_8143,N_7418,N_7287);
nand U8144 (N_8144,N_6919,N_6828);
or U8145 (N_8145,N_7484,N_7191);
and U8146 (N_8146,N_6255,N_7182);
or U8147 (N_8147,N_7070,N_6503);
and U8148 (N_8148,N_6528,N_7083);
or U8149 (N_8149,N_7155,N_6440);
nor U8150 (N_8150,N_6146,N_6604);
nor U8151 (N_8151,N_6415,N_6075);
or U8152 (N_8152,N_6093,N_6073);
and U8153 (N_8153,N_6949,N_7361);
or U8154 (N_8154,N_7021,N_7248);
and U8155 (N_8155,N_6931,N_7430);
or U8156 (N_8156,N_6520,N_6639);
and U8157 (N_8157,N_6660,N_7197);
nand U8158 (N_8158,N_6143,N_6720);
or U8159 (N_8159,N_6218,N_6233);
nand U8160 (N_8160,N_7295,N_6037);
nand U8161 (N_8161,N_6975,N_6327);
or U8162 (N_8162,N_6106,N_7247);
xor U8163 (N_8163,N_6592,N_6420);
nor U8164 (N_8164,N_6775,N_6406);
nor U8165 (N_8165,N_6024,N_6449);
xor U8166 (N_8166,N_7116,N_6317);
nand U8167 (N_8167,N_6253,N_6402);
and U8168 (N_8168,N_6136,N_6150);
and U8169 (N_8169,N_7449,N_7468);
nand U8170 (N_8170,N_6477,N_6238);
nor U8171 (N_8171,N_6799,N_6837);
and U8172 (N_8172,N_6552,N_7253);
nand U8173 (N_8173,N_6529,N_6729);
xor U8174 (N_8174,N_6891,N_6096);
or U8175 (N_8175,N_7364,N_6121);
nor U8176 (N_8176,N_6435,N_7047);
nand U8177 (N_8177,N_6625,N_6611);
nand U8178 (N_8178,N_7224,N_6716);
and U8179 (N_8179,N_7059,N_7268);
nand U8180 (N_8180,N_6743,N_6889);
nand U8181 (N_8181,N_7363,N_6633);
and U8182 (N_8182,N_7304,N_7204);
and U8183 (N_8183,N_7080,N_6626);
xnor U8184 (N_8184,N_6607,N_7408);
and U8185 (N_8185,N_6620,N_7390);
nor U8186 (N_8186,N_7423,N_7082);
or U8187 (N_8187,N_6062,N_6385);
nand U8188 (N_8188,N_6550,N_7351);
or U8189 (N_8189,N_6815,N_7404);
and U8190 (N_8190,N_6632,N_6100);
nand U8191 (N_8191,N_6285,N_6366);
and U8192 (N_8192,N_7466,N_7161);
or U8193 (N_8193,N_6025,N_6513);
nor U8194 (N_8194,N_7289,N_7023);
nor U8195 (N_8195,N_6941,N_6514);
or U8196 (N_8196,N_6912,N_6018);
or U8197 (N_8197,N_6827,N_6102);
or U8198 (N_8198,N_6854,N_7175);
and U8199 (N_8199,N_7103,N_6613);
nand U8200 (N_8200,N_7312,N_6624);
nor U8201 (N_8201,N_6480,N_7439);
and U8202 (N_8202,N_6580,N_6665);
nor U8203 (N_8203,N_7479,N_6488);
and U8204 (N_8204,N_6076,N_6181);
and U8205 (N_8205,N_6005,N_6142);
or U8206 (N_8206,N_6272,N_7112);
nor U8207 (N_8207,N_6015,N_7447);
or U8208 (N_8208,N_7409,N_6638);
or U8209 (N_8209,N_7168,N_6926);
or U8210 (N_8210,N_7063,N_6053);
and U8211 (N_8211,N_7416,N_6532);
and U8212 (N_8212,N_6333,N_6712);
nor U8213 (N_8213,N_6494,N_6205);
nand U8214 (N_8214,N_6276,N_6946);
or U8215 (N_8215,N_7014,N_6598);
or U8216 (N_8216,N_7388,N_7299);
and U8217 (N_8217,N_7236,N_6553);
nand U8218 (N_8218,N_7098,N_7044);
or U8219 (N_8219,N_6969,N_6938);
nor U8220 (N_8220,N_6640,N_7013);
nand U8221 (N_8221,N_7469,N_6614);
nor U8222 (N_8222,N_6426,N_6769);
and U8223 (N_8223,N_6958,N_6314);
nor U8224 (N_8224,N_6615,N_6895);
or U8225 (N_8225,N_7152,N_7291);
nor U8226 (N_8226,N_6250,N_7037);
or U8227 (N_8227,N_6801,N_7373);
nand U8228 (N_8228,N_6241,N_6839);
nand U8229 (N_8229,N_6788,N_6334);
and U8230 (N_8230,N_6568,N_6779);
and U8231 (N_8231,N_6742,N_7129);
nand U8232 (N_8232,N_6046,N_6445);
nor U8233 (N_8233,N_7141,N_6144);
nor U8234 (N_8234,N_6791,N_6064);
nand U8235 (N_8235,N_6860,N_6354);
nor U8236 (N_8236,N_6443,N_6446);
nor U8237 (N_8237,N_6501,N_7054);
nand U8238 (N_8238,N_6275,N_7134);
nand U8239 (N_8239,N_6648,N_6968);
nor U8240 (N_8240,N_6562,N_6997);
nand U8241 (N_8241,N_6315,N_6022);
nor U8242 (N_8242,N_6132,N_6838);
xnor U8243 (N_8243,N_7211,N_6049);
or U8244 (N_8244,N_6226,N_6133);
nand U8245 (N_8245,N_6673,N_6922);
or U8246 (N_8246,N_6980,N_6887);
nand U8247 (N_8247,N_7370,N_6871);
or U8248 (N_8248,N_6128,N_7029);
and U8249 (N_8249,N_6269,N_7086);
nor U8250 (N_8250,N_6274,N_7355);
nand U8251 (N_8251,N_7142,N_6177);
or U8252 (N_8252,N_6390,N_7023);
and U8253 (N_8253,N_7395,N_7138);
nor U8254 (N_8254,N_7397,N_7459);
and U8255 (N_8255,N_7495,N_6239);
nor U8256 (N_8256,N_6193,N_6673);
and U8257 (N_8257,N_7166,N_7227);
nor U8258 (N_8258,N_6006,N_6955);
nand U8259 (N_8259,N_6494,N_7316);
or U8260 (N_8260,N_7442,N_6247);
nor U8261 (N_8261,N_6770,N_6717);
nor U8262 (N_8262,N_6242,N_6903);
or U8263 (N_8263,N_7353,N_6126);
or U8264 (N_8264,N_6955,N_7185);
nand U8265 (N_8265,N_7374,N_7348);
nor U8266 (N_8266,N_6425,N_6046);
nor U8267 (N_8267,N_6693,N_6675);
or U8268 (N_8268,N_6666,N_6867);
or U8269 (N_8269,N_7176,N_6836);
or U8270 (N_8270,N_6353,N_6333);
and U8271 (N_8271,N_6847,N_7067);
and U8272 (N_8272,N_6683,N_6938);
or U8273 (N_8273,N_7354,N_6825);
nand U8274 (N_8274,N_7271,N_6235);
nand U8275 (N_8275,N_6346,N_7358);
or U8276 (N_8276,N_6213,N_6443);
nand U8277 (N_8277,N_6551,N_6150);
nand U8278 (N_8278,N_7340,N_6724);
nor U8279 (N_8279,N_7169,N_7277);
or U8280 (N_8280,N_6358,N_7081);
nor U8281 (N_8281,N_6819,N_7196);
and U8282 (N_8282,N_6114,N_6524);
or U8283 (N_8283,N_6358,N_7498);
nand U8284 (N_8284,N_6610,N_6953);
and U8285 (N_8285,N_7197,N_7316);
nor U8286 (N_8286,N_7455,N_6608);
nor U8287 (N_8287,N_6376,N_7272);
nor U8288 (N_8288,N_6299,N_6796);
nor U8289 (N_8289,N_6643,N_7086);
nand U8290 (N_8290,N_6681,N_7379);
nand U8291 (N_8291,N_6462,N_6241);
nand U8292 (N_8292,N_7492,N_6975);
nand U8293 (N_8293,N_7199,N_6536);
nand U8294 (N_8294,N_7494,N_6313);
and U8295 (N_8295,N_6906,N_7203);
and U8296 (N_8296,N_6017,N_6831);
or U8297 (N_8297,N_6914,N_6678);
nand U8298 (N_8298,N_6742,N_6859);
or U8299 (N_8299,N_6713,N_6754);
or U8300 (N_8300,N_7460,N_6479);
nand U8301 (N_8301,N_6206,N_7317);
nand U8302 (N_8302,N_6723,N_6609);
nand U8303 (N_8303,N_6901,N_6013);
and U8304 (N_8304,N_6084,N_6324);
or U8305 (N_8305,N_7211,N_6866);
and U8306 (N_8306,N_6546,N_7279);
or U8307 (N_8307,N_6949,N_6581);
or U8308 (N_8308,N_6468,N_7081);
and U8309 (N_8309,N_6274,N_6282);
nand U8310 (N_8310,N_7111,N_6045);
and U8311 (N_8311,N_6342,N_6893);
nand U8312 (N_8312,N_7302,N_6842);
nand U8313 (N_8313,N_6573,N_7308);
and U8314 (N_8314,N_7327,N_6355);
xor U8315 (N_8315,N_7366,N_7007);
nor U8316 (N_8316,N_7288,N_6407);
nor U8317 (N_8317,N_7085,N_6529);
and U8318 (N_8318,N_7430,N_6448);
nand U8319 (N_8319,N_6761,N_7468);
and U8320 (N_8320,N_6931,N_7382);
and U8321 (N_8321,N_7003,N_6578);
nand U8322 (N_8322,N_6435,N_6103);
nor U8323 (N_8323,N_6816,N_6521);
nand U8324 (N_8324,N_6224,N_6190);
and U8325 (N_8325,N_6917,N_6564);
nand U8326 (N_8326,N_6263,N_7349);
nor U8327 (N_8327,N_7330,N_6555);
and U8328 (N_8328,N_6468,N_6675);
or U8329 (N_8329,N_6453,N_6538);
and U8330 (N_8330,N_6258,N_6668);
nand U8331 (N_8331,N_7240,N_7121);
or U8332 (N_8332,N_6582,N_7446);
nand U8333 (N_8333,N_6264,N_6931);
and U8334 (N_8334,N_7228,N_7208);
nor U8335 (N_8335,N_7197,N_6504);
and U8336 (N_8336,N_7128,N_6827);
nand U8337 (N_8337,N_6739,N_7366);
nor U8338 (N_8338,N_6808,N_7386);
nand U8339 (N_8339,N_6206,N_6289);
and U8340 (N_8340,N_7231,N_7314);
nand U8341 (N_8341,N_6390,N_6645);
nor U8342 (N_8342,N_6458,N_6715);
and U8343 (N_8343,N_6120,N_6872);
or U8344 (N_8344,N_6539,N_7024);
and U8345 (N_8345,N_6779,N_6754);
nor U8346 (N_8346,N_6583,N_6024);
nor U8347 (N_8347,N_6921,N_6063);
or U8348 (N_8348,N_7002,N_6548);
nand U8349 (N_8349,N_6911,N_6898);
or U8350 (N_8350,N_7208,N_7286);
nor U8351 (N_8351,N_6612,N_6362);
or U8352 (N_8352,N_6072,N_6258);
or U8353 (N_8353,N_6223,N_6255);
nor U8354 (N_8354,N_6195,N_7092);
and U8355 (N_8355,N_6295,N_6212);
nand U8356 (N_8356,N_6865,N_6653);
or U8357 (N_8357,N_7490,N_6645);
nor U8358 (N_8358,N_7401,N_6819);
nand U8359 (N_8359,N_7426,N_6749);
nand U8360 (N_8360,N_6134,N_6966);
nor U8361 (N_8361,N_7179,N_7410);
or U8362 (N_8362,N_6030,N_6049);
nand U8363 (N_8363,N_6257,N_7298);
nor U8364 (N_8364,N_6350,N_6243);
or U8365 (N_8365,N_6287,N_6177);
nand U8366 (N_8366,N_6699,N_6257);
nand U8367 (N_8367,N_7116,N_6367);
nand U8368 (N_8368,N_7411,N_6627);
nand U8369 (N_8369,N_6723,N_6069);
or U8370 (N_8370,N_7325,N_7182);
nor U8371 (N_8371,N_6663,N_6356);
xor U8372 (N_8372,N_7113,N_6969);
nor U8373 (N_8373,N_6071,N_7444);
nor U8374 (N_8374,N_6231,N_7421);
and U8375 (N_8375,N_6667,N_7025);
or U8376 (N_8376,N_6966,N_6788);
nor U8377 (N_8377,N_7089,N_7305);
nand U8378 (N_8378,N_7092,N_7379);
nor U8379 (N_8379,N_7375,N_6221);
nor U8380 (N_8380,N_7422,N_7060);
and U8381 (N_8381,N_6946,N_6857);
nor U8382 (N_8382,N_6269,N_6476);
nor U8383 (N_8383,N_7409,N_7334);
or U8384 (N_8384,N_6530,N_6451);
nand U8385 (N_8385,N_7085,N_6223);
and U8386 (N_8386,N_6378,N_6610);
nand U8387 (N_8387,N_7431,N_6926);
or U8388 (N_8388,N_7290,N_7392);
or U8389 (N_8389,N_7464,N_6432);
or U8390 (N_8390,N_7113,N_6251);
nor U8391 (N_8391,N_6137,N_6057);
nand U8392 (N_8392,N_6837,N_6087);
or U8393 (N_8393,N_6983,N_7197);
or U8394 (N_8394,N_6901,N_6082);
nor U8395 (N_8395,N_6226,N_7178);
or U8396 (N_8396,N_7140,N_6198);
or U8397 (N_8397,N_6021,N_7337);
and U8398 (N_8398,N_6303,N_7179);
or U8399 (N_8399,N_7187,N_6840);
nor U8400 (N_8400,N_7049,N_7016);
and U8401 (N_8401,N_6629,N_6559);
nand U8402 (N_8402,N_6134,N_6567);
or U8403 (N_8403,N_6569,N_6674);
nand U8404 (N_8404,N_7332,N_6380);
nand U8405 (N_8405,N_6226,N_6946);
nand U8406 (N_8406,N_6806,N_6782);
nand U8407 (N_8407,N_6045,N_6598);
and U8408 (N_8408,N_7344,N_7355);
or U8409 (N_8409,N_6249,N_7449);
nand U8410 (N_8410,N_6550,N_7140);
and U8411 (N_8411,N_6579,N_6719);
nand U8412 (N_8412,N_7480,N_7116);
nor U8413 (N_8413,N_6827,N_6154);
nand U8414 (N_8414,N_6159,N_6995);
and U8415 (N_8415,N_6434,N_6260);
nor U8416 (N_8416,N_6987,N_6292);
nand U8417 (N_8417,N_6645,N_6571);
and U8418 (N_8418,N_6688,N_7094);
nor U8419 (N_8419,N_7357,N_7048);
and U8420 (N_8420,N_6226,N_6081);
nand U8421 (N_8421,N_7176,N_7001);
nand U8422 (N_8422,N_6926,N_7435);
and U8423 (N_8423,N_6977,N_6586);
or U8424 (N_8424,N_6279,N_6764);
nand U8425 (N_8425,N_7031,N_6885);
nand U8426 (N_8426,N_6097,N_6012);
nor U8427 (N_8427,N_6835,N_7391);
nor U8428 (N_8428,N_6196,N_6231);
and U8429 (N_8429,N_6249,N_6940);
nor U8430 (N_8430,N_6255,N_6096);
nor U8431 (N_8431,N_7027,N_6567);
and U8432 (N_8432,N_6401,N_6580);
nor U8433 (N_8433,N_6691,N_6103);
nor U8434 (N_8434,N_6667,N_7155);
and U8435 (N_8435,N_7006,N_7225);
and U8436 (N_8436,N_6925,N_6675);
and U8437 (N_8437,N_6111,N_7378);
nor U8438 (N_8438,N_6511,N_6880);
nor U8439 (N_8439,N_6443,N_6786);
or U8440 (N_8440,N_6441,N_6892);
or U8441 (N_8441,N_6663,N_6170);
nor U8442 (N_8442,N_6768,N_6515);
nand U8443 (N_8443,N_7137,N_7294);
nand U8444 (N_8444,N_7070,N_6232);
or U8445 (N_8445,N_6868,N_7055);
nand U8446 (N_8446,N_6408,N_7324);
or U8447 (N_8447,N_6849,N_7037);
nor U8448 (N_8448,N_6489,N_7097);
or U8449 (N_8449,N_7162,N_7204);
or U8450 (N_8450,N_6142,N_6085);
or U8451 (N_8451,N_6310,N_6335);
or U8452 (N_8452,N_7088,N_7299);
and U8453 (N_8453,N_6156,N_7212);
and U8454 (N_8454,N_6066,N_7007);
nor U8455 (N_8455,N_6244,N_6596);
and U8456 (N_8456,N_7253,N_6721);
and U8457 (N_8457,N_6852,N_7288);
nand U8458 (N_8458,N_6757,N_7422);
nand U8459 (N_8459,N_6645,N_6408);
nand U8460 (N_8460,N_7135,N_6246);
nand U8461 (N_8461,N_7275,N_6158);
nand U8462 (N_8462,N_6819,N_7389);
nor U8463 (N_8463,N_6460,N_6535);
nor U8464 (N_8464,N_6858,N_7152);
nand U8465 (N_8465,N_6389,N_7450);
or U8466 (N_8466,N_7010,N_7287);
and U8467 (N_8467,N_7115,N_6616);
and U8468 (N_8468,N_6009,N_6301);
nand U8469 (N_8469,N_6331,N_6621);
nor U8470 (N_8470,N_7265,N_6926);
or U8471 (N_8471,N_7271,N_6147);
nor U8472 (N_8472,N_6963,N_6084);
xor U8473 (N_8473,N_7470,N_7187);
or U8474 (N_8474,N_6246,N_6263);
and U8475 (N_8475,N_6368,N_7387);
nor U8476 (N_8476,N_6083,N_6970);
or U8477 (N_8477,N_6332,N_7117);
or U8478 (N_8478,N_6761,N_7414);
nor U8479 (N_8479,N_6858,N_7478);
nor U8480 (N_8480,N_6833,N_6581);
or U8481 (N_8481,N_6871,N_6970);
nand U8482 (N_8482,N_7453,N_6243);
nor U8483 (N_8483,N_6100,N_6543);
or U8484 (N_8484,N_7132,N_6413);
and U8485 (N_8485,N_6894,N_7318);
or U8486 (N_8486,N_6092,N_7284);
nand U8487 (N_8487,N_6837,N_6843);
nand U8488 (N_8488,N_7254,N_7236);
nor U8489 (N_8489,N_7421,N_6045);
and U8490 (N_8490,N_7241,N_7462);
and U8491 (N_8491,N_6475,N_6477);
and U8492 (N_8492,N_6557,N_6426);
and U8493 (N_8493,N_6314,N_6501);
and U8494 (N_8494,N_6854,N_7429);
nand U8495 (N_8495,N_6235,N_6602);
nor U8496 (N_8496,N_6647,N_6176);
and U8497 (N_8497,N_6247,N_7264);
nand U8498 (N_8498,N_7153,N_6018);
nand U8499 (N_8499,N_7125,N_7373);
and U8500 (N_8500,N_6536,N_6907);
nor U8501 (N_8501,N_6267,N_7034);
and U8502 (N_8502,N_7283,N_6939);
nand U8503 (N_8503,N_6338,N_6597);
and U8504 (N_8504,N_6903,N_6691);
nand U8505 (N_8505,N_7255,N_6842);
nor U8506 (N_8506,N_7368,N_6699);
and U8507 (N_8507,N_7406,N_6266);
nor U8508 (N_8508,N_6367,N_6337);
or U8509 (N_8509,N_6398,N_6751);
nor U8510 (N_8510,N_6394,N_7318);
nand U8511 (N_8511,N_7146,N_7148);
nand U8512 (N_8512,N_7073,N_6095);
and U8513 (N_8513,N_7041,N_6874);
and U8514 (N_8514,N_7221,N_6737);
or U8515 (N_8515,N_6052,N_6032);
and U8516 (N_8516,N_7305,N_6215);
or U8517 (N_8517,N_6728,N_6399);
nor U8518 (N_8518,N_6402,N_7456);
nor U8519 (N_8519,N_7084,N_6969);
and U8520 (N_8520,N_7430,N_6003);
or U8521 (N_8521,N_6247,N_7335);
nand U8522 (N_8522,N_7168,N_6413);
and U8523 (N_8523,N_7156,N_6253);
or U8524 (N_8524,N_6882,N_7228);
nor U8525 (N_8525,N_6742,N_6175);
nor U8526 (N_8526,N_6682,N_6427);
nor U8527 (N_8527,N_6974,N_6679);
nor U8528 (N_8528,N_7066,N_7200);
or U8529 (N_8529,N_6163,N_7279);
or U8530 (N_8530,N_6573,N_6984);
or U8531 (N_8531,N_6179,N_6530);
nand U8532 (N_8532,N_7236,N_7214);
and U8533 (N_8533,N_6445,N_6481);
or U8534 (N_8534,N_6997,N_6804);
and U8535 (N_8535,N_7313,N_6661);
and U8536 (N_8536,N_6914,N_6094);
and U8537 (N_8537,N_6503,N_6828);
and U8538 (N_8538,N_6772,N_6230);
or U8539 (N_8539,N_6229,N_6341);
or U8540 (N_8540,N_7293,N_7012);
and U8541 (N_8541,N_6250,N_6633);
nor U8542 (N_8542,N_7108,N_6962);
and U8543 (N_8543,N_6593,N_6105);
or U8544 (N_8544,N_7062,N_7036);
or U8545 (N_8545,N_7040,N_6711);
or U8546 (N_8546,N_6891,N_6503);
and U8547 (N_8547,N_6961,N_6330);
or U8548 (N_8548,N_7005,N_6767);
and U8549 (N_8549,N_7399,N_6541);
and U8550 (N_8550,N_7333,N_6381);
nand U8551 (N_8551,N_7029,N_6975);
or U8552 (N_8552,N_6415,N_7142);
or U8553 (N_8553,N_6065,N_6366);
nand U8554 (N_8554,N_6555,N_6449);
nand U8555 (N_8555,N_6679,N_6941);
or U8556 (N_8556,N_6708,N_7181);
nor U8557 (N_8557,N_6950,N_7221);
and U8558 (N_8558,N_6118,N_6620);
nand U8559 (N_8559,N_6095,N_6638);
and U8560 (N_8560,N_6754,N_6609);
nor U8561 (N_8561,N_7307,N_7415);
nor U8562 (N_8562,N_6963,N_6104);
nor U8563 (N_8563,N_6339,N_6344);
or U8564 (N_8564,N_7126,N_7359);
nor U8565 (N_8565,N_7104,N_7348);
and U8566 (N_8566,N_7105,N_6306);
or U8567 (N_8567,N_7009,N_7429);
nand U8568 (N_8568,N_7398,N_7478);
or U8569 (N_8569,N_7299,N_7421);
nand U8570 (N_8570,N_6409,N_6929);
nor U8571 (N_8571,N_6818,N_7030);
nor U8572 (N_8572,N_6615,N_7267);
nor U8573 (N_8573,N_7179,N_7487);
or U8574 (N_8574,N_7261,N_7264);
and U8575 (N_8575,N_6643,N_7403);
and U8576 (N_8576,N_6545,N_6848);
or U8577 (N_8577,N_6887,N_7039);
nor U8578 (N_8578,N_6355,N_6661);
or U8579 (N_8579,N_6433,N_7250);
nand U8580 (N_8580,N_6993,N_6414);
or U8581 (N_8581,N_6459,N_6489);
and U8582 (N_8582,N_6138,N_6719);
nand U8583 (N_8583,N_7317,N_6615);
nand U8584 (N_8584,N_7225,N_6251);
and U8585 (N_8585,N_7167,N_6414);
and U8586 (N_8586,N_6530,N_7073);
and U8587 (N_8587,N_7445,N_7175);
nand U8588 (N_8588,N_6754,N_6811);
nor U8589 (N_8589,N_6766,N_7020);
and U8590 (N_8590,N_6482,N_6381);
xnor U8591 (N_8591,N_7263,N_6850);
and U8592 (N_8592,N_6684,N_6925);
or U8593 (N_8593,N_6012,N_6477);
nand U8594 (N_8594,N_6062,N_7063);
and U8595 (N_8595,N_6035,N_6565);
nand U8596 (N_8596,N_6699,N_6798);
xor U8597 (N_8597,N_6834,N_6728);
or U8598 (N_8598,N_7157,N_6480);
and U8599 (N_8599,N_6204,N_6604);
nand U8600 (N_8600,N_6141,N_7103);
or U8601 (N_8601,N_6351,N_7017);
or U8602 (N_8602,N_6371,N_7377);
or U8603 (N_8603,N_6680,N_7350);
or U8604 (N_8604,N_6088,N_7257);
nor U8605 (N_8605,N_7288,N_7048);
or U8606 (N_8606,N_7041,N_6819);
and U8607 (N_8607,N_6607,N_6034);
nand U8608 (N_8608,N_6965,N_7069);
nor U8609 (N_8609,N_7161,N_7315);
nor U8610 (N_8610,N_6960,N_6932);
or U8611 (N_8611,N_7199,N_6808);
nand U8612 (N_8612,N_6110,N_7151);
nand U8613 (N_8613,N_6942,N_6675);
nor U8614 (N_8614,N_6774,N_7142);
or U8615 (N_8615,N_6190,N_6456);
nor U8616 (N_8616,N_6264,N_6285);
and U8617 (N_8617,N_6033,N_6585);
nand U8618 (N_8618,N_6001,N_6868);
xnor U8619 (N_8619,N_6049,N_7149);
nand U8620 (N_8620,N_6578,N_6726);
or U8621 (N_8621,N_6445,N_6656);
or U8622 (N_8622,N_6770,N_6230);
or U8623 (N_8623,N_6625,N_6469);
and U8624 (N_8624,N_7337,N_6332);
or U8625 (N_8625,N_7123,N_6184);
nor U8626 (N_8626,N_6806,N_6983);
nor U8627 (N_8627,N_6405,N_7488);
and U8628 (N_8628,N_7067,N_7199);
or U8629 (N_8629,N_7274,N_7133);
nand U8630 (N_8630,N_6189,N_6899);
and U8631 (N_8631,N_6008,N_6836);
nor U8632 (N_8632,N_6796,N_6024);
or U8633 (N_8633,N_7033,N_6677);
nand U8634 (N_8634,N_6088,N_6502);
or U8635 (N_8635,N_6507,N_7355);
nor U8636 (N_8636,N_6641,N_6250);
nor U8637 (N_8637,N_6957,N_6048);
nand U8638 (N_8638,N_6628,N_7084);
nand U8639 (N_8639,N_7240,N_6941);
or U8640 (N_8640,N_6084,N_7358);
nand U8641 (N_8641,N_6265,N_6894);
nand U8642 (N_8642,N_7225,N_6519);
nor U8643 (N_8643,N_6974,N_6324);
nor U8644 (N_8644,N_7146,N_6995);
nor U8645 (N_8645,N_7239,N_6792);
nor U8646 (N_8646,N_6013,N_6338);
and U8647 (N_8647,N_6587,N_6086);
or U8648 (N_8648,N_6854,N_7143);
or U8649 (N_8649,N_6333,N_7157);
and U8650 (N_8650,N_7053,N_7260);
nand U8651 (N_8651,N_7113,N_7274);
and U8652 (N_8652,N_7351,N_6631);
and U8653 (N_8653,N_7002,N_6396);
nor U8654 (N_8654,N_6380,N_6167);
or U8655 (N_8655,N_6001,N_6313);
nor U8656 (N_8656,N_7129,N_7245);
nand U8657 (N_8657,N_6767,N_6650);
and U8658 (N_8658,N_6771,N_7143);
and U8659 (N_8659,N_6140,N_7017);
nand U8660 (N_8660,N_6424,N_6440);
or U8661 (N_8661,N_6700,N_7400);
and U8662 (N_8662,N_6765,N_6910);
xnor U8663 (N_8663,N_6218,N_6841);
nor U8664 (N_8664,N_6997,N_6507);
nor U8665 (N_8665,N_7044,N_6273);
nand U8666 (N_8666,N_6288,N_7161);
nor U8667 (N_8667,N_6350,N_6323);
and U8668 (N_8668,N_6957,N_6359);
and U8669 (N_8669,N_6800,N_6980);
nor U8670 (N_8670,N_6931,N_6085);
and U8671 (N_8671,N_7124,N_7419);
and U8672 (N_8672,N_6206,N_6339);
nor U8673 (N_8673,N_6386,N_7158);
and U8674 (N_8674,N_7461,N_6505);
or U8675 (N_8675,N_7228,N_6521);
nand U8676 (N_8676,N_7204,N_7141);
or U8677 (N_8677,N_6157,N_6809);
or U8678 (N_8678,N_6782,N_6058);
nand U8679 (N_8679,N_6466,N_6169);
and U8680 (N_8680,N_6681,N_6228);
and U8681 (N_8681,N_6654,N_7315);
nand U8682 (N_8682,N_6607,N_7482);
nand U8683 (N_8683,N_6085,N_7136);
or U8684 (N_8684,N_6734,N_6862);
nor U8685 (N_8685,N_6238,N_7127);
or U8686 (N_8686,N_7430,N_7125);
or U8687 (N_8687,N_6320,N_7348);
or U8688 (N_8688,N_6451,N_6261);
or U8689 (N_8689,N_6317,N_6825);
nor U8690 (N_8690,N_6269,N_6369);
or U8691 (N_8691,N_7206,N_6849);
and U8692 (N_8692,N_6313,N_6839);
nand U8693 (N_8693,N_6126,N_7324);
nor U8694 (N_8694,N_6592,N_6988);
and U8695 (N_8695,N_6654,N_6640);
nor U8696 (N_8696,N_6063,N_7294);
nand U8697 (N_8697,N_7382,N_6681);
and U8698 (N_8698,N_6327,N_6282);
and U8699 (N_8699,N_6372,N_7261);
nor U8700 (N_8700,N_6055,N_6884);
and U8701 (N_8701,N_6307,N_6215);
and U8702 (N_8702,N_7474,N_6563);
nand U8703 (N_8703,N_6336,N_6255);
nor U8704 (N_8704,N_6647,N_7008);
or U8705 (N_8705,N_7120,N_7263);
or U8706 (N_8706,N_6625,N_7068);
nor U8707 (N_8707,N_7139,N_6792);
nor U8708 (N_8708,N_6816,N_6413);
and U8709 (N_8709,N_6391,N_7133);
nor U8710 (N_8710,N_6310,N_6963);
or U8711 (N_8711,N_7349,N_6404);
nand U8712 (N_8712,N_7319,N_7053);
and U8713 (N_8713,N_6322,N_6120);
nand U8714 (N_8714,N_6193,N_6674);
nor U8715 (N_8715,N_7419,N_6233);
or U8716 (N_8716,N_6085,N_6265);
nor U8717 (N_8717,N_7110,N_6570);
or U8718 (N_8718,N_7388,N_6609);
nor U8719 (N_8719,N_6857,N_6279);
nand U8720 (N_8720,N_7288,N_7410);
xnor U8721 (N_8721,N_6309,N_6552);
or U8722 (N_8722,N_7326,N_6540);
nor U8723 (N_8723,N_6385,N_7492);
or U8724 (N_8724,N_6084,N_7227);
nor U8725 (N_8725,N_7344,N_7486);
and U8726 (N_8726,N_6674,N_6421);
nand U8727 (N_8727,N_6020,N_6720);
nand U8728 (N_8728,N_6752,N_6799);
or U8729 (N_8729,N_7329,N_6697);
nand U8730 (N_8730,N_7319,N_6300);
nor U8731 (N_8731,N_6515,N_6136);
or U8732 (N_8732,N_6555,N_6237);
or U8733 (N_8733,N_6437,N_7224);
and U8734 (N_8734,N_7452,N_7344);
nand U8735 (N_8735,N_6529,N_6784);
nor U8736 (N_8736,N_6225,N_6119);
and U8737 (N_8737,N_6051,N_6574);
nor U8738 (N_8738,N_6616,N_6948);
nand U8739 (N_8739,N_6126,N_6853);
nand U8740 (N_8740,N_6144,N_7270);
and U8741 (N_8741,N_6120,N_7078);
nand U8742 (N_8742,N_6189,N_6073);
and U8743 (N_8743,N_7289,N_7467);
and U8744 (N_8744,N_7139,N_7177);
or U8745 (N_8745,N_7065,N_6613);
nand U8746 (N_8746,N_7366,N_7483);
or U8747 (N_8747,N_7144,N_7478);
nand U8748 (N_8748,N_7151,N_6779);
nor U8749 (N_8749,N_6278,N_7206);
nand U8750 (N_8750,N_7330,N_7403);
nand U8751 (N_8751,N_6633,N_6535);
or U8752 (N_8752,N_6349,N_6732);
nor U8753 (N_8753,N_6607,N_6957);
nand U8754 (N_8754,N_6408,N_6052);
xor U8755 (N_8755,N_6198,N_7019);
xnor U8756 (N_8756,N_7167,N_6484);
nand U8757 (N_8757,N_6286,N_7227);
or U8758 (N_8758,N_7206,N_6168);
nand U8759 (N_8759,N_6475,N_7210);
and U8760 (N_8760,N_6975,N_6811);
nand U8761 (N_8761,N_7279,N_6119);
or U8762 (N_8762,N_6247,N_6266);
or U8763 (N_8763,N_6763,N_6161);
and U8764 (N_8764,N_6592,N_7067);
or U8765 (N_8765,N_7138,N_6176);
nor U8766 (N_8766,N_6183,N_7003);
nand U8767 (N_8767,N_6766,N_6356);
and U8768 (N_8768,N_7311,N_7078);
and U8769 (N_8769,N_6217,N_7068);
nor U8770 (N_8770,N_6535,N_6094);
and U8771 (N_8771,N_7197,N_6042);
or U8772 (N_8772,N_6096,N_6078);
nand U8773 (N_8773,N_7354,N_7308);
and U8774 (N_8774,N_6082,N_6245);
xor U8775 (N_8775,N_6511,N_7015);
nand U8776 (N_8776,N_6751,N_6934);
nand U8777 (N_8777,N_7480,N_7207);
nand U8778 (N_8778,N_6423,N_6070);
nand U8779 (N_8779,N_7426,N_7321);
nor U8780 (N_8780,N_7304,N_7098);
nand U8781 (N_8781,N_6531,N_6144);
and U8782 (N_8782,N_6117,N_6293);
and U8783 (N_8783,N_6685,N_7088);
nand U8784 (N_8784,N_6080,N_6835);
nand U8785 (N_8785,N_6852,N_6270);
nor U8786 (N_8786,N_7294,N_6079);
nand U8787 (N_8787,N_6004,N_6023);
nor U8788 (N_8788,N_6521,N_6702);
or U8789 (N_8789,N_7218,N_6632);
nor U8790 (N_8790,N_6915,N_6879);
or U8791 (N_8791,N_6374,N_7170);
and U8792 (N_8792,N_7355,N_6627);
nand U8793 (N_8793,N_6632,N_6405);
nor U8794 (N_8794,N_7481,N_6187);
nand U8795 (N_8795,N_6631,N_6188);
nand U8796 (N_8796,N_6589,N_6529);
xor U8797 (N_8797,N_7440,N_6688);
and U8798 (N_8798,N_6979,N_6705);
or U8799 (N_8799,N_6976,N_6313);
nor U8800 (N_8800,N_6060,N_7431);
and U8801 (N_8801,N_6000,N_7332);
or U8802 (N_8802,N_7374,N_6604);
and U8803 (N_8803,N_7298,N_6092);
and U8804 (N_8804,N_6497,N_7458);
and U8805 (N_8805,N_7244,N_7470);
nand U8806 (N_8806,N_7175,N_6579);
or U8807 (N_8807,N_6811,N_7044);
and U8808 (N_8808,N_7230,N_6984);
nand U8809 (N_8809,N_6566,N_6089);
nand U8810 (N_8810,N_6394,N_6404);
or U8811 (N_8811,N_6403,N_7321);
and U8812 (N_8812,N_6280,N_7098);
and U8813 (N_8813,N_7181,N_6113);
nor U8814 (N_8814,N_7390,N_7135);
nor U8815 (N_8815,N_6074,N_6605);
and U8816 (N_8816,N_6887,N_7267);
or U8817 (N_8817,N_7298,N_6876);
or U8818 (N_8818,N_6410,N_6917);
and U8819 (N_8819,N_7338,N_7258);
nor U8820 (N_8820,N_6418,N_6175);
nor U8821 (N_8821,N_6346,N_6532);
or U8822 (N_8822,N_7368,N_6094);
and U8823 (N_8823,N_6485,N_6165);
and U8824 (N_8824,N_7276,N_6442);
or U8825 (N_8825,N_7432,N_6891);
nand U8826 (N_8826,N_7419,N_7258);
or U8827 (N_8827,N_6184,N_6383);
or U8828 (N_8828,N_6740,N_7292);
or U8829 (N_8829,N_6920,N_7334);
nand U8830 (N_8830,N_6755,N_6871);
nor U8831 (N_8831,N_7233,N_6999);
or U8832 (N_8832,N_7450,N_7119);
nand U8833 (N_8833,N_6478,N_6750);
nor U8834 (N_8834,N_6964,N_6500);
nand U8835 (N_8835,N_6242,N_7331);
xor U8836 (N_8836,N_7486,N_7007);
or U8837 (N_8837,N_6819,N_6354);
nand U8838 (N_8838,N_7006,N_6334);
or U8839 (N_8839,N_6584,N_6365);
nor U8840 (N_8840,N_7444,N_7238);
nor U8841 (N_8841,N_6013,N_6099);
and U8842 (N_8842,N_6434,N_7150);
xnor U8843 (N_8843,N_6332,N_7086);
and U8844 (N_8844,N_7160,N_6751);
and U8845 (N_8845,N_6274,N_6487);
or U8846 (N_8846,N_6805,N_7370);
nand U8847 (N_8847,N_6955,N_7188);
and U8848 (N_8848,N_6514,N_7180);
or U8849 (N_8849,N_6021,N_7152);
and U8850 (N_8850,N_6957,N_7174);
nor U8851 (N_8851,N_6535,N_6284);
nand U8852 (N_8852,N_7307,N_6048);
or U8853 (N_8853,N_6385,N_6098);
and U8854 (N_8854,N_7390,N_7436);
and U8855 (N_8855,N_6850,N_7136);
nor U8856 (N_8856,N_6895,N_6208);
nand U8857 (N_8857,N_6812,N_6413);
nor U8858 (N_8858,N_6960,N_6178);
and U8859 (N_8859,N_6317,N_6756);
and U8860 (N_8860,N_6478,N_6973);
or U8861 (N_8861,N_6711,N_6151);
nand U8862 (N_8862,N_7274,N_6139);
nor U8863 (N_8863,N_7358,N_6427);
and U8864 (N_8864,N_6769,N_7372);
and U8865 (N_8865,N_6009,N_6704);
nand U8866 (N_8866,N_6217,N_7195);
or U8867 (N_8867,N_7097,N_6703);
nand U8868 (N_8868,N_6897,N_6943);
or U8869 (N_8869,N_7287,N_7061);
nor U8870 (N_8870,N_7108,N_7012);
and U8871 (N_8871,N_6965,N_6981);
or U8872 (N_8872,N_6296,N_6350);
or U8873 (N_8873,N_6709,N_7089);
or U8874 (N_8874,N_7093,N_6566);
nand U8875 (N_8875,N_7134,N_6552);
and U8876 (N_8876,N_6780,N_7223);
or U8877 (N_8877,N_6972,N_7177);
or U8878 (N_8878,N_6193,N_7219);
and U8879 (N_8879,N_6366,N_6390);
nor U8880 (N_8880,N_6830,N_7316);
nor U8881 (N_8881,N_6238,N_6721);
or U8882 (N_8882,N_6293,N_6027);
or U8883 (N_8883,N_6001,N_7490);
nand U8884 (N_8884,N_6434,N_6323);
and U8885 (N_8885,N_6020,N_7036);
or U8886 (N_8886,N_7494,N_7013);
nand U8887 (N_8887,N_6247,N_6522);
and U8888 (N_8888,N_6910,N_6546);
nor U8889 (N_8889,N_6312,N_6426);
or U8890 (N_8890,N_7322,N_6541);
or U8891 (N_8891,N_7138,N_6001);
and U8892 (N_8892,N_6164,N_6287);
nand U8893 (N_8893,N_6211,N_6424);
and U8894 (N_8894,N_6833,N_7363);
nor U8895 (N_8895,N_6085,N_6594);
or U8896 (N_8896,N_7230,N_6310);
nand U8897 (N_8897,N_7392,N_7167);
and U8898 (N_8898,N_6000,N_7292);
nand U8899 (N_8899,N_7261,N_7222);
or U8900 (N_8900,N_7453,N_7488);
and U8901 (N_8901,N_7249,N_6242);
or U8902 (N_8902,N_6708,N_6950);
or U8903 (N_8903,N_6510,N_7429);
nand U8904 (N_8904,N_7067,N_6264);
and U8905 (N_8905,N_6271,N_7467);
and U8906 (N_8906,N_6706,N_7121);
and U8907 (N_8907,N_7292,N_7097);
nand U8908 (N_8908,N_6206,N_6376);
nor U8909 (N_8909,N_7253,N_6139);
nand U8910 (N_8910,N_6225,N_7309);
nor U8911 (N_8911,N_7384,N_7040);
or U8912 (N_8912,N_7186,N_7261);
and U8913 (N_8913,N_6649,N_6848);
nor U8914 (N_8914,N_7020,N_6020);
nor U8915 (N_8915,N_6020,N_6018);
nand U8916 (N_8916,N_6171,N_6302);
nand U8917 (N_8917,N_7212,N_6519);
and U8918 (N_8918,N_6199,N_6499);
and U8919 (N_8919,N_6346,N_6242);
and U8920 (N_8920,N_6684,N_7286);
or U8921 (N_8921,N_6646,N_6174);
xor U8922 (N_8922,N_7369,N_7319);
nor U8923 (N_8923,N_7309,N_6859);
nand U8924 (N_8924,N_7329,N_7416);
or U8925 (N_8925,N_6940,N_6365);
nor U8926 (N_8926,N_6382,N_6939);
and U8927 (N_8927,N_6000,N_7082);
or U8928 (N_8928,N_7368,N_6611);
nor U8929 (N_8929,N_6962,N_7104);
and U8930 (N_8930,N_6084,N_6706);
or U8931 (N_8931,N_6537,N_6187);
and U8932 (N_8932,N_6997,N_6026);
or U8933 (N_8933,N_6945,N_6805);
xor U8934 (N_8934,N_7452,N_6280);
nand U8935 (N_8935,N_6830,N_6852);
nor U8936 (N_8936,N_6085,N_6698);
and U8937 (N_8937,N_7187,N_7162);
nor U8938 (N_8938,N_6459,N_6899);
or U8939 (N_8939,N_6573,N_6176);
nand U8940 (N_8940,N_6397,N_6781);
nand U8941 (N_8941,N_7128,N_7423);
and U8942 (N_8942,N_7062,N_6196);
or U8943 (N_8943,N_6365,N_7339);
nor U8944 (N_8944,N_6655,N_6656);
or U8945 (N_8945,N_7413,N_6041);
nand U8946 (N_8946,N_7031,N_6669);
or U8947 (N_8947,N_6313,N_7315);
nand U8948 (N_8948,N_6014,N_7299);
or U8949 (N_8949,N_7267,N_6276);
or U8950 (N_8950,N_6769,N_6314);
nand U8951 (N_8951,N_6752,N_6002);
nand U8952 (N_8952,N_6934,N_6555);
nor U8953 (N_8953,N_7307,N_6764);
or U8954 (N_8954,N_6052,N_6433);
or U8955 (N_8955,N_6010,N_6603);
and U8956 (N_8956,N_7049,N_6932);
nor U8957 (N_8957,N_6918,N_6289);
or U8958 (N_8958,N_6562,N_6081);
and U8959 (N_8959,N_6475,N_7417);
nor U8960 (N_8960,N_6503,N_7332);
and U8961 (N_8961,N_7038,N_6782);
and U8962 (N_8962,N_6047,N_7246);
or U8963 (N_8963,N_6750,N_7396);
or U8964 (N_8964,N_6390,N_7070);
nand U8965 (N_8965,N_7168,N_7463);
nand U8966 (N_8966,N_7033,N_6113);
or U8967 (N_8967,N_6675,N_6512);
or U8968 (N_8968,N_6862,N_6837);
nand U8969 (N_8969,N_7053,N_6949);
nand U8970 (N_8970,N_6041,N_6293);
and U8971 (N_8971,N_6516,N_7349);
nor U8972 (N_8972,N_6900,N_6682);
and U8973 (N_8973,N_7412,N_6734);
or U8974 (N_8974,N_6616,N_7493);
nor U8975 (N_8975,N_6925,N_6620);
nor U8976 (N_8976,N_6557,N_7105);
or U8977 (N_8977,N_7391,N_6667);
nand U8978 (N_8978,N_6768,N_6874);
or U8979 (N_8979,N_7351,N_6060);
and U8980 (N_8980,N_6541,N_6243);
or U8981 (N_8981,N_6132,N_6016);
and U8982 (N_8982,N_7253,N_6768);
and U8983 (N_8983,N_6889,N_6956);
and U8984 (N_8984,N_6555,N_6748);
nand U8985 (N_8985,N_6467,N_6413);
nor U8986 (N_8986,N_6763,N_6397);
and U8987 (N_8987,N_6232,N_7469);
and U8988 (N_8988,N_6740,N_7353);
or U8989 (N_8989,N_6790,N_6074);
nand U8990 (N_8990,N_7234,N_6827);
and U8991 (N_8991,N_7260,N_7254);
nor U8992 (N_8992,N_6449,N_7310);
and U8993 (N_8993,N_6314,N_7134);
nand U8994 (N_8994,N_6329,N_7346);
or U8995 (N_8995,N_6456,N_6291);
nand U8996 (N_8996,N_6677,N_6281);
and U8997 (N_8997,N_6029,N_6944);
or U8998 (N_8998,N_6714,N_7415);
and U8999 (N_8999,N_6952,N_7345);
or U9000 (N_9000,N_7717,N_7928);
or U9001 (N_9001,N_8828,N_8688);
nand U9002 (N_9002,N_8633,N_7672);
and U9003 (N_9003,N_8477,N_8091);
nand U9004 (N_9004,N_8721,N_7675);
nand U9005 (N_9005,N_7557,N_7660);
nor U9006 (N_9006,N_8664,N_7598);
and U9007 (N_9007,N_7701,N_8755);
or U9008 (N_9008,N_7593,N_8385);
or U9009 (N_9009,N_7524,N_8580);
and U9010 (N_9010,N_8946,N_7694);
xnor U9011 (N_9011,N_7937,N_8445);
or U9012 (N_9012,N_8398,N_7974);
nand U9013 (N_9013,N_8678,N_7778);
and U9014 (N_9014,N_8720,N_7715);
nor U9015 (N_9015,N_7570,N_7682);
nor U9016 (N_9016,N_8594,N_7959);
nand U9017 (N_9017,N_7727,N_8314);
or U9018 (N_9018,N_7765,N_8389);
nand U9019 (N_9019,N_8916,N_8702);
nand U9020 (N_9020,N_7732,N_8951);
nand U9021 (N_9021,N_8456,N_8076);
nor U9022 (N_9022,N_8358,N_7507);
nor U9023 (N_9023,N_8793,N_7637);
and U9024 (N_9024,N_8514,N_8260);
and U9025 (N_9025,N_8166,N_8188);
nand U9026 (N_9026,N_8681,N_8629);
nor U9027 (N_9027,N_8805,N_7877);
nor U9028 (N_9028,N_8247,N_8691);
and U9029 (N_9029,N_8997,N_7806);
xor U9030 (N_9030,N_8203,N_8989);
and U9031 (N_9031,N_8801,N_8868);
and U9032 (N_9032,N_8795,N_7782);
and U9033 (N_9033,N_8264,N_8584);
or U9034 (N_9034,N_7686,N_8438);
nand U9035 (N_9035,N_8854,N_7746);
or U9036 (N_9036,N_8865,N_7638);
and U9037 (N_9037,N_7831,N_7662);
or U9038 (N_9038,N_8948,N_7671);
or U9039 (N_9039,N_8888,N_7670);
or U9040 (N_9040,N_8544,N_7560);
or U9041 (N_9041,N_8243,N_8796);
or U9042 (N_9042,N_8409,N_8446);
nor U9043 (N_9043,N_8448,N_8545);
nand U9044 (N_9044,N_7777,N_8523);
and U9045 (N_9045,N_8839,N_7876);
nand U9046 (N_9046,N_8503,N_7572);
and U9047 (N_9047,N_7601,N_8637);
nor U9048 (N_9048,N_8296,N_8427);
or U9049 (N_9049,N_8936,N_7734);
nor U9050 (N_9050,N_7610,N_7951);
nand U9051 (N_9051,N_7828,N_8950);
and U9052 (N_9052,N_7906,N_8207);
nor U9053 (N_9053,N_8890,N_8275);
or U9054 (N_9054,N_8489,N_8541);
xnor U9055 (N_9055,N_8507,N_8624);
or U9056 (N_9056,N_8288,N_7956);
nand U9057 (N_9057,N_8789,N_8792);
xor U9058 (N_9058,N_7626,N_8769);
and U9059 (N_9059,N_8092,N_8324);
and U9060 (N_9060,N_8454,N_8830);
and U9061 (N_9061,N_7779,N_8869);
or U9062 (N_9062,N_7904,N_8995);
or U9063 (N_9063,N_7833,N_8248);
nand U9064 (N_9064,N_8138,N_8042);
or U9065 (N_9065,N_7995,N_8947);
or U9066 (N_9066,N_8983,N_7647);
and U9067 (N_9067,N_8832,N_7826);
nand U9068 (N_9068,N_8812,N_8778);
and U9069 (N_9069,N_7788,N_7958);
nor U9070 (N_9070,N_8232,N_7905);
nand U9071 (N_9071,N_8718,N_7976);
and U9072 (N_9072,N_7830,N_8053);
or U9073 (N_9073,N_7936,N_8298);
nor U9074 (N_9074,N_7939,N_8016);
nand U9075 (N_9075,N_7564,N_8158);
and U9076 (N_9076,N_7718,N_8791);
nor U9077 (N_9077,N_8128,N_8172);
and U9078 (N_9078,N_8729,N_8988);
or U9079 (N_9079,N_7836,N_7934);
and U9080 (N_9080,N_8597,N_7563);
nor U9081 (N_9081,N_8293,N_8099);
nand U9082 (N_9082,N_8743,N_8312);
nor U9083 (N_9083,N_8899,N_7613);
nand U9084 (N_9084,N_7528,N_7850);
nor U9085 (N_9085,N_8674,N_7907);
or U9086 (N_9086,N_8308,N_7993);
nand U9087 (N_9087,N_8601,N_8177);
or U9088 (N_9088,N_7978,N_8538);
nor U9089 (N_9089,N_7573,N_7886);
nor U9090 (N_9090,N_8018,N_8039);
nand U9091 (N_9091,N_8998,N_8222);
nand U9092 (N_9092,N_7791,N_7699);
nor U9093 (N_9093,N_7733,N_7720);
nand U9094 (N_9094,N_8441,N_7611);
and U9095 (N_9095,N_7621,N_8282);
nand U9096 (N_9096,N_8253,N_7971);
xnor U9097 (N_9097,N_8539,N_8161);
nand U9098 (N_9098,N_7960,N_7918);
or U9099 (N_9099,N_8840,N_7762);
nand U9100 (N_9100,N_8263,N_7986);
nor U9101 (N_9101,N_8551,N_7933);
or U9102 (N_9102,N_8716,N_8131);
nand U9103 (N_9103,N_8414,N_7917);
or U9104 (N_9104,N_8517,N_7988);
nand U9105 (N_9105,N_8698,N_8030);
or U9106 (N_9106,N_8150,N_8440);
and U9107 (N_9107,N_8134,N_8364);
or U9108 (N_9108,N_8707,N_8415);
nor U9109 (N_9109,N_8021,N_7827);
nand U9110 (N_9110,N_8962,N_8422);
or U9111 (N_9111,N_7767,N_7712);
or U9112 (N_9112,N_7596,N_8014);
or U9113 (N_9113,N_7947,N_8818);
and U9114 (N_9114,N_8197,N_8867);
and U9115 (N_9115,N_7711,N_7780);
nor U9116 (N_9116,N_8225,N_8887);
nand U9117 (N_9117,N_7883,N_8349);
or U9118 (N_9118,N_8505,N_7750);
nor U9119 (N_9119,N_8648,N_8802);
and U9120 (N_9120,N_8960,N_7967);
nor U9121 (N_9121,N_8776,N_8547);
and U9122 (N_9122,N_7838,N_8659);
and U9123 (N_9123,N_8245,N_8110);
or U9124 (N_9124,N_8770,N_7758);
and U9125 (N_9125,N_8240,N_8301);
nand U9126 (N_9126,N_7693,N_8763);
nand U9127 (N_9127,N_7808,N_8100);
or U9128 (N_9128,N_8752,N_7914);
nor U9129 (N_9129,N_8094,N_8564);
nand U9130 (N_9130,N_8346,N_8531);
and U9131 (N_9131,N_7798,N_8844);
nor U9132 (N_9132,N_8403,N_7664);
or U9133 (N_9133,N_8910,N_8165);
and U9134 (N_9134,N_8462,N_7603);
or U9135 (N_9135,N_8993,N_7931);
or U9136 (N_9136,N_8286,N_8746);
and U9137 (N_9137,N_8426,N_7789);
or U9138 (N_9138,N_8347,N_8618);
nand U9139 (N_9139,N_8751,N_8089);
xnor U9140 (N_9140,N_7530,N_8004);
or U9141 (N_9141,N_7867,N_8670);
nand U9142 (N_9142,N_7982,N_7639);
or U9143 (N_9143,N_8874,N_8304);
nor U9144 (N_9144,N_8057,N_8749);
nor U9145 (N_9145,N_8327,N_7716);
nor U9146 (N_9146,N_7961,N_8316);
and U9147 (N_9147,N_8259,N_8090);
or U9148 (N_9148,N_8954,N_8406);
or U9149 (N_9149,N_8130,N_8423);
or U9150 (N_9150,N_8373,N_8086);
and U9151 (N_9151,N_8804,N_8405);
and U9152 (N_9152,N_8322,N_8236);
and U9153 (N_9153,N_8493,N_8933);
or U9154 (N_9154,N_8838,N_8764);
and U9155 (N_9155,N_7846,N_8449);
nor U9156 (N_9156,N_7977,N_7805);
nor U9157 (N_9157,N_8725,N_8699);
nand U9158 (N_9158,N_8291,N_8809);
nor U9159 (N_9159,N_7837,N_8783);
nor U9160 (N_9160,N_8816,N_8256);
and U9161 (N_9161,N_8336,N_8550);
and U9162 (N_9162,N_8574,N_7683);
nor U9163 (N_9163,N_7996,N_7745);
or U9164 (N_9164,N_7756,N_8020);
and U9165 (N_9165,N_8905,N_8957);
or U9166 (N_9166,N_7678,N_8156);
and U9167 (N_9167,N_7829,N_7751);
and U9168 (N_9168,N_8155,N_8395);
nor U9169 (N_9169,N_8829,N_8961);
and U9170 (N_9170,N_8118,N_8434);
nor U9171 (N_9171,N_8435,N_7612);
and U9172 (N_9172,N_8619,N_8622);
xnor U9173 (N_9173,N_7901,N_8025);
or U9174 (N_9174,N_8380,N_8964);
or U9175 (N_9175,N_7817,N_7552);
and U9176 (N_9176,N_8515,N_7842);
nand U9177 (N_9177,N_8965,N_7668);
or U9178 (N_9178,N_7633,N_8175);
nor U9179 (N_9179,N_8756,N_8953);
nand U9180 (N_9180,N_8290,N_7900);
nand U9181 (N_9181,N_8891,N_8148);
nor U9182 (N_9182,N_8239,N_7700);
and U9183 (N_9183,N_8062,N_8003);
and U9184 (N_9184,N_7880,N_8596);
or U9185 (N_9185,N_7508,N_8628);
and U9186 (N_9186,N_8252,N_8268);
nand U9187 (N_9187,N_7856,N_8781);
or U9188 (N_9188,N_8602,N_8520);
xnor U9189 (N_9189,N_8595,N_8714);
nor U9190 (N_9190,N_8483,N_7747);
or U9191 (N_9191,N_8083,N_8973);
xnor U9192 (N_9192,N_8902,N_8591);
nand U9193 (N_9193,N_8491,N_8904);
and U9194 (N_9194,N_8051,N_7571);
nand U9195 (N_9195,N_7763,N_7546);
nand U9196 (N_9196,N_8490,N_8536);
nor U9197 (N_9197,N_8318,N_8060);
and U9198 (N_9198,N_8666,N_8433);
or U9199 (N_9199,N_8254,N_8990);
or U9200 (N_9200,N_8966,N_8095);
or U9201 (N_9201,N_8392,N_8579);
or U9202 (N_9202,N_7903,N_8819);
and U9203 (N_9203,N_8853,N_7736);
and U9204 (N_9204,N_7609,N_7955);
nand U9205 (N_9205,N_8706,N_8991);
and U9206 (N_9206,N_8817,N_8534);
nor U9207 (N_9207,N_8696,N_8937);
or U9208 (N_9208,N_8881,N_8354);
nand U9209 (N_9209,N_8238,N_8889);
or U9210 (N_9210,N_8469,N_7814);
and U9211 (N_9211,N_8041,N_8709);
and U9212 (N_9212,N_8001,N_7981);
nor U9213 (N_9213,N_7600,N_8588);
or U9214 (N_9214,N_7743,N_8692);
and U9215 (N_9215,N_7599,N_7871);
nand U9216 (N_9216,N_7659,N_7898);
nor U9217 (N_9217,N_8654,N_8986);
nand U9218 (N_9218,N_8180,N_8310);
nand U9219 (N_9219,N_8339,N_8393);
nand U9220 (N_9220,N_7764,N_8736);
or U9221 (N_9221,N_8122,N_8639);
nor U9222 (N_9222,N_8944,N_8269);
nand U9223 (N_9223,N_8162,N_8636);
nand U9224 (N_9224,N_8072,N_7690);
nand U9225 (N_9225,N_8191,N_8790);
and U9226 (N_9226,N_8450,N_8968);
nor U9227 (N_9227,N_7945,N_7793);
nor U9228 (N_9228,N_8497,N_8082);
and U9229 (N_9229,N_8187,N_8476);
nor U9230 (N_9230,N_8930,N_8333);
nand U9231 (N_9231,N_8183,N_7890);
or U9232 (N_9232,N_8771,N_8416);
and U9233 (N_9233,N_8657,N_8919);
and U9234 (N_9234,N_8583,N_8810);
nand U9235 (N_9235,N_7726,N_8388);
or U9236 (N_9236,N_8821,N_8974);
and U9237 (N_9237,N_8896,N_7766);
nor U9238 (N_9238,N_7991,N_8927);
or U9239 (N_9239,N_7893,N_8443);
nand U9240 (N_9240,N_7769,N_7619);
and U9241 (N_9241,N_8460,N_8012);
or U9242 (N_9242,N_8593,N_8361);
and U9243 (N_9243,N_7516,N_8221);
nor U9244 (N_9244,N_7691,N_8599);
and U9245 (N_9245,N_8151,N_8303);
nor U9246 (N_9246,N_8360,N_8920);
nor U9247 (N_9247,N_8642,N_7569);
nor U9248 (N_9248,N_7790,N_7957);
nand U9249 (N_9249,N_8132,N_8411);
nand U9250 (N_9250,N_7894,N_7994);
and U9251 (N_9251,N_8367,N_7577);
nor U9252 (N_9252,N_8007,N_8143);
or U9253 (N_9253,N_7608,N_8124);
nand U9254 (N_9254,N_8682,N_7964);
nand U9255 (N_9255,N_8938,N_8061);
or U9256 (N_9256,N_8262,N_7781);
nand U9257 (N_9257,N_8017,N_8056);
nor U9258 (N_9258,N_8186,N_7863);
or U9259 (N_9259,N_8578,N_7689);
and U9260 (N_9260,N_7744,N_8685);
nor U9261 (N_9261,N_8949,N_8570);
or U9262 (N_9262,N_8442,N_7812);
nand U9263 (N_9263,N_8885,N_7645);
or U9264 (N_9264,N_7741,N_8608);
or U9265 (N_9265,N_8759,N_8532);
nand U9266 (N_9266,N_8703,N_7587);
nand U9267 (N_9267,N_7655,N_8171);
or U9268 (N_9268,N_8429,N_8350);
or U9269 (N_9269,N_7753,N_8147);
nor U9270 (N_9270,N_8344,N_8571);
or U9271 (N_9271,N_8586,N_8842);
nor U9272 (N_9272,N_8813,N_8480);
or U9273 (N_9273,N_7792,N_8548);
nand U9274 (N_9274,N_8713,N_7872);
nand U9275 (N_9275,N_8472,N_8294);
and U9276 (N_9276,N_7652,N_8560);
or U9277 (N_9277,N_8369,N_8875);
nor U9278 (N_9278,N_8048,N_8641);
and U9279 (N_9279,N_8137,N_8727);
nand U9280 (N_9280,N_7811,N_8022);
nand U9281 (N_9281,N_7553,N_8465);
and U9282 (N_9282,N_7935,N_8750);
or U9283 (N_9283,N_8066,N_7803);
or U9284 (N_9284,N_7580,N_8246);
nor U9285 (N_9285,N_7628,N_8856);
and U9286 (N_9286,N_8765,N_8690);
nor U9287 (N_9287,N_8307,N_7708);
nand U9288 (N_9288,N_8032,N_8033);
and U9289 (N_9289,N_7632,N_8529);
nor U9290 (N_9290,N_7558,N_7707);
nor U9291 (N_9291,N_8391,N_7999);
nor U9292 (N_9292,N_8975,N_7706);
nor U9293 (N_9293,N_8332,N_7604);
and U9294 (N_9294,N_8537,N_8535);
and U9295 (N_9295,N_7650,N_7679);
or U9296 (N_9296,N_8466,N_8215);
nand U9297 (N_9297,N_8087,N_8609);
and U9298 (N_9298,N_8234,N_7921);
nand U9299 (N_9299,N_8357,N_8977);
and U9300 (N_9300,N_8277,N_8058);
and U9301 (N_9301,N_8371,N_7523);
nor U9302 (N_9302,N_7859,N_7926);
and U9303 (N_9303,N_8634,N_8644);
and U9304 (N_9304,N_7940,N_8474);
nand U9305 (N_9305,N_8492,N_8157);
nand U9306 (N_9306,N_8283,N_8194);
nor U9307 (N_9307,N_8375,N_8084);
nor U9308 (N_9308,N_8144,N_8181);
xor U9309 (N_9309,N_8184,N_8273);
nor U9310 (N_9310,N_7759,N_8451);
and U9311 (N_9311,N_8669,N_7949);
nand U9312 (N_9312,N_7797,N_8774);
and U9313 (N_9313,N_8400,N_7556);
nor U9314 (N_9314,N_7550,N_8626);
nor U9315 (N_9315,N_8285,N_8363);
nand U9316 (N_9316,N_8680,N_8141);
or U9317 (N_9317,N_7821,N_8195);
nor U9318 (N_9318,N_8261,N_7695);
nor U9319 (N_9319,N_7506,N_8649);
or U9320 (N_9320,N_8168,N_8811);
nand U9321 (N_9321,N_8733,N_7980);
and U9322 (N_9322,N_8281,N_8705);
or U9323 (N_9323,N_8915,N_8498);
nand U9324 (N_9324,N_7515,N_8035);
nand U9325 (N_9325,N_8331,N_8211);
nand U9326 (N_9326,N_7616,N_8129);
or U9327 (N_9327,N_8127,N_8204);
nor U9328 (N_9328,N_7518,N_8835);
nand U9329 (N_9329,N_8849,N_8009);
and U9330 (N_9330,N_8070,N_8237);
and U9331 (N_9331,N_7924,N_8834);
nor U9332 (N_9332,N_7820,N_7879);
and U9333 (N_9333,N_8573,N_8108);
nand U9334 (N_9334,N_7529,N_7540);
or U9335 (N_9335,N_8911,N_7889);
nand U9336 (N_9336,N_8023,N_7585);
and U9337 (N_9337,N_8464,N_7946);
or U9338 (N_9338,N_8071,N_8803);
and U9339 (N_9339,N_8559,N_7617);
or U9340 (N_9340,N_8824,N_7920);
and U9341 (N_9341,N_8860,N_8971);
and U9342 (N_9342,N_8908,N_7622);
nor U9343 (N_9343,N_8431,N_8098);
nor U9344 (N_9344,N_8745,N_8368);
nand U9345 (N_9345,N_8800,N_8255);
nand U9346 (N_9346,N_7983,N_8552);
or U9347 (N_9347,N_8436,N_7887);
and U9348 (N_9348,N_7627,N_8979);
nand U9349 (N_9349,N_8027,N_8921);
nor U9350 (N_9350,N_7860,N_8043);
or U9351 (N_9351,N_8452,N_8976);
nor U9352 (N_9352,N_8823,N_7899);
or U9353 (N_9353,N_7642,N_7509);
and U9354 (N_9354,N_8748,N_7768);
nor U9355 (N_9355,N_7990,N_7930);
and U9356 (N_9356,N_8967,N_8722);
or U9357 (N_9357,N_8996,N_8107);
or U9358 (N_9358,N_8831,N_7653);
nand U9359 (N_9359,N_8982,N_8463);
nor U9360 (N_9360,N_7688,N_7729);
or U9361 (N_9361,N_7500,N_8723);
or U9362 (N_9362,N_7669,N_7752);
nand U9363 (N_9363,N_8542,N_7888);
and U9364 (N_9364,N_7559,N_7562);
nor U9365 (N_9365,N_8677,N_8216);
nor U9366 (N_9366,N_8069,N_7885);
nor U9367 (N_9367,N_8926,N_7629);
nor U9368 (N_9368,N_7503,N_7548);
or U9369 (N_9369,N_7586,N_7987);
or U9370 (N_9370,N_8825,N_8640);
or U9371 (N_9371,N_7802,N_7950);
nor U9372 (N_9372,N_8555,N_8511);
or U9373 (N_9373,N_7870,N_8121);
nor U9374 (N_9374,N_7667,N_8120);
and U9375 (N_9375,N_8437,N_8126);
nand U9376 (N_9376,N_8064,N_8562);
nand U9377 (N_9377,N_8337,N_8329);
and U9378 (N_9378,N_7938,N_7724);
or U9379 (N_9379,N_8879,N_8687);
or U9380 (N_9380,N_8019,N_8851);
nand U9381 (N_9381,N_8201,N_7684);
nand U9382 (N_9382,N_8683,N_8900);
or U9383 (N_9383,N_7800,N_8173);
nand U9384 (N_9384,N_7922,N_8762);
and U9385 (N_9385,N_8600,N_7687);
and U9386 (N_9386,N_8568,N_7602);
and U9387 (N_9387,N_8617,N_8338);
nand U9388 (N_9388,N_8972,N_8146);
nand U9389 (N_9389,N_8424,N_7635);
nand U9390 (N_9390,N_8567,N_8112);
and U9391 (N_9391,N_8418,N_8390);
nand U9392 (N_9392,N_7835,N_8251);
and U9393 (N_9393,N_8855,N_8111);
or U9394 (N_9394,N_8739,N_8543);
xor U9395 (N_9395,N_7644,N_8665);
and U9396 (N_9396,N_8328,N_8508);
nand U9397 (N_9397,N_8419,N_8113);
nand U9398 (N_9398,N_8178,N_8934);
and U9399 (N_9399,N_8980,N_8724);
and U9400 (N_9400,N_8223,N_8952);
and U9401 (N_9401,N_8199,N_8872);
and U9402 (N_9402,N_7725,N_7641);
and U9403 (N_9403,N_8036,N_8309);
nor U9404 (N_9404,N_8026,N_8413);
nor U9405 (N_9405,N_7545,N_8808);
or U9406 (N_9406,N_8826,N_8969);
nand U9407 (N_9407,N_8566,N_8540);
or U9408 (N_9408,N_8737,N_7630);
and U9409 (N_9409,N_7919,N_8598);
nand U9410 (N_9410,N_7719,N_8708);
or U9411 (N_9411,N_8799,N_7588);
nor U9412 (N_9412,N_8939,N_8340);
and U9413 (N_9413,N_8031,N_8351);
xnor U9414 (N_9414,N_8381,N_8845);
or U9415 (N_9415,N_8067,N_7722);
nor U9416 (N_9416,N_8372,N_8510);
nand U9417 (N_9417,N_8686,N_8894);
and U9418 (N_9418,N_7542,N_8822);
and U9419 (N_9419,N_7501,N_7873);
nand U9420 (N_9420,N_7623,N_8710);
nand U9421 (N_9421,N_8715,N_8097);
nand U9422 (N_9422,N_8123,N_7840);
nand U9423 (N_9423,N_8359,N_7676);
nor U9424 (N_9424,N_7785,N_7698);
and U9425 (N_9425,N_8176,N_8085);
nor U9426 (N_9426,N_7584,N_7582);
or U9427 (N_9427,N_8494,N_8297);
nor U9428 (N_9428,N_8695,N_8650);
and U9429 (N_9429,N_7574,N_7853);
or U9430 (N_9430,N_8228,N_8295);
nand U9431 (N_9431,N_8412,N_8065);
nand U9432 (N_9432,N_8719,N_7576);
and U9433 (N_9433,N_8565,N_7551);
xnor U9434 (N_9434,N_8163,N_7544);
and U9435 (N_9435,N_7998,N_7787);
nand U9436 (N_9436,N_7575,N_8777);
nand U9437 (N_9437,N_8313,N_7902);
nor U9438 (N_9438,N_8028,N_7841);
or U9439 (N_9439,N_8488,N_7985);
or U9440 (N_9440,N_7819,N_7607);
nand U9441 (N_9441,N_7929,N_8645);
or U9442 (N_9442,N_8788,N_8174);
nor U9443 (N_9443,N_8002,N_8738);
nor U9444 (N_9444,N_8487,N_7561);
nor U9445 (N_9445,N_8348,N_7844);
nor U9446 (N_9446,N_7723,N_7851);
nand U9447 (N_9447,N_8052,N_8928);
nor U9448 (N_9448,N_8914,N_8728);
nor U9449 (N_9449,N_8455,N_8500);
nor U9450 (N_9450,N_7892,N_7845);
or U9451 (N_9451,N_7538,N_8942);
nor U9452 (N_9452,N_8658,N_7761);
or U9453 (N_9453,N_7656,N_7896);
and U9454 (N_9454,N_8898,N_7760);
nor U9455 (N_9455,N_7526,N_8563);
nor U9456 (N_9456,N_7874,N_8485);
and U9457 (N_9457,N_7813,N_8320);
nor U9458 (N_9458,N_7786,N_8209);
and U9459 (N_9459,N_8077,N_8153);
or U9460 (N_9460,N_8768,N_7807);
xor U9461 (N_9461,N_7954,N_7620);
nand U9462 (N_9462,N_8079,N_7912);
or U9463 (N_9463,N_7855,N_8940);
or U9464 (N_9464,N_8623,N_8850);
nand U9465 (N_9465,N_7661,N_7923);
and U9466 (N_9466,N_8958,N_7925);
and U9467 (N_9467,N_8558,N_8272);
nor U9468 (N_9468,N_8673,N_7696);
nor U9469 (N_9469,N_8139,N_7738);
nor U9470 (N_9470,N_8913,N_8786);
nor U9471 (N_9471,N_8182,N_8334);
nor U9472 (N_9472,N_7504,N_8766);
and U9473 (N_9473,N_8185,N_8164);
nor U9474 (N_9474,N_8342,N_8206);
and U9475 (N_9475,N_8922,N_8459);
or U9476 (N_9476,N_8675,N_7801);
and U9477 (N_9477,N_8394,N_8661);
nor U9478 (N_9478,N_7615,N_7685);
or U9479 (N_9479,N_8561,N_7631);
nand U9480 (N_9480,N_7776,N_8496);
nor U9481 (N_9481,N_8244,N_7692);
nand U9482 (N_9482,N_7895,N_8994);
or U9483 (N_9483,N_7865,N_8249);
xor U9484 (N_9484,N_8420,N_8046);
or U9485 (N_9485,N_8820,N_8135);
nor U9486 (N_9486,N_7972,N_8689);
and U9487 (N_9487,N_8522,N_7703);
nor U9488 (N_9488,N_8884,N_7713);
nor U9489 (N_9489,N_8352,N_8731);
nand U9490 (N_9490,N_8833,N_8453);
or U9491 (N_9491,N_8909,N_8159);
nand U9492 (N_9492,N_7849,N_8484);
nand U9493 (N_9493,N_8732,N_7625);
nor U9494 (N_9494,N_7513,N_7825);
nor U9495 (N_9495,N_7824,N_8684);
and U9496 (N_9496,N_8284,N_8676);
or U9497 (N_9497,N_8384,N_7681);
nor U9498 (N_9498,N_8606,N_8461);
nor U9499 (N_9499,N_7882,N_7749);
nor U9500 (N_9500,N_8630,N_8401);
or U9501 (N_9501,N_8467,N_8524);
and U9502 (N_9502,N_8073,N_8858);
nor U9503 (N_9503,N_8471,N_7646);
nand U9504 (N_9504,N_7794,N_7772);
and U9505 (N_9505,N_8192,N_8546);
nor U9506 (N_9506,N_8475,N_8585);
nor U9507 (N_9507,N_7735,N_8589);
and U9508 (N_9508,N_8353,N_8005);
xor U9509 (N_9509,N_8343,N_8047);
nand U9510 (N_9510,N_7649,N_8744);
nand U9511 (N_9511,N_8509,N_8773);
or U9512 (N_9512,N_7868,N_8154);
or U9513 (N_9513,N_7783,N_8815);
nand U9514 (N_9514,N_7597,N_8697);
nor U9515 (N_9515,N_8740,N_8444);
nor U9516 (N_9516,N_8499,N_8772);
nand U9517 (N_9517,N_7754,N_7784);
and U9518 (N_9518,N_7680,N_8142);
nand U9519 (N_9519,N_8145,N_8292);
nand U9520 (N_9520,N_7624,N_8863);
nor U9521 (N_9521,N_7737,N_7910);
nand U9522 (N_9522,N_8742,N_8049);
or U9523 (N_9523,N_7665,N_8747);
or U9524 (N_9524,N_8068,N_7531);
or U9525 (N_9525,N_8258,N_7804);
nor U9526 (N_9526,N_8170,N_8037);
and U9527 (N_9527,N_8235,N_8553);
nor U9528 (N_9528,N_8883,N_8906);
or U9529 (N_9529,N_8712,N_8482);
nand U9530 (N_9530,N_8457,N_8470);
or U9531 (N_9531,N_7731,N_8378);
nand U9532 (N_9532,N_8383,N_8149);
and U9533 (N_9533,N_8267,N_8078);
or U9534 (N_9534,N_7966,N_8093);
or U9535 (N_9535,N_7654,N_7677);
and U9536 (N_9536,N_8193,N_8785);
nor U9537 (N_9537,N_8501,N_8700);
or U9538 (N_9538,N_7927,N_8355);
nor U9539 (N_9539,N_8468,N_7710);
nor U9540 (N_9540,N_7963,N_7636);
nand U9541 (N_9541,N_8241,N_8662);
nor U9542 (N_9542,N_7984,N_8101);
xor U9543 (N_9543,N_8323,N_7566);
nand U9544 (N_9544,N_8402,N_8582);
nand U9545 (N_9545,N_7704,N_7852);
and U9546 (N_9546,N_7740,N_8907);
nor U9547 (N_9547,N_8653,N_8878);
nand U9548 (N_9548,N_7875,N_8701);
nor U9549 (N_9549,N_8011,N_7858);
nand U9550 (N_9550,N_8208,N_8923);
or U9551 (N_9551,N_8616,N_8362);
nor U9552 (N_9552,N_8189,N_8169);
nor U9553 (N_9553,N_7555,N_8620);
nand U9554 (N_9554,N_7519,N_8447);
and U9555 (N_9555,N_8784,N_8880);
and U9556 (N_9556,N_7755,N_8886);
and U9557 (N_9557,N_8311,N_8668);
nor U9558 (N_9558,N_8569,N_7714);
nand U9559 (N_9559,N_8133,N_8760);
or U9560 (N_9560,N_8876,N_8230);
and U9561 (N_9561,N_8848,N_8837);
and U9562 (N_9562,N_7997,N_7605);
and U9563 (N_9563,N_7942,N_7522);
and U9564 (N_9564,N_7932,N_8807);
nand U9565 (N_9565,N_7527,N_8397);
nor U9566 (N_9566,N_8300,N_7864);
and U9567 (N_9567,N_8660,N_8655);
or U9568 (N_9568,N_8918,N_8379);
or U9569 (N_9569,N_8912,N_8210);
nand U9570 (N_9570,N_8611,N_7512);
nor U9571 (N_9571,N_8374,N_7857);
or U9572 (N_9572,N_8667,N_7843);
and U9573 (N_9573,N_8321,N_8212);
nand U9574 (N_9574,N_7915,N_8711);
and U9575 (N_9575,N_8603,N_8704);
nor U9576 (N_9576,N_7965,N_8693);
and U9577 (N_9577,N_8512,N_8059);
nor U9578 (N_9578,N_7535,N_7590);
nand U9579 (N_9579,N_7539,N_8767);
or U9580 (N_9580,N_8190,N_8612);
or U9581 (N_9581,N_8631,N_8502);
nand U9582 (N_9582,N_7543,N_7944);
nor U9583 (N_9583,N_8981,N_8119);
xnor U9584 (N_9584,N_7968,N_8717);
or U9585 (N_9585,N_7567,N_8276);
or U9586 (N_9586,N_8365,N_8943);
nor U9587 (N_9587,N_7541,N_8530);
or U9588 (N_9588,N_7774,N_8999);
and U9589 (N_9589,N_8604,N_8278);
and U9590 (N_9590,N_8088,N_8866);
xor U9591 (N_9591,N_7992,N_7823);
or U9592 (N_9592,N_8859,N_8407);
xnor U9593 (N_9593,N_8428,N_7651);
or U9594 (N_9594,N_7657,N_8096);
or U9595 (N_9595,N_8289,N_8115);
and U9596 (N_9596,N_7618,N_8136);
nor U9597 (N_9597,N_8386,N_8315);
nor U9598 (N_9598,N_8495,N_8478);
and U9599 (N_9599,N_8577,N_7909);
or U9600 (N_9600,N_7834,N_7848);
nand U9601 (N_9601,N_7773,N_7952);
nor U9602 (N_9602,N_8104,N_8873);
nor U9603 (N_9603,N_8330,N_8217);
or U9604 (N_9604,N_8008,N_8080);
or U9605 (N_9605,N_7534,N_8109);
or U9606 (N_9606,N_7565,N_8063);
and U9607 (N_9607,N_8125,N_8607);
and U9608 (N_9608,N_7510,N_7948);
nor U9609 (N_9609,N_8615,N_8345);
nor U9610 (N_9610,N_8651,N_8556);
nor U9611 (N_9611,N_7839,N_7606);
nor U9612 (N_9612,N_7878,N_7648);
nand U9613 (N_9613,N_8775,N_8726);
or U9614 (N_9614,N_7969,N_8992);
nand U9615 (N_9615,N_8218,N_8040);
and U9616 (N_9616,N_8554,N_8200);
and U9617 (N_9617,N_7589,N_8935);
nor U9618 (N_9618,N_8399,N_7989);
nor U9619 (N_9619,N_8226,N_8526);
or U9620 (N_9620,N_7818,N_7697);
or U9621 (N_9621,N_8214,N_8054);
and U9622 (N_9622,N_8892,N_8592);
nand U9623 (N_9623,N_8794,N_8882);
and U9624 (N_9624,N_8000,N_8167);
or U9625 (N_9625,N_8549,N_8279);
and U9626 (N_9626,N_8075,N_7891);
or U9627 (N_9627,N_7517,N_8533);
and U9628 (N_9628,N_8335,N_7815);
and U9629 (N_9629,N_8827,N_7854);
nand U9630 (N_9630,N_8116,N_8780);
nor U9631 (N_9631,N_8638,N_8430);
or U9632 (N_9632,N_7869,N_8152);
nand U9633 (N_9633,N_8055,N_8274);
nor U9634 (N_9634,N_8984,N_8179);
and U9635 (N_9635,N_8730,N_7810);
and U9636 (N_9636,N_8787,N_8306);
nor U9637 (N_9637,N_7673,N_8970);
nand U9638 (N_9638,N_8439,N_8233);
nor U9639 (N_9639,N_7549,N_8635);
or U9640 (N_9640,N_8325,N_8857);
and U9641 (N_9641,N_8160,N_8525);
nand U9642 (N_9642,N_8029,N_8924);
or U9643 (N_9643,N_7775,N_7536);
xnor U9644 (N_9644,N_8366,N_8528);
nor U9645 (N_9645,N_7796,N_7666);
nor U9646 (N_9646,N_7757,N_7970);
and U9647 (N_9647,N_8782,N_8106);
or U9648 (N_9648,N_8250,N_7943);
nor U9649 (N_9649,N_8006,N_7916);
nand U9650 (N_9650,N_8224,N_8871);
and U9651 (N_9651,N_8861,N_7640);
or U9652 (N_9652,N_7881,N_8843);
nand U9653 (N_9653,N_8757,N_8231);
and U9654 (N_9654,N_8806,N_7816);
nand U9655 (N_9655,N_8581,N_7847);
nor U9656 (N_9656,N_7705,N_8074);
nor U9657 (N_9657,N_7941,N_7771);
nor U9658 (N_9658,N_8956,N_8643);
nand U9659 (N_9659,N_7643,N_8761);
nor U9660 (N_9660,N_8610,N_8081);
and U9661 (N_9661,N_8798,N_8932);
nor U9662 (N_9662,N_7799,N_8117);
or U9663 (N_9663,N_8613,N_7728);
and U9664 (N_9664,N_8202,N_8326);
and U9665 (N_9665,N_7634,N_7911);
nand U9666 (N_9666,N_8557,N_8925);
or U9667 (N_9667,N_8302,N_8516);
nor U9668 (N_9668,N_7594,N_7595);
nor U9669 (N_9669,N_7514,N_8013);
or U9670 (N_9670,N_8257,N_7739);
and U9671 (N_9671,N_7532,N_8213);
nor U9672 (N_9672,N_7866,N_8299);
nand U9673 (N_9673,N_8852,N_7908);
or U9674 (N_9674,N_8797,N_8387);
and U9675 (N_9675,N_8735,N_8198);
nor U9676 (N_9676,N_8458,N_7742);
and U9677 (N_9677,N_8396,N_7822);
nand U9678 (N_9678,N_7709,N_8196);
nand U9679 (N_9679,N_8102,N_8044);
and U9680 (N_9680,N_8038,N_8265);
nand U9681 (N_9681,N_8877,N_8955);
and U9682 (N_9682,N_8219,N_8382);
or U9683 (N_9683,N_7973,N_7953);
and U9684 (N_9684,N_7581,N_8903);
nor U9685 (N_9685,N_8590,N_8432);
nor U9686 (N_9686,N_8504,N_8572);
and U9687 (N_9687,N_8632,N_8270);
or U9688 (N_9688,N_7975,N_7979);
or U9689 (N_9689,N_8103,N_8621);
and U9690 (N_9690,N_7862,N_8417);
or U9691 (N_9691,N_8753,N_8758);
and U9692 (N_9692,N_8341,N_8656);
or U9693 (N_9693,N_7770,N_7505);
nand U9694 (N_9694,N_8518,N_8671);
nor U9695 (N_9695,N_8741,N_8987);
nand U9696 (N_9696,N_8931,N_7913);
nor U9697 (N_9697,N_7520,N_8870);
or U9698 (N_9698,N_8846,N_7583);
and U9699 (N_9699,N_8527,N_8506);
and U9700 (N_9700,N_8647,N_7511);
nand U9701 (N_9701,N_8754,N_8408);
nor U9702 (N_9702,N_8481,N_8929);
or U9703 (N_9703,N_8024,N_8864);
and U9704 (N_9704,N_8473,N_8679);
or U9705 (N_9705,N_8672,N_8229);
nand U9706 (N_9706,N_8734,N_8814);
nor U9707 (N_9707,N_8513,N_7962);
nor U9708 (N_9708,N_8280,N_8841);
or U9709 (N_9709,N_7525,N_7579);
nand U9710 (N_9710,N_8034,N_7578);
or U9711 (N_9711,N_8317,N_8587);
nand U9712 (N_9712,N_8901,N_8895);
nand U9713 (N_9713,N_8897,N_8862);
nand U9714 (N_9714,N_8893,N_8114);
and U9715 (N_9715,N_8356,N_7658);
nor U9716 (N_9716,N_8486,N_8266);
and U9717 (N_9717,N_8521,N_7674);
nand U9718 (N_9718,N_7533,N_8627);
nand U9719 (N_9719,N_7663,N_8242);
and U9720 (N_9720,N_8963,N_8694);
nand U9721 (N_9721,N_8421,N_8287);
and U9722 (N_9722,N_8978,N_8410);
or U9723 (N_9723,N_8519,N_7521);
and U9724 (N_9724,N_7884,N_7702);
xnor U9725 (N_9725,N_8663,N_8941);
and U9726 (N_9726,N_8575,N_8050);
and U9727 (N_9727,N_7809,N_7748);
xor U9728 (N_9728,N_8305,N_8479);
and U9729 (N_9729,N_8646,N_7547);
nor U9730 (N_9730,N_8404,N_7897);
nor U9731 (N_9731,N_7832,N_8959);
and U9732 (N_9732,N_8605,N_8220);
xnor U9733 (N_9733,N_8945,N_8652);
nand U9734 (N_9734,N_8779,N_8205);
nor U9735 (N_9735,N_8377,N_7592);
nand U9736 (N_9736,N_7861,N_8045);
nor U9737 (N_9737,N_8015,N_8227);
nor U9738 (N_9738,N_7568,N_8614);
and U9739 (N_9739,N_8370,N_8625);
and U9740 (N_9740,N_8105,N_8425);
nor U9741 (N_9741,N_8836,N_8271);
and U9742 (N_9742,N_7721,N_8140);
nor U9743 (N_9743,N_8917,N_7502);
and U9744 (N_9744,N_8847,N_8576);
nor U9745 (N_9745,N_8985,N_7730);
or U9746 (N_9746,N_8319,N_7614);
and U9747 (N_9747,N_7591,N_7554);
nand U9748 (N_9748,N_7795,N_8376);
or U9749 (N_9749,N_8010,N_7537);
and U9750 (N_9750,N_8115,N_8420);
nand U9751 (N_9751,N_8854,N_8899);
and U9752 (N_9752,N_8422,N_8717);
nor U9753 (N_9753,N_7613,N_7615);
or U9754 (N_9754,N_7884,N_7789);
nand U9755 (N_9755,N_8624,N_8917);
nor U9756 (N_9756,N_8237,N_7733);
or U9757 (N_9757,N_7957,N_7817);
nand U9758 (N_9758,N_8723,N_8876);
or U9759 (N_9759,N_8577,N_8632);
or U9760 (N_9760,N_8537,N_7918);
nor U9761 (N_9761,N_8180,N_7791);
and U9762 (N_9762,N_8685,N_8058);
or U9763 (N_9763,N_7554,N_8240);
nor U9764 (N_9764,N_8043,N_8548);
and U9765 (N_9765,N_8342,N_7984);
or U9766 (N_9766,N_8046,N_7544);
or U9767 (N_9767,N_8015,N_8343);
nor U9768 (N_9768,N_7797,N_8046);
nand U9769 (N_9769,N_8809,N_8089);
nand U9770 (N_9770,N_8175,N_8201);
nor U9771 (N_9771,N_8235,N_7505);
nor U9772 (N_9772,N_8851,N_8776);
or U9773 (N_9773,N_8599,N_8953);
and U9774 (N_9774,N_8628,N_7815);
nor U9775 (N_9775,N_8531,N_8891);
or U9776 (N_9776,N_8179,N_8790);
and U9777 (N_9777,N_7912,N_8473);
or U9778 (N_9778,N_8681,N_8588);
xor U9779 (N_9779,N_8847,N_8990);
and U9780 (N_9780,N_8240,N_8988);
nand U9781 (N_9781,N_7529,N_8322);
nand U9782 (N_9782,N_8853,N_8258);
nand U9783 (N_9783,N_8247,N_7761);
nor U9784 (N_9784,N_8005,N_8637);
and U9785 (N_9785,N_8750,N_8370);
or U9786 (N_9786,N_8087,N_8919);
nor U9787 (N_9787,N_8027,N_7622);
nor U9788 (N_9788,N_8863,N_7599);
nand U9789 (N_9789,N_7711,N_8331);
and U9790 (N_9790,N_7768,N_7543);
nor U9791 (N_9791,N_8894,N_7596);
and U9792 (N_9792,N_7839,N_7966);
or U9793 (N_9793,N_7606,N_7646);
nand U9794 (N_9794,N_8125,N_8662);
nor U9795 (N_9795,N_8526,N_8081);
nor U9796 (N_9796,N_7705,N_8054);
nor U9797 (N_9797,N_7539,N_8869);
or U9798 (N_9798,N_7832,N_8574);
and U9799 (N_9799,N_8431,N_8444);
nand U9800 (N_9800,N_8120,N_7505);
or U9801 (N_9801,N_8474,N_7702);
and U9802 (N_9802,N_8799,N_7690);
nand U9803 (N_9803,N_8952,N_8465);
nor U9804 (N_9804,N_8727,N_8387);
or U9805 (N_9805,N_8724,N_8761);
nor U9806 (N_9806,N_8503,N_7748);
nor U9807 (N_9807,N_8415,N_8939);
or U9808 (N_9808,N_8710,N_8241);
nor U9809 (N_9809,N_8871,N_8483);
and U9810 (N_9810,N_8499,N_7674);
nor U9811 (N_9811,N_8952,N_8225);
nor U9812 (N_9812,N_8029,N_7827);
nand U9813 (N_9813,N_7879,N_8805);
and U9814 (N_9814,N_7781,N_7796);
nand U9815 (N_9815,N_8627,N_8462);
or U9816 (N_9816,N_8616,N_8565);
nand U9817 (N_9817,N_8625,N_7539);
nand U9818 (N_9818,N_7566,N_7934);
and U9819 (N_9819,N_8498,N_8842);
nand U9820 (N_9820,N_8206,N_7587);
or U9821 (N_9821,N_8420,N_7695);
nor U9822 (N_9822,N_8660,N_8019);
or U9823 (N_9823,N_8403,N_8230);
or U9824 (N_9824,N_7658,N_8294);
and U9825 (N_9825,N_8443,N_7815);
and U9826 (N_9826,N_8418,N_8153);
nor U9827 (N_9827,N_8154,N_8816);
and U9828 (N_9828,N_8479,N_7981);
or U9829 (N_9829,N_8840,N_8573);
nor U9830 (N_9830,N_8456,N_7581);
xor U9831 (N_9831,N_7651,N_8384);
and U9832 (N_9832,N_8500,N_7526);
nor U9833 (N_9833,N_8880,N_7694);
nor U9834 (N_9834,N_8070,N_8147);
nor U9835 (N_9835,N_8278,N_7743);
or U9836 (N_9836,N_8958,N_8494);
nor U9837 (N_9837,N_8088,N_7920);
or U9838 (N_9838,N_7915,N_8255);
nand U9839 (N_9839,N_7745,N_7785);
nor U9840 (N_9840,N_8177,N_8497);
nor U9841 (N_9841,N_8976,N_7559);
and U9842 (N_9842,N_8194,N_8097);
and U9843 (N_9843,N_7872,N_7629);
nor U9844 (N_9844,N_7865,N_7651);
nor U9845 (N_9845,N_8961,N_8499);
nand U9846 (N_9846,N_8339,N_8211);
nand U9847 (N_9847,N_7722,N_7715);
or U9848 (N_9848,N_8063,N_8382);
nand U9849 (N_9849,N_8321,N_8367);
and U9850 (N_9850,N_8296,N_7696);
nor U9851 (N_9851,N_8008,N_8711);
nand U9852 (N_9852,N_7826,N_8371);
nor U9853 (N_9853,N_8016,N_8950);
nand U9854 (N_9854,N_8852,N_8409);
nor U9855 (N_9855,N_8392,N_8504);
or U9856 (N_9856,N_7853,N_8773);
and U9857 (N_9857,N_8020,N_8029);
or U9858 (N_9858,N_8818,N_8534);
nor U9859 (N_9859,N_8489,N_7540);
and U9860 (N_9860,N_7918,N_8976);
and U9861 (N_9861,N_8245,N_7969);
and U9862 (N_9862,N_8420,N_8769);
nand U9863 (N_9863,N_8302,N_8387);
nor U9864 (N_9864,N_7764,N_7536);
or U9865 (N_9865,N_7583,N_7786);
or U9866 (N_9866,N_7819,N_7647);
or U9867 (N_9867,N_7785,N_7541);
nor U9868 (N_9868,N_8568,N_7697);
nand U9869 (N_9869,N_8846,N_8557);
and U9870 (N_9870,N_8712,N_8974);
or U9871 (N_9871,N_8833,N_7898);
nand U9872 (N_9872,N_7887,N_8054);
nor U9873 (N_9873,N_7941,N_8285);
or U9874 (N_9874,N_7530,N_8555);
or U9875 (N_9875,N_8705,N_7868);
nor U9876 (N_9876,N_8606,N_8095);
nor U9877 (N_9877,N_8971,N_7969);
or U9878 (N_9878,N_8473,N_8884);
or U9879 (N_9879,N_8081,N_8312);
or U9880 (N_9880,N_7536,N_8238);
or U9881 (N_9881,N_8039,N_7737);
nor U9882 (N_9882,N_8797,N_8643);
nor U9883 (N_9883,N_7654,N_7556);
or U9884 (N_9884,N_8182,N_8292);
nand U9885 (N_9885,N_8051,N_8607);
or U9886 (N_9886,N_8654,N_8554);
and U9887 (N_9887,N_7977,N_8918);
nand U9888 (N_9888,N_8746,N_8127);
nand U9889 (N_9889,N_8303,N_8737);
and U9890 (N_9890,N_7595,N_8154);
nor U9891 (N_9891,N_7965,N_7702);
or U9892 (N_9892,N_7555,N_8531);
or U9893 (N_9893,N_8635,N_7679);
nor U9894 (N_9894,N_8614,N_7680);
and U9895 (N_9895,N_8341,N_8393);
nand U9896 (N_9896,N_7817,N_8352);
nand U9897 (N_9897,N_7675,N_8580);
nand U9898 (N_9898,N_8682,N_8377);
or U9899 (N_9899,N_8758,N_8796);
or U9900 (N_9900,N_8578,N_8883);
and U9901 (N_9901,N_8901,N_7993);
nand U9902 (N_9902,N_8069,N_8667);
or U9903 (N_9903,N_8557,N_7796);
nand U9904 (N_9904,N_8571,N_8740);
nand U9905 (N_9905,N_8783,N_7510);
nor U9906 (N_9906,N_8094,N_7618);
and U9907 (N_9907,N_8673,N_7785);
or U9908 (N_9908,N_8005,N_8218);
nand U9909 (N_9909,N_7890,N_8380);
or U9910 (N_9910,N_8261,N_8891);
or U9911 (N_9911,N_7646,N_8917);
or U9912 (N_9912,N_8015,N_8071);
or U9913 (N_9913,N_8698,N_8024);
nand U9914 (N_9914,N_8050,N_8355);
nand U9915 (N_9915,N_8769,N_7893);
nor U9916 (N_9916,N_8088,N_8106);
and U9917 (N_9917,N_8598,N_8269);
nor U9918 (N_9918,N_7687,N_8583);
and U9919 (N_9919,N_8229,N_8315);
or U9920 (N_9920,N_7934,N_8075);
nand U9921 (N_9921,N_8697,N_8807);
or U9922 (N_9922,N_8909,N_8816);
and U9923 (N_9923,N_8997,N_7684);
nand U9924 (N_9924,N_8101,N_8745);
nand U9925 (N_9925,N_8338,N_8183);
nor U9926 (N_9926,N_7529,N_8885);
or U9927 (N_9927,N_7738,N_7646);
or U9928 (N_9928,N_8404,N_8555);
and U9929 (N_9929,N_7606,N_7523);
and U9930 (N_9930,N_8322,N_8203);
nand U9931 (N_9931,N_8293,N_7799);
or U9932 (N_9932,N_8650,N_7858);
and U9933 (N_9933,N_8465,N_8369);
and U9934 (N_9934,N_8284,N_8486);
nand U9935 (N_9935,N_7648,N_8896);
nor U9936 (N_9936,N_8641,N_7576);
nand U9937 (N_9937,N_8221,N_8360);
nand U9938 (N_9938,N_8740,N_8362);
and U9939 (N_9939,N_7876,N_8009);
nand U9940 (N_9940,N_8788,N_7614);
or U9941 (N_9941,N_8404,N_7741);
and U9942 (N_9942,N_8916,N_8817);
nor U9943 (N_9943,N_7841,N_8733);
or U9944 (N_9944,N_7645,N_8461);
nand U9945 (N_9945,N_8784,N_8467);
and U9946 (N_9946,N_8330,N_7570);
nor U9947 (N_9947,N_8885,N_7725);
nor U9948 (N_9948,N_8948,N_7625);
or U9949 (N_9949,N_8728,N_8261);
or U9950 (N_9950,N_8588,N_8754);
or U9951 (N_9951,N_8644,N_8226);
nor U9952 (N_9952,N_8400,N_8326);
and U9953 (N_9953,N_8979,N_7780);
or U9954 (N_9954,N_7758,N_8905);
nor U9955 (N_9955,N_8404,N_8736);
and U9956 (N_9956,N_7868,N_7830);
or U9957 (N_9957,N_7516,N_8048);
or U9958 (N_9958,N_8157,N_8318);
nor U9959 (N_9959,N_8118,N_8159);
and U9960 (N_9960,N_7636,N_8995);
nor U9961 (N_9961,N_7620,N_8565);
xnor U9962 (N_9962,N_7906,N_8691);
or U9963 (N_9963,N_8572,N_8175);
nand U9964 (N_9964,N_7914,N_7735);
nand U9965 (N_9965,N_8790,N_8638);
nand U9966 (N_9966,N_8194,N_8675);
xor U9967 (N_9967,N_7551,N_8394);
nor U9968 (N_9968,N_8277,N_8164);
and U9969 (N_9969,N_7525,N_8804);
and U9970 (N_9970,N_8612,N_8306);
nand U9971 (N_9971,N_8719,N_8058);
and U9972 (N_9972,N_8390,N_8204);
or U9973 (N_9973,N_7807,N_8167);
or U9974 (N_9974,N_7897,N_8348);
and U9975 (N_9975,N_8667,N_7604);
nand U9976 (N_9976,N_7620,N_8681);
or U9977 (N_9977,N_7618,N_8633);
or U9978 (N_9978,N_8037,N_8798);
nor U9979 (N_9979,N_7636,N_7515);
nand U9980 (N_9980,N_8091,N_8478);
nor U9981 (N_9981,N_8101,N_8726);
or U9982 (N_9982,N_7904,N_7536);
nand U9983 (N_9983,N_7519,N_8225);
nor U9984 (N_9984,N_7666,N_8668);
nor U9985 (N_9985,N_7685,N_7894);
nand U9986 (N_9986,N_8631,N_7734);
or U9987 (N_9987,N_7888,N_7565);
nand U9988 (N_9988,N_8299,N_8447);
nor U9989 (N_9989,N_7551,N_8270);
nor U9990 (N_9990,N_7681,N_8555);
nand U9991 (N_9991,N_7504,N_7741);
nand U9992 (N_9992,N_7975,N_8238);
nor U9993 (N_9993,N_8652,N_8413);
nor U9994 (N_9994,N_8260,N_8772);
nor U9995 (N_9995,N_8935,N_8811);
or U9996 (N_9996,N_7577,N_8780);
nor U9997 (N_9997,N_8357,N_8020);
nor U9998 (N_9998,N_8106,N_8431);
nand U9999 (N_9999,N_8946,N_8954);
and U10000 (N_10000,N_8106,N_7817);
or U10001 (N_10001,N_7662,N_8540);
or U10002 (N_10002,N_7813,N_8259);
or U10003 (N_10003,N_8277,N_7662);
nand U10004 (N_10004,N_8018,N_8252);
or U10005 (N_10005,N_7730,N_8940);
nand U10006 (N_10006,N_8414,N_8087);
nor U10007 (N_10007,N_8521,N_7992);
nor U10008 (N_10008,N_7740,N_7743);
and U10009 (N_10009,N_8300,N_7545);
or U10010 (N_10010,N_7891,N_8566);
and U10011 (N_10011,N_8013,N_7657);
or U10012 (N_10012,N_8596,N_8969);
nor U10013 (N_10013,N_8349,N_7877);
nand U10014 (N_10014,N_8977,N_8788);
nand U10015 (N_10015,N_7685,N_8791);
nor U10016 (N_10016,N_8268,N_7773);
or U10017 (N_10017,N_7896,N_7804);
nand U10018 (N_10018,N_8007,N_8543);
and U10019 (N_10019,N_7773,N_8889);
nor U10020 (N_10020,N_8314,N_8978);
or U10021 (N_10021,N_8853,N_7845);
and U10022 (N_10022,N_8050,N_8847);
nand U10023 (N_10023,N_8971,N_8153);
and U10024 (N_10024,N_8950,N_8855);
or U10025 (N_10025,N_8902,N_8326);
or U10026 (N_10026,N_8149,N_7502);
or U10027 (N_10027,N_7566,N_8392);
or U10028 (N_10028,N_8095,N_7659);
and U10029 (N_10029,N_8521,N_7922);
or U10030 (N_10030,N_7829,N_7763);
nand U10031 (N_10031,N_8169,N_7621);
nand U10032 (N_10032,N_7947,N_7502);
nor U10033 (N_10033,N_8693,N_8209);
or U10034 (N_10034,N_8008,N_7791);
nand U10035 (N_10035,N_8293,N_8976);
or U10036 (N_10036,N_8737,N_8500);
nand U10037 (N_10037,N_7744,N_7997);
and U10038 (N_10038,N_7710,N_8524);
nor U10039 (N_10039,N_7811,N_8424);
and U10040 (N_10040,N_7892,N_8779);
nor U10041 (N_10041,N_8715,N_8428);
nor U10042 (N_10042,N_8390,N_8937);
nor U10043 (N_10043,N_7992,N_7504);
or U10044 (N_10044,N_8760,N_8870);
and U10045 (N_10045,N_8715,N_8270);
and U10046 (N_10046,N_7855,N_8495);
nand U10047 (N_10047,N_8874,N_8934);
nor U10048 (N_10048,N_7923,N_7503);
nor U10049 (N_10049,N_7611,N_8570);
nand U10050 (N_10050,N_8913,N_8781);
or U10051 (N_10051,N_7984,N_8319);
and U10052 (N_10052,N_7814,N_7775);
nor U10053 (N_10053,N_8694,N_8013);
and U10054 (N_10054,N_8831,N_7804);
nor U10055 (N_10055,N_8541,N_7624);
or U10056 (N_10056,N_7771,N_7571);
or U10057 (N_10057,N_7985,N_7678);
nor U10058 (N_10058,N_7904,N_8817);
or U10059 (N_10059,N_8350,N_7753);
nor U10060 (N_10060,N_7572,N_8957);
nor U10061 (N_10061,N_8254,N_7837);
nand U10062 (N_10062,N_8379,N_8477);
nand U10063 (N_10063,N_7880,N_8643);
or U10064 (N_10064,N_7786,N_8674);
nor U10065 (N_10065,N_8343,N_7993);
or U10066 (N_10066,N_8413,N_8483);
and U10067 (N_10067,N_8670,N_8199);
nand U10068 (N_10068,N_8722,N_8650);
nand U10069 (N_10069,N_8060,N_8494);
nor U10070 (N_10070,N_7781,N_8440);
and U10071 (N_10071,N_7786,N_8480);
or U10072 (N_10072,N_8906,N_8310);
or U10073 (N_10073,N_8363,N_7756);
nor U10074 (N_10074,N_8340,N_8893);
and U10075 (N_10075,N_7934,N_7888);
nor U10076 (N_10076,N_8110,N_8982);
or U10077 (N_10077,N_8940,N_8166);
nor U10078 (N_10078,N_7925,N_8533);
nand U10079 (N_10079,N_8082,N_8893);
xnor U10080 (N_10080,N_7575,N_7827);
or U10081 (N_10081,N_8222,N_8182);
and U10082 (N_10082,N_7800,N_7515);
nor U10083 (N_10083,N_8843,N_7536);
nor U10084 (N_10084,N_7672,N_8095);
nor U10085 (N_10085,N_7687,N_7995);
and U10086 (N_10086,N_8335,N_7532);
nand U10087 (N_10087,N_8711,N_8266);
and U10088 (N_10088,N_7740,N_8665);
nor U10089 (N_10089,N_7696,N_8009);
nand U10090 (N_10090,N_8843,N_8492);
nor U10091 (N_10091,N_8057,N_7881);
and U10092 (N_10092,N_7930,N_8224);
nor U10093 (N_10093,N_8854,N_8738);
nand U10094 (N_10094,N_8418,N_8299);
or U10095 (N_10095,N_8168,N_8184);
and U10096 (N_10096,N_8858,N_8965);
nand U10097 (N_10097,N_7823,N_7952);
nor U10098 (N_10098,N_8844,N_8449);
nor U10099 (N_10099,N_8274,N_8703);
and U10100 (N_10100,N_8120,N_8096);
nand U10101 (N_10101,N_8966,N_7540);
or U10102 (N_10102,N_8854,N_7865);
nor U10103 (N_10103,N_8854,N_8747);
nor U10104 (N_10104,N_7967,N_7577);
nor U10105 (N_10105,N_7789,N_7972);
nor U10106 (N_10106,N_8328,N_8042);
nor U10107 (N_10107,N_7635,N_8584);
nor U10108 (N_10108,N_8837,N_8550);
and U10109 (N_10109,N_8010,N_7692);
or U10110 (N_10110,N_8810,N_7527);
nor U10111 (N_10111,N_8083,N_8571);
nor U10112 (N_10112,N_7986,N_8302);
nor U10113 (N_10113,N_7662,N_8058);
nor U10114 (N_10114,N_7910,N_7639);
nand U10115 (N_10115,N_8062,N_8024);
nand U10116 (N_10116,N_8356,N_7824);
nand U10117 (N_10117,N_7999,N_7759);
or U10118 (N_10118,N_8481,N_7518);
or U10119 (N_10119,N_8380,N_8032);
or U10120 (N_10120,N_8667,N_8847);
nand U10121 (N_10121,N_8752,N_7545);
or U10122 (N_10122,N_8805,N_8236);
nor U10123 (N_10123,N_8593,N_8776);
nor U10124 (N_10124,N_7716,N_8424);
and U10125 (N_10125,N_8403,N_8369);
or U10126 (N_10126,N_8536,N_7663);
and U10127 (N_10127,N_7830,N_8097);
nor U10128 (N_10128,N_8840,N_7782);
xnor U10129 (N_10129,N_7635,N_8171);
nor U10130 (N_10130,N_7848,N_7707);
nand U10131 (N_10131,N_8697,N_8770);
and U10132 (N_10132,N_7883,N_8162);
and U10133 (N_10133,N_8680,N_8770);
nand U10134 (N_10134,N_8035,N_8260);
nor U10135 (N_10135,N_7821,N_7685);
nand U10136 (N_10136,N_8131,N_8332);
nor U10137 (N_10137,N_8828,N_7768);
nor U10138 (N_10138,N_7531,N_8752);
or U10139 (N_10139,N_8572,N_8474);
nand U10140 (N_10140,N_8964,N_8645);
and U10141 (N_10141,N_8921,N_8124);
nand U10142 (N_10142,N_8640,N_8623);
and U10143 (N_10143,N_7994,N_7584);
nand U10144 (N_10144,N_8547,N_7830);
nor U10145 (N_10145,N_7799,N_8175);
or U10146 (N_10146,N_7763,N_8912);
or U10147 (N_10147,N_8069,N_8738);
xor U10148 (N_10148,N_8789,N_8287);
and U10149 (N_10149,N_8140,N_8431);
nand U10150 (N_10150,N_8993,N_8476);
and U10151 (N_10151,N_8973,N_8211);
and U10152 (N_10152,N_8132,N_7893);
or U10153 (N_10153,N_8304,N_8733);
and U10154 (N_10154,N_8253,N_7500);
nand U10155 (N_10155,N_7803,N_8488);
nand U10156 (N_10156,N_8680,N_8415);
nor U10157 (N_10157,N_8466,N_8795);
nand U10158 (N_10158,N_7976,N_8852);
nand U10159 (N_10159,N_7701,N_8057);
or U10160 (N_10160,N_8470,N_8923);
nor U10161 (N_10161,N_7537,N_8012);
nand U10162 (N_10162,N_8244,N_7561);
nor U10163 (N_10163,N_8462,N_8543);
or U10164 (N_10164,N_7790,N_8287);
nand U10165 (N_10165,N_8331,N_7634);
xnor U10166 (N_10166,N_8896,N_8495);
nor U10167 (N_10167,N_8220,N_8498);
nor U10168 (N_10168,N_7697,N_7906);
or U10169 (N_10169,N_8328,N_7966);
and U10170 (N_10170,N_8795,N_8147);
or U10171 (N_10171,N_7604,N_8829);
and U10172 (N_10172,N_7815,N_7889);
and U10173 (N_10173,N_8721,N_8269);
and U10174 (N_10174,N_7870,N_8181);
nand U10175 (N_10175,N_8830,N_8373);
or U10176 (N_10176,N_8110,N_8957);
or U10177 (N_10177,N_8226,N_7901);
and U10178 (N_10178,N_8595,N_8118);
or U10179 (N_10179,N_8675,N_8972);
and U10180 (N_10180,N_8688,N_8747);
and U10181 (N_10181,N_8736,N_8599);
nand U10182 (N_10182,N_8824,N_8021);
or U10183 (N_10183,N_7668,N_8312);
and U10184 (N_10184,N_8989,N_7821);
nor U10185 (N_10185,N_8668,N_8038);
and U10186 (N_10186,N_7675,N_7810);
and U10187 (N_10187,N_7670,N_7764);
nand U10188 (N_10188,N_7580,N_8996);
and U10189 (N_10189,N_8409,N_7817);
nor U10190 (N_10190,N_7718,N_7766);
or U10191 (N_10191,N_7843,N_8175);
and U10192 (N_10192,N_8219,N_8178);
or U10193 (N_10193,N_7690,N_7731);
nand U10194 (N_10194,N_8058,N_8091);
nand U10195 (N_10195,N_8876,N_7806);
and U10196 (N_10196,N_8319,N_7978);
or U10197 (N_10197,N_8650,N_8503);
or U10198 (N_10198,N_7596,N_8638);
nand U10199 (N_10199,N_7645,N_8929);
and U10200 (N_10200,N_8560,N_8167);
nand U10201 (N_10201,N_7564,N_8321);
nor U10202 (N_10202,N_7720,N_7961);
and U10203 (N_10203,N_7839,N_8154);
or U10204 (N_10204,N_8197,N_7621);
nand U10205 (N_10205,N_7952,N_8663);
or U10206 (N_10206,N_8079,N_7761);
or U10207 (N_10207,N_8878,N_8511);
or U10208 (N_10208,N_7770,N_8612);
and U10209 (N_10209,N_8135,N_8023);
or U10210 (N_10210,N_8443,N_7747);
nand U10211 (N_10211,N_8290,N_8477);
and U10212 (N_10212,N_7748,N_8810);
and U10213 (N_10213,N_8761,N_8912);
and U10214 (N_10214,N_8158,N_8876);
nor U10215 (N_10215,N_8121,N_8266);
nor U10216 (N_10216,N_8791,N_7603);
or U10217 (N_10217,N_8274,N_8454);
and U10218 (N_10218,N_7977,N_8564);
nand U10219 (N_10219,N_8734,N_7576);
and U10220 (N_10220,N_7880,N_8511);
or U10221 (N_10221,N_8704,N_7703);
nand U10222 (N_10222,N_8442,N_8478);
or U10223 (N_10223,N_7684,N_7924);
nand U10224 (N_10224,N_8672,N_8763);
nand U10225 (N_10225,N_8788,N_7598);
nand U10226 (N_10226,N_8948,N_8432);
and U10227 (N_10227,N_8524,N_8391);
nor U10228 (N_10228,N_7800,N_7654);
nand U10229 (N_10229,N_7971,N_7938);
nor U10230 (N_10230,N_7815,N_8393);
and U10231 (N_10231,N_8553,N_8436);
and U10232 (N_10232,N_7781,N_7609);
nand U10233 (N_10233,N_8383,N_7971);
or U10234 (N_10234,N_7832,N_8819);
nand U10235 (N_10235,N_7660,N_8647);
nor U10236 (N_10236,N_7833,N_8833);
nand U10237 (N_10237,N_8805,N_8960);
nand U10238 (N_10238,N_7818,N_7588);
or U10239 (N_10239,N_8810,N_8425);
or U10240 (N_10240,N_8893,N_7885);
and U10241 (N_10241,N_8606,N_8778);
nor U10242 (N_10242,N_8834,N_8645);
nor U10243 (N_10243,N_7506,N_8679);
nor U10244 (N_10244,N_8815,N_8564);
nor U10245 (N_10245,N_8902,N_8559);
nor U10246 (N_10246,N_8180,N_8090);
or U10247 (N_10247,N_8817,N_7947);
or U10248 (N_10248,N_7561,N_8965);
or U10249 (N_10249,N_8192,N_8423);
nand U10250 (N_10250,N_8767,N_7975);
and U10251 (N_10251,N_8577,N_7947);
or U10252 (N_10252,N_8054,N_8286);
and U10253 (N_10253,N_7982,N_8706);
and U10254 (N_10254,N_7868,N_8422);
nand U10255 (N_10255,N_7819,N_7960);
or U10256 (N_10256,N_8467,N_7650);
or U10257 (N_10257,N_8991,N_7925);
and U10258 (N_10258,N_7791,N_7548);
nor U10259 (N_10259,N_8072,N_8894);
nand U10260 (N_10260,N_7564,N_7688);
nor U10261 (N_10261,N_8081,N_8865);
nand U10262 (N_10262,N_7665,N_8045);
and U10263 (N_10263,N_7979,N_8950);
nor U10264 (N_10264,N_8310,N_7584);
nor U10265 (N_10265,N_8710,N_8074);
and U10266 (N_10266,N_7635,N_8062);
and U10267 (N_10267,N_8708,N_8616);
and U10268 (N_10268,N_8070,N_8839);
nor U10269 (N_10269,N_8343,N_8613);
and U10270 (N_10270,N_8030,N_7715);
or U10271 (N_10271,N_8567,N_7624);
nor U10272 (N_10272,N_7820,N_8961);
or U10273 (N_10273,N_7545,N_8637);
and U10274 (N_10274,N_8818,N_7830);
and U10275 (N_10275,N_8308,N_8562);
nand U10276 (N_10276,N_8618,N_7733);
nand U10277 (N_10277,N_8329,N_8392);
and U10278 (N_10278,N_8798,N_8450);
nand U10279 (N_10279,N_8550,N_7734);
and U10280 (N_10280,N_8735,N_8450);
nor U10281 (N_10281,N_8108,N_8190);
and U10282 (N_10282,N_7665,N_8919);
nand U10283 (N_10283,N_8140,N_7736);
nand U10284 (N_10284,N_8114,N_8269);
nand U10285 (N_10285,N_8628,N_8178);
nand U10286 (N_10286,N_8254,N_8335);
xor U10287 (N_10287,N_7641,N_8499);
and U10288 (N_10288,N_8860,N_8585);
nor U10289 (N_10289,N_8303,N_8258);
or U10290 (N_10290,N_8126,N_8402);
or U10291 (N_10291,N_8629,N_7972);
nor U10292 (N_10292,N_7837,N_7936);
and U10293 (N_10293,N_7887,N_8699);
nand U10294 (N_10294,N_7834,N_7588);
or U10295 (N_10295,N_8062,N_7840);
and U10296 (N_10296,N_8483,N_8119);
and U10297 (N_10297,N_8661,N_8886);
and U10298 (N_10298,N_8903,N_8384);
or U10299 (N_10299,N_7908,N_7839);
or U10300 (N_10300,N_8952,N_8537);
nor U10301 (N_10301,N_7672,N_7713);
nand U10302 (N_10302,N_7521,N_8687);
nor U10303 (N_10303,N_8792,N_7877);
nor U10304 (N_10304,N_7587,N_7571);
or U10305 (N_10305,N_8157,N_7819);
nand U10306 (N_10306,N_8944,N_7898);
nand U10307 (N_10307,N_8773,N_8556);
and U10308 (N_10308,N_7879,N_8589);
nor U10309 (N_10309,N_8221,N_8101);
nor U10310 (N_10310,N_8422,N_8436);
and U10311 (N_10311,N_8728,N_8168);
nand U10312 (N_10312,N_8858,N_7812);
and U10313 (N_10313,N_7502,N_7725);
and U10314 (N_10314,N_8421,N_8929);
and U10315 (N_10315,N_7883,N_8187);
or U10316 (N_10316,N_8000,N_8385);
and U10317 (N_10317,N_7714,N_8380);
and U10318 (N_10318,N_7978,N_7757);
nand U10319 (N_10319,N_7885,N_8616);
nor U10320 (N_10320,N_8557,N_8829);
or U10321 (N_10321,N_8653,N_8616);
or U10322 (N_10322,N_7855,N_8507);
and U10323 (N_10323,N_8326,N_8077);
and U10324 (N_10324,N_8013,N_8255);
nor U10325 (N_10325,N_8418,N_8401);
and U10326 (N_10326,N_7721,N_8935);
nand U10327 (N_10327,N_8315,N_7799);
nand U10328 (N_10328,N_8468,N_8819);
nand U10329 (N_10329,N_7734,N_8712);
or U10330 (N_10330,N_8006,N_8024);
nor U10331 (N_10331,N_7508,N_8985);
nand U10332 (N_10332,N_8100,N_8220);
or U10333 (N_10333,N_7854,N_8450);
or U10334 (N_10334,N_7869,N_7949);
and U10335 (N_10335,N_8098,N_8971);
nor U10336 (N_10336,N_7951,N_8278);
and U10337 (N_10337,N_8250,N_7541);
nor U10338 (N_10338,N_7833,N_7754);
nand U10339 (N_10339,N_8166,N_8989);
nor U10340 (N_10340,N_8222,N_8584);
nand U10341 (N_10341,N_7555,N_7532);
nand U10342 (N_10342,N_7801,N_8778);
nand U10343 (N_10343,N_7571,N_8935);
nor U10344 (N_10344,N_8549,N_8135);
nor U10345 (N_10345,N_7792,N_7737);
or U10346 (N_10346,N_7730,N_8896);
nor U10347 (N_10347,N_7868,N_8944);
or U10348 (N_10348,N_8046,N_7595);
or U10349 (N_10349,N_8010,N_8715);
and U10350 (N_10350,N_8871,N_7841);
or U10351 (N_10351,N_7779,N_8197);
and U10352 (N_10352,N_7848,N_7546);
nand U10353 (N_10353,N_8041,N_8859);
nand U10354 (N_10354,N_7625,N_7589);
nand U10355 (N_10355,N_8098,N_7621);
nand U10356 (N_10356,N_8310,N_8126);
nor U10357 (N_10357,N_8419,N_7834);
and U10358 (N_10358,N_8883,N_7584);
nor U10359 (N_10359,N_8574,N_8094);
nand U10360 (N_10360,N_8731,N_8575);
nor U10361 (N_10361,N_8502,N_7616);
or U10362 (N_10362,N_8421,N_8619);
nor U10363 (N_10363,N_8083,N_8049);
or U10364 (N_10364,N_7932,N_8334);
nand U10365 (N_10365,N_8890,N_7526);
and U10366 (N_10366,N_8860,N_7945);
and U10367 (N_10367,N_7502,N_8486);
or U10368 (N_10368,N_8923,N_8874);
and U10369 (N_10369,N_8836,N_8815);
and U10370 (N_10370,N_7992,N_8929);
or U10371 (N_10371,N_7853,N_8546);
or U10372 (N_10372,N_8051,N_8770);
nand U10373 (N_10373,N_8504,N_8507);
nand U10374 (N_10374,N_7604,N_8436);
nor U10375 (N_10375,N_7933,N_7545);
nand U10376 (N_10376,N_8603,N_8251);
nand U10377 (N_10377,N_8770,N_7554);
or U10378 (N_10378,N_8191,N_7936);
nor U10379 (N_10379,N_8257,N_7901);
nand U10380 (N_10380,N_7598,N_8981);
nor U10381 (N_10381,N_8980,N_8977);
and U10382 (N_10382,N_7520,N_8376);
nand U10383 (N_10383,N_8346,N_8602);
nand U10384 (N_10384,N_8680,N_7802);
nand U10385 (N_10385,N_7917,N_8146);
and U10386 (N_10386,N_7609,N_7817);
and U10387 (N_10387,N_8328,N_8250);
nor U10388 (N_10388,N_8142,N_8120);
and U10389 (N_10389,N_8758,N_7867);
nor U10390 (N_10390,N_8154,N_7812);
nand U10391 (N_10391,N_8160,N_7925);
nor U10392 (N_10392,N_8762,N_8371);
nand U10393 (N_10393,N_7548,N_8775);
or U10394 (N_10394,N_8832,N_7888);
and U10395 (N_10395,N_7855,N_8384);
and U10396 (N_10396,N_7769,N_7895);
and U10397 (N_10397,N_8073,N_7954);
nor U10398 (N_10398,N_8661,N_8046);
nor U10399 (N_10399,N_8105,N_7631);
nor U10400 (N_10400,N_8065,N_7720);
or U10401 (N_10401,N_7870,N_7585);
nor U10402 (N_10402,N_8847,N_7802);
or U10403 (N_10403,N_7609,N_8302);
or U10404 (N_10404,N_7647,N_7779);
nand U10405 (N_10405,N_7608,N_8037);
nand U10406 (N_10406,N_8132,N_8890);
nand U10407 (N_10407,N_7964,N_8820);
and U10408 (N_10408,N_8127,N_7674);
and U10409 (N_10409,N_8405,N_7943);
or U10410 (N_10410,N_8317,N_8907);
and U10411 (N_10411,N_7886,N_8570);
or U10412 (N_10412,N_8448,N_8113);
and U10413 (N_10413,N_8732,N_8167);
and U10414 (N_10414,N_7564,N_8332);
or U10415 (N_10415,N_8682,N_8852);
and U10416 (N_10416,N_8178,N_7835);
and U10417 (N_10417,N_7513,N_7777);
nand U10418 (N_10418,N_8955,N_8543);
or U10419 (N_10419,N_7983,N_8110);
nor U10420 (N_10420,N_8447,N_8388);
and U10421 (N_10421,N_8126,N_7782);
nor U10422 (N_10422,N_8291,N_8231);
and U10423 (N_10423,N_8513,N_8131);
and U10424 (N_10424,N_8215,N_8015);
or U10425 (N_10425,N_7972,N_8100);
xnor U10426 (N_10426,N_8602,N_7793);
and U10427 (N_10427,N_8773,N_8034);
and U10428 (N_10428,N_8845,N_7707);
nor U10429 (N_10429,N_7735,N_7639);
nor U10430 (N_10430,N_8120,N_8084);
or U10431 (N_10431,N_8758,N_8027);
nor U10432 (N_10432,N_8748,N_8845);
nand U10433 (N_10433,N_7619,N_7503);
or U10434 (N_10434,N_8928,N_8455);
nand U10435 (N_10435,N_8735,N_8725);
nor U10436 (N_10436,N_7530,N_8537);
or U10437 (N_10437,N_8716,N_8622);
or U10438 (N_10438,N_7965,N_7505);
nand U10439 (N_10439,N_8225,N_7691);
or U10440 (N_10440,N_8207,N_8728);
and U10441 (N_10441,N_7810,N_8743);
and U10442 (N_10442,N_8751,N_7892);
and U10443 (N_10443,N_7909,N_7666);
or U10444 (N_10444,N_8163,N_7629);
and U10445 (N_10445,N_8413,N_8498);
nand U10446 (N_10446,N_8668,N_7543);
nor U10447 (N_10447,N_7750,N_8343);
xnor U10448 (N_10448,N_8768,N_8405);
and U10449 (N_10449,N_7728,N_8445);
and U10450 (N_10450,N_8061,N_8513);
nor U10451 (N_10451,N_8176,N_8001);
nand U10452 (N_10452,N_8648,N_7623);
or U10453 (N_10453,N_8787,N_7767);
nand U10454 (N_10454,N_8420,N_8958);
and U10455 (N_10455,N_8335,N_7590);
nor U10456 (N_10456,N_7503,N_8621);
nand U10457 (N_10457,N_8398,N_7601);
nor U10458 (N_10458,N_7555,N_7672);
or U10459 (N_10459,N_7548,N_7745);
nand U10460 (N_10460,N_8259,N_7835);
or U10461 (N_10461,N_8898,N_8847);
nor U10462 (N_10462,N_7661,N_8794);
and U10463 (N_10463,N_8378,N_7646);
or U10464 (N_10464,N_8766,N_8117);
and U10465 (N_10465,N_8973,N_7605);
or U10466 (N_10466,N_8863,N_8498);
and U10467 (N_10467,N_8509,N_7747);
nor U10468 (N_10468,N_8684,N_8868);
or U10469 (N_10469,N_8419,N_7804);
and U10470 (N_10470,N_7679,N_7923);
nand U10471 (N_10471,N_8121,N_7671);
and U10472 (N_10472,N_8465,N_7980);
and U10473 (N_10473,N_7875,N_8444);
or U10474 (N_10474,N_7863,N_7864);
nand U10475 (N_10475,N_7785,N_8531);
or U10476 (N_10476,N_8740,N_8508);
and U10477 (N_10477,N_8235,N_8197);
nand U10478 (N_10478,N_8168,N_7878);
nand U10479 (N_10479,N_8357,N_8299);
nor U10480 (N_10480,N_7893,N_8678);
or U10481 (N_10481,N_8997,N_8714);
or U10482 (N_10482,N_8731,N_8141);
and U10483 (N_10483,N_7640,N_8807);
nand U10484 (N_10484,N_7566,N_7520);
or U10485 (N_10485,N_8741,N_8134);
and U10486 (N_10486,N_8446,N_8406);
or U10487 (N_10487,N_8900,N_8650);
nor U10488 (N_10488,N_8032,N_8505);
and U10489 (N_10489,N_7957,N_8481);
or U10490 (N_10490,N_7614,N_7655);
nand U10491 (N_10491,N_8857,N_8815);
nand U10492 (N_10492,N_8074,N_8716);
and U10493 (N_10493,N_7524,N_8039);
or U10494 (N_10494,N_8086,N_8253);
nor U10495 (N_10495,N_8623,N_8219);
and U10496 (N_10496,N_7937,N_8210);
nor U10497 (N_10497,N_8405,N_8715);
nor U10498 (N_10498,N_7762,N_8894);
nand U10499 (N_10499,N_8137,N_8038);
nor U10500 (N_10500,N_10197,N_9739);
nand U10501 (N_10501,N_9844,N_9288);
nand U10502 (N_10502,N_9995,N_9886);
nor U10503 (N_10503,N_9525,N_9847);
nand U10504 (N_10504,N_9348,N_9273);
nor U10505 (N_10505,N_10133,N_10092);
nor U10506 (N_10506,N_9204,N_10240);
nor U10507 (N_10507,N_10216,N_9323);
or U10508 (N_10508,N_9430,N_10081);
and U10509 (N_10509,N_10299,N_9583);
and U10510 (N_10510,N_9282,N_10336);
nand U10511 (N_10511,N_10297,N_10064);
and U10512 (N_10512,N_9118,N_10466);
and U10513 (N_10513,N_10010,N_10429);
nand U10514 (N_10514,N_10249,N_9837);
and U10515 (N_10515,N_9668,N_9636);
and U10516 (N_10516,N_10091,N_9817);
and U10517 (N_10517,N_10014,N_9326);
nand U10518 (N_10518,N_10199,N_10219);
nor U10519 (N_10519,N_9381,N_10002);
or U10520 (N_10520,N_10251,N_9445);
nor U10521 (N_10521,N_9045,N_10395);
or U10522 (N_10522,N_9728,N_9604);
nor U10523 (N_10523,N_9364,N_9090);
or U10524 (N_10524,N_10163,N_9352);
nand U10525 (N_10525,N_10190,N_9310);
nor U10526 (N_10526,N_9664,N_10481);
and U10527 (N_10527,N_10356,N_9005);
nand U10528 (N_10528,N_9626,N_10454);
nor U10529 (N_10529,N_10017,N_10156);
or U10530 (N_10530,N_10161,N_9457);
and U10531 (N_10531,N_10252,N_9599);
or U10532 (N_10532,N_9635,N_9785);
nand U10533 (N_10533,N_9486,N_10460);
nand U10534 (N_10534,N_9201,N_9949);
nor U10535 (N_10535,N_9932,N_9126);
nand U10536 (N_10536,N_9577,N_9796);
and U10537 (N_10537,N_9605,N_9451);
nand U10538 (N_10538,N_10257,N_9329);
nand U10539 (N_10539,N_10269,N_9734);
nor U10540 (N_10540,N_9829,N_9539);
nand U10541 (N_10541,N_10462,N_9174);
or U10542 (N_10542,N_10048,N_10205);
or U10543 (N_10543,N_9614,N_10228);
and U10544 (N_10544,N_10185,N_9939);
or U10545 (N_10545,N_9193,N_10420);
nor U10546 (N_10546,N_10265,N_10130);
or U10547 (N_10547,N_10174,N_9906);
nand U10548 (N_10548,N_9633,N_9562);
and U10549 (N_10549,N_9259,N_9362);
nand U10550 (N_10550,N_10142,N_9954);
xnor U10551 (N_10551,N_10270,N_10381);
nand U10552 (N_10552,N_10346,N_9615);
nand U10553 (N_10553,N_9570,N_9320);
nor U10554 (N_10554,N_9440,N_9957);
or U10555 (N_10555,N_10065,N_9152);
or U10556 (N_10556,N_9600,N_9754);
or U10557 (N_10557,N_9942,N_10282);
nand U10558 (N_10558,N_10062,N_10117);
and U10559 (N_10559,N_9142,N_9770);
nor U10560 (N_10560,N_9564,N_9137);
nor U10561 (N_10561,N_10098,N_9285);
and U10562 (N_10562,N_10424,N_10242);
nand U10563 (N_10563,N_9062,N_9280);
or U10564 (N_10564,N_9850,N_10331);
nand U10565 (N_10565,N_10340,N_9104);
and U10566 (N_10566,N_9656,N_9861);
and U10567 (N_10567,N_10215,N_10207);
nand U10568 (N_10568,N_9233,N_9033);
or U10569 (N_10569,N_10070,N_10468);
nor U10570 (N_10570,N_9298,N_10001);
nand U10571 (N_10571,N_9928,N_9719);
nor U10572 (N_10572,N_9946,N_10068);
and U10573 (N_10573,N_9907,N_9257);
or U10574 (N_10574,N_10223,N_9023);
or U10575 (N_10575,N_9867,N_9370);
nor U10576 (N_10576,N_9998,N_10123);
and U10577 (N_10577,N_9400,N_9549);
or U10578 (N_10578,N_9331,N_10260);
nor U10579 (N_10579,N_9220,N_9253);
nand U10580 (N_10580,N_10353,N_9077);
or U10581 (N_10581,N_9456,N_10406);
or U10582 (N_10582,N_9027,N_9689);
and U10583 (N_10583,N_9517,N_9043);
and U10584 (N_10584,N_9736,N_10097);
nor U10585 (N_10585,N_9640,N_9088);
nor U10586 (N_10586,N_9411,N_10300);
or U10587 (N_10587,N_9303,N_9497);
nand U10588 (N_10588,N_9685,N_10321);
nand U10589 (N_10589,N_10060,N_10140);
nor U10590 (N_10590,N_9908,N_10035);
nand U10591 (N_10591,N_10482,N_9985);
nand U10592 (N_10592,N_10128,N_10271);
nor U10593 (N_10593,N_10499,N_10108);
nand U10594 (N_10594,N_9710,N_9649);
nor U10595 (N_10595,N_9302,N_9530);
nand U10596 (N_10596,N_10218,N_9569);
nor U10597 (N_10597,N_10054,N_10415);
xnor U10598 (N_10598,N_9912,N_10279);
nor U10599 (N_10599,N_10289,N_9556);
and U10600 (N_10600,N_9172,N_9572);
nor U10601 (N_10601,N_9346,N_9264);
nor U10602 (N_10602,N_9116,N_9763);
nor U10603 (N_10603,N_9226,N_9522);
or U10604 (N_10604,N_10389,N_9543);
nor U10605 (N_10605,N_9811,N_10203);
nand U10606 (N_10606,N_9859,N_10339);
nand U10607 (N_10607,N_9744,N_9474);
and U10608 (N_10608,N_9792,N_10397);
or U10609 (N_10609,N_10447,N_10405);
nor U10610 (N_10610,N_9654,N_10029);
and U10611 (N_10611,N_9720,N_9631);
nor U10612 (N_10612,N_9214,N_9444);
and U10613 (N_10613,N_9742,N_10224);
or U10614 (N_10614,N_9422,N_9794);
nand U10615 (N_10615,N_9831,N_9977);
nand U10616 (N_10616,N_9363,N_10487);
nand U10617 (N_10617,N_10044,N_10398);
or U10618 (N_10618,N_9112,N_10493);
and U10619 (N_10619,N_9666,N_9997);
nor U10620 (N_10620,N_9435,N_9820);
nand U10621 (N_10621,N_9805,N_9904);
nand U10622 (N_10622,N_10354,N_10359);
and U10623 (N_10623,N_9948,N_10072);
or U10624 (N_10624,N_9771,N_10438);
nand U10625 (N_10625,N_10226,N_9925);
or U10626 (N_10626,N_9495,N_9874);
or U10627 (N_10627,N_10086,N_9822);
and U10628 (N_10628,N_10032,N_9501);
nor U10629 (N_10629,N_9095,N_10426);
nor U10630 (N_10630,N_9171,N_9246);
or U10631 (N_10631,N_10194,N_9415);
nor U10632 (N_10632,N_9568,N_10109);
nand U10633 (N_10633,N_9718,N_10452);
and U10634 (N_10634,N_10372,N_9038);
nor U10635 (N_10635,N_9416,N_10248);
nand U10636 (N_10636,N_10285,N_9813);
nand U10637 (N_10637,N_9341,N_9084);
or U10638 (N_10638,N_9863,N_9202);
and U10639 (N_10639,N_9970,N_10115);
nand U10640 (N_10640,N_10030,N_9947);
nor U10641 (N_10641,N_9487,N_10166);
nand U10642 (N_10642,N_9842,N_9756);
nor U10643 (N_10643,N_10083,N_10134);
and U10644 (N_10644,N_9231,N_9165);
nor U10645 (N_10645,N_10446,N_9513);
nor U10646 (N_10646,N_9296,N_10085);
nor U10647 (N_10647,N_9943,N_9625);
nor U10648 (N_10648,N_9458,N_10192);
nand U10649 (N_10649,N_10434,N_9268);
and U10650 (N_10650,N_9052,N_9012);
nand U10651 (N_10651,N_9559,N_9723);
or U10652 (N_10652,N_9067,N_9824);
and U10653 (N_10653,N_9671,N_10052);
or U10654 (N_10654,N_10178,N_9592);
or U10655 (N_10655,N_9597,N_10168);
or U10656 (N_10656,N_9237,N_9176);
or U10657 (N_10657,N_9294,N_10102);
nand U10658 (N_10658,N_10319,N_10419);
and U10659 (N_10659,N_10293,N_9937);
or U10660 (N_10660,N_9894,N_9630);
and U10661 (N_10661,N_9755,N_9029);
nand U10662 (N_10662,N_10079,N_10058);
nor U10663 (N_10663,N_9629,N_10479);
or U10664 (N_10664,N_9546,N_10416);
nand U10665 (N_10665,N_9853,N_9648);
nand U10666 (N_10666,N_10306,N_9120);
nand U10667 (N_10667,N_9490,N_9524);
nand U10668 (N_10668,N_10088,N_9211);
and U10669 (N_10669,N_9743,N_10361);
and U10670 (N_10670,N_10041,N_9421);
and U10671 (N_10671,N_10276,N_9827);
or U10672 (N_10672,N_9160,N_10394);
nor U10673 (N_10673,N_10028,N_9013);
nand U10674 (N_10674,N_10009,N_9965);
nor U10675 (N_10675,N_9892,N_9958);
nor U10676 (N_10676,N_9727,N_10188);
nor U10677 (N_10677,N_10322,N_9836);
or U10678 (N_10678,N_9810,N_9747);
nor U10679 (N_10679,N_10124,N_9207);
and U10680 (N_10680,N_9395,N_9070);
nor U10681 (N_10681,N_9278,N_9425);
or U10682 (N_10682,N_9047,N_9167);
nor U10683 (N_10683,N_9040,N_10314);
nand U10684 (N_10684,N_9493,N_9980);
and U10685 (N_10685,N_9984,N_10440);
xnor U10686 (N_10686,N_10329,N_9235);
and U10687 (N_10687,N_9146,N_10266);
nand U10688 (N_10688,N_9638,N_10409);
or U10689 (N_10689,N_9586,N_10318);
nand U10690 (N_10690,N_9818,N_9927);
and U10691 (N_10691,N_9574,N_10316);
nand U10692 (N_10692,N_10323,N_9001);
or U10693 (N_10693,N_9950,N_9641);
and U10694 (N_10694,N_9851,N_10018);
or U10695 (N_10695,N_9065,N_9439);
nand U10696 (N_10696,N_9905,N_9979);
or U10697 (N_10697,N_9145,N_9482);
or U10698 (N_10698,N_9313,N_10061);
or U10699 (N_10699,N_9159,N_10090);
nor U10700 (N_10700,N_9433,N_9494);
nand U10701 (N_10701,N_10268,N_9807);
nand U10702 (N_10702,N_10013,N_9598);
xor U10703 (N_10703,N_9974,N_9035);
and U10704 (N_10704,N_9772,N_9918);
and U10705 (N_10705,N_9377,N_10475);
nor U10706 (N_10706,N_9042,N_9491);
nand U10707 (N_10707,N_9702,N_9308);
or U10708 (N_10708,N_9085,N_9617);
nand U10709 (N_10709,N_9469,N_10315);
and U10710 (N_10710,N_10000,N_9355);
nand U10711 (N_10711,N_9558,N_10187);
and U10712 (N_10712,N_9579,N_9188);
or U10713 (N_10713,N_10392,N_10101);
nor U10714 (N_10714,N_10368,N_9437);
nor U10715 (N_10715,N_10349,N_10444);
nand U10716 (N_10716,N_9519,N_10333);
and U10717 (N_10717,N_9930,N_9109);
nor U10718 (N_10718,N_9748,N_9639);
or U10719 (N_10719,N_10459,N_9752);
nor U10720 (N_10720,N_9209,N_10135);
and U10721 (N_10721,N_9356,N_10179);
nand U10722 (N_10722,N_10427,N_9384);
nand U10723 (N_10723,N_9389,N_10150);
or U10724 (N_10724,N_9473,N_10127);
and U10725 (N_10725,N_9299,N_9647);
nor U10726 (N_10726,N_9520,N_9976);
and U10727 (N_10727,N_9170,N_10141);
and U10728 (N_10728,N_10267,N_10023);
nor U10729 (N_10729,N_10171,N_9114);
or U10730 (N_10730,N_9774,N_10131);
or U10731 (N_10731,N_10334,N_9156);
or U10732 (N_10732,N_9858,N_9607);
and U10733 (N_10733,N_9373,N_9982);
nor U10734 (N_10734,N_9420,N_9452);
and U10735 (N_10735,N_10256,N_10042);
or U10736 (N_10736,N_9499,N_9397);
or U10737 (N_10737,N_10132,N_10272);
and U10738 (N_10738,N_10206,N_9642);
or U10739 (N_10739,N_10378,N_9484);
and U10740 (N_10740,N_9483,N_9011);
nand U10741 (N_10741,N_9022,N_9870);
and U10742 (N_10742,N_9127,N_10495);
nand U10743 (N_10743,N_9398,N_10414);
nand U10744 (N_10744,N_10437,N_9407);
or U10745 (N_10745,N_10089,N_10432);
and U10746 (N_10746,N_9210,N_9178);
nor U10747 (N_10747,N_9149,N_9677);
or U10748 (N_10748,N_9344,N_9821);
and U10749 (N_10749,N_9215,N_10004);
nor U10750 (N_10750,N_9884,N_9441);
nand U10751 (N_10751,N_9401,N_9595);
or U10752 (N_10752,N_9737,N_9131);
nand U10753 (N_10753,N_9554,N_9512);
nand U10754 (N_10754,N_10037,N_9103);
and U10755 (N_10755,N_10073,N_9369);
and U10756 (N_10756,N_9304,N_10019);
or U10757 (N_10757,N_9080,N_9276);
or U10758 (N_10758,N_10464,N_10183);
and U10759 (N_10759,N_9895,N_10213);
or U10760 (N_10760,N_9923,N_10374);
nor U10761 (N_10761,N_9387,N_10158);
nor U10762 (N_10762,N_9448,N_9250);
nand U10763 (N_10763,N_9661,N_9391);
nor U10764 (N_10764,N_9372,N_9694);
nand U10765 (N_10765,N_10049,N_10116);
or U10766 (N_10766,N_10488,N_9882);
nand U10767 (N_10767,N_10317,N_9988);
nor U10768 (N_10768,N_9267,N_10347);
nor U10769 (N_10769,N_10380,N_9291);
and U10770 (N_10770,N_9509,N_9550);
nand U10771 (N_10771,N_9478,N_10386);
nor U10772 (N_10772,N_9347,N_9069);
nand U10773 (N_10773,N_9975,N_9361);
nand U10774 (N_10774,N_10253,N_9972);
nand U10775 (N_10775,N_9318,N_10175);
or U10776 (N_10776,N_9196,N_10153);
nor U10777 (N_10777,N_9696,N_9026);
nor U10778 (N_10778,N_10084,N_10275);
or U10779 (N_10779,N_10087,N_9812);
and U10780 (N_10780,N_9699,N_9585);
nand U10781 (N_10781,N_9540,N_9472);
and U10782 (N_10782,N_9964,N_10144);
nor U10783 (N_10783,N_10177,N_9060);
nor U10784 (N_10784,N_10208,N_9968);
or U10785 (N_10785,N_10401,N_9242);
nor U10786 (N_10786,N_10477,N_10055);
nor U10787 (N_10787,N_9132,N_10232);
nand U10788 (N_10788,N_10463,N_9135);
and U10789 (N_10789,N_10107,N_10182);
nor U10790 (N_10790,N_9724,N_9826);
and U10791 (N_10791,N_10362,N_9480);
and U10792 (N_10792,N_9404,N_9833);
nand U10793 (N_10793,N_10180,N_9388);
nor U10794 (N_10794,N_9751,N_9460);
or U10795 (N_10795,N_9097,N_9999);
or U10796 (N_10796,N_10121,N_9672);
nor U10797 (N_10797,N_10484,N_9703);
and U10798 (N_10798,N_9529,N_9295);
or U10799 (N_10799,N_9305,N_9393);
and U10800 (N_10800,N_9681,N_9766);
and U10801 (N_10801,N_9613,N_10118);
nand U10802 (N_10802,N_9555,N_9228);
nand U10803 (N_10803,N_9248,N_10006);
or U10804 (N_10804,N_10114,N_9891);
nor U10805 (N_10805,N_9275,N_9862);
nand U10806 (N_10806,N_10411,N_10413);
and U10807 (N_10807,N_9101,N_9477);
and U10808 (N_10808,N_10129,N_10231);
nor U10809 (N_10809,N_9868,N_9732);
nand U10810 (N_10810,N_9423,N_10137);
or U10811 (N_10811,N_9717,N_9147);
or U10812 (N_10812,N_10154,N_10443);
and U10813 (N_10813,N_9809,N_9213);
nand U10814 (N_10814,N_10393,N_9914);
nor U10815 (N_10815,N_9306,N_9096);
nand U10816 (N_10816,N_10008,N_10012);
and U10817 (N_10817,N_9762,N_10011);
nor U10818 (N_10818,N_10288,N_10383);
nor U10819 (N_10819,N_10407,N_9986);
or U10820 (N_10820,N_9992,N_9663);
or U10821 (N_10821,N_9079,N_9406);
nand U10822 (N_10822,N_9889,N_9399);
nor U10823 (N_10823,N_9117,N_9136);
nor U10824 (N_10824,N_9144,N_9777);
nor U10825 (N_10825,N_9197,N_9655);
or U10826 (N_10826,N_9931,N_9050);
nor U10827 (N_10827,N_9578,N_9704);
or U10828 (N_10828,N_9073,N_9236);
or U10829 (N_10829,N_9686,N_10038);
and U10830 (N_10830,N_9588,N_9297);
or U10831 (N_10831,N_10186,N_10326);
nor U10832 (N_10832,N_10096,N_10422);
nor U10833 (N_10833,N_9910,N_9878);
nand U10834 (N_10834,N_10465,N_9669);
nand U10835 (N_10835,N_9279,N_9338);
and U10836 (N_10836,N_9838,N_9773);
or U10837 (N_10837,N_9087,N_9611);
or U10838 (N_10838,N_9716,N_9092);
nor U10839 (N_10839,N_10243,N_9767);
nor U10840 (N_10840,N_9667,N_10230);
nand U10841 (N_10841,N_9270,N_9322);
xnor U10842 (N_10842,N_9860,N_9746);
nor U10843 (N_10843,N_9072,N_9620);
nor U10844 (N_10844,N_9919,N_9383);
nor U10845 (N_10845,N_10149,N_9856);
nand U10846 (N_10846,N_9317,N_9098);
and U10847 (N_10847,N_10382,N_10496);
or U10848 (N_10848,N_9637,N_9485);
xnor U10849 (N_10849,N_10435,N_9100);
and U10850 (N_10850,N_9428,N_9498);
nand U10851 (N_10851,N_9223,N_10139);
or U10852 (N_10852,N_9075,N_9106);
or U10853 (N_10853,N_10364,N_9557);
or U10854 (N_10854,N_9769,N_9885);
or U10855 (N_10855,N_9573,N_9177);
nand U10856 (N_10856,N_9234,N_9518);
or U10857 (N_10857,N_9189,N_9725);
or U10858 (N_10858,N_9057,N_10273);
nand U10859 (N_10859,N_9453,N_9528);
nand U10860 (N_10860,N_9500,N_10335);
nand U10861 (N_10861,N_9349,N_10157);
and U10862 (N_10862,N_9224,N_9429);
or U10863 (N_10863,N_9778,N_9527);
nand U10864 (N_10864,N_9107,N_10441);
xor U10865 (N_10865,N_9018,N_9151);
nor U10866 (N_10866,N_10067,N_9263);
nor U10867 (N_10867,N_9459,N_9108);
nor U10868 (N_10868,N_10222,N_9463);
nand U10869 (N_10869,N_10418,N_10050);
nor U10870 (N_10870,N_10365,N_9646);
nor U10871 (N_10871,N_9194,N_9333);
nand U10872 (N_10872,N_9883,N_10369);
and U10873 (N_10873,N_9799,N_10312);
or U10874 (N_10874,N_9665,N_10066);
and U10875 (N_10875,N_10296,N_9800);
or U10876 (N_10876,N_10220,N_10113);
nor U10877 (N_10877,N_9261,N_9502);
nand U10878 (N_10878,N_9709,N_9786);
nor U10879 (N_10879,N_9738,N_10033);
nand U10880 (N_10880,N_9571,N_9157);
nand U10881 (N_10881,N_9768,N_10280);
or U10882 (N_10882,N_9798,N_10425);
or U10883 (N_10883,N_9782,N_10093);
xnor U10884 (N_10884,N_9247,N_9366);
or U10885 (N_10885,N_10304,N_10221);
nand U10886 (N_10886,N_9651,N_9921);
or U10887 (N_10887,N_10286,N_9195);
or U10888 (N_10888,N_10100,N_9314);
nand U10889 (N_10889,N_9410,N_9535);
or U10890 (N_10890,N_9621,N_10167);
or U10891 (N_10891,N_10120,N_9922);
or U10892 (N_10892,N_9541,N_10490);
and U10893 (N_10893,N_9424,N_9697);
and U10894 (N_10894,N_9447,N_10210);
or U10895 (N_10895,N_10095,N_9099);
nand U10896 (N_10896,N_9749,N_9783);
or U10897 (N_10897,N_9693,N_9081);
and U10898 (N_10898,N_10445,N_9877);
xor U10899 (N_10899,N_9622,N_9956);
and U10900 (N_10900,N_9712,N_10053);
nand U10901 (N_10901,N_9835,N_9565);
nor U10902 (N_10902,N_10217,N_9653);
and U10903 (N_10903,N_9113,N_9074);
or U10904 (N_10904,N_9125,N_9028);
or U10905 (N_10905,N_9606,N_9841);
or U10906 (N_10906,N_9688,N_10498);
and U10907 (N_10907,N_9828,N_9037);
and U10908 (N_10908,N_9283,N_9514);
or U10909 (N_10909,N_10046,N_9616);
and U10910 (N_10910,N_9492,N_10305);
nor U10911 (N_10911,N_9489,N_9274);
nor U10912 (N_10912,N_9680,N_9593);
or U10913 (N_10913,N_10237,N_10325);
nand U10914 (N_10914,N_9053,N_9007);
nand U10915 (N_10915,N_9203,N_10483);
nand U10916 (N_10916,N_9337,N_9627);
nand U10917 (N_10917,N_9030,N_9155);
or U10918 (N_10918,N_10417,N_9232);
nor U10919 (N_10919,N_9969,N_9186);
nand U10920 (N_10920,N_10351,N_10172);
nor U10921 (N_10921,N_9678,N_9690);
and U10922 (N_10922,N_10338,N_10025);
nand U10923 (N_10923,N_9902,N_10471);
nand U10924 (N_10924,N_9547,N_9086);
or U10925 (N_10925,N_10045,N_9544);
or U10926 (N_10926,N_9417,N_9580);
or U10927 (N_10927,N_10355,N_9219);
and U10928 (N_10928,N_9345,N_9687);
and U10929 (N_10929,N_9260,N_10181);
nor U10930 (N_10930,N_9707,N_9582);
nand U10931 (N_10931,N_9272,N_9059);
and U10932 (N_10932,N_9335,N_10262);
or U10933 (N_10933,N_9455,N_9192);
nor U10934 (N_10934,N_10377,N_9515);
nand U10935 (N_10935,N_10489,N_10330);
nor U10936 (N_10936,N_9183,N_9900);
and U10937 (N_10937,N_9983,N_9632);
nand U10938 (N_10938,N_9576,N_9368);
and U10939 (N_10939,N_10457,N_9840);
and U10940 (N_10940,N_9412,N_10461);
and U10941 (N_10941,N_9408,N_10152);
nand U10942 (N_10942,N_9789,N_9581);
nor U10943 (N_10943,N_9801,N_9190);
nor U10944 (N_10944,N_9516,N_9000);
nand U10945 (N_10945,N_10176,N_9990);
nor U10946 (N_10946,N_10027,N_9360);
or U10947 (N_10947,N_9596,N_10458);
nand U10948 (N_10948,N_9325,N_9924);
or U10949 (N_10949,N_9802,N_9164);
nor U10950 (N_10950,N_9873,N_9340);
nand U10951 (N_10951,N_9021,N_9134);
or U10952 (N_10952,N_9169,N_10403);
nand U10953 (N_10953,N_10442,N_9761);
nand U10954 (N_10954,N_9695,N_9915);
and U10955 (N_10955,N_9701,N_9130);
and U10956 (N_10956,N_10345,N_9692);
and U10957 (N_10957,N_9449,N_9803);
nand U10958 (N_10958,N_10358,N_10026);
or U10959 (N_10959,N_9143,N_9198);
nand U10960 (N_10960,N_9993,N_9832);
nand U10961 (N_10961,N_9312,N_9775);
and U10962 (N_10962,N_9048,N_9951);
and U10963 (N_10963,N_10404,N_9071);
and U10964 (N_10964,N_9934,N_9713);
and U10965 (N_10965,N_10069,N_9123);
and U10966 (N_10966,N_10020,N_10308);
nor U10967 (N_10967,N_9255,N_9779);
and U10968 (N_10968,N_9468,N_9508);
or U10969 (N_10969,N_9293,N_9307);
and U10970 (N_10970,N_10313,N_10193);
or U10971 (N_10971,N_9350,N_9465);
or U10972 (N_10972,N_10337,N_10467);
nand U10973 (N_10973,N_10080,N_9032);
nand U10974 (N_10974,N_10076,N_9705);
or U10975 (N_10975,N_9020,N_9036);
nand U10976 (N_10976,N_9505,N_9561);
or U10977 (N_10977,N_10448,N_10202);
nor U10978 (N_10978,N_9227,N_9454);
and U10979 (N_10979,N_9676,N_9175);
and U10980 (N_10980,N_9981,N_10453);
nand U10981 (N_10981,N_9590,N_10122);
nand U10982 (N_10982,N_9652,N_9823);
and U10983 (N_10983,N_9241,N_10332);
nor U10984 (N_10984,N_10348,N_9839);
and U10985 (N_10985,N_10151,N_10492);
nor U10986 (N_10986,N_10169,N_9650);
nand U10987 (N_10987,N_10341,N_10343);
nand U10988 (N_10988,N_9121,N_9367);
nand U10989 (N_10989,N_9898,N_9758);
nand U10990 (N_10990,N_9238,N_9531);
or U10991 (N_10991,N_9936,N_9920);
and U10992 (N_10992,N_10396,N_10494);
or U10993 (N_10993,N_9034,N_9140);
or U10994 (N_10994,N_10255,N_10162);
nand U10995 (N_10995,N_9618,N_10043);
or U10996 (N_10996,N_9358,N_10016);
and U10997 (N_10997,N_10039,N_10258);
nor U10998 (N_10998,N_9760,N_9684);
nor U10999 (N_10999,N_9991,N_10204);
nand U11000 (N_11000,N_9380,N_9797);
and U11001 (N_11001,N_10303,N_9733);
and U11002 (N_11002,N_9945,N_9154);
and U11003 (N_11003,N_9376,N_10384);
or U11004 (N_11004,N_9432,N_9218);
and U11005 (N_11005,N_10198,N_9199);
nor U11006 (N_11006,N_9251,N_9722);
and U11007 (N_11007,N_9128,N_9041);
and U11008 (N_11008,N_9619,N_9691);
and U11009 (N_11009,N_10366,N_10164);
and U11010 (N_11010,N_10034,N_9258);
nor U11011 (N_11011,N_9185,N_9708);
nand U11012 (N_11012,N_10473,N_9019);
nand U11013 (N_11013,N_10373,N_9216);
and U11014 (N_11014,N_9063,N_9466);
nand U11015 (N_11015,N_10147,N_9857);
nor U11016 (N_11016,N_9787,N_10244);
and U11017 (N_11017,N_9804,N_10450);
nand U11018 (N_11018,N_9419,N_9316);
and U11019 (N_11019,N_9962,N_9292);
nand U11020 (N_11020,N_9119,N_9624);
nand U11021 (N_11021,N_9311,N_10209);
nand U11022 (N_11022,N_9819,N_9010);
nor U11023 (N_11023,N_10212,N_9634);
or U11024 (N_11024,N_9963,N_10350);
or U11025 (N_11025,N_9507,N_9017);
or U11026 (N_11026,N_9846,N_10078);
nor U11027 (N_11027,N_9989,N_10485);
nand U11028 (N_11028,N_9481,N_10497);
and U11029 (N_11029,N_10105,N_9643);
nand U11030 (N_11030,N_10469,N_9301);
nor U11031 (N_11031,N_9953,N_9609);
nor U11032 (N_11032,N_10099,N_9068);
xor U11033 (N_11033,N_10376,N_9240);
and U11034 (N_11034,N_9321,N_9475);
nor U11035 (N_11035,N_9025,N_10201);
nor U11036 (N_11036,N_10196,N_9888);
and U11037 (N_11037,N_9996,N_9479);
nand U11038 (N_11038,N_9351,N_9729);
nor U11039 (N_11039,N_10233,N_9082);
nand U11040 (N_11040,N_10388,N_10238);
or U11041 (N_11041,N_9660,N_9536);
nand U11042 (N_11042,N_9269,N_9941);
and U11043 (N_11043,N_10015,N_10370);
nor U11044 (N_11044,N_10363,N_9971);
and U11045 (N_11045,N_10480,N_10412);
or U11046 (N_11046,N_9243,N_9700);
and U11047 (N_11047,N_9815,N_9414);
nand U11048 (N_11048,N_9488,N_10428);
or U11049 (N_11049,N_9212,N_9180);
or U11050 (N_11050,N_9105,N_9089);
and U11051 (N_11051,N_10352,N_9168);
nor U11052 (N_11052,N_9006,N_10094);
nand U11053 (N_11053,N_9141,N_10136);
nand U11054 (N_11054,N_10309,N_9431);
nor U11055 (N_11055,N_9327,N_9115);
nor U11056 (N_11056,N_10456,N_9324);
nor U11057 (N_11057,N_10005,N_9575);
and U11058 (N_11058,N_9139,N_10476);
and U11059 (N_11059,N_9750,N_10059);
nand U11060 (N_11060,N_10342,N_9816);
nand U11061 (N_11061,N_10486,N_9955);
nand U11062 (N_11062,N_9780,N_10189);
or U11063 (N_11063,N_9058,N_9793);
and U11064 (N_11064,N_10379,N_10307);
and U11065 (N_11065,N_10320,N_9277);
and U11066 (N_11066,N_10082,N_9864);
and U11067 (N_11067,N_10478,N_10165);
nand U11068 (N_11068,N_9467,N_9462);
nand U11069 (N_11069,N_10298,N_9008);
nand U11070 (N_11070,N_10143,N_9051);
nor U11071 (N_11071,N_9589,N_9674);
nor U11072 (N_11072,N_9003,N_10281);
nor U11073 (N_11073,N_10278,N_9731);
nand U11074 (N_11074,N_9890,N_9776);
nor U11075 (N_11075,N_9553,N_9933);
and U11076 (N_11076,N_9336,N_9426);
nand U11077 (N_11077,N_9266,N_9181);
or U11078 (N_11078,N_9434,N_9470);
or U11079 (N_11079,N_9623,N_9683);
nand U11080 (N_11080,N_10146,N_9332);
nand U11081 (N_11081,N_9790,N_10410);
or U11082 (N_11082,N_9161,N_10051);
nand U11083 (N_11083,N_9254,N_9402);
and U11084 (N_11084,N_9808,N_9994);
nor U11085 (N_11085,N_9865,N_9061);
and U11086 (N_11086,N_9715,N_9711);
nor U11087 (N_11087,N_9788,N_9608);
and U11088 (N_11088,N_9093,N_9158);
nor U11089 (N_11089,N_9952,N_10236);
nand U11090 (N_11090,N_9532,N_10110);
and U11091 (N_11091,N_9076,N_9973);
nand U11092 (N_11092,N_9806,N_10294);
and U11093 (N_11093,N_9730,N_9644);
or U11094 (N_11094,N_9959,N_10310);
or U11095 (N_11095,N_9405,N_9427);
or U11096 (N_11096,N_10491,N_9111);
nand U11097 (N_11097,N_9024,N_10170);
or U11098 (N_11098,N_9814,N_9173);
and U11099 (N_11099,N_9386,N_9319);
nor U11100 (N_11100,N_9413,N_10103);
and U11101 (N_11101,N_9365,N_10063);
nand U11102 (N_11102,N_9354,N_10470);
or U11103 (N_11103,N_9064,N_9265);
or U11104 (N_11104,N_9926,N_10261);
or U11105 (N_11105,N_9471,N_9901);
and U11106 (N_11106,N_9300,N_9866);
nand U11107 (N_11107,N_9548,N_9403);
nor U11108 (N_11108,N_9602,N_9339);
and U11109 (N_11109,N_9221,N_10071);
and U11110 (N_11110,N_10003,N_9852);
or U11111 (N_11111,N_9764,N_9418);
or U11112 (N_11112,N_9757,N_10451);
and U11113 (N_11113,N_9110,N_10375);
nand U11114 (N_11114,N_9869,N_9496);
or U11115 (N_11115,N_9503,N_9897);
and U11116 (N_11116,N_9133,N_10106);
nor U11117 (N_11117,N_9309,N_9014);
and U11118 (N_11118,N_10119,N_10385);
nand U11119 (N_11119,N_9256,N_9587);
or U11120 (N_11120,N_9357,N_10360);
and U11121 (N_11121,N_10250,N_9659);
nor U11122 (N_11122,N_9271,N_9745);
or U11123 (N_11123,N_9016,N_9443);
nand U11124 (N_11124,N_10367,N_10254);
or U11125 (N_11125,N_9166,N_9909);
nand U11126 (N_11126,N_9791,N_9978);
or U11127 (N_11127,N_9584,N_9610);
nor U11128 (N_11128,N_9382,N_9450);
and U11129 (N_11129,N_10173,N_9184);
and U11130 (N_11130,N_10234,N_9552);
or U11131 (N_11131,N_10274,N_10474);
nor U11132 (N_11132,N_9191,N_9940);
and U11133 (N_11133,N_9880,N_9881);
or U11134 (N_11134,N_9476,N_9179);
nor U11135 (N_11135,N_9628,N_10111);
or U11136 (N_11136,N_10390,N_9015);
nand U11137 (N_11137,N_10387,N_9698);
nand U11138 (N_11138,N_9148,N_9879);
nor U11139 (N_11139,N_9855,N_10057);
nor U11140 (N_11140,N_10302,N_9124);
nor U11141 (N_11141,N_9394,N_9315);
nand U11142 (N_11142,N_10191,N_9286);
nand U11143 (N_11143,N_9675,N_9987);
or U11144 (N_11144,N_9938,N_9871);
and U11145 (N_11145,N_9245,N_10074);
and U11146 (N_11146,N_9150,N_9916);
nor U11147 (N_11147,N_9287,N_10007);
nor U11148 (N_11148,N_9784,N_9002);
or U11149 (N_11149,N_9262,N_9741);
nor U11150 (N_11150,N_10235,N_9229);
nor U11151 (N_11151,N_10159,N_10402);
nor U11152 (N_11152,N_9781,N_9896);
nand U11153 (N_11153,N_9046,N_9903);
and U11154 (N_11154,N_9843,N_9721);
or U11155 (N_11155,N_9560,N_9162);
nor U11156 (N_11156,N_9670,N_9534);
nor U11157 (N_11157,N_9371,N_9759);
and U11158 (N_11158,N_9966,N_9875);
xor U11159 (N_11159,N_9658,N_9353);
and U11160 (N_11160,N_10290,N_9612);
nand U11161 (N_11161,N_9182,N_9706);
nor U11162 (N_11162,N_9396,N_9944);
nand U11163 (N_11163,N_9726,N_10371);
nor U11164 (N_11164,N_10160,N_9375);
nand U11165 (N_11165,N_10327,N_9601);
and U11166 (N_11166,N_10295,N_9244);
or U11167 (N_11167,N_9385,N_9392);
or U11168 (N_11168,N_10287,N_9281);
and U11169 (N_11169,N_9379,N_9409);
nor U11170 (N_11170,N_9893,N_10263);
nand U11171 (N_11171,N_9545,N_9551);
and U11172 (N_11172,N_10155,N_10211);
or U11173 (N_11173,N_9504,N_10184);
nor U11174 (N_11174,N_9510,N_9078);
and U11175 (N_11175,N_10148,N_10047);
or U11176 (N_11176,N_10229,N_9594);
or U11177 (N_11177,N_9845,N_10247);
and U11178 (N_11178,N_9682,N_9960);
nand U11179 (N_11179,N_9163,N_10077);
or U11180 (N_11180,N_9290,N_9523);
and U11181 (N_11181,N_10125,N_10225);
and U11182 (N_11182,N_10399,N_9230);
nand U11183 (N_11183,N_9252,N_9834);
xnor U11184 (N_11184,N_9049,N_10246);
or U11185 (N_11185,N_9153,N_9044);
and U11186 (N_11186,N_9342,N_10056);
or U11187 (N_11187,N_10324,N_10239);
nor U11188 (N_11188,N_9967,N_9359);
nor U11189 (N_11189,N_9031,N_9446);
nor U11190 (N_11190,N_10104,N_9795);
and U11191 (N_11191,N_9208,N_9899);
and U11192 (N_11192,N_9679,N_10112);
and U11193 (N_11193,N_9289,N_9438);
and U11194 (N_11194,N_9825,N_9872);
and U11195 (N_11195,N_9603,N_9538);
or U11196 (N_11196,N_9537,N_9442);
nor U11197 (N_11197,N_9343,N_10421);
nand U11198 (N_11198,N_9887,N_9935);
or U11199 (N_11199,N_9009,N_9206);
nor U11200 (N_11200,N_10021,N_9464);
or U11201 (N_11201,N_9566,N_9849);
or U11202 (N_11202,N_9714,N_9122);
or U11203 (N_11203,N_9083,N_9521);
and U11204 (N_11204,N_9239,N_9740);
nor U11205 (N_11205,N_10075,N_10245);
nor U11206 (N_11206,N_10328,N_9657);
nand U11207 (N_11207,N_10391,N_9542);
and U11208 (N_11208,N_10284,N_10138);
nand U11209 (N_11209,N_10472,N_10357);
nand U11210 (N_11210,N_10431,N_9591);
nand U11211 (N_11211,N_10022,N_9205);
and U11212 (N_11212,N_9735,N_9056);
or U11213 (N_11213,N_9526,N_10036);
nand U11214 (N_11214,N_9911,N_10455);
and U11215 (N_11215,N_9830,N_9673);
and U11216 (N_11216,N_10344,N_9511);
nor U11217 (N_11217,N_9567,N_9249);
nor U11218 (N_11218,N_10400,N_10430);
nand U11219 (N_11219,N_10031,N_10195);
nor U11220 (N_11220,N_9563,N_10241);
nand U11221 (N_11221,N_10227,N_10311);
and U11222 (N_11222,N_10145,N_9094);
nor U11223 (N_11223,N_10408,N_10024);
nand U11224 (N_11224,N_10283,N_9187);
or U11225 (N_11225,N_10439,N_9461);
or U11226 (N_11226,N_9374,N_9913);
and U11227 (N_11227,N_9753,N_9929);
and U11228 (N_11228,N_9330,N_9004);
or U11229 (N_11229,N_9054,N_9662);
nand U11230 (N_11230,N_9961,N_10291);
nor U11231 (N_11231,N_9765,N_9436);
nand U11232 (N_11232,N_10040,N_10259);
nor U11233 (N_11233,N_9138,N_9876);
nand U11234 (N_11234,N_9129,N_9328);
or U11235 (N_11235,N_9055,N_9102);
or U11236 (N_11236,N_10264,N_9533);
or U11237 (N_11237,N_10449,N_10433);
nand U11238 (N_11238,N_9217,N_9225);
and U11239 (N_11239,N_9645,N_10277);
nor U11240 (N_11240,N_9039,N_9222);
or U11241 (N_11241,N_9378,N_9284);
nand U11242 (N_11242,N_9917,N_10423);
or U11243 (N_11243,N_10126,N_10200);
and U11244 (N_11244,N_9848,N_10436);
or U11245 (N_11245,N_9091,N_9854);
or U11246 (N_11246,N_10214,N_9390);
xor U11247 (N_11247,N_10292,N_9334);
nand U11248 (N_11248,N_9506,N_10301);
nor U11249 (N_11249,N_9066,N_9200);
and U11250 (N_11250,N_9647,N_9298);
and U11251 (N_11251,N_9494,N_9179);
or U11252 (N_11252,N_10120,N_9592);
or U11253 (N_11253,N_9992,N_10113);
nand U11254 (N_11254,N_9919,N_9698);
or U11255 (N_11255,N_9559,N_10216);
nand U11256 (N_11256,N_9053,N_9666);
nor U11257 (N_11257,N_9855,N_9423);
and U11258 (N_11258,N_9240,N_9488);
nand U11259 (N_11259,N_10091,N_9696);
and U11260 (N_11260,N_9722,N_9135);
and U11261 (N_11261,N_9783,N_10267);
and U11262 (N_11262,N_10161,N_9236);
and U11263 (N_11263,N_10373,N_10191);
and U11264 (N_11264,N_10209,N_9821);
and U11265 (N_11265,N_10142,N_9466);
or U11266 (N_11266,N_9011,N_9604);
and U11267 (N_11267,N_10328,N_9649);
or U11268 (N_11268,N_10010,N_9661);
nand U11269 (N_11269,N_10403,N_9518);
and U11270 (N_11270,N_9265,N_10140);
or U11271 (N_11271,N_9872,N_10447);
xor U11272 (N_11272,N_9828,N_10210);
or U11273 (N_11273,N_10021,N_9321);
nor U11274 (N_11274,N_10230,N_10022);
nand U11275 (N_11275,N_9645,N_10493);
and U11276 (N_11276,N_10192,N_9264);
nor U11277 (N_11277,N_9494,N_9247);
or U11278 (N_11278,N_9634,N_9288);
and U11279 (N_11279,N_9486,N_9642);
nor U11280 (N_11280,N_10415,N_9384);
nor U11281 (N_11281,N_10183,N_10392);
nand U11282 (N_11282,N_10465,N_9876);
nor U11283 (N_11283,N_10178,N_9900);
or U11284 (N_11284,N_9260,N_9224);
nand U11285 (N_11285,N_9812,N_9336);
nand U11286 (N_11286,N_10113,N_9526);
and U11287 (N_11287,N_9312,N_9665);
and U11288 (N_11288,N_9984,N_10079);
and U11289 (N_11289,N_9873,N_10498);
or U11290 (N_11290,N_9792,N_10323);
or U11291 (N_11291,N_10232,N_9017);
nand U11292 (N_11292,N_9244,N_9998);
nor U11293 (N_11293,N_9929,N_9915);
and U11294 (N_11294,N_9118,N_9725);
xnor U11295 (N_11295,N_10176,N_9677);
and U11296 (N_11296,N_9622,N_9274);
or U11297 (N_11297,N_10437,N_9887);
and U11298 (N_11298,N_9312,N_9478);
or U11299 (N_11299,N_9855,N_9527);
nand U11300 (N_11300,N_9738,N_10314);
and U11301 (N_11301,N_9263,N_9102);
and U11302 (N_11302,N_9498,N_9290);
and U11303 (N_11303,N_9699,N_9590);
or U11304 (N_11304,N_10294,N_9843);
or U11305 (N_11305,N_9444,N_10407);
xnor U11306 (N_11306,N_10302,N_9433);
and U11307 (N_11307,N_10405,N_9299);
nand U11308 (N_11308,N_10076,N_9493);
or U11309 (N_11309,N_9796,N_9916);
or U11310 (N_11310,N_9979,N_9994);
or U11311 (N_11311,N_10041,N_9946);
nand U11312 (N_11312,N_9105,N_9599);
nor U11313 (N_11313,N_10464,N_10389);
and U11314 (N_11314,N_10282,N_9748);
nor U11315 (N_11315,N_9506,N_10310);
nor U11316 (N_11316,N_9270,N_10141);
nand U11317 (N_11317,N_10228,N_10315);
and U11318 (N_11318,N_9416,N_9665);
and U11319 (N_11319,N_10252,N_9492);
and U11320 (N_11320,N_9811,N_10482);
nor U11321 (N_11321,N_9053,N_10175);
or U11322 (N_11322,N_10311,N_10344);
or U11323 (N_11323,N_9473,N_9171);
or U11324 (N_11324,N_10175,N_9244);
nor U11325 (N_11325,N_9492,N_10286);
nand U11326 (N_11326,N_9176,N_9011);
or U11327 (N_11327,N_9971,N_10280);
or U11328 (N_11328,N_9055,N_9312);
and U11329 (N_11329,N_9703,N_10481);
or U11330 (N_11330,N_9829,N_9784);
or U11331 (N_11331,N_9544,N_9513);
nand U11332 (N_11332,N_9652,N_10421);
xor U11333 (N_11333,N_9272,N_9807);
nand U11334 (N_11334,N_9094,N_9679);
nand U11335 (N_11335,N_10221,N_10132);
and U11336 (N_11336,N_9719,N_10483);
or U11337 (N_11337,N_9811,N_9873);
or U11338 (N_11338,N_10234,N_9954);
nand U11339 (N_11339,N_10320,N_10232);
and U11340 (N_11340,N_9288,N_9022);
nor U11341 (N_11341,N_9330,N_10177);
nand U11342 (N_11342,N_9902,N_9202);
or U11343 (N_11343,N_9340,N_9016);
xor U11344 (N_11344,N_9128,N_9459);
nor U11345 (N_11345,N_9988,N_9166);
and U11346 (N_11346,N_10354,N_9618);
nor U11347 (N_11347,N_9363,N_9358);
nor U11348 (N_11348,N_10002,N_10243);
nor U11349 (N_11349,N_9443,N_10337);
and U11350 (N_11350,N_9916,N_9494);
or U11351 (N_11351,N_10216,N_9184);
or U11352 (N_11352,N_9188,N_9641);
and U11353 (N_11353,N_9803,N_9065);
nor U11354 (N_11354,N_9258,N_9666);
nand U11355 (N_11355,N_9403,N_10280);
or U11356 (N_11356,N_9274,N_9172);
nand U11357 (N_11357,N_9768,N_9347);
nand U11358 (N_11358,N_9927,N_10047);
and U11359 (N_11359,N_9923,N_9822);
nand U11360 (N_11360,N_9238,N_9734);
and U11361 (N_11361,N_10207,N_9159);
or U11362 (N_11362,N_9253,N_9506);
or U11363 (N_11363,N_9103,N_9911);
nand U11364 (N_11364,N_10244,N_10384);
nand U11365 (N_11365,N_9799,N_9394);
and U11366 (N_11366,N_9918,N_10325);
nor U11367 (N_11367,N_10068,N_9061);
or U11368 (N_11368,N_9848,N_9039);
nand U11369 (N_11369,N_9197,N_9874);
or U11370 (N_11370,N_10148,N_10403);
nand U11371 (N_11371,N_9449,N_10373);
and U11372 (N_11372,N_9478,N_9261);
and U11373 (N_11373,N_9495,N_9871);
and U11374 (N_11374,N_9130,N_9021);
or U11375 (N_11375,N_9318,N_9486);
or U11376 (N_11376,N_9878,N_9332);
nand U11377 (N_11377,N_10411,N_9971);
nor U11378 (N_11378,N_9500,N_9335);
or U11379 (N_11379,N_9483,N_10157);
and U11380 (N_11380,N_9148,N_9825);
nand U11381 (N_11381,N_9227,N_10085);
nor U11382 (N_11382,N_9520,N_9736);
or U11383 (N_11383,N_9187,N_9912);
nand U11384 (N_11384,N_10363,N_10387);
or U11385 (N_11385,N_9623,N_9391);
nand U11386 (N_11386,N_9559,N_9651);
or U11387 (N_11387,N_9684,N_10376);
and U11388 (N_11388,N_9941,N_10267);
nor U11389 (N_11389,N_10406,N_10434);
nor U11390 (N_11390,N_9738,N_9181);
and U11391 (N_11391,N_9434,N_10199);
nor U11392 (N_11392,N_9151,N_9461);
or U11393 (N_11393,N_9859,N_9278);
nand U11394 (N_11394,N_9931,N_9373);
nor U11395 (N_11395,N_10272,N_9178);
nand U11396 (N_11396,N_9797,N_10170);
nand U11397 (N_11397,N_9763,N_10424);
or U11398 (N_11398,N_10071,N_10274);
or U11399 (N_11399,N_10084,N_10246);
or U11400 (N_11400,N_9834,N_10061);
nand U11401 (N_11401,N_9223,N_9068);
nand U11402 (N_11402,N_9955,N_9823);
and U11403 (N_11403,N_9545,N_9146);
or U11404 (N_11404,N_9778,N_9674);
nor U11405 (N_11405,N_9113,N_10473);
or U11406 (N_11406,N_9730,N_9240);
and U11407 (N_11407,N_9479,N_9385);
or U11408 (N_11408,N_9813,N_10014);
and U11409 (N_11409,N_9912,N_9231);
nand U11410 (N_11410,N_9819,N_9814);
nor U11411 (N_11411,N_9638,N_9456);
nand U11412 (N_11412,N_9919,N_9790);
and U11413 (N_11413,N_10425,N_9290);
or U11414 (N_11414,N_9814,N_10093);
or U11415 (N_11415,N_9766,N_10357);
nor U11416 (N_11416,N_9325,N_9404);
or U11417 (N_11417,N_9637,N_10316);
nand U11418 (N_11418,N_9226,N_9592);
or U11419 (N_11419,N_9618,N_9044);
or U11420 (N_11420,N_9881,N_9648);
nor U11421 (N_11421,N_9352,N_9465);
and U11422 (N_11422,N_10409,N_9255);
and U11423 (N_11423,N_10156,N_9973);
and U11424 (N_11424,N_9580,N_9855);
nand U11425 (N_11425,N_10360,N_9939);
nor U11426 (N_11426,N_10004,N_10412);
or U11427 (N_11427,N_10024,N_9279);
nor U11428 (N_11428,N_10459,N_10121);
nor U11429 (N_11429,N_10314,N_10340);
xnor U11430 (N_11430,N_10204,N_9205);
nand U11431 (N_11431,N_9490,N_9035);
nand U11432 (N_11432,N_9339,N_10307);
and U11433 (N_11433,N_9936,N_10026);
and U11434 (N_11434,N_9795,N_9108);
and U11435 (N_11435,N_9268,N_9069);
or U11436 (N_11436,N_9980,N_10277);
nand U11437 (N_11437,N_9158,N_10167);
or U11438 (N_11438,N_9764,N_9651);
nor U11439 (N_11439,N_9120,N_9656);
and U11440 (N_11440,N_10193,N_10316);
and U11441 (N_11441,N_9613,N_9361);
nand U11442 (N_11442,N_10233,N_9874);
nand U11443 (N_11443,N_9653,N_9625);
nor U11444 (N_11444,N_9116,N_9319);
nand U11445 (N_11445,N_10377,N_9258);
nor U11446 (N_11446,N_10495,N_9711);
nand U11447 (N_11447,N_9665,N_9947);
nor U11448 (N_11448,N_9986,N_9232);
or U11449 (N_11449,N_9637,N_9044);
nand U11450 (N_11450,N_10390,N_10043);
and U11451 (N_11451,N_10485,N_10078);
nand U11452 (N_11452,N_10381,N_9677);
nand U11453 (N_11453,N_9855,N_9641);
or U11454 (N_11454,N_9720,N_10223);
nor U11455 (N_11455,N_9621,N_10494);
or U11456 (N_11456,N_9203,N_10148);
and U11457 (N_11457,N_9490,N_10318);
or U11458 (N_11458,N_9278,N_9441);
nor U11459 (N_11459,N_9874,N_9116);
nand U11460 (N_11460,N_10344,N_10227);
nand U11461 (N_11461,N_9942,N_9605);
or U11462 (N_11462,N_9503,N_9446);
nand U11463 (N_11463,N_10346,N_9908);
and U11464 (N_11464,N_10134,N_10059);
nand U11465 (N_11465,N_10378,N_9488);
and U11466 (N_11466,N_9447,N_9196);
nor U11467 (N_11467,N_9445,N_9775);
nand U11468 (N_11468,N_9777,N_10360);
or U11469 (N_11469,N_10241,N_9136);
nand U11470 (N_11470,N_10312,N_9230);
nor U11471 (N_11471,N_10213,N_10138);
or U11472 (N_11472,N_10496,N_9264);
or U11473 (N_11473,N_10131,N_9855);
nor U11474 (N_11474,N_9371,N_9994);
nand U11475 (N_11475,N_10241,N_9649);
or U11476 (N_11476,N_9018,N_9649);
nand U11477 (N_11477,N_10301,N_9363);
xor U11478 (N_11478,N_10390,N_10084);
and U11479 (N_11479,N_9931,N_9178);
nor U11480 (N_11480,N_9714,N_9516);
nor U11481 (N_11481,N_9980,N_9866);
and U11482 (N_11482,N_9867,N_10142);
or U11483 (N_11483,N_9158,N_9502);
or U11484 (N_11484,N_10203,N_10498);
and U11485 (N_11485,N_9825,N_9138);
nor U11486 (N_11486,N_9174,N_9035);
and U11487 (N_11487,N_9314,N_10213);
and U11488 (N_11488,N_9552,N_9566);
or U11489 (N_11489,N_9580,N_9019);
and U11490 (N_11490,N_9181,N_10410);
nand U11491 (N_11491,N_10022,N_9836);
nand U11492 (N_11492,N_10413,N_9798);
and U11493 (N_11493,N_9797,N_9739);
and U11494 (N_11494,N_9836,N_9802);
and U11495 (N_11495,N_10368,N_9791);
nor U11496 (N_11496,N_10152,N_9371);
or U11497 (N_11497,N_10182,N_9895);
nand U11498 (N_11498,N_10445,N_9468);
and U11499 (N_11499,N_9092,N_9551);
or U11500 (N_11500,N_9640,N_10026);
nand U11501 (N_11501,N_9563,N_9640);
and U11502 (N_11502,N_10226,N_10386);
or U11503 (N_11503,N_9143,N_10429);
nand U11504 (N_11504,N_9102,N_9490);
nor U11505 (N_11505,N_10324,N_9677);
and U11506 (N_11506,N_9188,N_10315);
nor U11507 (N_11507,N_9739,N_9727);
nor U11508 (N_11508,N_9927,N_10417);
and U11509 (N_11509,N_10022,N_10321);
nand U11510 (N_11510,N_9931,N_9695);
or U11511 (N_11511,N_9291,N_9504);
or U11512 (N_11512,N_9298,N_9317);
and U11513 (N_11513,N_9450,N_9705);
and U11514 (N_11514,N_9247,N_9369);
or U11515 (N_11515,N_10452,N_9948);
nor U11516 (N_11516,N_9845,N_9461);
or U11517 (N_11517,N_10214,N_10057);
or U11518 (N_11518,N_10454,N_9516);
nor U11519 (N_11519,N_9100,N_9356);
or U11520 (N_11520,N_10481,N_9810);
nand U11521 (N_11521,N_10233,N_9573);
nand U11522 (N_11522,N_10030,N_9257);
nor U11523 (N_11523,N_9973,N_9797);
or U11524 (N_11524,N_9373,N_9690);
and U11525 (N_11525,N_9373,N_10361);
nor U11526 (N_11526,N_9146,N_10073);
nor U11527 (N_11527,N_9258,N_10298);
or U11528 (N_11528,N_9005,N_9346);
or U11529 (N_11529,N_10051,N_9930);
nand U11530 (N_11530,N_9705,N_9704);
nor U11531 (N_11531,N_10365,N_10362);
and U11532 (N_11532,N_9558,N_9504);
and U11533 (N_11533,N_9132,N_9005);
and U11534 (N_11534,N_9436,N_9355);
and U11535 (N_11535,N_10218,N_9353);
nor U11536 (N_11536,N_9414,N_9333);
nand U11537 (N_11537,N_9709,N_10216);
nor U11538 (N_11538,N_9102,N_9408);
nand U11539 (N_11539,N_9679,N_9454);
nor U11540 (N_11540,N_9642,N_10365);
or U11541 (N_11541,N_9348,N_9421);
nand U11542 (N_11542,N_10396,N_9131);
or U11543 (N_11543,N_9089,N_10333);
nand U11544 (N_11544,N_10071,N_9139);
and U11545 (N_11545,N_9432,N_9632);
nor U11546 (N_11546,N_9362,N_9501);
or U11547 (N_11547,N_9836,N_10200);
and U11548 (N_11548,N_10048,N_9680);
nand U11549 (N_11549,N_10413,N_10343);
and U11550 (N_11550,N_9040,N_10379);
or U11551 (N_11551,N_9377,N_9292);
nor U11552 (N_11552,N_9149,N_9017);
and U11553 (N_11553,N_10373,N_9264);
and U11554 (N_11554,N_9324,N_9757);
and U11555 (N_11555,N_9280,N_9408);
xnor U11556 (N_11556,N_9773,N_10250);
and U11557 (N_11557,N_9872,N_9119);
nand U11558 (N_11558,N_9683,N_9961);
nor U11559 (N_11559,N_10042,N_9135);
or U11560 (N_11560,N_9257,N_10170);
or U11561 (N_11561,N_9851,N_10048);
and U11562 (N_11562,N_10242,N_9043);
nand U11563 (N_11563,N_9746,N_9095);
nor U11564 (N_11564,N_10169,N_10268);
and U11565 (N_11565,N_9724,N_10302);
nor U11566 (N_11566,N_9625,N_9490);
xnor U11567 (N_11567,N_10301,N_9525);
and U11568 (N_11568,N_10263,N_10417);
and U11569 (N_11569,N_10075,N_9954);
and U11570 (N_11570,N_9864,N_10087);
and U11571 (N_11571,N_10254,N_9815);
or U11572 (N_11572,N_9497,N_10418);
nor U11573 (N_11573,N_10043,N_9492);
or U11574 (N_11574,N_9976,N_10046);
nand U11575 (N_11575,N_10290,N_9093);
nand U11576 (N_11576,N_9594,N_9838);
or U11577 (N_11577,N_10444,N_9501);
nand U11578 (N_11578,N_9850,N_9424);
nand U11579 (N_11579,N_10041,N_9526);
and U11580 (N_11580,N_9885,N_10359);
nor U11581 (N_11581,N_9580,N_9795);
nor U11582 (N_11582,N_10060,N_9167);
and U11583 (N_11583,N_10121,N_9106);
nor U11584 (N_11584,N_9624,N_9911);
and U11585 (N_11585,N_10212,N_9194);
nand U11586 (N_11586,N_10172,N_9172);
nor U11587 (N_11587,N_10395,N_10372);
nand U11588 (N_11588,N_10085,N_10173);
nor U11589 (N_11589,N_10407,N_9889);
nand U11590 (N_11590,N_10182,N_9332);
and U11591 (N_11591,N_9486,N_10038);
nand U11592 (N_11592,N_10123,N_9947);
nor U11593 (N_11593,N_9915,N_10087);
nand U11594 (N_11594,N_9266,N_9618);
nand U11595 (N_11595,N_9425,N_10136);
or U11596 (N_11596,N_9994,N_10481);
nand U11597 (N_11597,N_9425,N_9198);
nand U11598 (N_11598,N_9533,N_10263);
nand U11599 (N_11599,N_9445,N_9123);
and U11600 (N_11600,N_10262,N_10209);
nand U11601 (N_11601,N_9876,N_9253);
nor U11602 (N_11602,N_9464,N_10154);
or U11603 (N_11603,N_9785,N_9948);
and U11604 (N_11604,N_10371,N_9928);
nor U11605 (N_11605,N_10367,N_9329);
or U11606 (N_11606,N_9266,N_10303);
and U11607 (N_11607,N_10344,N_9539);
or U11608 (N_11608,N_9439,N_9781);
nor U11609 (N_11609,N_9532,N_9849);
and U11610 (N_11610,N_9494,N_10168);
or U11611 (N_11611,N_9218,N_9850);
nor U11612 (N_11612,N_9813,N_9319);
and U11613 (N_11613,N_10007,N_9130);
nor U11614 (N_11614,N_10492,N_9649);
and U11615 (N_11615,N_9995,N_10015);
nand U11616 (N_11616,N_10195,N_9972);
nand U11617 (N_11617,N_9686,N_9870);
nand U11618 (N_11618,N_9776,N_9908);
and U11619 (N_11619,N_10459,N_9136);
or U11620 (N_11620,N_9847,N_10185);
nand U11621 (N_11621,N_10441,N_10174);
xnor U11622 (N_11622,N_10245,N_9878);
and U11623 (N_11623,N_9643,N_10247);
and U11624 (N_11624,N_9646,N_9533);
nor U11625 (N_11625,N_9517,N_9285);
and U11626 (N_11626,N_9131,N_10442);
nand U11627 (N_11627,N_10058,N_9848);
nor U11628 (N_11628,N_10398,N_9183);
and U11629 (N_11629,N_9360,N_9310);
and U11630 (N_11630,N_9516,N_9883);
nand U11631 (N_11631,N_9935,N_9326);
or U11632 (N_11632,N_10440,N_10377);
xnor U11633 (N_11633,N_9482,N_9257);
and U11634 (N_11634,N_10433,N_9962);
nand U11635 (N_11635,N_9874,N_9023);
nor U11636 (N_11636,N_10399,N_9307);
nor U11637 (N_11637,N_9855,N_9592);
nor U11638 (N_11638,N_9966,N_10003);
or U11639 (N_11639,N_9819,N_9026);
nor U11640 (N_11640,N_9550,N_9072);
nand U11641 (N_11641,N_9964,N_9004);
and U11642 (N_11642,N_10378,N_9874);
nand U11643 (N_11643,N_9938,N_9844);
nor U11644 (N_11644,N_9265,N_10027);
nand U11645 (N_11645,N_10186,N_9856);
nor U11646 (N_11646,N_9315,N_9551);
or U11647 (N_11647,N_9913,N_9651);
nor U11648 (N_11648,N_10306,N_9791);
nand U11649 (N_11649,N_9752,N_10334);
nand U11650 (N_11650,N_10115,N_9482);
nor U11651 (N_11651,N_10301,N_10456);
nor U11652 (N_11652,N_9097,N_9341);
nand U11653 (N_11653,N_9690,N_10266);
or U11654 (N_11654,N_9104,N_9965);
and U11655 (N_11655,N_10293,N_9408);
and U11656 (N_11656,N_9960,N_9428);
nor U11657 (N_11657,N_10362,N_10169);
and U11658 (N_11658,N_9159,N_10071);
nor U11659 (N_11659,N_9024,N_10294);
or U11660 (N_11660,N_9436,N_9001);
nand U11661 (N_11661,N_9153,N_9465);
or U11662 (N_11662,N_10428,N_9558);
nand U11663 (N_11663,N_9134,N_9872);
nor U11664 (N_11664,N_9348,N_9514);
nor U11665 (N_11665,N_9748,N_10115);
nor U11666 (N_11666,N_10008,N_10328);
nand U11667 (N_11667,N_10090,N_10427);
nand U11668 (N_11668,N_9538,N_9262);
nand U11669 (N_11669,N_9946,N_9423);
nand U11670 (N_11670,N_10001,N_9503);
and U11671 (N_11671,N_9572,N_10206);
nor U11672 (N_11672,N_9875,N_10104);
and U11673 (N_11673,N_9933,N_9014);
and U11674 (N_11674,N_9411,N_10218);
nor U11675 (N_11675,N_9013,N_10172);
nor U11676 (N_11676,N_9683,N_10315);
nor U11677 (N_11677,N_9659,N_9235);
and U11678 (N_11678,N_9162,N_10169);
nand U11679 (N_11679,N_10491,N_9256);
and U11680 (N_11680,N_9100,N_9832);
or U11681 (N_11681,N_9068,N_9887);
nor U11682 (N_11682,N_10394,N_9497);
or U11683 (N_11683,N_9501,N_9624);
and U11684 (N_11684,N_9252,N_9212);
or U11685 (N_11685,N_10320,N_9684);
nor U11686 (N_11686,N_9761,N_9292);
nor U11687 (N_11687,N_9869,N_9475);
nand U11688 (N_11688,N_9970,N_10199);
and U11689 (N_11689,N_9755,N_10045);
nand U11690 (N_11690,N_10132,N_9376);
nor U11691 (N_11691,N_9170,N_10005);
nor U11692 (N_11692,N_9942,N_9683);
and U11693 (N_11693,N_9678,N_9209);
nand U11694 (N_11694,N_9189,N_10199);
nor U11695 (N_11695,N_9803,N_10118);
or U11696 (N_11696,N_10252,N_9195);
nand U11697 (N_11697,N_10363,N_9603);
nand U11698 (N_11698,N_10215,N_10204);
or U11699 (N_11699,N_10223,N_10369);
and U11700 (N_11700,N_10210,N_10133);
and U11701 (N_11701,N_10125,N_10047);
and U11702 (N_11702,N_9117,N_9497);
nor U11703 (N_11703,N_9609,N_9498);
or U11704 (N_11704,N_9503,N_9693);
or U11705 (N_11705,N_9026,N_9312);
or U11706 (N_11706,N_9705,N_10312);
nand U11707 (N_11707,N_9940,N_10318);
nand U11708 (N_11708,N_9256,N_9330);
nand U11709 (N_11709,N_9562,N_9667);
and U11710 (N_11710,N_9037,N_9330);
nand U11711 (N_11711,N_10449,N_9402);
and U11712 (N_11712,N_9145,N_9344);
or U11713 (N_11713,N_10067,N_9095);
or U11714 (N_11714,N_9038,N_9977);
nand U11715 (N_11715,N_9040,N_9334);
nor U11716 (N_11716,N_9640,N_9585);
and U11717 (N_11717,N_10189,N_9025);
nor U11718 (N_11718,N_9160,N_9487);
or U11719 (N_11719,N_9794,N_9136);
nor U11720 (N_11720,N_9887,N_9383);
and U11721 (N_11721,N_9444,N_9662);
nand U11722 (N_11722,N_9745,N_10305);
nand U11723 (N_11723,N_10201,N_10257);
and U11724 (N_11724,N_9171,N_9525);
nand U11725 (N_11725,N_9539,N_10391);
nor U11726 (N_11726,N_9828,N_10200);
or U11727 (N_11727,N_9553,N_9299);
or U11728 (N_11728,N_10328,N_9068);
nor U11729 (N_11729,N_9273,N_10074);
nor U11730 (N_11730,N_10042,N_9682);
and U11731 (N_11731,N_10386,N_9110);
or U11732 (N_11732,N_10225,N_9756);
and U11733 (N_11733,N_9750,N_9896);
nand U11734 (N_11734,N_9800,N_9727);
or U11735 (N_11735,N_9877,N_9563);
or U11736 (N_11736,N_9159,N_10164);
nand U11737 (N_11737,N_9098,N_10076);
xor U11738 (N_11738,N_9760,N_9444);
nand U11739 (N_11739,N_9102,N_10475);
nand U11740 (N_11740,N_9156,N_10492);
or U11741 (N_11741,N_9893,N_10087);
or U11742 (N_11742,N_9683,N_9687);
or U11743 (N_11743,N_10135,N_9497);
or U11744 (N_11744,N_9414,N_9263);
nor U11745 (N_11745,N_10328,N_9584);
or U11746 (N_11746,N_9436,N_10399);
and U11747 (N_11747,N_9759,N_10146);
or U11748 (N_11748,N_9453,N_9299);
nor U11749 (N_11749,N_10040,N_9033);
or U11750 (N_11750,N_9876,N_9317);
and U11751 (N_11751,N_10188,N_10320);
nor U11752 (N_11752,N_9647,N_10366);
and U11753 (N_11753,N_10453,N_9889);
and U11754 (N_11754,N_10117,N_9291);
and U11755 (N_11755,N_10191,N_9681);
nand U11756 (N_11756,N_9394,N_9631);
and U11757 (N_11757,N_9794,N_10431);
or U11758 (N_11758,N_9314,N_9246);
nand U11759 (N_11759,N_10011,N_10185);
nor U11760 (N_11760,N_9059,N_9782);
nor U11761 (N_11761,N_9233,N_10416);
nor U11762 (N_11762,N_9084,N_9537);
nor U11763 (N_11763,N_9527,N_9207);
or U11764 (N_11764,N_9680,N_9748);
or U11765 (N_11765,N_10429,N_9886);
or U11766 (N_11766,N_10223,N_10304);
nand U11767 (N_11767,N_9138,N_10114);
and U11768 (N_11768,N_9012,N_10001);
and U11769 (N_11769,N_10267,N_9167);
or U11770 (N_11770,N_10130,N_9669);
or U11771 (N_11771,N_10212,N_9255);
or U11772 (N_11772,N_9041,N_9218);
or U11773 (N_11773,N_10363,N_9106);
or U11774 (N_11774,N_9551,N_9033);
or U11775 (N_11775,N_9073,N_9963);
and U11776 (N_11776,N_9772,N_9161);
and U11777 (N_11777,N_10163,N_9820);
nand U11778 (N_11778,N_9980,N_9673);
nand U11779 (N_11779,N_9968,N_10012);
or U11780 (N_11780,N_9917,N_10137);
or U11781 (N_11781,N_9151,N_9716);
nor U11782 (N_11782,N_10474,N_10497);
or U11783 (N_11783,N_9934,N_9886);
and U11784 (N_11784,N_9394,N_10230);
nor U11785 (N_11785,N_9371,N_10129);
or U11786 (N_11786,N_10366,N_9225);
and U11787 (N_11787,N_10234,N_9778);
nor U11788 (N_11788,N_10245,N_10470);
and U11789 (N_11789,N_9794,N_10404);
nor U11790 (N_11790,N_9848,N_9449);
and U11791 (N_11791,N_9994,N_10086);
and U11792 (N_11792,N_9277,N_9302);
nor U11793 (N_11793,N_9102,N_10209);
nand U11794 (N_11794,N_9033,N_9686);
nand U11795 (N_11795,N_9040,N_10238);
nor U11796 (N_11796,N_10300,N_9142);
nand U11797 (N_11797,N_9881,N_9345);
or U11798 (N_11798,N_10249,N_9492);
nand U11799 (N_11799,N_9715,N_9745);
nand U11800 (N_11800,N_9124,N_9513);
and U11801 (N_11801,N_10130,N_9650);
and U11802 (N_11802,N_9085,N_10425);
or U11803 (N_11803,N_10034,N_9961);
and U11804 (N_11804,N_9158,N_9948);
nor U11805 (N_11805,N_9065,N_9862);
or U11806 (N_11806,N_9945,N_9208);
nand U11807 (N_11807,N_10299,N_9647);
and U11808 (N_11808,N_10405,N_9903);
and U11809 (N_11809,N_9800,N_9209);
or U11810 (N_11810,N_9437,N_9747);
nor U11811 (N_11811,N_9654,N_9808);
or U11812 (N_11812,N_9983,N_9503);
or U11813 (N_11813,N_9943,N_9791);
and U11814 (N_11814,N_9653,N_9237);
nor U11815 (N_11815,N_9787,N_9114);
nor U11816 (N_11816,N_9174,N_9658);
or U11817 (N_11817,N_10380,N_9401);
or U11818 (N_11818,N_10256,N_9101);
nand U11819 (N_11819,N_9823,N_10261);
nand U11820 (N_11820,N_10384,N_9891);
or U11821 (N_11821,N_9556,N_9199);
or U11822 (N_11822,N_9572,N_10158);
or U11823 (N_11823,N_9834,N_9371);
and U11824 (N_11824,N_9097,N_10022);
or U11825 (N_11825,N_10047,N_10114);
or U11826 (N_11826,N_9880,N_10465);
or U11827 (N_11827,N_9958,N_10216);
nand U11828 (N_11828,N_9469,N_10197);
nand U11829 (N_11829,N_10253,N_9997);
nand U11830 (N_11830,N_9434,N_10046);
and U11831 (N_11831,N_9298,N_9001);
and U11832 (N_11832,N_9305,N_9197);
nand U11833 (N_11833,N_10065,N_9036);
nor U11834 (N_11834,N_9838,N_10482);
and U11835 (N_11835,N_9267,N_10275);
nor U11836 (N_11836,N_9593,N_9321);
and U11837 (N_11837,N_9737,N_9043);
nand U11838 (N_11838,N_10024,N_9488);
and U11839 (N_11839,N_10435,N_9048);
nor U11840 (N_11840,N_9272,N_9187);
nand U11841 (N_11841,N_9210,N_9154);
and U11842 (N_11842,N_9134,N_9506);
nor U11843 (N_11843,N_9713,N_9159);
nor U11844 (N_11844,N_9301,N_10405);
and U11845 (N_11845,N_9886,N_9013);
nor U11846 (N_11846,N_9785,N_10403);
nor U11847 (N_11847,N_9682,N_9763);
nor U11848 (N_11848,N_9004,N_10462);
and U11849 (N_11849,N_9608,N_9977);
nand U11850 (N_11850,N_9153,N_9642);
nand U11851 (N_11851,N_9779,N_9612);
or U11852 (N_11852,N_10284,N_9883);
nor U11853 (N_11853,N_9790,N_9874);
nor U11854 (N_11854,N_9936,N_9961);
nand U11855 (N_11855,N_9071,N_10360);
nor U11856 (N_11856,N_10241,N_9359);
nor U11857 (N_11857,N_10319,N_9168);
nor U11858 (N_11858,N_9378,N_9400);
nor U11859 (N_11859,N_9762,N_9743);
and U11860 (N_11860,N_10486,N_9460);
nor U11861 (N_11861,N_9771,N_9153);
nor U11862 (N_11862,N_10187,N_10216);
or U11863 (N_11863,N_10284,N_9215);
nand U11864 (N_11864,N_10499,N_10101);
nor U11865 (N_11865,N_9714,N_9551);
and U11866 (N_11866,N_9054,N_9996);
and U11867 (N_11867,N_10377,N_9488);
nand U11868 (N_11868,N_10274,N_10288);
or U11869 (N_11869,N_10312,N_9703);
nand U11870 (N_11870,N_9268,N_9095);
nand U11871 (N_11871,N_9232,N_9201);
or U11872 (N_11872,N_10032,N_9147);
and U11873 (N_11873,N_10356,N_9400);
nand U11874 (N_11874,N_9864,N_9138);
nand U11875 (N_11875,N_9706,N_10064);
and U11876 (N_11876,N_10335,N_9929);
and U11877 (N_11877,N_9583,N_9016);
nor U11878 (N_11878,N_9542,N_9676);
or U11879 (N_11879,N_10427,N_9749);
nand U11880 (N_11880,N_10245,N_9734);
nor U11881 (N_11881,N_9241,N_9041);
nor U11882 (N_11882,N_9050,N_9667);
or U11883 (N_11883,N_10243,N_9793);
nand U11884 (N_11884,N_9367,N_9737);
or U11885 (N_11885,N_10282,N_9569);
or U11886 (N_11886,N_9787,N_9236);
nand U11887 (N_11887,N_10413,N_10140);
nand U11888 (N_11888,N_10005,N_10434);
and U11889 (N_11889,N_9897,N_10393);
nor U11890 (N_11890,N_9285,N_9691);
or U11891 (N_11891,N_10421,N_10096);
nand U11892 (N_11892,N_10314,N_9633);
or U11893 (N_11893,N_10343,N_9186);
nor U11894 (N_11894,N_9733,N_9417);
nand U11895 (N_11895,N_9057,N_10266);
nand U11896 (N_11896,N_10060,N_10383);
or U11897 (N_11897,N_9853,N_9323);
and U11898 (N_11898,N_9368,N_9513);
nand U11899 (N_11899,N_9687,N_9968);
nor U11900 (N_11900,N_10071,N_10379);
nand U11901 (N_11901,N_9989,N_9059);
nor U11902 (N_11902,N_9413,N_9063);
and U11903 (N_11903,N_9468,N_10289);
nor U11904 (N_11904,N_9814,N_9189);
nor U11905 (N_11905,N_10167,N_9729);
nor U11906 (N_11906,N_10354,N_10353);
and U11907 (N_11907,N_10334,N_9360);
and U11908 (N_11908,N_10085,N_10228);
nor U11909 (N_11909,N_9970,N_9206);
and U11910 (N_11910,N_9276,N_10400);
nor U11911 (N_11911,N_10494,N_9790);
or U11912 (N_11912,N_9806,N_9052);
and U11913 (N_11913,N_9158,N_10481);
or U11914 (N_11914,N_9474,N_9598);
nand U11915 (N_11915,N_9008,N_9524);
nand U11916 (N_11916,N_9499,N_10146);
or U11917 (N_11917,N_9468,N_9917);
nor U11918 (N_11918,N_9720,N_9754);
xor U11919 (N_11919,N_9239,N_10121);
nand U11920 (N_11920,N_10417,N_9580);
nand U11921 (N_11921,N_9034,N_9945);
or U11922 (N_11922,N_9685,N_9607);
and U11923 (N_11923,N_9614,N_9615);
nor U11924 (N_11924,N_9202,N_9783);
and U11925 (N_11925,N_10368,N_9162);
and U11926 (N_11926,N_9038,N_10009);
or U11927 (N_11927,N_9362,N_10416);
nor U11928 (N_11928,N_9776,N_9108);
nor U11929 (N_11929,N_9450,N_10290);
or U11930 (N_11930,N_9398,N_9260);
or U11931 (N_11931,N_10130,N_9834);
nand U11932 (N_11932,N_10023,N_10429);
or U11933 (N_11933,N_9833,N_10252);
nor U11934 (N_11934,N_9793,N_9546);
or U11935 (N_11935,N_9637,N_9718);
and U11936 (N_11936,N_9582,N_9423);
and U11937 (N_11937,N_10016,N_9153);
and U11938 (N_11938,N_10041,N_10223);
nand U11939 (N_11939,N_9077,N_9809);
nand U11940 (N_11940,N_9036,N_9012);
or U11941 (N_11941,N_9957,N_9675);
nor U11942 (N_11942,N_9627,N_9480);
and U11943 (N_11943,N_10303,N_9044);
and U11944 (N_11944,N_9512,N_9704);
xor U11945 (N_11945,N_10435,N_9942);
or U11946 (N_11946,N_9519,N_10444);
nor U11947 (N_11947,N_9953,N_9006);
or U11948 (N_11948,N_9949,N_10399);
and U11949 (N_11949,N_9706,N_9860);
nand U11950 (N_11950,N_10066,N_9179);
nor U11951 (N_11951,N_9503,N_9546);
and U11952 (N_11952,N_9137,N_10169);
nor U11953 (N_11953,N_9351,N_9524);
nor U11954 (N_11954,N_9819,N_9094);
nand U11955 (N_11955,N_9747,N_10432);
and U11956 (N_11956,N_9766,N_10250);
nor U11957 (N_11957,N_9470,N_9967);
nor U11958 (N_11958,N_10060,N_9252);
or U11959 (N_11959,N_10367,N_10118);
nand U11960 (N_11960,N_9882,N_9941);
nand U11961 (N_11961,N_10110,N_9301);
and U11962 (N_11962,N_9428,N_10117);
and U11963 (N_11963,N_10320,N_9777);
and U11964 (N_11964,N_9373,N_9535);
nor U11965 (N_11965,N_10344,N_9026);
and U11966 (N_11966,N_9092,N_9392);
and U11967 (N_11967,N_9965,N_9163);
nand U11968 (N_11968,N_9362,N_9922);
and U11969 (N_11969,N_10033,N_10200);
nor U11970 (N_11970,N_9367,N_9138);
or U11971 (N_11971,N_9637,N_9083);
nand U11972 (N_11972,N_10277,N_9332);
nand U11973 (N_11973,N_9985,N_9708);
nor U11974 (N_11974,N_9768,N_9424);
or U11975 (N_11975,N_10254,N_10487);
nand U11976 (N_11976,N_10263,N_10036);
nand U11977 (N_11977,N_10166,N_9505);
or U11978 (N_11978,N_9580,N_9746);
or U11979 (N_11979,N_9352,N_9063);
and U11980 (N_11980,N_9426,N_9458);
nor U11981 (N_11981,N_10206,N_9250);
nand U11982 (N_11982,N_9793,N_9979);
nand U11983 (N_11983,N_9402,N_9982);
and U11984 (N_11984,N_9096,N_10305);
and U11985 (N_11985,N_9636,N_10247);
nor U11986 (N_11986,N_10242,N_10251);
nand U11987 (N_11987,N_9267,N_10430);
nor U11988 (N_11988,N_9619,N_9348);
nand U11989 (N_11989,N_9510,N_9319);
nand U11990 (N_11990,N_10269,N_9209);
or U11991 (N_11991,N_9899,N_9648);
and U11992 (N_11992,N_9337,N_10309);
or U11993 (N_11993,N_9581,N_10036);
nand U11994 (N_11994,N_9631,N_9419);
nand U11995 (N_11995,N_9231,N_9970);
and U11996 (N_11996,N_9982,N_9002);
and U11997 (N_11997,N_9977,N_10306);
and U11998 (N_11998,N_9239,N_10143);
or U11999 (N_11999,N_10203,N_9690);
and U12000 (N_12000,N_11333,N_11045);
nor U12001 (N_12001,N_10502,N_11811);
nor U12002 (N_12002,N_11013,N_11159);
nor U12003 (N_12003,N_10619,N_11626);
or U12004 (N_12004,N_10984,N_10683);
or U12005 (N_12005,N_11497,N_10797);
or U12006 (N_12006,N_11128,N_11971);
nor U12007 (N_12007,N_11384,N_11369);
nand U12008 (N_12008,N_11118,N_11003);
and U12009 (N_12009,N_10778,N_11817);
and U12010 (N_12010,N_10539,N_10857);
nor U12011 (N_12011,N_10662,N_11737);
or U12012 (N_12012,N_11580,N_11896);
and U12013 (N_12013,N_11078,N_11813);
and U12014 (N_12014,N_10574,N_11031);
or U12015 (N_12015,N_11995,N_10896);
nor U12016 (N_12016,N_11082,N_11177);
or U12017 (N_12017,N_11394,N_11714);
and U12018 (N_12018,N_10583,N_10565);
nand U12019 (N_12019,N_11435,N_10591);
and U12020 (N_12020,N_10518,N_10844);
or U12021 (N_12021,N_11519,N_11019);
or U12022 (N_12022,N_11994,N_11196);
or U12023 (N_12023,N_11720,N_10846);
nor U12024 (N_12024,N_10722,N_11332);
and U12025 (N_12025,N_11719,N_10986);
or U12026 (N_12026,N_10514,N_11467);
nand U12027 (N_12027,N_11047,N_11952);
or U12028 (N_12028,N_11253,N_10646);
and U12029 (N_12029,N_10859,N_11761);
nand U12030 (N_12030,N_11699,N_11595);
nand U12031 (N_12031,N_10620,N_10530);
or U12032 (N_12032,N_11404,N_11695);
or U12033 (N_12033,N_11751,N_11499);
or U12034 (N_12034,N_11429,N_11573);
and U12035 (N_12035,N_11911,N_11116);
or U12036 (N_12036,N_11053,N_11521);
and U12037 (N_12037,N_10815,N_10605);
and U12038 (N_12038,N_11001,N_10876);
nor U12039 (N_12039,N_10601,N_11703);
nand U12040 (N_12040,N_11598,N_10692);
nand U12041 (N_12041,N_11412,N_11549);
nand U12042 (N_12042,N_10682,N_11302);
nor U12043 (N_12043,N_11388,N_11924);
or U12044 (N_12044,N_11599,N_11892);
or U12045 (N_12045,N_11974,N_11740);
nand U12046 (N_12046,N_11567,N_11509);
and U12047 (N_12047,N_10705,N_10974);
and U12048 (N_12048,N_11849,N_10536);
xnor U12049 (N_12049,N_11818,N_11681);
nor U12050 (N_12050,N_11421,N_11335);
nor U12051 (N_12051,N_10871,N_11837);
or U12052 (N_12052,N_11861,N_11864);
nand U12053 (N_12053,N_11096,N_10588);
and U12054 (N_12054,N_10639,N_11209);
and U12055 (N_12055,N_11512,N_11997);
or U12056 (N_12056,N_11434,N_10660);
or U12057 (N_12057,N_10556,N_10901);
nor U12058 (N_12058,N_11713,N_10762);
nand U12059 (N_12059,N_11328,N_10863);
nand U12060 (N_12060,N_11273,N_10929);
nor U12061 (N_12061,N_11980,N_11417);
nand U12062 (N_12062,N_10575,N_11642);
and U12063 (N_12063,N_11822,N_10718);
nand U12064 (N_12064,N_11016,N_11535);
or U12065 (N_12065,N_11339,N_11688);
or U12066 (N_12066,N_11297,N_10719);
nor U12067 (N_12067,N_11073,N_11205);
or U12068 (N_12068,N_10892,N_11176);
or U12069 (N_12069,N_10845,N_10817);
nand U12070 (N_12070,N_10782,N_10586);
and U12071 (N_12071,N_11587,N_10653);
and U12072 (N_12072,N_11292,N_11092);
nand U12073 (N_12073,N_11941,N_10814);
and U12074 (N_12074,N_10763,N_11025);
or U12075 (N_12075,N_10630,N_11401);
or U12076 (N_12076,N_11189,N_11767);
or U12077 (N_12077,N_11359,N_10736);
or U12078 (N_12078,N_11743,N_11560);
nor U12079 (N_12079,N_11570,N_10663);
or U12080 (N_12080,N_11794,N_10548);
and U12081 (N_12081,N_11372,N_11242);
nand U12082 (N_12082,N_11569,N_10911);
nor U12083 (N_12083,N_10991,N_10979);
nor U12084 (N_12084,N_11330,N_11385);
nor U12085 (N_12085,N_11575,N_11261);
nor U12086 (N_12086,N_11141,N_10989);
or U12087 (N_12087,N_11825,N_10973);
nor U12088 (N_12088,N_10878,N_11250);
or U12089 (N_12089,N_11111,N_10724);
nand U12090 (N_12090,N_11789,N_10975);
and U12091 (N_12091,N_11293,N_11773);
nand U12092 (N_12092,N_10920,N_11363);
nor U12093 (N_12093,N_10573,N_11879);
nand U12094 (N_12094,N_11863,N_11915);
nand U12095 (N_12095,N_11114,N_10507);
nor U12096 (N_12096,N_10524,N_10712);
nor U12097 (N_12097,N_11286,N_11926);
or U12098 (N_12098,N_10527,N_11392);
and U12099 (N_12099,N_11156,N_11472);
nand U12100 (N_12100,N_11457,N_10790);
xor U12101 (N_12101,N_11508,N_11545);
nor U12102 (N_12102,N_11329,N_11059);
and U12103 (N_12103,N_10667,N_11393);
nand U12104 (N_12104,N_10943,N_10908);
nand U12105 (N_12105,N_11682,N_10604);
or U12106 (N_12106,N_11014,N_11083);
and U12107 (N_12107,N_10862,N_11762);
and U12108 (N_12108,N_10999,N_11677);
or U12109 (N_12109,N_11975,N_11972);
nand U12110 (N_12110,N_11913,N_10675);
and U12111 (N_12111,N_10829,N_10642);
nor U12112 (N_12112,N_10671,N_11797);
or U12113 (N_12113,N_11692,N_11364);
or U12114 (N_12114,N_11925,N_11077);
nor U12115 (N_12115,N_10884,N_10729);
or U12116 (N_12116,N_11396,N_11938);
and U12117 (N_12117,N_10950,N_10831);
nor U12118 (N_12118,N_11976,N_11462);
nor U12119 (N_12119,N_11338,N_11400);
and U12120 (N_12120,N_11481,N_11300);
and U12121 (N_12121,N_11162,N_11216);
and U12122 (N_12122,N_10776,N_10579);
nand U12123 (N_12123,N_11255,N_10633);
nor U12124 (N_12124,N_10644,N_11548);
nand U12125 (N_12125,N_10874,N_11226);
or U12126 (N_12126,N_10978,N_11653);
and U12127 (N_12127,N_11876,N_11660);
or U12128 (N_12128,N_11854,N_10664);
nand U12129 (N_12129,N_11693,N_10938);
and U12130 (N_12130,N_10750,N_11571);
nand U12131 (N_12131,N_11129,N_11288);
nand U12132 (N_12132,N_11442,N_11357);
nand U12133 (N_12133,N_11717,N_11064);
xor U12134 (N_12134,N_10947,N_11377);
nand U12135 (N_12135,N_11744,N_11781);
and U12136 (N_12136,N_10540,N_10847);
or U12137 (N_12137,N_11147,N_10504);
nor U12138 (N_12138,N_11379,N_10710);
nand U12139 (N_12139,N_11042,N_10593);
or U12140 (N_12140,N_10669,N_10657);
nor U12141 (N_12141,N_10964,N_10753);
and U12142 (N_12142,N_11314,N_10900);
and U12143 (N_12143,N_11919,N_10651);
or U12144 (N_12144,N_10515,N_11528);
and U12145 (N_12145,N_10558,N_11920);
nand U12146 (N_12146,N_11191,N_10658);
nor U12147 (N_12147,N_11436,N_11778);
or U12148 (N_12148,N_11270,N_11043);
or U12149 (N_12149,N_10632,N_11875);
or U12150 (N_12150,N_10732,N_11373);
and U12151 (N_12151,N_11175,N_10924);
or U12152 (N_12152,N_11859,N_11000);
or U12153 (N_12153,N_11865,N_10500);
nand U12154 (N_12154,N_11124,N_11468);
and U12155 (N_12155,N_11414,N_11440);
nor U12156 (N_12156,N_11904,N_10703);
xor U12157 (N_12157,N_11718,N_10802);
or U12158 (N_12158,N_11673,N_11562);
nor U12159 (N_12159,N_11893,N_11786);
or U12160 (N_12160,N_11843,N_11168);
nand U12161 (N_12161,N_10899,N_11945);
and U12162 (N_12162,N_11074,N_10550);
nand U12163 (N_12163,N_11826,N_11172);
and U12164 (N_12164,N_11476,N_11607);
and U12165 (N_12165,N_10582,N_11622);
or U12166 (N_12166,N_11011,N_11613);
nand U12167 (N_12167,N_10806,N_10925);
and U12168 (N_12168,N_11827,N_11135);
nand U12169 (N_12169,N_10873,N_10905);
nand U12170 (N_12170,N_10728,N_10656);
or U12171 (N_12171,N_11711,N_10826);
or U12172 (N_12172,N_10723,N_11221);
nor U12173 (N_12173,N_10824,N_10693);
nor U12174 (N_12174,N_11397,N_11935);
nor U12175 (N_12175,N_11685,N_11746);
or U12176 (N_12176,N_11258,N_11726);
nand U12177 (N_12177,N_11593,N_11235);
or U12178 (N_12178,N_11696,N_10785);
and U12179 (N_12179,N_10680,N_10501);
xor U12180 (N_12180,N_11728,N_11227);
nand U12181 (N_12181,N_11783,N_11006);
or U12182 (N_12182,N_11891,N_11763);
nor U12183 (N_12183,N_11670,N_10607);
nand U12184 (N_12184,N_10739,N_11679);
nor U12185 (N_12185,N_11094,N_10560);
nand U12186 (N_12186,N_11540,N_11929);
xnor U12187 (N_12187,N_10535,N_11610);
or U12188 (N_12188,N_11530,N_10903);
nand U12189 (N_12189,N_11219,N_10760);
nor U12190 (N_12190,N_11950,N_10623);
nor U12191 (N_12191,N_10807,N_11104);
nand U12192 (N_12192,N_11050,N_10870);
or U12193 (N_12193,N_11448,N_11839);
or U12194 (N_12194,N_10821,N_11170);
nor U12195 (N_12195,N_11493,N_11239);
nor U12196 (N_12196,N_11597,N_10521);
or U12197 (N_12197,N_10914,N_11039);
nor U12198 (N_12198,N_11174,N_11779);
and U12199 (N_12199,N_11782,N_10625);
and U12200 (N_12200,N_11947,N_10571);
and U12201 (N_12201,N_11590,N_11367);
nor U12202 (N_12202,N_11712,N_11061);
and U12203 (N_12203,N_11731,N_11160);
nor U12204 (N_12204,N_11858,N_11192);
and U12205 (N_12205,N_11769,N_11091);
and U12206 (N_12206,N_10505,N_11878);
nand U12207 (N_12207,N_11510,N_11171);
nand U12208 (N_12208,N_10684,N_11152);
or U12209 (N_12209,N_11868,N_11993);
or U12210 (N_12210,N_10742,N_10946);
nor U12211 (N_12211,N_11620,N_10510);
and U12212 (N_12212,N_10637,N_11999);
nand U12213 (N_12213,N_11916,N_10603);
or U12214 (N_12214,N_11466,N_11289);
or U12215 (N_12215,N_11574,N_10805);
nor U12216 (N_12216,N_11424,N_11507);
or U12217 (N_12217,N_10823,N_11028);
or U12218 (N_12218,N_11041,N_10592);
or U12219 (N_12219,N_11029,N_11139);
nand U12220 (N_12220,N_11518,N_11948);
and U12221 (N_12221,N_11634,N_11852);
and U12222 (N_12222,N_10944,N_11988);
and U12223 (N_12223,N_11121,N_11534);
or U12224 (N_12224,N_11636,N_11697);
or U12225 (N_12225,N_11882,N_10523);
nor U12226 (N_12226,N_11957,N_10688);
or U12227 (N_12227,N_10833,N_10928);
and U12228 (N_12228,N_10977,N_11841);
and U12229 (N_12229,N_11949,N_11166);
or U12230 (N_12230,N_10727,N_11986);
and U12231 (N_12231,N_11275,N_10567);
nor U12232 (N_12232,N_10600,N_11900);
or U12233 (N_12233,N_11604,N_11772);
nand U12234 (N_12234,N_10864,N_10860);
and U12235 (N_12235,N_10503,N_10696);
nand U12236 (N_12236,N_11241,N_11730);
nor U12237 (N_12237,N_11532,N_11020);
and U12238 (N_12238,N_11629,N_11867);
and U12239 (N_12239,N_11909,N_11097);
nor U12240 (N_12240,N_11109,N_11150);
and U12241 (N_12241,N_10794,N_10981);
or U12242 (N_12242,N_11155,N_10961);
or U12243 (N_12243,N_10512,N_10881);
xnor U12244 (N_12244,N_11093,N_11352);
and U12245 (N_12245,N_11350,N_11004);
and U12246 (N_12246,N_10704,N_10645);
or U12247 (N_12247,N_10725,N_10879);
nor U12248 (N_12248,N_11420,N_11299);
or U12249 (N_12249,N_11674,N_11306);
nor U12250 (N_12250,N_11021,N_11356);
or U12251 (N_12251,N_10922,N_11017);
nor U12252 (N_12252,N_11186,N_11844);
nor U12253 (N_12253,N_11551,N_10545);
nand U12254 (N_12254,N_11298,N_11054);
nor U12255 (N_12255,N_11079,N_10720);
nor U12256 (N_12256,N_10966,N_10554);
nor U12257 (N_12257,N_10906,N_11774);
and U12258 (N_12258,N_10976,N_11395);
nand U12259 (N_12259,N_10547,N_11568);
nor U12260 (N_12260,N_10990,N_11280);
or U12261 (N_12261,N_10559,N_11546);
nor U12262 (N_12262,N_10534,N_10994);
and U12263 (N_12263,N_10668,N_11458);
nor U12264 (N_12264,N_10542,N_11617);
nor U12265 (N_12265,N_11075,N_10759);
and U12266 (N_12266,N_11931,N_11832);
nand U12267 (N_12267,N_10552,N_11895);
or U12268 (N_12268,N_10855,N_11490);
or U12269 (N_12269,N_10808,N_11795);
nand U12270 (N_12270,N_11263,N_11315);
or U12271 (N_12271,N_10538,N_10549);
nand U12272 (N_12272,N_11382,N_10774);
or U12273 (N_12273,N_11203,N_10717);
or U12274 (N_12274,N_11391,N_11355);
or U12275 (N_12275,N_11724,N_11638);
or U12276 (N_12276,N_11310,N_11556);
nand U12277 (N_12277,N_10626,N_11960);
or U12278 (N_12278,N_11431,N_11552);
or U12279 (N_12279,N_10741,N_11482);
and U12280 (N_12280,N_11542,N_11643);
and U12281 (N_12281,N_11349,N_11589);
or U12282 (N_12282,N_10882,N_11183);
nor U12283 (N_12283,N_11473,N_10919);
or U12284 (N_12284,N_11577,N_11256);
or U12285 (N_12285,N_11672,N_10980);
nand U12286 (N_12286,N_10880,N_11403);
or U12287 (N_12287,N_10793,N_11759);
or U12288 (N_12288,N_11471,N_11433);
nor U12289 (N_12289,N_10764,N_10854);
nand U12290 (N_12290,N_10913,N_11234);
nand U12291 (N_12291,N_10618,N_11765);
nor U12292 (N_12292,N_11721,N_11513);
nor U12293 (N_12293,N_10945,N_10921);
or U12294 (N_12294,N_11823,N_10767);
nand U12295 (N_12295,N_11912,N_11416);
nand U12296 (N_12296,N_10949,N_10522);
nand U12297 (N_12297,N_11501,N_10963);
nand U12298 (N_12298,N_11600,N_11543);
nand U12299 (N_12299,N_10621,N_11698);
nand U12300 (N_12300,N_10751,N_10533);
nor U12301 (N_12301,N_11057,N_10590);
and U12302 (N_12302,N_11026,N_11807);
and U12303 (N_12303,N_11276,N_11821);
and U12304 (N_12304,N_11428,N_11820);
nor U12305 (N_12305,N_11007,N_11977);
and U12306 (N_12306,N_10801,N_11967);
or U12307 (N_12307,N_10714,N_11970);
and U12308 (N_12308,N_11410,N_11112);
and U12309 (N_12309,N_11491,N_11370);
nand U12310 (N_12310,N_11684,N_10756);
xor U12311 (N_12311,N_11398,N_11961);
nor U12312 (N_12312,N_11087,N_10996);
nand U12313 (N_12313,N_11866,N_11488);
nor U12314 (N_12314,N_11231,N_11855);
nor U12315 (N_12315,N_11153,N_11753);
nor U12316 (N_12316,N_11650,N_10868);
and U12317 (N_12317,N_10576,N_11405);
and U12318 (N_12318,N_10689,N_11799);
xnor U12319 (N_12319,N_11027,N_10818);
and U12320 (N_12320,N_11046,N_11954);
nand U12321 (N_12321,N_11294,N_10869);
or U12322 (N_12322,N_11873,N_11602);
or U12323 (N_12323,N_11449,N_10551);
or U12324 (N_12324,N_11343,N_10796);
and U12325 (N_12325,N_10634,N_10706);
and U12326 (N_12326,N_11103,N_11065);
nor U12327 (N_12327,N_11430,N_10789);
and U12328 (N_12328,N_11368,N_10528);
nand U12329 (N_12329,N_11951,N_11274);
or U12330 (N_12330,N_11741,N_11324);
nor U12331 (N_12331,N_10948,N_11179);
nand U12332 (N_12332,N_11898,N_11654);
nand U12333 (N_12333,N_10596,N_10754);
nor U12334 (N_12334,N_11635,N_10798);
nor U12335 (N_12335,N_11375,N_11119);
and U12336 (N_12336,N_11138,N_10609);
nand U12337 (N_12337,N_11437,N_11225);
nor U12338 (N_12338,N_10834,N_11145);
nand U12339 (N_12339,N_11584,N_11374);
and U12340 (N_12340,N_10531,N_10813);
and U12341 (N_12341,N_10895,N_11908);
and U12342 (N_12342,N_10711,N_11308);
or U12343 (N_12343,N_11644,N_10721);
and U12344 (N_12344,N_11564,N_11281);
nand U12345 (N_12345,N_11106,N_11295);
nand U12346 (N_12346,N_10792,N_10968);
and U12347 (N_12347,N_11834,N_11550);
or U12348 (N_12348,N_11283,N_10516);
nand U12349 (N_12349,N_11914,N_10838);
nand U12350 (N_12350,N_11637,N_11755);
and U12351 (N_12351,N_10569,N_11748);
nor U12352 (N_12352,N_11903,N_11591);
nand U12353 (N_12353,N_11804,N_11705);
or U12354 (N_12354,N_11130,N_11793);
or U12355 (N_12355,N_11766,N_11805);
and U12356 (N_12356,N_11100,N_10934);
xnor U12357 (N_12357,N_10936,N_10971);
or U12358 (N_12358,N_11639,N_10772);
or U12359 (N_12359,N_11102,N_11533);
or U12360 (N_12360,N_11760,N_10602);
or U12361 (N_12361,N_11022,N_11689);
and U12362 (N_12362,N_10581,N_11800);
or U12363 (N_12363,N_11701,N_10698);
or U12364 (N_12364,N_11495,N_11850);
and U12365 (N_12365,N_10595,N_11008);
nor U12366 (N_12366,N_11459,N_10923);
and U12367 (N_12367,N_11051,N_10606);
nand U12368 (N_12368,N_11030,N_11857);
or U12369 (N_12369,N_11985,N_11426);
or U12370 (N_12370,N_10781,N_11667);
nand U12371 (N_12371,N_11067,N_10636);
nand U12372 (N_12372,N_10967,N_11739);
and U12373 (N_12373,N_11002,N_11872);
nor U12374 (N_12374,N_11454,N_10932);
and U12375 (N_12375,N_11101,N_11185);
and U12376 (N_12376,N_11120,N_10768);
and U12377 (N_12377,N_11252,N_11902);
or U12378 (N_12378,N_11009,N_11956);
nand U12379 (N_12379,N_11136,N_11048);
and U12380 (N_12380,N_11631,N_11690);
nor U12381 (N_12381,N_10917,N_10532);
or U12382 (N_12382,N_11583,N_11452);
nand U12383 (N_12383,N_11215,N_11791);
and U12384 (N_12384,N_11944,N_11715);
xnor U12385 (N_12385,N_11413,N_11344);
nand U12386 (N_12386,N_10894,N_10902);
nor U12387 (N_12387,N_11337,N_11323);
and U12388 (N_12388,N_11619,N_11307);
or U12389 (N_12389,N_11489,N_11538);
and U12390 (N_12390,N_11853,N_11301);
nand U12391 (N_12391,N_10631,N_11089);
nand U12392 (N_12392,N_10962,N_11107);
and U12393 (N_12393,N_11835,N_10775);
or U12394 (N_12394,N_11646,N_11987);
nand U12395 (N_12395,N_11291,N_11611);
nand U12396 (N_12396,N_11886,N_11056);
and U12397 (N_12397,N_10942,N_10640);
and U12398 (N_12398,N_10701,N_11259);
nand U12399 (N_12399,N_11668,N_11516);
nor U12400 (N_12400,N_10677,N_11651);
and U12401 (N_12401,N_10643,N_11210);
nand U12402 (N_12402,N_11279,N_10610);
nand U12403 (N_12403,N_11080,N_10745);
nor U12404 (N_12404,N_11680,N_11784);
and U12405 (N_12405,N_10678,N_11484);
or U12406 (N_12406,N_11438,N_10877);
nand U12407 (N_12407,N_11366,N_11206);
nand U12408 (N_12408,N_11842,N_10783);
or U12409 (N_12409,N_11402,N_11733);
or U12410 (N_12410,N_11012,N_11981);
nand U12411 (N_12411,N_11918,N_11633);
or U12412 (N_12412,N_11905,N_11319);
nand U12413 (N_12413,N_11511,N_11140);
nor U12414 (N_12414,N_11143,N_11505);
nor U12415 (N_12415,N_11485,N_10852);
nor U12416 (N_12416,N_11523,N_11833);
nand U12417 (N_12417,N_10650,N_11190);
or U12418 (N_12418,N_10955,N_10679);
and U12419 (N_12419,N_11184,N_11456);
nor U12420 (N_12420,N_10506,N_11188);
or U12421 (N_12421,N_11264,N_10715);
nor U12422 (N_12422,N_11563,N_10853);
and U12423 (N_12423,N_11586,N_10766);
nand U12424 (N_12424,N_11953,N_10930);
nand U12425 (N_12425,N_11224,N_11040);
or U12426 (N_12426,N_11474,N_10562);
nand U12427 (N_12427,N_11055,N_10546);
and U12428 (N_12428,N_11326,N_11742);
nand U12429 (N_12429,N_11327,N_11345);
and U12430 (N_12430,N_11502,N_11536);
nor U12431 (N_12431,N_10841,N_11851);
and U12432 (N_12432,N_11802,N_11500);
nor U12433 (N_12433,N_11415,N_11069);
nor U12434 (N_12434,N_11038,N_11465);
and U12435 (N_12435,N_10563,N_10959);
nand U12436 (N_12436,N_11998,N_10557);
nor U12437 (N_12437,N_11110,N_11671);
nor U12438 (N_12438,N_10819,N_11716);
or U12439 (N_12439,N_11024,N_11940);
and U12440 (N_12440,N_11775,N_10707);
or U12441 (N_12441,N_11579,N_11282);
nor U12442 (N_12442,N_11325,N_11578);
and U12443 (N_12443,N_11381,N_11658);
and U12444 (N_12444,N_11444,N_11460);
nor U12445 (N_12445,N_11498,N_10992);
and U12446 (N_12446,N_10755,N_11943);
and U12447 (N_12447,N_10954,N_11445);
and U12448 (N_12448,N_10757,N_10708);
or U12449 (N_12449,N_11959,N_11645);
nand U12450 (N_12450,N_11910,N_10770);
or U12451 (N_12451,N_10803,N_11334);
nand U12452 (N_12452,N_11180,N_11142);
and U12453 (N_12453,N_11888,N_10835);
xnor U12454 (N_12454,N_10594,N_10820);
nor U12455 (N_12455,N_10952,N_11923);
nand U12456 (N_12456,N_11378,N_11194);
or U12457 (N_12457,N_11582,N_11870);
nor U12458 (N_12458,N_10743,N_10780);
or U12459 (N_12459,N_10566,N_10761);
nor U12460 (N_12460,N_10769,N_11163);
nand U12461 (N_12461,N_10887,N_11313);
nand U12462 (N_12462,N_11085,N_11230);
or U12463 (N_12463,N_11169,N_10665);
nand U12464 (N_12464,N_10825,N_11787);
and U12465 (N_12465,N_11647,N_10695);
and U12466 (N_12466,N_10773,N_10672);
and U12467 (N_12467,N_11517,N_11630);
nor U12468 (N_12468,N_11809,N_11504);
xor U12469 (N_12469,N_10740,N_11266);
and U12470 (N_12470,N_10747,N_10956);
or U12471 (N_12471,N_10843,N_11422);
or U12472 (N_12472,N_10673,N_11702);
and U12473 (N_12473,N_11871,N_11346);
nor U12474 (N_12474,N_11615,N_11088);
nand U12475 (N_12475,N_10858,N_10691);
nand U12476 (N_12476,N_10779,N_10700);
nand U12477 (N_12477,N_11249,N_11686);
nand U12478 (N_12478,N_10697,N_11113);
and U12479 (N_12479,N_11860,N_10918);
and U12480 (N_12480,N_10795,N_10733);
and U12481 (N_12481,N_10907,N_11232);
or U12482 (N_12482,N_10832,N_11164);
and U12483 (N_12483,N_10758,N_10589);
or U12484 (N_12484,N_11127,N_11808);
nor U12485 (N_12485,N_10752,N_11461);
and U12486 (N_12486,N_10970,N_11676);
or U12487 (N_12487,N_11628,N_10525);
or U12488 (N_12488,N_11389,N_10670);
or U12489 (N_12489,N_10926,N_11195);
nand U12490 (N_12490,N_11233,N_11869);
nand U12491 (N_12491,N_11907,N_11780);
nor U12492 (N_12492,N_10628,N_11322);
or U12493 (N_12493,N_11425,N_10655);
nand U12494 (N_12494,N_11887,N_10812);
nor U12495 (N_12495,N_11796,N_11627);
or U12496 (N_12496,N_10578,N_10985);
nor U12497 (N_12497,N_11487,N_11240);
nand U12498 (N_12498,N_10555,N_11470);
nor U12499 (N_12499,N_10837,N_11049);
or U12500 (N_12500,N_11084,N_10836);
or U12501 (N_12501,N_10553,N_11840);
nor U12502 (N_12502,N_10649,N_11978);
or U12503 (N_12503,N_11524,N_11483);
or U12504 (N_12504,N_10622,N_11525);
nor U12505 (N_12505,N_10866,N_11447);
and U12506 (N_12506,N_10699,N_11922);
and U12507 (N_12507,N_11515,N_11845);
nand U12508 (N_12508,N_11312,N_10685);
nand U12509 (N_12509,N_11704,N_11260);
or U12510 (N_12510,N_10840,N_11149);
nor U12511 (N_12511,N_11559,N_10509);
or U12512 (N_12512,N_10737,N_11934);
or U12513 (N_12513,N_11480,N_11657);
nor U12514 (N_12514,N_10511,N_11070);
and U12515 (N_12515,N_10580,N_11228);
nand U12516 (N_12516,N_11331,N_11181);
nor U12517 (N_12517,N_10953,N_10786);
nor U12518 (N_12518,N_11360,N_11750);
and U12519 (N_12519,N_11641,N_11899);
and U12520 (N_12520,N_11539,N_11455);
or U12521 (N_12521,N_11035,N_10951);
or U12522 (N_12522,N_11729,N_11958);
and U12523 (N_12523,N_11531,N_11664);
and U12524 (N_12524,N_11603,N_11208);
or U12525 (N_12525,N_11754,N_11063);
and U12526 (N_12526,N_11296,N_11182);
and U12527 (N_12527,N_11144,N_10957);
nand U12528 (N_12528,N_10988,N_11649);
nor U12529 (N_12529,N_11081,N_11336);
nand U12530 (N_12530,N_11847,N_11640);
and U12531 (N_12531,N_10850,N_10661);
or U12532 (N_12532,N_11555,N_11146);
nand U12533 (N_12533,N_10654,N_11752);
nor U12534 (N_12534,N_10648,N_10972);
nand U12535 (N_12535,N_11675,N_11238);
nor U12536 (N_12536,N_11200,N_11133);
or U12537 (N_12537,N_11566,N_11132);
nand U12538 (N_12538,N_11201,N_11451);
and U12539 (N_12539,N_11340,N_11648);
nand U12540 (N_12540,N_11906,N_11005);
and U12541 (N_12541,N_11015,N_10822);
nor U12542 (N_12542,N_11212,N_10744);
nor U12543 (N_12543,N_10927,N_10526);
nand U12544 (N_12544,N_10616,N_10784);
nor U12545 (N_12545,N_11265,N_11496);
nor U12546 (N_12546,N_11706,N_11376);
nand U12547 (N_12547,N_11735,N_11463);
or U12548 (N_12548,N_11277,N_10735);
and U12549 (N_12549,N_10599,N_11165);
nor U12550 (N_12550,N_11173,N_11193);
and U12551 (N_12551,N_11927,N_11529);
nand U12552 (N_12552,N_11246,N_11236);
and U12553 (N_12553,N_11342,N_11351);
nor U12554 (N_12554,N_11527,N_11756);
and U12555 (N_12555,N_11305,N_11757);
nor U12556 (N_12556,N_11117,N_11199);
and U12557 (N_12557,N_11072,N_10544);
and U12558 (N_12558,N_11897,N_11311);
nor U12559 (N_12559,N_10931,N_11803);
or U12560 (N_12560,N_10577,N_10861);
or U12561 (N_12561,N_10997,N_10816);
nand U12562 (N_12562,N_11884,N_11245);
nand U12563 (N_12563,N_11625,N_10570);
nor U12564 (N_12564,N_10652,N_10537);
nand U12565 (N_12565,N_10731,N_11624);
nand U12566 (N_12566,N_11278,N_11362);
and U12567 (N_12567,N_10647,N_11792);
nand U12568 (N_12568,N_11601,N_11178);
and U12569 (N_12569,N_11167,N_11921);
and U12570 (N_12570,N_11032,N_11828);
or U12571 (N_12571,N_11318,N_11992);
nor U12572 (N_12572,N_11213,N_11076);
nand U12573 (N_12573,N_11477,N_11561);
or U12574 (N_12574,N_11862,N_11939);
nand U12575 (N_12575,N_11290,N_10613);
nand U12576 (N_12576,N_10749,N_11553);
nor U12577 (N_12577,N_11095,N_11776);
and U12578 (N_12578,N_11387,N_11303);
nor U12579 (N_12579,N_10777,N_11411);
nor U12580 (N_12580,N_11747,N_11347);
nor U12581 (N_12581,N_11937,N_11247);
nor U12582 (N_12582,N_11592,N_11211);
nand U12583 (N_12583,N_11588,N_10872);
or U12584 (N_12584,N_11220,N_11557);
and U12585 (N_12585,N_11764,N_11514);
or U12586 (N_12586,N_11777,N_11450);
and U12587 (N_12587,N_10865,N_11439);
nand U12588 (N_12588,N_10830,N_10960);
nand U12589 (N_12589,N_10849,N_11594);
or U12590 (N_12590,N_11708,N_10983);
and U12591 (N_12591,N_11830,N_10716);
and U12592 (N_12592,N_10543,N_11503);
and U12593 (N_12593,N_11836,N_11158);
or U12594 (N_12594,N_10940,N_11885);
or U12595 (N_12595,N_11969,N_11520);
or U12596 (N_12596,N_10517,N_10987);
or U12597 (N_12597,N_11612,N_11616);
nor U12598 (N_12598,N_11815,N_11605);
or U12599 (N_12599,N_11126,N_10564);
and U12600 (N_12600,N_11320,N_10889);
nor U12601 (N_12601,N_11284,N_11996);
nand U12602 (N_12602,N_10608,N_10941);
nor U12603 (N_12603,N_10738,N_10856);
and U12604 (N_12604,N_11202,N_10916);
and U12605 (N_12605,N_10937,N_11659);
and U12606 (N_12606,N_11810,N_10638);
nand U12607 (N_12607,N_11933,N_11237);
or U12608 (N_12608,N_11432,N_11722);
or U12609 (N_12609,N_10681,N_10508);
or U12610 (N_12610,N_11122,N_10694);
nor U12611 (N_12611,N_11262,N_11829);
nand U12612 (N_12612,N_11790,N_11134);
nand U12613 (N_12613,N_10912,N_10748);
or U12614 (N_12614,N_11732,N_11745);
or U12615 (N_12615,N_11443,N_11788);
nand U12616 (N_12616,N_11881,N_11655);
nor U12617 (N_12617,N_11157,N_11123);
or U12618 (N_12618,N_10893,N_11137);
nor U12619 (N_12619,N_11819,N_10627);
or U12620 (N_12620,N_11738,N_10851);
and U12621 (N_12621,N_11198,N_11883);
nor U12622 (N_12622,N_10875,N_11154);
nor U12623 (N_12623,N_11770,N_11071);
nor U12624 (N_12624,N_11386,N_11272);
nand U12625 (N_12625,N_11963,N_11749);
or U12626 (N_12626,N_11427,N_11316);
or U12627 (N_12627,N_11469,N_10597);
nor U12628 (N_12628,N_11131,N_11419);
and U12629 (N_12629,N_11023,N_11257);
nand U12630 (N_12630,N_10598,N_11723);
or U12631 (N_12631,N_11285,N_11108);
or U12632 (N_12632,N_11678,N_11229);
and U12633 (N_12633,N_11727,N_11962);
nand U12634 (N_12634,N_10585,N_11691);
or U12635 (N_12635,N_10886,N_11890);
nand U12636 (N_12636,N_11197,N_10561);
nor U12637 (N_12637,N_11917,N_11608);
and U12638 (N_12638,N_11243,N_10520);
and U12639 (N_12639,N_11354,N_10615);
nand U12640 (N_12640,N_10674,N_10709);
and U12641 (N_12641,N_11984,N_11661);
or U12642 (N_12642,N_11785,N_10935);
and U12643 (N_12643,N_11353,N_10788);
nand U12644 (N_12644,N_11812,N_10898);
nand U12645 (N_12645,N_11365,N_10765);
nor U12646 (N_12646,N_11446,N_11856);
nor U12647 (N_12647,N_11614,N_11928);
nand U12648 (N_12648,N_10939,N_10883);
nor U12649 (N_12649,N_10787,N_11965);
or U12650 (N_12650,N_11725,N_11479);
nand U12651 (N_12651,N_11901,N_11522);
or U12652 (N_12652,N_11218,N_11068);
nand U12653 (N_12653,N_11652,N_11894);
nor U12654 (N_12654,N_11222,N_11418);
nor U12655 (N_12655,N_11409,N_11044);
nand U12656 (N_12656,N_10810,N_10885);
nand U12657 (N_12657,N_11380,N_11148);
nor U12658 (N_12658,N_10811,N_11453);
or U12659 (N_12659,N_11304,N_10791);
nand U12660 (N_12660,N_11267,N_11105);
and U12661 (N_12661,N_11341,N_11478);
or U12662 (N_12662,N_10848,N_10702);
nor U12663 (N_12663,N_11090,N_11623);
or U12664 (N_12664,N_11506,N_11806);
and U12665 (N_12665,N_11709,N_11669);
or U12666 (N_12666,N_11254,N_11758);
or U12667 (N_12667,N_11585,N_11838);
and U12668 (N_12668,N_11801,N_11537);
nor U12669 (N_12669,N_10842,N_10958);
nor U12670 (N_12670,N_11544,N_10612);
nand U12671 (N_12671,N_11034,N_11161);
nand U12672 (N_12672,N_10982,N_11390);
and U12673 (N_12673,N_11151,N_10513);
nand U12674 (N_12674,N_11441,N_10888);
xor U12675 (N_12675,N_11494,N_10897);
and U12676 (N_12676,N_11687,N_11831);
or U12677 (N_12677,N_11086,N_11979);
and U12678 (N_12678,N_11268,N_11964);
nand U12679 (N_12679,N_11018,N_11983);
or U12680 (N_12680,N_10687,N_11406);
or U12681 (N_12681,N_10904,N_10915);
or U12682 (N_12682,N_11814,N_10746);
and U12683 (N_12683,N_10726,N_11361);
nor U12684 (N_12684,N_11989,N_10713);
nor U12685 (N_12685,N_11632,N_11251);
nand U12686 (N_12686,N_11955,N_11710);
nor U12687 (N_12687,N_11269,N_11816);
or U12688 (N_12688,N_10659,N_10828);
nor U12689 (N_12689,N_10635,N_11558);
and U12690 (N_12690,N_11936,N_11407);
nand U12691 (N_12691,N_10614,N_11217);
or U12692 (N_12692,N_11547,N_11736);
and U12693 (N_12693,N_10804,N_10827);
or U12694 (N_12694,N_11621,N_10867);
and U12695 (N_12695,N_11033,N_11383);
nand U12696 (N_12696,N_11098,N_10587);
or U12697 (N_12697,N_11874,N_11824);
nor U12698 (N_12698,N_10641,N_11052);
and U12699 (N_12699,N_11990,N_11889);
or U12700 (N_12700,N_11576,N_11475);
and U12701 (N_12701,N_11609,N_11946);
and U12702 (N_12702,N_10568,N_10629);
nand U12703 (N_12703,N_11968,N_11125);
nor U12704 (N_12704,N_11244,N_10969);
nand U12705 (N_12705,N_11062,N_10771);
and U12706 (N_12706,N_11408,N_10611);
or U12707 (N_12707,N_11010,N_11798);
or U12708 (N_12708,N_10965,N_11541);
and U12709 (N_12709,N_11846,N_10676);
or U12710 (N_12710,N_11099,N_11991);
and U12711 (N_12711,N_10891,N_10624);
or U12712 (N_12712,N_10933,N_11966);
and U12713 (N_12713,N_11662,N_11771);
nor U12714 (N_12714,N_11973,N_10799);
and U12715 (N_12715,N_11492,N_11596);
and U12716 (N_12716,N_10909,N_11606);
nor U12717 (N_12717,N_11321,N_11207);
or U12718 (N_12718,N_11734,N_11618);
or U12719 (N_12719,N_10910,N_11187);
or U12720 (N_12720,N_10572,N_11942);
nor U12721 (N_12721,N_11877,N_10734);
or U12722 (N_12722,N_11060,N_10686);
and U12723 (N_12723,N_10541,N_11930);
nor U12724 (N_12724,N_11423,N_11271);
xnor U12725 (N_12725,N_10890,N_11932);
or U12726 (N_12726,N_10993,N_10666);
or U12727 (N_12727,N_11848,N_11572);
nand U12728 (N_12728,N_10800,N_10617);
and U12729 (N_12729,N_11248,N_11700);
and U12730 (N_12730,N_11223,N_11464);
and U12731 (N_12731,N_11663,N_11665);
nor U12732 (N_12732,N_11204,N_11554);
nor U12733 (N_12733,N_10690,N_11526);
nand U12734 (N_12734,N_11348,N_11309);
and U12735 (N_12735,N_11358,N_11581);
and U12736 (N_12736,N_11707,N_10730);
or U12737 (N_12737,N_10995,N_11371);
and U12738 (N_12738,N_10809,N_11287);
and U12739 (N_12739,N_11399,N_10839);
nand U12740 (N_12740,N_11115,N_11565);
nand U12741 (N_12741,N_11058,N_11214);
nand U12742 (N_12742,N_10529,N_11036);
or U12743 (N_12743,N_11656,N_10584);
and U12744 (N_12744,N_11666,N_11768);
or U12745 (N_12745,N_10998,N_11880);
and U12746 (N_12746,N_11982,N_11066);
or U12747 (N_12747,N_11037,N_11694);
xor U12748 (N_12748,N_11486,N_11317);
and U12749 (N_12749,N_10519,N_11683);
nor U12750 (N_12750,N_11578,N_11468);
nand U12751 (N_12751,N_11145,N_11863);
or U12752 (N_12752,N_11464,N_11253);
nor U12753 (N_12753,N_11304,N_11554);
and U12754 (N_12754,N_11619,N_10640);
nor U12755 (N_12755,N_10727,N_11649);
or U12756 (N_12756,N_11496,N_10718);
and U12757 (N_12757,N_10766,N_11555);
or U12758 (N_12758,N_11305,N_11872);
nor U12759 (N_12759,N_11869,N_11310);
nand U12760 (N_12760,N_11081,N_11240);
and U12761 (N_12761,N_10733,N_10522);
and U12762 (N_12762,N_10741,N_10832);
nor U12763 (N_12763,N_10500,N_11189);
nand U12764 (N_12764,N_10921,N_10937);
and U12765 (N_12765,N_11026,N_11581);
nand U12766 (N_12766,N_11816,N_11657);
nand U12767 (N_12767,N_11024,N_11184);
and U12768 (N_12768,N_11809,N_11038);
nor U12769 (N_12769,N_11768,N_11432);
and U12770 (N_12770,N_11465,N_10824);
and U12771 (N_12771,N_10658,N_11240);
nor U12772 (N_12772,N_10547,N_11110);
or U12773 (N_12773,N_11560,N_11200);
or U12774 (N_12774,N_10825,N_11981);
xnor U12775 (N_12775,N_11171,N_10922);
nand U12776 (N_12776,N_10842,N_11439);
and U12777 (N_12777,N_10822,N_11538);
nor U12778 (N_12778,N_10527,N_11186);
nand U12779 (N_12779,N_11692,N_11327);
and U12780 (N_12780,N_11782,N_11159);
or U12781 (N_12781,N_10949,N_10501);
and U12782 (N_12782,N_11599,N_11127);
or U12783 (N_12783,N_11403,N_11299);
and U12784 (N_12784,N_11867,N_10698);
or U12785 (N_12785,N_10875,N_11102);
nor U12786 (N_12786,N_11579,N_11850);
nor U12787 (N_12787,N_11309,N_10532);
nor U12788 (N_12788,N_10843,N_10637);
and U12789 (N_12789,N_11949,N_10783);
nor U12790 (N_12790,N_10628,N_11040);
or U12791 (N_12791,N_11474,N_11658);
and U12792 (N_12792,N_10983,N_11781);
nor U12793 (N_12793,N_11573,N_11434);
or U12794 (N_12794,N_10500,N_11672);
and U12795 (N_12795,N_11271,N_11128);
nor U12796 (N_12796,N_11750,N_11727);
and U12797 (N_12797,N_10630,N_10510);
xor U12798 (N_12798,N_11214,N_11930);
nand U12799 (N_12799,N_11976,N_10688);
nand U12800 (N_12800,N_11890,N_11588);
or U12801 (N_12801,N_11675,N_11270);
and U12802 (N_12802,N_11147,N_11058);
and U12803 (N_12803,N_11474,N_11500);
nor U12804 (N_12804,N_11954,N_10501);
nand U12805 (N_12805,N_11456,N_11011);
and U12806 (N_12806,N_11548,N_10581);
and U12807 (N_12807,N_10877,N_10943);
or U12808 (N_12808,N_11990,N_10643);
and U12809 (N_12809,N_10522,N_11662);
nor U12810 (N_12810,N_10521,N_11316);
nor U12811 (N_12811,N_10842,N_11154);
or U12812 (N_12812,N_11907,N_11788);
and U12813 (N_12813,N_10572,N_10540);
or U12814 (N_12814,N_11676,N_11096);
or U12815 (N_12815,N_11974,N_10513);
or U12816 (N_12816,N_11863,N_10736);
nor U12817 (N_12817,N_11588,N_11202);
and U12818 (N_12818,N_10670,N_10975);
nor U12819 (N_12819,N_11555,N_11585);
nand U12820 (N_12820,N_10771,N_11459);
or U12821 (N_12821,N_11905,N_11719);
nand U12822 (N_12822,N_11845,N_10943);
nand U12823 (N_12823,N_11287,N_11185);
or U12824 (N_12824,N_10608,N_11906);
nor U12825 (N_12825,N_10558,N_11606);
and U12826 (N_12826,N_11292,N_11971);
nor U12827 (N_12827,N_10505,N_10891);
nand U12828 (N_12828,N_11115,N_10869);
and U12829 (N_12829,N_11162,N_11560);
or U12830 (N_12830,N_11727,N_10870);
or U12831 (N_12831,N_11701,N_11344);
or U12832 (N_12832,N_10842,N_11836);
nand U12833 (N_12833,N_11768,N_10614);
or U12834 (N_12834,N_11301,N_11112);
or U12835 (N_12835,N_11218,N_11376);
nor U12836 (N_12836,N_11721,N_11931);
or U12837 (N_12837,N_11328,N_11838);
nand U12838 (N_12838,N_10864,N_10575);
nand U12839 (N_12839,N_11781,N_10580);
or U12840 (N_12840,N_11824,N_11074);
nor U12841 (N_12841,N_11448,N_11435);
and U12842 (N_12842,N_10507,N_10561);
nor U12843 (N_12843,N_10918,N_10521);
or U12844 (N_12844,N_10630,N_11266);
or U12845 (N_12845,N_11108,N_10994);
and U12846 (N_12846,N_11233,N_11331);
nand U12847 (N_12847,N_10835,N_10504);
nor U12848 (N_12848,N_11669,N_10631);
nor U12849 (N_12849,N_10592,N_11680);
or U12850 (N_12850,N_11671,N_11118);
or U12851 (N_12851,N_11021,N_11734);
or U12852 (N_12852,N_10894,N_11100);
and U12853 (N_12853,N_11312,N_10675);
and U12854 (N_12854,N_11899,N_11695);
nor U12855 (N_12855,N_10531,N_10768);
nor U12856 (N_12856,N_11733,N_10811);
or U12857 (N_12857,N_11535,N_11611);
nor U12858 (N_12858,N_11137,N_10792);
nand U12859 (N_12859,N_10515,N_10942);
nor U12860 (N_12860,N_10687,N_11086);
and U12861 (N_12861,N_11277,N_10513);
nand U12862 (N_12862,N_10957,N_10925);
nor U12863 (N_12863,N_11290,N_11966);
nor U12864 (N_12864,N_11504,N_11224);
or U12865 (N_12865,N_11123,N_11382);
and U12866 (N_12866,N_11836,N_10779);
or U12867 (N_12867,N_10596,N_11817);
or U12868 (N_12868,N_11897,N_10702);
nand U12869 (N_12869,N_11054,N_11855);
nand U12870 (N_12870,N_10506,N_10799);
or U12871 (N_12871,N_10790,N_11042);
nor U12872 (N_12872,N_11816,N_11591);
nand U12873 (N_12873,N_11248,N_11163);
nand U12874 (N_12874,N_11666,N_10857);
or U12875 (N_12875,N_11574,N_11957);
and U12876 (N_12876,N_11828,N_11559);
nor U12877 (N_12877,N_11605,N_10693);
or U12878 (N_12878,N_11150,N_11580);
nand U12879 (N_12879,N_11361,N_10599);
nor U12880 (N_12880,N_11631,N_10555);
nand U12881 (N_12881,N_11632,N_11719);
and U12882 (N_12882,N_11652,N_11432);
or U12883 (N_12883,N_11814,N_10859);
and U12884 (N_12884,N_11208,N_10629);
nand U12885 (N_12885,N_11977,N_10742);
nand U12886 (N_12886,N_11576,N_11323);
nor U12887 (N_12887,N_10607,N_10573);
nor U12888 (N_12888,N_10708,N_11514);
and U12889 (N_12889,N_10608,N_11260);
nand U12890 (N_12890,N_10942,N_11578);
and U12891 (N_12891,N_10770,N_10756);
or U12892 (N_12892,N_11872,N_10725);
nor U12893 (N_12893,N_11716,N_11906);
or U12894 (N_12894,N_10720,N_11946);
or U12895 (N_12895,N_11252,N_11342);
and U12896 (N_12896,N_11901,N_10587);
or U12897 (N_12897,N_11413,N_11121);
nor U12898 (N_12898,N_11091,N_10829);
and U12899 (N_12899,N_10912,N_11796);
xor U12900 (N_12900,N_10559,N_11434);
or U12901 (N_12901,N_11653,N_11694);
nor U12902 (N_12902,N_11386,N_11889);
nand U12903 (N_12903,N_11258,N_11097);
nand U12904 (N_12904,N_11770,N_11540);
nor U12905 (N_12905,N_10837,N_11250);
or U12906 (N_12906,N_11866,N_11676);
or U12907 (N_12907,N_11324,N_11725);
nor U12908 (N_12908,N_11119,N_11470);
or U12909 (N_12909,N_11900,N_11525);
nor U12910 (N_12910,N_10864,N_10970);
nor U12911 (N_12911,N_11023,N_11910);
and U12912 (N_12912,N_10948,N_11746);
or U12913 (N_12913,N_10812,N_11067);
or U12914 (N_12914,N_10557,N_10722);
nor U12915 (N_12915,N_10657,N_11126);
nand U12916 (N_12916,N_10783,N_10564);
nor U12917 (N_12917,N_10954,N_11552);
nand U12918 (N_12918,N_10906,N_10545);
nor U12919 (N_12919,N_11620,N_11971);
or U12920 (N_12920,N_11665,N_11687);
and U12921 (N_12921,N_10995,N_11972);
and U12922 (N_12922,N_10570,N_11943);
nand U12923 (N_12923,N_11769,N_10793);
and U12924 (N_12924,N_11195,N_10526);
nor U12925 (N_12925,N_11461,N_11455);
nand U12926 (N_12926,N_10561,N_11676);
nand U12927 (N_12927,N_11646,N_11498);
nand U12928 (N_12928,N_11413,N_11537);
nand U12929 (N_12929,N_11214,N_11743);
or U12930 (N_12930,N_11213,N_11350);
xnor U12931 (N_12931,N_11232,N_11719);
and U12932 (N_12932,N_11604,N_10545);
nor U12933 (N_12933,N_11957,N_11830);
and U12934 (N_12934,N_11685,N_11582);
or U12935 (N_12935,N_11381,N_11750);
or U12936 (N_12936,N_11664,N_10929);
nor U12937 (N_12937,N_10827,N_11662);
or U12938 (N_12938,N_11224,N_11720);
nand U12939 (N_12939,N_11733,N_11210);
nand U12940 (N_12940,N_11587,N_11515);
nor U12941 (N_12941,N_11901,N_11482);
and U12942 (N_12942,N_11820,N_11810);
or U12943 (N_12943,N_11766,N_10743);
and U12944 (N_12944,N_11698,N_10649);
or U12945 (N_12945,N_11281,N_11792);
and U12946 (N_12946,N_11776,N_10574);
nor U12947 (N_12947,N_11213,N_10671);
or U12948 (N_12948,N_11588,N_10957);
and U12949 (N_12949,N_11756,N_11741);
and U12950 (N_12950,N_11937,N_11232);
nor U12951 (N_12951,N_11782,N_11373);
or U12952 (N_12952,N_11148,N_11643);
nor U12953 (N_12953,N_10696,N_11917);
nor U12954 (N_12954,N_11081,N_10505);
or U12955 (N_12955,N_10610,N_10700);
and U12956 (N_12956,N_10743,N_11085);
and U12957 (N_12957,N_10722,N_10507);
nor U12958 (N_12958,N_10980,N_11228);
nand U12959 (N_12959,N_10702,N_11250);
nor U12960 (N_12960,N_11127,N_11204);
xnor U12961 (N_12961,N_11789,N_11108);
or U12962 (N_12962,N_11875,N_10519);
nand U12963 (N_12963,N_11553,N_10745);
nor U12964 (N_12964,N_11030,N_11108);
nor U12965 (N_12965,N_11785,N_11800);
nor U12966 (N_12966,N_11996,N_11900);
or U12967 (N_12967,N_10597,N_10941);
or U12968 (N_12968,N_11772,N_11773);
nand U12969 (N_12969,N_10745,N_11975);
nor U12970 (N_12970,N_10929,N_11831);
and U12971 (N_12971,N_11263,N_11339);
nor U12972 (N_12972,N_11414,N_11376);
nor U12973 (N_12973,N_11882,N_10987);
nor U12974 (N_12974,N_10840,N_10778);
nor U12975 (N_12975,N_11810,N_11297);
or U12976 (N_12976,N_11715,N_10595);
or U12977 (N_12977,N_10531,N_11788);
nand U12978 (N_12978,N_10930,N_10615);
and U12979 (N_12979,N_11523,N_11247);
or U12980 (N_12980,N_11834,N_11525);
and U12981 (N_12981,N_11763,N_11272);
and U12982 (N_12982,N_11386,N_10830);
and U12983 (N_12983,N_11482,N_11568);
nand U12984 (N_12984,N_11643,N_10904);
or U12985 (N_12985,N_10810,N_10851);
or U12986 (N_12986,N_11461,N_11218);
nand U12987 (N_12987,N_10952,N_11578);
nand U12988 (N_12988,N_11131,N_11610);
nand U12989 (N_12989,N_10841,N_10979);
nor U12990 (N_12990,N_11922,N_11978);
nand U12991 (N_12991,N_10545,N_11425);
nand U12992 (N_12992,N_10631,N_10536);
nor U12993 (N_12993,N_11416,N_10603);
and U12994 (N_12994,N_11794,N_10686);
nor U12995 (N_12995,N_11401,N_11700);
and U12996 (N_12996,N_11722,N_11294);
nand U12997 (N_12997,N_11046,N_10504);
and U12998 (N_12998,N_11948,N_11660);
and U12999 (N_12999,N_11438,N_10938);
and U13000 (N_13000,N_11426,N_10574);
or U13001 (N_13001,N_11435,N_11455);
nand U13002 (N_13002,N_11079,N_11603);
nor U13003 (N_13003,N_10866,N_11846);
or U13004 (N_13004,N_11144,N_11444);
nand U13005 (N_13005,N_11496,N_10872);
nor U13006 (N_13006,N_11408,N_10903);
or U13007 (N_13007,N_10508,N_11789);
or U13008 (N_13008,N_11488,N_11043);
xnor U13009 (N_13009,N_11772,N_11408);
and U13010 (N_13010,N_11205,N_11474);
or U13011 (N_13011,N_11940,N_11128);
nand U13012 (N_13012,N_10779,N_11042);
nand U13013 (N_13013,N_11580,N_11505);
nor U13014 (N_13014,N_11437,N_11869);
and U13015 (N_13015,N_10519,N_10928);
nor U13016 (N_13016,N_10986,N_10670);
nand U13017 (N_13017,N_11657,N_11827);
nand U13018 (N_13018,N_10651,N_11099);
nand U13019 (N_13019,N_11409,N_11492);
and U13020 (N_13020,N_11358,N_11065);
nor U13021 (N_13021,N_11084,N_11709);
nor U13022 (N_13022,N_11164,N_10736);
or U13023 (N_13023,N_10640,N_11745);
and U13024 (N_13024,N_11711,N_10527);
or U13025 (N_13025,N_11421,N_11216);
nor U13026 (N_13026,N_11492,N_10910);
and U13027 (N_13027,N_11114,N_11616);
and U13028 (N_13028,N_11053,N_11361);
or U13029 (N_13029,N_11219,N_10908);
nor U13030 (N_13030,N_10818,N_11682);
nand U13031 (N_13031,N_11405,N_10850);
or U13032 (N_13032,N_10579,N_11499);
or U13033 (N_13033,N_10716,N_10860);
or U13034 (N_13034,N_11435,N_11697);
and U13035 (N_13035,N_11988,N_10865);
and U13036 (N_13036,N_10573,N_11839);
nand U13037 (N_13037,N_11317,N_11195);
nand U13038 (N_13038,N_11448,N_11582);
nand U13039 (N_13039,N_11107,N_10922);
and U13040 (N_13040,N_11186,N_11443);
nor U13041 (N_13041,N_11303,N_11260);
nor U13042 (N_13042,N_10696,N_10842);
and U13043 (N_13043,N_11606,N_11734);
nor U13044 (N_13044,N_10755,N_10506);
nor U13045 (N_13045,N_10861,N_11470);
nand U13046 (N_13046,N_11172,N_11892);
and U13047 (N_13047,N_10884,N_10984);
nand U13048 (N_13048,N_10700,N_10683);
nor U13049 (N_13049,N_11038,N_10737);
nor U13050 (N_13050,N_10578,N_11450);
nor U13051 (N_13051,N_11477,N_11122);
nor U13052 (N_13052,N_10706,N_11696);
nand U13053 (N_13053,N_11428,N_11034);
nor U13054 (N_13054,N_10759,N_11983);
xnor U13055 (N_13055,N_11909,N_11657);
or U13056 (N_13056,N_11149,N_11638);
or U13057 (N_13057,N_11131,N_11893);
or U13058 (N_13058,N_11573,N_10758);
nand U13059 (N_13059,N_11767,N_11758);
xor U13060 (N_13060,N_11778,N_10592);
and U13061 (N_13061,N_11705,N_11577);
or U13062 (N_13062,N_11624,N_10836);
nor U13063 (N_13063,N_11471,N_11484);
and U13064 (N_13064,N_10869,N_11555);
or U13065 (N_13065,N_11005,N_11982);
xnor U13066 (N_13066,N_10971,N_11664);
nor U13067 (N_13067,N_10579,N_10678);
nand U13068 (N_13068,N_10540,N_11763);
and U13069 (N_13069,N_11117,N_11106);
or U13070 (N_13070,N_10852,N_11323);
nor U13071 (N_13071,N_11482,N_11164);
nor U13072 (N_13072,N_10653,N_11588);
and U13073 (N_13073,N_10671,N_11166);
and U13074 (N_13074,N_11733,N_11766);
nand U13075 (N_13075,N_11628,N_11080);
nor U13076 (N_13076,N_11543,N_11333);
nand U13077 (N_13077,N_11065,N_11567);
or U13078 (N_13078,N_11805,N_10781);
nand U13079 (N_13079,N_10942,N_11237);
nor U13080 (N_13080,N_11875,N_10709);
nor U13081 (N_13081,N_10910,N_11882);
and U13082 (N_13082,N_11303,N_10783);
or U13083 (N_13083,N_11392,N_10695);
nor U13084 (N_13084,N_11620,N_11036);
nand U13085 (N_13085,N_11759,N_10625);
nand U13086 (N_13086,N_11772,N_11495);
and U13087 (N_13087,N_11495,N_11892);
nor U13088 (N_13088,N_11803,N_11774);
or U13089 (N_13089,N_10762,N_11844);
and U13090 (N_13090,N_10585,N_10822);
or U13091 (N_13091,N_11286,N_10504);
nor U13092 (N_13092,N_11451,N_11176);
or U13093 (N_13093,N_10776,N_10638);
or U13094 (N_13094,N_11591,N_11289);
or U13095 (N_13095,N_10990,N_10577);
nand U13096 (N_13096,N_11704,N_11110);
nand U13097 (N_13097,N_11564,N_10854);
and U13098 (N_13098,N_11334,N_10762);
and U13099 (N_13099,N_11225,N_11192);
nor U13100 (N_13100,N_10569,N_10697);
xnor U13101 (N_13101,N_11356,N_11451);
and U13102 (N_13102,N_10755,N_11325);
nor U13103 (N_13103,N_11818,N_10949);
or U13104 (N_13104,N_11714,N_11777);
xor U13105 (N_13105,N_10616,N_11041);
and U13106 (N_13106,N_11338,N_11231);
and U13107 (N_13107,N_10721,N_11431);
nor U13108 (N_13108,N_11691,N_10807);
nand U13109 (N_13109,N_10514,N_10589);
nand U13110 (N_13110,N_10738,N_10879);
nor U13111 (N_13111,N_10611,N_11768);
or U13112 (N_13112,N_11948,N_11253);
or U13113 (N_13113,N_11197,N_11267);
nor U13114 (N_13114,N_10910,N_11655);
nand U13115 (N_13115,N_10532,N_10977);
nor U13116 (N_13116,N_11233,N_11853);
or U13117 (N_13117,N_10510,N_11104);
or U13118 (N_13118,N_10800,N_10831);
and U13119 (N_13119,N_11243,N_10687);
nor U13120 (N_13120,N_10646,N_11007);
or U13121 (N_13121,N_11030,N_11982);
xor U13122 (N_13122,N_10663,N_10503);
xnor U13123 (N_13123,N_11332,N_11898);
nor U13124 (N_13124,N_11057,N_11416);
or U13125 (N_13125,N_11962,N_11557);
nand U13126 (N_13126,N_11604,N_10848);
nor U13127 (N_13127,N_10622,N_11051);
nand U13128 (N_13128,N_11416,N_11544);
or U13129 (N_13129,N_11656,N_11622);
or U13130 (N_13130,N_11867,N_11241);
nand U13131 (N_13131,N_11907,N_11359);
or U13132 (N_13132,N_11877,N_11129);
nand U13133 (N_13133,N_10871,N_11242);
nand U13134 (N_13134,N_11154,N_10960);
nor U13135 (N_13135,N_10647,N_11954);
nor U13136 (N_13136,N_11374,N_10563);
nand U13137 (N_13137,N_10617,N_10681);
or U13138 (N_13138,N_11217,N_11540);
nand U13139 (N_13139,N_11325,N_10556);
nor U13140 (N_13140,N_11030,N_11344);
and U13141 (N_13141,N_11231,N_10764);
nor U13142 (N_13142,N_11125,N_10849);
and U13143 (N_13143,N_11266,N_11673);
or U13144 (N_13144,N_10615,N_11840);
nand U13145 (N_13145,N_10638,N_10708);
nand U13146 (N_13146,N_11193,N_10690);
nand U13147 (N_13147,N_11551,N_11146);
or U13148 (N_13148,N_11832,N_11097);
or U13149 (N_13149,N_11477,N_11342);
and U13150 (N_13150,N_11300,N_10806);
nor U13151 (N_13151,N_11246,N_11418);
nand U13152 (N_13152,N_11669,N_10783);
nor U13153 (N_13153,N_10667,N_11327);
or U13154 (N_13154,N_11290,N_11007);
nand U13155 (N_13155,N_11077,N_11409);
nor U13156 (N_13156,N_11610,N_11273);
nor U13157 (N_13157,N_11882,N_10963);
nand U13158 (N_13158,N_10764,N_10740);
xor U13159 (N_13159,N_11893,N_11861);
or U13160 (N_13160,N_11983,N_11198);
and U13161 (N_13161,N_10858,N_11729);
and U13162 (N_13162,N_11207,N_11403);
or U13163 (N_13163,N_11883,N_11828);
nand U13164 (N_13164,N_11273,N_11354);
nor U13165 (N_13165,N_11216,N_11611);
or U13166 (N_13166,N_11487,N_11463);
or U13167 (N_13167,N_11050,N_11994);
or U13168 (N_13168,N_11690,N_10593);
and U13169 (N_13169,N_11988,N_11461);
or U13170 (N_13170,N_10622,N_10506);
or U13171 (N_13171,N_10529,N_11161);
nand U13172 (N_13172,N_11899,N_11400);
nor U13173 (N_13173,N_11242,N_11235);
xor U13174 (N_13174,N_10826,N_11895);
and U13175 (N_13175,N_11713,N_10891);
or U13176 (N_13176,N_11188,N_11688);
nor U13177 (N_13177,N_11982,N_11621);
and U13178 (N_13178,N_11229,N_11395);
nor U13179 (N_13179,N_10740,N_11148);
and U13180 (N_13180,N_10993,N_10603);
nand U13181 (N_13181,N_11506,N_10545);
nand U13182 (N_13182,N_11396,N_10880);
nor U13183 (N_13183,N_11239,N_11757);
and U13184 (N_13184,N_10910,N_10997);
and U13185 (N_13185,N_11572,N_10995);
nand U13186 (N_13186,N_11725,N_11883);
and U13187 (N_13187,N_11345,N_10567);
and U13188 (N_13188,N_10761,N_11333);
nand U13189 (N_13189,N_11600,N_11055);
or U13190 (N_13190,N_11511,N_11918);
nand U13191 (N_13191,N_11752,N_10837);
or U13192 (N_13192,N_10601,N_10855);
nand U13193 (N_13193,N_11839,N_11696);
or U13194 (N_13194,N_11073,N_10923);
or U13195 (N_13195,N_10504,N_10684);
or U13196 (N_13196,N_11835,N_11230);
nand U13197 (N_13197,N_11968,N_11819);
or U13198 (N_13198,N_11457,N_11079);
nor U13199 (N_13199,N_11102,N_10822);
nand U13200 (N_13200,N_11391,N_11416);
nand U13201 (N_13201,N_10683,N_11936);
or U13202 (N_13202,N_11668,N_11899);
or U13203 (N_13203,N_10554,N_11578);
nor U13204 (N_13204,N_11941,N_11535);
nand U13205 (N_13205,N_10543,N_10531);
and U13206 (N_13206,N_10728,N_11897);
nand U13207 (N_13207,N_11249,N_11092);
xnor U13208 (N_13208,N_11540,N_11533);
nand U13209 (N_13209,N_11277,N_10727);
nand U13210 (N_13210,N_11935,N_10936);
nor U13211 (N_13211,N_11083,N_11721);
or U13212 (N_13212,N_10671,N_10598);
and U13213 (N_13213,N_11486,N_10509);
nor U13214 (N_13214,N_11526,N_11325);
and U13215 (N_13215,N_11736,N_10631);
or U13216 (N_13216,N_11824,N_10926);
and U13217 (N_13217,N_10650,N_11585);
and U13218 (N_13218,N_10532,N_11317);
and U13219 (N_13219,N_10710,N_10624);
nand U13220 (N_13220,N_11243,N_11016);
nor U13221 (N_13221,N_11757,N_11032);
nand U13222 (N_13222,N_11895,N_11601);
and U13223 (N_13223,N_11242,N_11128);
nor U13224 (N_13224,N_11440,N_11624);
nor U13225 (N_13225,N_11906,N_11077);
or U13226 (N_13226,N_11400,N_11983);
and U13227 (N_13227,N_10865,N_10599);
or U13228 (N_13228,N_10816,N_11807);
or U13229 (N_13229,N_10547,N_11934);
nor U13230 (N_13230,N_11908,N_11646);
and U13231 (N_13231,N_10972,N_10662);
and U13232 (N_13232,N_11030,N_11954);
or U13233 (N_13233,N_11476,N_10508);
and U13234 (N_13234,N_11053,N_11267);
nand U13235 (N_13235,N_11345,N_10671);
or U13236 (N_13236,N_11385,N_10851);
or U13237 (N_13237,N_10748,N_11069);
nand U13238 (N_13238,N_11224,N_11229);
and U13239 (N_13239,N_10871,N_11039);
nand U13240 (N_13240,N_10694,N_11225);
nand U13241 (N_13241,N_11726,N_11102);
nor U13242 (N_13242,N_10619,N_11049);
or U13243 (N_13243,N_10817,N_11278);
nor U13244 (N_13244,N_11001,N_10857);
nand U13245 (N_13245,N_11150,N_10897);
or U13246 (N_13246,N_11212,N_11213);
or U13247 (N_13247,N_10551,N_11488);
and U13248 (N_13248,N_10776,N_11483);
and U13249 (N_13249,N_11466,N_10681);
nand U13250 (N_13250,N_10541,N_11981);
and U13251 (N_13251,N_11796,N_11090);
nor U13252 (N_13252,N_11240,N_10839);
and U13253 (N_13253,N_10893,N_11720);
nor U13254 (N_13254,N_10874,N_10941);
and U13255 (N_13255,N_11286,N_10882);
nor U13256 (N_13256,N_10810,N_11537);
nor U13257 (N_13257,N_10652,N_10657);
nand U13258 (N_13258,N_11334,N_10602);
nor U13259 (N_13259,N_11384,N_11632);
or U13260 (N_13260,N_10906,N_11280);
or U13261 (N_13261,N_11940,N_10743);
and U13262 (N_13262,N_11639,N_11369);
and U13263 (N_13263,N_11021,N_11314);
nand U13264 (N_13264,N_10709,N_11194);
and U13265 (N_13265,N_10933,N_11321);
nand U13266 (N_13266,N_11531,N_10695);
nand U13267 (N_13267,N_11447,N_11061);
nand U13268 (N_13268,N_11580,N_10689);
or U13269 (N_13269,N_10787,N_11689);
nor U13270 (N_13270,N_11047,N_11252);
nor U13271 (N_13271,N_11050,N_11609);
nor U13272 (N_13272,N_11524,N_10717);
or U13273 (N_13273,N_11559,N_10978);
nand U13274 (N_13274,N_11971,N_10591);
or U13275 (N_13275,N_10964,N_10715);
nor U13276 (N_13276,N_11246,N_11177);
xor U13277 (N_13277,N_11560,N_10767);
or U13278 (N_13278,N_11566,N_10651);
nand U13279 (N_13279,N_11196,N_11619);
or U13280 (N_13280,N_10899,N_10848);
or U13281 (N_13281,N_10535,N_11926);
nand U13282 (N_13282,N_11079,N_10628);
nand U13283 (N_13283,N_11212,N_10794);
nand U13284 (N_13284,N_11084,N_10855);
and U13285 (N_13285,N_11406,N_10858);
nand U13286 (N_13286,N_11163,N_11712);
nand U13287 (N_13287,N_11351,N_10876);
nor U13288 (N_13288,N_11363,N_11154);
and U13289 (N_13289,N_10722,N_10779);
nor U13290 (N_13290,N_11229,N_10572);
nor U13291 (N_13291,N_11640,N_11214);
or U13292 (N_13292,N_10926,N_11794);
nand U13293 (N_13293,N_10789,N_11894);
nor U13294 (N_13294,N_10645,N_11753);
nor U13295 (N_13295,N_11866,N_11772);
and U13296 (N_13296,N_11461,N_11689);
nor U13297 (N_13297,N_11565,N_11110);
or U13298 (N_13298,N_11520,N_11140);
or U13299 (N_13299,N_11089,N_11623);
and U13300 (N_13300,N_11159,N_10845);
or U13301 (N_13301,N_10767,N_10595);
or U13302 (N_13302,N_11939,N_11179);
nand U13303 (N_13303,N_11881,N_10795);
or U13304 (N_13304,N_11445,N_11244);
nor U13305 (N_13305,N_11514,N_11882);
nor U13306 (N_13306,N_10606,N_11118);
nor U13307 (N_13307,N_11993,N_11635);
nand U13308 (N_13308,N_10551,N_11943);
or U13309 (N_13309,N_10744,N_11943);
nand U13310 (N_13310,N_11891,N_10519);
nor U13311 (N_13311,N_11670,N_11533);
nand U13312 (N_13312,N_11232,N_10983);
or U13313 (N_13313,N_11091,N_11762);
nand U13314 (N_13314,N_11077,N_11529);
nand U13315 (N_13315,N_11763,N_11610);
nor U13316 (N_13316,N_11388,N_10541);
nand U13317 (N_13317,N_11181,N_11126);
and U13318 (N_13318,N_10982,N_11662);
and U13319 (N_13319,N_11665,N_11557);
nor U13320 (N_13320,N_11650,N_11228);
nor U13321 (N_13321,N_10661,N_11702);
and U13322 (N_13322,N_10576,N_11541);
nor U13323 (N_13323,N_11202,N_10804);
and U13324 (N_13324,N_10530,N_11927);
nor U13325 (N_13325,N_11067,N_10821);
nor U13326 (N_13326,N_11712,N_11349);
or U13327 (N_13327,N_11552,N_11574);
and U13328 (N_13328,N_10518,N_10601);
nand U13329 (N_13329,N_11457,N_10943);
nand U13330 (N_13330,N_10984,N_11983);
nand U13331 (N_13331,N_11502,N_11993);
or U13332 (N_13332,N_10946,N_10534);
nor U13333 (N_13333,N_11528,N_10807);
and U13334 (N_13334,N_11279,N_11345);
or U13335 (N_13335,N_11786,N_10853);
nand U13336 (N_13336,N_10823,N_10727);
nand U13337 (N_13337,N_10501,N_10744);
or U13338 (N_13338,N_11890,N_11055);
nand U13339 (N_13339,N_10662,N_11356);
or U13340 (N_13340,N_11922,N_11603);
nand U13341 (N_13341,N_10783,N_10521);
and U13342 (N_13342,N_11378,N_11799);
and U13343 (N_13343,N_11308,N_11092);
nand U13344 (N_13344,N_11323,N_11862);
or U13345 (N_13345,N_11495,N_10850);
nand U13346 (N_13346,N_10698,N_11354);
nand U13347 (N_13347,N_11104,N_10827);
nor U13348 (N_13348,N_10754,N_11381);
nand U13349 (N_13349,N_11958,N_11696);
nand U13350 (N_13350,N_10564,N_11985);
or U13351 (N_13351,N_10843,N_11178);
nand U13352 (N_13352,N_11837,N_10788);
nand U13353 (N_13353,N_11843,N_10978);
nand U13354 (N_13354,N_11599,N_11098);
and U13355 (N_13355,N_11589,N_10996);
or U13356 (N_13356,N_11558,N_11689);
or U13357 (N_13357,N_10769,N_11389);
or U13358 (N_13358,N_11344,N_10610);
nor U13359 (N_13359,N_10735,N_11020);
or U13360 (N_13360,N_10942,N_11081);
or U13361 (N_13361,N_11230,N_10805);
nor U13362 (N_13362,N_11066,N_11405);
nand U13363 (N_13363,N_11235,N_11588);
and U13364 (N_13364,N_10912,N_11355);
nand U13365 (N_13365,N_11628,N_11604);
or U13366 (N_13366,N_11769,N_11298);
nor U13367 (N_13367,N_11096,N_10545);
nand U13368 (N_13368,N_11476,N_11241);
nand U13369 (N_13369,N_11194,N_11233);
or U13370 (N_13370,N_11505,N_11481);
nand U13371 (N_13371,N_11288,N_11862);
or U13372 (N_13372,N_11811,N_10972);
or U13373 (N_13373,N_11366,N_11677);
and U13374 (N_13374,N_10688,N_10875);
nand U13375 (N_13375,N_10628,N_11746);
or U13376 (N_13376,N_11746,N_11269);
nor U13377 (N_13377,N_11040,N_10556);
nor U13378 (N_13378,N_10997,N_11195);
nand U13379 (N_13379,N_10504,N_11967);
nor U13380 (N_13380,N_11081,N_11841);
nand U13381 (N_13381,N_10708,N_11703);
nand U13382 (N_13382,N_11854,N_10868);
nor U13383 (N_13383,N_10601,N_10967);
nor U13384 (N_13384,N_11580,N_11954);
and U13385 (N_13385,N_11468,N_10513);
or U13386 (N_13386,N_11558,N_11567);
and U13387 (N_13387,N_11242,N_11194);
nand U13388 (N_13388,N_11082,N_11417);
nand U13389 (N_13389,N_10892,N_11561);
or U13390 (N_13390,N_11105,N_10516);
or U13391 (N_13391,N_11800,N_10560);
nand U13392 (N_13392,N_11028,N_10826);
and U13393 (N_13393,N_11017,N_10577);
and U13394 (N_13394,N_10724,N_10842);
or U13395 (N_13395,N_11978,N_11536);
and U13396 (N_13396,N_11204,N_10768);
or U13397 (N_13397,N_11324,N_11043);
or U13398 (N_13398,N_10951,N_10611);
nand U13399 (N_13399,N_11927,N_10766);
nand U13400 (N_13400,N_11845,N_10593);
nand U13401 (N_13401,N_11027,N_11239);
and U13402 (N_13402,N_10752,N_10560);
nor U13403 (N_13403,N_11321,N_11656);
and U13404 (N_13404,N_10642,N_10727);
nor U13405 (N_13405,N_11297,N_10954);
nand U13406 (N_13406,N_10755,N_11036);
xnor U13407 (N_13407,N_10503,N_11480);
and U13408 (N_13408,N_11506,N_11422);
nor U13409 (N_13409,N_11272,N_11302);
or U13410 (N_13410,N_11227,N_10913);
and U13411 (N_13411,N_11689,N_11836);
and U13412 (N_13412,N_10561,N_10970);
nor U13413 (N_13413,N_11881,N_11350);
nand U13414 (N_13414,N_11512,N_11546);
or U13415 (N_13415,N_11947,N_11220);
nor U13416 (N_13416,N_10756,N_10518);
nand U13417 (N_13417,N_11393,N_10506);
and U13418 (N_13418,N_11591,N_11809);
and U13419 (N_13419,N_11873,N_10805);
nand U13420 (N_13420,N_11155,N_10790);
nand U13421 (N_13421,N_10907,N_10542);
and U13422 (N_13422,N_10665,N_11966);
and U13423 (N_13423,N_11322,N_10534);
nor U13424 (N_13424,N_11900,N_10610);
or U13425 (N_13425,N_11695,N_11617);
nor U13426 (N_13426,N_11427,N_10804);
or U13427 (N_13427,N_11142,N_10763);
nor U13428 (N_13428,N_10612,N_10634);
nand U13429 (N_13429,N_11242,N_10518);
and U13430 (N_13430,N_11647,N_10755);
nand U13431 (N_13431,N_11561,N_10700);
and U13432 (N_13432,N_11855,N_11423);
and U13433 (N_13433,N_11736,N_10531);
nor U13434 (N_13434,N_10875,N_11835);
nor U13435 (N_13435,N_11322,N_11002);
or U13436 (N_13436,N_11904,N_11090);
and U13437 (N_13437,N_10796,N_10839);
nor U13438 (N_13438,N_10665,N_11706);
and U13439 (N_13439,N_11267,N_11265);
or U13440 (N_13440,N_11050,N_11645);
and U13441 (N_13441,N_10970,N_11696);
or U13442 (N_13442,N_11958,N_11317);
nor U13443 (N_13443,N_11941,N_11537);
nor U13444 (N_13444,N_11490,N_10715);
or U13445 (N_13445,N_10535,N_10521);
nand U13446 (N_13446,N_10559,N_11105);
nor U13447 (N_13447,N_10964,N_11662);
and U13448 (N_13448,N_11251,N_11383);
and U13449 (N_13449,N_11767,N_10794);
nor U13450 (N_13450,N_10663,N_11077);
or U13451 (N_13451,N_10732,N_10782);
or U13452 (N_13452,N_11432,N_10923);
or U13453 (N_13453,N_11033,N_11556);
nor U13454 (N_13454,N_11190,N_11011);
and U13455 (N_13455,N_10734,N_11843);
or U13456 (N_13456,N_11720,N_11971);
and U13457 (N_13457,N_11393,N_11573);
nor U13458 (N_13458,N_10674,N_11929);
nor U13459 (N_13459,N_10889,N_11223);
nor U13460 (N_13460,N_10745,N_11778);
nand U13461 (N_13461,N_11258,N_10812);
and U13462 (N_13462,N_11152,N_11253);
or U13463 (N_13463,N_11575,N_11024);
nand U13464 (N_13464,N_10902,N_11635);
or U13465 (N_13465,N_11542,N_10551);
nor U13466 (N_13466,N_10983,N_11627);
and U13467 (N_13467,N_10699,N_11180);
nor U13468 (N_13468,N_10967,N_11156);
nand U13469 (N_13469,N_10640,N_10687);
and U13470 (N_13470,N_11429,N_10649);
and U13471 (N_13471,N_11559,N_10989);
and U13472 (N_13472,N_11679,N_10680);
and U13473 (N_13473,N_10920,N_11236);
and U13474 (N_13474,N_11440,N_11546);
nand U13475 (N_13475,N_11975,N_11410);
and U13476 (N_13476,N_10821,N_10710);
nand U13477 (N_13477,N_11097,N_10873);
nor U13478 (N_13478,N_11979,N_10703);
and U13479 (N_13479,N_11233,N_11687);
nand U13480 (N_13480,N_11797,N_11848);
nor U13481 (N_13481,N_11656,N_11894);
nand U13482 (N_13482,N_10800,N_11339);
or U13483 (N_13483,N_10554,N_10856);
nor U13484 (N_13484,N_11617,N_10952);
nor U13485 (N_13485,N_10742,N_11991);
and U13486 (N_13486,N_10830,N_11151);
nand U13487 (N_13487,N_10797,N_11564);
nand U13488 (N_13488,N_11692,N_10649);
and U13489 (N_13489,N_10885,N_11683);
nand U13490 (N_13490,N_11746,N_11106);
and U13491 (N_13491,N_11142,N_10638);
xnor U13492 (N_13492,N_11508,N_10558);
nor U13493 (N_13493,N_10985,N_11100);
nor U13494 (N_13494,N_10696,N_11829);
or U13495 (N_13495,N_11896,N_10595);
and U13496 (N_13496,N_11442,N_11072);
nand U13497 (N_13497,N_11665,N_11500);
nand U13498 (N_13498,N_10905,N_11409);
nand U13499 (N_13499,N_11237,N_11542);
or U13500 (N_13500,N_12958,N_12297);
nand U13501 (N_13501,N_12032,N_12571);
nor U13502 (N_13502,N_12284,N_13439);
nor U13503 (N_13503,N_13253,N_12556);
and U13504 (N_13504,N_12871,N_12679);
nand U13505 (N_13505,N_12662,N_13410);
and U13506 (N_13506,N_13178,N_13122);
nor U13507 (N_13507,N_12031,N_13312);
xnor U13508 (N_13508,N_12083,N_12670);
nand U13509 (N_13509,N_13269,N_12413);
nor U13510 (N_13510,N_12071,N_12534);
nor U13511 (N_13511,N_13016,N_12653);
or U13512 (N_13512,N_12680,N_12451);
and U13513 (N_13513,N_13405,N_12993);
nand U13514 (N_13514,N_12580,N_12587);
nand U13515 (N_13515,N_13204,N_12875);
nor U13516 (N_13516,N_12314,N_13195);
or U13517 (N_13517,N_13088,N_12940);
and U13518 (N_13518,N_12305,N_12120);
nor U13519 (N_13519,N_12187,N_13048);
nor U13520 (N_13520,N_12595,N_13198);
or U13521 (N_13521,N_12416,N_13089);
nor U13522 (N_13522,N_12540,N_13466);
nand U13523 (N_13523,N_12462,N_12574);
and U13524 (N_13524,N_12447,N_13235);
nor U13525 (N_13525,N_12743,N_12589);
and U13526 (N_13526,N_12911,N_13185);
nor U13527 (N_13527,N_12172,N_13396);
xnor U13528 (N_13528,N_12912,N_12964);
and U13529 (N_13529,N_13033,N_12597);
or U13530 (N_13530,N_12735,N_12861);
nand U13531 (N_13531,N_12970,N_13031);
or U13532 (N_13532,N_12042,N_12768);
nand U13533 (N_13533,N_12212,N_12576);
nor U13534 (N_13534,N_13479,N_12424);
and U13535 (N_13535,N_12164,N_13177);
or U13536 (N_13536,N_13052,N_12019);
nand U13537 (N_13537,N_12084,N_12693);
nand U13538 (N_13538,N_12238,N_12064);
or U13539 (N_13539,N_12752,N_12464);
nand U13540 (N_13540,N_12866,N_12717);
or U13541 (N_13541,N_13142,N_13165);
and U13542 (N_13542,N_12517,N_13167);
and U13543 (N_13543,N_12489,N_13041);
nor U13544 (N_13544,N_12793,N_12005);
and U13545 (N_13545,N_12332,N_12971);
or U13546 (N_13546,N_13050,N_12343);
nand U13547 (N_13547,N_12420,N_12758);
nor U13548 (N_13548,N_13112,N_12727);
nor U13549 (N_13549,N_12180,N_12355);
nand U13550 (N_13550,N_13153,N_12431);
nand U13551 (N_13551,N_12062,N_13444);
or U13552 (N_13552,N_12614,N_12224);
nand U13553 (N_13553,N_12381,N_12272);
and U13554 (N_13554,N_12117,N_12983);
or U13555 (N_13555,N_12454,N_12530);
or U13556 (N_13556,N_12754,N_12926);
and U13557 (N_13557,N_13302,N_13378);
nor U13558 (N_13558,N_13124,N_13111);
or U13559 (N_13559,N_12229,N_12857);
or U13560 (N_13560,N_12661,N_12873);
nand U13561 (N_13561,N_13386,N_12476);
nor U13562 (N_13562,N_13313,N_12006);
nand U13563 (N_13563,N_13193,N_12022);
and U13564 (N_13564,N_12444,N_12872);
nor U13565 (N_13565,N_13242,N_13243);
nand U13566 (N_13566,N_12979,N_13449);
nor U13567 (N_13567,N_12880,N_13373);
or U13568 (N_13568,N_12591,N_12546);
or U13569 (N_13569,N_13435,N_12050);
nor U13570 (N_13570,N_12613,N_12354);
nand U13571 (N_13571,N_13331,N_13343);
or U13572 (N_13572,N_13416,N_12065);
and U13573 (N_13573,N_12425,N_13457);
xnor U13574 (N_13574,N_12992,N_12706);
and U13575 (N_13575,N_13446,N_12897);
nor U13576 (N_13576,N_12646,N_12266);
nor U13577 (N_13577,N_12584,N_13398);
or U13578 (N_13578,N_12103,N_13200);
nor U13579 (N_13579,N_13319,N_12449);
or U13580 (N_13580,N_12577,N_13003);
nor U13581 (N_13581,N_13450,N_12667);
nor U13582 (N_13582,N_12426,N_13379);
and U13583 (N_13583,N_12533,N_13275);
nand U13584 (N_13584,N_12058,N_12977);
nor U13585 (N_13585,N_12835,N_12500);
nor U13586 (N_13586,N_12807,N_13158);
nand U13587 (N_13587,N_13082,N_13293);
nor U13588 (N_13588,N_12891,N_12815);
nand U13589 (N_13589,N_13064,N_12460);
and U13590 (N_13590,N_12157,N_12719);
or U13591 (N_13591,N_12326,N_12626);
and U13592 (N_13592,N_12619,N_13186);
or U13593 (N_13593,N_12986,N_12487);
nand U13594 (N_13594,N_12887,N_13072);
nand U13595 (N_13595,N_12568,N_12852);
or U13596 (N_13596,N_12927,N_12257);
or U13597 (N_13597,N_13078,N_12353);
and U13598 (N_13598,N_12731,N_12784);
or U13599 (N_13599,N_13197,N_13125);
nand U13600 (N_13600,N_13203,N_12602);
or U13601 (N_13601,N_12292,N_12247);
or U13602 (N_13602,N_12030,N_13277);
or U13603 (N_13603,N_13465,N_12664);
and U13604 (N_13604,N_12683,N_13094);
or U13605 (N_13605,N_12124,N_12078);
nor U13606 (N_13606,N_12913,N_12729);
nor U13607 (N_13607,N_13256,N_13037);
nand U13608 (N_13608,N_13014,N_13029);
nor U13609 (N_13609,N_13406,N_12672);
or U13610 (N_13610,N_12269,N_13420);
nand U13611 (N_13611,N_12041,N_13495);
and U13612 (N_13612,N_12251,N_12328);
nand U13613 (N_13613,N_12561,N_13464);
or U13614 (N_13614,N_13104,N_12834);
nor U13615 (N_13615,N_12162,N_12601);
nor U13616 (N_13616,N_12151,N_13325);
nand U13617 (N_13617,N_12175,N_13120);
and U13618 (N_13618,N_12053,N_12287);
and U13619 (N_13619,N_12553,N_12982);
nand U13620 (N_13620,N_12099,N_12944);
and U13621 (N_13621,N_12824,N_12308);
nand U13622 (N_13622,N_13443,N_13447);
and U13623 (N_13623,N_12557,N_12712);
xnor U13624 (N_13624,N_12169,N_12551);
and U13625 (N_13625,N_12780,N_13494);
nor U13626 (N_13626,N_12787,N_12294);
nor U13627 (N_13627,N_13413,N_13338);
nor U13628 (N_13628,N_12635,N_13482);
and U13629 (N_13629,N_12480,N_12973);
nor U13630 (N_13630,N_12318,N_13045);
xor U13631 (N_13631,N_13423,N_12077);
nor U13632 (N_13632,N_12087,N_12773);
and U13633 (N_13633,N_12627,N_12119);
or U13634 (N_13634,N_13210,N_12737);
and U13635 (N_13635,N_12280,N_12265);
nor U13636 (N_13636,N_12324,N_13425);
and U13637 (N_13637,N_13141,N_12583);
and U13638 (N_13638,N_12378,N_13005);
or U13639 (N_13639,N_12302,N_12252);
nand U13640 (N_13640,N_12230,N_12094);
or U13641 (N_13641,N_12437,N_13261);
and U13642 (N_13642,N_12611,N_13404);
or U13643 (N_13643,N_12446,N_12313);
nand U13644 (N_13644,N_13222,N_13147);
or U13645 (N_13645,N_12904,N_13365);
or U13646 (N_13646,N_13062,N_12366);
or U13647 (N_13647,N_13012,N_12732);
nor U13648 (N_13648,N_13421,N_12137);
and U13649 (N_13649,N_12849,N_12772);
nor U13650 (N_13650,N_12063,N_13305);
or U13651 (N_13651,N_13021,N_12610);
and U13652 (N_13652,N_12967,N_13399);
nor U13653 (N_13653,N_12928,N_12660);
or U13654 (N_13654,N_13392,N_13179);
nor U13655 (N_13655,N_13192,N_12337);
and U13656 (N_13656,N_12586,N_12696);
or U13657 (N_13657,N_12937,N_13170);
and U13658 (N_13658,N_12036,N_12359);
nor U13659 (N_13659,N_12996,N_12742);
and U13660 (N_13660,N_12703,N_13451);
and U13661 (N_13661,N_12908,N_12502);
or U13662 (N_13662,N_13300,N_12300);
nor U13663 (N_13663,N_13391,N_12628);
nor U13664 (N_13664,N_12917,N_12612);
and U13665 (N_13665,N_12794,N_12692);
or U13666 (N_13666,N_12396,N_12014);
xor U13667 (N_13667,N_12532,N_12310);
or U13668 (N_13668,N_12263,N_12342);
and U13669 (N_13669,N_12514,N_12216);
nor U13670 (N_13670,N_12286,N_12725);
nor U13671 (N_13671,N_13131,N_12405);
nand U13672 (N_13672,N_12105,N_12980);
nor U13673 (N_13673,N_12631,N_12878);
and U13674 (N_13674,N_12622,N_12235);
and U13675 (N_13675,N_13267,N_13206);
nor U13676 (N_13676,N_12192,N_12419);
nor U13677 (N_13677,N_13299,N_12903);
nand U13678 (N_13678,N_13220,N_13426);
nand U13679 (N_13679,N_12461,N_12828);
nor U13680 (N_13680,N_12620,N_12002);
and U13681 (N_13681,N_12633,N_12141);
nand U13682 (N_13682,N_12562,N_13344);
nand U13683 (N_13683,N_12255,N_13481);
or U13684 (N_13684,N_12630,N_12649);
nand U13685 (N_13685,N_13184,N_12285);
or U13686 (N_13686,N_13057,N_13250);
nor U13687 (N_13687,N_12325,N_12496);
or U13688 (N_13688,N_12097,N_13237);
nand U13689 (N_13689,N_12320,N_12290);
nand U13690 (N_13690,N_12443,N_12629);
nand U13691 (N_13691,N_13294,N_12155);
and U13692 (N_13692,N_12091,N_12775);
nor U13693 (N_13693,N_13211,N_13321);
or U13694 (N_13694,N_12185,N_12881);
nand U13695 (N_13695,N_12985,N_12563);
or U13696 (N_13696,N_12380,N_13164);
nor U13697 (N_13697,N_13295,N_12195);
or U13698 (N_13698,N_13252,N_12723);
and U13699 (N_13699,N_12015,N_13334);
and U13700 (N_13700,N_13232,N_13341);
nor U13701 (N_13701,N_13355,N_12767);
and U13702 (N_13702,N_12067,N_12851);
or U13703 (N_13703,N_12746,N_12573);
nand U13704 (N_13704,N_12104,N_13049);
and U13705 (N_13705,N_13118,N_12037);
and U13706 (N_13706,N_12818,N_12375);
or U13707 (N_13707,N_13219,N_12177);
nand U13708 (N_13708,N_13051,N_12919);
nand U13709 (N_13709,N_12499,N_12778);
nand U13710 (N_13710,N_12412,N_12028);
or U13711 (N_13711,N_12435,N_12469);
or U13712 (N_13712,N_12946,N_12156);
and U13713 (N_13713,N_13463,N_12060);
nand U13714 (N_13714,N_12678,N_12808);
nand U13715 (N_13715,N_12289,N_12181);
nor U13716 (N_13716,N_12239,N_12007);
nand U13717 (N_13717,N_13440,N_12669);
xor U13718 (N_13718,N_12021,N_13485);
nand U13719 (N_13719,N_12508,N_13226);
and U13720 (N_13720,N_13079,N_12429);
nor U13721 (N_13721,N_12962,N_13090);
nand U13722 (N_13722,N_13159,N_13462);
and U13723 (N_13723,N_12483,N_12167);
nand U13724 (N_13724,N_12704,N_12129);
nor U13725 (N_13725,N_12714,N_13401);
and U13726 (N_13726,N_13239,N_13214);
or U13727 (N_13727,N_13453,N_12080);
nor U13728 (N_13728,N_12760,N_12234);
and U13729 (N_13729,N_12459,N_12865);
or U13730 (N_13730,N_12074,N_12275);
nor U13731 (N_13731,N_12625,N_12995);
nor U13732 (N_13732,N_13070,N_12186);
nand U13733 (N_13733,N_12513,N_13017);
nand U13734 (N_13734,N_13286,N_12659);
or U13735 (N_13735,N_13136,N_12505);
nor U13736 (N_13736,N_13077,N_12322);
nand U13737 (N_13737,N_12855,N_13417);
nand U13738 (N_13738,N_12733,N_12932);
xnor U13739 (N_13739,N_13081,N_13455);
and U13740 (N_13740,N_13004,N_12203);
or U13741 (N_13741,N_12999,N_12319);
nor U13742 (N_13742,N_13274,N_12018);
nand U13743 (N_13743,N_12945,N_12528);
or U13744 (N_13744,N_12825,N_12895);
nor U13745 (N_13745,N_13486,N_13139);
and U13746 (N_13746,N_13095,N_12641);
and U13747 (N_13747,N_13032,N_13329);
or U13748 (N_13748,N_12843,N_12406);
or U13749 (N_13749,N_12930,N_12814);
nand U13750 (N_13750,N_13058,N_13236);
nor U13751 (N_13751,N_13161,N_13388);
or U13752 (N_13752,N_12552,N_13061);
or U13753 (N_13753,N_13225,N_12484);
nor U13754 (N_13754,N_12038,N_12700);
nand U13755 (N_13755,N_13075,N_12228);
and U13756 (N_13756,N_12914,N_12202);
or U13757 (N_13757,N_12312,N_12535);
xor U13758 (N_13758,N_12541,N_12456);
or U13759 (N_13759,N_12076,N_13475);
and U13760 (N_13760,N_12518,N_12997);
or U13761 (N_13761,N_12373,N_13359);
nand U13762 (N_13762,N_13209,N_12841);
and U13763 (N_13763,N_12095,N_12766);
nor U13764 (N_13764,N_12596,N_13469);
nor U13765 (N_13765,N_13011,N_12870);
and U13766 (N_13766,N_13007,N_12923);
nand U13767 (N_13767,N_12522,N_12278);
nand U13768 (N_13768,N_13073,N_12968);
nand U13769 (N_13769,N_12386,N_12369);
and U13770 (N_13770,N_12242,N_12165);
nand U13771 (N_13771,N_13454,N_12890);
nand U13772 (N_13772,N_12604,N_12829);
nor U13773 (N_13773,N_12013,N_12127);
or U13774 (N_13774,N_12194,N_12182);
and U13775 (N_13775,N_12267,N_13411);
nand U13776 (N_13776,N_13370,N_13493);
or U13777 (N_13777,N_12298,N_12368);
or U13778 (N_13778,N_12581,N_12491);
nand U13779 (N_13779,N_12455,N_13148);
and U13780 (N_13780,N_13318,N_12174);
nand U13781 (N_13781,N_12889,N_12020);
and U13782 (N_13782,N_12391,N_12309);
nand U13783 (N_13783,N_12774,N_12362);
nor U13784 (N_13784,N_13445,N_12045);
nor U13785 (N_13785,N_12140,N_12722);
nand U13786 (N_13786,N_13102,N_13489);
nor U13787 (N_13787,N_12833,N_13162);
and U13788 (N_13788,N_12521,N_12385);
and U13789 (N_13789,N_13208,N_12874);
nor U13790 (N_13790,N_12902,N_12218);
and U13791 (N_13791,N_12321,N_12184);
nand U13792 (N_13792,N_13149,N_12920);
or U13793 (N_13793,N_13430,N_12507);
nand U13794 (N_13794,N_12941,N_13452);
and U13795 (N_13795,N_12658,N_12179);
nor U13796 (N_13796,N_13163,N_13393);
nor U13797 (N_13797,N_12283,N_12981);
nor U13798 (N_13798,N_12801,N_13157);
nor U13799 (N_13799,N_13096,N_12954);
or U13800 (N_13800,N_13191,N_12131);
or U13801 (N_13801,N_13087,N_13020);
nand U13802 (N_13802,N_12204,N_12044);
nand U13803 (N_13803,N_12671,N_12868);
and U13804 (N_13804,N_12243,N_12423);
nand U13805 (N_13805,N_13205,N_13327);
nor U13806 (N_13806,N_12106,N_12757);
or U13807 (N_13807,N_13030,N_12748);
or U13808 (N_13808,N_12466,N_13431);
and U13809 (N_13809,N_13044,N_13459);
nor U13810 (N_13810,N_12279,N_13074);
nand U13811 (N_13811,N_12925,N_13255);
nand U13812 (N_13812,N_12519,N_13429);
nand U13813 (N_13813,N_12952,N_12142);
and U13814 (N_13814,N_13212,N_12883);
nand U13815 (N_13815,N_12682,N_12107);
nor U13816 (N_13816,N_13105,N_13369);
or U13817 (N_13817,N_13437,N_12860);
nor U13818 (N_13818,N_13434,N_12809);
and U13819 (N_13819,N_12598,N_12295);
nor U13820 (N_13820,N_12245,N_13085);
nor U13821 (N_13821,N_12751,N_12512);
nor U13822 (N_13822,N_12492,N_12072);
and U13823 (N_13823,N_13172,N_12341);
or U13824 (N_13824,N_12531,N_12388);
and U13825 (N_13825,N_12850,N_12728);
nor U13826 (N_13826,N_13291,N_13251);
and U13827 (N_13827,N_13320,N_12158);
xor U13828 (N_13828,N_12804,N_12178);
or U13829 (N_13829,N_12356,N_13332);
nand U13830 (N_13830,N_12989,N_12008);
and U13831 (N_13831,N_12351,N_12035);
nor U13832 (N_13832,N_12197,N_12972);
and U13833 (N_13833,N_12544,N_12974);
nand U13834 (N_13834,N_12582,N_12088);
or U13835 (N_13835,N_13173,N_12494);
nor U13836 (N_13836,N_13477,N_13352);
nor U13837 (N_13837,N_12839,N_12066);
and U13838 (N_13838,N_13397,N_13015);
or U13839 (N_13839,N_12826,N_12009);
or U13840 (N_13840,N_12436,N_12741);
or U13841 (N_13841,N_12542,N_13377);
nand U13842 (N_13842,N_12593,N_12191);
or U13843 (N_13843,N_12608,N_12948);
nand U13844 (N_13844,N_12276,N_13068);
nand U13845 (N_13845,N_12303,N_12951);
or U13846 (N_13846,N_12707,N_12208);
nand U13847 (N_13847,N_13385,N_12526);
nand U13848 (N_13848,N_13035,N_12575);
nor U13849 (N_13849,N_12905,N_12811);
and U13850 (N_13850,N_12372,N_12410);
or U13851 (N_13851,N_12475,N_13171);
nor U13852 (N_13852,N_12114,N_12585);
nor U13853 (N_13853,N_12827,N_13137);
and U13854 (N_13854,N_12331,N_12984);
or U13855 (N_13855,N_13353,N_12070);
and U13856 (N_13856,N_12567,N_12588);
and U13857 (N_13857,N_13133,N_13436);
nand U13858 (N_13858,N_12349,N_12665);
and U13859 (N_13859,N_13376,N_12956);
nor U13860 (N_13860,N_13174,N_12893);
and U13861 (N_13861,N_13292,N_12219);
and U13862 (N_13862,N_12291,N_12632);
and U13863 (N_13863,N_13038,N_13263);
or U13864 (N_13864,N_13117,N_12790);
nand U13865 (N_13865,N_13474,N_13483);
nor U13866 (N_13866,N_12404,N_13181);
nor U13867 (N_13867,N_13428,N_12691);
nor U13868 (N_13868,N_13375,N_13180);
nor U13869 (N_13869,N_12441,N_13116);
nand U13870 (N_13870,N_12501,N_12495);
nor U13871 (N_13871,N_12138,N_13264);
and U13872 (N_13872,N_12490,N_12763);
and U13873 (N_13873,N_12323,N_12188);
nand U13874 (N_13874,N_12040,N_12756);
and U13875 (N_13875,N_12493,N_12217);
nor U13876 (N_13876,N_12110,N_12987);
and U13877 (N_13877,N_13281,N_12086);
or U13878 (N_13878,N_12916,N_12953);
nand U13879 (N_13879,N_12547,N_13478);
nor U13880 (N_13880,N_13254,N_13340);
nor U13881 (N_13881,N_12685,N_12001);
or U13882 (N_13882,N_13298,N_12761);
nand U13883 (N_13883,N_12000,N_12467);
or U13884 (N_13884,N_12259,N_12102);
and U13885 (N_13885,N_12736,N_12716);
or U13886 (N_13886,N_13339,N_13187);
nand U13887 (N_13887,N_12592,N_12783);
nor U13888 (N_13888,N_12856,N_12233);
and U13889 (N_13889,N_12214,N_13155);
nand U13890 (N_13890,N_13154,N_12200);
nand U13891 (N_13891,N_12688,N_12838);
nor U13892 (N_13892,N_12145,N_12039);
and U13893 (N_13893,N_12689,N_13488);
nor U13894 (N_13894,N_13306,N_12821);
nand U13895 (N_13895,N_12207,N_13093);
nand U13896 (N_13896,N_13019,N_12847);
and U13897 (N_13897,N_12432,N_12133);
or U13898 (N_13898,N_12618,N_12663);
and U13899 (N_13899,N_12211,N_12550);
nor U13900 (N_13900,N_13227,N_12643);
or U13901 (N_13901,N_12894,N_12777);
and U13902 (N_13902,N_13394,N_12477);
nor U13903 (N_13903,N_12786,N_13498);
nand U13904 (N_13904,N_12428,N_12089);
nand U13905 (N_13905,N_13266,N_12740);
or U13906 (N_13906,N_13099,N_13301);
nor U13907 (N_13907,N_12198,N_13207);
nand U13908 (N_13908,N_12196,N_12049);
nand U13909 (N_13909,N_13188,N_12651);
nor U13910 (N_13910,N_13107,N_12918);
nor U13911 (N_13911,N_12260,N_12832);
nor U13912 (N_13912,N_12150,N_13040);
and U13913 (N_13913,N_12118,N_12422);
and U13914 (N_13914,N_12885,N_12011);
nor U13915 (N_13915,N_13309,N_12527);
and U13916 (N_13916,N_12896,N_13471);
and U13917 (N_13917,N_12055,N_12674);
or U13918 (N_13918,N_13328,N_12112);
xor U13919 (N_13919,N_12402,N_12176);
nand U13920 (N_13920,N_12210,N_13336);
nor U13921 (N_13921,N_13092,N_12148);
nor U13922 (N_13922,N_12485,N_12092);
and U13923 (N_13923,N_13345,N_12609);
nand U13924 (N_13924,N_13333,N_13350);
nand U13925 (N_13925,N_12430,N_12572);
nor U13926 (N_13926,N_12976,N_13043);
and U13927 (N_13927,N_13221,N_12545);
nor U13928 (N_13928,N_12082,N_12636);
nor U13929 (N_13929,N_13067,N_13348);
or U13930 (N_13930,N_12046,N_13432);
or U13931 (N_13931,N_12166,N_12606);
nand U13932 (N_13932,N_12858,N_12458);
nand U13933 (N_13933,N_12085,N_13366);
nand U13934 (N_13934,N_13395,N_12788);
xor U13935 (N_13935,N_12034,N_13156);
nor U13936 (N_13936,N_12600,N_12753);
nand U13937 (N_13937,N_12258,N_13260);
nor U13938 (N_13938,N_13065,N_13458);
xnor U13939 (N_13939,N_12048,N_13484);
and U13940 (N_13940,N_13280,N_12509);
nor U13941 (N_13941,N_12241,N_12327);
or U13942 (N_13942,N_12959,N_12549);
and U13943 (N_13943,N_12755,N_13314);
nor U13944 (N_13944,N_13060,N_12524);
nand U13945 (N_13945,N_12950,N_12189);
nor U13946 (N_13946,N_12361,N_12069);
or U13947 (N_13947,N_12296,N_13361);
and U13948 (N_13948,N_12307,N_12739);
and U13949 (N_13949,N_13130,N_12853);
nand U13950 (N_13950,N_12061,N_13380);
and U13951 (N_13951,N_13407,N_12957);
nand U13952 (N_13952,N_13080,N_13389);
or U13953 (N_13953,N_13316,N_13135);
nor U13954 (N_13954,N_12122,N_12975);
nand U13955 (N_13955,N_12384,N_13113);
and U13956 (N_13956,N_12599,N_12473);
nand U13957 (N_13957,N_13091,N_13084);
nand U13958 (N_13958,N_13476,N_12900);
nor U13959 (N_13959,N_12656,N_12299);
or U13960 (N_13960,N_13330,N_13472);
or U13961 (N_13961,N_13390,N_13169);
or U13962 (N_13962,N_12666,N_12935);
nor U13963 (N_13963,N_12539,N_12075);
nand U13964 (N_13964,N_13103,N_12647);
and U13965 (N_13965,N_12223,N_13216);
nand U13966 (N_13966,N_12393,N_12877);
nor U13967 (N_13967,N_12374,N_12910);
nor U13968 (N_13968,N_12803,N_12650);
and U13969 (N_13969,N_13363,N_13461);
nor U13970 (N_13970,N_12781,N_13114);
nand U13971 (N_13971,N_13145,N_13128);
or U13972 (N_13972,N_12261,N_12338);
nand U13973 (N_13973,N_12639,N_12056);
nand U13974 (N_13974,N_13046,N_13190);
or U13975 (N_13975,N_12498,N_13490);
nor U13976 (N_13976,N_12859,N_13354);
nand U13977 (N_13977,N_12816,N_12411);
and U13978 (N_13978,N_13071,N_13276);
or U13979 (N_13979,N_12677,N_12559);
and U13980 (N_13980,N_12281,N_13231);
and U13981 (N_13981,N_13422,N_12370);
or U13982 (N_13982,N_12511,N_13168);
and U13983 (N_13983,N_13056,N_12115);
and U13984 (N_13984,N_12068,N_12869);
or U13985 (N_13985,N_13047,N_12699);
or U13986 (N_13986,N_12565,N_13460);
or U13987 (N_13987,N_12607,N_12594);
or U13988 (N_13988,N_12470,N_13244);
and U13989 (N_13989,N_13194,N_12147);
and U13990 (N_13990,N_13418,N_12364);
or U13991 (N_13991,N_12315,N_13335);
xor U13992 (N_13992,N_13438,N_12906);
or U13993 (N_13993,N_13287,N_12515);
and U13994 (N_13994,N_13109,N_12796);
and U13995 (N_13995,N_12603,N_13022);
and U13996 (N_13996,N_13217,N_12116);
or U13997 (N_13997,N_13097,N_12392);
nor U13998 (N_13998,N_13372,N_12701);
nor U13999 (N_13999,N_13403,N_13262);
nand U14000 (N_14000,N_13360,N_12134);
or U14001 (N_14001,N_13152,N_12543);
or U14002 (N_14002,N_12990,N_12390);
nor U14003 (N_14003,N_12317,N_13289);
nor U14004 (N_14004,N_12398,N_12170);
nor U14005 (N_14005,N_12109,N_12724);
nand U14006 (N_14006,N_12352,N_12497);
nor U14007 (N_14007,N_13034,N_12350);
or U14008 (N_14008,N_12854,N_12282);
and U14009 (N_14009,N_12798,N_13166);
and U14010 (N_14010,N_12418,N_13183);
and U14011 (N_14011,N_13101,N_13025);
nand U14012 (N_14012,N_12249,N_13042);
and U14013 (N_14013,N_12765,N_12132);
and U14014 (N_14014,N_13026,N_12795);
nand U14015 (N_14015,N_12898,N_13229);
and U14016 (N_14016,N_12668,N_12744);
and U14017 (N_14017,N_13356,N_13351);
nand U14018 (N_14018,N_12879,N_12867);
or U14019 (N_14019,N_12270,N_13146);
or U14020 (N_14020,N_12655,N_12504);
or U14021 (N_14021,N_12478,N_12942);
nor U14022 (N_14022,N_13224,N_12922);
or U14023 (N_14023,N_12394,N_12779);
and U14024 (N_14024,N_12383,N_12407);
and U14025 (N_14025,N_12143,N_13241);
and U14026 (N_14026,N_12250,N_12336);
and U14027 (N_14027,N_13382,N_13108);
and U14028 (N_14028,N_12471,N_12654);
nor U14029 (N_14029,N_12335,N_12448);
or U14030 (N_14030,N_12345,N_13134);
and U14031 (N_14031,N_12222,N_12797);
and U14032 (N_14032,N_13246,N_12966);
and U14033 (N_14033,N_12876,N_12246);
nand U14034 (N_14034,N_12749,N_13470);
nand U14035 (N_14035,N_12360,N_12025);
or U14036 (N_14036,N_13324,N_13265);
and U14037 (N_14037,N_12991,N_12316);
and U14038 (N_14038,N_12227,N_12738);
nand U14039 (N_14039,N_13018,N_12111);
nand U14040 (N_14040,N_12033,N_12311);
nand U14041 (N_14041,N_12558,N_12820);
and U14042 (N_14042,N_12718,N_12408);
and U14043 (N_14043,N_13381,N_13115);
nand U14044 (N_14044,N_12560,N_13315);
or U14045 (N_14045,N_13303,N_12884);
nand U14046 (N_14046,N_12745,N_12657);
and U14047 (N_14047,N_12135,N_12256);
nand U14048 (N_14048,N_12482,N_12004);
and U14049 (N_14049,N_13409,N_13002);
nor U14050 (N_14050,N_12205,N_12675);
or U14051 (N_14051,N_12776,N_12268);
and U14052 (N_14052,N_12330,N_12367);
or U14053 (N_14053,N_12254,N_12943);
nand U14054 (N_14054,N_13419,N_13346);
or U14055 (N_14055,N_13027,N_13240);
or U14056 (N_14056,N_12822,N_13233);
nor U14057 (N_14057,N_13467,N_12506);
nor U14058 (N_14058,N_12273,N_13283);
nand U14059 (N_14059,N_13000,N_13151);
or U14060 (N_14060,N_13342,N_13066);
and U14061 (N_14061,N_12523,N_13387);
and U14062 (N_14062,N_13001,N_13383);
nor U14063 (N_14063,N_12800,N_12277);
or U14064 (N_14064,N_12438,N_12810);
or U14065 (N_14065,N_12376,N_13371);
nand U14066 (N_14066,N_13491,N_12427);
or U14067 (N_14067,N_12555,N_12329);
or U14068 (N_14068,N_12149,N_12481);
or U14069 (N_14069,N_13121,N_12785);
and U14070 (N_14070,N_13028,N_12848);
or U14071 (N_14071,N_13023,N_13110);
xor U14072 (N_14072,N_12802,N_13083);
nand U14073 (N_14073,N_12813,N_13189);
or U14074 (N_14074,N_12347,N_13323);
and U14075 (N_14075,N_12488,N_13347);
nand U14076 (N_14076,N_12965,N_12173);
and U14077 (N_14077,N_12711,N_13278);
or U14078 (N_14078,N_12949,N_12845);
and U14079 (N_14079,N_12715,N_13234);
or U14080 (N_14080,N_12365,N_12590);
nand U14081 (N_14081,N_12792,N_12823);
and U14082 (N_14082,N_12433,N_12623);
and U14083 (N_14083,N_13473,N_13296);
or U14084 (N_14084,N_12193,N_12747);
or U14085 (N_14085,N_13076,N_12403);
and U14086 (N_14086,N_12634,N_12371);
nor U14087 (N_14087,N_12171,N_12769);
nand U14088 (N_14088,N_12024,N_12452);
and U14089 (N_14089,N_12817,N_12998);
nand U14090 (N_14090,N_12450,N_13364);
and U14091 (N_14091,N_13009,N_12921);
or U14092 (N_14092,N_13055,N_12840);
nand U14093 (N_14093,N_12750,N_13129);
and U14094 (N_14094,N_12789,N_12695);
xnor U14095 (N_14095,N_12253,N_12694);
and U14096 (N_14096,N_12421,N_12215);
nor U14097 (N_14097,N_12615,N_12348);
or U14098 (N_14098,N_12225,N_12882);
or U14099 (N_14099,N_12924,N_12358);
or U14100 (N_14100,N_12782,N_13322);
nor U14101 (N_14101,N_12762,N_13215);
or U14102 (N_14102,N_13272,N_12554);
or U14103 (N_14103,N_12676,N_12096);
xnor U14104 (N_14104,N_13349,N_12529);
or U14105 (N_14105,N_12201,N_13326);
nor U14106 (N_14106,N_12862,N_12909);
nand U14107 (N_14107,N_12363,N_12648);
and U14108 (N_14108,N_12486,N_13006);
nor U14109 (N_14109,N_12791,N_13127);
nor U14110 (N_14110,N_13268,N_12548);
and U14111 (N_14111,N_12579,N_12799);
nand U14112 (N_14112,N_12244,N_13468);
or U14113 (N_14113,N_12346,N_12136);
nor U14114 (N_14114,N_13213,N_12090);
nand U14115 (N_14115,N_13400,N_13245);
nor U14116 (N_14116,N_12934,N_13013);
nor U14117 (N_14117,N_12113,N_12831);
nor U14118 (N_14118,N_13288,N_12213);
and U14119 (N_14119,N_12713,N_12726);
nand U14120 (N_14120,N_12963,N_13448);
and U14121 (N_14121,N_12183,N_12538);
or U14122 (N_14122,N_12933,N_13140);
nand U14123 (N_14123,N_12415,N_13238);
or U14124 (N_14124,N_13182,N_13308);
nand U14125 (N_14125,N_12293,N_12100);
nand U14126 (N_14126,N_13259,N_13499);
nor U14127 (N_14127,N_13492,N_12616);
nand U14128 (N_14128,N_12969,N_13271);
nand U14129 (N_14129,N_13441,N_13039);
nor U14130 (N_14130,N_12929,N_12644);
and U14131 (N_14131,N_12520,N_12720);
nand U14132 (N_14132,N_12624,N_12079);
or U14133 (N_14133,N_12463,N_12721);
and U14134 (N_14134,N_12709,N_13427);
nand U14135 (N_14135,N_12029,N_12566);
nand U14136 (N_14136,N_12051,N_12027);
or U14137 (N_14137,N_12231,N_12026);
or U14138 (N_14138,N_12901,N_12387);
nand U14139 (N_14139,N_13414,N_12564);
or U14140 (N_14140,N_12168,N_12805);
or U14141 (N_14141,N_12771,N_12569);
or U14142 (N_14142,N_13100,N_12409);
nand U14143 (N_14143,N_12395,N_12144);
and U14144 (N_14144,N_13098,N_12240);
nand U14145 (N_14145,N_13456,N_12708);
nor U14146 (N_14146,N_12130,N_13010);
or U14147 (N_14147,N_12899,N_13201);
nand U14148 (N_14148,N_12237,N_12988);
nand U14149 (N_14149,N_12264,N_12578);
and U14150 (N_14150,N_12047,N_13230);
and U14151 (N_14151,N_12907,N_12819);
and U14152 (N_14152,N_12125,N_13358);
nand U14153 (N_14153,N_13059,N_12764);
nand U14154 (N_14154,N_13284,N_12401);
nor U14155 (N_14155,N_12262,N_12479);
and U14156 (N_14156,N_12734,N_12536);
or U14157 (N_14157,N_12888,N_12012);
nor U14158 (N_14158,N_12864,N_12093);
or U14159 (N_14159,N_13176,N_12161);
and U14160 (N_14160,N_12468,N_12377);
and U14161 (N_14161,N_12304,N_12414);
nor U14162 (N_14162,N_12570,N_13160);
nand U14163 (N_14163,N_13218,N_12994);
nand U14164 (N_14164,N_12121,N_12209);
or U14165 (N_14165,N_13496,N_13487);
nor U14166 (N_14166,N_13384,N_12961);
nand U14167 (N_14167,N_13368,N_12759);
nor U14168 (N_14168,N_12221,N_12842);
or U14169 (N_14169,N_13270,N_12220);
and U14170 (N_14170,N_13279,N_12503);
and U14171 (N_14171,N_12640,N_13126);
or U14172 (N_14172,N_12730,N_12915);
nand U14173 (N_14173,N_12206,N_12417);
or U14174 (N_14174,N_12434,N_12248);
or U14175 (N_14175,N_12139,N_12770);
and U14176 (N_14176,N_13442,N_12698);
nor U14177 (N_14177,N_13036,N_13196);
or U14178 (N_14178,N_12152,N_13337);
nor U14179 (N_14179,N_13424,N_13285);
nor U14180 (N_14180,N_12806,N_12016);
nand U14181 (N_14181,N_13412,N_12003);
or U14182 (N_14182,N_12023,N_13024);
or U14183 (N_14183,N_13273,N_12525);
nand U14184 (N_14184,N_12445,N_12108);
nor U14185 (N_14185,N_12605,N_12710);
or U14186 (N_14186,N_13199,N_12637);
nor U14187 (N_14187,N_12306,N_13175);
nand U14188 (N_14188,N_12081,N_13053);
and U14189 (N_14189,N_13480,N_13063);
nor U14190 (N_14190,N_12043,N_13317);
nand U14191 (N_14191,N_12397,N_12516);
nor U14192 (N_14192,N_12334,N_12936);
nand U14193 (N_14193,N_12271,N_12153);
or U14194 (N_14194,N_13304,N_12339);
nand U14195 (N_14195,N_12098,N_13249);
nand U14196 (N_14196,N_12690,N_12301);
and U14197 (N_14197,N_12379,N_13144);
nand U14198 (N_14198,N_13311,N_13290);
or U14199 (N_14199,N_13282,N_13106);
nor U14200 (N_14200,N_13202,N_12190);
nor U14201 (N_14201,N_12126,N_12389);
nor U14202 (N_14202,N_12621,N_12681);
or U14203 (N_14203,N_12465,N_12931);
nor U14204 (N_14204,N_12159,N_12673);
or U14205 (N_14205,N_13069,N_12010);
and U14206 (N_14206,N_12978,N_12123);
nand U14207 (N_14207,N_12199,N_12645);
nand U14208 (N_14208,N_12160,N_12892);
or U14209 (N_14209,N_12340,N_12705);
and U14210 (N_14210,N_12947,N_12686);
nor U14211 (N_14211,N_12382,N_13132);
nand U14212 (N_14212,N_12537,N_12344);
or U14213 (N_14213,N_13086,N_12453);
nand U14214 (N_14214,N_12236,N_12146);
and U14215 (N_14215,N_13054,N_12702);
nor U14216 (N_14216,N_12163,N_13258);
nor U14217 (N_14217,N_12333,N_12684);
and U14218 (N_14218,N_13357,N_12812);
and U14219 (N_14219,N_12510,N_12642);
or U14220 (N_14220,N_12638,N_13362);
and U14221 (N_14221,N_12288,N_12844);
and U14222 (N_14222,N_12274,N_12128);
and U14223 (N_14223,N_12054,N_12955);
nor U14224 (N_14224,N_13408,N_13223);
nor U14225 (N_14225,N_12399,N_12960);
or U14226 (N_14226,N_13150,N_13374);
and U14227 (N_14227,N_12457,N_12442);
and U14228 (N_14228,N_12830,N_12697);
or U14229 (N_14229,N_13402,N_12440);
and U14230 (N_14230,N_12226,N_12439);
or U14231 (N_14231,N_13143,N_13257);
or U14232 (N_14232,N_12472,N_12073);
and U14233 (N_14233,N_13307,N_13415);
or U14234 (N_14234,N_13228,N_12400);
nand U14235 (N_14235,N_12154,N_13138);
nor U14236 (N_14236,N_12652,N_12939);
or U14237 (N_14237,N_13433,N_13247);
nor U14238 (N_14238,N_12017,N_12886);
and U14239 (N_14239,N_12836,N_12474);
or U14240 (N_14240,N_12863,N_12357);
and U14241 (N_14241,N_12846,N_12057);
nor U14242 (N_14242,N_13367,N_13497);
or U14243 (N_14243,N_13008,N_12837);
nand U14244 (N_14244,N_12059,N_13310);
or U14245 (N_14245,N_12617,N_12232);
nand U14246 (N_14246,N_13119,N_12101);
or U14247 (N_14247,N_12687,N_13248);
nor U14248 (N_14248,N_12938,N_12052);
nor U14249 (N_14249,N_13297,N_13123);
and U14250 (N_14250,N_13017,N_12484);
nor U14251 (N_14251,N_13091,N_12845);
nand U14252 (N_14252,N_12139,N_12466);
and U14253 (N_14253,N_13218,N_13481);
and U14254 (N_14254,N_12256,N_13493);
nand U14255 (N_14255,N_12091,N_13295);
or U14256 (N_14256,N_12843,N_12231);
or U14257 (N_14257,N_12001,N_12407);
nand U14258 (N_14258,N_12410,N_12235);
nand U14259 (N_14259,N_12273,N_13360);
nor U14260 (N_14260,N_12857,N_12812);
nand U14261 (N_14261,N_12843,N_12174);
or U14262 (N_14262,N_12575,N_12912);
or U14263 (N_14263,N_12577,N_12482);
nand U14264 (N_14264,N_13026,N_13086);
nor U14265 (N_14265,N_12503,N_12542);
nand U14266 (N_14266,N_13469,N_12667);
or U14267 (N_14267,N_12665,N_12086);
and U14268 (N_14268,N_13126,N_12146);
nand U14269 (N_14269,N_12020,N_13346);
and U14270 (N_14270,N_13063,N_12498);
and U14271 (N_14271,N_13391,N_12902);
or U14272 (N_14272,N_12821,N_13058);
nand U14273 (N_14273,N_12781,N_13397);
nand U14274 (N_14274,N_12661,N_12392);
or U14275 (N_14275,N_13223,N_12064);
nand U14276 (N_14276,N_12947,N_12195);
and U14277 (N_14277,N_13444,N_13352);
nand U14278 (N_14278,N_12240,N_12650);
nand U14279 (N_14279,N_12607,N_13032);
or U14280 (N_14280,N_12600,N_13355);
and U14281 (N_14281,N_12152,N_12849);
nand U14282 (N_14282,N_12296,N_12401);
or U14283 (N_14283,N_12517,N_12664);
xor U14284 (N_14284,N_12079,N_13258);
nand U14285 (N_14285,N_12041,N_13001);
or U14286 (N_14286,N_12174,N_12665);
nor U14287 (N_14287,N_13472,N_12547);
or U14288 (N_14288,N_13155,N_13369);
or U14289 (N_14289,N_12010,N_12722);
nor U14290 (N_14290,N_12147,N_12089);
or U14291 (N_14291,N_12652,N_12947);
and U14292 (N_14292,N_12940,N_12619);
nand U14293 (N_14293,N_12417,N_12957);
and U14294 (N_14294,N_12662,N_13041);
nand U14295 (N_14295,N_13047,N_12790);
nand U14296 (N_14296,N_12478,N_13050);
nor U14297 (N_14297,N_13021,N_12684);
and U14298 (N_14298,N_12212,N_12676);
or U14299 (N_14299,N_12893,N_12663);
xnor U14300 (N_14300,N_12103,N_13330);
nand U14301 (N_14301,N_12770,N_12530);
nor U14302 (N_14302,N_13083,N_12060);
or U14303 (N_14303,N_12007,N_12457);
xor U14304 (N_14304,N_12688,N_13182);
nand U14305 (N_14305,N_13420,N_13403);
nor U14306 (N_14306,N_13187,N_12992);
nor U14307 (N_14307,N_12886,N_12372);
nand U14308 (N_14308,N_12499,N_12560);
nor U14309 (N_14309,N_12464,N_12380);
or U14310 (N_14310,N_12531,N_12562);
nand U14311 (N_14311,N_12878,N_13177);
nand U14312 (N_14312,N_12102,N_12957);
xnor U14313 (N_14313,N_12307,N_12362);
nand U14314 (N_14314,N_12004,N_12283);
or U14315 (N_14315,N_12101,N_12756);
nand U14316 (N_14316,N_12408,N_12021);
or U14317 (N_14317,N_12895,N_12026);
nor U14318 (N_14318,N_12569,N_12571);
and U14319 (N_14319,N_13033,N_13462);
nand U14320 (N_14320,N_12707,N_13224);
nor U14321 (N_14321,N_12949,N_13206);
and U14322 (N_14322,N_12947,N_12570);
nand U14323 (N_14323,N_12739,N_12205);
and U14324 (N_14324,N_12348,N_13046);
nand U14325 (N_14325,N_13010,N_12573);
nand U14326 (N_14326,N_12292,N_13146);
and U14327 (N_14327,N_12297,N_12819);
nand U14328 (N_14328,N_12551,N_12243);
or U14329 (N_14329,N_12244,N_13495);
or U14330 (N_14330,N_12399,N_12970);
nand U14331 (N_14331,N_13209,N_13405);
and U14332 (N_14332,N_12079,N_12930);
nor U14333 (N_14333,N_12720,N_12026);
and U14334 (N_14334,N_12945,N_12572);
and U14335 (N_14335,N_12227,N_12398);
or U14336 (N_14336,N_12279,N_13309);
and U14337 (N_14337,N_12389,N_13229);
nor U14338 (N_14338,N_12110,N_13409);
nor U14339 (N_14339,N_12331,N_12430);
nand U14340 (N_14340,N_12845,N_13193);
or U14341 (N_14341,N_12112,N_12732);
nor U14342 (N_14342,N_12324,N_13100);
or U14343 (N_14343,N_12331,N_12247);
nor U14344 (N_14344,N_12149,N_13317);
and U14345 (N_14345,N_12786,N_12963);
and U14346 (N_14346,N_12204,N_12700);
and U14347 (N_14347,N_12244,N_12998);
nor U14348 (N_14348,N_12097,N_12308);
or U14349 (N_14349,N_12211,N_13314);
or U14350 (N_14350,N_12375,N_12837);
or U14351 (N_14351,N_12670,N_12036);
and U14352 (N_14352,N_13047,N_12199);
nor U14353 (N_14353,N_12688,N_12651);
and U14354 (N_14354,N_12682,N_13192);
nand U14355 (N_14355,N_12929,N_13406);
nor U14356 (N_14356,N_12915,N_12696);
or U14357 (N_14357,N_12494,N_13086);
nor U14358 (N_14358,N_13072,N_12650);
and U14359 (N_14359,N_12520,N_12183);
or U14360 (N_14360,N_12861,N_12964);
or U14361 (N_14361,N_13411,N_12678);
and U14362 (N_14362,N_12347,N_12224);
or U14363 (N_14363,N_13383,N_12013);
nand U14364 (N_14364,N_13488,N_12843);
or U14365 (N_14365,N_13448,N_12648);
nand U14366 (N_14366,N_12358,N_13151);
nor U14367 (N_14367,N_12217,N_12702);
and U14368 (N_14368,N_12244,N_12561);
nor U14369 (N_14369,N_12824,N_12527);
or U14370 (N_14370,N_12551,N_12536);
and U14371 (N_14371,N_13292,N_13259);
xor U14372 (N_14372,N_12839,N_13436);
and U14373 (N_14373,N_12028,N_12915);
nor U14374 (N_14374,N_13456,N_12724);
nand U14375 (N_14375,N_13426,N_12382);
nand U14376 (N_14376,N_12208,N_12424);
nand U14377 (N_14377,N_13194,N_12730);
and U14378 (N_14378,N_12012,N_13360);
nand U14379 (N_14379,N_12662,N_12537);
and U14380 (N_14380,N_13014,N_12712);
and U14381 (N_14381,N_13317,N_12489);
xnor U14382 (N_14382,N_12839,N_12828);
nor U14383 (N_14383,N_13114,N_12747);
nor U14384 (N_14384,N_12902,N_12842);
or U14385 (N_14385,N_13389,N_12179);
xor U14386 (N_14386,N_13155,N_13147);
and U14387 (N_14387,N_12996,N_13130);
nor U14388 (N_14388,N_13467,N_12587);
and U14389 (N_14389,N_12207,N_12564);
nor U14390 (N_14390,N_12395,N_12877);
nand U14391 (N_14391,N_13495,N_13014);
or U14392 (N_14392,N_13073,N_12607);
nor U14393 (N_14393,N_12001,N_13213);
or U14394 (N_14394,N_12971,N_12167);
and U14395 (N_14395,N_12461,N_12632);
nor U14396 (N_14396,N_13010,N_13069);
and U14397 (N_14397,N_12916,N_13363);
and U14398 (N_14398,N_12862,N_13062);
or U14399 (N_14399,N_12960,N_12774);
nand U14400 (N_14400,N_12436,N_13248);
nand U14401 (N_14401,N_12314,N_13283);
nand U14402 (N_14402,N_12157,N_13357);
or U14403 (N_14403,N_12205,N_12727);
nand U14404 (N_14404,N_12073,N_12654);
or U14405 (N_14405,N_13302,N_13259);
or U14406 (N_14406,N_13197,N_12651);
or U14407 (N_14407,N_12064,N_12116);
nand U14408 (N_14408,N_12062,N_13350);
nor U14409 (N_14409,N_12641,N_12949);
and U14410 (N_14410,N_13006,N_12787);
and U14411 (N_14411,N_12745,N_12453);
or U14412 (N_14412,N_12227,N_13214);
and U14413 (N_14413,N_13480,N_13279);
and U14414 (N_14414,N_13093,N_13461);
and U14415 (N_14415,N_12672,N_13425);
or U14416 (N_14416,N_12683,N_13259);
nor U14417 (N_14417,N_12903,N_13016);
nand U14418 (N_14418,N_12209,N_13320);
or U14419 (N_14419,N_12348,N_12814);
nor U14420 (N_14420,N_13473,N_13028);
and U14421 (N_14421,N_12993,N_12409);
or U14422 (N_14422,N_12591,N_12231);
or U14423 (N_14423,N_12099,N_12098);
nand U14424 (N_14424,N_12888,N_12446);
or U14425 (N_14425,N_13140,N_12962);
and U14426 (N_14426,N_12448,N_12712);
nand U14427 (N_14427,N_12207,N_13156);
nor U14428 (N_14428,N_13269,N_12965);
nor U14429 (N_14429,N_12334,N_12881);
nand U14430 (N_14430,N_13051,N_13128);
and U14431 (N_14431,N_12406,N_12419);
nor U14432 (N_14432,N_12908,N_12557);
nand U14433 (N_14433,N_13038,N_12100);
and U14434 (N_14434,N_12874,N_12926);
nor U14435 (N_14435,N_12722,N_12243);
nor U14436 (N_14436,N_13456,N_13286);
or U14437 (N_14437,N_12667,N_12409);
and U14438 (N_14438,N_12346,N_12283);
nor U14439 (N_14439,N_12766,N_13395);
and U14440 (N_14440,N_12718,N_12084);
and U14441 (N_14441,N_13365,N_12626);
or U14442 (N_14442,N_12141,N_12040);
and U14443 (N_14443,N_13164,N_12997);
or U14444 (N_14444,N_12651,N_12149);
xnor U14445 (N_14445,N_12389,N_13242);
nor U14446 (N_14446,N_13188,N_13001);
and U14447 (N_14447,N_13016,N_12480);
nor U14448 (N_14448,N_12269,N_13426);
nor U14449 (N_14449,N_12042,N_12408);
or U14450 (N_14450,N_13478,N_13278);
nand U14451 (N_14451,N_12451,N_12849);
or U14452 (N_14452,N_13445,N_13284);
and U14453 (N_14453,N_12466,N_12486);
nor U14454 (N_14454,N_12139,N_12563);
and U14455 (N_14455,N_12631,N_12643);
or U14456 (N_14456,N_12145,N_12399);
nor U14457 (N_14457,N_12740,N_12292);
xnor U14458 (N_14458,N_12856,N_12300);
nor U14459 (N_14459,N_13218,N_12552);
nor U14460 (N_14460,N_13291,N_13104);
nand U14461 (N_14461,N_13207,N_12070);
and U14462 (N_14462,N_13015,N_12970);
or U14463 (N_14463,N_12111,N_12022);
nor U14464 (N_14464,N_12200,N_13158);
nand U14465 (N_14465,N_13452,N_13092);
and U14466 (N_14466,N_12991,N_13351);
nand U14467 (N_14467,N_12062,N_12026);
nand U14468 (N_14468,N_12375,N_12111);
or U14469 (N_14469,N_12056,N_12864);
and U14470 (N_14470,N_12850,N_12088);
nand U14471 (N_14471,N_12765,N_13079);
nand U14472 (N_14472,N_12275,N_12544);
nor U14473 (N_14473,N_12656,N_12694);
xor U14474 (N_14474,N_13201,N_12942);
nand U14475 (N_14475,N_13206,N_12019);
nand U14476 (N_14476,N_12933,N_12279);
nor U14477 (N_14477,N_12185,N_12555);
nand U14478 (N_14478,N_12393,N_12180);
nor U14479 (N_14479,N_12128,N_12937);
or U14480 (N_14480,N_12751,N_12853);
and U14481 (N_14481,N_12522,N_12813);
and U14482 (N_14482,N_12146,N_13253);
nand U14483 (N_14483,N_12258,N_13043);
and U14484 (N_14484,N_12121,N_12145);
nand U14485 (N_14485,N_13422,N_13171);
nand U14486 (N_14486,N_13319,N_12943);
nor U14487 (N_14487,N_13057,N_12934);
or U14488 (N_14488,N_12898,N_12841);
or U14489 (N_14489,N_13380,N_12281);
nand U14490 (N_14490,N_12499,N_12783);
and U14491 (N_14491,N_13119,N_12805);
and U14492 (N_14492,N_13399,N_12855);
and U14493 (N_14493,N_12466,N_13022);
and U14494 (N_14494,N_13271,N_12178);
nand U14495 (N_14495,N_12309,N_13384);
or U14496 (N_14496,N_12183,N_12612);
nand U14497 (N_14497,N_12315,N_13226);
or U14498 (N_14498,N_12878,N_12316);
nand U14499 (N_14499,N_13349,N_12337);
nand U14500 (N_14500,N_12169,N_12045);
and U14501 (N_14501,N_13416,N_12197);
and U14502 (N_14502,N_13465,N_12185);
nand U14503 (N_14503,N_12758,N_12807);
and U14504 (N_14504,N_12563,N_12176);
nand U14505 (N_14505,N_12206,N_12281);
nor U14506 (N_14506,N_12718,N_12358);
nor U14507 (N_14507,N_12788,N_13110);
or U14508 (N_14508,N_12424,N_12640);
nor U14509 (N_14509,N_12486,N_13244);
and U14510 (N_14510,N_12027,N_12001);
nor U14511 (N_14511,N_12763,N_12484);
nand U14512 (N_14512,N_12691,N_12972);
nor U14513 (N_14513,N_12281,N_12580);
or U14514 (N_14514,N_13364,N_13238);
nand U14515 (N_14515,N_12723,N_12024);
and U14516 (N_14516,N_13050,N_12291);
nand U14517 (N_14517,N_13050,N_12465);
nand U14518 (N_14518,N_13432,N_12824);
and U14519 (N_14519,N_12838,N_12729);
nor U14520 (N_14520,N_12905,N_13365);
and U14521 (N_14521,N_12139,N_12686);
nor U14522 (N_14522,N_12436,N_13469);
and U14523 (N_14523,N_12944,N_13287);
nand U14524 (N_14524,N_13462,N_13343);
nand U14525 (N_14525,N_12266,N_12374);
or U14526 (N_14526,N_12648,N_12336);
nor U14527 (N_14527,N_13035,N_12781);
nor U14528 (N_14528,N_12900,N_13496);
and U14529 (N_14529,N_12674,N_12178);
nor U14530 (N_14530,N_13018,N_12995);
nand U14531 (N_14531,N_12768,N_13139);
nand U14532 (N_14532,N_13310,N_12079);
and U14533 (N_14533,N_12008,N_12504);
nor U14534 (N_14534,N_12376,N_13038);
nand U14535 (N_14535,N_12191,N_13273);
nor U14536 (N_14536,N_12744,N_13104);
nand U14537 (N_14537,N_12064,N_13095);
nand U14538 (N_14538,N_12383,N_12691);
or U14539 (N_14539,N_12015,N_13452);
nor U14540 (N_14540,N_12533,N_13376);
nor U14541 (N_14541,N_13429,N_13143);
and U14542 (N_14542,N_12982,N_12022);
nor U14543 (N_14543,N_12436,N_13353);
and U14544 (N_14544,N_12893,N_12110);
and U14545 (N_14545,N_13071,N_12257);
nor U14546 (N_14546,N_12376,N_12578);
and U14547 (N_14547,N_13083,N_12194);
or U14548 (N_14548,N_12119,N_12892);
nand U14549 (N_14549,N_12956,N_12726);
or U14550 (N_14550,N_12885,N_13082);
nand U14551 (N_14551,N_12169,N_12717);
or U14552 (N_14552,N_13243,N_13059);
and U14553 (N_14553,N_12604,N_12749);
nand U14554 (N_14554,N_12485,N_12705);
and U14555 (N_14555,N_13028,N_12529);
or U14556 (N_14556,N_12837,N_13130);
nor U14557 (N_14557,N_12264,N_12839);
nand U14558 (N_14558,N_12741,N_12497);
or U14559 (N_14559,N_12070,N_12693);
and U14560 (N_14560,N_12470,N_12126);
nor U14561 (N_14561,N_12423,N_12061);
nand U14562 (N_14562,N_12033,N_12625);
and U14563 (N_14563,N_13165,N_12676);
or U14564 (N_14564,N_13341,N_12153);
nor U14565 (N_14565,N_12182,N_12412);
or U14566 (N_14566,N_13365,N_12732);
or U14567 (N_14567,N_13338,N_12792);
nand U14568 (N_14568,N_12521,N_13145);
and U14569 (N_14569,N_12002,N_13209);
nand U14570 (N_14570,N_13168,N_12797);
nor U14571 (N_14571,N_12810,N_12476);
nand U14572 (N_14572,N_12267,N_12036);
or U14573 (N_14573,N_12231,N_13061);
nor U14574 (N_14574,N_12074,N_12854);
or U14575 (N_14575,N_12144,N_12380);
nand U14576 (N_14576,N_13348,N_13038);
nand U14577 (N_14577,N_12644,N_13226);
nand U14578 (N_14578,N_12791,N_13272);
or U14579 (N_14579,N_13044,N_12721);
nand U14580 (N_14580,N_13323,N_12888);
or U14581 (N_14581,N_13118,N_13487);
or U14582 (N_14582,N_12330,N_13474);
nand U14583 (N_14583,N_12421,N_13355);
nor U14584 (N_14584,N_13048,N_12009);
and U14585 (N_14585,N_12679,N_12089);
and U14586 (N_14586,N_13002,N_13068);
nor U14587 (N_14587,N_12571,N_12697);
nand U14588 (N_14588,N_12225,N_12409);
nand U14589 (N_14589,N_12363,N_12758);
nand U14590 (N_14590,N_13283,N_12037);
nand U14591 (N_14591,N_13389,N_12431);
nor U14592 (N_14592,N_12622,N_13100);
nor U14593 (N_14593,N_13447,N_12802);
and U14594 (N_14594,N_12736,N_12788);
nor U14595 (N_14595,N_12594,N_13268);
nand U14596 (N_14596,N_13226,N_12872);
nand U14597 (N_14597,N_13012,N_13479);
or U14598 (N_14598,N_13276,N_12388);
nand U14599 (N_14599,N_13152,N_13241);
nor U14600 (N_14600,N_13240,N_12352);
and U14601 (N_14601,N_12449,N_12054);
or U14602 (N_14602,N_12061,N_12107);
or U14603 (N_14603,N_12336,N_13381);
or U14604 (N_14604,N_12701,N_12463);
or U14605 (N_14605,N_12206,N_12726);
and U14606 (N_14606,N_13299,N_13492);
nand U14607 (N_14607,N_13454,N_12013);
nand U14608 (N_14608,N_12541,N_13405);
nor U14609 (N_14609,N_12108,N_12019);
and U14610 (N_14610,N_12275,N_12490);
nand U14611 (N_14611,N_12348,N_12464);
xnor U14612 (N_14612,N_13485,N_13474);
nor U14613 (N_14613,N_12965,N_12302);
and U14614 (N_14614,N_13012,N_13407);
nor U14615 (N_14615,N_12648,N_12428);
nand U14616 (N_14616,N_13004,N_12143);
and U14617 (N_14617,N_12604,N_12168);
or U14618 (N_14618,N_13069,N_13040);
or U14619 (N_14619,N_12320,N_13483);
or U14620 (N_14620,N_13396,N_13349);
nor U14621 (N_14621,N_12477,N_12059);
and U14622 (N_14622,N_12922,N_12919);
nor U14623 (N_14623,N_12904,N_13123);
or U14624 (N_14624,N_12624,N_12877);
nor U14625 (N_14625,N_12291,N_13072);
nor U14626 (N_14626,N_12856,N_12581);
and U14627 (N_14627,N_13376,N_12413);
and U14628 (N_14628,N_13329,N_12916);
nand U14629 (N_14629,N_12213,N_13100);
nand U14630 (N_14630,N_12134,N_13040);
or U14631 (N_14631,N_13315,N_12893);
or U14632 (N_14632,N_12045,N_13068);
or U14633 (N_14633,N_12939,N_13072);
or U14634 (N_14634,N_12388,N_12485);
nor U14635 (N_14635,N_13238,N_12219);
or U14636 (N_14636,N_12418,N_12810);
or U14637 (N_14637,N_12105,N_13080);
and U14638 (N_14638,N_12354,N_12054);
or U14639 (N_14639,N_12990,N_12043);
and U14640 (N_14640,N_12697,N_12444);
or U14641 (N_14641,N_12672,N_13098);
or U14642 (N_14642,N_12087,N_12932);
nand U14643 (N_14643,N_12438,N_13159);
nor U14644 (N_14644,N_12685,N_12471);
nor U14645 (N_14645,N_12948,N_12745);
or U14646 (N_14646,N_12463,N_13078);
or U14647 (N_14647,N_13140,N_13201);
or U14648 (N_14648,N_12487,N_12818);
and U14649 (N_14649,N_13178,N_12872);
nor U14650 (N_14650,N_12979,N_12486);
or U14651 (N_14651,N_12671,N_12541);
nor U14652 (N_14652,N_13314,N_12077);
or U14653 (N_14653,N_13360,N_12901);
nand U14654 (N_14654,N_13313,N_12877);
or U14655 (N_14655,N_12358,N_13191);
nor U14656 (N_14656,N_12303,N_13217);
or U14657 (N_14657,N_13062,N_12050);
or U14658 (N_14658,N_12969,N_12534);
nand U14659 (N_14659,N_12515,N_12959);
and U14660 (N_14660,N_12523,N_13141);
nand U14661 (N_14661,N_12590,N_12721);
nand U14662 (N_14662,N_12595,N_13076);
or U14663 (N_14663,N_12377,N_12978);
and U14664 (N_14664,N_12618,N_13190);
nor U14665 (N_14665,N_12512,N_12492);
nand U14666 (N_14666,N_12700,N_12899);
or U14667 (N_14667,N_12663,N_12869);
nor U14668 (N_14668,N_12025,N_13378);
nand U14669 (N_14669,N_12581,N_13235);
and U14670 (N_14670,N_12441,N_12724);
nor U14671 (N_14671,N_12856,N_12909);
nand U14672 (N_14672,N_12333,N_12867);
nor U14673 (N_14673,N_12153,N_12787);
nand U14674 (N_14674,N_13448,N_12888);
and U14675 (N_14675,N_12929,N_12643);
or U14676 (N_14676,N_13461,N_12102);
nor U14677 (N_14677,N_12323,N_13038);
nand U14678 (N_14678,N_12781,N_12412);
and U14679 (N_14679,N_12423,N_12273);
nand U14680 (N_14680,N_12095,N_13490);
nor U14681 (N_14681,N_13333,N_13301);
and U14682 (N_14682,N_13183,N_13387);
nand U14683 (N_14683,N_12595,N_12100);
and U14684 (N_14684,N_12297,N_12606);
or U14685 (N_14685,N_13263,N_12932);
or U14686 (N_14686,N_12862,N_12213);
or U14687 (N_14687,N_12900,N_13065);
nand U14688 (N_14688,N_13000,N_12535);
and U14689 (N_14689,N_12184,N_12537);
and U14690 (N_14690,N_12433,N_13022);
and U14691 (N_14691,N_12326,N_13117);
or U14692 (N_14692,N_13463,N_13492);
nor U14693 (N_14693,N_12888,N_12715);
nor U14694 (N_14694,N_12629,N_13335);
and U14695 (N_14695,N_13262,N_13166);
or U14696 (N_14696,N_12695,N_12366);
nor U14697 (N_14697,N_13248,N_12303);
nand U14698 (N_14698,N_12804,N_12026);
or U14699 (N_14699,N_13199,N_12399);
or U14700 (N_14700,N_13105,N_12795);
nor U14701 (N_14701,N_12195,N_13169);
or U14702 (N_14702,N_12426,N_13185);
and U14703 (N_14703,N_12672,N_12510);
nand U14704 (N_14704,N_12609,N_12199);
and U14705 (N_14705,N_12749,N_12410);
and U14706 (N_14706,N_12688,N_12186);
or U14707 (N_14707,N_12001,N_12474);
nor U14708 (N_14708,N_12420,N_12176);
xnor U14709 (N_14709,N_13339,N_13159);
nand U14710 (N_14710,N_12230,N_12173);
or U14711 (N_14711,N_12487,N_12237);
and U14712 (N_14712,N_12686,N_12725);
nor U14713 (N_14713,N_13117,N_12734);
nand U14714 (N_14714,N_12951,N_13430);
nand U14715 (N_14715,N_12422,N_13315);
nor U14716 (N_14716,N_12572,N_12411);
and U14717 (N_14717,N_13054,N_12697);
nand U14718 (N_14718,N_12316,N_12600);
or U14719 (N_14719,N_13197,N_13143);
or U14720 (N_14720,N_12792,N_12398);
nor U14721 (N_14721,N_12068,N_13267);
and U14722 (N_14722,N_13036,N_13258);
nor U14723 (N_14723,N_12437,N_12080);
nand U14724 (N_14724,N_12285,N_13477);
nor U14725 (N_14725,N_13287,N_12293);
or U14726 (N_14726,N_12261,N_12503);
and U14727 (N_14727,N_12087,N_12011);
and U14728 (N_14728,N_13162,N_12564);
nand U14729 (N_14729,N_13194,N_12914);
and U14730 (N_14730,N_12841,N_12998);
nor U14731 (N_14731,N_12448,N_12857);
and U14732 (N_14732,N_12287,N_13397);
and U14733 (N_14733,N_12802,N_13363);
or U14734 (N_14734,N_13318,N_12838);
nor U14735 (N_14735,N_12687,N_13345);
and U14736 (N_14736,N_12838,N_12582);
or U14737 (N_14737,N_12240,N_12119);
or U14738 (N_14738,N_12874,N_12747);
nand U14739 (N_14739,N_12129,N_12385);
and U14740 (N_14740,N_12009,N_12858);
or U14741 (N_14741,N_12133,N_13358);
and U14742 (N_14742,N_13482,N_12165);
and U14743 (N_14743,N_12123,N_12072);
and U14744 (N_14744,N_12428,N_12459);
nand U14745 (N_14745,N_13152,N_12377);
nor U14746 (N_14746,N_12418,N_12351);
nand U14747 (N_14747,N_13127,N_12231);
nand U14748 (N_14748,N_13011,N_12122);
or U14749 (N_14749,N_13107,N_12149);
nand U14750 (N_14750,N_12048,N_13387);
and U14751 (N_14751,N_12150,N_12601);
and U14752 (N_14752,N_13453,N_12963);
or U14753 (N_14753,N_13371,N_12032);
or U14754 (N_14754,N_12671,N_13286);
nand U14755 (N_14755,N_12564,N_12602);
nor U14756 (N_14756,N_13305,N_12057);
and U14757 (N_14757,N_12402,N_12364);
and U14758 (N_14758,N_12204,N_13428);
nor U14759 (N_14759,N_12338,N_13158);
nand U14760 (N_14760,N_12990,N_12258);
and U14761 (N_14761,N_12911,N_12254);
or U14762 (N_14762,N_12235,N_12299);
or U14763 (N_14763,N_12639,N_13112);
nand U14764 (N_14764,N_12880,N_12144);
and U14765 (N_14765,N_12655,N_12332);
or U14766 (N_14766,N_13304,N_12486);
nor U14767 (N_14767,N_13167,N_12813);
or U14768 (N_14768,N_12776,N_13280);
or U14769 (N_14769,N_12475,N_12287);
or U14770 (N_14770,N_12466,N_13402);
nand U14771 (N_14771,N_12355,N_12839);
nand U14772 (N_14772,N_12456,N_12880);
nor U14773 (N_14773,N_13247,N_13454);
nor U14774 (N_14774,N_13179,N_12188);
nor U14775 (N_14775,N_12595,N_12720);
and U14776 (N_14776,N_12922,N_12270);
and U14777 (N_14777,N_13390,N_12196);
and U14778 (N_14778,N_13006,N_12093);
or U14779 (N_14779,N_12735,N_12620);
nor U14780 (N_14780,N_12104,N_13492);
and U14781 (N_14781,N_12283,N_12010);
nand U14782 (N_14782,N_12323,N_12197);
or U14783 (N_14783,N_12938,N_12831);
and U14784 (N_14784,N_13276,N_12066);
and U14785 (N_14785,N_13074,N_13381);
or U14786 (N_14786,N_12773,N_12410);
or U14787 (N_14787,N_13012,N_12922);
or U14788 (N_14788,N_12419,N_12801);
nand U14789 (N_14789,N_13063,N_12262);
nor U14790 (N_14790,N_12925,N_12591);
nor U14791 (N_14791,N_12346,N_12781);
nor U14792 (N_14792,N_12146,N_12083);
nor U14793 (N_14793,N_12091,N_13272);
and U14794 (N_14794,N_12619,N_12997);
or U14795 (N_14795,N_13136,N_12077);
and U14796 (N_14796,N_13232,N_12723);
or U14797 (N_14797,N_13018,N_12622);
nor U14798 (N_14798,N_13444,N_12576);
and U14799 (N_14799,N_13310,N_12447);
and U14800 (N_14800,N_13396,N_12989);
nand U14801 (N_14801,N_12945,N_13491);
nor U14802 (N_14802,N_12825,N_13357);
or U14803 (N_14803,N_13291,N_13393);
nor U14804 (N_14804,N_12098,N_12008);
or U14805 (N_14805,N_12205,N_12489);
and U14806 (N_14806,N_12760,N_13425);
nor U14807 (N_14807,N_12600,N_13326);
nor U14808 (N_14808,N_12880,N_13032);
or U14809 (N_14809,N_13030,N_13119);
nand U14810 (N_14810,N_12177,N_12184);
nor U14811 (N_14811,N_13145,N_12981);
and U14812 (N_14812,N_13011,N_12461);
and U14813 (N_14813,N_13301,N_12337);
and U14814 (N_14814,N_12886,N_12921);
and U14815 (N_14815,N_12103,N_12525);
nand U14816 (N_14816,N_12869,N_12073);
nor U14817 (N_14817,N_13266,N_12487);
nor U14818 (N_14818,N_12588,N_12614);
nor U14819 (N_14819,N_13033,N_12365);
or U14820 (N_14820,N_12845,N_12138);
nand U14821 (N_14821,N_12597,N_13097);
nand U14822 (N_14822,N_12306,N_12873);
or U14823 (N_14823,N_13221,N_13248);
nor U14824 (N_14824,N_12419,N_13247);
and U14825 (N_14825,N_13279,N_12312);
nand U14826 (N_14826,N_12743,N_12289);
nor U14827 (N_14827,N_13283,N_13012);
nand U14828 (N_14828,N_13258,N_12177);
xnor U14829 (N_14829,N_12000,N_12299);
nor U14830 (N_14830,N_12305,N_12396);
nand U14831 (N_14831,N_13345,N_12794);
nand U14832 (N_14832,N_12029,N_12811);
or U14833 (N_14833,N_12154,N_12194);
or U14834 (N_14834,N_12487,N_12527);
and U14835 (N_14835,N_12722,N_12107);
nand U14836 (N_14836,N_12692,N_13495);
nor U14837 (N_14837,N_13418,N_12275);
nand U14838 (N_14838,N_12975,N_12114);
or U14839 (N_14839,N_12503,N_12124);
nand U14840 (N_14840,N_12102,N_13207);
or U14841 (N_14841,N_12953,N_12411);
or U14842 (N_14842,N_12244,N_12331);
xnor U14843 (N_14843,N_13387,N_12429);
and U14844 (N_14844,N_13373,N_13467);
nor U14845 (N_14845,N_12089,N_13404);
nor U14846 (N_14846,N_13325,N_13250);
or U14847 (N_14847,N_12047,N_13233);
or U14848 (N_14848,N_12948,N_13125);
nor U14849 (N_14849,N_13141,N_13022);
nor U14850 (N_14850,N_13461,N_12836);
nand U14851 (N_14851,N_13085,N_13158);
and U14852 (N_14852,N_12797,N_13146);
nor U14853 (N_14853,N_13309,N_12651);
nor U14854 (N_14854,N_12961,N_13404);
xnor U14855 (N_14855,N_12601,N_12096);
nand U14856 (N_14856,N_13241,N_12272);
or U14857 (N_14857,N_13110,N_12941);
nor U14858 (N_14858,N_13189,N_12644);
and U14859 (N_14859,N_12712,N_12922);
nand U14860 (N_14860,N_12475,N_12932);
nor U14861 (N_14861,N_12411,N_12442);
nor U14862 (N_14862,N_12114,N_12710);
nand U14863 (N_14863,N_12608,N_12129);
nor U14864 (N_14864,N_12407,N_13298);
and U14865 (N_14865,N_13317,N_13384);
nor U14866 (N_14866,N_13432,N_12893);
and U14867 (N_14867,N_12278,N_13437);
and U14868 (N_14868,N_12450,N_13114);
and U14869 (N_14869,N_12205,N_12552);
or U14870 (N_14870,N_12336,N_13186);
nor U14871 (N_14871,N_12931,N_13258);
nand U14872 (N_14872,N_12127,N_12132);
nor U14873 (N_14873,N_13345,N_13010);
nand U14874 (N_14874,N_12925,N_13003);
nor U14875 (N_14875,N_13046,N_12267);
or U14876 (N_14876,N_12247,N_13200);
or U14877 (N_14877,N_12635,N_13067);
or U14878 (N_14878,N_12641,N_13194);
nand U14879 (N_14879,N_12061,N_12225);
and U14880 (N_14880,N_13287,N_12292);
or U14881 (N_14881,N_12418,N_13264);
or U14882 (N_14882,N_12065,N_12948);
and U14883 (N_14883,N_12494,N_12999);
or U14884 (N_14884,N_12801,N_12207);
nor U14885 (N_14885,N_13477,N_12705);
nand U14886 (N_14886,N_12742,N_12643);
nor U14887 (N_14887,N_12364,N_13434);
or U14888 (N_14888,N_12007,N_13136);
nand U14889 (N_14889,N_12570,N_13222);
nor U14890 (N_14890,N_12488,N_12049);
nor U14891 (N_14891,N_12418,N_13093);
nand U14892 (N_14892,N_13463,N_12801);
nor U14893 (N_14893,N_12104,N_12518);
or U14894 (N_14894,N_13430,N_12838);
nor U14895 (N_14895,N_12128,N_13021);
nor U14896 (N_14896,N_12124,N_12779);
nand U14897 (N_14897,N_13090,N_12640);
or U14898 (N_14898,N_12072,N_12333);
nor U14899 (N_14899,N_12922,N_12355);
and U14900 (N_14900,N_12604,N_12910);
xnor U14901 (N_14901,N_12895,N_12700);
nand U14902 (N_14902,N_12521,N_13085);
or U14903 (N_14903,N_12499,N_12453);
or U14904 (N_14904,N_12154,N_12641);
and U14905 (N_14905,N_13227,N_13454);
nor U14906 (N_14906,N_13041,N_12719);
and U14907 (N_14907,N_13158,N_12366);
nor U14908 (N_14908,N_12033,N_13449);
and U14909 (N_14909,N_12512,N_12084);
nand U14910 (N_14910,N_12405,N_13036);
nand U14911 (N_14911,N_12979,N_12616);
and U14912 (N_14912,N_12962,N_12229);
and U14913 (N_14913,N_12099,N_12038);
nor U14914 (N_14914,N_13011,N_12984);
nor U14915 (N_14915,N_12268,N_13231);
nor U14916 (N_14916,N_12037,N_12277);
nand U14917 (N_14917,N_12859,N_12765);
and U14918 (N_14918,N_12073,N_13129);
or U14919 (N_14919,N_13036,N_12716);
or U14920 (N_14920,N_12131,N_12656);
and U14921 (N_14921,N_12790,N_12157);
nand U14922 (N_14922,N_12286,N_13035);
nand U14923 (N_14923,N_13096,N_12813);
nand U14924 (N_14924,N_12691,N_12771);
or U14925 (N_14925,N_12496,N_12598);
and U14926 (N_14926,N_12648,N_12987);
nand U14927 (N_14927,N_13202,N_12578);
nand U14928 (N_14928,N_13441,N_13366);
or U14929 (N_14929,N_12962,N_13309);
and U14930 (N_14930,N_13133,N_12428);
and U14931 (N_14931,N_13233,N_13499);
nor U14932 (N_14932,N_12400,N_12241);
nor U14933 (N_14933,N_13271,N_13309);
nand U14934 (N_14934,N_12413,N_12173);
and U14935 (N_14935,N_12770,N_12388);
and U14936 (N_14936,N_13330,N_13223);
or U14937 (N_14937,N_13469,N_13258);
or U14938 (N_14938,N_13312,N_12117);
nor U14939 (N_14939,N_12257,N_13188);
or U14940 (N_14940,N_12614,N_13360);
nand U14941 (N_14941,N_13390,N_13155);
nand U14942 (N_14942,N_12045,N_12084);
nand U14943 (N_14943,N_12736,N_13044);
or U14944 (N_14944,N_12196,N_12844);
nor U14945 (N_14945,N_12564,N_12021);
and U14946 (N_14946,N_12944,N_13272);
nor U14947 (N_14947,N_12885,N_13333);
nor U14948 (N_14948,N_12991,N_13193);
and U14949 (N_14949,N_13407,N_12682);
and U14950 (N_14950,N_12064,N_12884);
nor U14951 (N_14951,N_13333,N_12366);
nand U14952 (N_14952,N_12241,N_12779);
or U14953 (N_14953,N_12998,N_12447);
or U14954 (N_14954,N_12371,N_12575);
or U14955 (N_14955,N_12737,N_13017);
nand U14956 (N_14956,N_13468,N_12501);
or U14957 (N_14957,N_13304,N_13188);
or U14958 (N_14958,N_13236,N_13159);
and U14959 (N_14959,N_12296,N_13328);
and U14960 (N_14960,N_12949,N_12538);
nor U14961 (N_14961,N_13206,N_12944);
and U14962 (N_14962,N_12629,N_12402);
and U14963 (N_14963,N_13181,N_13077);
nand U14964 (N_14964,N_13268,N_12260);
nand U14965 (N_14965,N_13036,N_13397);
or U14966 (N_14966,N_12208,N_12371);
nor U14967 (N_14967,N_13024,N_12272);
xor U14968 (N_14968,N_12447,N_13039);
or U14969 (N_14969,N_12537,N_13097);
nor U14970 (N_14970,N_13266,N_12342);
nand U14971 (N_14971,N_12089,N_12456);
or U14972 (N_14972,N_12392,N_12100);
and U14973 (N_14973,N_12147,N_12515);
nand U14974 (N_14974,N_13204,N_13488);
or U14975 (N_14975,N_12911,N_13020);
nand U14976 (N_14976,N_13290,N_12189);
nor U14977 (N_14977,N_12345,N_12676);
or U14978 (N_14978,N_12380,N_13377);
or U14979 (N_14979,N_13163,N_12125);
nand U14980 (N_14980,N_13021,N_12410);
nand U14981 (N_14981,N_13405,N_12432);
nor U14982 (N_14982,N_13435,N_12513);
nor U14983 (N_14983,N_12539,N_12015);
nand U14984 (N_14984,N_12347,N_12262);
and U14985 (N_14985,N_12067,N_12771);
nand U14986 (N_14986,N_12323,N_12021);
and U14987 (N_14987,N_12786,N_12923);
nor U14988 (N_14988,N_12666,N_12503);
nand U14989 (N_14989,N_12605,N_13144);
or U14990 (N_14990,N_12901,N_12559);
nand U14991 (N_14991,N_13387,N_12809);
nor U14992 (N_14992,N_13312,N_13134);
or U14993 (N_14993,N_13297,N_12820);
and U14994 (N_14994,N_12569,N_12924);
or U14995 (N_14995,N_12535,N_12722);
and U14996 (N_14996,N_12004,N_13228);
nand U14997 (N_14997,N_12825,N_13199);
nor U14998 (N_14998,N_12978,N_12111);
and U14999 (N_14999,N_12418,N_13215);
and UO_0 (O_0,N_13572,N_14066);
nor UO_1 (O_1,N_14391,N_13626);
nor UO_2 (O_2,N_14551,N_13919);
nor UO_3 (O_3,N_14029,N_14601);
and UO_4 (O_4,N_13522,N_13765);
or UO_5 (O_5,N_13956,N_13543);
or UO_6 (O_6,N_14536,N_14765);
xor UO_7 (O_7,N_13717,N_14556);
nand UO_8 (O_8,N_14844,N_14670);
or UO_9 (O_9,N_13900,N_14181);
nor UO_10 (O_10,N_13961,N_14374);
nand UO_11 (O_11,N_13716,N_14015);
nor UO_12 (O_12,N_14101,N_14806);
nand UO_13 (O_13,N_13944,N_14998);
or UO_14 (O_14,N_13506,N_14183);
and UO_15 (O_15,N_14873,N_13786);
or UO_16 (O_16,N_13503,N_13530);
nand UO_17 (O_17,N_14744,N_14853);
or UO_18 (O_18,N_14741,N_14582);
nand UO_19 (O_19,N_13945,N_13697);
nand UO_20 (O_20,N_13650,N_14353);
and UO_21 (O_21,N_13865,N_14386);
nand UO_22 (O_22,N_14552,N_14492);
nand UO_23 (O_23,N_13646,N_13728);
or UO_24 (O_24,N_13953,N_14487);
xnor UO_25 (O_25,N_13709,N_13850);
nor UO_26 (O_26,N_14159,N_13782);
and UO_27 (O_27,N_14784,N_14919);
or UO_28 (O_28,N_14977,N_14686);
nor UO_29 (O_29,N_13653,N_14795);
and UO_30 (O_30,N_13556,N_13502);
or UO_31 (O_31,N_13525,N_13630);
and UO_32 (O_32,N_14688,N_14389);
nor UO_33 (O_33,N_14093,N_14849);
nand UO_34 (O_34,N_14877,N_13742);
or UO_35 (O_35,N_14063,N_13802);
and UO_36 (O_36,N_13749,N_14016);
or UO_37 (O_37,N_13715,N_13514);
nand UO_38 (O_38,N_13739,N_13960);
nor UO_39 (O_39,N_14893,N_14489);
or UO_40 (O_40,N_14398,N_13969);
nor UO_41 (O_41,N_14141,N_14572);
or UO_42 (O_42,N_14148,N_13567);
or UO_43 (O_43,N_13753,N_14336);
or UO_44 (O_44,N_14171,N_14416);
nor UO_45 (O_45,N_13970,N_14982);
and UO_46 (O_46,N_14925,N_14023);
nor UO_47 (O_47,N_13771,N_13901);
nand UO_48 (O_48,N_13624,N_14476);
and UO_49 (O_49,N_13760,N_13821);
or UO_50 (O_50,N_14668,N_14026);
and UO_51 (O_51,N_14583,N_14772);
nand UO_52 (O_52,N_13833,N_14960);
nand UO_53 (O_53,N_14862,N_13776);
or UO_54 (O_54,N_13822,N_14248);
and UO_55 (O_55,N_14285,N_14498);
nand UO_56 (O_56,N_14387,N_14434);
or UO_57 (O_57,N_13762,N_14813);
and UO_58 (O_58,N_14190,N_14576);
or UO_59 (O_59,N_14037,N_14523);
nand UO_60 (O_60,N_14952,N_14515);
or UO_61 (O_61,N_14217,N_14196);
nand UO_62 (O_62,N_13955,N_13857);
nor UO_63 (O_63,N_13580,N_13851);
nand UO_64 (O_64,N_14699,N_14521);
nor UO_65 (O_65,N_13818,N_14033);
nand UO_66 (O_66,N_14007,N_14214);
or UO_67 (O_67,N_14432,N_13596);
or UO_68 (O_68,N_14624,N_14994);
and UO_69 (O_69,N_13702,N_14958);
nand UO_70 (O_70,N_14564,N_13829);
or UO_71 (O_71,N_14155,N_14828);
or UO_72 (O_72,N_14458,N_14511);
or UO_73 (O_73,N_14143,N_14865);
and UO_74 (O_74,N_13923,N_14247);
or UO_75 (O_75,N_13838,N_14036);
nor UO_76 (O_76,N_13814,N_14928);
and UO_77 (O_77,N_13625,N_13873);
or UO_78 (O_78,N_13748,N_13500);
or UO_79 (O_79,N_13768,N_13544);
nand UO_80 (O_80,N_14810,N_13531);
xor UO_81 (O_81,N_14628,N_14149);
and UO_82 (O_82,N_13523,N_13659);
nor UO_83 (O_83,N_14393,N_14533);
nor UO_84 (O_84,N_14461,N_14917);
nand UO_85 (O_85,N_14038,N_14139);
nor UO_86 (O_86,N_13517,N_13971);
or UO_87 (O_87,N_14047,N_14030);
or UO_88 (O_88,N_14068,N_14943);
and UO_89 (O_89,N_14537,N_13591);
nand UO_90 (O_90,N_14570,N_14832);
nand UO_91 (O_91,N_13640,N_14395);
and UO_92 (O_92,N_13780,N_14463);
nand UO_93 (O_93,N_13685,N_14587);
nor UO_94 (O_94,N_14920,N_14845);
nor UO_95 (O_95,N_14375,N_14403);
and UO_96 (O_96,N_13858,N_13976);
nand UO_97 (O_97,N_13806,N_14292);
nand UO_98 (O_98,N_13555,N_13991);
and UO_99 (O_99,N_14157,N_13869);
nor UO_100 (O_100,N_13711,N_13639);
and UO_101 (O_101,N_14225,N_14579);
or UO_102 (O_102,N_14716,N_14289);
nand UO_103 (O_103,N_14715,N_14158);
nor UO_104 (O_104,N_14619,N_14860);
or UO_105 (O_105,N_14776,N_14745);
or UO_106 (O_106,N_14774,N_14257);
or UO_107 (O_107,N_14867,N_14909);
nor UO_108 (O_108,N_14105,N_14335);
and UO_109 (O_109,N_13550,N_14614);
nand UO_110 (O_110,N_14044,N_14035);
or UO_111 (O_111,N_14805,N_14617);
nand UO_112 (O_112,N_13566,N_14651);
or UO_113 (O_113,N_14456,N_14750);
and UO_114 (O_114,N_14004,N_14114);
nand UO_115 (O_115,N_13589,N_14469);
nand UO_116 (O_116,N_14694,N_13964);
nor UO_117 (O_117,N_13593,N_14242);
or UO_118 (O_118,N_14811,N_14665);
and UO_119 (O_119,N_13670,N_13537);
nand UO_120 (O_120,N_14163,N_14525);
nand UO_121 (O_121,N_14174,N_13852);
or UO_122 (O_122,N_14493,N_13657);
or UO_123 (O_123,N_14124,N_13827);
nor UO_124 (O_124,N_14192,N_14526);
nand UO_125 (O_125,N_13870,N_14550);
nor UO_126 (O_126,N_14755,N_14747);
xnor UO_127 (O_127,N_14791,N_14528);
or UO_128 (O_128,N_14441,N_13518);
or UO_129 (O_129,N_14485,N_13618);
nor UO_130 (O_130,N_14589,N_14334);
and UO_131 (O_131,N_14782,N_13766);
and UO_132 (O_132,N_14527,N_13601);
and UO_133 (O_133,N_13721,N_14201);
nand UO_134 (O_134,N_13884,N_14838);
nand UO_135 (O_135,N_14687,N_14307);
and UO_136 (O_136,N_13545,N_14275);
and UO_137 (O_137,N_14310,N_13823);
and UO_138 (O_138,N_14969,N_14554);
and UO_139 (O_139,N_14679,N_14206);
nand UO_140 (O_140,N_14597,N_13983);
and UO_141 (O_141,N_14126,N_14912);
and UO_142 (O_142,N_14298,N_13908);
xnor UO_143 (O_143,N_14717,N_14540);
and UO_144 (O_144,N_14859,N_13936);
or UO_145 (O_145,N_14112,N_14987);
or UO_146 (O_146,N_14720,N_13787);
nand UO_147 (O_147,N_13773,N_14074);
or UO_148 (O_148,N_14276,N_14459);
and UO_149 (O_149,N_13927,N_13605);
nand UO_150 (O_150,N_14736,N_13967);
and UO_151 (O_151,N_14889,N_14993);
nand UO_152 (O_152,N_14885,N_14645);
or UO_153 (O_153,N_14759,N_14238);
and UO_154 (O_154,N_14955,N_14305);
nand UO_155 (O_155,N_14559,N_14472);
nand UO_156 (O_156,N_14700,N_14881);
nand UO_157 (O_157,N_13904,N_13779);
nand UO_158 (O_158,N_14503,N_14988);
nand UO_159 (O_159,N_14706,N_14359);
nand UO_160 (O_160,N_13541,N_13999);
and UO_161 (O_161,N_14954,N_14253);
nand UO_162 (O_162,N_13575,N_14671);
xnor UO_163 (O_163,N_14083,N_14975);
or UO_164 (O_164,N_13830,N_14421);
nor UO_165 (O_165,N_14075,N_14486);
nand UO_166 (O_166,N_14728,N_14634);
nand UO_167 (O_167,N_13810,N_13651);
nand UO_168 (O_168,N_14496,N_14823);
or UO_169 (O_169,N_13701,N_14259);
nor UO_170 (O_170,N_14172,N_14924);
and UO_171 (O_171,N_14228,N_14731);
nand UO_172 (O_172,N_13563,N_14205);
nor UO_173 (O_173,N_13602,N_13800);
nor UO_174 (O_174,N_13649,N_14470);
nand UO_175 (O_175,N_14945,N_14830);
and UO_176 (O_176,N_13980,N_14479);
and UO_177 (O_177,N_14117,N_13910);
and UO_178 (O_178,N_13939,N_13914);
nand UO_179 (O_179,N_13511,N_13824);
nand UO_180 (O_180,N_14640,N_14581);
nor UO_181 (O_181,N_14048,N_14468);
nand UO_182 (O_182,N_13738,N_13707);
nor UO_183 (O_183,N_14641,N_14786);
nor UO_184 (O_184,N_13747,N_13557);
or UO_185 (O_185,N_13791,N_14133);
or UO_186 (O_186,N_14709,N_13801);
nor UO_187 (O_187,N_14032,N_13615);
nor UO_188 (O_188,N_13941,N_13859);
or UO_189 (O_189,N_13671,N_13770);
nand UO_190 (O_190,N_14146,N_14367);
nand UO_191 (O_191,N_14145,N_13688);
nand UO_192 (O_192,N_13636,N_14095);
nand UO_193 (O_193,N_14968,N_14907);
nand UO_194 (O_194,N_14457,N_14057);
and UO_195 (O_195,N_13737,N_14990);
nand UO_196 (O_196,N_13609,N_14481);
nand UO_197 (O_197,N_14027,N_13816);
nand UO_198 (O_198,N_13846,N_14073);
nor UO_199 (O_199,N_14613,N_13794);
and UO_200 (O_200,N_14545,N_13933);
or UO_201 (O_201,N_13896,N_13735);
and UO_202 (O_202,N_14883,N_13889);
and UO_203 (O_203,N_13644,N_14742);
or UO_204 (O_204,N_13894,N_13968);
and UO_205 (O_205,N_13654,N_14077);
and UO_206 (O_206,N_13928,N_14454);
nand UO_207 (O_207,N_14065,N_14346);
or UO_208 (O_208,N_14655,N_14340);
nor UO_209 (O_209,N_13995,N_13621);
and UO_210 (O_210,N_14164,N_14136);
and UO_211 (O_211,N_14031,N_13883);
or UO_212 (O_212,N_13558,N_14178);
and UO_213 (O_213,N_14423,N_14976);
nor UO_214 (O_214,N_14739,N_14147);
nand UO_215 (O_215,N_13902,N_14251);
nor UO_216 (O_216,N_14111,N_14288);
nor UO_217 (O_217,N_13655,N_14783);
nand UO_218 (O_218,N_14256,N_13718);
nor UO_219 (O_219,N_13611,N_14377);
or UO_220 (O_220,N_14236,N_14212);
and UO_221 (O_221,N_14188,N_14711);
nor UO_222 (O_222,N_13632,N_13704);
and UO_223 (O_223,N_13694,N_14078);
nand UO_224 (O_224,N_14268,N_14422);
and UO_225 (O_225,N_14590,N_14356);
and UO_226 (O_226,N_14763,N_14300);
and UO_227 (O_227,N_14401,N_14892);
nand UO_228 (O_228,N_14344,N_14544);
or UO_229 (O_229,N_14549,N_14371);
or UO_230 (O_230,N_13783,N_13836);
and UO_231 (O_231,N_14072,N_14986);
nor UO_232 (O_232,N_14333,N_14315);
nand UO_233 (O_233,N_14611,N_14100);
and UO_234 (O_234,N_14918,N_13899);
nand UO_235 (O_235,N_13696,N_14080);
or UO_236 (O_236,N_13638,N_13635);
or UO_237 (O_237,N_13731,N_14766);
and UO_238 (O_238,N_14518,N_14412);
and UO_239 (O_239,N_14964,N_13957);
nor UO_240 (O_240,N_14465,N_14802);
nor UO_241 (O_241,N_14390,N_14569);
or UO_242 (O_242,N_14748,N_14233);
and UO_243 (O_243,N_13573,N_14703);
or UO_244 (O_244,N_14270,N_14324);
nor UO_245 (O_245,N_14524,N_14705);
and UO_246 (O_246,N_14639,N_14293);
nor UO_247 (O_247,N_14685,N_14675);
nand UO_248 (O_248,N_14087,N_13699);
nor UO_249 (O_249,N_14635,N_14547);
nand UO_250 (O_250,N_13740,N_14915);
nand UO_251 (O_251,N_14102,N_13774);
or UO_252 (O_252,N_14483,N_14596);
nand UO_253 (O_253,N_13730,N_13796);
xnor UO_254 (O_254,N_14760,N_14254);
or UO_255 (O_255,N_14674,N_14956);
and UO_256 (O_256,N_13965,N_14692);
or UO_257 (O_257,N_14283,N_14160);
nand UO_258 (O_258,N_14473,N_14051);
or UO_259 (O_259,N_14768,N_14824);
nand UO_260 (O_260,N_14950,N_14939);
and UO_261 (O_261,N_13710,N_14186);
and UO_262 (O_262,N_14999,N_14682);
nand UO_263 (O_263,N_14466,N_14382);
and UO_264 (O_264,N_14131,N_14656);
or UO_265 (O_265,N_14792,N_14904);
or UO_266 (O_266,N_14005,N_14252);
and UO_267 (O_267,N_14517,N_13994);
and UO_268 (O_268,N_14680,N_14600);
or UO_269 (O_269,N_14992,N_14280);
nand UO_270 (O_270,N_13940,N_14932);
nor UO_271 (O_271,N_14819,N_14109);
xnor UO_272 (O_272,N_14851,N_14013);
xor UO_273 (O_273,N_14757,N_13661);
nand UO_274 (O_274,N_14874,N_14847);
nor UO_275 (O_275,N_14495,N_14347);
nand UO_276 (O_276,N_14447,N_14663);
nor UO_277 (O_277,N_14642,N_13706);
and UO_278 (O_278,N_14729,N_14378);
or UO_279 (O_279,N_14098,N_13629);
and UO_280 (O_280,N_13917,N_13535);
or UO_281 (O_281,N_14296,N_14654);
nor UO_282 (O_282,N_14210,N_14876);
nand UO_283 (O_283,N_14435,N_14970);
and UO_284 (O_284,N_14740,N_14603);
nor UO_285 (O_285,N_14648,N_14452);
or UO_286 (O_286,N_14399,N_13958);
nor UO_287 (O_287,N_14779,N_14506);
nor UO_288 (O_288,N_14249,N_14529);
or UO_289 (O_289,N_14235,N_14935);
nand UO_290 (O_290,N_14957,N_13977);
or UO_291 (O_291,N_14546,N_13990);
or UO_292 (O_292,N_14258,N_14420);
nand UO_293 (O_293,N_14563,N_13819);
and UO_294 (O_294,N_14905,N_14852);
nand UO_295 (O_295,N_13607,N_14631);
nand UO_296 (O_296,N_14501,N_14076);
or UO_297 (O_297,N_14383,N_13687);
nor UO_298 (O_298,N_14303,N_13714);
nor UO_299 (O_299,N_13682,N_13569);
nor UO_300 (O_300,N_14433,N_14341);
or UO_301 (O_301,N_14232,N_14239);
nand UO_302 (O_302,N_14983,N_14250);
and UO_303 (O_303,N_13516,N_14974);
nor UO_304 (O_304,N_14010,N_14138);
nor UO_305 (O_305,N_14927,N_14354);
and UO_306 (O_306,N_14834,N_14410);
xor UO_307 (O_307,N_13963,N_13686);
and UO_308 (O_308,N_13798,N_14942);
nand UO_309 (O_309,N_14949,N_13564);
nand UO_310 (O_310,N_14185,N_14702);
nand UO_311 (O_311,N_14272,N_14829);
nand UO_312 (O_312,N_14429,N_14710);
and UO_313 (O_313,N_13785,N_14963);
and UO_314 (O_314,N_13512,N_14593);
nand UO_315 (O_315,N_14756,N_14636);
nor UO_316 (O_316,N_13826,N_14908);
nor UO_317 (O_317,N_13723,N_14125);
or UO_318 (O_318,N_13856,N_14175);
nand UO_319 (O_319,N_14319,N_14869);
nor UO_320 (O_320,N_13628,N_14464);
nor UO_321 (O_321,N_14577,N_14245);
nor UO_322 (O_322,N_14261,N_13559);
or UO_323 (O_323,N_14132,N_13734);
nand UO_324 (O_324,N_14129,N_14000);
or UO_325 (O_325,N_14571,N_14020);
nor UO_326 (O_326,N_13993,N_14327);
and UO_327 (O_327,N_14734,N_14749);
and UO_328 (O_328,N_13757,N_14153);
nand UO_329 (O_329,N_13799,N_14022);
or UO_330 (O_330,N_13526,N_14989);
nor UO_331 (O_331,N_14722,N_13524);
and UO_332 (O_332,N_13538,N_14012);
or UO_333 (O_333,N_14265,N_14610);
nor UO_334 (O_334,N_13845,N_14723);
or UO_335 (O_335,N_13736,N_14696);
and UO_336 (O_336,N_14708,N_14946);
nand UO_337 (O_337,N_13966,N_14002);
nand UO_338 (O_338,N_14453,N_13608);
and UO_339 (O_339,N_14650,N_14514);
nand UO_340 (O_340,N_14681,N_14197);
nor UO_341 (O_341,N_14903,N_14947);
and UO_342 (O_342,N_13684,N_14598);
and UO_343 (O_343,N_14623,N_14854);
nor UO_344 (O_344,N_14940,N_14902);
and UO_345 (O_345,N_14162,N_14182);
or UO_346 (O_346,N_14052,N_13708);
nand UO_347 (O_347,N_14368,N_14516);
and UO_348 (O_348,N_14099,N_14234);
or UO_349 (O_349,N_14202,N_13981);
nand UO_350 (O_350,N_13947,N_14595);
nand UO_351 (O_351,N_14649,N_14643);
nand UO_352 (O_352,N_13585,N_13658);
nor UO_353 (O_353,N_14263,N_14796);
nand UO_354 (O_354,N_14825,N_14531);
nor UO_355 (O_355,N_14058,N_13534);
or UO_356 (O_356,N_14001,N_14769);
nor UO_357 (O_357,N_14380,N_13666);
nand UO_358 (O_358,N_13729,N_13892);
xor UO_359 (O_359,N_14041,N_14227);
nor UO_360 (O_360,N_13510,N_13909);
and UO_361 (O_361,N_14284,N_14009);
nand UO_362 (O_362,N_13886,N_14666);
nand UO_363 (O_363,N_14532,N_14025);
nand UO_364 (O_364,N_14553,N_14490);
nand UO_365 (O_365,N_13532,N_14764);
and UO_366 (O_366,N_14165,N_14978);
nand UO_367 (O_367,N_14875,N_14237);
or UO_368 (O_368,N_13668,N_14788);
or UO_369 (O_369,N_14067,N_14173);
and UO_370 (O_370,N_14615,N_14054);
or UO_371 (O_371,N_13832,N_14510);
and UO_372 (O_372,N_13903,N_14309);
nand UO_373 (O_373,N_14379,N_13700);
nor UO_374 (O_374,N_14392,N_14690);
nand UO_375 (O_375,N_14156,N_14204);
nand UO_376 (O_376,N_14211,N_13552);
or UO_377 (O_377,N_13866,N_13916);
and UO_378 (O_378,N_13582,N_13820);
and UO_379 (O_379,N_14625,N_14633);
nand UO_380 (O_380,N_13867,N_14848);
or UO_381 (O_381,N_14176,N_13508);
and UO_382 (O_382,N_14343,N_13606);
nor UO_383 (O_383,N_13576,N_14797);
or UO_384 (O_384,N_14480,N_13578);
nand UO_385 (O_385,N_14712,N_14088);
and UO_386 (O_386,N_13844,N_14115);
or UO_387 (O_387,N_14439,N_14438);
nor UO_388 (O_388,N_13574,N_13631);
or UO_389 (O_389,N_14450,N_14638);
nand UO_390 (O_390,N_14814,N_14014);
nand UO_391 (O_391,N_13614,N_14291);
or UO_392 (O_392,N_14269,N_14350);
nor UO_393 (O_393,N_14314,N_14170);
nand UO_394 (O_394,N_14436,N_13691);
or UO_395 (O_395,N_14984,N_13777);
nor UO_396 (O_396,N_13906,N_14372);
nand UO_397 (O_397,N_14475,N_14944);
and UO_398 (O_398,N_14169,N_14820);
nand UO_399 (O_399,N_13652,N_14896);
nor UO_400 (O_400,N_14091,N_14168);
or UO_401 (O_401,N_14406,N_14500);
or UO_402 (O_402,N_14934,N_14231);
nand UO_403 (O_403,N_14384,N_13667);
nand UO_404 (O_404,N_14142,N_14789);
xor UO_405 (O_405,N_13898,N_14555);
nor UO_406 (O_406,N_14807,N_14130);
nand UO_407 (O_407,N_13577,N_13619);
and UO_408 (O_408,N_13813,N_14428);
nand UO_409 (O_409,N_14732,N_13925);
nand UO_410 (O_410,N_14053,N_13676);
and UO_411 (O_411,N_14230,N_13812);
and UO_412 (O_412,N_13954,N_13643);
and UO_413 (O_413,N_14474,N_13584);
nor UO_414 (O_414,N_14542,N_14637);
nor UO_415 (O_415,N_14355,N_14721);
nand UO_416 (O_416,N_13772,N_13872);
and UO_417 (O_417,N_14297,N_13592);
and UO_418 (O_418,N_14278,N_14321);
nor UO_419 (O_419,N_14069,N_13952);
and UO_420 (O_420,N_13840,N_14404);
or UO_421 (O_421,N_13895,N_14396);
and UO_422 (O_422,N_14482,N_13597);
nor UO_423 (O_423,N_14411,N_13727);
and UO_424 (O_424,N_13912,N_14426);
nand UO_425 (O_425,N_14322,N_13835);
nor UO_426 (O_426,N_13509,N_13874);
or UO_427 (O_427,N_13612,N_14302);
nor UO_428 (O_428,N_14407,N_14916);
nor UO_429 (O_429,N_14266,N_14264);
nand UO_430 (O_430,N_13656,N_13674);
and UO_431 (O_431,N_13946,N_14840);
nor UO_432 (O_432,N_14697,N_14505);
or UO_433 (O_433,N_14857,N_14827);
nor UO_434 (O_434,N_14923,N_14677);
and UO_435 (O_435,N_13663,N_14352);
nand UO_436 (O_436,N_13529,N_14448);
or UO_437 (O_437,N_14290,N_13761);
nand UO_438 (O_438,N_14121,N_13501);
nand UO_439 (O_439,N_13789,N_14971);
and UO_440 (O_440,N_13897,N_14092);
nor UO_441 (O_441,N_14084,N_14771);
nor UO_442 (O_442,N_14445,N_13863);
nor UO_443 (O_443,N_13672,N_13839);
nand UO_444 (O_444,N_14714,N_14329);
and UO_445 (O_445,N_13759,N_14442);
or UO_446 (O_446,N_13797,N_14082);
nor UO_447 (O_447,N_13795,N_14241);
or UO_448 (O_448,N_14400,N_14737);
or UO_449 (O_449,N_14704,N_14301);
nand UO_450 (O_450,N_14730,N_14761);
nor UO_451 (O_451,N_14661,N_14207);
nand UO_452 (O_452,N_13693,N_13973);
nand UO_453 (O_453,N_14509,N_14842);
nor UO_454 (O_454,N_14931,N_14325);
nand UO_455 (O_455,N_14888,N_13943);
nand UO_456 (O_456,N_13885,N_13683);
nor UO_457 (O_457,N_14122,N_13972);
nand UO_458 (O_458,N_14866,N_13617);
nor UO_459 (O_459,N_14566,N_13587);
and UO_460 (O_460,N_13533,N_13637);
nor UO_461 (O_461,N_14906,N_14558);
or UO_462 (O_462,N_14573,N_14758);
nand UO_463 (O_463,N_14094,N_13918);
xnor UO_464 (O_464,N_14961,N_13712);
and UO_465 (O_465,N_13633,N_14951);
nand UO_466 (O_466,N_13689,N_13720);
nand UO_467 (O_467,N_13673,N_13950);
nand UO_468 (O_468,N_14519,N_14780);
nor UO_469 (O_469,N_14179,N_14962);
nor UO_470 (O_470,N_14221,N_14484);
nand UO_471 (O_471,N_14886,N_14914);
nand UO_472 (O_472,N_14930,N_14308);
nand UO_473 (O_473,N_14348,N_14180);
nor UO_474 (O_474,N_13861,N_13784);
and UO_475 (O_475,N_14794,N_14817);
nor UO_476 (O_476,N_13627,N_14751);
nand UO_477 (O_477,N_14365,N_13938);
and UO_478 (O_478,N_14006,N_14331);
xor UO_479 (O_479,N_14870,N_14520);
nand UO_480 (O_480,N_14096,N_14752);
and UO_481 (O_481,N_13769,N_14208);
and UO_482 (O_482,N_13803,N_14804);
nand UO_483 (O_483,N_14762,N_14455);
or UO_484 (O_484,N_14085,N_14800);
nor UO_485 (O_485,N_14535,N_14575);
nand UO_486 (O_486,N_14622,N_13805);
and UO_487 (O_487,N_14313,N_13583);
or UO_488 (O_488,N_14043,N_14167);
and UO_489 (O_489,N_14922,N_13528);
nand UO_490 (O_490,N_14733,N_14910);
and UO_491 (O_491,N_13951,N_13893);
nor UO_492 (O_492,N_14882,N_14223);
nor UO_493 (O_493,N_14086,N_14801);
nand UO_494 (O_494,N_14604,N_14491);
nand UO_495 (O_495,N_13561,N_14816);
or UO_496 (O_496,N_13598,N_14659);
and UO_497 (O_497,N_14864,N_14921);
and UO_498 (O_498,N_14653,N_13767);
nor UO_499 (O_499,N_14754,N_13882);
nor UO_500 (O_500,N_13590,N_13610);
or UO_501 (O_501,N_14991,N_14071);
nand UO_502 (O_502,N_13807,N_13842);
nor UO_503 (O_503,N_14209,N_14358);
nor UO_504 (O_504,N_13959,N_14127);
nand UO_505 (O_505,N_13679,N_14586);
nor UO_506 (O_506,N_14833,N_14775);
nor UO_507 (O_507,N_13986,N_13540);
or UO_508 (O_508,N_13725,N_14815);
nand UO_509 (O_509,N_14224,N_14134);
and UO_510 (O_510,N_14630,N_14591);
nand UO_511 (O_511,N_14548,N_14370);
nor UO_512 (O_512,N_14166,N_14929);
or UO_513 (O_513,N_14376,N_14727);
and UO_514 (O_514,N_13793,N_14981);
nor UO_515 (O_515,N_13600,N_14738);
nand UO_516 (O_516,N_13594,N_14229);
and UO_517 (O_517,N_14028,N_14691);
or UO_518 (O_518,N_13703,N_13778);
nand UO_519 (O_519,N_13743,N_13905);
and UO_520 (O_520,N_13764,N_13536);
nand UO_521 (O_521,N_13520,N_13875);
or UO_522 (O_522,N_14785,N_14200);
and UO_523 (O_523,N_14911,N_14725);
nand UO_524 (O_524,N_14045,N_13924);
and UO_525 (O_525,N_14812,N_14402);
or UO_526 (O_526,N_13560,N_13741);
or UO_527 (O_527,N_14110,N_14419);
or UO_528 (O_528,N_14538,N_13680);
nand UO_529 (O_529,N_14089,N_14953);
or UO_530 (O_530,N_14831,N_13876);
or UO_531 (O_531,N_14152,N_13549);
nand UO_532 (O_532,N_13755,N_13815);
or UO_533 (O_533,N_13507,N_14616);
nand UO_534 (O_534,N_14718,N_14822);
nand UO_535 (O_535,N_13879,N_14856);
and UO_536 (O_536,N_14446,N_14787);
or UO_537 (O_537,N_13604,N_14693);
and UO_538 (O_538,N_13929,N_14444);
or UO_539 (O_539,N_13669,N_14996);
nand UO_540 (O_540,N_14676,N_14295);
nand UO_541 (O_541,N_14437,N_14652);
nor UO_542 (O_542,N_14108,N_14507);
nand UO_543 (O_543,N_14046,N_13942);
and UO_544 (O_544,N_13675,N_14588);
nor UO_545 (O_545,N_14488,N_14567);
and UO_546 (O_546,N_13603,N_14627);
or UO_547 (O_547,N_14913,N_13978);
nor UO_548 (O_548,N_14534,N_14417);
or UO_549 (O_549,N_14667,N_13752);
or UO_550 (O_550,N_14713,N_14724);
nor UO_551 (O_551,N_14271,N_14260);
nand UO_552 (O_552,N_14151,N_14837);
or UO_553 (O_553,N_14339,N_14618);
nor UO_554 (O_554,N_13831,N_13849);
nand UO_555 (O_555,N_13841,N_13792);
and UO_556 (O_556,N_14050,N_14021);
and UO_557 (O_557,N_13521,N_14707);
nand UO_558 (O_558,N_14199,N_13988);
nor UO_559 (O_559,N_13754,N_13878);
xnor UO_560 (O_560,N_13571,N_14040);
or UO_561 (O_561,N_14557,N_14154);
or UO_562 (O_562,N_14144,N_14351);
or UO_563 (O_563,N_13890,N_14369);
nor UO_564 (O_564,N_14900,N_13505);
nand UO_565 (O_565,N_13599,N_14607);
nand UO_566 (O_566,N_13911,N_14502);
and UO_567 (O_567,N_14119,N_14478);
nor UO_568 (O_568,N_14240,N_14669);
and UO_569 (O_569,N_14767,N_14312);
and UO_570 (O_570,N_14409,N_14608);
nand UO_571 (O_571,N_13515,N_14081);
nor UO_572 (O_572,N_14735,N_14626);
nand UO_573 (O_573,N_13932,N_14338);
nor UO_574 (O_574,N_13565,N_13979);
or UO_575 (O_575,N_14863,N_14431);
or UO_576 (O_576,N_14471,N_14846);
and UO_577 (O_577,N_13997,N_14055);
and UO_578 (O_578,N_13745,N_13616);
or UO_579 (O_579,N_13920,N_14948);
nor UO_580 (O_580,N_14695,N_14632);
nor UO_581 (O_581,N_14781,N_13746);
and UO_582 (O_582,N_13987,N_14890);
xnor UO_583 (O_583,N_14213,N_14195);
and UO_584 (O_584,N_13984,N_14042);
and UO_585 (O_585,N_14218,N_14460);
and UO_586 (O_586,N_14821,N_14884);
nor UO_587 (O_587,N_13732,N_14449);
nor UO_588 (O_588,N_14839,N_13982);
nor UO_589 (O_589,N_13808,N_14899);
and UO_590 (O_590,N_13692,N_14244);
and UO_591 (O_591,N_14941,N_13775);
and UO_592 (O_592,N_14364,N_14793);
xnor UO_593 (O_593,N_14079,N_14373);
xnor UO_594 (O_594,N_13756,N_13542);
nand UO_595 (O_595,N_14499,N_14363);
nor UO_596 (O_596,N_13613,N_14609);
and UO_597 (O_597,N_14294,N_13698);
nand UO_598 (O_598,N_14592,N_14539);
and UO_599 (O_599,N_14361,N_14388);
nand UO_600 (O_600,N_14644,N_13719);
and UO_601 (O_601,N_13921,N_13562);
and UO_602 (O_602,N_14574,N_14059);
nand UO_603 (O_603,N_14980,N_13837);
or UO_604 (O_604,N_13758,N_13724);
nor UO_605 (O_605,N_14560,N_14097);
nor UO_606 (O_606,N_14128,N_14328);
or UO_607 (O_607,N_14451,N_14311);
nor UO_608 (O_608,N_14405,N_14060);
and UO_609 (O_609,N_14316,N_14282);
nor UO_610 (O_610,N_13926,N_14345);
and UO_611 (O_611,N_14019,N_14443);
nand UO_612 (O_612,N_14894,N_13843);
or UO_613 (O_613,N_13985,N_14878);
nand UO_614 (O_614,N_14879,N_14039);
and UO_615 (O_615,N_14120,N_14320);
nand UO_616 (O_616,N_14602,N_13922);
nand UO_617 (O_617,N_14522,N_13641);
nand UO_618 (O_618,N_13665,N_14056);
nor UO_619 (O_619,N_14061,N_13804);
or UO_620 (O_620,N_13937,N_13817);
and UO_621 (O_621,N_14494,N_14664);
and UO_622 (O_622,N_14565,N_13751);
nand UO_623 (O_623,N_14809,N_13513);
and UO_624 (O_624,N_14194,N_13527);
and UO_625 (O_625,N_14778,N_14965);
nand UO_626 (O_626,N_14530,N_14497);
nand UO_627 (O_627,N_14872,N_14107);
or UO_628 (O_628,N_14287,N_14599);
and UO_629 (O_629,N_14467,N_13568);
nor UO_630 (O_630,N_14580,N_13546);
nand UO_631 (O_631,N_13553,N_13622);
or UO_632 (O_632,N_14317,N_14281);
and UO_633 (O_633,N_14323,N_14198);
nor UO_634 (O_634,N_14425,N_14477);
and UO_635 (O_635,N_14689,N_14594);
or UO_636 (O_636,N_14541,N_14871);
and UO_637 (O_637,N_14349,N_14818);
nor UO_638 (O_638,N_14770,N_14408);
nor UO_639 (O_639,N_14678,N_14187);
nor UO_640 (O_640,N_13860,N_14394);
nor UO_641 (O_641,N_14850,N_14150);
or UO_642 (O_642,N_13588,N_13948);
and UO_643 (O_643,N_13790,N_14332);
and UO_644 (O_644,N_14937,N_13931);
and UO_645 (O_645,N_13847,N_14219);
nor UO_646 (O_646,N_14898,N_14972);
and UO_647 (O_647,N_14222,N_14959);
and UO_648 (O_648,N_14683,N_13554);
nor UO_649 (O_649,N_14985,N_14773);
and UO_650 (O_650,N_14701,N_14360);
or UO_651 (O_651,N_14273,N_14090);
nor UO_652 (O_652,N_13989,N_14584);
nand UO_653 (O_653,N_14220,N_14568);
nand UO_654 (O_654,N_13853,N_13935);
or UO_655 (O_655,N_14243,N_13548);
nor UO_656 (O_656,N_14135,N_14123);
or UO_657 (O_657,N_13930,N_14462);
or UO_658 (O_658,N_14512,N_14008);
and UO_659 (O_659,N_13828,N_14841);
or UO_660 (O_660,N_14508,N_14997);
nand UO_661 (O_661,N_14938,N_14397);
or UO_662 (O_662,N_14673,N_13781);
or UO_663 (O_663,N_14606,N_14362);
and UO_664 (O_664,N_14262,N_14418);
nand UO_665 (O_665,N_13887,N_14424);
and UO_666 (O_666,N_14858,N_14177);
and UO_667 (O_667,N_14034,N_14306);
and UO_668 (O_668,N_14161,N_14672);
nor UO_669 (O_669,N_14966,N_14790);
nor UO_670 (O_670,N_14753,N_14427);
nor UO_671 (O_671,N_14414,N_13763);
and UO_672 (O_672,N_13713,N_14719);
nand UO_673 (O_673,N_13539,N_14933);
nor UO_674 (O_674,N_13623,N_14226);
or UO_675 (O_675,N_14777,N_14246);
nor UO_676 (O_676,N_14660,N_13788);
nor UO_677 (O_677,N_14562,N_14011);
nand UO_678 (O_678,N_14385,N_14104);
nor UO_679 (O_679,N_14605,N_14103);
nor UO_680 (O_680,N_14299,N_14726);
nor UO_681 (O_681,N_14070,N_14843);
nor UO_682 (O_682,N_13825,N_13996);
or UO_683 (O_683,N_13664,N_14895);
and UO_684 (O_684,N_14255,N_13586);
nand UO_685 (O_685,N_14342,N_13705);
nor UO_686 (O_686,N_13733,N_14585);
and UO_687 (O_687,N_14698,N_14646);
or UO_688 (O_688,N_14274,N_13871);
nand UO_689 (O_689,N_13888,N_14621);
nor UO_690 (O_690,N_14973,N_14191);
nand UO_691 (O_691,N_14746,N_13880);
nand UO_692 (O_692,N_14868,N_14337);
and UO_693 (O_693,N_13744,N_13647);
or UO_694 (O_694,N_13913,N_13974);
nand UO_695 (O_695,N_13877,N_14279);
and UO_696 (O_696,N_13678,N_14137);
nor UO_697 (O_697,N_14064,N_14967);
and UO_698 (O_698,N_14049,N_14891);
nand UO_699 (O_699,N_14979,N_14513);
nand UO_700 (O_700,N_13695,N_14620);
or UO_701 (O_701,N_14657,N_13660);
nand UO_702 (O_702,N_14140,N_14018);
nor UO_703 (O_703,N_14304,N_14216);
nor UO_704 (O_704,N_14880,N_14113);
nand UO_705 (O_705,N_13750,N_14887);
nand UO_706 (O_706,N_13634,N_14835);
nor UO_707 (O_707,N_14215,N_14799);
nand UO_708 (O_708,N_14106,N_13690);
or UO_709 (O_709,N_14504,N_14647);
and UO_710 (O_710,N_14415,N_14936);
or UO_711 (O_711,N_14357,N_14743);
and UO_712 (O_712,N_14024,N_14440);
nor UO_713 (O_713,N_14901,N_13855);
nor UO_714 (O_714,N_14318,N_14798);
xor UO_715 (O_715,N_13891,N_13504);
and UO_716 (O_716,N_14995,N_14330);
nand UO_717 (O_717,N_14277,N_13834);
nor UO_718 (O_718,N_13547,N_13645);
and UO_719 (O_719,N_14326,N_13868);
and UO_720 (O_720,N_13809,N_13915);
and UO_721 (O_721,N_13848,N_14855);
nor UO_722 (O_722,N_14003,N_14062);
and UO_723 (O_723,N_13681,N_13595);
nand UO_724 (O_724,N_14017,N_13934);
or UO_725 (O_725,N_14658,N_13962);
and UO_726 (O_726,N_13862,N_13620);
nor UO_727 (O_727,N_13907,N_13992);
nand UO_728 (O_728,N_14189,N_14193);
nand UO_729 (O_729,N_13998,N_13881);
nand UO_730 (O_730,N_14629,N_13811);
nand UO_731 (O_731,N_14543,N_14366);
and UO_732 (O_732,N_13579,N_13519);
or UO_733 (O_733,N_13581,N_14662);
nand UO_734 (O_734,N_13642,N_13854);
nand UO_735 (O_735,N_13570,N_14286);
and UO_736 (O_736,N_13551,N_14578);
nor UO_737 (O_737,N_14561,N_14803);
nand UO_738 (O_738,N_14430,N_14826);
and UO_739 (O_739,N_14381,N_13975);
or UO_740 (O_740,N_14267,N_13662);
and UO_741 (O_741,N_14861,N_13677);
xnor UO_742 (O_742,N_14118,N_14413);
nand UO_743 (O_743,N_13949,N_14684);
nor UO_744 (O_744,N_14116,N_14897);
or UO_745 (O_745,N_13726,N_13648);
nor UO_746 (O_746,N_14184,N_13722);
and UO_747 (O_747,N_14836,N_13864);
nor UO_748 (O_748,N_14808,N_14612);
nand UO_749 (O_749,N_14203,N_14926);
nor UO_750 (O_750,N_14720,N_14201);
or UO_751 (O_751,N_14014,N_14216);
xnor UO_752 (O_752,N_14557,N_14519);
or UO_753 (O_753,N_14039,N_14667);
and UO_754 (O_754,N_14118,N_14193);
or UO_755 (O_755,N_14847,N_14073);
nand UO_756 (O_756,N_13997,N_13939);
and UO_757 (O_757,N_14936,N_14174);
nand UO_758 (O_758,N_14929,N_14087);
nor UO_759 (O_759,N_14727,N_14884);
and UO_760 (O_760,N_14518,N_14237);
or UO_761 (O_761,N_14471,N_13692);
or UO_762 (O_762,N_14673,N_14575);
nor UO_763 (O_763,N_14718,N_14780);
nand UO_764 (O_764,N_14066,N_14911);
or UO_765 (O_765,N_13659,N_14794);
nor UO_766 (O_766,N_14536,N_13871);
nand UO_767 (O_767,N_14508,N_13624);
nor UO_768 (O_768,N_13637,N_14477);
or UO_769 (O_769,N_13706,N_14294);
and UO_770 (O_770,N_13826,N_14746);
or UO_771 (O_771,N_14709,N_14686);
or UO_772 (O_772,N_14398,N_13617);
nor UO_773 (O_773,N_14081,N_14976);
or UO_774 (O_774,N_14990,N_13561);
nor UO_775 (O_775,N_13930,N_13855);
or UO_776 (O_776,N_14333,N_13915);
and UO_777 (O_777,N_13724,N_14904);
or UO_778 (O_778,N_13932,N_14865);
or UO_779 (O_779,N_13838,N_13722);
nor UO_780 (O_780,N_14235,N_13780);
or UO_781 (O_781,N_13785,N_14103);
nor UO_782 (O_782,N_14360,N_14673);
and UO_783 (O_783,N_14493,N_14653);
or UO_784 (O_784,N_13762,N_14057);
or UO_785 (O_785,N_14230,N_13987);
nand UO_786 (O_786,N_13964,N_14904);
nor UO_787 (O_787,N_14279,N_14588);
nand UO_788 (O_788,N_14525,N_14446);
nand UO_789 (O_789,N_14493,N_14612);
or UO_790 (O_790,N_14009,N_14311);
or UO_791 (O_791,N_14600,N_14493);
nor UO_792 (O_792,N_14591,N_14730);
nor UO_793 (O_793,N_14383,N_13541);
nor UO_794 (O_794,N_14916,N_13845);
nand UO_795 (O_795,N_14934,N_14188);
nor UO_796 (O_796,N_14010,N_14898);
and UO_797 (O_797,N_14846,N_13825);
nand UO_798 (O_798,N_13786,N_13946);
or UO_799 (O_799,N_13558,N_14785);
nor UO_800 (O_800,N_13637,N_13666);
and UO_801 (O_801,N_14643,N_14320);
and UO_802 (O_802,N_14829,N_13829);
nor UO_803 (O_803,N_14109,N_14127);
nor UO_804 (O_804,N_13738,N_14513);
xor UO_805 (O_805,N_14513,N_14232);
and UO_806 (O_806,N_13718,N_14282);
nand UO_807 (O_807,N_14294,N_14295);
or UO_808 (O_808,N_14879,N_13708);
nor UO_809 (O_809,N_13536,N_14952);
or UO_810 (O_810,N_14810,N_14125);
nor UO_811 (O_811,N_14029,N_13807);
and UO_812 (O_812,N_14769,N_14544);
or UO_813 (O_813,N_13556,N_14002);
or UO_814 (O_814,N_13736,N_13660);
and UO_815 (O_815,N_14695,N_13883);
and UO_816 (O_816,N_13550,N_14992);
or UO_817 (O_817,N_14578,N_13530);
nor UO_818 (O_818,N_14296,N_13845);
or UO_819 (O_819,N_14144,N_13986);
or UO_820 (O_820,N_13834,N_14402);
nand UO_821 (O_821,N_13617,N_13747);
or UO_822 (O_822,N_14583,N_14783);
or UO_823 (O_823,N_14616,N_14302);
and UO_824 (O_824,N_14498,N_13719);
nor UO_825 (O_825,N_14446,N_14688);
and UO_826 (O_826,N_13545,N_14463);
and UO_827 (O_827,N_14006,N_14466);
nor UO_828 (O_828,N_14170,N_13569);
and UO_829 (O_829,N_14815,N_13961);
and UO_830 (O_830,N_14152,N_14149);
or UO_831 (O_831,N_13949,N_13654);
nor UO_832 (O_832,N_14780,N_13812);
nor UO_833 (O_833,N_14212,N_14191);
xnor UO_834 (O_834,N_14459,N_13994);
nand UO_835 (O_835,N_14652,N_14176);
nand UO_836 (O_836,N_14717,N_13515);
and UO_837 (O_837,N_14388,N_13616);
and UO_838 (O_838,N_14811,N_13992);
and UO_839 (O_839,N_13765,N_14814);
or UO_840 (O_840,N_14398,N_14882);
or UO_841 (O_841,N_13699,N_14422);
or UO_842 (O_842,N_14114,N_13904);
and UO_843 (O_843,N_14722,N_14328);
or UO_844 (O_844,N_14876,N_13991);
nand UO_845 (O_845,N_13830,N_14598);
nor UO_846 (O_846,N_14223,N_14840);
nor UO_847 (O_847,N_14261,N_14291);
nor UO_848 (O_848,N_14528,N_13960);
and UO_849 (O_849,N_14911,N_14095);
or UO_850 (O_850,N_13550,N_13693);
and UO_851 (O_851,N_13693,N_14766);
nor UO_852 (O_852,N_14397,N_14463);
or UO_853 (O_853,N_14970,N_14105);
or UO_854 (O_854,N_14817,N_13524);
nor UO_855 (O_855,N_14311,N_13764);
and UO_856 (O_856,N_14605,N_13963);
and UO_857 (O_857,N_13581,N_14887);
and UO_858 (O_858,N_14993,N_14872);
nor UO_859 (O_859,N_14778,N_13666);
or UO_860 (O_860,N_13691,N_14253);
or UO_861 (O_861,N_14675,N_14385);
nand UO_862 (O_862,N_14418,N_13984);
nand UO_863 (O_863,N_14067,N_13915);
or UO_864 (O_864,N_14980,N_14835);
and UO_865 (O_865,N_14314,N_13759);
nor UO_866 (O_866,N_14658,N_13701);
nand UO_867 (O_867,N_14694,N_13620);
nor UO_868 (O_868,N_14301,N_14792);
nand UO_869 (O_869,N_14462,N_14658);
nand UO_870 (O_870,N_14064,N_13707);
nand UO_871 (O_871,N_14076,N_14202);
and UO_872 (O_872,N_14215,N_14622);
nor UO_873 (O_873,N_14125,N_14548);
and UO_874 (O_874,N_14660,N_14022);
and UO_875 (O_875,N_14300,N_13768);
and UO_876 (O_876,N_14496,N_14374);
nand UO_877 (O_877,N_14717,N_14511);
nand UO_878 (O_878,N_14052,N_14809);
nand UO_879 (O_879,N_14061,N_14774);
and UO_880 (O_880,N_13788,N_13718);
nand UO_881 (O_881,N_14726,N_14461);
and UO_882 (O_882,N_13820,N_14310);
and UO_883 (O_883,N_14966,N_13947);
nand UO_884 (O_884,N_14049,N_13837);
nand UO_885 (O_885,N_14371,N_14200);
nor UO_886 (O_886,N_14594,N_14158);
nor UO_887 (O_887,N_14897,N_13752);
nand UO_888 (O_888,N_14962,N_13958);
nor UO_889 (O_889,N_14972,N_14046);
nand UO_890 (O_890,N_14492,N_14258);
and UO_891 (O_891,N_13671,N_14839);
nand UO_892 (O_892,N_13840,N_13505);
and UO_893 (O_893,N_14838,N_14069);
and UO_894 (O_894,N_14989,N_13754);
nor UO_895 (O_895,N_14399,N_14876);
nor UO_896 (O_896,N_14568,N_14330);
or UO_897 (O_897,N_14040,N_14520);
nor UO_898 (O_898,N_14264,N_13518);
and UO_899 (O_899,N_14919,N_14611);
nor UO_900 (O_900,N_13580,N_14337);
nor UO_901 (O_901,N_14373,N_13657);
nor UO_902 (O_902,N_14455,N_13943);
nand UO_903 (O_903,N_14047,N_14467);
or UO_904 (O_904,N_14174,N_14494);
nor UO_905 (O_905,N_14408,N_14821);
or UO_906 (O_906,N_13701,N_14204);
nor UO_907 (O_907,N_14145,N_14631);
nand UO_908 (O_908,N_14884,N_13728);
nor UO_909 (O_909,N_14127,N_14126);
and UO_910 (O_910,N_14715,N_14760);
xnor UO_911 (O_911,N_14292,N_13528);
nand UO_912 (O_912,N_14645,N_14454);
or UO_913 (O_913,N_14098,N_14663);
or UO_914 (O_914,N_14230,N_14250);
and UO_915 (O_915,N_14484,N_13578);
or UO_916 (O_916,N_13950,N_13532);
or UO_917 (O_917,N_14062,N_14960);
or UO_918 (O_918,N_14680,N_13993);
nor UO_919 (O_919,N_14340,N_13719);
nand UO_920 (O_920,N_14132,N_14593);
or UO_921 (O_921,N_14470,N_14595);
or UO_922 (O_922,N_14379,N_14831);
xnor UO_923 (O_923,N_14340,N_14973);
and UO_924 (O_924,N_13748,N_14342);
nor UO_925 (O_925,N_13743,N_14179);
xor UO_926 (O_926,N_14087,N_14524);
nor UO_927 (O_927,N_14901,N_13527);
and UO_928 (O_928,N_14793,N_13816);
and UO_929 (O_929,N_14278,N_13923);
and UO_930 (O_930,N_14130,N_14760);
nand UO_931 (O_931,N_14873,N_14066);
and UO_932 (O_932,N_14111,N_14860);
or UO_933 (O_933,N_14933,N_14459);
nor UO_934 (O_934,N_14502,N_13732);
nor UO_935 (O_935,N_14082,N_13995);
nand UO_936 (O_936,N_13680,N_14196);
and UO_937 (O_937,N_14607,N_14590);
or UO_938 (O_938,N_14879,N_14145);
and UO_939 (O_939,N_13555,N_14106);
nand UO_940 (O_940,N_14284,N_13649);
nand UO_941 (O_941,N_14956,N_14513);
nand UO_942 (O_942,N_13687,N_14169);
or UO_943 (O_943,N_13654,N_14648);
or UO_944 (O_944,N_14613,N_13691);
or UO_945 (O_945,N_13636,N_14010);
and UO_946 (O_946,N_14348,N_14092);
nor UO_947 (O_947,N_13883,N_14246);
nor UO_948 (O_948,N_14342,N_13812);
and UO_949 (O_949,N_14529,N_14764);
nand UO_950 (O_950,N_13975,N_13842);
nand UO_951 (O_951,N_14357,N_14966);
or UO_952 (O_952,N_14678,N_14499);
nor UO_953 (O_953,N_14256,N_13630);
nor UO_954 (O_954,N_14919,N_14020);
nor UO_955 (O_955,N_14902,N_14135);
and UO_956 (O_956,N_14930,N_14065);
nor UO_957 (O_957,N_14800,N_14951);
or UO_958 (O_958,N_14683,N_14758);
or UO_959 (O_959,N_13554,N_14037);
nor UO_960 (O_960,N_14690,N_14898);
and UO_961 (O_961,N_14742,N_14200);
nor UO_962 (O_962,N_14719,N_13882);
nand UO_963 (O_963,N_14124,N_13754);
nand UO_964 (O_964,N_13736,N_14922);
nand UO_965 (O_965,N_14843,N_13904);
nor UO_966 (O_966,N_13851,N_14921);
nand UO_967 (O_967,N_14697,N_14975);
xor UO_968 (O_968,N_14272,N_14387);
nand UO_969 (O_969,N_14917,N_14372);
and UO_970 (O_970,N_14299,N_13973);
nand UO_971 (O_971,N_14311,N_14584);
or UO_972 (O_972,N_14826,N_14006);
nor UO_973 (O_973,N_13612,N_14526);
and UO_974 (O_974,N_13902,N_13959);
nand UO_975 (O_975,N_14043,N_14047);
or UO_976 (O_976,N_14035,N_14449);
or UO_977 (O_977,N_14041,N_13934);
nor UO_978 (O_978,N_14533,N_13697);
nor UO_979 (O_979,N_13938,N_13654);
nand UO_980 (O_980,N_14773,N_14094);
or UO_981 (O_981,N_13967,N_14500);
nor UO_982 (O_982,N_14910,N_14708);
nor UO_983 (O_983,N_14086,N_14263);
and UO_984 (O_984,N_14606,N_14984);
nand UO_985 (O_985,N_14176,N_14051);
nor UO_986 (O_986,N_14511,N_13947);
nand UO_987 (O_987,N_14446,N_14325);
nand UO_988 (O_988,N_14391,N_13992);
and UO_989 (O_989,N_14966,N_13868);
and UO_990 (O_990,N_14777,N_13707);
or UO_991 (O_991,N_14997,N_14760);
nand UO_992 (O_992,N_14736,N_14980);
and UO_993 (O_993,N_13600,N_14108);
nor UO_994 (O_994,N_14987,N_13978);
and UO_995 (O_995,N_14561,N_14600);
and UO_996 (O_996,N_14597,N_14533);
or UO_997 (O_997,N_14837,N_13950);
nor UO_998 (O_998,N_13780,N_14327);
nand UO_999 (O_999,N_14781,N_14422);
and UO_1000 (O_1000,N_14879,N_14711);
and UO_1001 (O_1001,N_14629,N_14285);
or UO_1002 (O_1002,N_14788,N_14306);
or UO_1003 (O_1003,N_14092,N_13579);
nor UO_1004 (O_1004,N_14161,N_13564);
and UO_1005 (O_1005,N_13719,N_14515);
and UO_1006 (O_1006,N_14473,N_14137);
and UO_1007 (O_1007,N_13834,N_13634);
or UO_1008 (O_1008,N_14550,N_14467);
or UO_1009 (O_1009,N_13883,N_14128);
nand UO_1010 (O_1010,N_13689,N_13657);
nand UO_1011 (O_1011,N_14437,N_13840);
nand UO_1012 (O_1012,N_14443,N_14249);
and UO_1013 (O_1013,N_14271,N_14903);
nand UO_1014 (O_1014,N_14137,N_14130);
and UO_1015 (O_1015,N_13773,N_14210);
nor UO_1016 (O_1016,N_13796,N_14711);
or UO_1017 (O_1017,N_14238,N_14029);
nor UO_1018 (O_1018,N_14384,N_14850);
and UO_1019 (O_1019,N_14614,N_14037);
or UO_1020 (O_1020,N_13749,N_13865);
nor UO_1021 (O_1021,N_14260,N_14971);
nand UO_1022 (O_1022,N_13611,N_14004);
nor UO_1023 (O_1023,N_14930,N_13697);
nand UO_1024 (O_1024,N_14662,N_14569);
nor UO_1025 (O_1025,N_14166,N_14054);
or UO_1026 (O_1026,N_14720,N_13694);
and UO_1027 (O_1027,N_14273,N_14529);
nand UO_1028 (O_1028,N_13994,N_13738);
or UO_1029 (O_1029,N_14274,N_14245);
xnor UO_1030 (O_1030,N_14238,N_14502);
nor UO_1031 (O_1031,N_14764,N_14049);
and UO_1032 (O_1032,N_14361,N_13596);
or UO_1033 (O_1033,N_14478,N_13757);
nand UO_1034 (O_1034,N_14903,N_13547);
or UO_1035 (O_1035,N_14200,N_14122);
or UO_1036 (O_1036,N_14910,N_13906);
nand UO_1037 (O_1037,N_13798,N_13623);
and UO_1038 (O_1038,N_14815,N_14039);
or UO_1039 (O_1039,N_14165,N_14973);
or UO_1040 (O_1040,N_13757,N_14320);
and UO_1041 (O_1041,N_13974,N_13938);
nor UO_1042 (O_1042,N_13913,N_14018);
nor UO_1043 (O_1043,N_14540,N_14671);
or UO_1044 (O_1044,N_14409,N_13609);
nand UO_1045 (O_1045,N_13901,N_13668);
nor UO_1046 (O_1046,N_13897,N_14689);
nor UO_1047 (O_1047,N_13877,N_14391);
nor UO_1048 (O_1048,N_14948,N_13815);
nand UO_1049 (O_1049,N_14757,N_14332);
nor UO_1050 (O_1050,N_14327,N_13835);
nor UO_1051 (O_1051,N_14422,N_13804);
or UO_1052 (O_1052,N_14052,N_13809);
or UO_1053 (O_1053,N_14403,N_14138);
nand UO_1054 (O_1054,N_13573,N_13958);
nand UO_1055 (O_1055,N_14486,N_14878);
or UO_1056 (O_1056,N_14048,N_14684);
nand UO_1057 (O_1057,N_14311,N_14927);
nor UO_1058 (O_1058,N_14835,N_14460);
nand UO_1059 (O_1059,N_14433,N_14987);
nand UO_1060 (O_1060,N_14090,N_14026);
nor UO_1061 (O_1061,N_13941,N_14394);
nand UO_1062 (O_1062,N_14647,N_13714);
nor UO_1063 (O_1063,N_14914,N_14577);
nor UO_1064 (O_1064,N_14948,N_14265);
nor UO_1065 (O_1065,N_13759,N_14133);
nor UO_1066 (O_1066,N_14217,N_13638);
and UO_1067 (O_1067,N_14603,N_13927);
and UO_1068 (O_1068,N_13834,N_14701);
and UO_1069 (O_1069,N_14436,N_14285);
or UO_1070 (O_1070,N_14459,N_14466);
nand UO_1071 (O_1071,N_14409,N_14624);
nand UO_1072 (O_1072,N_14561,N_14595);
nor UO_1073 (O_1073,N_14592,N_14128);
nand UO_1074 (O_1074,N_14353,N_13879);
nand UO_1075 (O_1075,N_14082,N_13682);
and UO_1076 (O_1076,N_13967,N_13957);
or UO_1077 (O_1077,N_14063,N_14335);
xor UO_1078 (O_1078,N_14238,N_13735);
and UO_1079 (O_1079,N_14725,N_14826);
nor UO_1080 (O_1080,N_14561,N_14184);
or UO_1081 (O_1081,N_13633,N_14180);
nor UO_1082 (O_1082,N_13700,N_13848);
or UO_1083 (O_1083,N_14002,N_14433);
nand UO_1084 (O_1084,N_14024,N_14802);
or UO_1085 (O_1085,N_14113,N_13505);
nand UO_1086 (O_1086,N_13590,N_13718);
and UO_1087 (O_1087,N_14189,N_14949);
nor UO_1088 (O_1088,N_14959,N_14269);
nor UO_1089 (O_1089,N_14162,N_14097);
nor UO_1090 (O_1090,N_13697,N_14151);
nand UO_1091 (O_1091,N_14626,N_14605);
and UO_1092 (O_1092,N_14500,N_14308);
and UO_1093 (O_1093,N_14973,N_13886);
and UO_1094 (O_1094,N_14581,N_14058);
or UO_1095 (O_1095,N_14827,N_14896);
nand UO_1096 (O_1096,N_14398,N_13623);
or UO_1097 (O_1097,N_14143,N_14180);
and UO_1098 (O_1098,N_14180,N_14481);
nand UO_1099 (O_1099,N_13815,N_13745);
nand UO_1100 (O_1100,N_14041,N_13532);
and UO_1101 (O_1101,N_14545,N_14266);
or UO_1102 (O_1102,N_13823,N_14652);
nand UO_1103 (O_1103,N_14378,N_13966);
nand UO_1104 (O_1104,N_13636,N_14037);
and UO_1105 (O_1105,N_14665,N_13988);
and UO_1106 (O_1106,N_13849,N_14541);
nor UO_1107 (O_1107,N_14655,N_13619);
and UO_1108 (O_1108,N_14735,N_14452);
and UO_1109 (O_1109,N_14888,N_14378);
nand UO_1110 (O_1110,N_14808,N_13866);
nand UO_1111 (O_1111,N_14470,N_14363);
and UO_1112 (O_1112,N_14395,N_13633);
or UO_1113 (O_1113,N_14088,N_14741);
nand UO_1114 (O_1114,N_13630,N_13971);
and UO_1115 (O_1115,N_13536,N_13605);
nor UO_1116 (O_1116,N_14659,N_14509);
and UO_1117 (O_1117,N_14461,N_14312);
or UO_1118 (O_1118,N_14035,N_14460);
or UO_1119 (O_1119,N_13915,N_14851);
nor UO_1120 (O_1120,N_14398,N_14905);
nand UO_1121 (O_1121,N_14700,N_14211);
and UO_1122 (O_1122,N_14860,N_14490);
nand UO_1123 (O_1123,N_13569,N_13965);
nand UO_1124 (O_1124,N_14188,N_13535);
nand UO_1125 (O_1125,N_13730,N_13535);
nand UO_1126 (O_1126,N_13953,N_14028);
and UO_1127 (O_1127,N_14852,N_14048);
or UO_1128 (O_1128,N_13619,N_14168);
or UO_1129 (O_1129,N_14636,N_14410);
and UO_1130 (O_1130,N_13869,N_14582);
nand UO_1131 (O_1131,N_14745,N_13691);
and UO_1132 (O_1132,N_14668,N_14939);
nand UO_1133 (O_1133,N_14896,N_14557);
and UO_1134 (O_1134,N_13982,N_14747);
nand UO_1135 (O_1135,N_14992,N_14803);
nor UO_1136 (O_1136,N_13805,N_13961);
or UO_1137 (O_1137,N_14788,N_13922);
nor UO_1138 (O_1138,N_14034,N_13761);
nor UO_1139 (O_1139,N_14559,N_13995);
nand UO_1140 (O_1140,N_14981,N_13875);
nor UO_1141 (O_1141,N_13751,N_14648);
nor UO_1142 (O_1142,N_14813,N_14114);
or UO_1143 (O_1143,N_13676,N_13971);
nor UO_1144 (O_1144,N_14617,N_13643);
and UO_1145 (O_1145,N_14657,N_14558);
nand UO_1146 (O_1146,N_13822,N_14460);
nand UO_1147 (O_1147,N_14127,N_14411);
nand UO_1148 (O_1148,N_14482,N_14455);
nand UO_1149 (O_1149,N_13871,N_14902);
and UO_1150 (O_1150,N_13900,N_14013);
and UO_1151 (O_1151,N_14043,N_14236);
or UO_1152 (O_1152,N_13551,N_14296);
or UO_1153 (O_1153,N_14059,N_13927);
or UO_1154 (O_1154,N_13540,N_13583);
and UO_1155 (O_1155,N_13784,N_13748);
nor UO_1156 (O_1156,N_14507,N_13816);
and UO_1157 (O_1157,N_14541,N_14158);
and UO_1158 (O_1158,N_14740,N_14756);
or UO_1159 (O_1159,N_14924,N_14921);
nor UO_1160 (O_1160,N_14267,N_14432);
nor UO_1161 (O_1161,N_14025,N_14506);
nand UO_1162 (O_1162,N_14462,N_13801);
nor UO_1163 (O_1163,N_14778,N_14203);
nand UO_1164 (O_1164,N_14570,N_14393);
nand UO_1165 (O_1165,N_14448,N_14258);
or UO_1166 (O_1166,N_13590,N_14549);
or UO_1167 (O_1167,N_14575,N_13798);
and UO_1168 (O_1168,N_14723,N_13631);
or UO_1169 (O_1169,N_14940,N_14302);
nand UO_1170 (O_1170,N_14993,N_13520);
nor UO_1171 (O_1171,N_14908,N_14333);
or UO_1172 (O_1172,N_14057,N_13708);
nand UO_1173 (O_1173,N_14367,N_14075);
nor UO_1174 (O_1174,N_14151,N_13986);
nor UO_1175 (O_1175,N_14426,N_14578);
or UO_1176 (O_1176,N_14015,N_14115);
or UO_1177 (O_1177,N_14111,N_14657);
and UO_1178 (O_1178,N_13876,N_14935);
or UO_1179 (O_1179,N_13776,N_13823);
xor UO_1180 (O_1180,N_14960,N_14179);
nor UO_1181 (O_1181,N_13509,N_14545);
and UO_1182 (O_1182,N_13545,N_14714);
and UO_1183 (O_1183,N_13972,N_14888);
and UO_1184 (O_1184,N_14678,N_14672);
nor UO_1185 (O_1185,N_14884,N_14590);
nand UO_1186 (O_1186,N_14581,N_13667);
nand UO_1187 (O_1187,N_13802,N_13769);
and UO_1188 (O_1188,N_14473,N_14997);
and UO_1189 (O_1189,N_14757,N_13677);
and UO_1190 (O_1190,N_14977,N_14098);
and UO_1191 (O_1191,N_14635,N_13724);
nand UO_1192 (O_1192,N_14870,N_14848);
or UO_1193 (O_1193,N_14521,N_14799);
or UO_1194 (O_1194,N_13799,N_13660);
nand UO_1195 (O_1195,N_13943,N_13912);
nor UO_1196 (O_1196,N_13897,N_13945);
nand UO_1197 (O_1197,N_14804,N_14114);
or UO_1198 (O_1198,N_14351,N_14069);
nand UO_1199 (O_1199,N_14763,N_13670);
nor UO_1200 (O_1200,N_14643,N_13936);
or UO_1201 (O_1201,N_14135,N_14603);
nor UO_1202 (O_1202,N_13664,N_14116);
nor UO_1203 (O_1203,N_14604,N_14024);
nor UO_1204 (O_1204,N_14032,N_14535);
or UO_1205 (O_1205,N_13676,N_14278);
and UO_1206 (O_1206,N_14537,N_14096);
nor UO_1207 (O_1207,N_13992,N_14330);
xor UO_1208 (O_1208,N_13847,N_14536);
nor UO_1209 (O_1209,N_13537,N_14297);
nand UO_1210 (O_1210,N_13995,N_13588);
and UO_1211 (O_1211,N_13979,N_14162);
and UO_1212 (O_1212,N_14412,N_14616);
or UO_1213 (O_1213,N_14564,N_13941);
nor UO_1214 (O_1214,N_13711,N_14901);
nand UO_1215 (O_1215,N_13797,N_13659);
nand UO_1216 (O_1216,N_14828,N_13807);
nand UO_1217 (O_1217,N_14859,N_14643);
nand UO_1218 (O_1218,N_14822,N_14182);
nand UO_1219 (O_1219,N_14440,N_14386);
or UO_1220 (O_1220,N_14661,N_13563);
nand UO_1221 (O_1221,N_13715,N_14910);
xnor UO_1222 (O_1222,N_13922,N_13839);
nor UO_1223 (O_1223,N_13517,N_14203);
and UO_1224 (O_1224,N_14147,N_14275);
nand UO_1225 (O_1225,N_14538,N_14206);
and UO_1226 (O_1226,N_14279,N_14136);
and UO_1227 (O_1227,N_13686,N_14308);
and UO_1228 (O_1228,N_13814,N_13626);
or UO_1229 (O_1229,N_14579,N_13907);
nand UO_1230 (O_1230,N_14368,N_14674);
nor UO_1231 (O_1231,N_14540,N_14891);
or UO_1232 (O_1232,N_14216,N_14835);
or UO_1233 (O_1233,N_14995,N_14787);
nand UO_1234 (O_1234,N_14268,N_13685);
nor UO_1235 (O_1235,N_13647,N_14685);
nor UO_1236 (O_1236,N_14129,N_14350);
or UO_1237 (O_1237,N_14941,N_13536);
nand UO_1238 (O_1238,N_14971,N_14669);
and UO_1239 (O_1239,N_13656,N_13738);
or UO_1240 (O_1240,N_14564,N_13607);
and UO_1241 (O_1241,N_13609,N_13635);
nand UO_1242 (O_1242,N_14681,N_13817);
or UO_1243 (O_1243,N_13860,N_14715);
or UO_1244 (O_1244,N_14514,N_13855);
nand UO_1245 (O_1245,N_13813,N_14283);
nor UO_1246 (O_1246,N_14646,N_13872);
nor UO_1247 (O_1247,N_14150,N_14233);
nand UO_1248 (O_1248,N_14806,N_14328);
and UO_1249 (O_1249,N_14829,N_14648);
and UO_1250 (O_1250,N_14437,N_14481);
and UO_1251 (O_1251,N_14716,N_14757);
nand UO_1252 (O_1252,N_13973,N_13991);
or UO_1253 (O_1253,N_14216,N_14751);
and UO_1254 (O_1254,N_14794,N_13737);
or UO_1255 (O_1255,N_13640,N_14134);
nand UO_1256 (O_1256,N_14980,N_14011);
or UO_1257 (O_1257,N_14415,N_13692);
and UO_1258 (O_1258,N_14207,N_14849);
and UO_1259 (O_1259,N_14486,N_14777);
nor UO_1260 (O_1260,N_14740,N_13583);
nor UO_1261 (O_1261,N_14741,N_14803);
and UO_1262 (O_1262,N_13782,N_13901);
nand UO_1263 (O_1263,N_14634,N_14520);
and UO_1264 (O_1264,N_14896,N_14935);
or UO_1265 (O_1265,N_14732,N_14913);
nand UO_1266 (O_1266,N_14793,N_13980);
or UO_1267 (O_1267,N_14656,N_14951);
nor UO_1268 (O_1268,N_14061,N_14972);
nor UO_1269 (O_1269,N_14527,N_14007);
and UO_1270 (O_1270,N_14572,N_14254);
or UO_1271 (O_1271,N_14290,N_14280);
nand UO_1272 (O_1272,N_14448,N_14176);
and UO_1273 (O_1273,N_13854,N_13936);
nand UO_1274 (O_1274,N_13867,N_14961);
nor UO_1275 (O_1275,N_13692,N_14480);
nor UO_1276 (O_1276,N_14262,N_13865);
or UO_1277 (O_1277,N_14787,N_14237);
nand UO_1278 (O_1278,N_13509,N_14657);
or UO_1279 (O_1279,N_14416,N_13610);
or UO_1280 (O_1280,N_14980,N_14631);
or UO_1281 (O_1281,N_14554,N_14401);
nand UO_1282 (O_1282,N_13840,N_14907);
or UO_1283 (O_1283,N_13893,N_13781);
nor UO_1284 (O_1284,N_13817,N_13674);
nand UO_1285 (O_1285,N_13631,N_14020);
nand UO_1286 (O_1286,N_14691,N_14303);
or UO_1287 (O_1287,N_14088,N_14355);
nor UO_1288 (O_1288,N_13674,N_14097);
and UO_1289 (O_1289,N_13751,N_13709);
nor UO_1290 (O_1290,N_14915,N_13552);
or UO_1291 (O_1291,N_14716,N_14926);
nor UO_1292 (O_1292,N_13717,N_14458);
nor UO_1293 (O_1293,N_13662,N_14655);
nand UO_1294 (O_1294,N_13932,N_14405);
or UO_1295 (O_1295,N_13626,N_13911);
nand UO_1296 (O_1296,N_13688,N_14757);
nand UO_1297 (O_1297,N_14053,N_14002);
and UO_1298 (O_1298,N_14581,N_14908);
nor UO_1299 (O_1299,N_14073,N_13965);
and UO_1300 (O_1300,N_14073,N_14670);
nor UO_1301 (O_1301,N_14873,N_14454);
or UO_1302 (O_1302,N_14889,N_14016);
nor UO_1303 (O_1303,N_13589,N_13862);
or UO_1304 (O_1304,N_13962,N_14847);
or UO_1305 (O_1305,N_13617,N_13859);
nor UO_1306 (O_1306,N_14308,N_14583);
or UO_1307 (O_1307,N_14470,N_14610);
xor UO_1308 (O_1308,N_14763,N_14936);
or UO_1309 (O_1309,N_13634,N_14086);
and UO_1310 (O_1310,N_13526,N_14905);
or UO_1311 (O_1311,N_14632,N_14415);
and UO_1312 (O_1312,N_13659,N_13967);
and UO_1313 (O_1313,N_13769,N_13519);
nor UO_1314 (O_1314,N_14646,N_13909);
nand UO_1315 (O_1315,N_13935,N_14151);
nand UO_1316 (O_1316,N_13506,N_14640);
and UO_1317 (O_1317,N_14391,N_14643);
nor UO_1318 (O_1318,N_14760,N_13685);
and UO_1319 (O_1319,N_13666,N_14948);
nand UO_1320 (O_1320,N_14785,N_14471);
or UO_1321 (O_1321,N_13970,N_14088);
or UO_1322 (O_1322,N_14844,N_14042);
and UO_1323 (O_1323,N_14747,N_14438);
or UO_1324 (O_1324,N_14754,N_13964);
nand UO_1325 (O_1325,N_14694,N_13724);
and UO_1326 (O_1326,N_14860,N_14764);
nor UO_1327 (O_1327,N_14013,N_14575);
nand UO_1328 (O_1328,N_13673,N_13906);
and UO_1329 (O_1329,N_13737,N_14926);
xor UO_1330 (O_1330,N_14822,N_13756);
or UO_1331 (O_1331,N_14526,N_14470);
nand UO_1332 (O_1332,N_14428,N_14058);
nand UO_1333 (O_1333,N_13882,N_13686);
nor UO_1334 (O_1334,N_14254,N_13645);
or UO_1335 (O_1335,N_14853,N_14277);
or UO_1336 (O_1336,N_14037,N_14506);
nand UO_1337 (O_1337,N_14152,N_13929);
and UO_1338 (O_1338,N_14886,N_14413);
or UO_1339 (O_1339,N_14776,N_14544);
and UO_1340 (O_1340,N_14884,N_13754);
nor UO_1341 (O_1341,N_13887,N_13849);
nor UO_1342 (O_1342,N_14045,N_14914);
or UO_1343 (O_1343,N_14082,N_14924);
or UO_1344 (O_1344,N_13801,N_14179);
nand UO_1345 (O_1345,N_14470,N_14008);
or UO_1346 (O_1346,N_14784,N_14910);
and UO_1347 (O_1347,N_14258,N_14174);
nor UO_1348 (O_1348,N_14242,N_14409);
nor UO_1349 (O_1349,N_13511,N_13932);
or UO_1350 (O_1350,N_13806,N_14772);
or UO_1351 (O_1351,N_13589,N_13761);
nand UO_1352 (O_1352,N_13915,N_13539);
nand UO_1353 (O_1353,N_14507,N_14311);
or UO_1354 (O_1354,N_13825,N_14428);
nand UO_1355 (O_1355,N_14961,N_14149);
or UO_1356 (O_1356,N_13681,N_14133);
nor UO_1357 (O_1357,N_13716,N_14185);
and UO_1358 (O_1358,N_13907,N_14476);
nor UO_1359 (O_1359,N_14730,N_14066);
or UO_1360 (O_1360,N_13711,N_14039);
nor UO_1361 (O_1361,N_14637,N_14724);
and UO_1362 (O_1362,N_13760,N_13503);
and UO_1363 (O_1363,N_14752,N_14897);
and UO_1364 (O_1364,N_14189,N_14633);
and UO_1365 (O_1365,N_14412,N_13916);
or UO_1366 (O_1366,N_13944,N_14201);
and UO_1367 (O_1367,N_14927,N_13572);
and UO_1368 (O_1368,N_13821,N_13722);
nand UO_1369 (O_1369,N_13703,N_14337);
and UO_1370 (O_1370,N_13855,N_14523);
nand UO_1371 (O_1371,N_14129,N_13691);
nor UO_1372 (O_1372,N_14174,N_14883);
or UO_1373 (O_1373,N_13959,N_14857);
and UO_1374 (O_1374,N_14334,N_14894);
xor UO_1375 (O_1375,N_14481,N_13901);
or UO_1376 (O_1376,N_14454,N_14086);
and UO_1377 (O_1377,N_14033,N_13788);
and UO_1378 (O_1378,N_13915,N_13890);
nand UO_1379 (O_1379,N_14237,N_14261);
or UO_1380 (O_1380,N_14135,N_14453);
or UO_1381 (O_1381,N_13854,N_14203);
and UO_1382 (O_1382,N_14006,N_14444);
or UO_1383 (O_1383,N_13766,N_14793);
nor UO_1384 (O_1384,N_14832,N_13924);
and UO_1385 (O_1385,N_13898,N_13747);
nand UO_1386 (O_1386,N_13561,N_13848);
and UO_1387 (O_1387,N_14107,N_14954);
nand UO_1388 (O_1388,N_14612,N_13745);
or UO_1389 (O_1389,N_14013,N_14705);
and UO_1390 (O_1390,N_13583,N_13960);
or UO_1391 (O_1391,N_14888,N_14111);
nor UO_1392 (O_1392,N_13840,N_14848);
or UO_1393 (O_1393,N_14958,N_13873);
or UO_1394 (O_1394,N_14066,N_13512);
or UO_1395 (O_1395,N_14368,N_14978);
nand UO_1396 (O_1396,N_13745,N_13906);
nor UO_1397 (O_1397,N_14132,N_14270);
nor UO_1398 (O_1398,N_13743,N_13990);
nor UO_1399 (O_1399,N_14812,N_14570);
or UO_1400 (O_1400,N_14966,N_14013);
nor UO_1401 (O_1401,N_13743,N_14539);
nand UO_1402 (O_1402,N_14087,N_14735);
and UO_1403 (O_1403,N_14979,N_14409);
nor UO_1404 (O_1404,N_14790,N_13941);
or UO_1405 (O_1405,N_14372,N_14939);
or UO_1406 (O_1406,N_14600,N_14890);
nand UO_1407 (O_1407,N_13610,N_14138);
nor UO_1408 (O_1408,N_13788,N_14333);
and UO_1409 (O_1409,N_13979,N_13525);
nand UO_1410 (O_1410,N_14109,N_13563);
nor UO_1411 (O_1411,N_14154,N_13850);
or UO_1412 (O_1412,N_14759,N_13550);
and UO_1413 (O_1413,N_14998,N_13555);
nor UO_1414 (O_1414,N_13657,N_13982);
nand UO_1415 (O_1415,N_13685,N_14712);
or UO_1416 (O_1416,N_13941,N_14550);
or UO_1417 (O_1417,N_14035,N_13727);
or UO_1418 (O_1418,N_13672,N_14127);
nor UO_1419 (O_1419,N_14110,N_14198);
nor UO_1420 (O_1420,N_13664,N_13889);
or UO_1421 (O_1421,N_13578,N_14707);
nand UO_1422 (O_1422,N_14607,N_13722);
or UO_1423 (O_1423,N_14259,N_13990);
or UO_1424 (O_1424,N_13724,N_14799);
or UO_1425 (O_1425,N_13768,N_13855);
nand UO_1426 (O_1426,N_14782,N_13555);
nor UO_1427 (O_1427,N_13767,N_14640);
or UO_1428 (O_1428,N_13790,N_14896);
and UO_1429 (O_1429,N_14343,N_14232);
and UO_1430 (O_1430,N_13557,N_13963);
or UO_1431 (O_1431,N_14240,N_13941);
and UO_1432 (O_1432,N_13819,N_13787);
or UO_1433 (O_1433,N_13730,N_14523);
nand UO_1434 (O_1434,N_14997,N_13550);
or UO_1435 (O_1435,N_13963,N_14716);
or UO_1436 (O_1436,N_13620,N_13732);
and UO_1437 (O_1437,N_14768,N_14729);
nand UO_1438 (O_1438,N_14642,N_14205);
nor UO_1439 (O_1439,N_13993,N_14865);
nor UO_1440 (O_1440,N_14528,N_13984);
nor UO_1441 (O_1441,N_14868,N_14716);
nand UO_1442 (O_1442,N_14147,N_14018);
and UO_1443 (O_1443,N_14062,N_14212);
nor UO_1444 (O_1444,N_14097,N_14239);
and UO_1445 (O_1445,N_14684,N_13882);
or UO_1446 (O_1446,N_14704,N_13582);
nor UO_1447 (O_1447,N_13887,N_13926);
or UO_1448 (O_1448,N_14576,N_13835);
or UO_1449 (O_1449,N_14325,N_14394);
nor UO_1450 (O_1450,N_13704,N_14756);
nand UO_1451 (O_1451,N_14761,N_13575);
nor UO_1452 (O_1452,N_14060,N_13658);
and UO_1453 (O_1453,N_13835,N_13680);
and UO_1454 (O_1454,N_14118,N_14418);
nor UO_1455 (O_1455,N_14608,N_14198);
xnor UO_1456 (O_1456,N_13964,N_13949);
nand UO_1457 (O_1457,N_13573,N_14498);
nand UO_1458 (O_1458,N_14056,N_14709);
or UO_1459 (O_1459,N_14121,N_14422);
and UO_1460 (O_1460,N_14999,N_13808);
and UO_1461 (O_1461,N_14633,N_14833);
nor UO_1462 (O_1462,N_14943,N_14688);
and UO_1463 (O_1463,N_14711,N_14060);
nor UO_1464 (O_1464,N_14383,N_14654);
nand UO_1465 (O_1465,N_14352,N_14434);
nor UO_1466 (O_1466,N_14464,N_14322);
or UO_1467 (O_1467,N_14597,N_14113);
nand UO_1468 (O_1468,N_14400,N_13949);
nor UO_1469 (O_1469,N_13574,N_13772);
nor UO_1470 (O_1470,N_14839,N_14429);
and UO_1471 (O_1471,N_14186,N_14981);
nor UO_1472 (O_1472,N_14380,N_14000);
nor UO_1473 (O_1473,N_13756,N_14739);
or UO_1474 (O_1474,N_14571,N_13588);
or UO_1475 (O_1475,N_13970,N_14309);
nor UO_1476 (O_1476,N_13679,N_14285);
and UO_1477 (O_1477,N_13959,N_14132);
or UO_1478 (O_1478,N_13719,N_14119);
nand UO_1479 (O_1479,N_14094,N_13967);
nor UO_1480 (O_1480,N_14684,N_14977);
nand UO_1481 (O_1481,N_14854,N_13879);
nand UO_1482 (O_1482,N_14106,N_13612);
or UO_1483 (O_1483,N_13989,N_13883);
or UO_1484 (O_1484,N_13811,N_14174);
and UO_1485 (O_1485,N_13865,N_14995);
nor UO_1486 (O_1486,N_14391,N_14853);
or UO_1487 (O_1487,N_13589,N_14846);
or UO_1488 (O_1488,N_13878,N_14171);
and UO_1489 (O_1489,N_14618,N_14492);
or UO_1490 (O_1490,N_14056,N_13538);
nor UO_1491 (O_1491,N_14757,N_13915);
nor UO_1492 (O_1492,N_13789,N_13865);
nand UO_1493 (O_1493,N_14356,N_14373);
and UO_1494 (O_1494,N_14486,N_13888);
nand UO_1495 (O_1495,N_14252,N_14141);
and UO_1496 (O_1496,N_13845,N_14875);
nand UO_1497 (O_1497,N_14774,N_14784);
nor UO_1498 (O_1498,N_14996,N_14333);
nor UO_1499 (O_1499,N_13652,N_13944);
nor UO_1500 (O_1500,N_13992,N_14816);
nand UO_1501 (O_1501,N_13696,N_14062);
or UO_1502 (O_1502,N_13988,N_13920);
nor UO_1503 (O_1503,N_14067,N_14192);
and UO_1504 (O_1504,N_14668,N_14602);
nand UO_1505 (O_1505,N_14714,N_14703);
nand UO_1506 (O_1506,N_14244,N_13514);
nor UO_1507 (O_1507,N_14885,N_14011);
nor UO_1508 (O_1508,N_14698,N_14809);
nor UO_1509 (O_1509,N_13766,N_14674);
and UO_1510 (O_1510,N_14317,N_14810);
and UO_1511 (O_1511,N_13703,N_13976);
nor UO_1512 (O_1512,N_14783,N_14031);
nor UO_1513 (O_1513,N_13692,N_14363);
and UO_1514 (O_1514,N_14265,N_14168);
and UO_1515 (O_1515,N_14217,N_13767);
nor UO_1516 (O_1516,N_14504,N_14600);
nor UO_1517 (O_1517,N_13954,N_14975);
nand UO_1518 (O_1518,N_14610,N_13939);
or UO_1519 (O_1519,N_14870,N_14667);
nand UO_1520 (O_1520,N_14928,N_14111);
nand UO_1521 (O_1521,N_14096,N_14630);
nand UO_1522 (O_1522,N_14960,N_14945);
nand UO_1523 (O_1523,N_14599,N_14414);
or UO_1524 (O_1524,N_14773,N_14744);
or UO_1525 (O_1525,N_13939,N_14942);
and UO_1526 (O_1526,N_14532,N_14120);
nand UO_1527 (O_1527,N_13927,N_14242);
and UO_1528 (O_1528,N_13902,N_14847);
nor UO_1529 (O_1529,N_14041,N_14699);
nand UO_1530 (O_1530,N_14733,N_14545);
nand UO_1531 (O_1531,N_14954,N_14121);
nand UO_1532 (O_1532,N_13689,N_14376);
nand UO_1533 (O_1533,N_14579,N_13548);
or UO_1534 (O_1534,N_14250,N_13550);
nor UO_1535 (O_1535,N_14951,N_14474);
nand UO_1536 (O_1536,N_13703,N_13602);
nor UO_1537 (O_1537,N_14036,N_13767);
or UO_1538 (O_1538,N_13628,N_13678);
and UO_1539 (O_1539,N_14060,N_13623);
or UO_1540 (O_1540,N_14542,N_14056);
nand UO_1541 (O_1541,N_14832,N_13772);
or UO_1542 (O_1542,N_13705,N_13939);
and UO_1543 (O_1543,N_14163,N_13747);
or UO_1544 (O_1544,N_13667,N_13899);
or UO_1545 (O_1545,N_14228,N_14682);
and UO_1546 (O_1546,N_14226,N_14848);
or UO_1547 (O_1547,N_14418,N_14296);
and UO_1548 (O_1548,N_14978,N_13802);
or UO_1549 (O_1549,N_13873,N_14416);
or UO_1550 (O_1550,N_14163,N_13759);
and UO_1551 (O_1551,N_14565,N_14135);
nor UO_1552 (O_1552,N_14595,N_13751);
nor UO_1553 (O_1553,N_14263,N_14344);
and UO_1554 (O_1554,N_13951,N_14292);
and UO_1555 (O_1555,N_14456,N_13551);
nor UO_1556 (O_1556,N_14732,N_14571);
or UO_1557 (O_1557,N_14875,N_14823);
or UO_1558 (O_1558,N_14507,N_13988);
or UO_1559 (O_1559,N_13718,N_14115);
nand UO_1560 (O_1560,N_14450,N_14190);
nor UO_1561 (O_1561,N_13909,N_14575);
or UO_1562 (O_1562,N_14982,N_14517);
or UO_1563 (O_1563,N_14974,N_13726);
nand UO_1564 (O_1564,N_14468,N_14289);
nand UO_1565 (O_1565,N_13704,N_14069);
or UO_1566 (O_1566,N_13876,N_14030);
or UO_1567 (O_1567,N_14869,N_13994);
and UO_1568 (O_1568,N_14345,N_13870);
nor UO_1569 (O_1569,N_13522,N_14770);
nand UO_1570 (O_1570,N_13634,N_13546);
or UO_1571 (O_1571,N_14093,N_13793);
nor UO_1572 (O_1572,N_14880,N_13757);
nor UO_1573 (O_1573,N_14199,N_14270);
and UO_1574 (O_1574,N_14385,N_14052);
and UO_1575 (O_1575,N_13912,N_14394);
nand UO_1576 (O_1576,N_14107,N_14699);
nor UO_1577 (O_1577,N_14382,N_13773);
and UO_1578 (O_1578,N_13792,N_14218);
nor UO_1579 (O_1579,N_14122,N_14370);
nand UO_1580 (O_1580,N_13672,N_13934);
nand UO_1581 (O_1581,N_14580,N_14759);
nand UO_1582 (O_1582,N_14122,N_14367);
nor UO_1583 (O_1583,N_14635,N_14297);
or UO_1584 (O_1584,N_13588,N_14717);
nor UO_1585 (O_1585,N_14779,N_13573);
or UO_1586 (O_1586,N_13658,N_14979);
nor UO_1587 (O_1587,N_13876,N_14750);
nor UO_1588 (O_1588,N_13773,N_14123);
and UO_1589 (O_1589,N_13943,N_13517);
or UO_1590 (O_1590,N_14475,N_14073);
or UO_1591 (O_1591,N_13930,N_13556);
nand UO_1592 (O_1592,N_13930,N_14331);
or UO_1593 (O_1593,N_14794,N_13853);
nor UO_1594 (O_1594,N_13607,N_13979);
and UO_1595 (O_1595,N_14498,N_14045);
nor UO_1596 (O_1596,N_13668,N_14625);
nor UO_1597 (O_1597,N_14523,N_13633);
or UO_1598 (O_1598,N_14778,N_13812);
nor UO_1599 (O_1599,N_14982,N_13690);
or UO_1600 (O_1600,N_14188,N_14176);
and UO_1601 (O_1601,N_14882,N_14963);
or UO_1602 (O_1602,N_13617,N_14842);
nand UO_1603 (O_1603,N_14080,N_14167);
nand UO_1604 (O_1604,N_14751,N_13849);
nor UO_1605 (O_1605,N_13930,N_14944);
nand UO_1606 (O_1606,N_13616,N_13971);
nand UO_1607 (O_1607,N_14130,N_14689);
nor UO_1608 (O_1608,N_14671,N_13792);
and UO_1609 (O_1609,N_14359,N_13719);
or UO_1610 (O_1610,N_14809,N_14203);
and UO_1611 (O_1611,N_14101,N_14301);
nand UO_1612 (O_1612,N_13688,N_14279);
nand UO_1613 (O_1613,N_14082,N_14774);
nand UO_1614 (O_1614,N_14022,N_13850);
or UO_1615 (O_1615,N_14266,N_14230);
or UO_1616 (O_1616,N_13782,N_14590);
and UO_1617 (O_1617,N_14961,N_14732);
nand UO_1618 (O_1618,N_14152,N_14517);
nand UO_1619 (O_1619,N_14964,N_13929);
nor UO_1620 (O_1620,N_13821,N_13999);
nor UO_1621 (O_1621,N_14832,N_14208);
nand UO_1622 (O_1622,N_14680,N_14786);
nor UO_1623 (O_1623,N_14851,N_13549);
or UO_1624 (O_1624,N_13759,N_14125);
nor UO_1625 (O_1625,N_14365,N_14273);
or UO_1626 (O_1626,N_13668,N_14480);
and UO_1627 (O_1627,N_13777,N_13648);
or UO_1628 (O_1628,N_14646,N_13988);
or UO_1629 (O_1629,N_14431,N_13786);
or UO_1630 (O_1630,N_14829,N_14197);
nor UO_1631 (O_1631,N_14999,N_13976);
nor UO_1632 (O_1632,N_13782,N_14246);
nor UO_1633 (O_1633,N_14519,N_14184);
and UO_1634 (O_1634,N_13527,N_14709);
or UO_1635 (O_1635,N_14551,N_14138);
nor UO_1636 (O_1636,N_14518,N_13502);
nand UO_1637 (O_1637,N_13874,N_14239);
nand UO_1638 (O_1638,N_14485,N_14576);
nor UO_1639 (O_1639,N_14509,N_14918);
nor UO_1640 (O_1640,N_14632,N_13670);
nand UO_1641 (O_1641,N_14839,N_14335);
nand UO_1642 (O_1642,N_13683,N_14563);
and UO_1643 (O_1643,N_14804,N_14043);
nand UO_1644 (O_1644,N_14238,N_14845);
nor UO_1645 (O_1645,N_13511,N_13649);
nand UO_1646 (O_1646,N_14246,N_14844);
and UO_1647 (O_1647,N_14361,N_13713);
and UO_1648 (O_1648,N_14995,N_14913);
and UO_1649 (O_1649,N_13652,N_13890);
or UO_1650 (O_1650,N_14579,N_14093);
or UO_1651 (O_1651,N_14072,N_13797);
and UO_1652 (O_1652,N_13865,N_13734);
nand UO_1653 (O_1653,N_14455,N_13781);
nor UO_1654 (O_1654,N_13601,N_14641);
nor UO_1655 (O_1655,N_14578,N_14301);
nor UO_1656 (O_1656,N_14782,N_13596);
nor UO_1657 (O_1657,N_13984,N_14011);
nor UO_1658 (O_1658,N_14906,N_14378);
nor UO_1659 (O_1659,N_13597,N_14606);
or UO_1660 (O_1660,N_14580,N_14464);
or UO_1661 (O_1661,N_13627,N_14680);
nand UO_1662 (O_1662,N_14351,N_14893);
and UO_1663 (O_1663,N_14925,N_14406);
nand UO_1664 (O_1664,N_13863,N_13796);
and UO_1665 (O_1665,N_14965,N_14642);
or UO_1666 (O_1666,N_14675,N_13862);
nand UO_1667 (O_1667,N_14013,N_14315);
and UO_1668 (O_1668,N_14389,N_14057);
nor UO_1669 (O_1669,N_14891,N_14066);
nand UO_1670 (O_1670,N_14942,N_14907);
and UO_1671 (O_1671,N_13646,N_14852);
nand UO_1672 (O_1672,N_14782,N_14309);
nor UO_1673 (O_1673,N_13911,N_13838);
nand UO_1674 (O_1674,N_14113,N_13977);
or UO_1675 (O_1675,N_14542,N_13987);
and UO_1676 (O_1676,N_13551,N_14012);
nor UO_1677 (O_1677,N_13740,N_13505);
and UO_1678 (O_1678,N_13635,N_14369);
nand UO_1679 (O_1679,N_14626,N_14215);
and UO_1680 (O_1680,N_13784,N_14469);
and UO_1681 (O_1681,N_14959,N_14729);
nand UO_1682 (O_1682,N_14158,N_14938);
and UO_1683 (O_1683,N_13618,N_14913);
nand UO_1684 (O_1684,N_13842,N_14344);
nor UO_1685 (O_1685,N_14037,N_14868);
and UO_1686 (O_1686,N_14947,N_13500);
and UO_1687 (O_1687,N_13668,N_13547);
or UO_1688 (O_1688,N_14913,N_14954);
nor UO_1689 (O_1689,N_14385,N_14108);
xor UO_1690 (O_1690,N_13974,N_14929);
nor UO_1691 (O_1691,N_14088,N_14226);
and UO_1692 (O_1692,N_13532,N_13894);
and UO_1693 (O_1693,N_14094,N_14037);
or UO_1694 (O_1694,N_13769,N_13716);
and UO_1695 (O_1695,N_13632,N_14571);
xnor UO_1696 (O_1696,N_14477,N_13614);
and UO_1697 (O_1697,N_14150,N_14366);
and UO_1698 (O_1698,N_14939,N_14643);
nand UO_1699 (O_1699,N_14352,N_13839);
and UO_1700 (O_1700,N_13989,N_14019);
nand UO_1701 (O_1701,N_14560,N_13661);
nand UO_1702 (O_1702,N_13575,N_13687);
and UO_1703 (O_1703,N_14450,N_14699);
and UO_1704 (O_1704,N_13556,N_13644);
and UO_1705 (O_1705,N_13621,N_14468);
or UO_1706 (O_1706,N_14612,N_13635);
or UO_1707 (O_1707,N_13807,N_14031);
nor UO_1708 (O_1708,N_14759,N_13909);
nand UO_1709 (O_1709,N_13942,N_13540);
and UO_1710 (O_1710,N_14472,N_13715);
or UO_1711 (O_1711,N_14322,N_14039);
and UO_1712 (O_1712,N_14541,N_14779);
and UO_1713 (O_1713,N_14150,N_13854);
and UO_1714 (O_1714,N_14578,N_13792);
nor UO_1715 (O_1715,N_14080,N_13927);
nor UO_1716 (O_1716,N_13878,N_14107);
and UO_1717 (O_1717,N_14354,N_13591);
and UO_1718 (O_1718,N_14138,N_14387);
nand UO_1719 (O_1719,N_14781,N_14629);
nand UO_1720 (O_1720,N_13763,N_13788);
nand UO_1721 (O_1721,N_14662,N_14936);
nor UO_1722 (O_1722,N_13752,N_14962);
or UO_1723 (O_1723,N_13503,N_14891);
nand UO_1724 (O_1724,N_14457,N_13712);
or UO_1725 (O_1725,N_14844,N_14374);
nor UO_1726 (O_1726,N_13727,N_14834);
or UO_1727 (O_1727,N_13807,N_13829);
or UO_1728 (O_1728,N_14919,N_14964);
or UO_1729 (O_1729,N_13798,N_13796);
and UO_1730 (O_1730,N_14380,N_13644);
nor UO_1731 (O_1731,N_13538,N_14735);
nor UO_1732 (O_1732,N_14482,N_14583);
or UO_1733 (O_1733,N_14444,N_14176);
nand UO_1734 (O_1734,N_14614,N_14475);
and UO_1735 (O_1735,N_13950,N_13852);
or UO_1736 (O_1736,N_13635,N_13947);
and UO_1737 (O_1737,N_13706,N_14778);
and UO_1738 (O_1738,N_14172,N_13718);
and UO_1739 (O_1739,N_14549,N_14919);
and UO_1740 (O_1740,N_14955,N_14082);
xor UO_1741 (O_1741,N_14937,N_13609);
and UO_1742 (O_1742,N_14921,N_14538);
nor UO_1743 (O_1743,N_13808,N_14512);
nor UO_1744 (O_1744,N_14326,N_14944);
and UO_1745 (O_1745,N_13750,N_14951);
and UO_1746 (O_1746,N_14720,N_14783);
nor UO_1747 (O_1747,N_14450,N_14542);
and UO_1748 (O_1748,N_14648,N_14327);
nor UO_1749 (O_1749,N_14951,N_14042);
or UO_1750 (O_1750,N_14235,N_14236);
or UO_1751 (O_1751,N_14300,N_13607);
nor UO_1752 (O_1752,N_14975,N_14024);
and UO_1753 (O_1753,N_13604,N_13611);
and UO_1754 (O_1754,N_13925,N_14061);
xnor UO_1755 (O_1755,N_14378,N_14900);
and UO_1756 (O_1756,N_13889,N_13954);
nand UO_1757 (O_1757,N_13507,N_13760);
nor UO_1758 (O_1758,N_13853,N_14755);
and UO_1759 (O_1759,N_14872,N_13714);
and UO_1760 (O_1760,N_14739,N_13868);
nor UO_1761 (O_1761,N_14745,N_13814);
or UO_1762 (O_1762,N_14305,N_13686);
or UO_1763 (O_1763,N_14399,N_13905);
and UO_1764 (O_1764,N_14912,N_14610);
or UO_1765 (O_1765,N_14344,N_13710);
nand UO_1766 (O_1766,N_13643,N_13841);
nor UO_1767 (O_1767,N_13707,N_13701);
xor UO_1768 (O_1768,N_14090,N_14977);
or UO_1769 (O_1769,N_13718,N_14283);
xor UO_1770 (O_1770,N_14118,N_14998);
nor UO_1771 (O_1771,N_13589,N_14995);
and UO_1772 (O_1772,N_13886,N_14850);
nor UO_1773 (O_1773,N_14523,N_14889);
nor UO_1774 (O_1774,N_13970,N_13551);
nor UO_1775 (O_1775,N_13985,N_14246);
nand UO_1776 (O_1776,N_13607,N_13708);
nand UO_1777 (O_1777,N_14757,N_13800);
nor UO_1778 (O_1778,N_14254,N_13948);
and UO_1779 (O_1779,N_14561,N_14976);
or UO_1780 (O_1780,N_13800,N_13930);
nor UO_1781 (O_1781,N_14618,N_14473);
and UO_1782 (O_1782,N_13954,N_14996);
or UO_1783 (O_1783,N_13645,N_13942);
nor UO_1784 (O_1784,N_14338,N_14170);
nor UO_1785 (O_1785,N_13948,N_14356);
nand UO_1786 (O_1786,N_14615,N_14949);
or UO_1787 (O_1787,N_14669,N_14535);
xnor UO_1788 (O_1788,N_13687,N_13943);
nor UO_1789 (O_1789,N_13898,N_14312);
nand UO_1790 (O_1790,N_14236,N_14209);
or UO_1791 (O_1791,N_14287,N_13702);
or UO_1792 (O_1792,N_14202,N_14293);
nor UO_1793 (O_1793,N_14449,N_13682);
nand UO_1794 (O_1794,N_14265,N_13823);
nor UO_1795 (O_1795,N_14652,N_14747);
or UO_1796 (O_1796,N_14122,N_13826);
nor UO_1797 (O_1797,N_13536,N_14089);
nand UO_1798 (O_1798,N_14219,N_14450);
or UO_1799 (O_1799,N_13649,N_14914);
nor UO_1800 (O_1800,N_13828,N_14419);
nor UO_1801 (O_1801,N_14796,N_13799);
and UO_1802 (O_1802,N_14297,N_14803);
nor UO_1803 (O_1803,N_14341,N_13733);
or UO_1804 (O_1804,N_14874,N_14900);
and UO_1805 (O_1805,N_14084,N_13543);
or UO_1806 (O_1806,N_14672,N_14504);
nand UO_1807 (O_1807,N_14655,N_14127);
nand UO_1808 (O_1808,N_13510,N_14113);
or UO_1809 (O_1809,N_14008,N_14858);
and UO_1810 (O_1810,N_13984,N_14592);
nor UO_1811 (O_1811,N_14282,N_14247);
or UO_1812 (O_1812,N_14589,N_14156);
nand UO_1813 (O_1813,N_14706,N_13555);
or UO_1814 (O_1814,N_13908,N_14023);
and UO_1815 (O_1815,N_13755,N_14687);
nand UO_1816 (O_1816,N_13788,N_14364);
and UO_1817 (O_1817,N_13976,N_14632);
nor UO_1818 (O_1818,N_13886,N_13539);
nand UO_1819 (O_1819,N_14877,N_14848);
nand UO_1820 (O_1820,N_13756,N_13987);
nand UO_1821 (O_1821,N_14312,N_14168);
xnor UO_1822 (O_1822,N_13767,N_14042);
or UO_1823 (O_1823,N_14595,N_13870);
and UO_1824 (O_1824,N_14924,N_13550);
and UO_1825 (O_1825,N_13826,N_14704);
or UO_1826 (O_1826,N_14877,N_14852);
and UO_1827 (O_1827,N_13993,N_14947);
or UO_1828 (O_1828,N_13524,N_14139);
and UO_1829 (O_1829,N_14085,N_14012);
and UO_1830 (O_1830,N_14921,N_14909);
and UO_1831 (O_1831,N_13888,N_14907);
nand UO_1832 (O_1832,N_13632,N_14699);
nand UO_1833 (O_1833,N_14737,N_13551);
and UO_1834 (O_1834,N_13575,N_14709);
or UO_1835 (O_1835,N_13706,N_13850);
and UO_1836 (O_1836,N_14412,N_14495);
nand UO_1837 (O_1837,N_14481,N_13563);
nor UO_1838 (O_1838,N_14738,N_14991);
nor UO_1839 (O_1839,N_14909,N_13863);
and UO_1840 (O_1840,N_13616,N_13900);
or UO_1841 (O_1841,N_13794,N_14759);
and UO_1842 (O_1842,N_13830,N_14002);
nor UO_1843 (O_1843,N_13817,N_14787);
nor UO_1844 (O_1844,N_14381,N_13582);
or UO_1845 (O_1845,N_14034,N_14894);
nand UO_1846 (O_1846,N_14493,N_14834);
nand UO_1847 (O_1847,N_13760,N_14395);
or UO_1848 (O_1848,N_14565,N_13899);
or UO_1849 (O_1849,N_14736,N_13706);
nor UO_1850 (O_1850,N_14820,N_14703);
or UO_1851 (O_1851,N_14339,N_13818);
nand UO_1852 (O_1852,N_14227,N_13512);
nand UO_1853 (O_1853,N_14505,N_14434);
or UO_1854 (O_1854,N_14835,N_14395);
nand UO_1855 (O_1855,N_14591,N_13513);
nand UO_1856 (O_1856,N_14586,N_14652);
or UO_1857 (O_1857,N_14982,N_14771);
nand UO_1858 (O_1858,N_14946,N_13564);
nand UO_1859 (O_1859,N_14127,N_14639);
and UO_1860 (O_1860,N_14606,N_13571);
nor UO_1861 (O_1861,N_13897,N_13857);
nor UO_1862 (O_1862,N_14739,N_13547);
or UO_1863 (O_1863,N_14761,N_13643);
nor UO_1864 (O_1864,N_13804,N_14574);
nor UO_1865 (O_1865,N_13621,N_14187);
and UO_1866 (O_1866,N_14645,N_14888);
or UO_1867 (O_1867,N_13607,N_14551);
nand UO_1868 (O_1868,N_13853,N_14236);
or UO_1869 (O_1869,N_14938,N_13645);
nor UO_1870 (O_1870,N_14635,N_13679);
or UO_1871 (O_1871,N_14708,N_14470);
or UO_1872 (O_1872,N_13633,N_14246);
nor UO_1873 (O_1873,N_13789,N_14311);
nand UO_1874 (O_1874,N_13924,N_13927);
nand UO_1875 (O_1875,N_14164,N_13727);
nor UO_1876 (O_1876,N_14934,N_14585);
nor UO_1877 (O_1877,N_14904,N_14272);
and UO_1878 (O_1878,N_14983,N_13619);
and UO_1879 (O_1879,N_14715,N_13641);
nand UO_1880 (O_1880,N_13532,N_14881);
and UO_1881 (O_1881,N_14121,N_14851);
or UO_1882 (O_1882,N_14917,N_14808);
and UO_1883 (O_1883,N_14105,N_13509);
or UO_1884 (O_1884,N_14303,N_14652);
xnor UO_1885 (O_1885,N_14334,N_14367);
nor UO_1886 (O_1886,N_13945,N_14555);
nor UO_1887 (O_1887,N_14768,N_14016);
nor UO_1888 (O_1888,N_14885,N_14936);
xor UO_1889 (O_1889,N_14995,N_14926);
nor UO_1890 (O_1890,N_14835,N_13946);
nand UO_1891 (O_1891,N_14157,N_13983);
or UO_1892 (O_1892,N_13881,N_14220);
nand UO_1893 (O_1893,N_14050,N_13702);
nor UO_1894 (O_1894,N_13924,N_14933);
nand UO_1895 (O_1895,N_13721,N_13791);
nor UO_1896 (O_1896,N_13698,N_14699);
nand UO_1897 (O_1897,N_14762,N_14544);
nor UO_1898 (O_1898,N_14946,N_13695);
nor UO_1899 (O_1899,N_14286,N_13729);
nor UO_1900 (O_1900,N_14331,N_13961);
nor UO_1901 (O_1901,N_14604,N_14336);
and UO_1902 (O_1902,N_14432,N_14204);
and UO_1903 (O_1903,N_13971,N_14945);
and UO_1904 (O_1904,N_14806,N_14556);
or UO_1905 (O_1905,N_14372,N_13627);
or UO_1906 (O_1906,N_14696,N_14064);
nor UO_1907 (O_1907,N_14180,N_14016);
and UO_1908 (O_1908,N_14663,N_13955);
nand UO_1909 (O_1909,N_14194,N_14418);
or UO_1910 (O_1910,N_14110,N_13748);
and UO_1911 (O_1911,N_14969,N_13504);
nor UO_1912 (O_1912,N_14689,N_13570);
and UO_1913 (O_1913,N_14436,N_14353);
nand UO_1914 (O_1914,N_13631,N_14305);
nand UO_1915 (O_1915,N_13546,N_13729);
xnor UO_1916 (O_1916,N_14268,N_13818);
and UO_1917 (O_1917,N_14843,N_13574);
and UO_1918 (O_1918,N_14886,N_14542);
nand UO_1919 (O_1919,N_13958,N_14353);
nor UO_1920 (O_1920,N_13942,N_14471);
and UO_1921 (O_1921,N_14731,N_14618);
or UO_1922 (O_1922,N_14897,N_14053);
and UO_1923 (O_1923,N_13649,N_13930);
nand UO_1924 (O_1924,N_14814,N_13757);
nand UO_1925 (O_1925,N_14980,N_14823);
and UO_1926 (O_1926,N_13643,N_14923);
nor UO_1927 (O_1927,N_14963,N_14524);
and UO_1928 (O_1928,N_13835,N_13568);
and UO_1929 (O_1929,N_14350,N_13875);
nand UO_1930 (O_1930,N_14023,N_14328);
and UO_1931 (O_1931,N_13824,N_14814);
nor UO_1932 (O_1932,N_13951,N_14421);
nand UO_1933 (O_1933,N_14292,N_14649);
nand UO_1934 (O_1934,N_14815,N_14641);
nor UO_1935 (O_1935,N_13758,N_13551);
nand UO_1936 (O_1936,N_13898,N_14939);
or UO_1937 (O_1937,N_14550,N_14871);
and UO_1938 (O_1938,N_14279,N_14667);
nor UO_1939 (O_1939,N_14789,N_14111);
nand UO_1940 (O_1940,N_13850,N_14390);
or UO_1941 (O_1941,N_14504,N_14459);
nor UO_1942 (O_1942,N_13739,N_13943);
nor UO_1943 (O_1943,N_14450,N_14976);
or UO_1944 (O_1944,N_14037,N_14234);
or UO_1945 (O_1945,N_14738,N_14312);
nor UO_1946 (O_1946,N_13714,N_14183);
nor UO_1947 (O_1947,N_14537,N_14089);
nor UO_1948 (O_1948,N_13719,N_14399);
or UO_1949 (O_1949,N_14923,N_14458);
xnor UO_1950 (O_1950,N_13546,N_14988);
nand UO_1951 (O_1951,N_13752,N_13621);
nand UO_1952 (O_1952,N_14016,N_14356);
nor UO_1953 (O_1953,N_14783,N_13964);
nor UO_1954 (O_1954,N_14415,N_13663);
nand UO_1955 (O_1955,N_14321,N_14606);
or UO_1956 (O_1956,N_13883,N_13906);
nor UO_1957 (O_1957,N_13850,N_14565);
or UO_1958 (O_1958,N_14705,N_13570);
and UO_1959 (O_1959,N_13547,N_14930);
and UO_1960 (O_1960,N_13537,N_13974);
nand UO_1961 (O_1961,N_14070,N_14347);
nand UO_1962 (O_1962,N_14970,N_14362);
nor UO_1963 (O_1963,N_14843,N_14667);
and UO_1964 (O_1964,N_13682,N_14748);
nand UO_1965 (O_1965,N_13626,N_14751);
and UO_1966 (O_1966,N_14258,N_14595);
nand UO_1967 (O_1967,N_14005,N_14161);
and UO_1968 (O_1968,N_13624,N_13887);
or UO_1969 (O_1969,N_13998,N_14453);
nand UO_1970 (O_1970,N_14066,N_14882);
and UO_1971 (O_1971,N_14198,N_14107);
or UO_1972 (O_1972,N_14904,N_14794);
or UO_1973 (O_1973,N_14858,N_14759);
and UO_1974 (O_1974,N_13503,N_13534);
nand UO_1975 (O_1975,N_14913,N_14971);
or UO_1976 (O_1976,N_14518,N_14541);
nand UO_1977 (O_1977,N_13571,N_13569);
or UO_1978 (O_1978,N_13667,N_14802);
nand UO_1979 (O_1979,N_14760,N_14087);
and UO_1980 (O_1980,N_13702,N_14796);
and UO_1981 (O_1981,N_14889,N_13925);
nand UO_1982 (O_1982,N_14184,N_14628);
and UO_1983 (O_1983,N_14626,N_13595);
or UO_1984 (O_1984,N_14237,N_14612);
or UO_1985 (O_1985,N_13517,N_14446);
nand UO_1986 (O_1986,N_13714,N_13716);
or UO_1987 (O_1987,N_13726,N_13724);
and UO_1988 (O_1988,N_14247,N_14879);
nand UO_1989 (O_1989,N_13767,N_14413);
and UO_1990 (O_1990,N_13675,N_14750);
and UO_1991 (O_1991,N_13735,N_14504);
nand UO_1992 (O_1992,N_13840,N_13635);
nor UO_1993 (O_1993,N_14409,N_13547);
nor UO_1994 (O_1994,N_13802,N_13887);
or UO_1995 (O_1995,N_14535,N_14788);
and UO_1996 (O_1996,N_13995,N_14530);
or UO_1997 (O_1997,N_14810,N_13593);
and UO_1998 (O_1998,N_13925,N_13798);
nand UO_1999 (O_1999,N_13527,N_14074);
endmodule