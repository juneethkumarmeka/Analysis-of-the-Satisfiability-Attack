module basic_5000_50000_5000_20_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_3113,In_797);
xor U1 (N_1,In_4236,In_1827);
or U2 (N_2,In_2811,In_211);
nand U3 (N_3,In_2444,In_847);
or U4 (N_4,In_379,In_908);
and U5 (N_5,In_3732,In_2001);
nand U6 (N_6,In_1906,In_1517);
nor U7 (N_7,In_1301,In_2504);
nor U8 (N_8,In_250,In_538);
nand U9 (N_9,In_1210,In_2961);
nor U10 (N_10,In_1936,In_3670);
nor U11 (N_11,In_3584,In_2766);
or U12 (N_12,In_2835,In_1529);
and U13 (N_13,In_785,In_4561);
xor U14 (N_14,In_4713,In_629);
or U15 (N_15,In_647,In_3734);
nand U16 (N_16,In_436,In_4565);
nand U17 (N_17,In_968,In_4690);
nand U18 (N_18,In_3335,In_3103);
xnor U19 (N_19,In_4364,In_1180);
nor U20 (N_20,In_4137,In_3737);
and U21 (N_21,In_525,In_2119);
nor U22 (N_22,In_1648,In_4042);
nand U23 (N_23,In_4608,In_4738);
xnor U24 (N_24,In_2344,In_4095);
or U25 (N_25,In_1119,In_2026);
or U26 (N_26,In_4186,In_2863);
nand U27 (N_27,In_2977,In_2713);
nor U28 (N_28,In_77,In_3470);
xnor U29 (N_29,In_425,In_2490);
nor U30 (N_30,In_511,In_2902);
nand U31 (N_31,In_1359,In_3169);
nor U32 (N_32,In_2017,In_1397);
nor U33 (N_33,In_2030,In_1787);
and U34 (N_34,In_2892,In_1866);
and U35 (N_35,In_1786,In_12);
and U36 (N_36,In_4058,In_1950);
and U37 (N_37,In_4409,In_2183);
xnor U38 (N_38,In_596,In_626);
or U39 (N_39,In_4056,In_3133);
xnor U40 (N_40,In_1942,In_249);
and U41 (N_41,In_1158,In_943);
nand U42 (N_42,In_3746,In_4488);
nor U43 (N_43,In_4864,In_4383);
xor U44 (N_44,In_3539,In_307);
and U45 (N_45,In_3339,In_2452);
nand U46 (N_46,In_328,In_3134);
and U47 (N_47,In_3475,In_2709);
nand U48 (N_48,In_2635,In_1524);
nand U49 (N_49,In_1033,In_813);
xnor U50 (N_50,In_4019,In_4792);
or U51 (N_51,In_3241,In_566);
nor U52 (N_52,In_1393,In_4707);
xor U53 (N_53,In_2919,In_2669);
nand U54 (N_54,In_1252,In_3625);
xnor U55 (N_55,In_197,In_4408);
xor U56 (N_56,In_3985,In_3177);
xnor U57 (N_57,In_979,In_3557);
nand U58 (N_58,In_1740,In_4572);
or U59 (N_59,In_3765,In_3333);
xnor U60 (N_60,In_385,In_401);
or U61 (N_61,In_903,In_2272);
nor U62 (N_62,In_627,In_1017);
and U63 (N_63,In_164,In_4845);
xnor U64 (N_64,In_1184,In_1098);
or U65 (N_65,In_3243,In_3917);
nand U66 (N_66,In_863,In_196);
nor U67 (N_67,In_3847,In_2787);
nand U68 (N_68,In_2665,In_192);
nor U69 (N_69,In_3118,In_4104);
nor U70 (N_70,In_4138,In_3364);
or U71 (N_71,In_2071,In_3190);
nand U72 (N_72,In_4793,In_2630);
xor U73 (N_73,In_3180,In_2899);
and U74 (N_74,In_1586,In_1658);
or U75 (N_75,In_1910,In_608);
nor U76 (N_76,In_235,In_2620);
nor U77 (N_77,In_4836,In_239);
and U78 (N_78,In_3690,In_3480);
nor U79 (N_79,In_2756,In_4703);
nand U80 (N_80,In_3669,In_218);
nor U81 (N_81,In_3037,In_2844);
xnor U82 (N_82,In_4813,In_1046);
or U83 (N_83,In_1028,In_4317);
and U84 (N_84,In_309,In_4988);
nor U85 (N_85,In_3941,In_3387);
or U86 (N_86,In_1746,In_1433);
nor U87 (N_87,In_68,In_4552);
nor U88 (N_88,In_4979,In_3075);
or U89 (N_89,In_4729,In_3189);
or U90 (N_90,In_1166,In_1702);
nand U91 (N_91,In_4045,In_2690);
nand U92 (N_92,In_1706,In_1582);
nand U93 (N_93,In_4772,In_1381);
nor U94 (N_94,In_4180,In_3081);
nor U95 (N_95,In_3990,In_4627);
nand U96 (N_96,In_3864,In_4351);
and U97 (N_97,In_2232,In_2430);
or U98 (N_98,In_1760,In_2423);
nand U99 (N_99,In_4966,In_3157);
and U100 (N_100,In_257,In_1010);
nor U101 (N_101,In_3451,In_1840);
nand U102 (N_102,In_4606,In_2805);
or U103 (N_103,In_1984,In_1789);
nand U104 (N_104,In_3022,In_4723);
or U105 (N_105,In_3378,In_2261);
or U106 (N_106,In_2162,In_3083);
nor U107 (N_107,In_4304,In_1135);
nand U108 (N_108,In_2707,In_1070);
or U109 (N_109,In_1430,In_4298);
nand U110 (N_110,In_2985,In_4008);
nor U111 (N_111,In_2900,In_712);
and U112 (N_112,In_1928,In_2334);
or U113 (N_113,In_1552,In_2930);
nand U114 (N_114,In_156,In_135);
and U115 (N_115,In_4136,In_1303);
xor U116 (N_116,In_1431,In_2600);
nand U117 (N_117,In_1891,In_773);
nand U118 (N_118,In_4101,In_555);
xnor U119 (N_119,In_4615,In_2851);
or U120 (N_120,In_2447,In_3640);
and U121 (N_121,In_3846,In_3982);
or U122 (N_122,In_3913,In_4512);
nor U123 (N_123,In_3162,In_1632);
nor U124 (N_124,In_1687,In_2385);
nand U125 (N_125,In_1131,In_4296);
nand U126 (N_126,In_1076,In_4425);
nor U127 (N_127,In_3306,In_808);
nand U128 (N_128,In_3761,In_646);
nand U129 (N_129,In_3459,In_4957);
nand U130 (N_130,In_3199,In_174);
nand U131 (N_131,In_3977,In_4821);
or U132 (N_132,In_973,In_747);
xor U133 (N_133,In_2159,In_879);
xnor U134 (N_134,In_910,In_2857);
nor U135 (N_135,In_3135,In_206);
nor U136 (N_136,In_2876,In_2443);
or U137 (N_137,In_3659,In_2538);
or U138 (N_138,In_1683,In_3676);
or U139 (N_139,In_2582,In_3918);
nor U140 (N_140,In_3267,In_838);
nand U141 (N_141,In_1515,In_490);
xnor U142 (N_142,In_3963,In_4519);
xor U143 (N_143,In_2056,In_1653);
xor U144 (N_144,In_2998,In_243);
nor U145 (N_145,In_1148,In_2924);
xnor U146 (N_146,In_119,In_2080);
nand U147 (N_147,In_3202,In_909);
or U148 (N_148,In_2414,In_3675);
nor U149 (N_149,In_4973,In_2445);
nand U150 (N_150,In_1607,In_2337);
and U151 (N_151,In_3866,In_2277);
nand U152 (N_152,In_4146,In_1236);
or U153 (N_153,In_1972,In_3286);
or U154 (N_154,In_3208,In_3366);
or U155 (N_155,In_3884,In_3163);
or U156 (N_156,In_4743,In_4069);
and U157 (N_157,In_3536,In_1132);
nor U158 (N_158,In_2358,In_4105);
or U159 (N_159,In_522,In_1473);
or U160 (N_160,In_4705,In_4165);
nand U161 (N_161,In_162,In_2522);
and U162 (N_162,In_3598,In_1302);
or U163 (N_163,In_128,In_3888);
and U164 (N_164,In_2319,In_3406);
or U165 (N_165,In_4230,In_2199);
xnor U166 (N_166,In_4135,In_4767);
or U167 (N_167,In_92,In_3412);
xor U168 (N_168,In_4529,In_4625);
nor U169 (N_169,In_2010,In_3280);
nand U170 (N_170,In_1977,In_440);
and U171 (N_171,In_3835,In_3956);
or U172 (N_172,In_2895,In_2533);
and U173 (N_173,In_3006,In_1697);
nand U174 (N_174,In_1168,In_4202);
or U175 (N_175,In_2146,In_2938);
or U176 (N_176,In_2173,In_3404);
or U177 (N_177,In_4046,In_2921);
nand U178 (N_178,In_2008,In_2382);
xnor U179 (N_179,In_2222,In_47);
or U180 (N_180,In_3423,In_2117);
and U181 (N_181,In_2150,In_4749);
nand U182 (N_182,In_3816,In_2350);
and U183 (N_183,In_4075,In_2554);
nand U184 (N_184,In_872,In_2916);
nor U185 (N_185,In_1187,In_2711);
and U186 (N_186,In_845,In_2722);
nor U187 (N_187,In_2790,In_2493);
or U188 (N_188,In_544,In_1206);
and U189 (N_189,In_2945,In_4970);
and U190 (N_190,In_2979,In_2518);
and U191 (N_191,In_3678,In_2181);
and U192 (N_192,In_4025,In_1345);
and U193 (N_193,In_2953,In_767);
or U194 (N_194,In_4873,In_2929);
xor U195 (N_195,In_3720,In_1528);
nor U196 (N_196,In_3698,In_3297);
nand U197 (N_197,In_1440,In_2018);
or U198 (N_198,In_4613,In_3776);
nand U199 (N_199,In_1402,In_2978);
xor U200 (N_200,In_2605,In_1090);
nor U201 (N_201,In_1902,In_315);
xor U202 (N_202,In_2079,In_638);
nand U203 (N_203,In_2413,In_2516);
nand U204 (N_204,In_189,In_2810);
or U205 (N_205,In_3370,In_2770);
nor U206 (N_206,In_225,In_4375);
or U207 (N_207,In_657,In_57);
xnor U208 (N_208,In_990,In_4328);
nand U209 (N_209,In_3934,In_957);
and U210 (N_210,In_2312,In_1635);
xor U211 (N_211,In_2282,In_2400);
and U212 (N_212,In_1356,In_2752);
and U213 (N_213,In_2389,In_622);
nor U214 (N_214,In_967,In_550);
xor U215 (N_215,In_3995,In_4459);
xor U216 (N_216,In_1734,In_1321);
nor U217 (N_217,In_3872,In_2940);
nor U218 (N_218,In_1491,In_147);
and U219 (N_219,In_724,In_2595);
xor U220 (N_220,In_3173,In_2510);
nor U221 (N_221,In_4289,In_2298);
nand U222 (N_222,In_2775,In_3547);
or U223 (N_223,In_765,In_3770);
nand U224 (N_224,In_2356,In_2796);
and U225 (N_225,In_1143,In_2498);
nand U226 (N_226,In_730,In_2492);
xor U227 (N_227,In_483,In_4403);
xnor U228 (N_228,In_1032,In_176);
nand U229 (N_229,In_1191,In_1019);
or U230 (N_230,In_2771,In_4361);
nand U231 (N_231,In_3837,In_2276);
nand U232 (N_232,In_1127,In_4593);
or U233 (N_233,In_3210,In_4528);
or U234 (N_234,In_2704,In_3350);
nor U235 (N_235,In_4762,In_2575);
or U236 (N_236,In_2963,In_2288);
nor U237 (N_237,In_1496,In_4866);
nand U238 (N_238,In_2724,In_1261);
nand U239 (N_239,In_3156,In_2890);
nor U240 (N_240,In_171,In_2061);
nor U241 (N_241,In_4223,In_4635);
or U242 (N_242,In_2609,In_4679);
nor U243 (N_243,In_2555,In_4828);
and U244 (N_244,In_1660,In_4807);
or U245 (N_245,In_3601,In_2561);
nor U246 (N_246,In_1504,In_1145);
nor U247 (N_247,In_4311,In_2618);
nand U248 (N_248,In_2827,In_3394);
or U249 (N_249,In_1351,In_4588);
or U250 (N_250,In_1712,In_2219);
xor U251 (N_251,In_969,In_4590);
nand U252 (N_252,In_4943,In_514);
nor U253 (N_253,In_1725,In_3744);
nand U254 (N_254,In_1919,In_1078);
nand U255 (N_255,In_3993,In_299);
or U256 (N_256,In_87,In_631);
nand U257 (N_257,In_1868,In_1719);
or U258 (N_258,In_4662,In_994);
and U259 (N_259,In_2788,In_1215);
nor U260 (N_260,In_3032,In_3603);
xnor U261 (N_261,In_904,In_2275);
or U262 (N_262,In_1531,In_4392);
nor U263 (N_263,In_2333,In_1344);
or U264 (N_264,In_3588,In_4843);
or U265 (N_265,In_413,In_3545);
nor U266 (N_266,In_4902,In_2155);
nor U267 (N_267,In_4888,In_3937);
nand U268 (N_268,In_1300,In_2647);
nor U269 (N_269,In_1565,In_978);
or U270 (N_270,In_1114,In_682);
nand U271 (N_271,In_3308,In_1384);
xnor U272 (N_272,In_2501,In_2207);
and U273 (N_273,In_1322,In_3221);
or U274 (N_274,In_1762,In_4342);
nor U275 (N_275,In_3962,In_883);
nand U276 (N_276,In_3143,In_3907);
or U277 (N_277,In_2314,In_635);
and U278 (N_278,In_2435,In_4515);
nand U279 (N_279,In_3779,In_2233);
and U280 (N_280,In_3455,In_4085);
nand U281 (N_281,In_4002,In_19);
or U282 (N_282,In_641,In_3044);
xor U283 (N_283,In_2983,In_3465);
nand U284 (N_284,In_2361,In_1869);
nor U285 (N_285,In_4855,In_3538);
or U286 (N_286,In_1887,In_1263);
nor U287 (N_287,In_4072,In_64);
and U288 (N_288,In_1548,In_222);
or U289 (N_289,In_4422,In_4868);
nand U290 (N_290,In_3078,In_3467);
nor U291 (N_291,In_4788,In_495);
nor U292 (N_292,In_984,In_3805);
xnor U293 (N_293,In_1324,In_1039);
and U294 (N_294,In_1536,In_1113);
or U295 (N_295,In_2523,In_2834);
and U296 (N_296,In_1513,In_554);
nor U297 (N_297,In_795,In_2572);
nand U298 (N_298,In_742,In_324);
and U299 (N_299,In_1974,In_3857);
nor U300 (N_300,In_4215,In_3940);
and U301 (N_301,In_4981,In_2147);
or U302 (N_302,In_661,In_1674);
nor U303 (N_303,In_3608,In_422);
xor U304 (N_304,In_4811,In_1364);
nor U305 (N_305,In_3175,In_3062);
nand U306 (N_306,In_3424,In_4466);
nand U307 (N_307,In_88,In_1458);
nor U308 (N_308,In_3365,In_4277);
or U309 (N_309,In_3363,In_2142);
nor U310 (N_310,In_216,In_577);
and U311 (N_311,In_2705,In_4456);
xor U312 (N_312,In_2320,In_1770);
nor U313 (N_313,In_1014,In_4168);
or U314 (N_314,In_4489,In_2187);
or U315 (N_315,In_634,In_4308);
nand U316 (N_316,In_104,In_3929);
nor U317 (N_317,In_950,In_3094);
xnor U318 (N_318,In_2727,In_4953);
or U319 (N_319,In_3144,In_2268);
nand U320 (N_320,In_4919,In_4726);
nand U321 (N_321,In_4835,In_2213);
nor U322 (N_322,In_2825,In_3259);
and U323 (N_323,In_4119,In_3886);
and U324 (N_324,In_1484,In_4397);
and U325 (N_325,In_691,In_3085);
nand U326 (N_326,In_1208,In_3607);
nor U327 (N_327,In_3871,In_4024);
nand U328 (N_328,In_820,In_667);
nand U329 (N_329,In_530,In_915);
and U330 (N_330,In_2599,In_1485);
nand U331 (N_331,In_1570,In_3326);
nand U332 (N_332,In_2802,In_1121);
nor U333 (N_333,In_393,In_3933);
and U334 (N_334,In_2567,In_1420);
or U335 (N_335,In_4126,In_3413);
xor U336 (N_336,In_829,In_2322);
xor U337 (N_337,In_4997,In_3775);
xor U338 (N_338,In_1030,In_2371);
or U339 (N_339,In_3043,In_462);
and U340 (N_340,In_4581,In_858);
and U341 (N_341,In_1554,In_788);
or U342 (N_342,In_2616,In_3250);
xor U343 (N_343,In_2308,In_4794);
nand U344 (N_344,In_2095,In_2295);
or U345 (N_345,In_3965,In_4541);
nor U346 (N_346,In_625,In_3942);
nand U347 (N_347,In_1235,In_383);
xor U348 (N_348,In_2715,In_1042);
or U349 (N_349,In_4717,In_3733);
xor U350 (N_350,In_598,In_2004);
xnor U351 (N_351,In_3705,In_728);
and U352 (N_352,In_11,In_4382);
and U353 (N_353,In_3100,In_2658);
nand U354 (N_354,In_938,In_824);
nand U355 (N_355,In_3804,In_3642);
xor U356 (N_356,In_4416,In_878);
nand U357 (N_357,In_1879,In_2044);
nand U358 (N_358,In_2980,In_1821);
nor U359 (N_359,In_443,In_652);
xor U360 (N_360,In_1476,In_2619);
or U361 (N_361,In_51,In_1782);
nor U362 (N_362,In_3471,In_3931);
or U363 (N_363,In_4132,In_3803);
nand U364 (N_364,In_4144,In_320);
nor U365 (N_365,In_3112,In_4381);
and U366 (N_366,In_3332,In_2657);
xor U367 (N_367,In_10,In_4127);
nand U368 (N_368,In_1157,In_246);
xor U369 (N_369,In_1228,In_3811);
xor U370 (N_370,In_1709,In_4735);
nor U371 (N_371,In_3236,In_2910);
nand U372 (N_372,In_3722,In_79);
and U373 (N_373,In_4450,In_66);
or U374 (N_374,In_4272,In_744);
nand U375 (N_375,In_2093,In_1317);
or U376 (N_376,In_3101,In_2193);
nand U377 (N_377,In_4491,In_2165);
or U378 (N_378,In_2966,In_1571);
nand U379 (N_379,In_18,In_378);
or U380 (N_380,In_4419,In_4758);
nor U381 (N_381,In_2458,In_561);
xnor U382 (N_382,In_2529,In_71);
or U383 (N_383,In_90,In_3595);
or U384 (N_384,In_4090,In_2376);
xnor U385 (N_385,In_337,In_4900);
nor U386 (N_386,In_1918,In_4673);
and U387 (N_387,In_289,In_3540);
and U388 (N_388,In_4432,In_2970);
nand U389 (N_389,In_3205,In_3499);
nand U390 (N_390,In_1488,In_4411);
xnor U391 (N_391,In_2374,In_3273);
and U392 (N_392,In_2459,In_4242);
xor U393 (N_393,In_4337,In_3555);
or U394 (N_394,In_59,In_2072);
nand U395 (N_395,In_1299,In_2210);
nor U396 (N_396,In_3461,In_3957);
and U397 (N_397,In_3095,In_4000);
or U398 (N_398,In_4141,In_2743);
and U399 (N_399,In_2216,In_1122);
xor U400 (N_400,In_2992,In_4268);
xnor U401 (N_401,In_2316,In_941);
nand U402 (N_402,In_3008,In_1796);
and U403 (N_403,In_1411,In_3108);
nand U404 (N_404,In_4737,In_1971);
nand U405 (N_405,In_1027,In_1308);
nand U406 (N_406,In_2132,In_2380);
nand U407 (N_407,In_3828,In_2474);
nor U408 (N_408,In_1893,In_807);
nand U409 (N_409,In_935,In_2917);
xnor U410 (N_410,In_1412,In_1243);
or U411 (N_411,In_2935,In_656);
xor U412 (N_412,In_1054,In_3503);
xnor U413 (N_413,In_4632,In_4210);
nand U414 (N_414,In_2329,In_615);
xor U415 (N_415,In_3662,In_1556);
nor U416 (N_416,In_1282,In_911);
and U417 (N_417,In_4314,In_4643);
nor U418 (N_418,In_1779,In_168);
or U419 (N_419,In_1550,In_4384);
nor U420 (N_420,In_2343,In_112);
xor U421 (N_421,In_567,In_2073);
nand U422 (N_422,In_774,In_860);
or U423 (N_423,In_1067,In_170);
xnor U424 (N_424,In_1991,In_2696);
xor U425 (N_425,In_520,In_3105);
and U426 (N_426,In_1045,In_1043);
nor U427 (N_427,In_3198,In_3091);
xnor U428 (N_428,In_3025,In_3748);
or U429 (N_429,In_2139,In_1567);
or U430 (N_430,In_4142,In_551);
or U431 (N_431,In_4891,In_1810);
or U432 (N_432,In_3481,In_201);
nor U433 (N_433,In_690,In_4226);
xor U434 (N_434,In_431,In_1241);
or U435 (N_435,In_3768,In_3000);
and U436 (N_436,In_7,In_906);
nand U437 (N_437,In_565,In_1589);
nor U438 (N_438,In_893,In_4899);
and U439 (N_439,In_2390,In_2123);
or U440 (N_440,In_2596,In_449);
xnor U441 (N_441,In_166,In_2497);
xor U442 (N_442,In_470,In_3244);
and U443 (N_443,In_809,In_4336);
or U444 (N_444,In_3260,In_578);
nand U445 (N_445,In_4294,In_3206);
and U446 (N_446,In_3473,In_696);
or U447 (N_447,In_1818,In_2606);
nand U448 (N_448,In_1058,In_653);
or U449 (N_449,In_1756,In_1149);
xor U450 (N_450,In_3498,In_372);
nor U451 (N_451,In_2296,In_752);
and U452 (N_452,In_1759,In_2368);
nand U453 (N_453,In_3558,In_1847);
and U454 (N_454,In_3253,In_3204);
xnor U455 (N_455,In_3246,In_93);
nand U456 (N_456,In_1451,In_2663);
or U457 (N_457,In_404,In_1735);
nor U458 (N_458,In_1335,In_1854);
and U459 (N_459,In_995,In_3841);
nand U460 (N_460,In_4494,In_2815);
nor U461 (N_461,In_2748,In_1943);
xnor U462 (N_462,In_2250,In_2901);
and U463 (N_463,In_3336,In_44);
or U464 (N_464,In_1376,In_349);
xor U465 (N_465,In_2776,In_4374);
nand U466 (N_466,In_4054,In_3216);
nor U467 (N_467,In_2418,In_1419);
and U468 (N_468,In_1886,In_2807);
and U469 (N_469,In_297,In_1105);
or U470 (N_470,In_506,In_2564);
and U471 (N_471,In_254,In_343);
and U472 (N_472,In_1945,In_3054);
nor U473 (N_473,In_1276,In_4218);
xor U474 (N_474,In_1245,In_2393);
or U475 (N_475,In_1863,In_2158);
xor U476 (N_476,In_3930,In_966);
xnor U477 (N_477,In_1454,In_412);
xor U478 (N_478,In_2830,In_1609);
and U479 (N_479,In_2559,In_1898);
xor U480 (N_480,In_2597,In_1551);
and U481 (N_481,In_1792,In_1125);
xnor U482 (N_482,In_2311,In_3170);
or U483 (N_483,In_1997,In_4131);
and U484 (N_484,In_3311,In_3958);
or U485 (N_485,In_1009,In_3089);
and U486 (N_486,In_3002,In_2812);
nor U487 (N_487,In_2957,In_3673);
nand U488 (N_488,In_3602,In_1588);
nor U489 (N_489,In_2346,In_2131);
or U490 (N_490,In_517,In_3702);
or U491 (N_491,In_4417,In_1994);
and U492 (N_492,In_664,In_836);
nor U493 (N_493,In_2948,In_2101);
xor U494 (N_494,In_4660,In_727);
and U495 (N_495,In_4182,In_719);
and U496 (N_496,In_4229,In_1174);
and U497 (N_497,In_421,In_4516);
nor U498 (N_498,In_1337,In_3296);
or U499 (N_499,In_3009,In_725);
nor U500 (N_500,In_2891,In_2821);
nand U501 (N_501,In_2170,In_4400);
or U502 (N_502,In_15,In_758);
and U503 (N_503,In_1380,In_472);
or U504 (N_504,In_3624,In_367);
or U505 (N_505,In_4116,In_49);
nand U506 (N_506,In_916,In_1309);
xnor U507 (N_507,In_1633,In_4848);
nor U508 (N_508,In_1223,In_871);
xnor U509 (N_509,In_2396,In_3343);
nand U510 (N_510,In_2803,In_2383);
nand U511 (N_511,In_3790,In_1123);
nor U512 (N_512,In_308,In_2009);
and U513 (N_513,In_4537,In_1502);
nand U514 (N_514,In_2167,In_4221);
xor U515 (N_515,In_126,In_501);
nor U516 (N_516,In_4238,In_4978);
nand U517 (N_517,In_3400,In_569);
nor U518 (N_518,In_2204,In_1256);
nor U519 (N_519,In_141,In_686);
and U520 (N_520,In_921,In_1639);
nand U521 (N_521,In_4867,In_3058);
nand U522 (N_522,In_4571,In_2053);
and U523 (N_523,In_3014,In_3159);
and U524 (N_524,In_3685,In_3139);
xnor U525 (N_525,In_38,In_414);
xnor U526 (N_526,In_2036,In_1224);
nor U527 (N_527,In_3927,In_3252);
nor U528 (N_528,In_840,In_1825);
xor U529 (N_529,In_4080,In_3567);
nand U530 (N_530,In_4530,In_3533);
and U531 (N_531,In_4157,In_1229);
xor U532 (N_532,In_666,In_2043);
and U533 (N_533,In_2750,In_558);
nand U534 (N_534,In_539,In_2366);
and U535 (N_535,In_3721,In_3701);
and U536 (N_536,In_3368,In_2873);
nand U537 (N_537,In_3231,In_1025);
xnor U538 (N_538,In_406,In_3403);
nand U539 (N_539,In_4629,In_4313);
and U540 (N_540,In_338,In_548);
and U541 (N_541,In_1099,In_4578);
nand U542 (N_542,In_2310,In_304);
nand U543 (N_543,In_3469,In_1480);
xnor U544 (N_544,In_3687,In_2591);
and U545 (N_545,In_1395,In_4567);
xor U546 (N_546,In_4681,In_2969);
and U547 (N_547,In_3566,In_3682);
and U548 (N_548,In_3042,In_13);
xnor U549 (N_549,In_3388,In_4709);
and U550 (N_550,In_2426,In_3556);
or U551 (N_551,In_4909,In_4739);
and U552 (N_552,In_203,In_2266);
and U553 (N_553,In_543,In_1723);
nor U554 (N_554,In_869,In_4600);
nor U555 (N_555,In_513,In_1799);
and U556 (N_556,In_1409,In_4554);
xnor U557 (N_557,In_1170,In_2436);
or U558 (N_558,In_4558,In_2859);
xor U559 (N_559,In_741,In_2652);
and U560 (N_560,In_1631,In_499);
xnor U561 (N_561,In_2660,In_679);
nor U562 (N_562,In_4693,In_2741);
and U563 (N_563,In_4113,In_1304);
xnor U564 (N_564,In_286,In_4996);
nand U565 (N_565,In_4993,In_2634);
and U566 (N_566,In_1173,In_2415);
xor U567 (N_567,In_4394,In_269);
nand U568 (N_568,In_4833,In_1013);
nor U569 (N_569,In_4499,In_1271);
nand U570 (N_570,In_2995,In_4817);
xor U571 (N_571,In_2931,In_3582);
nand U572 (N_572,In_4619,In_2904);
or U573 (N_573,In_2850,In_3860);
and U574 (N_574,In_1883,In_1155);
and U575 (N_575,In_4803,In_4481);
xnor U576 (N_576,In_1479,In_1211);
nand U577 (N_577,In_2422,In_503);
nor U578 (N_578,In_4064,In_3925);
nor U579 (N_579,In_4701,In_3491);
nor U580 (N_580,In_1772,In_4160);
or U581 (N_581,In_1558,In_4842);
nor U582 (N_582,In_3446,In_4976);
xor U583 (N_583,In_476,In_4153);
nand U584 (N_584,In_3711,In_4465);
and U585 (N_585,In_2238,In_4405);
xnor U586 (N_586,In_3686,In_2189);
or U587 (N_587,In_2381,In_3815);
xor U588 (N_588,In_1970,In_4949);
nand U589 (N_589,In_3462,In_2789);
nor U590 (N_590,In_3793,In_3486);
or U591 (N_591,In_1284,In_1838);
nand U592 (N_592,In_4972,In_4551);
and U593 (N_593,In_2037,In_688);
xnor U594 (N_594,In_145,In_2176);
nor U595 (N_595,In_3136,In_4665);
xnor U596 (N_596,In_4748,In_3738);
and U597 (N_597,In_2801,In_4688);
nand U598 (N_598,In_3643,In_3649);
nand U599 (N_599,In_619,In_2479);
or U600 (N_600,In_3402,In_3851);
nand U601 (N_601,In_843,In_2515);
xnor U602 (N_602,In_3987,In_3905);
nand U603 (N_603,In_2840,In_1092);
and U604 (N_604,In_330,In_2300);
xor U605 (N_605,In_4082,In_648);
xnor U606 (N_606,In_2221,In_2172);
nand U607 (N_607,In_3596,In_2997);
nor U608 (N_608,In_1162,In_1248);
and U609 (N_609,In_480,In_1298);
nand U610 (N_610,In_39,In_2033);
and U611 (N_611,In_3021,In_3813);
nor U612 (N_612,In_4143,In_3519);
nor U613 (N_613,In_3693,In_4777);
nor U614 (N_614,In_2118,In_4933);
or U615 (N_615,In_778,In_2714);
or U616 (N_616,In_2885,In_37);
or U617 (N_617,In_2098,In_1824);
nor U618 (N_618,In_2560,In_4032);
xor U619 (N_619,In_4407,In_3454);
xnor U620 (N_620,In_2212,In_2197);
nor U621 (N_621,In_4335,In_368);
and U622 (N_622,In_601,In_1082);
nor U623 (N_623,In_4093,In_706);
xor U624 (N_624,In_2999,In_2215);
xnor U625 (N_625,In_2911,In_3484);
nand U626 (N_626,In_4776,In_209);
or U627 (N_627,In_4614,In_1091);
xor U628 (N_628,In_178,In_3110);
and U629 (N_629,In_1437,In_2739);
nand U630 (N_630,In_70,In_1722);
or U631 (N_631,In_1369,In_999);
or U632 (N_632,In_1445,In_1167);
nor U633 (N_633,In_3456,In_2512);
nand U634 (N_634,In_3119,In_2829);
xnor U635 (N_635,In_2237,In_779);
nor U636 (N_636,In_2767,In_4871);
or U637 (N_637,In_4323,In_2325);
nand U638 (N_638,In_4785,In_4444);
nand U639 (N_639,In_2055,In_2016);
or U640 (N_640,In_1773,In_3560);
xor U641 (N_641,In_2541,In_265);
xnor U642 (N_642,In_1761,In_4326);
or U643 (N_643,In_1222,In_4677);
xnor U644 (N_644,In_294,In_1783);
or U645 (N_645,In_1233,In_791);
and U646 (N_646,In_4921,In_3653);
nand U647 (N_647,In_4059,In_3304);
or U648 (N_648,In_4241,In_3448);
nor U649 (N_649,In_1336,In_3534);
nor U650 (N_650,In_3709,In_279);
xor U651 (N_651,In_4468,In_2011);
nand U652 (N_652,In_2482,In_4115);
xnor U653 (N_653,In_1897,In_1267);
xnor U654 (N_654,In_2535,In_429);
nor U655 (N_655,In_2905,In_4357);
and U656 (N_656,In_2692,In_900);
or U657 (N_657,In_3829,In_4252);
and U658 (N_658,In_4631,In_2816);
nor U659 (N_659,In_2936,In_274);
nand U660 (N_660,In_2476,In_2081);
nor U661 (N_661,In_291,In_3647);
nand U662 (N_662,In_4573,In_4227);
and U663 (N_663,In_1737,In_1713);
nor U664 (N_664,In_4373,In_1024);
nor U665 (N_665,In_2377,In_4942);
or U666 (N_666,In_2468,In_3735);
or U667 (N_667,In_2590,In_2256);
and U668 (N_668,In_1178,In_4977);
xor U669 (N_669,In_3810,In_157);
nor U670 (N_670,In_91,In_4246);
nor U671 (N_671,In_1985,In_1394);
and U672 (N_672,In_4556,In_4441);
and U673 (N_673,In_2481,In_3102);
or U674 (N_674,In_3040,In_3919);
or U675 (N_675,In_4293,In_4708);
and U676 (N_676,In_636,In_266);
xnor U677 (N_677,In_859,In_4617);
or U678 (N_678,In_427,In_2503);
or U679 (N_679,In_1416,In_3493);
and U680 (N_680,In_4544,In_97);
nor U681 (N_681,In_2861,In_1396);
or U682 (N_682,In_1069,In_710);
nand U683 (N_683,In_1920,In_3063);
nand U684 (N_684,In_1512,In_1230);
or U685 (N_685,In_314,In_1747);
nand U686 (N_686,In_4372,In_3096);
and U687 (N_687,In_288,In_4107);
nor U688 (N_688,In_3266,In_207);
nand U689 (N_689,In_4952,In_734);
or U690 (N_690,In_3131,In_1610);
xnor U691 (N_691,In_3039,In_2710);
nand U692 (N_692,In_4301,In_2291);
nor U693 (N_693,In_602,In_4527);
nand U694 (N_694,In_1749,In_2780);
nor U695 (N_695,In_2545,In_1695);
and U696 (N_696,In_2340,In_4079);
nand U697 (N_697,In_4802,In_2677);
nand U698 (N_698,In_4173,In_4765);
and U699 (N_699,In_4858,In_4546);
and U700 (N_700,In_1816,In_4534);
and U701 (N_701,In_2607,In_1475);
or U702 (N_702,In_1259,In_4930);
and U703 (N_703,In_4825,In_3497);
xor U704 (N_704,In_1986,In_521);
nand U705 (N_705,In_3500,In_85);
nor U706 (N_706,In_1642,In_1238);
and U707 (N_707,In_3909,In_2943);
and U708 (N_708,In_381,In_4756);
and U709 (N_709,In_1590,In_276);
and U710 (N_710,In_2480,In_1001);
and U711 (N_711,In_1146,In_3072);
or U712 (N_712,In_1,In_4247);
nor U713 (N_713,In_130,In_3145);
and U714 (N_714,In_317,In_4473);
and U715 (N_715,In_1990,In_1679);
nor U716 (N_716,In_1842,In_321);
and U717 (N_717,In_4609,In_1441);
nor U718 (N_718,In_3671,In_1339);
nor U719 (N_719,In_3782,In_1963);
nor U720 (N_720,In_1784,In_3033);
nand U721 (N_721,In_4706,In_1514);
nor U722 (N_722,In_1117,In_2460);
and U723 (N_723,In_3146,In_1096);
nand U724 (N_724,In_3045,In_4601);
nand U725 (N_725,In_574,In_67);
xor U726 (N_726,In_3478,In_3409);
nand U727 (N_727,In_100,In_1508);
nor U728 (N_728,In_2019,In_3548);
nor U729 (N_729,In_4533,In_376);
nor U730 (N_730,In_4369,In_3858);
nand U731 (N_731,In_885,In_1923);
nor U732 (N_732,In_1051,In_468);
nand U733 (N_733,In_2923,In_1802);
xnor U734 (N_734,In_3853,In_2781);
and U735 (N_735,In_3185,In_4029);
nand U736 (N_736,In_4410,In_3579);
nand U737 (N_737,In_3617,In_2457);
xor U738 (N_738,In_3463,In_2379);
xnor U739 (N_739,In_3809,In_1330);
or U740 (N_740,In_4994,In_989);
xnor U741 (N_741,In_4324,In_3627);
xnor U742 (N_742,In_4509,In_782);
xor U743 (N_743,In_3416,In_1975);
or U744 (N_744,In_4661,In_1745);
xnor U745 (N_745,In_3020,In_2122);
nand U746 (N_746,In_4652,In_4797);
xor U747 (N_747,In_2483,In_2754);
nor U748 (N_748,In_2336,In_1801);
nand U749 (N_749,In_2286,In_4746);
or U750 (N_750,In_753,In_3996);
nor U751 (N_751,In_3968,In_3861);
nand U752 (N_752,In_121,In_4827);
nand U753 (N_753,In_1771,In_4645);
xor U754 (N_754,In_3196,In_1845);
or U755 (N_755,In_1296,In_1636);
or U756 (N_756,In_3183,In_939);
nand U757 (N_757,In_738,In_3610);
and U758 (N_758,In_3511,In_4089);
nor U759 (N_759,In_1549,In_4406);
xnor U760 (N_760,In_3706,In_2675);
xor U761 (N_761,In_2543,In_952);
and U762 (N_762,In_955,In_1643);
or U763 (N_763,In_1961,In_3867);
xor U764 (N_764,In_2562,In_3338);
or U765 (N_765,In_4086,In_4271);
nor U766 (N_766,In_300,In_3314);
or U767 (N_767,In_4334,In_2862);
nand U768 (N_768,In_72,In_4013);
nor U769 (N_769,In_1080,In_3615);
and U770 (N_770,In_120,In_3910);
or U771 (N_771,In_2421,In_2868);
xor U772 (N_772,In_3612,In_570);
nand U773 (N_773,In_267,In_1200);
nand U774 (N_774,In_3902,In_1179);
nor U775 (N_775,In_4057,In_2645);
or U776 (N_776,In_4251,In_3542);
and U777 (N_777,In_1428,In_1405);
or U778 (N_778,In_2598,In_4685);
nor U779 (N_779,In_2870,In_2097);
and U780 (N_780,In_3527,In_1843);
or U781 (N_781,In_2220,In_3305);
xnor U782 (N_782,In_4721,In_748);
xnor U783 (N_783,In_1273,In_4694);
and U784 (N_784,In_2417,In_2200);
xor U785 (N_785,In_2580,In_4634);
xor U786 (N_786,In_351,In_3035);
or U787 (N_787,In_4098,In_3224);
or U788 (N_788,In_4641,In_3408);
nor U789 (N_789,In_2066,In_2764);
and U790 (N_790,In_818,In_3019);
and U791 (N_791,In_3896,In_1780);
or U792 (N_792,In_2571,In_515);
and U793 (N_793,In_2610,In_510);
or U794 (N_794,In_188,In_1715);
xor U795 (N_795,In_1134,In_4389);
nand U796 (N_796,In_1050,In_3172);
nor U797 (N_797,In_1881,In_4460);
or U798 (N_798,In_3794,In_4595);
xnor U799 (N_799,In_1940,In_1915);
or U800 (N_800,In_4256,In_4110);
nand U801 (N_801,In_4875,In_184);
nor U802 (N_802,In_586,In_153);
or U803 (N_803,In_2190,In_4819);
xnor U804 (N_804,In_945,In_3723);
or U805 (N_805,In_2718,In_1666);
nand U806 (N_806,In_1814,In_3611);
nor U807 (N_807,In_3654,In_4910);
nand U808 (N_808,In_4365,In_4622);
or U809 (N_809,In_179,In_2683);
nor U810 (N_810,In_1853,In_4960);
or U811 (N_811,In_4678,In_4770);
nand U812 (N_812,In_2544,In_1752);
and U813 (N_813,In_4155,In_4354);
and U814 (N_814,In_2087,In_1373);
nand U815 (N_815,In_2225,In_2786);
or U816 (N_816,In_3115,In_1763);
or U817 (N_817,In_182,In_2032);
nand U818 (N_818,In_3681,In_4214);
and U819 (N_819,In_4780,In_2779);
or U820 (N_820,In_2363,In_3971);
or U821 (N_821,In_4061,In_4814);
and U822 (N_822,In_3707,In_1382);
nand U823 (N_823,In_2438,In_1340);
xor U824 (N_824,In_4549,In_4290);
or U825 (N_825,In_1139,In_1358);
nor U826 (N_826,In_715,In_4099);
nand U827 (N_827,In_5,In_854);
nor U828 (N_828,In_2686,In_3310);
and U829 (N_829,In_2989,In_303);
xnor U830 (N_830,In_1016,In_2894);
nand U831 (N_831,In_4992,In_1182);
nand U832 (N_832,In_2694,In_4442);
or U833 (N_833,In_146,In_1965);
nand U834 (N_834,In_2768,In_2138);
nor U835 (N_835,In_1234,In_1360);
xor U836 (N_836,In_1160,In_1574);
and U837 (N_837,In_2993,In_4922);
xnor U838 (N_838,In_2462,In_3277);
nand U839 (N_839,In_749,In_4918);
nand U840 (N_840,In_1768,In_1597);
nor U841 (N_841,In_3319,In_452);
and U842 (N_842,In_4284,In_3411);
nor U843 (N_843,In_3391,In_3005);
and U844 (N_844,In_2271,In_2867);
xor U845 (N_845,In_1217,In_4961);
or U846 (N_846,In_3051,In_3609);
nand U847 (N_847,In_2410,In_731);
or U848 (N_848,In_3882,In_3704);
and U849 (N_849,In_1670,In_787);
nor U850 (N_850,In_478,In_4663);
or U851 (N_851,In_1257,In_2070);
nor U852 (N_852,In_1120,In_21);
xnor U853 (N_853,In_3466,In_1199);
or U854 (N_854,In_777,In_3807);
nand U855 (N_855,In_481,In_2099);
nand U856 (N_856,In_2294,In_1820);
nand U857 (N_857,In_4431,In_132);
xor U858 (N_858,In_3730,In_3651);
and U859 (N_859,In_3516,In_743);
and U860 (N_860,In_4414,In_1622);
xnor U861 (N_861,In_2029,In_124);
nor U862 (N_862,In_2025,In_3715);
or U863 (N_863,In_3275,In_2355);
nor U864 (N_864,In_927,In_1710);
and U865 (N_865,In_2226,In_2148);
nand U866 (N_866,In_839,In_199);
xor U867 (N_867,In_451,In_3614);
or U868 (N_868,In_672,In_1493);
and U869 (N_869,In_1603,In_3580);
xnor U870 (N_870,In_4194,In_931);
or U871 (N_871,In_4589,In_2283);
nor U872 (N_872,In_1649,In_2279);
and U873 (N_873,In_2747,In_2267);
or U874 (N_874,In_970,In_35);
or U875 (N_875,In_2446,In_3798);
or U876 (N_876,In_3453,In_913);
xnor U877 (N_877,In_512,In_1141);
xor U878 (N_878,In_4740,In_1951);
and U879 (N_879,In_3831,In_2407);
nand U880 (N_880,In_1708,In_3575);
nand U881 (N_881,In_1732,In_2318);
nand U882 (N_882,In_2005,In_2046);
xnor U883 (N_883,In_3291,In_2939);
nor U884 (N_884,In_3031,In_1218);
and U885 (N_885,In_721,In_334);
and U886 (N_886,In_2513,In_2526);
or U887 (N_887,In_1934,In_2278);
or U888 (N_888,In_2478,In_3160);
nor U889 (N_889,In_1608,In_3123);
nand U890 (N_890,In_1519,In_3382);
or U891 (N_891,In_2627,In_2726);
or U892 (N_892,In_873,In_2313);
nand U893 (N_893,In_2934,In_1391);
or U894 (N_894,In_3517,In_160);
and U895 (N_895,In_1673,In_4925);
nor U896 (N_896,In_4449,In_2394);
nor U897 (N_897,In_2514,In_2331);
nor U898 (N_898,In_3849,In_814);
nor U899 (N_899,In_2691,In_2494);
nand U900 (N_900,In_3667,In_3522);
nand U901 (N_901,In_1652,In_3442);
and U902 (N_902,In_4426,In_2206);
or U903 (N_903,In_4053,In_3531);
and U904 (N_904,In_1355,In_3832);
nand U905 (N_905,In_4923,In_3915);
nor U906 (N_906,In_3347,In_1501);
nand U907 (N_907,In_793,In_1540);
nor U908 (N_908,In_1138,In_500);
nand U909 (N_909,In_2587,In_3577);
and U910 (N_910,In_4163,In_1944);
or U911 (N_911,In_1442,In_53);
or U912 (N_912,In_3141,In_4094);
or U913 (N_913,In_4832,In_232);
nand U914 (N_914,In_702,In_2289);
xor U915 (N_915,In_4637,In_3868);
nor U916 (N_916,In_3240,In_3830);
xor U917 (N_917,In_4225,In_1283);
nor U918 (N_918,In_1864,In_2027);
and U919 (N_919,In_1855,In_675);
nor U920 (N_920,In_487,In_4404);
xnor U921 (N_921,In_3070,In_438);
or U922 (N_922,In_1406,In_4786);
and U923 (N_923,In_1896,In_4169);
nor U924 (N_924,In_256,In_2496);
xor U925 (N_925,In_3792,In_4211);
nor U926 (N_926,In_2878,In_3476);
xnor U927 (N_927,In_1487,In_4511);
or U928 (N_928,In_240,In_2499);
nor U929 (N_929,In_2171,In_341);
xnor U930 (N_930,In_1386,In_2461);
or U931 (N_931,In_4052,In_3574);
xnor U932 (N_932,In_1757,In_4380);
xnor U933 (N_933,In_1279,In_1102);
nor U934 (N_934,In_3578,In_4287);
nand U935 (N_935,In_3482,In_1086);
xnor U936 (N_936,In_1056,In_370);
and U937 (N_937,In_477,In_2849);
nor U938 (N_938,In_2409,In_2205);
nor U939 (N_939,In_4682,In_4111);
or U940 (N_940,In_3742,In_4623);
or U941 (N_941,In_1275,In_804);
and U942 (N_942,In_1293,In_2813);
xor U943 (N_943,In_318,In_3334);
or U944 (N_944,In_3836,In_3759);
nand U945 (N_945,In_992,In_200);
and U946 (N_946,In_2129,In_2617);
or U947 (N_947,In_889,In_1978);
or U948 (N_948,In_502,In_154);
nand U949 (N_949,In_3228,In_287);
xor U950 (N_950,In_1623,In_3512);
and U951 (N_951,In_4669,In_4676);
or U952 (N_952,In_1137,In_552);
nor U953 (N_953,In_4733,In_4288);
nor U954 (N_954,In_3766,In_3801);
nand U955 (N_955,In_3529,In_4798);
nand U956 (N_956,In_4498,In_3568);
nand U957 (N_957,In_4696,In_2104);
and U958 (N_958,In_1880,In_630);
nand U959 (N_959,In_2676,In_3360);
xor U960 (N_960,In_3895,In_2623);
and U961 (N_961,In_2604,In_825);
xor U962 (N_962,In_3232,In_4014);
xnor U963 (N_963,In_1453,In_4931);
xnor U964 (N_964,In_3834,In_764);
nor U965 (N_965,In_4890,In_2339);
xor U966 (N_966,In_1979,In_4911);
and U967 (N_967,In_4587,In_1465);
and U968 (N_968,In_2006,In_1865);
xnor U969 (N_969,In_4616,In_1265);
or U970 (N_970,In_3371,In_3695);
xnor U971 (N_971,In_592,In_1791);
and U972 (N_972,In_3953,In_4340);
xnor U973 (N_973,In_3606,In_1741);
or U974 (N_974,In_4683,In_4217);
nand U975 (N_975,In_3791,In_3506);
xor U976 (N_976,In_3920,In_1711);
nor U977 (N_977,In_3041,In_1546);
nand U978 (N_978,In_262,In_327);
nor U979 (N_979,In_4483,In_2845);
xnor U980 (N_980,In_2416,In_4804);
and U981 (N_981,In_36,In_3261);
nand U982 (N_982,In_1250,In_76);
and U983 (N_983,In_4121,In_3697);
xnor U984 (N_984,In_52,In_4897);
xor U985 (N_985,In_1927,In_2738);
xor U986 (N_986,In_628,In_1718);
nor U987 (N_987,In_1242,In_4237);
nor U988 (N_988,In_1000,In_1987);
nand U989 (N_989,In_2783,In_1733);
nor U990 (N_990,In_3410,In_3716);
nand U991 (N_991,In_144,In_4071);
or U992 (N_992,In_1212,In_4480);
and U993 (N_993,In_1085,In_2373);
nor U994 (N_994,In_3327,In_2542);
xnor U995 (N_995,In_3943,In_82);
nor U996 (N_996,In_2196,In_792);
nand U997 (N_997,In_4007,In_2024);
nor U998 (N_998,In_3289,In_1341);
xnor U999 (N_999,In_1518,In_3383);
nor U1000 (N_1000,In_3751,In_4006);
or U1001 (N_1001,In_1486,In_4539);
nand U1002 (N_1002,In_1933,In_3312);
or U1003 (N_1003,In_3521,In_4592);
and U1004 (N_1004,In_4174,In_2933);
and U1005 (N_1005,In_2839,In_163);
or U1006 (N_1006,In_4968,In_4907);
and U1007 (N_1007,In_2404,In_2451);
xor U1008 (N_1008,In_396,In_790);
xor U1009 (N_1009,In_138,In_3018);
nor U1010 (N_1010,In_2869,In_1192);
xor U1011 (N_1011,In_4760,In_541);
and U1012 (N_1012,In_2341,In_4951);
or U1013 (N_1013,In_993,In_2814);
nor U1014 (N_1014,In_3287,In_3251);
nor U1015 (N_1015,In_4212,In_32);
nand U1016 (N_1016,In_1545,In_33);
and U1017 (N_1017,In_1872,In_4401);
or U1018 (N_1018,In_3359,In_2611);
and U1019 (N_1019,In_1700,In_234);
nand U1020 (N_1020,In_397,In_937);
xnor U1021 (N_1021,In_3784,In_3543);
nor U1022 (N_1022,In_2749,In_45);
xor U1023 (N_1023,In_83,In_531);
or U1024 (N_1024,In_2534,In_3908);
and U1025 (N_1025,In_3212,In_670);
xor U1026 (N_1026,In_3254,In_2357);
or U1027 (N_1027,In_894,In_3290);
xnor U1028 (N_1028,In_4698,In_3313);
nor U1029 (N_1029,In_420,In_2896);
xnor U1030 (N_1030,In_2682,In_1472);
nor U1031 (N_1031,In_1657,In_1354);
and U1032 (N_1032,In_559,In_3785);
xnor U1033 (N_1033,In_3783,In_248);
xor U1034 (N_1034,In_1716,In_335);
and U1035 (N_1035,In_1999,In_4496);
nor U1036 (N_1036,In_3852,In_4959);
xnor U1037 (N_1037,In_400,In_613);
xor U1038 (N_1038,In_2112,In_771);
nor U1039 (N_1039,In_356,In_357);
nand U1040 (N_1040,In_1201,In_794);
xor U1041 (N_1041,In_997,In_369);
or U1042 (N_1042,In_4586,In_576);
xnor U1043 (N_1043,In_3298,In_3992);
nor U1044 (N_1044,In_2287,In_3502);
nand U1045 (N_1045,In_3367,In_2464);
nand U1046 (N_1046,In_1721,In_4265);
and U1047 (N_1047,In_545,In_3149);
xor U1048 (N_1048,In_3960,In_4926);
xor U1049 (N_1049,In_2625,In_4233);
and U1050 (N_1050,In_704,In_4467);
nor U1051 (N_1051,In_2700,In_4532);
nor U1052 (N_1052,In_3496,In_169);
nor U1053 (N_1053,In_4413,In_1436);
nand U1054 (N_1054,In_1057,In_2762);
or U1055 (N_1055,In_1829,In_1269);
xor U1056 (N_1056,In_3181,In_2981);
nor U1057 (N_1057,In_3150,In_4240);
nand U1058 (N_1058,In_1836,In_3724);
nand U1059 (N_1059,In_2484,In_2475);
and U1060 (N_1060,In_3787,In_3827);
nor U1061 (N_1061,In_4934,In_926);
nor U1062 (N_1062,In_3561,In_2638);
xnor U1063 (N_1063,In_2946,In_3258);
nor U1064 (N_1064,In_27,In_332);
xor U1065 (N_1065,In_1144,In_642);
and U1066 (N_1066,In_4531,In_1407);
or U1067 (N_1067,In_3590,In_2893);
nor U1068 (N_1068,In_185,In_1569);
nand U1069 (N_1069,In_2487,In_4646);
nor U1070 (N_1070,In_1161,In_4012);
or U1071 (N_1071,In_4250,In_1065);
and U1072 (N_1072,In_3401,In_621);
nor U1073 (N_1073,In_4497,In_4295);
nor U1074 (N_1074,In_2092,In_2622);
nor U1075 (N_1075,In_1500,In_651);
or U1076 (N_1076,In_1841,In_1370);
xor U1077 (N_1077,In_1537,In_1225);
or U1078 (N_1078,In_1696,In_3757);
and U1079 (N_1079,In_4206,In_3758);
or U1080 (N_1080,In_880,In_1834);
and U1081 (N_1081,In_226,In_96);
xnor U1082 (N_1082,In_1535,In_4766);
nor U1083 (N_1083,In_1462,In_251);
nand U1084 (N_1084,In_1562,In_290);
and U1085 (N_1085,In_2359,In_3998);
and U1086 (N_1086,In_4861,In_1835);
nand U1087 (N_1087,In_1828,In_1414);
nor U1088 (N_1088,In_4278,In_3954);
nor U1089 (N_1089,In_4575,In_4520);
nand U1090 (N_1090,In_2547,In_3988);
nor U1091 (N_1091,In_3745,In_473);
nor U1092 (N_1092,In_2509,In_2231);
xor U1093 (N_1093,In_1899,In_2408);
and U1094 (N_1094,In_2259,In_3991);
nor U1095 (N_1095,In_3591,In_3300);
and U1096 (N_1096,In_3679,In_4626);
nor U1097 (N_1097,In_3248,In_4428);
nand U1098 (N_1098,In_4624,In_4935);
or U1099 (N_1099,In_81,In_3840);
xor U1100 (N_1100,In_1917,In_1538);
nand U1101 (N_1101,In_4878,In_2315);
xnor U1102 (N_1102,In_193,In_213);
and U1103 (N_1103,In_1667,In_3357);
and U1104 (N_1104,In_976,In_4860);
nand U1105 (N_1105,In_344,In_2);
and U1106 (N_1106,In_3303,In_3324);
or U1107 (N_1107,In_2636,In_1363);
nand U1108 (N_1108,In_560,In_3983);
nor U1109 (N_1109,In_585,In_1654);
and U1110 (N_1110,In_2453,In_2988);
or U1111 (N_1111,In_3345,In_1460);
xnor U1112 (N_1112,In_1130,In_821);
nand U1113 (N_1113,In_1439,In_4461);
nor U1114 (N_1114,In_2257,In_4815);
nor U1115 (N_1115,In_3637,In_2052);
nand U1116 (N_1116,In_4612,In_964);
nor U1117 (N_1117,In_1031,In_3245);
or U1118 (N_1118,In_3507,In_612);
nand U1119 (N_1119,In_4189,In_700);
nor U1120 (N_1120,In_507,In_4010);
xor U1121 (N_1121,In_2120,In_584);
or U1122 (N_1122,In_1931,In_4570);
nor U1123 (N_1123,In_2662,In_516);
or U1124 (N_1124,In_1305,In_4905);
xor U1125 (N_1125,In_2841,In_25);
nand U1126 (N_1126,In_3989,In_4350);
or U1127 (N_1127,In_415,In_2068);
xor U1128 (N_1128,In_1352,In_3026);
nor U1129 (N_1129,In_350,In_708);
nor U1130 (N_1130,In_221,In_4699);
nand U1131 (N_1131,In_2285,In_605);
nand U1132 (N_1132,In_4839,In_2795);
xor U1133 (N_1133,In_775,In_2105);
or U1134 (N_1134,In_4862,In_3749);
or U1135 (N_1135,In_1948,In_4668);
and U1136 (N_1136,In_17,In_99);
or U1137 (N_1137,In_2877,In_895);
nand U1138 (N_1138,In_133,In_4083);
or U1139 (N_1139,In_1851,In_4171);
nor U1140 (N_1140,In_4964,In_3523);
or U1141 (N_1141,In_1837,In_3445);
nand U1142 (N_1142,In_4870,In_2309);
or U1143 (N_1143,In_3235,In_1680);
xor U1144 (N_1144,In_348,In_1587);
and U1145 (N_1145,In_1100,In_4670);
xor U1146 (N_1146,In_3762,In_2127);
and U1147 (N_1147,In_3855,In_471);
nand U1148 (N_1148,In_4114,In_1862);
and U1149 (N_1149,In_2403,In_2128);
or U1150 (N_1150,In_887,In_799);
nor U1151 (N_1151,In_624,In_4062);
nor U1152 (N_1152,In_3138,In_4611);
and U1153 (N_1153,In_3691,In_4259);
or U1154 (N_1154,In_2442,In_3222);
nor U1155 (N_1155,In_4454,In_4656);
xnor U1156 (N_1156,In_4779,In_4199);
nand U1157 (N_1157,In_447,In_3772);
and U1158 (N_1158,In_2402,In_3262);
nand U1159 (N_1159,In_4504,In_3814);
and U1160 (N_1160,In_881,In_1968);
nor U1161 (N_1161,In_3856,In_4164);
and U1162 (N_1162,In_2094,In_1526);
nor U1163 (N_1163,In_991,In_1738);
xor U1164 (N_1164,In_1023,In_159);
and U1165 (N_1165,In_4810,In_2136);
xor U1166 (N_1166,In_2108,In_1937);
or U1167 (N_1167,In_4249,In_2621);
or U1168 (N_1168,In_194,In_1988);
nor U1169 (N_1169,In_1611,In_1313);
and U1170 (N_1170,In_358,In_4027);
nand U1171 (N_1171,In_4583,In_2265);
xnor U1172 (N_1172,In_4346,In_3535);
and U1173 (N_1173,In_4003,In_2723);
nand U1174 (N_1174,In_3796,In_4120);
nor U1175 (N_1175,In_826,In_272);
nand U1176 (N_1176,In_3587,In_416);
xnor U1177 (N_1177,In_3583,In_277);
nor U1178 (N_1178,In_1483,In_1823);
xnor U1179 (N_1179,In_1286,In_2485);
or U1180 (N_1180,In_1289,In_4319);
xor U1181 (N_1181,In_4808,In_1641);
xnor U1182 (N_1182,In_1758,In_1118);
xor U1183 (N_1183,In_4490,In_3713);
nand U1184 (N_1184,In_498,In_1578);
nor U1185 (N_1185,In_4906,In_2145);
and U1186 (N_1186,In_2915,In_4628);
xor U1187 (N_1187,In_432,In_705);
nor U1188 (N_1188,In_3229,In_2305);
nor U1189 (N_1189,In_801,In_3257);
or U1190 (N_1190,In_1342,In_1185);
xor U1191 (N_1191,In_2067,In_2002);
and U1192 (N_1192,In_4,In_4547);
nand U1193 (N_1193,In_4145,In_4134);
or U1194 (N_1194,In_494,In_3419);
and U1195 (N_1195,In_4667,In_3530);
and U1196 (N_1196,In_1564,In_4781);
nor U1197 (N_1197,In_1103,In_4049);
xor U1198 (N_1198,In_3822,In_3355);
and U1199 (N_1199,In_3628,In_2378);
nor U1200 (N_1200,In_3823,In_3352);
xor U1201 (N_1201,In_1005,In_54);
nand U1202 (N_1202,In_2297,In_278);
and U1203 (N_1203,In_1954,In_4818);
and U1204 (N_1204,In_1980,In_2517);
xnor U1205 (N_1205,In_4385,In_3972);
or U1206 (N_1206,In_4347,In_2602);
xor U1207 (N_1207,In_2465,In_3819);
nor U1208 (N_1208,In_2540,In_3600);
xor U1209 (N_1209,In_4316,In_1297);
or U1210 (N_1210,In_1798,In_3421);
and U1211 (N_1211,In_2674,In_2569);
nand U1212 (N_1212,In_1101,In_282);
nand U1213 (N_1213,In_3226,In_977);
and U1214 (N_1214,In_1383,In_2239);
nor U1215 (N_1215,In_1214,In_1809);
and U1216 (N_1216,In_581,In_4269);
or U1217 (N_1217,In_4458,In_2847);
nand U1218 (N_1218,In_1953,In_1743);
nand U1219 (N_1219,In_3295,In_1181);
and U1220 (N_1220,In_1247,In_2433);
nor U1221 (N_1221,In_529,In_905);
nand U1222 (N_1222,In_643,In_2143);
and U1223 (N_1223,In_245,In_4603);
xnor U1224 (N_1224,In_3967,In_3923);
nand U1225 (N_1225,In_2639,In_1424);
nand U1226 (N_1226,In_2909,In_1253);
xor U1227 (N_1227,In_1690,In_3887);
nand U1228 (N_1228,In_4150,In_4262);
xor U1229 (N_1229,In_2881,In_2628);
nand U1230 (N_1230,In_4654,In_4903);
nand U1231 (N_1231,In_4159,In_1686);
nor U1232 (N_1232,In_1221,In_347);
or U1233 (N_1233,In_1318,In_3946);
or U1234 (N_1234,In_3317,In_1544);
nand U1235 (N_1235,In_275,In_3076);
nand U1236 (N_1236,In_4192,In_3898);
nand U1237 (N_1237,In_2048,In_1976);
xnor U1238 (N_1238,In_4379,In_3201);
and U1239 (N_1239,In_870,In_1939);
nand U1240 (N_1240,In_4402,In_4954);
or U1241 (N_1241,In_2321,In_4771);
nor U1242 (N_1242,In_1811,In_1015);
or U1243 (N_1243,In_2360,In_3986);
nand U1244 (N_1244,In_4893,In_3450);
xnor U1245 (N_1245,In_2022,In_949);
nor U1246 (N_1246,In_4938,In_2746);
nor U1247 (N_1247,In_4510,In_1805);
nand U1248 (N_1248,In_466,In_1426);
nand U1249 (N_1249,In_6,In_2858);
nor U1250 (N_1250,In_1343,In_1591);
xnor U1251 (N_1251,In_877,In_4886);
or U1252 (N_1252,In_3559,In_1422);
xor U1253 (N_1253,In_4686,In_1728);
xor U1254 (N_1254,In_2668,In_981);
and U1255 (N_1255,In_2059,In_3883);
or U1256 (N_1256,In_746,In_4281);
nor U1257 (N_1257,In_4722,In_2125);
nor U1258 (N_1258,In_609,In_2063);
nand U1259 (N_1259,In_4088,In_1966);
xnor U1260 (N_1260,In_4787,In_2049);
xnor U1261 (N_1261,In_2654,In_3255);
nor U1262 (N_1262,In_589,In_1520);
xor U1263 (N_1263,In_2824,In_4070);
and U1264 (N_1264,In_3053,In_3688);
and U1265 (N_1265,In_848,In_50);
nor U1266 (N_1266,In_528,In_3717);
xor U1267 (N_1267,In_703,In_1216);
nand U1268 (N_1268,In_247,In_1808);
xor U1269 (N_1269,In_4307,In_1717);
xor U1270 (N_1270,In_223,In_355);
or U1271 (N_1271,In_920,In_1053);
or U1272 (N_1272,In_640,In_1668);
xnor U1273 (N_1273,In_1691,In_3700);
nand U1274 (N_1274,In_3812,In_3740);
nand U1275 (N_1275,In_1338,In_227);
and U1276 (N_1276,In_1704,In_591);
xor U1277 (N_1277,In_806,In_4879);
nor U1278 (N_1278,In_2252,In_4636);
or U1279 (N_1279,In_3644,In_2051);
or U1280 (N_1280,In_4418,In_4724);
xnor U1281 (N_1281,In_1346,In_1839);
and U1282 (N_1282,In_3838,In_2702);
or U1283 (N_1283,In_4598,In_485);
nand U1284 (N_1284,In_1624,In_1227);
and U1285 (N_1285,In_535,In_4648);
nor U1286 (N_1286,In_2166,In_2918);
or U1287 (N_1287,In_1813,In_1295);
or U1288 (N_1288,In_4039,In_3576);
xnor U1289 (N_1289,In_2040,In_2473);
nand U1290 (N_1290,In_2990,In_2592);
xor U1291 (N_1291,In_1408,In_811);
and U1292 (N_1292,In_3826,In_4327);
nor U1293 (N_1293,In_1962,In_4299);
nand U1294 (N_1294,In_1751,In_323);
nor U1295 (N_1295,In_4882,In_3385);
nand U1296 (N_1296,In_4220,In_3379);
xor U1297 (N_1297,In_4055,In_695);
or U1298 (N_1298,In_1287,In_783);
and U1299 (N_1299,In_3966,In_4579);
nor U1300 (N_1300,In_2570,In_3952);
or U1301 (N_1301,In_2655,In_390);
and U1302 (N_1302,In_273,In_2427);
nor U1303 (N_1303,In_1739,In_962);
xor U1304 (N_1304,In_1656,In_2078);
xor U1305 (N_1305,In_1438,In_1150);
nor U1306 (N_1306,In_1904,In_114);
nor U1307 (N_1307,In_1684,In_2372);
xnor U1308 (N_1308,In_2399,In_4118);
and U1309 (N_1309,In_4305,In_1688);
nand U1310 (N_1310,In_1314,In_1434);
nor U1311 (N_1311,In_1681,In_448);
xnor U1312 (N_1312,In_1164,In_1750);
or U1313 (N_1313,In_3247,In_4362);
xor U1314 (N_1314,In_3924,In_2406);
nand U1315 (N_1315,In_2955,In_198);
xnor U1316 (N_1316,In_4166,In_737);
nor U1317 (N_1317,In_2880,In_2728);
or U1318 (N_1318,In_595,In_301);
and U1319 (N_1319,In_4112,In_1468);
or U1320 (N_1320,In_3921,In_363);
nor U1321 (N_1321,In_4109,In_2179);
or U1322 (N_1322,In_3712,In_3211);
and U1323 (N_1323,In_1644,In_3668);
and U1324 (N_1324,In_3127,In_1448);
xor U1325 (N_1325,In_3392,In_479);
nor U1326 (N_1326,In_3797,In_4947);
nand U1327 (N_1327,In_537,In_4476);
and U1328 (N_1328,In_3997,In_901);
or U1329 (N_1329,In_260,In_0);
nand U1330 (N_1330,In_1553,In_2557);
or U1331 (N_1331,In_4231,In_694);
nand U1332 (N_1332,In_1900,In_2846);
or U1333 (N_1333,In_2280,In_80);
nor U1334 (N_1334,In_1662,In_2612);
nor U1335 (N_1335,In_3223,In_296);
nor U1336 (N_1336,In_1270,In_1822);
or U1337 (N_1337,In_1848,In_2551);
nand U1338 (N_1338,In_2879,In_3432);
nor U1339 (N_1339,In_4139,In_572);
xor U1340 (N_1340,In_740,In_2303);
nand U1341 (N_1341,In_2744,In_1867);
or U1342 (N_1342,In_1525,In_3342);
and U1343 (N_1343,In_1581,In_258);
xor U1344 (N_1344,In_1804,In_3377);
nand U1345 (N_1345,In_2151,In_3407);
and U1346 (N_1346,In_2525,In_2797);
or U1347 (N_1347,In_3330,In_1981);
nand U1348 (N_1348,In_751,In_4368);
and U1349 (N_1349,In_2157,In_3015);
xnor U1350 (N_1350,In_3414,In_4995);
nor U1351 (N_1351,In_3666,In_918);
or U1352 (N_1352,In_2650,In_1788);
and U1353 (N_1353,In_1163,In_3164);
and U1354 (N_1354,In_1372,In_1871);
xor U1355 (N_1355,In_4178,In_2733);
nand U1356 (N_1356,In_3140,In_3626);
or U1357 (N_1357,In_3945,In_4457);
and U1358 (N_1358,In_3880,In_3850);
and U1359 (N_1359,In_1925,In_56);
and U1360 (N_1360,In_3104,In_3193);
or U1361 (N_1361,In_1806,In_4187);
xnor U1362 (N_1362,In_2304,In_2246);
xor U1363 (N_1363,In_4123,In_2062);
nor U1364 (N_1364,In_2086,In_4831);
and U1365 (N_1365,In_3036,In_1560);
nand U1366 (N_1366,In_1921,In_122);
and U1367 (N_1367,In_2264,In_4524);
xnor U1368 (N_1368,In_789,In_4816);
xnor U1369 (N_1369,In_2149,In_4791);
nor U1370 (N_1370,In_3249,In_2364);
and U1371 (N_1371,In_173,In_2395);
and U1372 (N_1372,In_1996,In_4248);
or U1373 (N_1373,In_1388,In_2653);
or U1374 (N_1374,In_4149,In_3689);
nand U1375 (N_1375,In_4037,In_433);
xnor U1376 (N_1376,In_3692,In_4376);
nand U1377 (N_1377,In_2505,In_191);
and U1378 (N_1378,In_3485,In_766);
nand U1379 (N_1379,In_3981,In_3369);
or U1380 (N_1380,In_3926,In_882);
nor U1381 (N_1381,In_4181,In_219);
and U1382 (N_1382,In_4297,In_3080);
xnor U1383 (N_1383,In_2100,In_850);
nor U1384 (N_1384,In_3309,In_4453);
nand U1385 (N_1385,In_2672,In_1319);
nand U1386 (N_1386,In_4604,In_4345);
nand U1387 (N_1387,In_3999,In_3356);
nand U1388 (N_1388,In_1803,In_1856);
and U1389 (N_1389,In_2103,In_2507);
nor U1390 (N_1390,In_3661,In_4924);
nand U1391 (N_1391,In_632,In_4257);
and U1392 (N_1392,In_161,In_4506);
xnor U1393 (N_1393,In_2932,In_1584);
or U1394 (N_1394,In_2198,In_75);
nand U1395 (N_1395,In_2552,In_2661);
nand U1396 (N_1396,In_1020,In_907);
and U1397 (N_1397,In_4846,In_1973);
nor U1398 (N_1398,In_310,In_459);
and U1399 (N_1399,In_4928,In_3349);
or U1400 (N_1400,In_1197,In_1671);
xor U1401 (N_1401,In_3935,In_1055);
xor U1402 (N_1402,In_1115,In_4731);
or U1403 (N_1403,In_1169,In_4078);
nor U1404 (N_1404,In_2432,In_3897);
and U1405 (N_1405,In_398,In_1600);
xor U1406 (N_1406,In_2223,In_2864);
and U1407 (N_1407,In_2889,In_3284);
or U1408 (N_1408,In_4849,In_3436);
and U1409 (N_1409,In_4560,In_1736);
or U1410 (N_1410,In_1650,In_1580);
and U1411 (N_1411,In_305,In_2532);
or U1412 (N_1412,In_125,In_733);
xor U1413 (N_1413,In_1561,In_1037);
nor U1414 (N_1414,In_3090,In_4675);
nor U1415 (N_1415,In_2208,In_3660);
nand U1416 (N_1416,In_1455,In_1901);
xnor U1417 (N_1417,In_723,In_1498);
xnor U1418 (N_1418,In_3802,In_669);
nand U1419 (N_1419,In_1969,In_3520);
and U1420 (N_1420,In_2370,In_1755);
and U1421 (N_1421,In_214,In_4203);
and U1422 (N_1422,In_2837,In_424);
nor U1423 (N_1423,In_2057,In_3028);
nor U1424 (N_1424,In_1914,In_593);
and U1425 (N_1425,In_2681,In_4732);
or U1426 (N_1426,In_536,In_2195);
nor U1427 (N_1427,In_1640,In_3589);
nand U1428 (N_1428,In_2441,In_3348);
nor U1429 (N_1429,In_4904,In_4941);
xnor U1430 (N_1430,In_614,In_3165);
and U1431 (N_1431,In_1960,In_1613);
nor U1432 (N_1432,In_3268,In_4975);
nor U1433 (N_1433,In_1489,In_252);
or U1434 (N_1434,In_3938,In_3621);
xnor U1435 (N_1435,In_2274,In_673);
or U1436 (N_1436,In_4783,In_611);
or U1437 (N_1437,In_1172,In_3551);
xnor U1438 (N_1438,In_2699,In_4117);
xnor U1439 (N_1439,In_3554,In_4128);
and U1440 (N_1440,In_3048,In_4333);
and U1441 (N_1441,In_4523,In_681);
xor U1442 (N_1442,In_3328,In_4610);
xnor U1443 (N_1443,In_1638,In_4026);
nor U1444 (N_1444,In_2096,In_3234);
and U1445 (N_1445,In_4018,In_2251);
xnor U1446 (N_1446,In_2327,In_3879);
nor U1447 (N_1447,In_3386,In_2549);
and U1448 (N_1448,In_865,In_680);
xnor U1449 (N_1449,In_720,In_4047);
and U1450 (N_1450,In_852,In_4711);
nand U1451 (N_1451,In_24,In_4399);
nand U1452 (N_1452,In_2644,In_2184);
nand U1453 (N_1453,In_4525,In_4687);
nand U1454 (N_1454,In_2679,In_1239);
nand U1455 (N_1455,In_1858,In_1154);
and U1456 (N_1456,In_4872,In_3599);
nand U1457 (N_1457,In_86,In_26);
and U1458 (N_1458,In_1410,In_4022);
nor U1459 (N_1459,In_4448,In_1481);
nor U1460 (N_1460,In_3581,In_1204);
and U1461 (N_1461,In_22,In_2244);
nand U1462 (N_1462,In_3362,In_4822);
nor U1463 (N_1463,In_3215,In_4720);
xnor U1464 (N_1464,In_1281,In_4989);
and U1465 (N_1465,In_3017,In_3817);
nor U1466 (N_1466,In_3443,In_391);
nand U1467 (N_1467,In_4349,In_2456);
nand U1468 (N_1468,In_1240,In_210);
nand U1469 (N_1469,In_3541,In_2967);
nand U1470 (N_1470,In_437,In_971);
nand U1471 (N_1471,In_446,In_3353);
nand U1472 (N_1472,In_4752,In_4585);
nor U1473 (N_1473,In_1592,In_684);
xor U1474 (N_1474,In_923,In_205);
and U1475 (N_1475,In_3233,In_4913);
and U1476 (N_1476,In_802,In_1368);
nor U1477 (N_1477,In_4718,In_1534);
nand U1478 (N_1478,In_2217,In_3440);
nor U1479 (N_1479,In_3489,In_3620);
nand U1480 (N_1480,In_4838,In_4363);
and U1481 (N_1481,In_1826,In_1655);
or U1482 (N_1482,In_2794,In_508);
or U1483 (N_1483,In_1916,In_2684);
and U1484 (N_1484,In_3331,In_1819);
or U1485 (N_1485,In_28,In_3641);
or U1486 (N_1486,In_912,In_204);
and U1487 (N_1487,In_857,In_603);
and U1488 (N_1488,In_582,In_3911);
nand U1489 (N_1489,In_2489,In_2520);
and U1490 (N_1490,In_2758,In_4148);
xnor U1491 (N_1491,In_1575,In_1490);
xnor U1492 (N_1492,In_3381,In_2928);
nor U1493 (N_1493,In_2972,In_1894);
and U1494 (N_1494,In_2760,In_3865);
or U1495 (N_1495,In_2984,In_2161);
nand U1496 (N_1496,In_2603,In_4495);
xnor U1497 (N_1497,In_3949,In_2855);
xnor U1498 (N_1498,In_3825,In_1398);
xor U1499 (N_1499,In_4768,In_3564);
or U1500 (N_1500,In_4747,In_523);
nor U1501 (N_1501,In_1703,In_1463);
nand U1502 (N_1502,In_3806,In_4429);
and U1503 (N_1503,In_665,In_3137);
nand U1504 (N_1504,In_4962,In_418);
nand U1505 (N_1505,In_319,In_3505);
xnor U1506 (N_1506,In_1630,In_3488);
xnor U1507 (N_1507,In_2856,In_4895);
nand U1508 (N_1508,In_4898,In_4883);
nand U1509 (N_1509,In_3288,In_2664);
nand U1510 (N_1510,In_902,In_4310);
nand U1511 (N_1511,In_4500,In_108);
xnor U1512 (N_1512,In_3064,In_3769);
nand U1513 (N_1513,In_953,In_2585);
and U1514 (N_1514,In_2074,In_4329);
nand U1515 (N_1515,In_4857,In_526);
nand U1516 (N_1516,In_2906,In_2351);
nand U1517 (N_1517,In_136,In_2434);
and U1518 (N_1518,In_671,In_4161);
or U1519 (N_1519,In_4757,In_1246);
nor U1520 (N_1520,In_546,In_828);
nand U1521 (N_1521,In_4602,In_2753);
nor U1522 (N_1522,In_4684,In_3427);
xor U1523 (N_1523,In_1074,In_165);
nor U1524 (N_1524,In_4998,In_3395);
and U1525 (N_1525,In_4607,In_4244);
xnor U1526 (N_1526,In_2968,In_2201);
or U1527 (N_1527,In_4091,In_1294);
xor U1528 (N_1528,In_4443,In_564);
or U1529 (N_1529,In_3777,In_1306);
or U1530 (N_1530,In_575,In_658);
nand U1531 (N_1531,In_4577,In_1955);
nor U1532 (N_1532,In_4325,In_4330);
nor U1533 (N_1533,In_1202,In_4991);
xor U1534 (N_1534,In_4447,In_2188);
xor U1535 (N_1535,In_986,In_2721);
and U1536 (N_1536,In_3256,In_1509);
or U1537 (N_1537,In_1832,In_4395);
and U1538 (N_1538,In_4015,In_2175);
nand U1539 (N_1539,In_1193,In_4493);
xor U1540 (N_1540,In_2133,In_2352);
and U1541 (N_1541,In_583,In_4060);
or U1542 (N_1542,In_2060,In_3483);
or U1543 (N_1543,In_442,In_4321);
nor U1544 (N_1544,In_4744,In_284);
nor U1545 (N_1545,In_3147,In_1620);
and U1546 (N_1546,In_1379,In_3881);
and U1547 (N_1547,In_1186,In_4884);
or U1548 (N_1548,In_2854,In_2614);
or U1549 (N_1549,In_1320,In_982);
nor U1550 (N_1550,In_3786,In_2950);
xor U1551 (N_1551,In_4477,In_1527);
nand U1552 (N_1552,In_1198,In_2716);
xnor U1553 (N_1553,In_1049,In_458);
xnor U1554 (N_1554,In_2241,In_371);
nor U1555 (N_1555,In_1362,In_4795);
nand U1556 (N_1556,In_2178,In_707);
nand U1557 (N_1557,In_4517,In_1365);
and U1558 (N_1558,In_4917,In_1846);
nand U1559 (N_1559,In_4658,In_4366);
xor U1560 (N_1560,In_1311,In_2629);
nand U1561 (N_1561,In_3218,In_2420);
or U1562 (N_1562,In_1505,In_1912);
nor U1563 (N_1563,In_1618,In_2160);
or U1564 (N_1564,In_2262,In_3374);
nor U1565 (N_1565,In_1264,In_1907);
nand U1566 (N_1566,In_4253,In_2793);
nand U1567 (N_1567,In_2089,In_46);
or U1568 (N_1568,In_3046,In_4338);
and U1569 (N_1569,In_2573,In_2818);
and U1570 (N_1570,In_2615,In_4657);
nand U1571 (N_1571,In_3016,In_1262);
nand U1572 (N_1572,In_3604,In_3220);
nand U1573 (N_1573,In_769,In_2088);
or U1574 (N_1574,In_1967,In_4801);
nand U1575 (N_1575,In_2769,In_1559);
nor U1576 (N_1576,In_3122,In_1645);
or U1577 (N_1577,In_4068,In_660);
xor U1578 (N_1578,In_714,In_4312);
nor U1579 (N_1579,In_2347,In_131);
xor U1580 (N_1580,In_2156,In_3024);
or U1581 (N_1581,In_292,In_2712);
nor U1582 (N_1582,In_4559,In_1885);
nor U1583 (N_1583,In_2137,In_4274);
and U1584 (N_1584,In_1601,In_3209);
nor U1585 (N_1585,In_1064,In_1506);
nor U1586 (N_1586,In_4108,In_3106);
nand U1587 (N_1587,In_3276,In_3398);
or U1588 (N_1588,In_444,In_3197);
nor U1589 (N_1589,In_181,In_1153);
nor U1590 (N_1590,In_2757,In_3767);
nor U1591 (N_1591,In_1794,In_2907);
nor U1592 (N_1592,In_3680,In_4216);
nor U1593 (N_1593,In_1547,In_2154);
xnor U1594 (N_1594,In_3979,In_1446);
xnor U1595 (N_1595,In_1415,In_947);
or U1596 (N_1596,In_4987,In_4455);
xnor U1597 (N_1597,In_3321,In_4753);
and U1598 (N_1598,In_2761,In_2843);
xnor U1599 (N_1599,In_364,In_1852);
nor U1600 (N_1600,In_2673,In_3699);
and U1601 (N_1601,In_610,In_3422);
or U1602 (N_1602,In_701,In_2397);
or U1603 (N_1603,In_2253,In_4784);
nor U1604 (N_1604,In_1165,In_4932);
and U1605 (N_1605,In_1913,In_241);
and U1606 (N_1606,In_644,In_594);
or U1607 (N_1607,In_867,In_1425);
or U1608 (N_1608,In_1040,In_457);
or U1609 (N_1609,In_4234,In_158);
and U1610 (N_1610,In_4300,In_2047);
xnor U1611 (N_1611,In_354,In_3914);
or U1612 (N_1612,In_3431,In_2065);
nor U1613 (N_1613,In_1348,In_533);
nor U1614 (N_1614,In_492,In_1568);
xor U1615 (N_1615,In_3060,In_4285);
or U1616 (N_1616,In_4255,In_4306);
nor U1617 (N_1617,In_3875,In_2809);
or U1618 (N_1618,In_697,In_103);
xnor U1619 (N_1619,In_739,In_4869);
xnor U1620 (N_1620,In_2448,In_1494);
xor U1621 (N_1621,In_933,In_2412);
or U1622 (N_1622,In_2258,In_1905);
nand U1623 (N_1623,In_2865,In_3225);
and U1624 (N_1624,In_4439,In_3518);
nor U1625 (N_1625,In_1285,In_1497);
and U1626 (N_1626,In_1128,In_2454);
or U1627 (N_1627,In_2021,In_678);
or U1628 (N_1628,In_4378,In_2956);
nand U1629 (N_1629,In_1435,In_2578);
and U1630 (N_1630,In_4937,In_2028);
and U1631 (N_1631,In_1707,In_1327);
or U1632 (N_1632,In_1237,In_2174);
and U1633 (N_1633,In_106,In_326);
nor U1634 (N_1634,In_2643,In_461);
xor U1635 (N_1635,In_4219,In_2041);
xor U1636 (N_1636,In_2951,In_4874);
or U1637 (N_1637,In_3179,In_2218);
nand U1638 (N_1638,In_3444,In_3859);
nand U1639 (N_1639,In_4184,In_1875);
and U1640 (N_1640,In_4208,In_3818);
or U1641 (N_1641,In_1048,In_750);
nor U1642 (N_1642,In_2586,In_4264);
nand U1643 (N_1643,In_1646,In_3633);
nand U1644 (N_1644,In_3904,In_726);
nand U1645 (N_1645,In_3013,In_2778);
nor U1646 (N_1646,In_817,In_65);
xnor U1647 (N_1647,In_387,In_1469);
or U1648 (N_1648,In_3552,In_4566);
or U1649 (N_1649,In_3457,In_1004);
or U1650 (N_1650,In_2362,In_4124);
and U1651 (N_1651,In_3061,In_3718);
nor U1652 (N_1652,In_3665,In_20);
xnor U1653 (N_1653,In_4475,In_762);
nand U1654 (N_1654,In_3301,In_454);
xor U1655 (N_1655,In_2345,In_3893);
nor U1656 (N_1656,In_1116,In_4630);
and U1657 (N_1657,In_3340,In_890);
xnor U1658 (N_1658,In_4302,In_637);
and U1659 (N_1659,In_1044,In_3474);
or U1660 (N_1660,In_1088,In_467);
xnor U1661 (N_1661,In_2290,In_4188);
and U1662 (N_1662,In_3800,In_2784);
or U1663 (N_1663,In_1777,In_1555);
xor U1664 (N_1664,In_3964,In_4390);
or U1665 (N_1665,In_974,In_3710);
or U1666 (N_1666,In_3263,In_1329);
and U1667 (N_1667,In_1884,In_1332);
nor U1668 (N_1668,In_2245,In_253);
xnor U1669 (N_1669,In_1602,In_4167);
and U1670 (N_1670,In_557,In_796);
or U1671 (N_1671,In_3741,In_841);
nor U1672 (N_1672,In_3130,In_1579);
xor U1673 (N_1673,In_2281,In_1255);
nor U1674 (N_1674,In_3346,In_599);
or U1675 (N_1675,In_1084,In_2367);
nor U1676 (N_1676,In_3086,In_3854);
xor U1677 (N_1677,In_1594,In_263);
nor U1678 (N_1678,In_94,In_3537);
nor U1679 (N_1679,In_2491,In_4005);
nor U1680 (N_1680,In_4097,In_3780);
or U1681 (N_1681,In_98,In_1989);
or U1682 (N_1682,In_4177,In_2975);
and U1683 (N_1683,In_1083,In_4655);
or U1684 (N_1684,In_1059,In_2182);
nor U1685 (N_1685,In_2759,In_2828);
nor U1686 (N_1686,In_958,In_4863);
and U1687 (N_1687,In_2502,In_1195);
and U1688 (N_1688,In_3120,In_851);
nand U1689 (N_1689,In_1374,In_2470);
or U1690 (N_1690,In_1466,In_333);
nand U1691 (N_1691,In_4030,In_919);
and U1692 (N_1692,In_322,In_2698);
nand U1693 (N_1693,In_2842,In_856);
or U1694 (N_1694,In_3166,In_4859);
or U1695 (N_1695,In_2626,In_4388);
nor U1696 (N_1696,In_4522,In_1541);
nand U1697 (N_1697,In_4436,In_668);
or U1698 (N_1698,In_830,In_4021);
nand U1699 (N_1699,In_4446,In_4944);
nor U1700 (N_1700,In_3487,In_568);
xor U1701 (N_1701,In_3912,In_402);
and U1702 (N_1702,In_3191,In_4806);
nor U1703 (N_1703,In_639,In_2973);
nor U1704 (N_1704,In_3645,In_654);
and U1705 (N_1705,In_484,In_2565);
nor U1706 (N_1706,In_3525,In_4621);
xnor U1707 (N_1707,In_1126,In_655);
nor U1708 (N_1708,In_2020,In_4837);
nor U1709 (N_1709,In_3728,In_325);
nor U1710 (N_1710,In_2424,In_616);
and U1711 (N_1711,In_2292,In_4999);
and U1712 (N_1712,In_3477,In_3549);
xor U1713 (N_1713,In_2666,In_4974);
nand U1714 (N_1714,In_215,In_2633);
and U1715 (N_1715,In_142,In_4044);
nand U1716 (N_1716,In_505,In_3439);
and U1717 (N_1717,In_3696,In_105);
xor U1718 (N_1718,In_1136,In_2987);
or U1719 (N_1719,In_2860,In_2952);
xor U1720 (N_1720,In_3572,In_4881);
and U1721 (N_1721,In_1349,In_1511);
nor U1722 (N_1722,In_3023,In_963);
or U1723 (N_1723,In_2798,In_186);
or U1724 (N_1724,In_419,In_553);
nor U1725 (N_1725,In_2914,In_1207);
or U1726 (N_1726,In_3684,In_346);
xnor U1727 (N_1727,In_2330,In_948);
xor U1728 (N_1728,In_2887,In_922);
or U1729 (N_1729,In_2826,In_426);
or U1730 (N_1730,In_772,In_1629);
xnor U1731 (N_1731,In_1522,In_3279);
and U1732 (N_1732,In_3213,In_4162);
xor U1733 (N_1733,In_4955,In_4618);
and U1734 (N_1734,In_1133,In_929);
and U1735 (N_1735,In_394,In_2085);
or U1736 (N_1736,In_1277,In_2455);
or U1737 (N_1737,In_2581,In_2388);
nor U1738 (N_1738,In_4542,In_3839);
or U1739 (N_1739,In_1219,In_1539);
nor U1740 (N_1740,In_1661,In_1797);
and U1741 (N_1741,In_3636,In_975);
nand U1742 (N_1742,In_4096,In_4830);
nor U1743 (N_1743,In_4092,In_3069);
or U1744 (N_1744,In_148,In_9);
or U1745 (N_1745,In_988,In_3890);
or U1746 (N_1746,In_606,In_1371);
and U1747 (N_1747,In_3873,In_2031);
nor U1748 (N_1748,In_3399,In_2254);
nand U1749 (N_1749,In_4322,In_4889);
and U1750 (N_1750,In_3616,In_3171);
nand U1751 (N_1751,In_34,In_4563);
xnor U1752 (N_1752,In_1129,In_1400);
or U1753 (N_1753,In_1375,In_3281);
nand U1754 (N_1754,In_1637,In_3093);
nand U1755 (N_1755,In_3593,In_674);
nor U1756 (N_1756,In_4691,In_1605);
or U1757 (N_1757,In_2566,In_3097);
or U1758 (N_1758,In_4122,In_527);
or U1759 (N_1759,In_4983,In_754);
or U1760 (N_1760,In_573,In_411);
nand U1761 (N_1761,In_1021,In_4513);
xor U1762 (N_1762,In_1232,In_2994);
and U1763 (N_1763,In_3452,In_2114);
or U1764 (N_1764,In_2263,In_4474);
and U1765 (N_1765,In_816,In_1047);
xor U1766 (N_1766,In_617,In_1844);
nand U1767 (N_1767,In_31,In_1326);
and U1768 (N_1768,In_74,In_4011);
and U1769 (N_1769,In_61,In_3605);
nor U1770 (N_1770,In_3874,In_2804);
nor U1771 (N_1771,In_1288,In_4672);
and U1772 (N_1772,In_298,In_2576);
nor U1773 (N_1773,In_776,In_556);
nand U1774 (N_1774,In_460,In_649);
xnor U1775 (N_1775,In_4545,In_465);
nor U1776 (N_1776,In_1935,In_2588);
xor U1777 (N_1777,In_4158,In_3674);
nand U1778 (N_1778,In_4176,In_4915);
or U1779 (N_1779,In_3727,In_2720);
or U1780 (N_1780,In_3969,In_1790);
xor U1781 (N_1781,In_1205,In_1882);
nand U1782 (N_1782,In_1038,In_1073);
and U1783 (N_1783,In_3900,In_110);
or U1784 (N_1784,In_2556,In_4472);
nor U1785 (N_1785,In_208,In_4876);
nor U1786 (N_1786,In_1290,In_3594);
nor U1787 (N_1787,In_3098,In_4901);
xor U1788 (N_1788,In_1124,In_2110);
nor U1789 (N_1789,In_3994,In_4984);
or U1790 (N_1790,In_1833,In_2255);
xnor U1791 (N_1791,In_469,In_4745);
and U1792 (N_1792,In_618,In_1634);
and U1793 (N_1793,In_340,In_4841);
or U1794 (N_1794,In_1323,In_2152);
nor U1795 (N_1795,In_4562,In_464);
or U1796 (N_1796,In_3168,In_58);
xnor U1797 (N_1797,In_3754,In_3514);
nor U1798 (N_1798,In_4492,In_2082);
and U1799 (N_1799,In_3435,In_3192);
nor U1800 (N_1800,In_930,In_884);
nor U1801 (N_1801,In_1413,In_972);
xor U1802 (N_1802,In_1366,In_4969);
nand U1803 (N_1803,In_1793,In_4982);
and U1804 (N_1804,In_3630,In_2488);
nor U1805 (N_1805,In_2680,In_4885);
and U1806 (N_1806,In_3906,In_2982);
nor U1807 (N_1807,In_2613,In_2450);
nor U1808 (N_1808,In_1585,In_1328);
or U1809 (N_1809,In_689,In_855);
and U1810 (N_1810,In_1908,In_4106);
and U1811 (N_1811,In_4505,In_1621);
and U1812 (N_1812,In_410,In_1307);
nand U1813 (N_1813,In_2306,In_4190);
and U1814 (N_1814,In_4358,In_1011);
nor U1815 (N_1815,In_4945,In_3337);
xnor U1816 (N_1816,In_8,In_1664);
nand U1817 (N_1817,In_1325,In_3570);
xor U1818 (N_1818,In_4704,In_1401);
or U1819 (N_1819,In_1576,In_524);
xnor U1820 (N_1820,In_149,In_2897);
and U1821 (N_1821,In_190,In_985);
or U1822 (N_1822,In_167,In_4036);
nand U1823 (N_1823,In_4009,In_3447);
nor U1824 (N_1824,In_1142,In_2439);
xnor U1825 (N_1825,In_4550,In_1244);
and U1826 (N_1826,In_946,In_2273);
and U1827 (N_1827,In_4469,In_786);
xnor U1828 (N_1828,In_1035,In_1002);
nand U1829 (N_1829,In_4343,In_4789);
xnor U1830 (N_1830,In_3082,In_1390);
xnor U1831 (N_1831,In_2670,In_940);
nor U1832 (N_1832,In_3509,In_1459);
nor U1833 (N_1833,In_3293,In_2163);
nand U1834 (N_1834,In_2772,In_336);
and U1835 (N_1835,In_3155,In_2069);
xnor U1836 (N_1836,In_2577,In_3274);
or U1837 (N_1837,In_2701,In_3079);
nand U1838 (N_1838,In_3437,In_48);
nand U1839 (N_1839,In_1418,In_1807);
xnor U1840 (N_1840,In_374,In_3656);
or U1841 (N_1841,In_1041,In_377);
nor U1842 (N_1842,In_3270,In_4478);
nor U1843 (N_1843,In_4642,In_3116);
xnor U1844 (N_1844,In_2584,In_732);
nand U1845 (N_1845,In_2734,In_2437);
and U1846 (N_1846,In_3178,In_4639);
xnor U1847 (N_1847,In_1533,In_1447);
or U1848 (N_1848,In_4840,In_4755);
or U1849 (N_1849,In_1112,In_3869);
nand U1850 (N_1850,In_4596,In_2678);
and U1851 (N_1851,In_4557,In_781);
xor U1852 (N_1852,In_1258,In_4318);
nor U1853 (N_1853,In_1598,In_1874);
xor U1854 (N_1854,In_3380,In_3207);
xnor U1855 (N_1855,In_3325,In_259);
nor U1856 (N_1856,In_4367,In_3799);
xor U1857 (N_1857,In_2054,In_4282);
nor U1858 (N_1858,In_2574,In_4445);
or U1859 (N_1859,In_917,In_4125);
nand U1860 (N_1860,In_1006,In_2224);
xor U1861 (N_1861,In_3417,In_3389);
nor U1862 (N_1862,In_3318,In_69);
and U1863 (N_1863,In_4971,In_3532);
or U1864 (N_1864,In_2202,In_230);
or U1865 (N_1865,In_2302,In_4066);
and U1866 (N_1866,In_2799,In_4484);
xnor U1867 (N_1867,In_4671,In_1417);
and U1868 (N_1868,In_4043,In_2976);
and U1869 (N_1869,In_3084,In_2425);
xnor U1870 (N_1870,In_4280,In_834);
and U1871 (N_1871,In_4424,In_579);
xor U1872 (N_1872,In_4452,In_3944);
and U1873 (N_1873,In_1521,In_810);
nor U1874 (N_1874,In_405,In_4267);
nand U1875 (N_1875,In_2667,In_942);
and U1876 (N_1876,In_2369,In_1147);
or U1877 (N_1877,In_2260,In_3862);
nor U1878 (N_1878,In_4582,In_2785);
nor U1879 (N_1879,In_3449,In_3950);
xnor U1880 (N_1880,In_3434,In_4243);
or U1881 (N_1881,In_683,In_2537);
or U1882 (N_1882,In_4435,In_1104);
xor U1883 (N_1883,In_3087,In_4535);
nand U1884 (N_1884,In_1982,In_519);
nor U1885 (N_1885,In_3959,In_3970);
nor U1886 (N_1886,In_2050,In_3638);
xnor U1887 (N_1887,In_2324,In_329);
or U1888 (N_1888,In_1625,In_770);
xor U1889 (N_1889,In_4824,In_2365);
or U1890 (N_1890,In_4396,In_2852);
or U1891 (N_1891,In_455,In_1617);
nor U1892 (N_1892,In_1873,In_1367);
and U1893 (N_1893,In_2531,In_2874);
xnor U1894 (N_1894,In_1022,In_3460);
or U1895 (N_1895,In_3059,In_2708);
and U1896 (N_1896,In_2965,In_2014);
nand U1897 (N_1897,In_874,In_837);
or U1898 (N_1898,In_3771,In_150);
xnor U1899 (N_1899,In_3635,In_4023);
xor U1900 (N_1900,In_676,In_2736);
xor U1901 (N_1901,In_822,In_1769);
and U1902 (N_1902,In_1861,In_1312);
and U1903 (N_1903,In_456,In_2737);
nand U1904 (N_1904,In_1079,In_4823);
and U1905 (N_1905,In_4778,In_4914);
and U1906 (N_1906,In_3683,In_441);
and U1907 (N_1907,In_934,In_2270);
nand U1908 (N_1908,In_3613,In_562);
xor U1909 (N_1909,In_1857,In_4568);
or U1910 (N_1910,In_718,In_475);
nor U1911 (N_1911,In_2942,In_2550);
or U1912 (N_1912,In_3655,In_3227);
nand U1913 (N_1913,In_2773,In_4536);
and U1914 (N_1914,In_2528,In_3663);
or U1915 (N_1915,In_540,In_3057);
nand U1916 (N_1916,In_1111,In_709);
xor U1917 (N_1917,In_4851,In_4908);
nand U1918 (N_1918,In_3214,In_1066);
nand U1919 (N_1919,In_2194,In_3778);
or U1920 (N_1920,In_361,In_518);
or U1921 (N_1921,In_375,In_2687);
nand U1922 (N_1922,In_4470,In_220);
and U1923 (N_1923,In_2107,In_4774);
and U1924 (N_1924,In_823,In_2477);
xnor U1925 (N_1925,In_3495,In_1183);
nor U1926 (N_1926,In_2511,In_3708);
and U1927 (N_1927,In_3984,In_3125);
nor U1928 (N_1928,In_3329,In_4633);
and U1929 (N_1929,In_2392,In_3152);
or U1930 (N_1930,In_3975,In_2671);
xnor U1931 (N_1931,In_2820,In_4725);
and U1932 (N_1932,In_1957,In_3973);
and U1933 (N_1933,In_4133,In_3586);
or U1934 (N_1934,In_3430,In_3158);
nor U1935 (N_1935,In_1781,In_1175);
xor U1936 (N_1936,In_3203,In_2875);
nor U1937 (N_1937,In_1628,In_1767);
xnor U1938 (N_1938,In_1429,In_2211);
and U1939 (N_1939,In_3230,In_3753);
nand U1940 (N_1940,In_2109,In_1647);
and U1941 (N_1941,In_597,In_4464);
or U1942 (N_1942,In_3219,In_3200);
or U1943 (N_1943,In_3947,In_238);
or U1944 (N_1944,In_1672,In_62);
or U1945 (N_1945,In_2428,In_1689);
and U1946 (N_1946,In_1077,In_956);
nor U1947 (N_1947,In_1699,In_172);
nand U1948 (N_1948,In_4292,In_434);
xor U1949 (N_1949,In_2960,In_3397);
or U1950 (N_1950,In_366,In_4854);
nand U1951 (N_1951,In_2866,In_4734);
xnor U1952 (N_1952,In_650,In_4339);
or U1953 (N_1953,In_2243,In_4651);
or U1954 (N_1954,In_1464,In_2012);
and U1955 (N_1955,In_1678,In_493);
or U1956 (N_1956,In_1993,In_590);
nand U1957 (N_1957,In_4812,In_4640);
or U1958 (N_1958,In_3619,In_3639);
nand U1959 (N_1959,In_2144,In_4201);
xnor U1960 (N_1960,In_831,In_4597);
and U1961 (N_1961,In_365,In_43);
and U1962 (N_1962,In_3315,In_2469);
nor U1963 (N_1963,In_392,In_1663);
xnor U1964 (N_1964,In_3186,In_4170);
nand U1965 (N_1965,In_3980,In_55);
nand U1966 (N_1966,In_2440,In_4273);
xor U1967 (N_1967,In_2269,In_4501);
xnor U1968 (N_1968,In_812,In_2642);
nand U1969 (N_1969,In_3597,In_4156);
nand U1970 (N_1970,In_2898,In_4440);
nor U1971 (N_1971,In_1859,In_1523);
nand U1972 (N_1972,In_1714,In_1421);
nand U1973 (N_1973,In_4263,In_1604);
and U1974 (N_1974,In_4434,In_3052);
or U1975 (N_1975,In_699,In_3129);
and U1976 (N_1976,In_4894,In_2115);
nand U1977 (N_1977,In_3650,In_1095);
nor U1978 (N_1978,In_1720,In_474);
nand U1979 (N_1979,In_2102,In_3652);
nand U1980 (N_1980,In_1499,In_1377);
xnor U1981 (N_1981,In_4016,In_2740);
nand U1982 (N_1982,In_1316,In_2908);
or U1983 (N_1983,In_261,In_42);
and U1984 (N_1984,In_3845,In_1280);
and U1985 (N_1985,In_2548,In_1831);
and U1986 (N_1986,In_1188,In_4175);
or U1987 (N_1987,In_134,In_3361);
nor U1988 (N_1988,In_423,In_1026);
and U1989 (N_1989,In_2819,In_4209);
xor U1990 (N_1990,In_4591,In_331);
or U1991 (N_1991,In_1203,In_3299);
nand U1992 (N_1992,In_1947,In_3429);
nor U1993 (N_1993,In_1876,In_1152);
xnor U1994 (N_1994,In_2203,In_3077);
and U1995 (N_1995,In_3099,In_4912);
nand U1996 (N_1996,In_4754,In_4196);
and U1997 (N_1997,In_2058,In_1599);
and U1998 (N_1998,In_998,In_2920);
or U1999 (N_1999,In_980,In_3479);
nand U2000 (N_2000,In_1063,In_4245);
or U2001 (N_2001,In_1890,In_3128);
nor U2002 (N_2002,In_3894,In_3396);
or U2003 (N_2003,In_4001,In_380);
and U2004 (N_2004,In_925,In_3631);
nor U2005 (N_2005,In_4759,In_217);
nor U2006 (N_2006,In_3899,In_4172);
nor U2007 (N_2007,In_3376,In_4041);
xor U2008 (N_2008,In_832,In_264);
or U2009 (N_2009,In_3951,In_4213);
xor U2010 (N_2010,In_1385,In_2240);
xnor U2011 (N_2011,In_924,In_3010);
nand U2012 (N_2012,In_761,In_4605);
xor U2013 (N_2013,In_4254,In_1478);
xor U2014 (N_2014,In_3034,In_3047);
and U2015 (N_2015,In_4710,In_3528);
nor U2016 (N_2016,In_3151,In_936);
xor U2017 (N_2017,In_2038,In_4270);
or U2018 (N_2018,In_3294,In_4782);
nor U2019 (N_2019,In_4102,In_4129);
xor U2020 (N_2020,In_4980,In_1572);
and U2021 (N_2021,In_4276,In_3731);
nand U2022 (N_2022,In_1778,In_1619);
nand U2023 (N_2023,In_4538,In_1427);
and U2024 (N_2024,In_113,In_4291);
or U2025 (N_2025,In_891,In_281);
nand U2026 (N_2026,In_4421,In_2872);
and U2027 (N_2027,In_2539,In_4033);
nand U2028 (N_2028,In_4360,In_2568);
nor U2029 (N_2029,In_3648,In_1068);
nand U2030 (N_2030,In_3892,In_285);
or U2031 (N_2031,In_1849,In_3903);
or U2032 (N_2032,In_4986,In_2034);
nor U2033 (N_2033,In_115,In_1089);
or U2034 (N_2034,In_3237,In_4650);
nor U2035 (N_2035,In_2954,In_3795);
nor U2036 (N_2036,In_1530,In_2735);
nor U2037 (N_2037,In_2632,In_4371);
nand U2038 (N_2038,In_2583,In_1334);
nor U2039 (N_2039,In_2023,In_2833);
nor U2040 (N_2040,In_3415,In_2697);
and U2041 (N_2041,In_1444,In_4920);
and U2042 (N_2042,In_2323,In_846);
or U2043 (N_2043,In_509,In_2234);
and U2044 (N_2044,In_1860,In_3955);
or U2045 (N_2045,In_3109,In_2235);
or U2046 (N_2046,In_2937,In_3007);
and U2047 (N_2047,In_735,In_2730);
and U2048 (N_2048,In_1189,In_3870);
and U2049 (N_2049,In_2791,In_40);
xor U2050 (N_2050,In_129,In_3285);
nor U2051 (N_2051,In_1911,In_1705);
or U2052 (N_2052,In_563,In_1087);
xnor U2053 (N_2053,In_2922,In_1776);
or U2054 (N_2054,In_4647,In_482);
and U2055 (N_2055,In_1895,In_140);
and U2056 (N_2056,In_1616,In_4521);
nand U2057 (N_2057,In_1959,In_1889);
and U2058 (N_2058,In_2751,In_137);
and U2059 (N_2059,In_2964,In_2732);
and U2060 (N_2060,In_996,In_3565);
or U2061 (N_2061,In_1378,In_3664);
nand U2062 (N_2062,In_488,In_102);
nor U2063 (N_2063,In_2242,In_3876);
nand U2064 (N_2064,In_3030,In_1698);
and U2065 (N_2065,In_1156,In_2090);
or U2066 (N_2066,In_4940,In_868);
or U2067 (N_2067,In_3916,In_987);
nor U2068 (N_2068,In_3194,In_4063);
or U2069 (N_2069,In_3510,In_4239);
and U2070 (N_2070,In_1958,In_2594);
and U2071 (N_2071,In_3238,In_1510);
nand U2072 (N_2072,In_2335,In_2888);
and U2073 (N_2073,In_2042,In_4712);
xor U2074 (N_2074,In_3781,In_2007);
or U2075 (N_2075,In_3148,In_4260);
or U2076 (N_2076,In_2884,In_835);
xnor U2077 (N_2077,In_4266,In_4103);
xor U2078 (N_2078,In_4950,In_4031);
or U2079 (N_2079,In_4763,In_1909);
or U2080 (N_2080,In_756,In_2836);
and U2081 (N_2081,In_2247,In_1194);
nor U2082 (N_2082,In_4004,In_3372);
nor U2083 (N_2083,In_4283,In_3729);
nand U2084 (N_2084,In_4569,In_1018);
or U2085 (N_2085,In_768,In_1892);
and U2086 (N_2086,In_4526,In_2466);
nor U2087 (N_2087,In_4659,In_1596);
and U2088 (N_2088,In_4769,In_3167);
xor U2089 (N_2089,In_1817,In_2495);
or U2090 (N_2090,In_2832,In_866);
nand U2091 (N_2091,In_2045,In_4664);
nor U2092 (N_2092,In_862,In_4574);
xnor U2093 (N_2093,In_693,In_2742);
nand U2094 (N_2094,In_983,In_2299);
and U2095 (N_2095,In_1563,In_633);
or U2096 (N_2096,In_1595,In_4393);
and U2097 (N_2097,In_1272,In_2913);
or U2098 (N_2098,In_212,In_729);
or U2099 (N_2099,In_928,In_3725);
and U2100 (N_2100,In_2974,In_4081);
and U2101 (N_2101,In_1176,In_2521);
nor U2102 (N_2102,In_63,In_78);
nand U2103 (N_2103,In_1685,In_4985);
nor U2104 (N_2104,In_4800,In_2326);
or U2105 (N_2105,In_1171,In_4315);
xnor U2106 (N_2106,In_1470,In_819);
xnor U2107 (N_2107,In_4773,In_4751);
xor U2108 (N_2108,In_1461,In_961);
nand U2109 (N_2109,In_373,In_944);
nor U2110 (N_2110,In_1353,In_3863);
nand U2111 (N_2111,In_4820,In_2391);
or U2112 (N_2112,In_388,In_3726);
nor U2113 (N_2113,In_4430,In_896);
and U2114 (N_2114,In_1052,In_3373);
xnor U2115 (N_2115,In_4834,In_4279);
or U2116 (N_2116,In_4887,In_2745);
xor U2117 (N_2117,In_1929,In_3375);
and U2118 (N_2118,In_4100,In_3);
nor U2119 (N_2119,In_352,In_408);
nand U2120 (N_2120,In_3182,In_1724);
nor U2121 (N_2121,In_1094,In_1995);
xnor U2122 (N_2122,In_3756,In_1292);
xnor U2123 (N_2123,In_1404,In_3719);
and U2124 (N_2124,In_428,In_359);
xor U2125 (N_2125,In_1274,In_3513);
xnor U2126 (N_2126,In_3891,In_2659);
and U2127 (N_2127,In_780,In_360);
xnor U2128 (N_2128,In_242,In_2164);
or U2129 (N_2129,In_4332,In_3124);
xor U2130 (N_2130,In_4207,In_2249);
nand U2131 (N_2131,In_3038,In_1952);
and U2132 (N_2132,In_430,In_2719);
xnor U2133 (N_2133,In_95,In_1949);
nor U2134 (N_2134,In_111,In_2191);
or U2135 (N_2135,In_3694,In_1107);
or U2136 (N_2136,In_1532,In_3107);
nand U2137 (N_2137,In_2685,In_1694);
nand U2138 (N_2138,In_4702,In_2429);
xor U2139 (N_2139,In_2015,In_4939);
nand U2140 (N_2140,In_395,In_3265);
or U2141 (N_2141,In_1072,In_2822);
xor U2142 (N_2142,In_1922,In_4193);
nor U2143 (N_2143,In_4034,In_4427);
nand U2144 (N_2144,In_3974,In_1495);
nand U2145 (N_2145,In_2648,In_3217);
xor U2146 (N_2146,In_3027,In_3418);
and U2147 (N_2147,In_4990,In_2076);
or U2148 (N_2148,In_255,In_4195);
or U2149 (N_2149,In_3750,In_4741);
nor U2150 (N_2150,In_2831,In_2949);
nor U2151 (N_2151,In_4352,In_1964);
and U2152 (N_2152,In_177,In_386);
or U2153 (N_2153,In_1109,In_1795);
nand U2154 (N_2154,In_3646,In_3932);
nor U2155 (N_2155,In_2135,In_4963);
and U2156 (N_2156,In_4412,In_534);
or U2157 (N_2157,In_3747,In_4067);
nand U2158 (N_2158,In_4946,In_2449);
nand U2159 (N_2159,In_4451,In_722);
xnor U2160 (N_2160,In_3184,In_1992);
or U2161 (N_2161,In_2886,In_224);
xor U2162 (N_2162,In_295,In_4050);
or U2163 (N_2163,In_4594,In_4829);
and U2164 (N_2164,In_342,In_3003);
xor U2165 (N_2165,In_1878,In_1730);
xor U2166 (N_2166,In_2169,In_3055);
nand U2167 (N_2167,In_183,In_2959);
nor U2168 (N_2168,In_3049,In_2384);
nand U2169 (N_2169,In_1543,In_3056);
and U2170 (N_2170,In_2140,In_3029);
or U2171 (N_2171,In_2926,In_3524);
or U2172 (N_2172,In_876,In_2640);
or U2173 (N_2173,In_2524,In_2134);
nor U2174 (N_2174,In_4370,In_4038);
xnor U2175 (N_2175,In_2848,In_4742);
and U2176 (N_2176,In_4948,In_316);
xor U2177 (N_2177,In_4775,In_4666);
nand U2178 (N_2178,In_409,In_73);
nor U2179 (N_2179,In_2500,In_2106);
and U2180 (N_2180,In_233,In_16);
nor U2181 (N_2181,In_4649,In_311);
nand U2182 (N_2182,In_1651,In_3458);
nand U2183 (N_2183,In_4191,In_3504);
nor U2184 (N_2184,In_1278,In_2624);
or U2185 (N_2185,In_4040,In_2121);
xor U2186 (N_2186,In_2035,In_2116);
xor U2187 (N_2187,In_542,In_4580);
and U2188 (N_2188,In_1941,In_1766);
nor U2189 (N_2189,In_4916,In_497);
and U2190 (N_2190,In_1093,In_3264);
nand U2191 (N_2191,In_2971,In_2817);
nand U2192 (N_2192,In_2084,In_844);
nand U2193 (N_2193,In_4320,In_2463);
and U2194 (N_2194,In_2546,In_1347);
and U2195 (N_2195,In_3188,In_1071);
nor U2196 (N_2196,In_30,In_3428);
nor U2197 (N_2197,In_4437,In_4387);
nand U2198 (N_2198,In_2688,In_1956);
xnor U2199 (N_2199,In_3065,In_1614);
nand U2200 (N_2200,In_4653,In_2536);
or U2201 (N_2201,In_4553,In_4147);
and U2202 (N_2202,In_965,In_4377);
nor U2203 (N_2203,In_899,In_3322);
and U2204 (N_2204,In_60,In_677);
nand U2205 (N_2205,In_698,In_123);
nand U2206 (N_2206,In_580,In_4028);
xor U2207 (N_2207,In_2731,In_1477);
nor U2208 (N_2208,In_759,In_3068);
nor U2209 (N_2209,In_3302,In_1888);
nor U2210 (N_2210,In_2064,In_4479);
nand U2211 (N_2211,In_2763,In_1606);
or U2212 (N_2212,In_155,In_3195);
xor U2213 (N_2213,In_152,In_3142);
or U2214 (N_2214,In_623,In_4847);
and U2215 (N_2215,In_2706,In_4844);
nor U2216 (N_2216,In_1830,In_2695);
nor U2217 (N_2217,In_3092,In_1742);
nand U2218 (N_2218,In_3634,In_84);
and U2219 (N_2219,In_486,In_2342);
and U2220 (N_2220,In_3433,In_3011);
and U2221 (N_2221,In_384,In_757);
nand U2222 (N_2222,In_463,In_2883);
xor U2223 (N_2223,In_362,In_2083);
nand U2224 (N_2224,In_1108,In_2637);
nor U2225 (N_2225,In_399,In_3553);
and U2226 (N_2226,In_2558,In_3004);
and U2227 (N_2227,In_3773,In_2338);
xnor U2228 (N_2228,In_692,In_4956);
nand U2229 (N_2229,In_4856,In_1677);
xor U2230 (N_2230,In_2725,In_1226);
or U2231 (N_2231,In_3351,In_1573);
xor U2232 (N_2232,In_607,In_1693);
xor U2233 (N_2233,In_1775,In_3760);
nor U2234 (N_2234,In_3501,In_2729);
and U2235 (N_2235,In_4087,In_833);
or U2236 (N_2236,In_662,In_1932);
and U2237 (N_2237,In_3928,In_3585);
xor U2238 (N_2238,In_3618,In_2755);
or U2239 (N_2239,In_1140,In_1075);
nand U2240 (N_2240,In_2126,In_3703);
nor U2241 (N_2241,In_2467,In_1626);
and U2242 (N_2242,In_1333,In_2293);
and U2243 (N_2243,In_175,In_645);
nand U2244 (N_2244,In_3354,In_4674);
and U2245 (N_2245,In_4438,In_2111);
xnor U2246 (N_2246,In_1361,In_3736);
nor U2247 (N_2247,In_2593,In_1110);
nand U2248 (N_2248,In_313,In_2646);
nor U2249 (N_2249,In_2168,In_1815);
nand U2250 (N_2250,In_280,In_4487);
nand U2251 (N_2251,In_1403,In_1357);
nor U2252 (N_2252,In_41,In_3550);
xor U2253 (N_2253,In_2387,In_2386);
or U2254 (N_2254,In_2991,In_4576);
or U2255 (N_2255,In_271,In_3569);
and U2256 (N_2256,In_180,In_244);
xor U2257 (N_2257,In_107,In_3763);
xnor U2258 (N_2258,In_2180,In_4507);
nand U2259 (N_2259,In_3278,In_3012);
xnor U2260 (N_2260,In_4727,In_4423);
nand U2261 (N_2261,In_1012,In_4865);
and U2262 (N_2262,In_3843,In_2353);
nor U2263 (N_2263,In_1754,In_2332);
and U2264 (N_2264,In_187,In_4680);
and U2265 (N_2265,In_1268,In_4518);
and U2266 (N_2266,In_4853,In_2765);
or U2267 (N_2267,In_4896,In_604);
or U2268 (N_2268,In_345,In_4880);
nand U2269 (N_2269,In_3405,In_1676);
nor U2270 (N_2270,In_4730,In_3426);
nand U2271 (N_2271,In_283,In_4228);
nand U2272 (N_2272,In_1482,In_450);
or U2273 (N_2273,In_1389,In_898);
nand U2274 (N_2274,In_3939,In_4183);
nand U2275 (N_2275,In_1350,In_3384);
and U2276 (N_2276,In_875,In_4644);
nor U2277 (N_2277,In_302,In_1593);
nand U2278 (N_2278,In_3114,In_960);
xnor U2279 (N_2279,In_2823,In_1812);
and U2280 (N_2280,In_2124,In_2472);
nand U2281 (N_2281,In_3111,In_2651);
nor U2282 (N_2282,In_1998,In_3922);
xor U2283 (N_2283,In_805,In_600);
and U2284 (N_2284,In_2230,In_4555);
nand U2285 (N_2285,In_886,In_4198);
or U2286 (N_2286,In_1034,In_3269);
xnor U2287 (N_2287,In_4761,In_2530);
nand U2288 (N_2288,In_4790,In_1081);
or U2289 (N_2289,In_3320,In_3344);
nand U2290 (N_2290,In_1291,In_1399);
nor U2291 (N_2291,In_3358,In_1387);
and U2292 (N_2292,In_2141,In_4386);
or U2293 (N_2293,In_4076,In_954);
nor U2294 (N_2294,In_4077,In_864);
and U2295 (N_2295,In_713,In_4051);
or U2296 (N_2296,In_1423,In_2579);
nand U2297 (N_2297,In_1331,In_2419);
nand U2298 (N_2298,In_202,In_4154);
xor U2299 (N_2299,In_4936,In_3562);
and U2300 (N_2300,In_4850,In_1903);
nand U2301 (N_2301,In_760,In_3161);
nor U2302 (N_2302,In_3961,In_4485);
or U2303 (N_2303,In_2349,In_4958);
nand U2304 (N_2304,In_4543,In_1726);
xnor U2305 (N_2305,In_1850,In_716);
or U2306 (N_2306,In_3420,In_504);
xnor U2307 (N_2307,In_1432,In_3316);
or U2308 (N_2308,In_4355,In_4799);
nor U2309 (N_2309,In_3282,In_4204);
xnor U2310 (N_2310,In_403,In_2774);
or U2311 (N_2311,In_3878,In_4514);
or U2312 (N_2312,In_4353,In_2348);
and U2313 (N_2313,In_1729,In_2431);
xnor U2314 (N_2314,In_3658,In_4462);
nand U2315 (N_2315,In_4929,In_4826);
or U2316 (N_2316,In_3187,In_293);
or U2317 (N_2317,In_143,In_4185);
nand U2318 (N_2318,In_4692,In_2589);
and U2319 (N_2319,In_3154,In_717);
and U2320 (N_2320,In_1924,In_1457);
nor U2321 (N_2321,In_2228,In_1516);
and U2322 (N_2322,In_1701,In_3117);
and U2323 (N_2323,In_4205,In_4017);
and U2324 (N_2324,In_1249,In_3271);
and U2325 (N_2325,In_2641,In_2792);
or U2326 (N_2326,In_1774,In_3494);
xor U2327 (N_2327,In_231,In_1946);
and U2328 (N_2328,In_2486,In_2236);
nand U2329 (N_2329,In_3820,In_1800);
xnor U2330 (N_2330,In_1452,In_2563);
and U2331 (N_2331,In_3743,In_2471);
and U2332 (N_2332,In_3492,In_151);
nand U2333 (N_2333,In_1062,In_3714);
nand U2334 (N_2334,In_1231,In_1765);
nor U2335 (N_2335,In_1870,In_547);
nor U2336 (N_2336,In_2229,In_2808);
nor U2337 (N_2337,In_3752,In_2553);
nor U2338 (N_2338,In_4309,In_4750);
nor U2339 (N_2339,In_1036,In_914);
and U2340 (N_2340,In_4764,In_4599);
nand U2341 (N_2341,In_195,In_4486);
or U2342 (N_2342,In_4303,In_389);
and U2343 (N_2343,In_1615,In_2405);
nand U2344 (N_2344,In_2077,In_2941);
nor U2345 (N_2345,In_3844,In_3121);
nand U2346 (N_2346,In_1557,In_3074);
nand U2347 (N_2347,In_1764,In_861);
nand U2348 (N_2348,In_3764,In_2703);
xnor U2349 (N_2349,In_1748,In_127);
and U2350 (N_2350,In_4584,In_4152);
nor U2351 (N_2351,In_2986,In_3808);
nor U2352 (N_2352,In_4020,In_496);
or U2353 (N_2353,In_588,In_4736);
nand U2354 (N_2354,In_3978,In_118);
or U2355 (N_2355,In_4197,In_4433);
and U2356 (N_2356,In_1220,In_2838);
and U2357 (N_2357,In_2996,In_763);
nand U2358 (N_2358,In_3948,In_3544);
xnor U2359 (N_2359,In_4540,In_116);
nand U2360 (N_2360,In_417,In_1151);
xor U2361 (N_2361,In_3877,In_4689);
or U2362 (N_2362,In_4258,In_4716);
or U2363 (N_2363,In_827,In_1659);
or U2364 (N_2364,In_4348,In_1213);
nand U2365 (N_2365,In_853,In_659);
nand U2366 (N_2366,In_687,In_3622);
xor U2367 (N_2367,In_1669,In_1612);
or U2368 (N_2368,In_4200,In_2075);
xor U2369 (N_2369,In_815,In_2508);
and U2370 (N_2370,In_4502,In_4620);
or U2371 (N_2371,In_1266,In_4927);
and U2372 (N_2372,In_711,In_2717);
and U2373 (N_2373,In_1260,In_532);
xnor U2374 (N_2374,In_3176,In_1177);
nand U2375 (N_2375,In_2871,In_4415);
and U2376 (N_2376,In_2000,In_4391);
or U2377 (N_2377,In_3242,In_4235);
nand U2378 (N_2378,In_2328,In_3323);
nand U2379 (N_2379,In_951,In_2806);
nand U2380 (N_2380,In_3088,In_4341);
and U2381 (N_2381,In_4179,In_237);
and U2382 (N_2382,In_1392,In_2689);
nor U2383 (N_2383,In_2401,In_3292);
or U2384 (N_2384,In_1785,In_842);
nor U2385 (N_2385,In_2317,In_445);
and U2386 (N_2386,In_2039,In_4697);
xnor U2387 (N_2387,In_3976,In_1106);
xor U2388 (N_2388,In_685,In_745);
nor U2389 (N_2389,In_888,In_2649);
and U2390 (N_2390,In_4286,In_1682);
xnor U2391 (N_2391,In_849,In_3824);
or U2392 (N_2392,In_736,In_2209);
and U2393 (N_2393,In_4420,In_4892);
or U2394 (N_2394,In_4852,In_4728);
or U2395 (N_2395,In_932,In_2777);
and U2396 (N_2396,In_4482,In_4398);
nor U2397 (N_2397,In_4232,In_2506);
nor U2398 (N_2398,In_2853,In_571);
and U2399 (N_2399,In_491,In_3441);
and U2400 (N_2400,In_3789,In_3067);
and U2401 (N_2401,In_3066,In_228);
and U2402 (N_2402,In_4224,In_1926);
and U2403 (N_2403,In_3788,In_1983);
nand U2404 (N_2404,In_2631,In_755);
nand U2405 (N_2405,In_3526,In_2227);
xnor U2406 (N_2406,In_1577,In_1443);
nor U2407 (N_2407,In_2527,In_798);
xnor U2408 (N_2408,In_3508,In_3623);
xnor U2409 (N_2409,In_3464,In_2091);
nor U2410 (N_2410,In_353,In_3833);
and U2411 (N_2411,In_2411,In_1003);
nor U2412 (N_2412,In_1159,In_4065);
and U2413 (N_2413,In_2398,In_3132);
and U2414 (N_2414,In_109,In_1938);
or U2415 (N_2415,In_2958,In_1566);
xor U2416 (N_2416,In_2214,In_89);
and U2417 (N_2417,In_4356,In_4130);
and U2418 (N_2418,In_2354,In_3073);
xnor U2419 (N_2419,In_4695,In_101);
nor U2420 (N_2420,In_3272,In_2656);
or U2421 (N_2421,In_800,In_1753);
xnor U2422 (N_2422,In_4700,In_1471);
or U2423 (N_2423,In_1503,In_1196);
xor U2424 (N_2424,In_4796,In_1542);
xnor U2425 (N_2425,In_1029,In_2375);
and U2426 (N_2426,In_4151,In_1507);
nor U2427 (N_2427,In_1254,In_2944);
nor U2428 (N_2428,In_3774,In_3632);
and U2429 (N_2429,In_663,In_549);
nand U2430 (N_2430,In_4638,In_3885);
nand U2431 (N_2431,In_784,In_4809);
nand U2432 (N_2432,In_3307,In_2693);
nor U2433 (N_2433,In_3573,In_3153);
xor U2434 (N_2434,In_2186,In_2130);
or U2435 (N_2435,In_489,In_29);
nand U2436 (N_2436,In_1209,In_1665);
and U2437 (N_2437,In_268,In_4965);
nand U2438 (N_2438,In_1310,In_4073);
and U2439 (N_2439,In_1450,In_2307);
nand U2440 (N_2440,In_3592,In_3571);
xor U2441 (N_2441,In_1930,In_2192);
xnor U2442 (N_2442,In_897,In_4222);
or U2443 (N_2443,In_1449,In_1061);
and U2444 (N_2444,In_1456,In_3393);
nand U2445 (N_2445,In_3672,In_587);
xor U2446 (N_2446,In_2947,In_3425);
nand U2447 (N_2447,In_2782,In_4967);
nand U2448 (N_2448,In_1731,In_4140);
nand U2449 (N_2449,In_1060,In_1627);
nor U2450 (N_2450,In_803,In_3071);
and U2451 (N_2451,In_3490,In_1190);
nand U2452 (N_2452,In_4503,In_4877);
nand U2453 (N_2453,In_1007,In_2912);
nor U2454 (N_2454,In_139,In_4471);
or U2455 (N_2455,In_1492,In_4344);
or U2456 (N_2456,In_236,In_3174);
and U2457 (N_2457,In_4331,In_2248);
nand U2458 (N_2458,In_4564,In_270);
xnor U2459 (N_2459,In_3001,In_3390);
nand U2460 (N_2460,In_3546,In_339);
nor U2461 (N_2461,In_2113,In_1251);
xor U2462 (N_2462,In_3341,In_1692);
and U2463 (N_2463,In_1675,In_4508);
or U2464 (N_2464,In_2882,In_3438);
and U2465 (N_2465,In_453,In_4084);
nor U2466 (N_2466,In_23,In_1727);
nand U2467 (N_2467,In_1474,In_229);
nor U2468 (N_2468,In_2177,In_3629);
xnor U2469 (N_2469,In_4714,In_1877);
nor U2470 (N_2470,In_3901,In_2153);
nand U2471 (N_2471,In_1467,In_117);
nor U2472 (N_2472,In_2800,In_3472);
nand U2473 (N_2473,In_4548,In_4359);
or U2474 (N_2474,In_3848,In_439);
nor U2475 (N_2475,In_2301,In_2608);
nor U2476 (N_2476,In_3515,In_959);
nand U2477 (N_2477,In_4261,In_3889);
and U2478 (N_2478,In_620,In_2601);
nand U2479 (N_2479,In_2013,In_3936);
xor U2480 (N_2480,In_2903,In_435);
nor U2481 (N_2481,In_3239,In_2519);
xor U2482 (N_2482,In_14,In_2927);
and U2483 (N_2483,In_3755,In_4074);
or U2484 (N_2484,In_312,In_382);
nand U2485 (N_2485,In_3657,In_1583);
xor U2486 (N_2486,In_3563,In_2925);
xor U2487 (N_2487,In_2284,In_3468);
xor U2488 (N_2488,In_2185,In_4463);
or U2489 (N_2489,In_4275,In_407);
and U2490 (N_2490,In_1008,In_1315);
nand U2491 (N_2491,In_4048,In_3050);
or U2492 (N_2492,In_3677,In_1744);
xnor U2493 (N_2493,In_4035,In_306);
nand U2494 (N_2494,In_2003,In_3126);
nor U2495 (N_2495,In_3283,In_4805);
and U2496 (N_2496,In_4715,In_2962);
nor U2497 (N_2497,In_892,In_4719);
or U2498 (N_2498,In_3842,In_3821);
nor U2499 (N_2499,In_1097,In_3739);
nor U2500 (N_2500,N_975,N_1881);
or U2501 (N_2501,N_138,N_417);
nor U2502 (N_2502,N_2111,N_2162);
or U2503 (N_2503,N_127,N_1096);
nand U2504 (N_2504,N_140,N_2046);
xnor U2505 (N_2505,N_1295,N_1600);
and U2506 (N_2506,N_591,N_2272);
nand U2507 (N_2507,N_2038,N_1041);
xor U2508 (N_2508,N_982,N_1297);
nand U2509 (N_2509,N_1685,N_2042);
nor U2510 (N_2510,N_128,N_45);
nand U2511 (N_2511,N_154,N_1320);
xor U2512 (N_2512,N_2348,N_748);
nand U2513 (N_2513,N_1520,N_1164);
nand U2514 (N_2514,N_1779,N_174);
nor U2515 (N_2515,N_443,N_965);
xor U2516 (N_2516,N_9,N_310);
nand U2517 (N_2517,N_1968,N_96);
nand U2518 (N_2518,N_2377,N_1375);
or U2519 (N_2519,N_509,N_215);
nor U2520 (N_2520,N_2082,N_1536);
and U2521 (N_2521,N_804,N_2045);
xnor U2522 (N_2522,N_2454,N_1459);
or U2523 (N_2523,N_2357,N_1347);
xor U2524 (N_2524,N_472,N_2391);
nor U2525 (N_2525,N_2117,N_321);
nand U2526 (N_2526,N_990,N_2474);
or U2527 (N_2527,N_1400,N_1609);
or U2528 (N_2528,N_1319,N_1996);
nand U2529 (N_2529,N_419,N_882);
nor U2530 (N_2530,N_367,N_258);
nand U2531 (N_2531,N_2356,N_364);
xnor U2532 (N_2532,N_162,N_176);
xor U2533 (N_2533,N_733,N_120);
nor U2534 (N_2534,N_622,N_78);
or U2535 (N_2535,N_1538,N_1848);
or U2536 (N_2536,N_1853,N_970);
or U2537 (N_2537,N_2483,N_1445);
or U2538 (N_2538,N_165,N_1831);
and U2539 (N_2539,N_1231,N_502);
nand U2540 (N_2540,N_1140,N_813);
nand U2541 (N_2541,N_2352,N_2192);
nand U2542 (N_2542,N_1434,N_1816);
nand U2543 (N_2543,N_119,N_1932);
xnor U2544 (N_2544,N_863,N_1606);
or U2545 (N_2545,N_1194,N_1732);
xor U2546 (N_2546,N_2137,N_61);
and U2547 (N_2547,N_163,N_1200);
nand U2548 (N_2548,N_70,N_341);
nand U2549 (N_2549,N_2021,N_7);
or U2550 (N_2550,N_2437,N_1329);
nor U2551 (N_2551,N_2423,N_1248);
nor U2552 (N_2552,N_701,N_1745);
nand U2553 (N_2553,N_1723,N_1302);
and U2554 (N_2554,N_2258,N_1604);
and U2555 (N_2555,N_1170,N_424);
and U2556 (N_2556,N_683,N_831);
nand U2557 (N_2557,N_2489,N_2448);
and U2558 (N_2558,N_1877,N_2224);
nor U2559 (N_2559,N_1417,N_345);
nand U2560 (N_2560,N_1250,N_550);
and U2561 (N_2561,N_1087,N_280);
and U2562 (N_2562,N_969,N_1212);
and U2563 (N_2563,N_2132,N_1098);
xor U2564 (N_2564,N_1102,N_1909);
and U2565 (N_2565,N_1947,N_855);
nand U2566 (N_2566,N_1174,N_1285);
xor U2567 (N_2567,N_522,N_1085);
and U2568 (N_2568,N_610,N_1450);
or U2569 (N_2569,N_1707,N_770);
and U2570 (N_2570,N_1639,N_494);
and U2571 (N_2571,N_1069,N_40);
nand U2572 (N_2572,N_526,N_1624);
or U2573 (N_2573,N_749,N_2435);
nand U2574 (N_2574,N_1662,N_1316);
xnor U2575 (N_2575,N_1587,N_1072);
and U2576 (N_2576,N_482,N_2424);
nand U2577 (N_2577,N_2163,N_943);
or U2578 (N_2578,N_8,N_2265);
xor U2579 (N_2579,N_0,N_2366);
or U2580 (N_2580,N_292,N_876);
xor U2581 (N_2581,N_158,N_387);
nand U2582 (N_2582,N_1339,N_866);
xor U2583 (N_2583,N_1610,N_2482);
nor U2584 (N_2584,N_711,N_1911);
xor U2585 (N_2585,N_1119,N_1418);
xnor U2586 (N_2586,N_1941,N_1734);
or U2587 (N_2587,N_1219,N_572);
nand U2588 (N_2588,N_1974,N_884);
nor U2589 (N_2589,N_243,N_166);
nand U2590 (N_2590,N_1821,N_1872);
and U2591 (N_2591,N_218,N_976);
nand U2592 (N_2592,N_2296,N_225);
nor U2593 (N_2593,N_2317,N_621);
xnor U2594 (N_2594,N_2419,N_2169);
nor U2595 (N_2595,N_1479,N_2232);
and U2596 (N_2596,N_756,N_1120);
nor U2597 (N_2597,N_2433,N_706);
xnor U2598 (N_2598,N_1257,N_1275);
and U2599 (N_2599,N_927,N_2223);
nand U2600 (N_2600,N_2480,N_1355);
nor U2601 (N_2601,N_1991,N_2142);
xor U2602 (N_2602,N_1233,N_480);
nor U2603 (N_2603,N_1573,N_1490);
or U2604 (N_2604,N_611,N_1065);
or U2605 (N_2605,N_1081,N_267);
or U2606 (N_2606,N_2314,N_382);
nor U2607 (N_2607,N_2109,N_1819);
nand U2608 (N_2608,N_1060,N_2288);
nand U2609 (N_2609,N_1280,N_567);
nand U2610 (N_2610,N_384,N_1493);
nor U2611 (N_2611,N_1691,N_34);
xnor U2612 (N_2612,N_736,N_1213);
and U2613 (N_2613,N_1618,N_714);
xor U2614 (N_2614,N_436,N_1207);
xnor U2615 (N_2615,N_10,N_104);
nand U2616 (N_2616,N_1839,N_1919);
xor U2617 (N_2617,N_2498,N_2218);
or U2618 (N_2618,N_1886,N_1483);
and U2619 (N_2619,N_1945,N_1616);
or U2620 (N_2620,N_2191,N_281);
nand U2621 (N_2621,N_1425,N_1547);
and U2622 (N_2622,N_836,N_2175);
and U2623 (N_2623,N_2475,N_2303);
and U2624 (N_2624,N_483,N_834);
nand U2625 (N_2625,N_2097,N_726);
nand U2626 (N_2626,N_689,N_1175);
nand U2627 (N_2627,N_202,N_2075);
and U2628 (N_2628,N_327,N_2236);
xnor U2629 (N_2629,N_2100,N_1173);
nor U2630 (N_2630,N_1736,N_2384);
and U2631 (N_2631,N_213,N_217);
xor U2632 (N_2632,N_644,N_2041);
and U2633 (N_2633,N_1845,N_1124);
nand U2634 (N_2634,N_348,N_363);
and U2635 (N_2635,N_1750,N_1153);
nand U2636 (N_2636,N_852,N_1004);
nor U2637 (N_2637,N_832,N_214);
and U2638 (N_2638,N_1992,N_875);
xnor U2639 (N_2639,N_1741,N_1626);
xnor U2640 (N_2640,N_1005,N_1546);
or U2641 (N_2641,N_2245,N_2057);
nand U2642 (N_2642,N_849,N_1594);
nor U2643 (N_2643,N_2270,N_1756);
nand U2644 (N_2644,N_2309,N_2129);
xnor U2645 (N_2645,N_923,N_1057);
nor U2646 (N_2646,N_2327,N_1395);
xor U2647 (N_2647,N_942,N_1002);
nor U2648 (N_2648,N_1887,N_2016);
xnor U2649 (N_2649,N_2299,N_121);
xnor U2650 (N_2650,N_785,N_2001);
or U2651 (N_2651,N_1883,N_2294);
nand U2652 (N_2652,N_233,N_136);
nand U2653 (N_2653,N_32,N_687);
nor U2654 (N_2654,N_767,N_2182);
nand U2655 (N_2655,N_775,N_1498);
nor U2656 (N_2656,N_1680,N_222);
or U2657 (N_2657,N_940,N_1894);
and U2658 (N_2658,N_91,N_1074);
nand U2659 (N_2659,N_288,N_1560);
xnor U2660 (N_2660,N_753,N_1156);
nand U2661 (N_2661,N_1323,N_1939);
or U2662 (N_2662,N_1163,N_1201);
nor U2663 (N_2663,N_1492,N_2014);
or U2664 (N_2664,N_766,N_907);
or U2665 (N_2665,N_1984,N_113);
or U2666 (N_2666,N_1635,N_27);
nor U2667 (N_2667,N_1776,N_872);
nand U2668 (N_2668,N_1149,N_73);
xnor U2669 (N_2669,N_1976,N_80);
or U2670 (N_2670,N_894,N_1773);
xor U2671 (N_2671,N_636,N_1092);
xnor U2672 (N_2672,N_1068,N_1273);
xnor U2673 (N_2673,N_2335,N_730);
xnor U2674 (N_2674,N_577,N_1895);
nor U2675 (N_2675,N_1117,N_449);
nor U2676 (N_2676,N_1407,N_1306);
nor U2677 (N_2677,N_1660,N_1398);
xnor U2678 (N_2678,N_1551,N_1566);
xnor U2679 (N_2679,N_251,N_1046);
xnor U2680 (N_2680,N_1749,N_1182);
nand U2681 (N_2681,N_2442,N_1867);
or U2682 (N_2682,N_1012,N_2170);
nand U2683 (N_2683,N_1011,N_1211);
nor U2684 (N_2684,N_1766,N_869);
or U2685 (N_2685,N_908,N_503);
and U2686 (N_2686,N_584,N_1882);
or U2687 (N_2687,N_264,N_913);
xnor U2688 (N_2688,N_2221,N_2092);
and U2689 (N_2689,N_393,N_2273);
or U2690 (N_2690,N_905,N_2071);
nor U2691 (N_2691,N_484,N_380);
xnor U2692 (N_2692,N_1020,N_523);
nor U2693 (N_2693,N_590,N_2237);
xor U2694 (N_2694,N_2096,N_703);
or U2695 (N_2695,N_2446,N_1565);
xor U2696 (N_2696,N_1671,N_1915);
nand U2697 (N_2697,N_955,N_2225);
or U2698 (N_2698,N_111,N_2430);
nand U2699 (N_2699,N_124,N_1127);
xor U2700 (N_2700,N_1478,N_334);
nand U2701 (N_2701,N_2230,N_2362);
xnor U2702 (N_2702,N_1451,N_302);
nand U2703 (N_2703,N_499,N_1583);
nor U2704 (N_2704,N_1852,N_1424);
nand U2705 (N_2705,N_470,N_650);
or U2706 (N_2706,N_385,N_972);
nor U2707 (N_2707,N_2462,N_1725);
nand U2708 (N_2708,N_1653,N_1966);
nor U2709 (N_2709,N_1298,N_333);
and U2710 (N_2710,N_169,N_411);
and U2711 (N_2711,N_1994,N_289);
nor U2712 (N_2712,N_651,N_81);
xnor U2713 (N_2713,N_487,N_2234);
xor U2714 (N_2714,N_1561,N_476);
nand U2715 (N_2715,N_1165,N_1061);
and U2716 (N_2716,N_2381,N_230);
nor U2717 (N_2717,N_2322,N_2243);
or U2718 (N_2718,N_1258,N_248);
nand U2719 (N_2719,N_1028,N_814);
xor U2720 (N_2720,N_1722,N_453);
nand U2721 (N_2721,N_320,N_1234);
nor U2722 (N_2722,N_514,N_149);
nand U2723 (N_2723,N_1623,N_822);
or U2724 (N_2724,N_1426,N_1111);
or U2725 (N_2725,N_987,N_1761);
or U2726 (N_2726,N_642,N_1078);
or U2727 (N_2727,N_861,N_1767);
xor U2728 (N_2728,N_244,N_2018);
or U2729 (N_2729,N_2083,N_2106);
or U2730 (N_2730,N_2107,N_1603);
or U2731 (N_2731,N_2434,N_959);
nand U2732 (N_2732,N_372,N_1925);
and U2733 (N_2733,N_1777,N_1452);
nand U2734 (N_2734,N_2319,N_1688);
nand U2735 (N_2735,N_886,N_1488);
or U2736 (N_2736,N_1818,N_840);
nor U2737 (N_2737,N_747,N_724);
nand U2738 (N_2738,N_1349,N_948);
and U2739 (N_2739,N_1611,N_2378);
and U2740 (N_2740,N_84,N_1710);
or U2741 (N_2741,N_1893,N_2425);
and U2742 (N_2742,N_2473,N_440);
nand U2743 (N_2743,N_582,N_2286);
nand U2744 (N_2744,N_2471,N_1093);
xor U2745 (N_2745,N_1588,N_192);
and U2746 (N_2746,N_1249,N_631);
and U2747 (N_2747,N_918,N_2359);
nor U2748 (N_2748,N_1897,N_457);
xnor U2749 (N_2749,N_1345,N_1690);
and U2750 (N_2750,N_1539,N_356);
and U2751 (N_2751,N_1787,N_2212);
xnor U2752 (N_2752,N_729,N_2093);
and U2753 (N_2753,N_339,N_518);
or U2754 (N_2754,N_1953,N_1462);
xnor U2755 (N_2755,N_1759,N_867);
and U2756 (N_2756,N_2338,N_1921);
or U2757 (N_2757,N_294,N_2008);
or U2758 (N_2758,N_2481,N_237);
nor U2759 (N_2759,N_2090,N_1333);
or U2760 (N_2760,N_1104,N_825);
xor U2761 (N_2761,N_2054,N_2113);
and U2762 (N_2762,N_376,N_988);
nor U2763 (N_2763,N_1924,N_185);
or U2764 (N_2764,N_699,N_1376);
xor U2765 (N_2765,N_238,N_2404);
nor U2766 (N_2766,N_2479,N_1361);
or U2767 (N_2767,N_966,N_186);
or U2768 (N_2768,N_1698,N_860);
nand U2769 (N_2769,N_859,N_1913);
xor U2770 (N_2770,N_1100,N_2158);
nor U2771 (N_2771,N_938,N_425);
or U2772 (N_2772,N_1393,N_2153);
nand U2773 (N_2773,N_910,N_1849);
xor U2774 (N_2774,N_1056,N_112);
or U2775 (N_2775,N_1365,N_1557);
or U2776 (N_2776,N_1956,N_2052);
xnor U2777 (N_2777,N_359,N_1528);
nand U2778 (N_2778,N_645,N_2456);
xnor U2779 (N_2779,N_2415,N_1979);
nand U2780 (N_2780,N_576,N_407);
and U2781 (N_2781,N_2470,N_52);
xnor U2782 (N_2782,N_490,N_2233);
nor U2783 (N_2783,N_780,N_731);
or U2784 (N_2784,N_2208,N_2247);
nor U2785 (N_2785,N_458,N_2323);
nor U2786 (N_2786,N_1254,N_911);
xnor U2787 (N_2787,N_1599,N_655);
nand U2788 (N_2788,N_2028,N_608);
nor U2789 (N_2789,N_679,N_269);
or U2790 (N_2790,N_1458,N_2070);
and U2791 (N_2791,N_1563,N_613);
xnor U2792 (N_2792,N_1755,N_1131);
xnor U2793 (N_2793,N_1040,N_993);
or U2794 (N_2794,N_1703,N_612);
or U2795 (N_2795,N_1847,N_2266);
xnor U2796 (N_2796,N_1066,N_1617);
nand U2797 (N_2797,N_473,N_1044);
or U2798 (N_2798,N_2036,N_2375);
xor U2799 (N_2799,N_2458,N_578);
nand U2800 (N_2800,N_2017,N_1474);
and U2801 (N_2801,N_330,N_719);
and U2802 (N_2802,N_207,N_2280);
and U2803 (N_2803,N_2382,N_2220);
or U2804 (N_2804,N_1500,N_1770);
xor U2805 (N_2805,N_2439,N_1531);
and U2806 (N_2806,N_1857,N_601);
or U2807 (N_2807,N_551,N_1942);
and U2808 (N_2808,N_581,N_681);
nor U2809 (N_2809,N_1412,N_2134);
xor U2810 (N_2810,N_62,N_426);
nor U2811 (N_2811,N_293,N_542);
nand U2812 (N_2812,N_141,N_2124);
nor U2813 (N_2813,N_1022,N_718);
or U2814 (N_2814,N_1471,N_2277);
and U2815 (N_2815,N_2497,N_2308);
xor U2816 (N_2816,N_257,N_125);
xnor U2817 (N_2817,N_772,N_2254);
nor U2818 (N_2818,N_558,N_28);
or U2819 (N_2819,N_231,N_2049);
nand U2820 (N_2820,N_447,N_998);
or U2821 (N_2821,N_1134,N_2328);
xnor U2822 (N_2822,N_1649,N_506);
nor U2823 (N_2823,N_160,N_1289);
nor U2824 (N_2824,N_2339,N_598);
nor U2825 (N_2825,N_802,N_1514);
nor U2826 (N_2826,N_1681,N_1346);
xnor U2827 (N_2827,N_618,N_2);
nand U2828 (N_2828,N_463,N_105);
nor U2829 (N_2829,N_2281,N_919);
nor U2830 (N_2830,N_2401,N_1372);
xnor U2831 (N_2831,N_1267,N_568);
xor U2832 (N_2832,N_707,N_2494);
nor U2833 (N_2833,N_830,N_984);
nor U2834 (N_2834,N_1875,N_1358);
nand U2835 (N_2835,N_1252,N_2108);
nand U2836 (N_2836,N_455,N_2073);
and U2837 (N_2837,N_2403,N_2340);
xnor U2838 (N_2838,N_2298,N_228);
or U2839 (N_2839,N_2098,N_1775);
or U2840 (N_2840,N_1047,N_1186);
xor U2841 (N_2841,N_805,N_1666);
nand U2842 (N_2842,N_1842,N_530);
nand U2843 (N_2843,N_2069,N_155);
or U2844 (N_2844,N_930,N_15);
or U2845 (N_2845,N_1754,N_1896);
nand U2846 (N_2846,N_389,N_1378);
nand U2847 (N_2847,N_1993,N_1862);
and U2848 (N_2848,N_1366,N_1215);
nand U2849 (N_2849,N_603,N_263);
nor U2850 (N_2850,N_2274,N_759);
xnor U2851 (N_2851,N_2094,N_381);
or U2852 (N_2852,N_1543,N_2418);
and U2853 (N_2853,N_761,N_2346);
nor U2854 (N_2854,N_2056,N_543);
xor U2855 (N_2855,N_1652,N_1287);
nor U2856 (N_2856,N_254,N_1657);
and U2857 (N_2857,N_2155,N_971);
nor U2858 (N_2858,N_1542,N_1608);
or U2859 (N_2859,N_1322,N_2431);
nor U2860 (N_2860,N_74,N_1946);
or U2861 (N_2861,N_1310,N_1097);
or U2862 (N_2862,N_1385,N_1261);
nand U2863 (N_2863,N_856,N_88);
or U2864 (N_2864,N_991,N_2461);
nand U2865 (N_2865,N_688,N_1985);
nand U2866 (N_2866,N_200,N_673);
and U2867 (N_2867,N_1453,N_891);
or U2868 (N_2868,N_1957,N_1391);
or U2869 (N_2869,N_229,N_1383);
nand U2870 (N_2870,N_1502,N_939);
and U2871 (N_2871,N_954,N_1381);
nand U2872 (N_2872,N_615,N_838);
nor U2873 (N_2873,N_1260,N_1283);
xnor U2874 (N_2874,N_783,N_896);
nand U2875 (N_2875,N_839,N_1961);
or U2876 (N_2876,N_1171,N_343);
nand U2877 (N_2877,N_1150,N_1769);
and U2878 (N_2878,N_843,N_2361);
xor U2879 (N_2879,N_515,N_2445);
xnor U2880 (N_2880,N_1006,N_501);
xnor U2881 (N_2881,N_2157,N_274);
xor U2882 (N_2882,N_2229,N_1571);
nand U2883 (N_2883,N_1147,N_1643);
xor U2884 (N_2884,N_1314,N_2079);
or U2885 (N_2885,N_452,N_709);
and U2886 (N_2886,N_143,N_1650);
or U2887 (N_2887,N_2257,N_2388);
or U2888 (N_2888,N_1826,N_2005);
nand U2889 (N_2889,N_1362,N_1299);
nor U2890 (N_2890,N_1679,N_2118);
xnor U2891 (N_2891,N_1811,N_2064);
or U2892 (N_2892,N_2013,N_774);
and U2893 (N_2893,N_890,N_1912);
xor U2894 (N_2894,N_1512,N_68);
nor U2895 (N_2895,N_1113,N_1324);
nor U2896 (N_2896,N_1486,N_2161);
xnor U2897 (N_2897,N_67,N_2179);
nand U2898 (N_2898,N_1332,N_1602);
nand U2899 (N_2899,N_2360,N_466);
xor U2900 (N_2900,N_732,N_2149);
nor U2901 (N_2901,N_817,N_549);
and U2902 (N_2902,N_720,N_1160);
and U2903 (N_2903,N_1700,N_2397);
or U2904 (N_2904,N_1654,N_2174);
or U2905 (N_2905,N_196,N_782);
xor U2906 (N_2906,N_1589,N_801);
xor U2907 (N_2907,N_1335,N_2414);
nand U2908 (N_2908,N_2402,N_725);
and U2909 (N_2909,N_1555,N_22);
or U2910 (N_2910,N_56,N_1664);
nand U2911 (N_2911,N_31,N_1612);
or U2912 (N_2912,N_170,N_2066);
xor U2913 (N_2913,N_556,N_1367);
nor U2914 (N_2914,N_989,N_1276);
or U2915 (N_2915,N_677,N_1930);
and U2916 (N_2916,N_1701,N_1438);
and U2917 (N_2917,N_1139,N_30);
and U2918 (N_2918,N_2264,N_1264);
and U2919 (N_2919,N_1711,N_2405);
nand U2920 (N_2920,N_1846,N_1647);
nor U2921 (N_2921,N_546,N_1136);
and U2922 (N_2922,N_134,N_1964);
or U2923 (N_2923,N_1824,N_1972);
nor U2924 (N_2924,N_325,N_445);
xnor U2925 (N_2925,N_2329,N_1308);
and U2926 (N_2926,N_1429,N_1533);
and U2927 (N_2927,N_1112,N_531);
xor U2928 (N_2928,N_692,N_1431);
and U2929 (N_2929,N_131,N_1670);
or U2930 (N_2930,N_171,N_2496);
xor U2931 (N_2931,N_456,N_794);
or U2932 (N_2932,N_818,N_1288);
and U2933 (N_2933,N_935,N_408);
and U2934 (N_2934,N_401,N_1661);
or U2935 (N_2935,N_1581,N_1771);
xnor U2936 (N_2936,N_997,N_1075);
nand U2937 (N_2937,N_1633,N_1035);
nor U2938 (N_2938,N_854,N_754);
or U2939 (N_2939,N_630,N_1789);
xor U2940 (N_2940,N_791,N_106);
nand U2941 (N_2941,N_1387,N_423);
nand U2942 (N_2942,N_620,N_1989);
xor U2943 (N_2943,N_2389,N_1336);
nor U2944 (N_2944,N_1592,N_1807);
xnor U2945 (N_2945,N_1045,N_1427);
xor U2946 (N_2946,N_1224,N_1523);
nor U2947 (N_2947,N_602,N_1491);
xor U2948 (N_2948,N_619,N_398);
nor U2949 (N_2949,N_2127,N_696);
nand U2950 (N_2950,N_42,N_2457);
nor U2951 (N_2951,N_628,N_1313);
nand U2952 (N_2952,N_2203,N_102);
xnor U2953 (N_2953,N_893,N_1586);
and U2954 (N_2954,N_1621,N_824);
and U2955 (N_2955,N_1879,N_2026);
nand U2956 (N_2956,N_432,N_1595);
nand U2957 (N_2957,N_1937,N_781);
or U2958 (N_2958,N_539,N_1860);
and U2959 (N_2959,N_369,N_307);
and U2960 (N_2960,N_2289,N_1294);
nand U2961 (N_2961,N_1572,N_1018);
nor U2962 (N_2962,N_776,N_864);
nand U2963 (N_2963,N_1067,N_1795);
nor U2964 (N_2964,N_1436,N_1803);
nor U2965 (N_2965,N_2067,N_1206);
and U2966 (N_2966,N_1596,N_1827);
nand U2967 (N_2967,N_1190,N_2350);
and U2968 (N_2968,N_261,N_206);
nor U2969 (N_2969,N_1977,N_1428);
and U2970 (N_2970,N_800,N_798);
xor U2971 (N_2971,N_1851,N_752);
and U2972 (N_2972,N_2209,N_159);
nor U2973 (N_2973,N_2334,N_633);
and U2974 (N_2974,N_1683,N_246);
xor U2975 (N_2975,N_1435,N_1556);
nor U2976 (N_2976,N_1138,N_1644);
and U2977 (N_2977,N_1526,N_2312);
nand U2978 (N_2978,N_1246,N_1185);
and U2979 (N_2979,N_1238,N_1752);
or U2980 (N_2980,N_1548,N_1494);
xnor U2981 (N_2981,N_1402,N_1751);
or U2982 (N_2982,N_72,N_1334);
and U2983 (N_2983,N_1341,N_1290);
and U2984 (N_2984,N_528,N_547);
xnor U2985 (N_2985,N_285,N_268);
or U2986 (N_2986,N_2128,N_1155);
or U2987 (N_2987,N_637,N_184);
xnor U2988 (N_2988,N_2032,N_2386);
and U2989 (N_2989,N_1278,N_1304);
xor U2990 (N_2990,N_1553,N_2040);
and U2991 (N_2991,N_2279,N_2358);
xor U2992 (N_2992,N_773,N_2320);
and U2993 (N_2993,N_2251,N_1419);
nand U2994 (N_2994,N_573,N_1950);
nand U2995 (N_2995,N_495,N_765);
nor U2996 (N_2996,N_1615,N_1199);
nor U2997 (N_2997,N_2148,N_906);
xnor U2998 (N_2998,N_1579,N_1676);
or U2999 (N_2999,N_1321,N_1177);
or U3000 (N_3000,N_871,N_107);
nor U3001 (N_3001,N_1986,N_2226);
nor U3002 (N_3002,N_1110,N_1439);
or U3003 (N_3003,N_2197,N_2326);
and U3004 (N_3004,N_589,N_1148);
or U3005 (N_3005,N_1796,N_1469);
xor U3006 (N_3006,N_668,N_1030);
xor U3007 (N_3007,N_1808,N_132);
and U3008 (N_3008,N_2499,N_89);
nor U3009 (N_3009,N_750,N_375);
nand U3010 (N_3010,N_2189,N_1399);
or U3011 (N_3011,N_1527,N_1051);
nand U3012 (N_3012,N_533,N_337);
nand U3013 (N_3013,N_1195,N_212);
or U3014 (N_3014,N_1187,N_2333);
or U3015 (N_3015,N_835,N_953);
and U3016 (N_3016,N_1782,N_715);
or U3017 (N_3017,N_1145,N_1935);
and U3018 (N_3018,N_2409,N_1386);
nand U3019 (N_3019,N_2105,N_1437);
and U3020 (N_3020,N_2330,N_1303);
and U3021 (N_3021,N_1226,N_2144);
or U3022 (N_3022,N_21,N_242);
or U3023 (N_3023,N_771,N_516);
nor U3024 (N_3024,N_232,N_3);
and U3025 (N_3025,N_1674,N_1516);
nand U3026 (N_3026,N_1634,N_2305);
and U3027 (N_3027,N_2488,N_1888);
nand U3028 (N_3028,N_1368,N_964);
nor U3029 (N_3029,N_2476,N_461);
nor U3030 (N_3030,N_1900,N_521);
nor U3031 (N_3031,N_978,N_1449);
or U3032 (N_3032,N_1379,N_1064);
and U3033 (N_3033,N_680,N_513);
or U3034 (N_3034,N_710,N_20);
nor U3035 (N_3035,N_1940,N_2487);
xor U3036 (N_3036,N_2394,N_2491);
nor U3037 (N_3037,N_979,N_1099);
xnor U3038 (N_3038,N_299,N_221);
or U3039 (N_3039,N_2302,N_76);
and U3040 (N_3040,N_1850,N_2428);
nand U3041 (N_3041,N_1286,N_2369);
or U3042 (N_3042,N_712,N_471);
nor U3043 (N_3043,N_133,N_1830);
nor U3044 (N_3044,N_1675,N_156);
xnor U3045 (N_3045,N_566,N_2166);
nand U3046 (N_3046,N_2353,N_1158);
nor U3047 (N_3047,N_442,N_2269);
nor U3048 (N_3048,N_2387,N_1441);
nand U3049 (N_3049,N_2207,N_451);
or U3050 (N_3050,N_1476,N_427);
nor U3051 (N_3051,N_181,N_2168);
and U3052 (N_3052,N_239,N_1269);
and U3053 (N_3053,N_535,N_788);
or U3054 (N_3054,N_779,N_1638);
nand U3055 (N_3055,N_63,N_757);
xnor U3056 (N_3056,N_1082,N_2199);
nor U3057 (N_3057,N_234,N_904);
nor U3058 (N_3058,N_1109,N_319);
nor U3059 (N_3059,N_1374,N_352);
or U3060 (N_3060,N_2164,N_1318);
nand U3061 (N_3061,N_1454,N_139);
xor U3062 (N_3062,N_335,N_983);
nand U3063 (N_3063,N_745,N_328);
and U3064 (N_3064,N_879,N_371);
xor U3065 (N_3065,N_1487,N_175);
nor U3066 (N_3066,N_2061,N_2325);
xor U3067 (N_3067,N_899,N_1470);
or U3068 (N_3068,N_926,N_1704);
and U3069 (N_3069,N_2410,N_1157);
and U3070 (N_3070,N_604,N_2407);
nor U3071 (N_3071,N_1590,N_1241);
and U3072 (N_3072,N_198,N_777);
nor U3073 (N_3073,N_1562,N_313);
nor U3074 (N_3074,N_2154,N_1780);
or U3075 (N_3075,N_1468,N_2146);
xor U3076 (N_3076,N_1636,N_842);
or U3077 (N_3077,N_342,N_2084);
or U3078 (N_3078,N_740,N_588);
xnor U3079 (N_3079,N_925,N_815);
or U3080 (N_3080,N_2053,N_1672);
nand U3081 (N_3081,N_2160,N_2114);
xnor U3082 (N_3082,N_101,N_1705);
nand U3083 (N_3083,N_1584,N_2116);
xor U3084 (N_3084,N_1015,N_837);
or U3085 (N_3085,N_1637,N_362);
and U3086 (N_3086,N_974,N_297);
or U3087 (N_3087,N_86,N_1049);
xor U3088 (N_3088,N_1737,N_826);
nand U3089 (N_3089,N_1694,N_1354);
or U3090 (N_3090,N_540,N_1960);
nor U3091 (N_3091,N_1377,N_2395);
nor U3092 (N_3092,N_1834,N_2227);
nand U3093 (N_3093,N_1760,N_2466);
nor U3094 (N_3094,N_2121,N_653);
and U3095 (N_3095,N_1938,N_309);
nor U3096 (N_3096,N_1166,N_1086);
nor U3097 (N_3097,N_1235,N_474);
or U3098 (N_3098,N_318,N_981);
nor U3099 (N_3099,N_1414,N_1965);
xnor U3100 (N_3100,N_1646,N_1326);
and U3101 (N_3101,N_931,N_178);
or U3102 (N_3102,N_2188,N_585);
xor U3103 (N_3103,N_145,N_646);
xnor U3104 (N_3104,N_1861,N_1292);
nor U3105 (N_3105,N_1916,N_2091);
and U3106 (N_3106,N_1980,N_1076);
nand U3107 (N_3107,N_2123,N_881);
nand U3108 (N_3108,N_2492,N_354);
or U3109 (N_3109,N_2235,N_1227);
nor U3110 (N_3110,N_1184,N_901);
xor U3111 (N_3111,N_1029,N_399);
nor U3112 (N_3112,N_403,N_760);
xnor U3113 (N_3113,N_147,N_643);
nor U3114 (N_3114,N_19,N_1343);
nand U3115 (N_3115,N_1863,N_137);
nand U3116 (N_3116,N_66,N_1340);
or U3117 (N_3117,N_557,N_368);
nor U3118 (N_3118,N_1790,N_1693);
xor U3119 (N_3119,N_662,N_2316);
nor U3120 (N_3120,N_1016,N_898);
and U3121 (N_3121,N_126,N_378);
nand U3122 (N_3122,N_397,N_167);
and U3123 (N_3123,N_190,N_2332);
nor U3124 (N_3124,N_928,N_350);
nor U3125 (N_3125,N_1669,N_1578);
and U3126 (N_3126,N_1866,N_405);
xor U3127 (N_3127,N_301,N_2048);
xor U3128 (N_3128,N_1765,N_1038);
xnor U3129 (N_3129,N_336,N_1176);
and U3130 (N_3130,N_168,N_1088);
nor U3131 (N_3131,N_1597,N_1331);
xor U3132 (N_3132,N_527,N_1856);
nor U3133 (N_3133,N_6,N_2125);
nor U3134 (N_3134,N_435,N_1764);
xor U3135 (N_3135,N_60,N_1037);
nand U3136 (N_3136,N_1161,N_1183);
nand U3137 (N_3137,N_2020,N_1209);
xor U3138 (N_3138,N_1116,N_262);
nand U3139 (N_3139,N_1892,N_1396);
and U3140 (N_3140,N_400,N_2283);
nand U3141 (N_3141,N_2263,N_694);
or U3142 (N_3142,N_59,N_2301);
or U3143 (N_3143,N_520,N_2469);
xor U3144 (N_3144,N_12,N_2460);
and U3145 (N_3145,N_1810,N_497);
nand U3146 (N_3146,N_324,N_827);
or U3147 (N_3147,N_315,N_1641);
nor U3148 (N_3148,N_1828,N_37);
xor U3149 (N_3149,N_900,N_272);
nor U3150 (N_3150,N_271,N_208);
xor U3151 (N_3151,N_1351,N_669);
or U3152 (N_3152,N_2313,N_1048);
nand U3153 (N_3153,N_2441,N_2307);
nor U3154 (N_3154,N_493,N_347);
and U3155 (N_3155,N_2341,N_1009);
or U3156 (N_3156,N_188,N_986);
or U3157 (N_3157,N_1836,N_402);
nand U3158 (N_3158,N_2248,N_564);
and U3159 (N_3159,N_2304,N_789);
nor U3160 (N_3160,N_996,N_1655);
nor U3161 (N_3161,N_2310,N_1103);
nor U3162 (N_3162,N_1651,N_199);
nor U3163 (N_3163,N_2171,N_1282);
xnor U3164 (N_3164,N_2165,N_1480);
or U3165 (N_3165,N_75,N_1899);
and U3166 (N_3166,N_583,N_2374);
and U3167 (N_3167,N_2138,N_5);
nand U3168 (N_3168,N_459,N_1914);
and U3169 (N_3169,N_2440,N_691);
nand U3170 (N_3170,N_1050,N_1495);
and U3171 (N_3171,N_100,N_2331);
and U3172 (N_3172,N_1141,N_2450);
nand U3173 (N_3173,N_656,N_1854);
and U3174 (N_3174,N_1389,N_1699);
xnor U3175 (N_3175,N_360,N_58);
xor U3176 (N_3176,N_575,N_1840);
and U3177 (N_3177,N_1309,N_2249);
and U3178 (N_3178,N_1822,N_211);
nand U3179 (N_3179,N_1239,N_1317);
or U3180 (N_3180,N_441,N_1815);
xnor U3181 (N_3181,N_1545,N_977);
xnor U3182 (N_3182,N_1798,N_2072);
nor U3183 (N_3183,N_2285,N_1410);
or U3184 (N_3184,N_2337,N_1151);
and U3185 (N_3185,N_2259,N_1746);
nor U3186 (N_3186,N_2453,N_2034);
and U3187 (N_3187,N_1763,N_1733);
nor U3188 (N_3188,N_2250,N_665);
nand U3189 (N_3189,N_1902,N_592);
xor U3190 (N_3190,N_429,N_1665);
nand U3191 (N_3191,N_2495,N_1159);
and U3192 (N_3192,N_2242,N_108);
or U3193 (N_3193,N_2010,N_90);
nand U3194 (N_3194,N_2416,N_1507);
or U3195 (N_3195,N_179,N_2029);
nor U3196 (N_3196,N_83,N_967);
and U3197 (N_3197,N_2467,N_1905);
nor U3198 (N_3198,N_2422,N_1511);
and U3199 (N_3199,N_2076,N_1791);
and U3200 (N_3200,N_1397,N_305);
nand U3201 (N_3201,N_2412,N_1146);
xor U3202 (N_3202,N_2324,N_1457);
and U3203 (N_3203,N_880,N_465);
nor U3204 (N_3204,N_647,N_1687);
and U3205 (N_3205,N_625,N_962);
xor U3206 (N_3206,N_1373,N_1864);
nor U3207 (N_3207,N_478,N_1251);
or U3208 (N_3208,N_428,N_444);
nand U3209 (N_3209,N_1277,N_916);
nand U3210 (N_3210,N_1835,N_2194);
nand U3211 (N_3211,N_2214,N_2241);
and U3212 (N_3212,N_877,N_1091);
or U3213 (N_3213,N_635,N_1605);
nand U3214 (N_3214,N_1792,N_1788);
nand U3215 (N_3215,N_2126,N_422);
nor U3216 (N_3216,N_1668,N_1812);
xor U3217 (N_3217,N_1095,N_999);
nand U3218 (N_3218,N_148,N_1001);
nand U3219 (N_3219,N_1833,N_410);
xor U3220 (N_3220,N_1577,N_1744);
and U3221 (N_3221,N_1422,N_1645);
or U3222 (N_3222,N_902,N_1325);
and U3223 (N_3223,N_2147,N_2287);
xor U3224 (N_3224,N_1353,N_2295);
nor U3225 (N_3225,N_609,N_157);
nand U3226 (N_3226,N_1013,N_41);
xnor U3227 (N_3227,N_300,N_1223);
and U3228 (N_3228,N_500,N_1077);
xor U3229 (N_3229,N_1420,N_1216);
or U3230 (N_3230,N_1245,N_1000);
nand U3231 (N_3231,N_1014,N_658);
nor U3232 (N_3232,N_1799,N_1401);
or U3233 (N_3233,N_182,N_1983);
nand U3234 (N_3234,N_1179,N_460);
and U3235 (N_3235,N_475,N_2451);
and U3236 (N_3236,N_796,N_587);
nor U3237 (N_3237,N_862,N_2390);
or U3238 (N_3238,N_1010,N_1205);
or U3239 (N_3239,N_1301,N_742);
nand U3240 (N_3240,N_2399,N_713);
xnor U3241 (N_3241,N_1043,N_1217);
or U3242 (N_3242,N_561,N_1181);
and U3243 (N_3243,N_690,N_49);
nand U3244 (N_3244,N_404,N_1126);
nor U3245 (N_3245,N_878,N_183);
and U3246 (N_3246,N_1342,N_738);
xnor U3247 (N_3247,N_1684,N_1293);
nor U3248 (N_3248,N_2152,N_1025);
nor U3249 (N_3249,N_722,N_2426);
xnor U3250 (N_3250,N_2315,N_331);
nand U3251 (N_3251,N_973,N_394);
nand U3252 (N_3252,N_1430,N_2490);
xor U3253 (N_3253,N_379,N_1715);
xor U3254 (N_3254,N_786,N_1786);
and U3255 (N_3255,N_1975,N_1959);
and U3256 (N_3256,N_614,N_2215);
or U3257 (N_3257,N_1948,N_1390);
and U3258 (N_3258,N_489,N_1598);
xor U3259 (N_3259,N_933,N_648);
and U3260 (N_3260,N_79,N_704);
xor U3261 (N_3261,N_1007,N_1003);
nand U3262 (N_3262,N_1501,N_117);
nor U3263 (N_3263,N_605,N_2449);
nor U3264 (N_3264,N_1525,N_1804);
xnor U3265 (N_3265,N_555,N_968);
and U3266 (N_3266,N_1797,N_1884);
nand U3267 (N_3267,N_252,N_1460);
xnor U3268 (N_3268,N_2078,N_2177);
and U3269 (N_3269,N_1415,N_2200);
xor U3270 (N_3270,N_1874,N_194);
xor U3271 (N_3271,N_1640,N_283);
or U3272 (N_3272,N_223,N_1969);
nand U3273 (N_3273,N_1878,N_1591);
nor U3274 (N_3274,N_2193,N_2421);
nor U3275 (N_3275,N_1918,N_2088);
nor U3276 (N_3276,N_340,N_1981);
or U3277 (N_3277,N_1255,N_1394);
xnor U3278 (N_3278,N_858,N_275);
or U3279 (N_3279,N_308,N_2371);
nor U3280 (N_3280,N_439,N_2022);
or U3281 (N_3281,N_1567,N_180);
nand U3282 (N_3282,N_1307,N_1967);
nor U3283 (N_3283,N_1482,N_1642);
nand U3284 (N_3284,N_723,N_1094);
nand U3285 (N_3285,N_1237,N_1291);
nand U3286 (N_3286,N_995,N_1413);
nand U3287 (N_3287,N_946,N_548);
nor U3288 (N_3288,N_1729,N_1716);
and U3289 (N_3289,N_1554,N_1885);
xor U3290 (N_3290,N_1444,N_1720);
nand U3291 (N_3291,N_1026,N_173);
nor U3292 (N_3292,N_1743,N_746);
xor U3293 (N_3293,N_421,N_1873);
nor U3294 (N_3294,N_201,N_1122);
or U3295 (N_3295,N_85,N_702);
or U3296 (N_3296,N_1510,N_1409);
xor U3297 (N_3297,N_2363,N_563);
xor U3298 (N_3298,N_1380,N_1955);
and U3299 (N_3299,N_1820,N_847);
nand U3300 (N_3300,N_1363,N_1135);
and U3301 (N_3301,N_1312,N_1625);
or U3302 (N_3302,N_153,N_596);
and U3303 (N_3303,N_1727,N_2143);
nor U3304 (N_3304,N_2455,N_1107);
nand U3305 (N_3305,N_1263,N_629);
nor U3306 (N_3306,N_1541,N_2024);
nand U3307 (N_3307,N_565,N_1017);
and U3308 (N_3308,N_1575,N_1504);
nand U3309 (N_3309,N_2432,N_291);
and U3310 (N_3310,N_390,N_2062);
or U3311 (N_3311,N_1825,N_1403);
nand U3312 (N_3312,N_828,N_2354);
nand U3313 (N_3313,N_1466,N_2074);
or U3314 (N_3314,N_358,N_2336);
and U3315 (N_3315,N_235,N_841);
nor U3316 (N_3316,N_197,N_505);
and U3317 (N_3317,N_737,N_1889);
and U3318 (N_3318,N_769,N_1034);
nand U3319 (N_3319,N_249,N_351);
nor U3320 (N_3320,N_1574,N_365);
or U3321 (N_3321,N_1713,N_1128);
and U3322 (N_3322,N_820,N_1118);
nand U3323 (N_3323,N_57,N_25);
and U3324 (N_3324,N_2342,N_758);
nor U3325 (N_3325,N_388,N_1496);
nand U3326 (N_3326,N_64,N_2130);
nor U3327 (N_3327,N_1330,N_1130);
nor U3328 (N_3328,N_1806,N_2183);
nor U3329 (N_3329,N_386,N_663);
xnor U3330 (N_3330,N_193,N_961);
xnor U3331 (N_3331,N_1198,N_1106);
nor U3332 (N_3332,N_914,N_329);
and U3333 (N_3333,N_97,N_510);
and U3334 (N_3334,N_55,N_1033);
nor U3335 (N_3335,N_311,N_741);
and U3336 (N_3336,N_1689,N_2477);
or U3337 (N_3337,N_344,N_17);
nor U3338 (N_3338,N_1300,N_129);
nand U3339 (N_3339,N_1696,N_1712);
nor U3340 (N_3340,N_1464,N_1270);
and U3341 (N_3341,N_1582,N_1485);
or U3342 (N_3342,N_332,N_468);
xnor U3343 (N_3343,N_287,N_1951);
nor U3344 (N_3344,N_672,N_2068);
nor U3345 (N_3345,N_298,N_897);
or U3346 (N_3346,N_488,N_1535);
or U3347 (N_3347,N_103,N_2140);
nor U3348 (N_3348,N_1929,N_1503);
or U3349 (N_3349,N_418,N_161);
and U3350 (N_3350,N_883,N_2459);
and U3351 (N_3351,N_109,N_36);
xnor U3352 (N_3352,N_498,N_537);
nor U3353 (N_3353,N_1607,N_2246);
nand U3354 (N_3354,N_616,N_2290);
nor U3355 (N_3355,N_1073,N_282);
or U3356 (N_3356,N_1230,N_851);
nand U3357 (N_3357,N_2478,N_2211);
or U3358 (N_3358,N_1188,N_1506);
nor U3359 (N_3359,N_496,N_1721);
xnor U3360 (N_3360,N_2131,N_2278);
nand U3361 (N_3361,N_1404,N_2447);
nor U3362 (N_3362,N_728,N_2260);
and U3363 (N_3363,N_1923,N_1858);
and U3364 (N_3364,N_2300,N_627);
nand U3365 (N_3365,N_77,N_695);
xnor U3366 (N_3366,N_952,N_1279);
xor U3367 (N_3367,N_1677,N_716);
or U3368 (N_3368,N_922,N_2035);
xor U3369 (N_3369,N_570,N_1123);
nand U3370 (N_3370,N_600,N_2345);
and U3371 (N_3371,N_1521,N_889);
xnor U3372 (N_3372,N_2376,N_903);
or U3373 (N_3373,N_1143,N_915);
nand U3374 (N_3374,N_1042,N_2030);
and U3375 (N_3375,N_227,N_1225);
xor U3376 (N_3376,N_1742,N_700);
nand U3377 (N_3377,N_357,N_1021);
or U3378 (N_3378,N_317,N_1898);
and U3379 (N_3379,N_1229,N_1125);
xnor U3380 (N_3380,N_626,N_203);
nand U3381 (N_3381,N_1580,N_2102);
nand U3382 (N_3382,N_2039,N_1728);
nor U3383 (N_3383,N_654,N_1196);
or U3384 (N_3384,N_912,N_396);
or U3385 (N_3385,N_1062,N_1534);
and U3386 (N_3386,N_1876,N_1296);
or U3387 (N_3387,N_1191,N_2196);
nor U3388 (N_3388,N_434,N_1739);
nor U3389 (N_3389,N_956,N_2408);
and U3390 (N_3390,N_1197,N_929);
xnor U3391 (N_3391,N_2493,N_1865);
and U3392 (N_3392,N_579,N_623);
nand U3393 (N_3393,N_2438,N_1774);
xor U3394 (N_3394,N_2139,N_829);
or U3395 (N_3395,N_797,N_2240);
nor U3396 (N_3396,N_1059,N_477);
and U3397 (N_3397,N_763,N_152);
xnor U3398 (N_3398,N_1659,N_553);
nor U3399 (N_3399,N_1686,N_2178);
xor U3400 (N_3400,N_338,N_1019);
and U3401 (N_3401,N_792,N_638);
nand U3402 (N_3402,N_1958,N_1802);
nor U3403 (N_3403,N_808,N_2156);
xor U3404 (N_3404,N_1540,N_1927);
nor U3405 (N_3405,N_209,N_1524);
and U3406 (N_3406,N_2222,N_224);
nor U3407 (N_3407,N_682,N_676);
nor U3408 (N_3408,N_247,N_135);
and U3409 (N_3409,N_1813,N_1505);
nand U3410 (N_3410,N_1058,N_743);
and U3411 (N_3411,N_1443,N_1998);
nand U3412 (N_3412,N_2112,N_1658);
nor U3413 (N_3413,N_1917,N_1663);
nand U3414 (N_3414,N_467,N_1692);
nor U3415 (N_3415,N_69,N_35);
xor U3416 (N_3416,N_1382,N_204);
nor U3417 (N_3417,N_2231,N_2012);
and U3418 (N_3418,N_481,N_1601);
nand U3419 (N_3419,N_1180,N_2472);
nor U3420 (N_3420,N_1406,N_1359);
nor U3421 (N_3421,N_414,N_960);
or U3422 (N_3422,N_684,N_941);
or U3423 (N_3423,N_95,N_1071);
or U3424 (N_3424,N_253,N_2050);
xnor U3425 (N_3425,N_433,N_1169);
xor U3426 (N_3426,N_1456,N_2198);
xor U3427 (N_3427,N_1132,N_1027);
nand U3428 (N_3428,N_1971,N_306);
and U3429 (N_3429,N_374,N_833);
nand U3430 (N_3430,N_1922,N_1718);
nand U3431 (N_3431,N_150,N_1311);
and U3432 (N_3432,N_220,N_1259);
nand U3433 (N_3433,N_674,N_2318);
xnor U3434 (N_3434,N_4,N_1628);
xnor U3435 (N_3435,N_1455,N_1805);
nor U3436 (N_3436,N_795,N_580);
nand U3437 (N_3437,N_1477,N_1228);
or U3438 (N_3438,N_1284,N_151);
and U3439 (N_3439,N_1433,N_529);
nand U3440 (N_3440,N_296,N_2120);
xor U3441 (N_3441,N_1868,N_2023);
nand U3442 (N_3442,N_819,N_2297);
or U3443 (N_3443,N_349,N_1108);
or U3444 (N_3444,N_1768,N_1202);
or U3445 (N_3445,N_1222,N_784);
nor U3446 (N_3446,N_2306,N_2239);
or U3447 (N_3447,N_1272,N_2238);
nor U3448 (N_3448,N_2003,N_2037);
nand U3449 (N_3449,N_1357,N_118);
nand U3450 (N_3450,N_2081,N_1890);
or U3451 (N_3451,N_2406,N_2452);
xor U3452 (N_3452,N_874,N_391);
nand U3453 (N_3453,N_2006,N_803);
nand U3454 (N_3454,N_1735,N_312);
nor U3455 (N_3455,N_1844,N_1133);
nand U3456 (N_3456,N_1593,N_853);
nor U3457 (N_3457,N_569,N_2089);
and U3458 (N_3458,N_845,N_1484);
xnor U3459 (N_3459,N_2044,N_1070);
xnor U3460 (N_3460,N_2172,N_735);
xor U3461 (N_3461,N_346,N_1448);
nand U3462 (N_3462,N_1987,N_304);
xnor U3463 (N_3463,N_2392,N_2349);
xnor U3464 (N_3464,N_437,N_1083);
or U3465 (N_3465,N_93,N_2201);
nand U3466 (N_3466,N_1928,N_286);
nor U3467 (N_3467,N_1256,N_1315);
or U3468 (N_3468,N_2344,N_2141);
nor U3469 (N_3469,N_1063,N_1697);
xor U3470 (N_3470,N_2463,N_811);
and U3471 (N_3471,N_844,N_664);
nand U3472 (N_3472,N_1467,N_1204);
xor U3473 (N_3473,N_2276,N_2255);
or U3474 (N_3474,N_594,N_265);
nand U3475 (N_3475,N_195,N_1843);
or U3476 (N_3476,N_2355,N_1281);
and U3477 (N_3477,N_2159,N_659);
or U3478 (N_3478,N_2370,N_39);
and U3479 (N_3479,N_462,N_71);
nand U3480 (N_3480,N_2031,N_1648);
or U3481 (N_3481,N_115,N_1841);
nand U3482 (N_3482,N_279,N_110);
or U3483 (N_3483,N_245,N_2420);
and U3484 (N_3484,N_2373,N_2095);
and U3485 (N_3485,N_1781,N_512);
xor U3486 (N_3486,N_1931,N_721);
or U3487 (N_3487,N_1709,N_536);
xnor U3488 (N_3488,N_2219,N_2176);
or U3489 (N_3489,N_2444,N_2051);
and U3490 (N_3490,N_353,N_43);
nand U3491 (N_3491,N_13,N_54);
xnor U3492 (N_3492,N_130,N_1039);
nand U3493 (N_3493,N_599,N_2104);
or U3494 (N_3494,N_1730,N_1508);
or U3495 (N_3495,N_98,N_1954);
nor U3496 (N_3496,N_1522,N_303);
and U3497 (N_3497,N_1268,N_219);
nand U3498 (N_3498,N_678,N_2217);
or U3499 (N_3499,N_1440,N_1632);
nand U3500 (N_3500,N_1871,N_226);
nor U3501 (N_3501,N_2187,N_2119);
xor U3502 (N_3502,N_1629,N_1008);
nand U3503 (N_3503,N_1114,N_2368);
xor U3504 (N_3504,N_1218,N_1793);
nor U3505 (N_3505,N_1757,N_1678);
and U3506 (N_3506,N_661,N_1152);
nor U3507 (N_3507,N_937,N_2252);
or U3508 (N_3508,N_1748,N_1168);
and U3509 (N_3509,N_2383,N_448);
xor U3510 (N_3510,N_479,N_2427);
or U3511 (N_3511,N_1829,N_1891);
xor U3512 (N_3512,N_1089,N_277);
xor U3513 (N_3513,N_892,N_469);
nor U3514 (N_3514,N_887,N_210);
and U3515 (N_3515,N_657,N_1558);
and U3516 (N_3516,N_82,N_1530);
and U3517 (N_3517,N_1369,N_1384);
nor U3518 (N_3518,N_807,N_164);
nand U3519 (N_3519,N_597,N_2261);
and U3520 (N_3520,N_768,N_2216);
nand U3521 (N_3521,N_1817,N_2151);
nand U3522 (N_3522,N_1327,N_559);
nand U3523 (N_3523,N_1904,N_1999);
or U3524 (N_3524,N_142,N_240);
or U3525 (N_3525,N_1192,N_697);
and U3526 (N_3526,N_1142,N_2385);
nor U3527 (N_3527,N_685,N_1447);
xor U3528 (N_3528,N_895,N_1023);
and U3529 (N_3529,N_541,N_2206);
or U3530 (N_3530,N_2033,N_412);
nand U3531 (N_3531,N_123,N_415);
and U3532 (N_3532,N_1167,N_1084);
nor U3533 (N_3533,N_1717,N_2103);
or U3534 (N_3534,N_816,N_2210);
xor U3535 (N_3535,N_534,N_1266);
and U3536 (N_3536,N_46,N_2015);
nand U3537 (N_3537,N_1509,N_11);
and U3538 (N_3538,N_532,N_787);
and U3539 (N_3539,N_172,N_739);
xnor U3540 (N_3540,N_1758,N_545);
nor U3541 (N_3541,N_1515,N_491);
nand U3542 (N_3542,N_2205,N_44);
xor U3543 (N_3543,N_2271,N_326);
nor U3544 (N_3544,N_2365,N_1305);
or U3545 (N_3545,N_1144,N_2486);
nor U3546 (N_3546,N_921,N_511);
nor U3547 (N_3547,N_1253,N_1926);
or U3548 (N_3548,N_1630,N_2058);
nor U3549 (N_3549,N_2321,N_2293);
nor U3550 (N_3550,N_216,N_1576);
or U3551 (N_3551,N_850,N_1772);
nand U3552 (N_3552,N_2185,N_1656);
or U3553 (N_3553,N_1907,N_1421);
nor U3554 (N_3554,N_2085,N_1800);
xor U3555 (N_3555,N_1970,N_1265);
or U3556 (N_3556,N_1344,N_806);
nand U3557 (N_3557,N_947,N_2043);
and U3558 (N_3558,N_1411,N_1990);
nor U3559 (N_3559,N_2485,N_366);
nand U3560 (N_3560,N_2135,N_1944);
nor U3561 (N_3561,N_595,N_2268);
nor U3562 (N_3562,N_2213,N_2025);
and U3563 (N_3563,N_2372,N_1360);
or U3564 (N_3564,N_1544,N_945);
and U3565 (N_3565,N_593,N_920);
or U3566 (N_3566,N_992,N_144);
xor U3567 (N_3567,N_764,N_2047);
and U3568 (N_3568,N_1232,N_2002);
nor U3569 (N_3569,N_1350,N_2063);
nor U3570 (N_3570,N_649,N_799);
nor U3571 (N_3571,N_2087,N_846);
nor U3572 (N_3572,N_446,N_1090);
nand U3573 (N_3573,N_957,N_936);
and U3574 (N_3574,N_1079,N_94);
or U3575 (N_3575,N_2413,N_1473);
nand U3576 (N_3576,N_870,N_1271);
xnor U3577 (N_3577,N_355,N_571);
xnor U3578 (N_3578,N_1518,N_1243);
or U3579 (N_3579,N_373,N_2282);
or U3580 (N_3580,N_1667,N_1753);
and U3581 (N_3581,N_2180,N_406);
and U3582 (N_3582,N_191,N_2343);
and U3583 (N_3583,N_1724,N_1442);
or U3584 (N_3584,N_2228,N_675);
or U3585 (N_3585,N_2468,N_38);
xnor U3586 (N_3586,N_1622,N_2204);
nand U3587 (N_3587,N_1337,N_2380);
nand U3588 (N_3588,N_48,N_544);
or U3589 (N_3589,N_413,N_361);
nand U3590 (N_3590,N_1416,N_2464);
nor U3591 (N_3591,N_1172,N_2202);
nand U3592 (N_3592,N_607,N_744);
and U3593 (N_3593,N_1101,N_1801);
and U3594 (N_3594,N_660,N_686);
nand U3595 (N_3595,N_727,N_848);
xor U3596 (N_3596,N_420,N_2027);
xor U3597 (N_3597,N_667,N_1348);
or U3598 (N_3598,N_1564,N_504);
or U3599 (N_3599,N_693,N_314);
xnor U3600 (N_3600,N_33,N_1129);
xor U3601 (N_3601,N_51,N_2379);
xnor U3602 (N_3602,N_295,N_1364);
nor U3603 (N_3603,N_1208,N_65);
xnor U3604 (N_3604,N_958,N_1920);
and U3605 (N_3605,N_2364,N_1446);
xnor U3606 (N_3606,N_524,N_624);
nand U3607 (N_3607,N_2101,N_26);
or U3608 (N_3608,N_2396,N_464);
nor U3609 (N_3609,N_963,N_1178);
xnor U3610 (N_3610,N_2011,N_1859);
xor U3611 (N_3611,N_809,N_554);
nor U3612 (N_3612,N_1262,N_1949);
nand U3613 (N_3613,N_1423,N_1784);
nor U3614 (N_3614,N_670,N_2060);
and U3615 (N_3615,N_888,N_485);
xnor U3616 (N_3616,N_2400,N_1475);
nor U3617 (N_3617,N_708,N_187);
or U3618 (N_3618,N_1569,N_1432);
and U3619 (N_3619,N_793,N_116);
nand U3620 (N_3620,N_698,N_431);
nand U3621 (N_3621,N_1115,N_1837);
and U3622 (N_3622,N_1619,N_1517);
nor U3623 (N_3623,N_87,N_1408);
or U3624 (N_3624,N_1154,N_1489);
nor U3625 (N_3625,N_1952,N_323);
xnor U3626 (N_3626,N_2351,N_1901);
or U3627 (N_3627,N_705,N_617);
xnor U3628 (N_3628,N_734,N_486);
or U3629 (N_3629,N_1121,N_454);
and U3630 (N_3630,N_507,N_2167);
and U3631 (N_3631,N_717,N_18);
xor U3632 (N_3632,N_560,N_2099);
xnor U3633 (N_3633,N_2000,N_1963);
nand U3634 (N_3634,N_1906,N_1463);
nand U3635 (N_3635,N_492,N_924);
nand U3636 (N_3636,N_177,N_1962);
xor U3637 (N_3637,N_1613,N_1934);
xor U3638 (N_3638,N_270,N_934);
or U3639 (N_3639,N_2009,N_409);
nor U3640 (N_3640,N_1499,N_2311);
xnor U3641 (N_3641,N_2077,N_1908);
xor U3642 (N_3642,N_47,N_652);
nand U3643 (N_3643,N_1338,N_1995);
nand U3644 (N_3644,N_1747,N_2436);
nand U3645 (N_3645,N_322,N_2484);
or U3646 (N_3646,N_266,N_1568);
xor U3647 (N_3647,N_1823,N_2059);
nand U3648 (N_3648,N_519,N_980);
xor U3649 (N_3649,N_2173,N_2398);
xor U3650 (N_3650,N_2115,N_2150);
xnor U3651 (N_3651,N_821,N_2055);
nor U3652 (N_3652,N_290,N_552);
or U3653 (N_3653,N_641,N_241);
or U3654 (N_3654,N_1371,N_1614);
nor U3655 (N_3655,N_1024,N_1933);
nand U3656 (N_3656,N_2465,N_1762);
and U3657 (N_3657,N_1080,N_1778);
or U3658 (N_3658,N_632,N_284);
nand U3659 (N_3659,N_606,N_1832);
nand U3660 (N_3660,N_1392,N_2007);
nand U3661 (N_3661,N_2145,N_430);
xor U3662 (N_3662,N_932,N_1214);
nand U3663 (N_3663,N_751,N_1726);
nand U3664 (N_3664,N_256,N_1388);
nand U3665 (N_3665,N_1,N_639);
nor U3666 (N_3666,N_2262,N_574);
xor U3667 (N_3667,N_1627,N_1052);
and U3668 (N_3668,N_260,N_2086);
nand U3669 (N_3669,N_2195,N_2253);
nor U3670 (N_3670,N_2136,N_1620);
nand U3671 (N_3671,N_1481,N_2429);
xnor U3672 (N_3672,N_2275,N_114);
nor U3673 (N_3673,N_1220,N_1673);
nand U3674 (N_3674,N_1943,N_2190);
or U3675 (N_3675,N_1031,N_1274);
or U3676 (N_3676,N_24,N_1880);
and U3677 (N_3677,N_2181,N_189);
or U3678 (N_3678,N_1550,N_1903);
xnor U3679 (N_3679,N_1513,N_810);
and U3680 (N_3680,N_2019,N_99);
xnor U3681 (N_3681,N_2133,N_634);
or U3682 (N_3682,N_205,N_1537);
nor U3683 (N_3683,N_92,N_1236);
xnor U3684 (N_3684,N_1529,N_508);
nor U3685 (N_3685,N_1714,N_250);
and U3686 (N_3686,N_1982,N_1203);
nor U3687 (N_3687,N_450,N_2256);
xor U3688 (N_3688,N_2244,N_2417);
nand U3689 (N_3689,N_865,N_917);
nor U3690 (N_3690,N_255,N_146);
or U3691 (N_3691,N_1405,N_1461);
xor U3692 (N_3692,N_2284,N_885);
nor U3693 (N_3693,N_1570,N_2186);
and U3694 (N_3694,N_1988,N_2411);
nor U3695 (N_3695,N_2080,N_857);
or U3696 (N_3696,N_2292,N_755);
or U3697 (N_3697,N_1053,N_16);
xnor U3698 (N_3698,N_873,N_1978);
and U3699 (N_3699,N_1910,N_2291);
or U3700 (N_3700,N_562,N_276);
or U3701 (N_3701,N_1682,N_2122);
nand U3702 (N_3702,N_1695,N_1702);
nand U3703 (N_3703,N_1814,N_259);
nor U3704 (N_3704,N_1352,N_1809);
and U3705 (N_3705,N_2110,N_1210);
nand U3706 (N_3706,N_1472,N_1783);
nand U3707 (N_3707,N_14,N_1552);
nor U3708 (N_3708,N_586,N_949);
or U3709 (N_3709,N_951,N_1631);
or U3710 (N_3710,N_438,N_762);
nor U3711 (N_3711,N_1838,N_1356);
nand U3712 (N_3712,N_2004,N_1740);
nand U3713 (N_3713,N_1240,N_640);
nand U3714 (N_3714,N_1719,N_1137);
and U3715 (N_3715,N_994,N_1242);
and U3716 (N_3716,N_370,N_1706);
nor U3717 (N_3717,N_1519,N_944);
xor U3718 (N_3718,N_1054,N_50);
and U3719 (N_3719,N_778,N_823);
nand U3720 (N_3720,N_1244,N_1731);
or U3721 (N_3721,N_790,N_985);
or U3722 (N_3722,N_53,N_23);
nor U3723 (N_3723,N_1032,N_236);
nor U3724 (N_3724,N_273,N_1465);
and U3725 (N_3725,N_395,N_29);
and U3726 (N_3726,N_1785,N_2443);
nor U3727 (N_3727,N_383,N_2347);
xnor U3728 (N_3728,N_1559,N_1036);
and U3729 (N_3729,N_1189,N_538);
nor U3730 (N_3730,N_122,N_666);
or U3731 (N_3731,N_1585,N_1162);
xnor U3732 (N_3732,N_1497,N_316);
nor U3733 (N_3733,N_2393,N_1870);
nor U3734 (N_3734,N_2184,N_868);
nand U3735 (N_3735,N_2267,N_1193);
or U3736 (N_3736,N_1869,N_1794);
nor U3737 (N_3737,N_525,N_1221);
or U3738 (N_3738,N_416,N_1936);
xor U3739 (N_3739,N_278,N_950);
and U3740 (N_3740,N_1532,N_1738);
nor U3741 (N_3741,N_2065,N_1328);
or U3742 (N_3742,N_2367,N_1247);
xor U3743 (N_3743,N_392,N_1105);
xor U3744 (N_3744,N_517,N_909);
xnor U3745 (N_3745,N_1055,N_1549);
nor U3746 (N_3746,N_1708,N_1997);
xor U3747 (N_3747,N_1855,N_671);
or U3748 (N_3748,N_812,N_377);
nand U3749 (N_3749,N_1973,N_1370);
or U3750 (N_3750,N_634,N_1343);
nor U3751 (N_3751,N_1096,N_2131);
and U3752 (N_3752,N_676,N_2383);
nand U3753 (N_3753,N_67,N_1186);
and U3754 (N_3754,N_818,N_1740);
nor U3755 (N_3755,N_1690,N_1677);
xnor U3756 (N_3756,N_1402,N_1620);
or U3757 (N_3757,N_1437,N_1909);
xnor U3758 (N_3758,N_1513,N_808);
and U3759 (N_3759,N_1521,N_2361);
and U3760 (N_3760,N_325,N_1579);
or U3761 (N_3761,N_2211,N_577);
nor U3762 (N_3762,N_330,N_656);
nor U3763 (N_3763,N_2018,N_1049);
and U3764 (N_3764,N_888,N_2492);
xnor U3765 (N_3765,N_76,N_2146);
or U3766 (N_3766,N_1987,N_769);
nand U3767 (N_3767,N_63,N_89);
and U3768 (N_3768,N_549,N_1319);
xnor U3769 (N_3769,N_1709,N_1961);
nand U3770 (N_3770,N_1701,N_826);
or U3771 (N_3771,N_2321,N_1751);
xor U3772 (N_3772,N_174,N_2170);
nand U3773 (N_3773,N_2126,N_1149);
or U3774 (N_3774,N_2127,N_1309);
nand U3775 (N_3775,N_143,N_1394);
nand U3776 (N_3776,N_5,N_596);
or U3777 (N_3777,N_883,N_1887);
nand U3778 (N_3778,N_1439,N_1939);
and U3779 (N_3779,N_987,N_2222);
or U3780 (N_3780,N_1205,N_494);
nor U3781 (N_3781,N_244,N_1376);
and U3782 (N_3782,N_2486,N_2332);
nand U3783 (N_3783,N_563,N_1379);
and U3784 (N_3784,N_2052,N_1670);
nand U3785 (N_3785,N_2065,N_2003);
and U3786 (N_3786,N_259,N_420);
nor U3787 (N_3787,N_2441,N_880);
nor U3788 (N_3788,N_1405,N_2437);
nor U3789 (N_3789,N_1336,N_814);
nor U3790 (N_3790,N_442,N_382);
or U3791 (N_3791,N_1179,N_879);
or U3792 (N_3792,N_482,N_2041);
nor U3793 (N_3793,N_120,N_2402);
xor U3794 (N_3794,N_469,N_2113);
nor U3795 (N_3795,N_1448,N_912);
nor U3796 (N_3796,N_1520,N_2413);
nor U3797 (N_3797,N_1647,N_2230);
or U3798 (N_3798,N_226,N_797);
or U3799 (N_3799,N_28,N_1666);
and U3800 (N_3800,N_335,N_1291);
or U3801 (N_3801,N_1612,N_437);
and U3802 (N_3802,N_2191,N_1066);
xor U3803 (N_3803,N_102,N_1364);
nand U3804 (N_3804,N_1334,N_1868);
nand U3805 (N_3805,N_890,N_532);
nor U3806 (N_3806,N_858,N_1806);
and U3807 (N_3807,N_2324,N_1782);
and U3808 (N_3808,N_1641,N_2340);
and U3809 (N_3809,N_862,N_2161);
or U3810 (N_3810,N_15,N_549);
nand U3811 (N_3811,N_2318,N_509);
nor U3812 (N_3812,N_703,N_962);
xnor U3813 (N_3813,N_232,N_2168);
nor U3814 (N_3814,N_1693,N_1123);
or U3815 (N_3815,N_1678,N_2470);
and U3816 (N_3816,N_924,N_1011);
xor U3817 (N_3817,N_888,N_2180);
and U3818 (N_3818,N_1614,N_103);
or U3819 (N_3819,N_2460,N_149);
or U3820 (N_3820,N_87,N_1179);
nand U3821 (N_3821,N_162,N_1052);
nand U3822 (N_3822,N_1034,N_2039);
and U3823 (N_3823,N_651,N_1744);
nand U3824 (N_3824,N_1829,N_1258);
nand U3825 (N_3825,N_1637,N_895);
xor U3826 (N_3826,N_1101,N_441);
xnor U3827 (N_3827,N_2329,N_719);
xnor U3828 (N_3828,N_1454,N_2058);
or U3829 (N_3829,N_558,N_1811);
nand U3830 (N_3830,N_394,N_1081);
and U3831 (N_3831,N_1717,N_2384);
and U3832 (N_3832,N_352,N_1484);
xor U3833 (N_3833,N_2495,N_1719);
and U3834 (N_3834,N_2235,N_2094);
xor U3835 (N_3835,N_1281,N_2311);
xor U3836 (N_3836,N_1979,N_1900);
or U3837 (N_3837,N_420,N_1430);
and U3838 (N_3838,N_517,N_1355);
or U3839 (N_3839,N_734,N_205);
nor U3840 (N_3840,N_1759,N_2208);
nand U3841 (N_3841,N_1675,N_187);
xor U3842 (N_3842,N_1859,N_757);
and U3843 (N_3843,N_195,N_2028);
nor U3844 (N_3844,N_236,N_1475);
and U3845 (N_3845,N_742,N_179);
xnor U3846 (N_3846,N_3,N_2038);
and U3847 (N_3847,N_455,N_634);
xor U3848 (N_3848,N_929,N_1191);
nor U3849 (N_3849,N_2379,N_928);
and U3850 (N_3850,N_1312,N_1826);
xor U3851 (N_3851,N_2314,N_1614);
nand U3852 (N_3852,N_235,N_2322);
xor U3853 (N_3853,N_1954,N_1595);
and U3854 (N_3854,N_2028,N_151);
and U3855 (N_3855,N_574,N_1514);
or U3856 (N_3856,N_1011,N_1610);
or U3857 (N_3857,N_1220,N_2423);
and U3858 (N_3858,N_1628,N_359);
nor U3859 (N_3859,N_625,N_2496);
or U3860 (N_3860,N_1970,N_1001);
nand U3861 (N_3861,N_2328,N_1315);
xor U3862 (N_3862,N_2381,N_723);
or U3863 (N_3863,N_2230,N_2313);
xnor U3864 (N_3864,N_1421,N_765);
and U3865 (N_3865,N_1527,N_350);
xor U3866 (N_3866,N_1940,N_2068);
and U3867 (N_3867,N_21,N_2034);
and U3868 (N_3868,N_295,N_319);
nor U3869 (N_3869,N_48,N_2320);
nand U3870 (N_3870,N_929,N_655);
or U3871 (N_3871,N_2320,N_962);
or U3872 (N_3872,N_2437,N_1650);
xor U3873 (N_3873,N_964,N_1349);
or U3874 (N_3874,N_611,N_2256);
nor U3875 (N_3875,N_2211,N_197);
or U3876 (N_3876,N_2471,N_454);
nand U3877 (N_3877,N_812,N_500);
xor U3878 (N_3878,N_755,N_1327);
or U3879 (N_3879,N_1824,N_745);
nor U3880 (N_3880,N_2005,N_12);
and U3881 (N_3881,N_2465,N_418);
xor U3882 (N_3882,N_531,N_1879);
or U3883 (N_3883,N_1359,N_1483);
xnor U3884 (N_3884,N_512,N_167);
or U3885 (N_3885,N_527,N_2398);
nor U3886 (N_3886,N_618,N_1084);
nor U3887 (N_3887,N_2186,N_635);
xor U3888 (N_3888,N_1741,N_1685);
and U3889 (N_3889,N_792,N_2038);
xor U3890 (N_3890,N_32,N_18);
nand U3891 (N_3891,N_864,N_2108);
xnor U3892 (N_3892,N_1163,N_961);
nor U3893 (N_3893,N_1737,N_708);
and U3894 (N_3894,N_902,N_60);
or U3895 (N_3895,N_1771,N_2126);
or U3896 (N_3896,N_159,N_2428);
xnor U3897 (N_3897,N_1765,N_2082);
xor U3898 (N_3898,N_1266,N_107);
or U3899 (N_3899,N_630,N_2334);
xor U3900 (N_3900,N_889,N_197);
and U3901 (N_3901,N_1538,N_346);
and U3902 (N_3902,N_56,N_1917);
and U3903 (N_3903,N_29,N_556);
xnor U3904 (N_3904,N_1143,N_2202);
and U3905 (N_3905,N_25,N_1892);
nand U3906 (N_3906,N_2084,N_1742);
xor U3907 (N_3907,N_1392,N_171);
or U3908 (N_3908,N_184,N_849);
xnor U3909 (N_3909,N_188,N_1944);
or U3910 (N_3910,N_1288,N_1509);
xnor U3911 (N_3911,N_2143,N_1280);
nand U3912 (N_3912,N_696,N_1895);
nand U3913 (N_3913,N_744,N_651);
nand U3914 (N_3914,N_1073,N_1521);
nor U3915 (N_3915,N_431,N_697);
xnor U3916 (N_3916,N_648,N_1320);
nor U3917 (N_3917,N_1806,N_1518);
xnor U3918 (N_3918,N_1856,N_424);
nor U3919 (N_3919,N_2376,N_550);
nand U3920 (N_3920,N_1432,N_1710);
xor U3921 (N_3921,N_695,N_74);
or U3922 (N_3922,N_1598,N_873);
or U3923 (N_3923,N_1433,N_396);
nor U3924 (N_3924,N_1643,N_1372);
xor U3925 (N_3925,N_2463,N_874);
nor U3926 (N_3926,N_1458,N_2015);
xnor U3927 (N_3927,N_1116,N_1568);
or U3928 (N_3928,N_1878,N_591);
nor U3929 (N_3929,N_1369,N_863);
xor U3930 (N_3930,N_1268,N_664);
xnor U3931 (N_3931,N_1070,N_1658);
nand U3932 (N_3932,N_1541,N_556);
xor U3933 (N_3933,N_1365,N_1341);
and U3934 (N_3934,N_1940,N_615);
or U3935 (N_3935,N_1347,N_1989);
nand U3936 (N_3936,N_489,N_2367);
and U3937 (N_3937,N_2098,N_37);
xnor U3938 (N_3938,N_15,N_1958);
and U3939 (N_3939,N_1158,N_8);
nor U3940 (N_3940,N_1618,N_2108);
nand U3941 (N_3941,N_208,N_2467);
nand U3942 (N_3942,N_702,N_1541);
or U3943 (N_3943,N_530,N_449);
nand U3944 (N_3944,N_966,N_1553);
xnor U3945 (N_3945,N_1083,N_2349);
nand U3946 (N_3946,N_1524,N_473);
and U3947 (N_3947,N_624,N_1996);
xnor U3948 (N_3948,N_2324,N_2446);
or U3949 (N_3949,N_1603,N_1161);
nor U3950 (N_3950,N_1639,N_2195);
nor U3951 (N_3951,N_418,N_542);
xnor U3952 (N_3952,N_2140,N_669);
nand U3953 (N_3953,N_574,N_1774);
xnor U3954 (N_3954,N_1069,N_559);
nand U3955 (N_3955,N_1822,N_93);
nand U3956 (N_3956,N_2175,N_1194);
xnor U3957 (N_3957,N_485,N_1684);
xnor U3958 (N_3958,N_1591,N_1533);
xor U3959 (N_3959,N_2339,N_264);
or U3960 (N_3960,N_242,N_1784);
and U3961 (N_3961,N_628,N_893);
nand U3962 (N_3962,N_2417,N_1886);
nand U3963 (N_3963,N_225,N_442);
nand U3964 (N_3964,N_1107,N_1430);
nor U3965 (N_3965,N_1863,N_453);
xnor U3966 (N_3966,N_553,N_2046);
nor U3967 (N_3967,N_2361,N_2329);
or U3968 (N_3968,N_884,N_1142);
nand U3969 (N_3969,N_2224,N_887);
and U3970 (N_3970,N_1853,N_1725);
nand U3971 (N_3971,N_1198,N_1008);
nand U3972 (N_3972,N_1264,N_2270);
xor U3973 (N_3973,N_1906,N_2121);
or U3974 (N_3974,N_284,N_981);
and U3975 (N_3975,N_2034,N_1428);
nand U3976 (N_3976,N_167,N_2056);
nand U3977 (N_3977,N_1462,N_396);
nand U3978 (N_3978,N_1120,N_372);
nor U3979 (N_3979,N_250,N_106);
xnor U3980 (N_3980,N_700,N_2419);
nor U3981 (N_3981,N_69,N_1381);
or U3982 (N_3982,N_1487,N_2033);
nand U3983 (N_3983,N_1927,N_476);
xnor U3984 (N_3984,N_1772,N_178);
nor U3985 (N_3985,N_747,N_1140);
nor U3986 (N_3986,N_1373,N_784);
xnor U3987 (N_3987,N_2404,N_1841);
xor U3988 (N_3988,N_2461,N_778);
nand U3989 (N_3989,N_684,N_848);
nor U3990 (N_3990,N_711,N_858);
nand U3991 (N_3991,N_1429,N_1244);
or U3992 (N_3992,N_2137,N_1649);
nand U3993 (N_3993,N_1205,N_273);
or U3994 (N_3994,N_277,N_249);
xor U3995 (N_3995,N_800,N_1582);
and U3996 (N_3996,N_1171,N_1233);
nand U3997 (N_3997,N_1063,N_1098);
xnor U3998 (N_3998,N_945,N_1511);
nand U3999 (N_3999,N_167,N_1760);
xnor U4000 (N_4000,N_186,N_532);
or U4001 (N_4001,N_458,N_418);
nand U4002 (N_4002,N_180,N_1120);
xor U4003 (N_4003,N_586,N_2354);
xor U4004 (N_4004,N_1156,N_308);
nand U4005 (N_4005,N_417,N_1594);
nor U4006 (N_4006,N_2082,N_1019);
or U4007 (N_4007,N_447,N_2266);
nand U4008 (N_4008,N_1446,N_163);
nor U4009 (N_4009,N_813,N_1689);
nor U4010 (N_4010,N_813,N_1429);
or U4011 (N_4011,N_1544,N_226);
or U4012 (N_4012,N_1305,N_1092);
xnor U4013 (N_4013,N_1684,N_1812);
nor U4014 (N_4014,N_77,N_16);
and U4015 (N_4015,N_368,N_341);
nand U4016 (N_4016,N_1854,N_1198);
nand U4017 (N_4017,N_1407,N_2403);
or U4018 (N_4018,N_1809,N_981);
nand U4019 (N_4019,N_1791,N_423);
nor U4020 (N_4020,N_2040,N_1952);
nand U4021 (N_4021,N_707,N_1617);
nor U4022 (N_4022,N_1554,N_131);
xor U4023 (N_4023,N_14,N_758);
xnor U4024 (N_4024,N_1953,N_440);
nand U4025 (N_4025,N_1953,N_1613);
or U4026 (N_4026,N_2098,N_209);
xnor U4027 (N_4027,N_2039,N_2413);
nor U4028 (N_4028,N_68,N_2148);
xor U4029 (N_4029,N_562,N_342);
nor U4030 (N_4030,N_1445,N_784);
nor U4031 (N_4031,N_859,N_1410);
xor U4032 (N_4032,N_2388,N_1606);
or U4033 (N_4033,N_1041,N_578);
xnor U4034 (N_4034,N_799,N_2293);
nor U4035 (N_4035,N_2330,N_1072);
nor U4036 (N_4036,N_594,N_476);
nand U4037 (N_4037,N_1869,N_538);
nand U4038 (N_4038,N_977,N_2196);
nor U4039 (N_4039,N_1639,N_368);
nor U4040 (N_4040,N_2408,N_2133);
and U4041 (N_4041,N_1933,N_1369);
xnor U4042 (N_4042,N_2163,N_1688);
nor U4043 (N_4043,N_506,N_215);
or U4044 (N_4044,N_2223,N_2332);
nand U4045 (N_4045,N_577,N_5);
and U4046 (N_4046,N_842,N_929);
and U4047 (N_4047,N_284,N_187);
or U4048 (N_4048,N_966,N_1688);
nand U4049 (N_4049,N_349,N_2454);
and U4050 (N_4050,N_2092,N_1984);
nor U4051 (N_4051,N_1098,N_1707);
or U4052 (N_4052,N_1564,N_497);
xor U4053 (N_4053,N_32,N_968);
or U4054 (N_4054,N_1461,N_2062);
xor U4055 (N_4055,N_2448,N_2409);
nand U4056 (N_4056,N_1894,N_1256);
xor U4057 (N_4057,N_75,N_863);
or U4058 (N_4058,N_1415,N_2269);
and U4059 (N_4059,N_869,N_698);
and U4060 (N_4060,N_515,N_605);
or U4061 (N_4061,N_2492,N_2024);
nand U4062 (N_4062,N_1436,N_2312);
nor U4063 (N_4063,N_1561,N_797);
nor U4064 (N_4064,N_1595,N_1634);
xnor U4065 (N_4065,N_2007,N_993);
or U4066 (N_4066,N_1650,N_1413);
xnor U4067 (N_4067,N_2324,N_1573);
nor U4068 (N_4068,N_2210,N_1450);
xnor U4069 (N_4069,N_1155,N_761);
xnor U4070 (N_4070,N_1416,N_830);
xnor U4071 (N_4071,N_1842,N_242);
and U4072 (N_4072,N_115,N_341);
xor U4073 (N_4073,N_1896,N_333);
xnor U4074 (N_4074,N_156,N_79);
or U4075 (N_4075,N_1867,N_1383);
xor U4076 (N_4076,N_1258,N_422);
or U4077 (N_4077,N_1949,N_136);
nand U4078 (N_4078,N_1910,N_835);
xnor U4079 (N_4079,N_2093,N_1965);
nand U4080 (N_4080,N_853,N_864);
xor U4081 (N_4081,N_1142,N_940);
nor U4082 (N_4082,N_680,N_1887);
nor U4083 (N_4083,N_2089,N_594);
and U4084 (N_4084,N_2155,N_2062);
nand U4085 (N_4085,N_396,N_1084);
nor U4086 (N_4086,N_1976,N_1639);
nor U4087 (N_4087,N_1638,N_1517);
xnor U4088 (N_4088,N_1248,N_1292);
nor U4089 (N_4089,N_1819,N_22);
nand U4090 (N_4090,N_250,N_1198);
nor U4091 (N_4091,N_2271,N_1212);
nand U4092 (N_4092,N_162,N_1790);
nand U4093 (N_4093,N_1833,N_1905);
or U4094 (N_4094,N_107,N_7);
xor U4095 (N_4095,N_292,N_349);
and U4096 (N_4096,N_2292,N_1323);
and U4097 (N_4097,N_1294,N_2109);
nor U4098 (N_4098,N_1461,N_2486);
nor U4099 (N_4099,N_511,N_174);
nand U4100 (N_4100,N_1626,N_774);
nand U4101 (N_4101,N_663,N_993);
xor U4102 (N_4102,N_667,N_1620);
or U4103 (N_4103,N_2048,N_2252);
nand U4104 (N_4104,N_1872,N_1743);
xnor U4105 (N_4105,N_1914,N_376);
nand U4106 (N_4106,N_410,N_431);
xnor U4107 (N_4107,N_1746,N_525);
and U4108 (N_4108,N_705,N_818);
and U4109 (N_4109,N_1266,N_100);
nand U4110 (N_4110,N_1493,N_1616);
and U4111 (N_4111,N_1253,N_1931);
and U4112 (N_4112,N_156,N_1549);
and U4113 (N_4113,N_1326,N_1937);
or U4114 (N_4114,N_573,N_1552);
nand U4115 (N_4115,N_2321,N_1178);
nand U4116 (N_4116,N_1399,N_75);
nor U4117 (N_4117,N_1979,N_872);
nand U4118 (N_4118,N_923,N_219);
nor U4119 (N_4119,N_1519,N_2307);
xnor U4120 (N_4120,N_1571,N_599);
or U4121 (N_4121,N_2372,N_1314);
or U4122 (N_4122,N_0,N_2038);
and U4123 (N_4123,N_2114,N_1136);
or U4124 (N_4124,N_956,N_908);
and U4125 (N_4125,N_106,N_1906);
and U4126 (N_4126,N_2300,N_751);
and U4127 (N_4127,N_488,N_142);
or U4128 (N_4128,N_1858,N_1532);
xnor U4129 (N_4129,N_950,N_1203);
or U4130 (N_4130,N_2332,N_2095);
nand U4131 (N_4131,N_737,N_91);
nor U4132 (N_4132,N_1313,N_1632);
nand U4133 (N_4133,N_2483,N_192);
or U4134 (N_4134,N_343,N_1842);
nand U4135 (N_4135,N_2212,N_423);
or U4136 (N_4136,N_1109,N_895);
and U4137 (N_4137,N_1547,N_2375);
and U4138 (N_4138,N_1228,N_2170);
and U4139 (N_4139,N_1878,N_409);
or U4140 (N_4140,N_2093,N_832);
nand U4141 (N_4141,N_107,N_1815);
xor U4142 (N_4142,N_768,N_698);
nand U4143 (N_4143,N_196,N_2211);
nor U4144 (N_4144,N_1681,N_1747);
or U4145 (N_4145,N_1250,N_1674);
nor U4146 (N_4146,N_1830,N_371);
and U4147 (N_4147,N_1169,N_715);
xor U4148 (N_4148,N_19,N_2470);
and U4149 (N_4149,N_1935,N_2139);
nor U4150 (N_4150,N_1675,N_873);
xor U4151 (N_4151,N_2402,N_1411);
or U4152 (N_4152,N_1450,N_1172);
nand U4153 (N_4153,N_763,N_1207);
nand U4154 (N_4154,N_470,N_1581);
nand U4155 (N_4155,N_2182,N_266);
nand U4156 (N_4156,N_65,N_21);
nand U4157 (N_4157,N_625,N_172);
nor U4158 (N_4158,N_2320,N_1382);
nor U4159 (N_4159,N_2254,N_1070);
nor U4160 (N_4160,N_1092,N_998);
nand U4161 (N_4161,N_2050,N_2278);
nand U4162 (N_4162,N_2400,N_2366);
and U4163 (N_4163,N_1630,N_1515);
or U4164 (N_4164,N_2338,N_2232);
nand U4165 (N_4165,N_1116,N_822);
nor U4166 (N_4166,N_1162,N_1557);
nand U4167 (N_4167,N_2198,N_1855);
xnor U4168 (N_4168,N_1083,N_2490);
nor U4169 (N_4169,N_199,N_1198);
or U4170 (N_4170,N_433,N_954);
or U4171 (N_4171,N_1621,N_777);
xor U4172 (N_4172,N_815,N_882);
nand U4173 (N_4173,N_179,N_2116);
xor U4174 (N_4174,N_378,N_2456);
xnor U4175 (N_4175,N_161,N_1468);
xnor U4176 (N_4176,N_656,N_2154);
nand U4177 (N_4177,N_2352,N_1207);
nand U4178 (N_4178,N_942,N_1452);
nand U4179 (N_4179,N_142,N_1456);
or U4180 (N_4180,N_834,N_2332);
nand U4181 (N_4181,N_1554,N_2323);
nand U4182 (N_4182,N_1602,N_536);
xor U4183 (N_4183,N_2483,N_1794);
nand U4184 (N_4184,N_394,N_2293);
and U4185 (N_4185,N_2009,N_676);
and U4186 (N_4186,N_1783,N_301);
xnor U4187 (N_4187,N_1850,N_477);
or U4188 (N_4188,N_744,N_1743);
and U4189 (N_4189,N_524,N_332);
nand U4190 (N_4190,N_1229,N_777);
xor U4191 (N_4191,N_548,N_2365);
or U4192 (N_4192,N_1012,N_1598);
xnor U4193 (N_4193,N_720,N_755);
and U4194 (N_4194,N_2328,N_721);
nand U4195 (N_4195,N_307,N_324);
xnor U4196 (N_4196,N_2480,N_2388);
xor U4197 (N_4197,N_51,N_866);
xnor U4198 (N_4198,N_2204,N_2389);
nand U4199 (N_4199,N_1867,N_1418);
and U4200 (N_4200,N_1447,N_1448);
or U4201 (N_4201,N_1134,N_1522);
xor U4202 (N_4202,N_1684,N_523);
nand U4203 (N_4203,N_1061,N_249);
xor U4204 (N_4204,N_1068,N_288);
nor U4205 (N_4205,N_279,N_1546);
nand U4206 (N_4206,N_2188,N_212);
nand U4207 (N_4207,N_2247,N_2267);
and U4208 (N_4208,N_2271,N_1130);
nand U4209 (N_4209,N_1012,N_663);
nand U4210 (N_4210,N_1832,N_1321);
or U4211 (N_4211,N_798,N_34);
or U4212 (N_4212,N_808,N_485);
nand U4213 (N_4213,N_1026,N_638);
or U4214 (N_4214,N_235,N_1667);
or U4215 (N_4215,N_1951,N_2332);
xor U4216 (N_4216,N_1559,N_609);
xor U4217 (N_4217,N_678,N_1663);
nand U4218 (N_4218,N_1451,N_2204);
and U4219 (N_4219,N_1468,N_439);
and U4220 (N_4220,N_65,N_823);
nor U4221 (N_4221,N_675,N_1642);
nand U4222 (N_4222,N_2171,N_2312);
or U4223 (N_4223,N_69,N_1763);
nor U4224 (N_4224,N_2205,N_2207);
nor U4225 (N_4225,N_684,N_1804);
nand U4226 (N_4226,N_729,N_2019);
or U4227 (N_4227,N_2441,N_1970);
and U4228 (N_4228,N_764,N_2344);
or U4229 (N_4229,N_2092,N_635);
nor U4230 (N_4230,N_349,N_287);
or U4231 (N_4231,N_2114,N_1544);
nor U4232 (N_4232,N_2174,N_454);
nor U4233 (N_4233,N_1217,N_178);
and U4234 (N_4234,N_2133,N_177);
nor U4235 (N_4235,N_2362,N_1352);
xor U4236 (N_4236,N_311,N_366);
and U4237 (N_4237,N_753,N_1880);
and U4238 (N_4238,N_405,N_1617);
or U4239 (N_4239,N_2409,N_1723);
or U4240 (N_4240,N_1003,N_1572);
and U4241 (N_4241,N_2137,N_867);
xnor U4242 (N_4242,N_1745,N_1953);
nand U4243 (N_4243,N_1574,N_1468);
nand U4244 (N_4244,N_991,N_274);
and U4245 (N_4245,N_1348,N_132);
xor U4246 (N_4246,N_602,N_676);
xor U4247 (N_4247,N_14,N_1779);
and U4248 (N_4248,N_281,N_2359);
xnor U4249 (N_4249,N_640,N_1799);
and U4250 (N_4250,N_509,N_1320);
nand U4251 (N_4251,N_1220,N_1147);
nand U4252 (N_4252,N_687,N_417);
nand U4253 (N_4253,N_2064,N_1263);
xor U4254 (N_4254,N_1021,N_287);
or U4255 (N_4255,N_1970,N_1876);
xnor U4256 (N_4256,N_1216,N_2405);
nor U4257 (N_4257,N_702,N_748);
xor U4258 (N_4258,N_1323,N_1541);
and U4259 (N_4259,N_666,N_1749);
xor U4260 (N_4260,N_1112,N_881);
and U4261 (N_4261,N_1891,N_1795);
xor U4262 (N_4262,N_285,N_761);
and U4263 (N_4263,N_1796,N_178);
nor U4264 (N_4264,N_1159,N_1722);
and U4265 (N_4265,N_975,N_849);
nor U4266 (N_4266,N_1316,N_2300);
and U4267 (N_4267,N_662,N_752);
and U4268 (N_4268,N_2427,N_1486);
nand U4269 (N_4269,N_779,N_690);
nor U4270 (N_4270,N_2188,N_361);
nor U4271 (N_4271,N_1631,N_235);
or U4272 (N_4272,N_1872,N_361);
or U4273 (N_4273,N_125,N_2217);
xor U4274 (N_4274,N_715,N_1852);
and U4275 (N_4275,N_1195,N_1091);
or U4276 (N_4276,N_1006,N_1863);
nand U4277 (N_4277,N_677,N_1133);
nand U4278 (N_4278,N_2401,N_1821);
or U4279 (N_4279,N_2027,N_914);
or U4280 (N_4280,N_737,N_1491);
nand U4281 (N_4281,N_1700,N_180);
or U4282 (N_4282,N_120,N_1880);
xnor U4283 (N_4283,N_1205,N_1809);
nor U4284 (N_4284,N_1957,N_1482);
or U4285 (N_4285,N_1679,N_120);
or U4286 (N_4286,N_60,N_88);
nand U4287 (N_4287,N_152,N_2320);
nor U4288 (N_4288,N_917,N_2475);
nand U4289 (N_4289,N_2331,N_1507);
nor U4290 (N_4290,N_2271,N_777);
nor U4291 (N_4291,N_32,N_1482);
and U4292 (N_4292,N_430,N_611);
nand U4293 (N_4293,N_679,N_2203);
and U4294 (N_4294,N_2361,N_1542);
xnor U4295 (N_4295,N_1938,N_749);
and U4296 (N_4296,N_613,N_2142);
nor U4297 (N_4297,N_2476,N_1544);
nand U4298 (N_4298,N_996,N_378);
nor U4299 (N_4299,N_1980,N_692);
nand U4300 (N_4300,N_2490,N_2445);
or U4301 (N_4301,N_1657,N_324);
or U4302 (N_4302,N_1234,N_1636);
nand U4303 (N_4303,N_2243,N_2102);
xnor U4304 (N_4304,N_1436,N_1937);
nand U4305 (N_4305,N_2122,N_987);
and U4306 (N_4306,N_837,N_2498);
or U4307 (N_4307,N_1903,N_1119);
xnor U4308 (N_4308,N_1723,N_1820);
nor U4309 (N_4309,N_1382,N_683);
or U4310 (N_4310,N_1323,N_1282);
or U4311 (N_4311,N_1465,N_699);
nand U4312 (N_4312,N_1328,N_1948);
and U4313 (N_4313,N_864,N_1850);
and U4314 (N_4314,N_1838,N_2450);
nand U4315 (N_4315,N_1815,N_1256);
or U4316 (N_4316,N_912,N_1711);
and U4317 (N_4317,N_34,N_203);
nand U4318 (N_4318,N_879,N_1523);
nor U4319 (N_4319,N_1182,N_1944);
nand U4320 (N_4320,N_145,N_1699);
nand U4321 (N_4321,N_973,N_1140);
or U4322 (N_4322,N_504,N_936);
nand U4323 (N_4323,N_1297,N_1903);
or U4324 (N_4324,N_1684,N_908);
nand U4325 (N_4325,N_1049,N_308);
or U4326 (N_4326,N_1386,N_1866);
nand U4327 (N_4327,N_1254,N_663);
xor U4328 (N_4328,N_1851,N_353);
xor U4329 (N_4329,N_849,N_196);
nor U4330 (N_4330,N_1210,N_625);
nor U4331 (N_4331,N_1342,N_1494);
and U4332 (N_4332,N_1570,N_2244);
xnor U4333 (N_4333,N_933,N_1901);
nor U4334 (N_4334,N_2012,N_232);
or U4335 (N_4335,N_166,N_1733);
xor U4336 (N_4336,N_759,N_2123);
xor U4337 (N_4337,N_505,N_462);
nand U4338 (N_4338,N_6,N_1451);
nand U4339 (N_4339,N_1504,N_552);
nor U4340 (N_4340,N_88,N_579);
xor U4341 (N_4341,N_238,N_1716);
and U4342 (N_4342,N_510,N_498);
or U4343 (N_4343,N_1103,N_471);
or U4344 (N_4344,N_2195,N_709);
nand U4345 (N_4345,N_1323,N_398);
or U4346 (N_4346,N_1555,N_858);
xnor U4347 (N_4347,N_373,N_841);
nor U4348 (N_4348,N_1614,N_736);
nor U4349 (N_4349,N_2310,N_312);
and U4350 (N_4350,N_1264,N_1197);
and U4351 (N_4351,N_2015,N_2020);
nand U4352 (N_4352,N_733,N_1178);
or U4353 (N_4353,N_125,N_1701);
nand U4354 (N_4354,N_1944,N_2142);
and U4355 (N_4355,N_2270,N_2301);
nor U4356 (N_4356,N_734,N_379);
or U4357 (N_4357,N_677,N_871);
or U4358 (N_4358,N_1696,N_904);
xnor U4359 (N_4359,N_245,N_242);
and U4360 (N_4360,N_1892,N_776);
nand U4361 (N_4361,N_2389,N_694);
or U4362 (N_4362,N_930,N_1116);
and U4363 (N_4363,N_1868,N_696);
nand U4364 (N_4364,N_2183,N_677);
xnor U4365 (N_4365,N_1323,N_974);
or U4366 (N_4366,N_869,N_1515);
nor U4367 (N_4367,N_128,N_636);
or U4368 (N_4368,N_55,N_511);
and U4369 (N_4369,N_2426,N_1320);
xor U4370 (N_4370,N_1957,N_1905);
nand U4371 (N_4371,N_506,N_18);
xnor U4372 (N_4372,N_1376,N_2388);
xor U4373 (N_4373,N_784,N_608);
and U4374 (N_4374,N_2047,N_1126);
and U4375 (N_4375,N_488,N_2009);
nor U4376 (N_4376,N_1663,N_906);
xor U4377 (N_4377,N_299,N_777);
nor U4378 (N_4378,N_2156,N_1513);
and U4379 (N_4379,N_1848,N_433);
nor U4380 (N_4380,N_1308,N_1408);
xnor U4381 (N_4381,N_2399,N_1517);
nand U4382 (N_4382,N_1444,N_2026);
xnor U4383 (N_4383,N_771,N_1260);
nand U4384 (N_4384,N_109,N_1077);
or U4385 (N_4385,N_1388,N_2000);
nor U4386 (N_4386,N_78,N_102);
and U4387 (N_4387,N_1018,N_46);
nor U4388 (N_4388,N_1734,N_1202);
nor U4389 (N_4389,N_694,N_1750);
and U4390 (N_4390,N_928,N_742);
nor U4391 (N_4391,N_536,N_2225);
nor U4392 (N_4392,N_889,N_616);
xnor U4393 (N_4393,N_287,N_1705);
or U4394 (N_4394,N_1729,N_1509);
xnor U4395 (N_4395,N_1726,N_2034);
and U4396 (N_4396,N_2489,N_1612);
nor U4397 (N_4397,N_1693,N_691);
xnor U4398 (N_4398,N_1973,N_2252);
xor U4399 (N_4399,N_753,N_1422);
or U4400 (N_4400,N_1577,N_1721);
and U4401 (N_4401,N_1397,N_2147);
nor U4402 (N_4402,N_1492,N_2242);
nor U4403 (N_4403,N_9,N_168);
nand U4404 (N_4404,N_2211,N_1483);
xor U4405 (N_4405,N_408,N_1994);
or U4406 (N_4406,N_988,N_407);
or U4407 (N_4407,N_1181,N_516);
and U4408 (N_4408,N_311,N_1743);
nand U4409 (N_4409,N_846,N_2436);
xnor U4410 (N_4410,N_210,N_1790);
nor U4411 (N_4411,N_1488,N_1418);
xor U4412 (N_4412,N_1173,N_1067);
xor U4413 (N_4413,N_1082,N_2221);
and U4414 (N_4414,N_2487,N_2040);
nor U4415 (N_4415,N_2467,N_2053);
xnor U4416 (N_4416,N_2375,N_2396);
or U4417 (N_4417,N_871,N_778);
nand U4418 (N_4418,N_736,N_843);
xor U4419 (N_4419,N_848,N_763);
and U4420 (N_4420,N_454,N_1383);
nand U4421 (N_4421,N_1568,N_823);
nor U4422 (N_4422,N_1043,N_1531);
xor U4423 (N_4423,N_1029,N_1307);
xor U4424 (N_4424,N_1032,N_2371);
or U4425 (N_4425,N_1565,N_2034);
nor U4426 (N_4426,N_925,N_1061);
nor U4427 (N_4427,N_1946,N_2063);
nor U4428 (N_4428,N_1610,N_356);
or U4429 (N_4429,N_1301,N_1238);
or U4430 (N_4430,N_431,N_2085);
xor U4431 (N_4431,N_2174,N_235);
and U4432 (N_4432,N_626,N_1234);
or U4433 (N_4433,N_823,N_1958);
and U4434 (N_4434,N_1332,N_1662);
and U4435 (N_4435,N_1436,N_1851);
nand U4436 (N_4436,N_1051,N_1094);
nor U4437 (N_4437,N_2391,N_190);
xor U4438 (N_4438,N_1621,N_377);
and U4439 (N_4439,N_2224,N_248);
nand U4440 (N_4440,N_950,N_532);
or U4441 (N_4441,N_2462,N_2102);
nand U4442 (N_4442,N_554,N_1944);
nor U4443 (N_4443,N_2057,N_296);
nor U4444 (N_4444,N_1450,N_2478);
nand U4445 (N_4445,N_2084,N_1255);
and U4446 (N_4446,N_966,N_1858);
or U4447 (N_4447,N_1020,N_1880);
and U4448 (N_4448,N_1280,N_31);
xnor U4449 (N_4449,N_1804,N_787);
or U4450 (N_4450,N_1010,N_840);
xor U4451 (N_4451,N_423,N_278);
and U4452 (N_4452,N_1193,N_413);
nand U4453 (N_4453,N_634,N_2320);
or U4454 (N_4454,N_368,N_1568);
xor U4455 (N_4455,N_1513,N_1222);
or U4456 (N_4456,N_54,N_2021);
nand U4457 (N_4457,N_44,N_1326);
or U4458 (N_4458,N_970,N_846);
or U4459 (N_4459,N_1240,N_1997);
and U4460 (N_4460,N_993,N_626);
nand U4461 (N_4461,N_199,N_970);
xor U4462 (N_4462,N_494,N_1046);
or U4463 (N_4463,N_1324,N_198);
xor U4464 (N_4464,N_612,N_1186);
nand U4465 (N_4465,N_324,N_2117);
nor U4466 (N_4466,N_684,N_208);
and U4467 (N_4467,N_2164,N_652);
nand U4468 (N_4468,N_1490,N_156);
nor U4469 (N_4469,N_1255,N_1137);
or U4470 (N_4470,N_1515,N_1457);
and U4471 (N_4471,N_1354,N_777);
and U4472 (N_4472,N_661,N_61);
nor U4473 (N_4473,N_765,N_818);
or U4474 (N_4474,N_1726,N_624);
and U4475 (N_4475,N_2209,N_1154);
nor U4476 (N_4476,N_2219,N_1039);
xnor U4477 (N_4477,N_2055,N_413);
nor U4478 (N_4478,N_1202,N_1586);
and U4479 (N_4479,N_207,N_2329);
nand U4480 (N_4480,N_2360,N_1175);
and U4481 (N_4481,N_547,N_894);
and U4482 (N_4482,N_2308,N_2367);
nor U4483 (N_4483,N_2392,N_377);
nor U4484 (N_4484,N_2320,N_2459);
xnor U4485 (N_4485,N_1350,N_844);
nor U4486 (N_4486,N_1838,N_1734);
or U4487 (N_4487,N_1214,N_993);
xnor U4488 (N_4488,N_913,N_1432);
or U4489 (N_4489,N_2044,N_728);
nand U4490 (N_4490,N_2406,N_1951);
or U4491 (N_4491,N_2047,N_1599);
and U4492 (N_4492,N_1856,N_886);
xor U4493 (N_4493,N_1330,N_230);
and U4494 (N_4494,N_689,N_2393);
xnor U4495 (N_4495,N_1068,N_792);
xnor U4496 (N_4496,N_989,N_2289);
nor U4497 (N_4497,N_2463,N_1198);
or U4498 (N_4498,N_280,N_168);
nor U4499 (N_4499,N_1396,N_1614);
and U4500 (N_4500,N_1152,N_711);
and U4501 (N_4501,N_417,N_203);
nor U4502 (N_4502,N_656,N_834);
or U4503 (N_4503,N_2033,N_1102);
and U4504 (N_4504,N_55,N_1174);
and U4505 (N_4505,N_2179,N_580);
nor U4506 (N_4506,N_1252,N_704);
nor U4507 (N_4507,N_1534,N_2210);
nand U4508 (N_4508,N_345,N_1828);
and U4509 (N_4509,N_2068,N_2120);
or U4510 (N_4510,N_1353,N_711);
or U4511 (N_4511,N_1390,N_268);
or U4512 (N_4512,N_2309,N_324);
nor U4513 (N_4513,N_1300,N_1493);
nand U4514 (N_4514,N_2491,N_1124);
or U4515 (N_4515,N_718,N_282);
xnor U4516 (N_4516,N_839,N_112);
nor U4517 (N_4517,N_655,N_2102);
nor U4518 (N_4518,N_205,N_1337);
nor U4519 (N_4519,N_1623,N_623);
nor U4520 (N_4520,N_849,N_2181);
nand U4521 (N_4521,N_1359,N_1909);
and U4522 (N_4522,N_1092,N_2144);
nand U4523 (N_4523,N_1052,N_2354);
xor U4524 (N_4524,N_2137,N_1552);
xor U4525 (N_4525,N_1097,N_864);
nor U4526 (N_4526,N_2139,N_2081);
xnor U4527 (N_4527,N_1472,N_480);
xnor U4528 (N_4528,N_1724,N_1840);
or U4529 (N_4529,N_1707,N_555);
and U4530 (N_4530,N_552,N_1354);
or U4531 (N_4531,N_1352,N_2498);
or U4532 (N_4532,N_1860,N_532);
nor U4533 (N_4533,N_1703,N_1821);
xnor U4534 (N_4534,N_215,N_2178);
nor U4535 (N_4535,N_742,N_507);
nor U4536 (N_4536,N_1365,N_1096);
or U4537 (N_4537,N_584,N_2267);
nor U4538 (N_4538,N_870,N_2257);
nand U4539 (N_4539,N_938,N_2328);
and U4540 (N_4540,N_796,N_1556);
or U4541 (N_4541,N_134,N_1628);
nand U4542 (N_4542,N_2114,N_507);
nor U4543 (N_4543,N_273,N_1764);
nor U4544 (N_4544,N_69,N_1483);
nand U4545 (N_4545,N_1876,N_960);
nand U4546 (N_4546,N_743,N_483);
nand U4547 (N_4547,N_6,N_1523);
and U4548 (N_4548,N_2383,N_1153);
or U4549 (N_4549,N_2012,N_674);
nor U4550 (N_4550,N_371,N_282);
nor U4551 (N_4551,N_639,N_1717);
nor U4552 (N_4552,N_2025,N_810);
nor U4553 (N_4553,N_361,N_1359);
nor U4554 (N_4554,N_2463,N_2195);
or U4555 (N_4555,N_1511,N_710);
or U4556 (N_4556,N_1310,N_1531);
nand U4557 (N_4557,N_1853,N_2309);
nand U4558 (N_4558,N_319,N_1813);
or U4559 (N_4559,N_1691,N_1897);
nor U4560 (N_4560,N_894,N_2125);
xnor U4561 (N_4561,N_1404,N_2430);
xor U4562 (N_4562,N_222,N_1763);
nand U4563 (N_4563,N_727,N_397);
nor U4564 (N_4564,N_2427,N_1998);
xnor U4565 (N_4565,N_1881,N_1082);
or U4566 (N_4566,N_421,N_2439);
or U4567 (N_4567,N_2146,N_1815);
nand U4568 (N_4568,N_201,N_192);
or U4569 (N_4569,N_1634,N_1101);
nor U4570 (N_4570,N_1161,N_1266);
and U4571 (N_4571,N_945,N_1211);
xnor U4572 (N_4572,N_940,N_1052);
nand U4573 (N_4573,N_1372,N_1059);
and U4574 (N_4574,N_278,N_244);
nor U4575 (N_4575,N_2175,N_574);
nand U4576 (N_4576,N_323,N_1523);
and U4577 (N_4577,N_1098,N_18);
and U4578 (N_4578,N_1054,N_1084);
nor U4579 (N_4579,N_1837,N_2275);
xnor U4580 (N_4580,N_2441,N_111);
nand U4581 (N_4581,N_22,N_624);
nor U4582 (N_4582,N_982,N_1597);
nor U4583 (N_4583,N_1884,N_1659);
and U4584 (N_4584,N_1614,N_2035);
xor U4585 (N_4585,N_1923,N_936);
and U4586 (N_4586,N_2328,N_188);
nand U4587 (N_4587,N_568,N_2127);
nand U4588 (N_4588,N_99,N_1721);
xor U4589 (N_4589,N_816,N_1203);
nor U4590 (N_4590,N_1238,N_197);
nand U4591 (N_4591,N_1843,N_428);
nand U4592 (N_4592,N_471,N_1751);
xnor U4593 (N_4593,N_947,N_2442);
nor U4594 (N_4594,N_794,N_2491);
and U4595 (N_4595,N_1529,N_2017);
and U4596 (N_4596,N_577,N_1738);
nand U4597 (N_4597,N_1461,N_137);
and U4598 (N_4598,N_2422,N_547);
nor U4599 (N_4599,N_1262,N_2006);
nor U4600 (N_4600,N_220,N_129);
nand U4601 (N_4601,N_1350,N_1836);
xnor U4602 (N_4602,N_1655,N_803);
xor U4603 (N_4603,N_708,N_1152);
or U4604 (N_4604,N_994,N_339);
and U4605 (N_4605,N_563,N_2217);
and U4606 (N_4606,N_1702,N_458);
nor U4607 (N_4607,N_2187,N_1503);
and U4608 (N_4608,N_944,N_1998);
xor U4609 (N_4609,N_279,N_642);
nand U4610 (N_4610,N_1993,N_1137);
xnor U4611 (N_4611,N_352,N_660);
or U4612 (N_4612,N_1051,N_660);
xor U4613 (N_4613,N_1513,N_2400);
nand U4614 (N_4614,N_841,N_2163);
and U4615 (N_4615,N_1995,N_272);
or U4616 (N_4616,N_459,N_1506);
nand U4617 (N_4617,N_2401,N_1708);
nand U4618 (N_4618,N_129,N_197);
xnor U4619 (N_4619,N_827,N_1502);
nand U4620 (N_4620,N_320,N_1535);
or U4621 (N_4621,N_1447,N_238);
or U4622 (N_4622,N_930,N_1832);
nand U4623 (N_4623,N_1791,N_1094);
and U4624 (N_4624,N_1934,N_865);
or U4625 (N_4625,N_2004,N_2021);
and U4626 (N_4626,N_1755,N_44);
and U4627 (N_4627,N_1700,N_1503);
and U4628 (N_4628,N_1354,N_1424);
xnor U4629 (N_4629,N_2010,N_124);
nor U4630 (N_4630,N_469,N_1942);
or U4631 (N_4631,N_253,N_363);
nor U4632 (N_4632,N_1707,N_2061);
or U4633 (N_4633,N_1313,N_509);
and U4634 (N_4634,N_2038,N_2179);
or U4635 (N_4635,N_647,N_898);
nor U4636 (N_4636,N_208,N_1250);
xnor U4637 (N_4637,N_1260,N_34);
xor U4638 (N_4638,N_1928,N_871);
or U4639 (N_4639,N_2118,N_1336);
and U4640 (N_4640,N_817,N_1242);
and U4641 (N_4641,N_966,N_1867);
and U4642 (N_4642,N_1372,N_1098);
and U4643 (N_4643,N_504,N_842);
and U4644 (N_4644,N_525,N_2183);
nor U4645 (N_4645,N_2281,N_2190);
nor U4646 (N_4646,N_830,N_1895);
nand U4647 (N_4647,N_1425,N_2466);
nand U4648 (N_4648,N_2328,N_836);
or U4649 (N_4649,N_2196,N_599);
nor U4650 (N_4650,N_89,N_1095);
nand U4651 (N_4651,N_291,N_1684);
or U4652 (N_4652,N_1517,N_1688);
xnor U4653 (N_4653,N_307,N_56);
and U4654 (N_4654,N_1830,N_1027);
nand U4655 (N_4655,N_2118,N_735);
nand U4656 (N_4656,N_1720,N_1634);
nand U4657 (N_4657,N_795,N_2394);
xor U4658 (N_4658,N_194,N_1550);
xor U4659 (N_4659,N_550,N_2226);
nor U4660 (N_4660,N_32,N_2040);
nor U4661 (N_4661,N_2177,N_582);
and U4662 (N_4662,N_84,N_431);
xor U4663 (N_4663,N_1830,N_1247);
xnor U4664 (N_4664,N_176,N_313);
nor U4665 (N_4665,N_1670,N_2090);
nor U4666 (N_4666,N_1846,N_1158);
or U4667 (N_4667,N_1161,N_1778);
nand U4668 (N_4668,N_577,N_1246);
and U4669 (N_4669,N_692,N_1732);
or U4670 (N_4670,N_1523,N_577);
nand U4671 (N_4671,N_1637,N_1288);
nand U4672 (N_4672,N_92,N_617);
nand U4673 (N_4673,N_1614,N_1990);
and U4674 (N_4674,N_163,N_1148);
nand U4675 (N_4675,N_1618,N_1005);
xor U4676 (N_4676,N_1884,N_466);
and U4677 (N_4677,N_178,N_328);
nand U4678 (N_4678,N_2058,N_1160);
and U4679 (N_4679,N_1795,N_2156);
nor U4680 (N_4680,N_1402,N_106);
or U4681 (N_4681,N_461,N_774);
nand U4682 (N_4682,N_2393,N_931);
xor U4683 (N_4683,N_711,N_1515);
xnor U4684 (N_4684,N_461,N_1851);
or U4685 (N_4685,N_2033,N_2468);
or U4686 (N_4686,N_1433,N_1154);
nand U4687 (N_4687,N_334,N_1699);
nor U4688 (N_4688,N_960,N_733);
nor U4689 (N_4689,N_931,N_1892);
nand U4690 (N_4690,N_843,N_2074);
or U4691 (N_4691,N_1302,N_390);
xor U4692 (N_4692,N_1364,N_1355);
nor U4693 (N_4693,N_1173,N_237);
and U4694 (N_4694,N_1958,N_548);
and U4695 (N_4695,N_1442,N_477);
xnor U4696 (N_4696,N_1566,N_1543);
nor U4697 (N_4697,N_731,N_292);
and U4698 (N_4698,N_1120,N_950);
xor U4699 (N_4699,N_975,N_1186);
and U4700 (N_4700,N_1434,N_2034);
nor U4701 (N_4701,N_1513,N_1096);
or U4702 (N_4702,N_1803,N_804);
xor U4703 (N_4703,N_1155,N_1797);
or U4704 (N_4704,N_2186,N_613);
nor U4705 (N_4705,N_34,N_2036);
and U4706 (N_4706,N_2406,N_1607);
or U4707 (N_4707,N_1687,N_1155);
nand U4708 (N_4708,N_649,N_315);
nor U4709 (N_4709,N_72,N_682);
and U4710 (N_4710,N_2112,N_1868);
nand U4711 (N_4711,N_1007,N_2013);
or U4712 (N_4712,N_1895,N_592);
nor U4713 (N_4713,N_1747,N_1376);
nor U4714 (N_4714,N_1372,N_884);
and U4715 (N_4715,N_2467,N_91);
nand U4716 (N_4716,N_1952,N_2483);
and U4717 (N_4717,N_1974,N_834);
nand U4718 (N_4718,N_743,N_845);
and U4719 (N_4719,N_798,N_1097);
and U4720 (N_4720,N_1961,N_2472);
nand U4721 (N_4721,N_2354,N_1745);
nand U4722 (N_4722,N_1765,N_1269);
xor U4723 (N_4723,N_63,N_1556);
and U4724 (N_4724,N_2000,N_1861);
xor U4725 (N_4725,N_1964,N_152);
xor U4726 (N_4726,N_1394,N_56);
and U4727 (N_4727,N_2295,N_372);
and U4728 (N_4728,N_437,N_2286);
or U4729 (N_4729,N_48,N_2234);
nor U4730 (N_4730,N_255,N_529);
xor U4731 (N_4731,N_594,N_2337);
nor U4732 (N_4732,N_1902,N_92);
and U4733 (N_4733,N_2154,N_892);
or U4734 (N_4734,N_1870,N_2431);
nor U4735 (N_4735,N_1516,N_1280);
and U4736 (N_4736,N_1460,N_2143);
or U4737 (N_4737,N_1969,N_1119);
nor U4738 (N_4738,N_1755,N_403);
or U4739 (N_4739,N_2313,N_744);
nor U4740 (N_4740,N_2408,N_1337);
xor U4741 (N_4741,N_1977,N_6);
nor U4742 (N_4742,N_112,N_187);
nand U4743 (N_4743,N_511,N_684);
or U4744 (N_4744,N_1978,N_2086);
and U4745 (N_4745,N_752,N_83);
and U4746 (N_4746,N_649,N_1418);
and U4747 (N_4747,N_2184,N_1904);
nand U4748 (N_4748,N_524,N_1422);
nand U4749 (N_4749,N_436,N_1799);
nand U4750 (N_4750,N_971,N_713);
nor U4751 (N_4751,N_1284,N_1736);
xor U4752 (N_4752,N_1162,N_744);
nand U4753 (N_4753,N_537,N_2069);
xnor U4754 (N_4754,N_1752,N_1002);
nand U4755 (N_4755,N_828,N_1816);
and U4756 (N_4756,N_147,N_1475);
xor U4757 (N_4757,N_2000,N_1731);
and U4758 (N_4758,N_370,N_380);
xnor U4759 (N_4759,N_2251,N_1847);
nand U4760 (N_4760,N_226,N_2232);
and U4761 (N_4761,N_1156,N_1544);
xnor U4762 (N_4762,N_218,N_194);
xor U4763 (N_4763,N_1689,N_1156);
nor U4764 (N_4764,N_1982,N_1942);
nand U4765 (N_4765,N_1086,N_526);
and U4766 (N_4766,N_1865,N_579);
nor U4767 (N_4767,N_227,N_281);
or U4768 (N_4768,N_1885,N_960);
nand U4769 (N_4769,N_610,N_1570);
nand U4770 (N_4770,N_2230,N_1833);
xor U4771 (N_4771,N_999,N_1015);
or U4772 (N_4772,N_2244,N_1436);
or U4773 (N_4773,N_1942,N_120);
nand U4774 (N_4774,N_644,N_502);
and U4775 (N_4775,N_368,N_789);
and U4776 (N_4776,N_2407,N_2387);
xnor U4777 (N_4777,N_421,N_1749);
or U4778 (N_4778,N_1008,N_965);
xor U4779 (N_4779,N_537,N_959);
and U4780 (N_4780,N_1573,N_1493);
and U4781 (N_4781,N_339,N_479);
nand U4782 (N_4782,N_577,N_2405);
or U4783 (N_4783,N_1972,N_1744);
and U4784 (N_4784,N_518,N_1425);
nand U4785 (N_4785,N_608,N_1128);
and U4786 (N_4786,N_657,N_1210);
xnor U4787 (N_4787,N_2238,N_747);
xnor U4788 (N_4788,N_1863,N_375);
xnor U4789 (N_4789,N_2369,N_1803);
xor U4790 (N_4790,N_1007,N_229);
nor U4791 (N_4791,N_2164,N_475);
xor U4792 (N_4792,N_482,N_1904);
nor U4793 (N_4793,N_431,N_1093);
xnor U4794 (N_4794,N_2064,N_160);
or U4795 (N_4795,N_1181,N_1793);
xnor U4796 (N_4796,N_327,N_68);
nand U4797 (N_4797,N_872,N_2484);
nand U4798 (N_4798,N_2382,N_387);
nor U4799 (N_4799,N_2412,N_859);
nand U4800 (N_4800,N_358,N_105);
nor U4801 (N_4801,N_1739,N_1980);
or U4802 (N_4802,N_742,N_2396);
and U4803 (N_4803,N_2491,N_1759);
nand U4804 (N_4804,N_2462,N_1523);
nor U4805 (N_4805,N_1143,N_556);
nand U4806 (N_4806,N_2258,N_1159);
nor U4807 (N_4807,N_2029,N_354);
and U4808 (N_4808,N_67,N_387);
xor U4809 (N_4809,N_300,N_1205);
nand U4810 (N_4810,N_1788,N_2205);
or U4811 (N_4811,N_1417,N_634);
xor U4812 (N_4812,N_2273,N_1231);
or U4813 (N_4813,N_1485,N_1665);
nand U4814 (N_4814,N_2192,N_608);
nor U4815 (N_4815,N_74,N_2269);
or U4816 (N_4816,N_333,N_2478);
nor U4817 (N_4817,N_2077,N_2280);
nand U4818 (N_4818,N_2,N_2171);
xor U4819 (N_4819,N_2472,N_709);
xnor U4820 (N_4820,N_93,N_61);
or U4821 (N_4821,N_2362,N_331);
or U4822 (N_4822,N_448,N_550);
nand U4823 (N_4823,N_125,N_677);
and U4824 (N_4824,N_1157,N_1572);
and U4825 (N_4825,N_309,N_2223);
nand U4826 (N_4826,N_2148,N_2149);
xor U4827 (N_4827,N_944,N_1701);
nand U4828 (N_4828,N_814,N_721);
nor U4829 (N_4829,N_1383,N_725);
or U4830 (N_4830,N_259,N_1236);
xor U4831 (N_4831,N_1520,N_961);
nand U4832 (N_4832,N_1555,N_1683);
or U4833 (N_4833,N_1470,N_2281);
xnor U4834 (N_4834,N_866,N_2160);
or U4835 (N_4835,N_545,N_2429);
and U4836 (N_4836,N_1402,N_2354);
xnor U4837 (N_4837,N_540,N_818);
xnor U4838 (N_4838,N_552,N_602);
xnor U4839 (N_4839,N_1825,N_1597);
and U4840 (N_4840,N_367,N_2182);
and U4841 (N_4841,N_978,N_443);
xnor U4842 (N_4842,N_119,N_33);
nor U4843 (N_4843,N_2256,N_1980);
nor U4844 (N_4844,N_598,N_2074);
and U4845 (N_4845,N_1124,N_757);
nand U4846 (N_4846,N_302,N_2383);
xor U4847 (N_4847,N_1927,N_752);
xnor U4848 (N_4848,N_1332,N_1999);
xor U4849 (N_4849,N_1819,N_394);
xor U4850 (N_4850,N_240,N_1709);
xnor U4851 (N_4851,N_1093,N_1931);
nor U4852 (N_4852,N_1519,N_1107);
and U4853 (N_4853,N_917,N_904);
or U4854 (N_4854,N_1697,N_351);
nand U4855 (N_4855,N_2477,N_2051);
and U4856 (N_4856,N_1630,N_1222);
nand U4857 (N_4857,N_1958,N_2281);
xor U4858 (N_4858,N_2022,N_2016);
or U4859 (N_4859,N_1996,N_791);
nand U4860 (N_4860,N_1471,N_2229);
nor U4861 (N_4861,N_300,N_2460);
nor U4862 (N_4862,N_1641,N_1221);
nor U4863 (N_4863,N_113,N_809);
xor U4864 (N_4864,N_455,N_2033);
nor U4865 (N_4865,N_1925,N_1704);
or U4866 (N_4866,N_1713,N_380);
or U4867 (N_4867,N_1813,N_1196);
xnor U4868 (N_4868,N_1035,N_1514);
or U4869 (N_4869,N_2094,N_2239);
nor U4870 (N_4870,N_1939,N_1175);
nand U4871 (N_4871,N_716,N_2088);
nand U4872 (N_4872,N_44,N_2448);
nand U4873 (N_4873,N_2035,N_2014);
and U4874 (N_4874,N_1444,N_1417);
nand U4875 (N_4875,N_2432,N_1294);
or U4876 (N_4876,N_1966,N_1313);
nor U4877 (N_4877,N_1408,N_1836);
nor U4878 (N_4878,N_1444,N_1655);
nand U4879 (N_4879,N_464,N_1583);
xor U4880 (N_4880,N_61,N_1865);
and U4881 (N_4881,N_967,N_59);
or U4882 (N_4882,N_2188,N_1160);
or U4883 (N_4883,N_571,N_917);
and U4884 (N_4884,N_1476,N_1420);
or U4885 (N_4885,N_375,N_1564);
nand U4886 (N_4886,N_2020,N_1834);
nor U4887 (N_4887,N_653,N_1562);
and U4888 (N_4888,N_503,N_329);
nand U4889 (N_4889,N_1796,N_1830);
nand U4890 (N_4890,N_987,N_1200);
xnor U4891 (N_4891,N_1430,N_1717);
nor U4892 (N_4892,N_1928,N_914);
nor U4893 (N_4893,N_212,N_12);
or U4894 (N_4894,N_158,N_2268);
nand U4895 (N_4895,N_284,N_673);
nor U4896 (N_4896,N_1694,N_1888);
nor U4897 (N_4897,N_2421,N_1414);
nand U4898 (N_4898,N_2329,N_1787);
nor U4899 (N_4899,N_771,N_2383);
nor U4900 (N_4900,N_2106,N_252);
nor U4901 (N_4901,N_1475,N_1962);
and U4902 (N_4902,N_719,N_1640);
nand U4903 (N_4903,N_1315,N_2275);
or U4904 (N_4904,N_341,N_1280);
or U4905 (N_4905,N_298,N_1871);
nor U4906 (N_4906,N_1611,N_150);
or U4907 (N_4907,N_1085,N_1188);
nor U4908 (N_4908,N_1867,N_1343);
nand U4909 (N_4909,N_1165,N_416);
and U4910 (N_4910,N_997,N_1463);
nor U4911 (N_4911,N_364,N_468);
and U4912 (N_4912,N_1109,N_554);
or U4913 (N_4913,N_1695,N_1918);
nor U4914 (N_4914,N_1414,N_2136);
nand U4915 (N_4915,N_439,N_1833);
xnor U4916 (N_4916,N_1120,N_498);
and U4917 (N_4917,N_1085,N_901);
or U4918 (N_4918,N_1900,N_2167);
or U4919 (N_4919,N_1894,N_535);
or U4920 (N_4920,N_2359,N_2072);
or U4921 (N_4921,N_591,N_2268);
or U4922 (N_4922,N_2470,N_359);
nand U4923 (N_4923,N_361,N_1558);
nand U4924 (N_4924,N_763,N_1491);
nor U4925 (N_4925,N_1468,N_1673);
and U4926 (N_4926,N_1295,N_327);
nor U4927 (N_4927,N_893,N_1055);
and U4928 (N_4928,N_1224,N_1070);
nor U4929 (N_4929,N_897,N_1999);
xnor U4930 (N_4930,N_346,N_582);
nor U4931 (N_4931,N_48,N_1649);
nor U4932 (N_4932,N_676,N_651);
or U4933 (N_4933,N_576,N_1915);
nor U4934 (N_4934,N_1905,N_321);
and U4935 (N_4935,N_582,N_1074);
xor U4936 (N_4936,N_2498,N_1548);
and U4937 (N_4937,N_1173,N_504);
xnor U4938 (N_4938,N_301,N_2134);
nand U4939 (N_4939,N_260,N_48);
nand U4940 (N_4940,N_794,N_2290);
and U4941 (N_4941,N_2140,N_860);
nor U4942 (N_4942,N_1971,N_2230);
or U4943 (N_4943,N_1412,N_1312);
or U4944 (N_4944,N_1175,N_685);
xor U4945 (N_4945,N_429,N_698);
xnor U4946 (N_4946,N_644,N_1844);
or U4947 (N_4947,N_1593,N_1493);
and U4948 (N_4948,N_2308,N_38);
and U4949 (N_4949,N_2494,N_77);
nor U4950 (N_4950,N_2232,N_569);
or U4951 (N_4951,N_1155,N_661);
nand U4952 (N_4952,N_1061,N_1737);
nor U4953 (N_4953,N_2280,N_322);
nor U4954 (N_4954,N_954,N_177);
nand U4955 (N_4955,N_2309,N_835);
and U4956 (N_4956,N_2151,N_867);
nand U4957 (N_4957,N_1582,N_2414);
nor U4958 (N_4958,N_582,N_1360);
xor U4959 (N_4959,N_1427,N_1299);
nor U4960 (N_4960,N_381,N_1405);
nor U4961 (N_4961,N_2130,N_301);
xnor U4962 (N_4962,N_2376,N_1958);
xnor U4963 (N_4963,N_619,N_1103);
xnor U4964 (N_4964,N_1684,N_172);
nand U4965 (N_4965,N_2478,N_153);
nor U4966 (N_4966,N_2029,N_2080);
or U4967 (N_4967,N_936,N_633);
or U4968 (N_4968,N_101,N_1609);
nand U4969 (N_4969,N_1934,N_1863);
nand U4970 (N_4970,N_1803,N_796);
nor U4971 (N_4971,N_2458,N_561);
or U4972 (N_4972,N_214,N_681);
or U4973 (N_4973,N_1624,N_2122);
nor U4974 (N_4974,N_1572,N_1354);
nand U4975 (N_4975,N_1597,N_614);
and U4976 (N_4976,N_2107,N_1724);
nand U4977 (N_4977,N_1347,N_629);
and U4978 (N_4978,N_2293,N_1041);
or U4979 (N_4979,N_1132,N_1255);
and U4980 (N_4980,N_780,N_272);
xor U4981 (N_4981,N_2236,N_1690);
nor U4982 (N_4982,N_856,N_898);
nand U4983 (N_4983,N_1215,N_1024);
or U4984 (N_4984,N_1200,N_896);
nand U4985 (N_4985,N_1305,N_1105);
xor U4986 (N_4986,N_150,N_1215);
or U4987 (N_4987,N_365,N_1644);
nand U4988 (N_4988,N_1147,N_2097);
xor U4989 (N_4989,N_1016,N_406);
and U4990 (N_4990,N_823,N_664);
xor U4991 (N_4991,N_331,N_73);
nor U4992 (N_4992,N_295,N_1032);
xnor U4993 (N_4993,N_2209,N_1383);
nor U4994 (N_4994,N_1744,N_2255);
nand U4995 (N_4995,N_455,N_1023);
and U4996 (N_4996,N_1264,N_1124);
or U4997 (N_4997,N_227,N_1798);
or U4998 (N_4998,N_2155,N_142);
nor U4999 (N_4999,N_2116,N_87);
nand U5000 (N_5000,N_4378,N_3177);
nor U5001 (N_5001,N_4044,N_3685);
nand U5002 (N_5002,N_4879,N_3100);
xnor U5003 (N_5003,N_4135,N_2754);
xor U5004 (N_5004,N_4920,N_3080);
xor U5005 (N_5005,N_4354,N_3014);
or U5006 (N_5006,N_2949,N_4919);
xor U5007 (N_5007,N_3839,N_3991);
nand U5008 (N_5008,N_3989,N_2525);
or U5009 (N_5009,N_3360,N_4750);
nor U5010 (N_5010,N_3190,N_3883);
nor U5011 (N_5011,N_3972,N_3879);
or U5012 (N_5012,N_2660,N_2783);
nand U5013 (N_5013,N_3663,N_4914);
nand U5014 (N_5014,N_4438,N_3760);
and U5015 (N_5015,N_2786,N_3001);
xnor U5016 (N_5016,N_2957,N_2685);
and U5017 (N_5017,N_3763,N_3158);
and U5018 (N_5018,N_4204,N_3726);
nand U5019 (N_5019,N_3370,N_2803);
xnor U5020 (N_5020,N_2999,N_4238);
and U5021 (N_5021,N_3417,N_3724);
nand U5022 (N_5022,N_2636,N_4801);
or U5023 (N_5023,N_3865,N_3297);
and U5024 (N_5024,N_4398,N_2751);
xnor U5025 (N_5025,N_4669,N_3157);
nand U5026 (N_5026,N_4065,N_4967);
and U5027 (N_5027,N_4397,N_4935);
nor U5028 (N_5028,N_3935,N_3076);
nand U5029 (N_5029,N_3302,N_4784);
and U5030 (N_5030,N_3867,N_3735);
and U5031 (N_5031,N_4089,N_3885);
or U5032 (N_5032,N_3727,N_3475);
and U5033 (N_5033,N_3889,N_4294);
or U5034 (N_5034,N_3494,N_3606);
and U5035 (N_5035,N_3139,N_4251);
xnor U5036 (N_5036,N_4757,N_4627);
nand U5037 (N_5037,N_3791,N_2665);
nor U5038 (N_5038,N_2694,N_2895);
xnor U5039 (N_5039,N_2628,N_4871);
xnor U5040 (N_5040,N_4979,N_3456);
xor U5041 (N_5041,N_3778,N_4907);
and U5042 (N_5042,N_4806,N_4410);
or U5043 (N_5043,N_4708,N_3504);
nor U5044 (N_5044,N_4675,N_2847);
or U5045 (N_5045,N_2517,N_4477);
nor U5046 (N_5046,N_4852,N_3786);
xnor U5047 (N_5047,N_3671,N_3143);
nor U5048 (N_5048,N_2811,N_3643);
nor U5049 (N_5049,N_2523,N_2977);
and U5050 (N_5050,N_4745,N_2789);
and U5051 (N_5051,N_4105,N_3353);
or U5052 (N_5052,N_3628,N_4250);
nand U5053 (N_5053,N_3955,N_3783);
xnor U5054 (N_5054,N_3126,N_3399);
nand U5055 (N_5055,N_4771,N_3924);
or U5056 (N_5056,N_4314,N_4962);
nand U5057 (N_5057,N_2520,N_4954);
nor U5058 (N_5058,N_4860,N_3197);
xor U5059 (N_5059,N_3163,N_2651);
or U5060 (N_5060,N_4830,N_4267);
xor U5061 (N_5061,N_4502,N_3765);
nor U5062 (N_5062,N_4787,N_4372);
or U5063 (N_5063,N_4448,N_4566);
xor U5064 (N_5064,N_2527,N_3669);
nor U5065 (N_5065,N_4318,N_3344);
nand U5066 (N_5066,N_2509,N_3994);
xor U5067 (N_5067,N_3249,N_4988);
nand U5068 (N_5068,N_4814,N_4032);
and U5069 (N_5069,N_4349,N_2863);
or U5070 (N_5070,N_4471,N_2878);
nor U5071 (N_5071,N_3603,N_3776);
nor U5072 (N_5072,N_2571,N_4129);
nor U5073 (N_5073,N_2641,N_4336);
and U5074 (N_5074,N_4703,N_4592);
nor U5075 (N_5075,N_3092,N_3950);
nor U5076 (N_5076,N_4216,N_3926);
and U5077 (N_5077,N_3292,N_4835);
nand U5078 (N_5078,N_3425,N_2701);
nor U5079 (N_5079,N_3421,N_4513);
xor U5080 (N_5080,N_4437,N_4021);
nand U5081 (N_5081,N_4290,N_4391);
nor U5082 (N_5082,N_4208,N_3293);
or U5083 (N_5083,N_3537,N_3945);
or U5084 (N_5084,N_2960,N_3079);
and U5085 (N_5085,N_4727,N_2876);
nor U5086 (N_5086,N_4951,N_2541);
nand U5087 (N_5087,N_3097,N_2668);
or U5088 (N_5088,N_3409,N_2968);
nor U5089 (N_5089,N_3944,N_3993);
nand U5090 (N_5090,N_4918,N_4087);
and U5091 (N_5091,N_3075,N_2779);
nor U5092 (N_5092,N_3265,N_2692);
xnor U5093 (N_5093,N_4066,N_3465);
nor U5094 (N_5094,N_3119,N_3648);
xor U5095 (N_5095,N_3961,N_4156);
nand U5096 (N_5096,N_4057,N_4371);
nand U5097 (N_5097,N_3308,N_4434);
and U5098 (N_5098,N_3857,N_3179);
nor U5099 (N_5099,N_4800,N_3151);
and U5100 (N_5100,N_3452,N_2686);
and U5101 (N_5101,N_4759,N_3689);
or U5102 (N_5102,N_3440,N_3533);
or U5103 (N_5103,N_3762,N_3929);
nand U5104 (N_5104,N_3911,N_3275);
nor U5105 (N_5105,N_3335,N_4744);
nand U5106 (N_5106,N_2870,N_4522);
nor U5107 (N_5107,N_3424,N_4539);
nand U5108 (N_5108,N_3806,N_3952);
nor U5109 (N_5109,N_4584,N_2965);
and U5110 (N_5110,N_4597,N_2549);
xor U5111 (N_5111,N_3212,N_3515);
or U5112 (N_5112,N_2943,N_3199);
and U5113 (N_5113,N_2621,N_4261);
nand U5114 (N_5114,N_3410,N_4339);
or U5115 (N_5115,N_4262,N_4640);
xnor U5116 (N_5116,N_2623,N_4224);
nand U5117 (N_5117,N_4258,N_3154);
and U5118 (N_5118,N_2890,N_2880);
or U5119 (N_5119,N_3394,N_2820);
or U5120 (N_5120,N_4666,N_4024);
nor U5121 (N_5121,N_2936,N_4244);
and U5122 (N_5122,N_4141,N_4520);
nor U5123 (N_5123,N_2563,N_3621);
or U5124 (N_5124,N_4850,N_4384);
and U5125 (N_5125,N_4615,N_2840);
xor U5126 (N_5126,N_4151,N_3650);
nand U5127 (N_5127,N_3875,N_3049);
xnor U5128 (N_5128,N_3884,N_4595);
and U5129 (N_5129,N_3542,N_4042);
or U5130 (N_5130,N_4439,N_3320);
and U5131 (N_5131,N_4181,N_3196);
and U5132 (N_5132,N_2532,N_3136);
nor U5133 (N_5133,N_2742,N_3958);
nor U5134 (N_5134,N_3240,N_4748);
and U5135 (N_5135,N_4512,N_4004);
and U5136 (N_5136,N_4901,N_3832);
or U5137 (N_5137,N_3539,N_4281);
or U5138 (N_5138,N_3691,N_4858);
xnor U5139 (N_5139,N_4588,N_3165);
or U5140 (N_5140,N_3607,N_4408);
nor U5141 (N_5141,N_2625,N_3705);
xnor U5142 (N_5142,N_4574,N_3990);
nand U5143 (N_5143,N_4223,N_2547);
or U5144 (N_5144,N_3433,N_3811);
nor U5145 (N_5145,N_4500,N_4980);
or U5146 (N_5146,N_3622,N_4711);
nor U5147 (N_5147,N_4594,N_4557);
nor U5148 (N_5148,N_4280,N_3849);
nand U5149 (N_5149,N_3728,N_2784);
nor U5150 (N_5150,N_4401,N_3784);
and U5151 (N_5151,N_4655,N_3574);
or U5152 (N_5152,N_3676,N_4106);
nor U5153 (N_5153,N_3432,N_3850);
and U5154 (N_5154,N_4934,N_3661);
and U5155 (N_5155,N_3534,N_3796);
nor U5156 (N_5156,N_2741,N_4684);
nand U5157 (N_5157,N_2806,N_3348);
xnor U5158 (N_5158,N_3658,N_2782);
xor U5159 (N_5159,N_4804,N_4517);
nand U5160 (N_5160,N_4012,N_3629);
and U5161 (N_5161,N_3655,N_3900);
or U5162 (N_5162,N_3920,N_3764);
xnor U5163 (N_5163,N_2848,N_2788);
nor U5164 (N_5164,N_3930,N_2639);
nor U5165 (N_5165,N_3323,N_3808);
xor U5166 (N_5166,N_4508,N_2767);
nor U5167 (N_5167,N_3802,N_4328);
and U5168 (N_5168,N_4710,N_4414);
xnor U5169 (N_5169,N_4900,N_3211);
xnor U5170 (N_5170,N_3054,N_3052);
and U5171 (N_5171,N_4386,N_3836);
nand U5172 (N_5172,N_3449,N_4734);
and U5173 (N_5173,N_3769,N_4310);
xnor U5174 (N_5174,N_2849,N_3687);
or U5175 (N_5175,N_4237,N_4605);
nor U5176 (N_5176,N_4768,N_4256);
nor U5177 (N_5177,N_3583,N_3656);
and U5178 (N_5178,N_2909,N_2629);
nor U5179 (N_5179,N_3375,N_4017);
and U5180 (N_5180,N_2927,N_4200);
xor U5181 (N_5181,N_2917,N_4071);
and U5182 (N_5182,N_4178,N_2898);
xor U5183 (N_5183,N_4957,N_4060);
and U5184 (N_5184,N_3463,N_4474);
nor U5185 (N_5185,N_4506,N_2940);
or U5186 (N_5186,N_3641,N_4287);
nor U5187 (N_5187,N_3005,N_4325);
nand U5188 (N_5188,N_2959,N_2902);
and U5189 (N_5189,N_3734,N_2558);
nor U5190 (N_5190,N_4777,N_2934);
nor U5191 (N_5191,N_4926,N_4149);
and U5192 (N_5192,N_4000,N_4046);
or U5193 (N_5193,N_3692,N_3238);
or U5194 (N_5194,N_4567,N_2687);
nor U5195 (N_5195,N_3332,N_4102);
nand U5196 (N_5196,N_3766,N_2944);
or U5197 (N_5197,N_3965,N_2883);
nand U5198 (N_5198,N_2529,N_3224);
xor U5199 (N_5199,N_3488,N_4035);
or U5200 (N_5200,N_4947,N_3619);
nor U5201 (N_5201,N_2746,N_2906);
nand U5202 (N_5202,N_4248,N_3416);
or U5203 (N_5203,N_4466,N_2618);
nand U5204 (N_5204,N_4998,N_3572);
and U5205 (N_5205,N_4356,N_2683);
nor U5206 (N_5206,N_4778,N_4292);
nand U5207 (N_5207,N_3191,N_4355);
and U5208 (N_5208,N_4515,N_3833);
and U5209 (N_5209,N_4240,N_3194);
nand U5210 (N_5210,N_3258,N_2877);
or U5211 (N_5211,N_2502,N_4387);
xnor U5212 (N_5212,N_4626,N_4765);
nor U5213 (N_5213,N_2827,N_2635);
and U5214 (N_5214,N_3273,N_4815);
and U5215 (N_5215,N_4925,N_4116);
nand U5216 (N_5216,N_3072,N_3142);
or U5217 (N_5217,N_2729,N_4169);
nand U5218 (N_5218,N_2607,N_2785);
xnor U5219 (N_5219,N_4819,N_3468);
nand U5220 (N_5220,N_3166,N_3963);
nor U5221 (N_5221,N_3343,N_2904);
and U5222 (N_5222,N_2610,N_3322);
xor U5223 (N_5223,N_4054,N_2673);
nor U5224 (N_5224,N_3493,N_3215);
xor U5225 (N_5225,N_3566,N_4442);
nor U5226 (N_5226,N_3120,N_3408);
or U5227 (N_5227,N_2775,N_3252);
and U5228 (N_5228,N_3248,N_4630);
nand U5229 (N_5229,N_4910,N_2584);
and U5230 (N_5230,N_4561,N_3666);
nor U5231 (N_5231,N_2736,N_4342);
xor U5232 (N_5232,N_3230,N_2723);
nor U5233 (N_5233,N_3761,N_4721);
nand U5234 (N_5234,N_4211,N_2631);
nand U5235 (N_5235,N_3321,N_2822);
nor U5236 (N_5236,N_3614,N_3437);
xnor U5237 (N_5237,N_4888,N_2914);
nand U5238 (N_5238,N_3774,N_3315);
and U5239 (N_5239,N_2583,N_3266);
nor U5240 (N_5240,N_2855,N_4521);
and U5241 (N_5241,N_3507,N_3086);
or U5242 (N_5242,N_2908,N_2556);
nand U5243 (N_5243,N_4959,N_3118);
or U5244 (N_5244,N_2738,N_3413);
nor U5245 (N_5245,N_4480,N_3514);
or U5246 (N_5246,N_4961,N_2709);
and U5247 (N_5247,N_2962,N_4505);
or U5248 (N_5248,N_2708,N_3999);
or U5249 (N_5249,N_2648,N_3890);
nand U5250 (N_5250,N_2797,N_3388);
nand U5251 (N_5251,N_3933,N_4831);
nand U5252 (N_5252,N_4866,N_2928);
or U5253 (N_5253,N_3182,N_3277);
nand U5254 (N_5254,N_4284,N_4572);
xnor U5255 (N_5255,N_2695,N_3284);
xor U5256 (N_5256,N_4656,N_2702);
and U5257 (N_5257,N_2579,N_4864);
nor U5258 (N_5258,N_3278,N_4589);
nor U5259 (N_5259,N_3474,N_4764);
or U5260 (N_5260,N_4533,N_4964);
and U5261 (N_5261,N_4317,N_2989);
or U5262 (N_5262,N_4324,N_2666);
xnor U5263 (N_5263,N_3088,N_4337);
or U5264 (N_5264,N_3376,N_3380);
xnor U5265 (N_5265,N_3827,N_3596);
nor U5266 (N_5266,N_4406,N_4345);
or U5267 (N_5267,N_3720,N_3820);
nor U5268 (N_5268,N_2537,N_2518);
nor U5269 (N_5269,N_4992,N_3519);
xor U5270 (N_5270,N_3812,N_3960);
nand U5271 (N_5271,N_4295,N_4699);
and U5272 (N_5272,N_3536,N_2511);
nand U5273 (N_5273,N_4917,N_4086);
nand U5274 (N_5274,N_4430,N_4111);
nor U5275 (N_5275,N_2812,N_3729);
and U5276 (N_5276,N_4476,N_3704);
nor U5277 (N_5277,N_3736,N_3527);
and U5278 (N_5278,N_3254,N_3132);
nor U5279 (N_5279,N_3912,N_3752);
nand U5280 (N_5280,N_4099,N_4068);
xnor U5281 (N_5281,N_3919,N_2577);
nor U5282 (N_5282,N_4762,N_3223);
nand U5283 (N_5283,N_3318,N_4887);
nor U5284 (N_5284,N_4293,N_4671);
or U5285 (N_5285,N_4174,N_3013);
and U5286 (N_5286,N_4763,N_2544);
xor U5287 (N_5287,N_3744,N_2717);
nor U5288 (N_5288,N_3947,N_4642);
nand U5289 (N_5289,N_3552,N_3684);
xnor U5290 (N_5290,N_4229,N_4658);
and U5291 (N_5291,N_4327,N_4045);
xnor U5292 (N_5292,N_3932,N_3516);
nand U5293 (N_5293,N_4534,N_4117);
xnor U5294 (N_5294,N_2550,N_4837);
nor U5295 (N_5295,N_4786,N_2769);
nand U5296 (N_5296,N_3567,N_4997);
and U5297 (N_5297,N_4591,N_3170);
nand U5298 (N_5298,N_4755,N_3931);
or U5299 (N_5299,N_2513,N_2508);
and U5300 (N_5300,N_2690,N_4526);
nor U5301 (N_5301,N_2516,N_2733);
nand U5302 (N_5302,N_4977,N_3334);
and U5303 (N_5303,N_4796,N_3585);
nor U5304 (N_5304,N_4373,N_3276);
nor U5305 (N_5305,N_3634,N_3372);
nand U5306 (N_5306,N_3698,N_4029);
nor U5307 (N_5307,N_4563,N_4532);
and U5308 (N_5308,N_3039,N_4118);
xnor U5309 (N_5309,N_3665,N_4633);
nand U5310 (N_5310,N_2752,N_3768);
or U5311 (N_5311,N_3202,N_2734);
and U5312 (N_5312,N_4014,N_3221);
xnor U5313 (N_5313,N_4230,N_3773);
nand U5314 (N_5314,N_2562,N_2698);
or U5315 (N_5315,N_3460,N_4537);
nor U5316 (N_5316,N_4958,N_4289);
nor U5317 (N_5317,N_3209,N_3184);
nor U5318 (N_5318,N_4899,N_3792);
or U5319 (N_5319,N_2875,N_4928);
or U5320 (N_5320,N_2582,N_4531);
and U5321 (N_5321,N_2930,N_2858);
and U5322 (N_5322,N_4485,N_4629);
xnor U5323 (N_5323,N_4164,N_3181);
and U5324 (N_5324,N_4080,N_4838);
nor U5325 (N_5325,N_3256,N_4746);
xor U5326 (N_5326,N_3436,N_2640);
and U5327 (N_5327,N_4647,N_4482);
nor U5328 (N_5328,N_3551,N_3490);
or U5329 (N_5329,N_2826,N_3451);
nor U5330 (N_5330,N_3770,N_4722);
nand U5331 (N_5331,N_3909,N_3847);
xor U5332 (N_5332,N_3844,N_3015);
xnor U5333 (N_5333,N_4535,N_2897);
nand U5334 (N_5334,N_2554,N_4090);
xor U5335 (N_5335,N_3070,N_2703);
nor U5336 (N_5336,N_4064,N_4217);
and U5337 (N_5337,N_3498,N_4509);
and U5338 (N_5338,N_4028,N_2800);
xnor U5339 (N_5339,N_2545,N_4756);
nor U5340 (N_5340,N_2590,N_4776);
or U5341 (N_5341,N_3759,N_3414);
nand U5342 (N_5342,N_2663,N_2990);
and U5343 (N_5343,N_4559,N_4375);
and U5344 (N_5344,N_3222,N_4683);
and U5345 (N_5345,N_3908,N_4396);
nor U5346 (N_5346,N_4486,N_3781);
xnor U5347 (N_5347,N_3134,N_4933);
xnor U5348 (N_5348,N_3591,N_3346);
xor U5349 (N_5349,N_2543,N_4225);
nand U5350 (N_5350,N_3733,N_4491);
nor U5351 (N_5351,N_3649,N_2514);
and U5352 (N_5352,N_2903,N_4754);
xnor U5353 (N_5353,N_4855,N_3986);
xor U5354 (N_5354,N_3180,N_3447);
nor U5355 (N_5355,N_4079,N_3294);
or U5356 (N_5356,N_3382,N_3517);
xor U5357 (N_5357,N_4740,N_3330);
xnor U5358 (N_5358,N_4076,N_4276);
or U5359 (N_5359,N_3810,N_4596);
xnor U5360 (N_5360,N_4826,N_4555);
and U5361 (N_5361,N_3793,N_3192);
or U5362 (N_5362,N_4395,N_4874);
nor U5363 (N_5363,N_3043,N_3189);
or U5364 (N_5364,N_2770,N_3943);
nand U5365 (N_5365,N_4185,N_4797);
nand U5366 (N_5366,N_3064,N_3444);
nor U5367 (N_5367,N_4377,N_2595);
nor U5368 (N_5368,N_4228,N_3545);
and U5369 (N_5369,N_3148,N_4875);
xor U5370 (N_5370,N_4709,N_3339);
nand U5371 (N_5371,N_4144,N_3429);
xor U5372 (N_5372,N_2731,N_2613);
or U5373 (N_5373,N_3483,N_2691);
nor U5374 (N_5374,N_4747,N_4530);
nor U5375 (N_5375,N_4645,N_3559);
and U5376 (N_5376,N_4351,N_3367);
nor U5377 (N_5377,N_4808,N_2598);
nand U5378 (N_5378,N_4867,N_2642);
nand U5379 (N_5379,N_2953,N_4872);
or U5380 (N_5380,N_4098,N_4186);
and U5381 (N_5381,N_2689,N_3616);
xnor U5382 (N_5382,N_2561,N_3809);
nand U5383 (N_5383,N_2743,N_3846);
nor U5384 (N_5384,N_4670,N_4677);
nand U5385 (N_5385,N_3681,N_3801);
nand U5386 (N_5386,N_3491,N_3862);
or U5387 (N_5387,N_4912,N_4807);
nor U5388 (N_5388,N_4383,N_3333);
nand U5389 (N_5389,N_4447,N_4197);
or U5390 (N_5390,N_3386,N_4547);
and U5391 (N_5391,N_3350,N_3149);
nor U5392 (N_5392,N_3081,N_4545);
and U5393 (N_5393,N_2867,N_2857);
and U5394 (N_5394,N_3109,N_2506);
and U5395 (N_5395,N_3268,N_4470);
xnor U5396 (N_5396,N_3922,N_3871);
nor U5397 (N_5397,N_4285,N_2656);
and U5398 (N_5398,N_2854,N_3547);
nand U5399 (N_5399,N_3031,N_4739);
nor U5400 (N_5400,N_3457,N_4277);
xor U5401 (N_5401,N_4162,N_3169);
xnor U5402 (N_5402,N_2842,N_4123);
xnor U5403 (N_5403,N_4033,N_3910);
or U5404 (N_5404,N_3422,N_4462);
and U5405 (N_5405,N_3565,N_4450);
nor U5406 (N_5406,N_2569,N_3518);
nor U5407 (N_5407,N_2958,N_4682);
nor U5408 (N_5408,N_4166,N_3264);
xnor U5409 (N_5409,N_3281,N_2873);
nor U5410 (N_5410,N_4027,N_2836);
xnor U5411 (N_5411,N_3745,N_4788);
and U5412 (N_5412,N_3026,N_2910);
and U5413 (N_5413,N_2713,N_3213);
xnor U5414 (N_5414,N_3611,N_4188);
nand U5415 (N_5415,N_3110,N_3313);
or U5416 (N_5416,N_3327,N_2553);
or U5417 (N_5417,N_4717,N_3966);
nand U5418 (N_5418,N_2852,N_3216);
xnor U5419 (N_5419,N_2596,N_3040);
and U5420 (N_5420,N_4503,N_3450);
and U5421 (N_5421,N_3535,N_2941);
nor U5422 (N_5422,N_3178,N_3398);
nor U5423 (N_5423,N_4891,N_4469);
or U5424 (N_5424,N_3021,N_2835);
or U5425 (N_5425,N_2916,N_3988);
nand U5426 (N_5426,N_4587,N_3501);
nor U5427 (N_5427,N_3601,N_2559);
xor U5428 (N_5428,N_3975,N_3306);
nand U5429 (N_5429,N_3680,N_3902);
and U5430 (N_5430,N_4581,N_2634);
xor U5431 (N_5431,N_4209,N_3311);
or U5432 (N_5432,N_4081,N_3512);
and U5433 (N_5433,N_4631,N_3442);
nor U5434 (N_5434,N_3948,N_2755);
nand U5435 (N_5435,N_3270,N_4965);
nand U5436 (N_5436,N_3642,N_4167);
and U5437 (N_5437,N_3395,N_4908);
nand U5438 (N_5438,N_4344,N_4736);
and U5439 (N_5439,N_4274,N_3918);
and U5440 (N_5440,N_3095,N_4636);
and U5441 (N_5441,N_4266,N_4222);
or U5442 (N_5442,N_2964,N_2974);
and U5443 (N_5443,N_2732,N_3805);
nand U5444 (N_5444,N_4301,N_4662);
or U5445 (N_5445,N_4131,N_3788);
nand U5446 (N_5446,N_4341,N_4825);
nor U5447 (N_5447,N_4619,N_4713);
nand U5448 (N_5448,N_3274,N_4036);
nor U5449 (N_5449,N_4031,N_3298);
xnor U5450 (N_5450,N_3369,N_3738);
nand U5451 (N_5451,N_3938,N_2627);
xor U5452 (N_5452,N_3868,N_3267);
nor U5453 (N_5453,N_4494,N_4782);
xnor U5454 (N_5454,N_4160,N_4063);
or U5455 (N_5455,N_3391,N_4904);
nand U5456 (N_5456,N_3419,N_4172);
nand U5457 (N_5457,N_3739,N_4243);
xnor U5458 (N_5458,N_4813,N_2860);
nor U5459 (N_5459,N_4307,N_2889);
xnor U5460 (N_5460,N_2967,N_4069);
or U5461 (N_5461,N_4618,N_4518);
xor U5462 (N_5462,N_3462,N_3795);
nor U5463 (N_5463,N_2716,N_4742);
xor U5464 (N_5464,N_3051,N_4170);
nand U5465 (N_5465,N_2825,N_3446);
nor U5466 (N_5466,N_3496,N_3017);
xnor U5467 (N_5467,N_3291,N_4404);
xor U5468 (N_5468,N_4420,N_4981);
or U5469 (N_5469,N_3779,N_4697);
and U5470 (N_5470,N_4302,N_3804);
and U5471 (N_5471,N_3528,N_4359);
nand U5472 (N_5472,N_3150,N_3328);
nand U5473 (N_5473,N_2500,N_4070);
or U5474 (N_5474,N_4286,N_4461);
and U5475 (N_5475,N_4921,N_3672);
or U5476 (N_5476,N_4270,N_2996);
xnor U5477 (N_5477,N_3405,N_3093);
or U5478 (N_5478,N_4305,N_3497);
and U5479 (N_5479,N_4475,N_3702);
or U5480 (N_5480,N_4025,N_3800);
nand U5481 (N_5481,N_2871,N_4492);
xor U5482 (N_5482,N_3122,N_3500);
nor U5483 (N_5483,N_4895,N_3467);
xor U5484 (N_5484,N_3006,N_4729);
nand U5485 (N_5485,N_3625,N_2893);
xor U5486 (N_5486,N_3623,N_4950);
and U5487 (N_5487,N_4429,N_4570);
xnor U5488 (N_5488,N_4418,N_2632);
xnor U5489 (N_5489,N_2913,N_4680);
nand U5490 (N_5490,N_3137,N_3167);
or U5491 (N_5491,N_4617,N_3124);
nor U5492 (N_5492,N_2805,N_4082);
or U5493 (N_5493,N_4865,N_3245);
xor U5494 (N_5494,N_3193,N_4995);
and U5495 (N_5495,N_4944,N_4767);
nand U5496 (N_5496,N_4741,N_2602);
nand U5497 (N_5497,N_4183,N_3753);
nor U5498 (N_5498,N_4146,N_3401);
nor U5499 (N_5499,N_4604,N_3546);
xor U5500 (N_5500,N_2542,N_4072);
xor U5501 (N_5501,N_4613,N_4393);
nand U5502 (N_5502,N_3061,N_4499);
or U5503 (N_5503,N_2661,N_4445);
and U5504 (N_5504,N_4093,N_2748);
xnor U5505 (N_5505,N_4366,N_3858);
nand U5506 (N_5506,N_4799,N_4859);
and U5507 (N_5507,N_3904,N_3892);
and U5508 (N_5508,N_3011,N_3084);
or U5509 (N_5509,N_2864,N_4189);
or U5510 (N_5510,N_3103,N_2591);
and U5511 (N_5511,N_3101,N_3571);
nor U5512 (N_5512,N_2711,N_3329);
nor U5513 (N_5513,N_3112,N_4575);
nor U5514 (N_5514,N_4542,N_2774);
xor U5515 (N_5515,N_4453,N_3699);
nor U5516 (N_5516,N_2969,N_3758);
nand U5517 (N_5517,N_4896,N_2900);
nand U5518 (N_5518,N_3825,N_4454);
nand U5519 (N_5519,N_3869,N_4472);
or U5520 (N_5520,N_2987,N_2802);
nor U5521 (N_5521,N_3581,N_4394);
nand U5522 (N_5522,N_3412,N_3478);
nor U5523 (N_5523,N_2810,N_4693);
and U5524 (N_5524,N_4565,N_4794);
nand U5525 (N_5525,N_2567,N_4380);
nand U5526 (N_5526,N_4043,N_4311);
nand U5527 (N_5527,N_3114,N_4369);
nor U5528 (N_5528,N_2667,N_2905);
or U5529 (N_5529,N_4971,N_3589);
xnor U5530 (N_5530,N_4668,N_3062);
and U5531 (N_5531,N_4443,N_4969);
or U5532 (N_5532,N_4015,N_3831);
nand U5533 (N_5533,N_4894,N_3654);
nand U5534 (N_5534,N_3675,N_4686);
nand U5535 (N_5535,N_2824,N_4478);
nor U5536 (N_5536,N_3555,N_3893);
nor U5537 (N_5537,N_3674,N_2728);
xnor U5538 (N_5538,N_4348,N_3789);
and U5539 (N_5539,N_2861,N_2979);
nor U5540 (N_5540,N_3817,N_4661);
xor U5541 (N_5541,N_3899,N_2766);
xnor U5542 (N_5542,N_2568,N_3089);
nand U5543 (N_5543,N_3807,N_4646);
nand U5544 (N_5544,N_3028,N_4844);
xnor U5545 (N_5545,N_4490,N_4019);
or U5546 (N_5546,N_3426,N_4110);
nor U5547 (N_5547,N_2580,N_3251);
nand U5548 (N_5548,N_4155,N_3349);
nand U5549 (N_5549,N_4673,N_2885);
nor U5550 (N_5550,N_2981,N_4863);
xnor U5551 (N_5551,N_3482,N_3056);
xor U5552 (N_5552,N_3141,N_4309);
xnor U5553 (N_5553,N_4580,N_4291);
xnor U5554 (N_5554,N_4145,N_4127);
nand U5555 (N_5555,N_4548,N_3657);
and U5556 (N_5556,N_4546,N_4026);
or U5557 (N_5557,N_2994,N_2539);
and U5558 (N_5558,N_4417,N_4939);
and U5559 (N_5559,N_2950,N_4034);
nand U5560 (N_5560,N_3253,N_2818);
and U5561 (N_5561,N_4452,N_4479);
and U5562 (N_5562,N_4828,N_3568);
xnor U5563 (N_5563,N_3411,N_3597);
nand U5564 (N_5564,N_3499,N_3840);
nand U5565 (N_5565,N_3624,N_4996);
or U5566 (N_5566,N_3550,N_4868);
xnor U5567 (N_5567,N_4495,N_3044);
xor U5568 (N_5568,N_3756,N_4018);
nor U5569 (N_5569,N_3673,N_3073);
nor U5570 (N_5570,N_4379,N_2724);
nor U5571 (N_5571,N_3074,N_3694);
nor U5572 (N_5572,N_3183,N_3289);
and U5573 (N_5573,N_3887,N_2653);
or U5574 (N_5574,N_3261,N_3959);
or U5575 (N_5575,N_2973,N_4022);
or U5576 (N_5576,N_4097,N_3204);
or U5577 (N_5577,N_4182,N_4664);
nor U5578 (N_5578,N_3697,N_3561);
or U5579 (N_5579,N_3479,N_3936);
or U5580 (N_5580,N_2605,N_3063);
nand U5581 (N_5581,N_3130,N_4818);
and U5582 (N_5582,N_3968,N_4073);
or U5583 (N_5583,N_4332,N_4902);
and U5584 (N_5584,N_4213,N_2637);
nand U5585 (N_5585,N_3459,N_3337);
xor U5586 (N_5586,N_2831,N_3476);
and U5587 (N_5587,N_3822,N_4774);
nand U5588 (N_5588,N_4400,N_4952);
or U5589 (N_5589,N_3260,N_4424);
xor U5590 (N_5590,N_4687,N_2633);
xnor U5591 (N_5591,N_4428,N_2740);
nand U5592 (N_5592,N_3985,N_2747);
nor U5593 (N_5593,N_3445,N_3331);
nand U5594 (N_5594,N_2899,N_4524);
nand U5595 (N_5595,N_2585,N_3631);
and U5596 (N_5596,N_3030,N_4365);
or U5597 (N_5597,N_4974,N_3470);
nor U5598 (N_5598,N_3543,N_2887);
nor U5599 (N_5599,N_3757,N_4052);
nor U5600 (N_5600,N_4190,N_4148);
xor U5601 (N_5601,N_3848,N_4220);
or U5602 (N_5602,N_2700,N_3864);
nor U5603 (N_5603,N_3992,N_3980);
or U5604 (N_5604,N_4361,N_3160);
or U5605 (N_5605,N_3618,N_4999);
or U5606 (N_5606,N_4249,N_3441);
xnor U5607 (N_5607,N_4810,N_4712);
nor U5608 (N_5608,N_3696,N_2844);
nand U5609 (N_5609,N_3345,N_4536);
xor U5610 (N_5610,N_3984,N_3896);
nand U5611 (N_5611,N_4039,N_2676);
xor U5612 (N_5612,N_4152,N_3861);
and U5613 (N_5613,N_4331,N_2984);
or U5614 (N_5614,N_4525,N_2839);
nor U5615 (N_5615,N_4579,N_4707);
and U5616 (N_5616,N_3782,N_4930);
xnor U5617 (N_5617,N_4923,N_4842);
xnor U5618 (N_5618,N_3821,N_3454);
nor U5619 (N_5619,N_3934,N_4991);
and U5620 (N_5620,N_4134,N_4803);
nand U5621 (N_5621,N_4966,N_3390);
nor U5622 (N_5622,N_2947,N_4836);
nor U5623 (N_5623,N_3226,N_4514);
xor U5624 (N_5624,N_2808,N_4625);
nand U5625 (N_5625,N_4573,N_3262);
and U5626 (N_5626,N_4440,N_3246);
and U5627 (N_5627,N_2597,N_3316);
nor U5628 (N_5628,N_4519,N_4501);
nor U5629 (N_5629,N_4367,N_4255);
nand U5630 (N_5630,N_2719,N_3269);
nor U5631 (N_5631,N_4870,N_3171);
and U5632 (N_5632,N_2828,N_4074);
and U5633 (N_5633,N_4308,N_3439);
nand U5634 (N_5634,N_3895,N_3125);
or U5635 (N_5635,N_4143,N_2654);
or U5636 (N_5636,N_3797,N_2510);
and U5637 (N_5637,N_2813,N_3032);
and U5638 (N_5638,N_3362,N_2926);
xor U5639 (N_5639,N_2920,N_2760);
nor U5640 (N_5640,N_3981,N_4463);
and U5641 (N_5641,N_3250,N_3008);
xnor U5642 (N_5642,N_4423,N_2603);
nand U5643 (N_5643,N_3020,N_4109);
nor U5644 (N_5644,N_2655,N_2753);
or U5645 (N_5645,N_4523,N_3489);
xor U5646 (N_5646,N_2599,N_2798);
xnor U5647 (N_5647,N_4840,N_3159);
nor U5648 (N_5648,N_3050,N_3228);
or U5649 (N_5649,N_4092,N_4688);
nor U5650 (N_5650,N_3048,N_3060);
nand U5651 (N_5651,N_4107,N_3835);
or U5652 (N_5652,N_2955,N_2681);
nor U5653 (N_5653,N_4956,N_4150);
nor U5654 (N_5654,N_3205,N_3255);
or U5655 (N_5655,N_4694,N_4426);
nor U5656 (N_5656,N_4323,N_2901);
nor U5657 (N_5657,N_4582,N_4275);
xor U5658 (N_5658,N_3588,N_3708);
and U5659 (N_5659,N_3147,N_3750);
nand U5660 (N_5660,N_3544,N_3094);
and U5661 (N_5661,N_3107,N_2972);
nor U5662 (N_5662,N_4473,N_4168);
and U5663 (N_5663,N_4622,N_4679);
nand U5664 (N_5664,N_4234,N_4753);
xnor U5665 (N_5665,N_3098,N_3091);
and U5666 (N_5666,N_3608,N_4381);
and U5667 (N_5667,N_4038,N_4569);
or U5668 (N_5668,N_4253,N_2814);
or U5669 (N_5669,N_4481,N_4199);
xor U5670 (N_5670,N_3877,N_3873);
nor U5671 (N_5671,N_3009,N_2649);
xor U5672 (N_5672,N_4811,N_4203);
nor U5673 (N_5673,N_4772,N_3024);
nand U5674 (N_5674,N_2697,N_3312);
nand U5675 (N_5675,N_4953,N_4207);
and U5676 (N_5676,N_4246,N_3434);
xor U5677 (N_5677,N_3913,N_4245);
xnor U5678 (N_5678,N_3880,N_3580);
xnor U5679 (N_5679,N_3220,N_4271);
nand U5680 (N_5680,N_4620,N_4639);
nand U5681 (N_5681,N_3838,N_3556);
and U5682 (N_5682,N_4306,N_3466);
nor U5683 (N_5683,N_4609,N_4464);
xor U5684 (N_5684,N_4577,N_2937);
and U5685 (N_5685,N_3630,N_4549);
and U5686 (N_5686,N_4094,N_4084);
xor U5687 (N_5687,N_3431,N_3780);
or U5688 (N_5688,N_4730,N_4053);
and U5689 (N_5689,N_3690,N_4139);
nor U5690 (N_5690,N_3065,N_3662);
and U5691 (N_5691,N_3921,N_3004);
and U5692 (N_5692,N_3560,N_2888);
or U5693 (N_5693,N_4970,N_3823);
and U5694 (N_5694,N_2817,N_4376);
and U5695 (N_5695,N_4733,N_4435);
nor U5696 (N_5696,N_4983,N_4412);
and U5697 (N_5697,N_4945,N_2536);
or U5698 (N_5698,N_2601,N_3995);
xor U5699 (N_5699,N_3746,N_4723);
nand U5700 (N_5700,N_2530,N_2843);
xnor U5701 (N_5701,N_2980,N_4614);
and U5702 (N_5702,N_2560,N_3161);
and U5703 (N_5703,N_2670,N_4780);
or U5704 (N_5704,N_4911,N_4691);
and U5705 (N_5705,N_3824,N_4987);
or U5706 (N_5706,N_4749,N_4205);
xor U5707 (N_5707,N_2715,N_2781);
nand U5708 (N_5708,N_3609,N_2868);
or U5709 (N_5709,N_2699,N_4388);
nand U5710 (N_5710,N_4003,N_2710);
nor U5711 (N_5711,N_3187,N_2912);
and U5712 (N_5712,N_3964,N_4137);
nor U5713 (N_5713,N_3071,N_2856);
and U5714 (N_5714,N_3198,N_3233);
or U5715 (N_5715,N_4663,N_4104);
nand U5716 (N_5716,N_4161,N_2617);
nand U5717 (N_5717,N_3731,N_2918);
and U5718 (N_5718,N_3876,N_3953);
or U5719 (N_5719,N_4165,N_3530);
or U5720 (N_5720,N_3325,N_3941);
xnor U5721 (N_5721,N_3718,N_4180);
or U5722 (N_5722,N_4724,N_4362);
nand U5723 (N_5723,N_4516,N_3813);
nand U5724 (N_5724,N_2594,N_4313);
nor U5725 (N_5725,N_3019,N_3430);
nand U5726 (N_5726,N_3140,N_4821);
and U5727 (N_5727,N_4347,N_3305);
xor U5728 (N_5728,N_3540,N_3837);
xor U5729 (N_5729,N_3969,N_4600);
nand U5730 (N_5730,N_3389,N_4173);
nor U5731 (N_5731,N_4889,N_4650);
and U5732 (N_5732,N_2942,N_3352);
and U5733 (N_5733,N_4564,N_4218);
and U5734 (N_5734,N_3635,N_3104);
nand U5735 (N_5735,N_4903,N_3487);
nand U5736 (N_5736,N_2922,N_4676);
xor U5737 (N_5737,N_3640,N_3852);
xor U5738 (N_5738,N_2954,N_3907);
and U5739 (N_5739,N_3927,N_2758);
xor U5740 (N_5740,N_2564,N_4158);
and U5741 (N_5741,N_4300,N_3400);
and U5742 (N_5742,N_3715,N_3029);
nand U5743 (N_5743,N_3593,N_4326);
or U5744 (N_5744,N_4415,N_2712);
and U5745 (N_5745,N_3740,N_3818);
nand U5746 (N_5746,N_3916,N_3799);
and U5747 (N_5747,N_4752,N_4932);
nor U5748 (N_5748,N_4496,N_2795);
xor U5749 (N_5749,N_2593,N_3721);
nor U5750 (N_5750,N_2589,N_4163);
and U5751 (N_5751,N_3897,N_4963);
and U5752 (N_5752,N_2572,N_2787);
nor U5753 (N_5753,N_3272,N_3455);
nand U5754 (N_5754,N_2720,N_4728);
or U5755 (N_5755,N_3237,N_4869);
and U5756 (N_5756,N_4201,N_3201);
xnor U5757 (N_5757,N_3703,N_4298);
nand U5758 (N_5758,N_3355,N_3872);
or U5759 (N_5759,N_3259,N_4527);
and U5760 (N_5760,N_3863,N_2761);
nor U5761 (N_5761,N_3035,N_4861);
and U5762 (N_5762,N_4674,N_2894);
and U5763 (N_5763,N_2945,N_3855);
nor U5764 (N_5764,N_2997,N_3287);
or U5765 (N_5765,N_3314,N_3087);
or U5766 (N_5766,N_2725,N_2845);
or U5767 (N_5767,N_4898,N_3242);
xnor U5768 (N_5768,N_4493,N_4929);
or U5769 (N_5769,N_3144,N_4061);
and U5770 (N_5770,N_4319,N_3626);
xnor U5771 (N_5771,N_2614,N_3573);
xor U5772 (N_5772,N_3477,N_3549);
xnor U5773 (N_5773,N_4411,N_4824);
or U5774 (N_5774,N_3610,N_4382);
and U5775 (N_5775,N_2570,N_3664);
and U5776 (N_5776,N_3594,N_4737);
xnor U5777 (N_5777,N_4363,N_3612);
xor U5778 (N_5778,N_2777,N_2799);
and U5779 (N_5779,N_4701,N_4050);
xor U5780 (N_5780,N_4002,N_4268);
and U5781 (N_5781,N_4095,N_4259);
xor U5782 (N_5782,N_3138,N_3282);
and U5783 (N_5783,N_4132,N_3003);
or U5784 (N_5784,N_4075,N_2992);
nor U5785 (N_5785,N_4779,N_3973);
nor U5786 (N_5786,N_3531,N_4088);
nand U5787 (N_5787,N_3173,N_2707);
nor U5788 (N_5788,N_3128,N_4839);
nor U5789 (N_5789,N_4511,N_3859);
nand U5790 (N_5790,N_2662,N_3319);
xor U5791 (N_5791,N_4578,N_4714);
nor U5792 (N_5792,N_4922,N_3775);
nand U5793 (N_5793,N_2600,N_4101);
nand U5794 (N_5794,N_3153,N_4321);
nor U5795 (N_5795,N_3716,N_3787);
nor U5796 (N_5796,N_3679,N_2759);
and U5797 (N_5797,N_4007,N_4715);
and U5798 (N_5798,N_3085,N_3651);
and U5799 (N_5799,N_4700,N_3870);
and U5800 (N_5800,N_2862,N_2531);
and U5801 (N_5801,N_2865,N_3378);
or U5802 (N_5802,N_3647,N_4938);
nand U5803 (N_5803,N_3244,N_3595);
and U5804 (N_5804,N_4960,N_3803);
xnor U5805 (N_5805,N_4936,N_4507);
nand U5806 (N_5806,N_4059,N_4040);
or U5807 (N_5807,N_3357,N_3123);
nor U5808 (N_5808,N_3208,N_2838);
nand U5809 (N_5809,N_2626,N_2765);
xnor U5810 (N_5810,N_3162,N_3473);
nand U5811 (N_5811,N_4718,N_3326);
xor U5812 (N_5812,N_4176,N_2650);
or U5813 (N_5813,N_3285,N_3653);
nor U5814 (N_5814,N_2978,N_2776);
nor U5815 (N_5815,N_3279,N_2993);
and U5816 (N_5816,N_4817,N_3977);
and U5817 (N_5817,N_3037,N_3997);
nand U5818 (N_5818,N_2931,N_2548);
nand U5819 (N_5819,N_4883,N_3529);
or U5820 (N_5820,N_4409,N_2923);
xnor U5821 (N_5821,N_4179,N_4497);
or U5822 (N_5822,N_4005,N_4226);
nand U5823 (N_5823,N_2919,N_3385);
nor U5824 (N_5824,N_3639,N_3785);
and U5825 (N_5825,N_4049,N_3706);
nor U5826 (N_5826,N_4358,N_3575);
nand U5827 (N_5827,N_3743,N_3365);
nor U5828 (N_5828,N_2756,N_2907);
or U5829 (N_5829,N_4407,N_4047);
nand U5830 (N_5830,N_4103,N_4611);
xor U5831 (N_5831,N_4416,N_3155);
xor U5832 (N_5832,N_3384,N_3767);
and U5833 (N_5833,N_4233,N_3971);
nor U5834 (N_5834,N_4335,N_4602);
and U5835 (N_5835,N_2677,N_4798);
or U5836 (N_5836,N_3338,N_3041);
nand U5837 (N_5837,N_4616,N_4009);
xor U5838 (N_5838,N_3300,N_4194);
xnor U5839 (N_5839,N_4368,N_4195);
nor U5840 (N_5840,N_2790,N_4598);
xor U5841 (N_5841,N_2604,N_4558);
or U5842 (N_5842,N_3336,N_2535);
nand U5843 (N_5843,N_3340,N_2566);
and U5844 (N_5844,N_4405,N_4489);
and U5845 (N_5845,N_4504,N_4451);
nand U5846 (N_5846,N_3843,N_4130);
nand U5847 (N_5847,N_3562,N_3722);
nor U5848 (N_5848,N_3121,N_4403);
and U5849 (N_5849,N_3683,N_4689);
and U5850 (N_5850,N_4138,N_4681);
nand U5851 (N_5851,N_3066,N_3794);
xnor U5852 (N_5852,N_3983,N_3058);
nor U5853 (N_5853,N_4623,N_4822);
and U5854 (N_5854,N_3210,N_2540);
nor U5855 (N_5855,N_3485,N_2643);
xnor U5856 (N_5856,N_3175,N_3135);
xor U5857 (N_5857,N_3036,N_3387);
nand U5858 (N_5858,N_3576,N_3717);
xnor U5859 (N_5859,N_3707,N_4881);
or U5860 (N_5860,N_4370,N_2680);
xor U5861 (N_5861,N_4455,N_4425);
nor U5862 (N_5862,N_2971,N_4760);
or U5863 (N_5863,N_4389,N_4644);
xor U5864 (N_5864,N_2578,N_4540);
nand U5865 (N_5865,N_3937,N_2671);
nor U5866 (N_5866,N_4607,N_4816);
or U5867 (N_5867,N_4743,N_3613);
nor U5868 (N_5868,N_3403,N_4785);
nor U5869 (N_5869,N_2961,N_2830);
xor U5870 (N_5870,N_2696,N_2565);
or U5871 (N_5871,N_3730,N_4576);
and U5872 (N_5872,N_2620,N_4283);
or U5873 (N_5873,N_2879,N_2646);
or U5874 (N_5874,N_4360,N_3363);
nand U5875 (N_5875,N_4541,N_4432);
or U5876 (N_5876,N_4385,N_4353);
nor U5877 (N_5877,N_4304,N_4692);
nor U5878 (N_5878,N_4154,N_3709);
nand U5879 (N_5879,N_3420,N_2866);
xor U5880 (N_5880,N_4374,N_4990);
and U5881 (N_5881,N_2551,N_3894);
nor U5882 (N_5882,N_4927,N_2615);
nand U5883 (N_5883,N_4467,N_2952);
nor U5884 (N_5884,N_3510,N_4242);
xnor U5885 (N_5885,N_2730,N_4766);
xnor U5886 (N_5886,N_4528,N_3214);
and U5887 (N_5887,N_4621,N_3448);
xnor U5888 (N_5888,N_2538,N_4937);
and U5889 (N_5889,N_4832,N_4834);
or U5890 (N_5890,N_3453,N_3295);
nand U5891 (N_5891,N_3053,N_3558);
and U5892 (N_5892,N_3538,N_3195);
xor U5893 (N_5893,N_2850,N_4985);
xnor U5894 (N_5894,N_3392,N_2524);
nand U5895 (N_5895,N_3834,N_3047);
nor U5896 (N_5896,N_2869,N_4770);
xor U5897 (N_5897,N_3532,N_3067);
xnor U5898 (N_5898,N_4560,N_3710);
nor U5899 (N_5899,N_2794,N_3903);
or U5900 (N_5900,N_3845,N_4876);
nor U5901 (N_5901,N_4122,N_4975);
xnor U5902 (N_5902,N_4638,N_2611);
xor U5903 (N_5903,N_4288,N_4637);
and U5904 (N_5904,N_4272,N_3513);
and U5905 (N_5905,N_3108,N_4833);
nor U5906 (N_5906,N_3670,N_4175);
and U5907 (N_5907,N_4008,N_3660);
or U5908 (N_5908,N_2929,N_3257);
xor U5909 (N_5909,N_3438,N_4468);
nor U5910 (N_5910,N_2841,N_3247);
or U5911 (N_5911,N_4820,N_3303);
xnor U5912 (N_5912,N_4419,N_3604);
nand U5913 (N_5913,N_4334,N_4299);
and U5914 (N_5914,N_3152,N_2652);
nand U5915 (N_5915,N_3579,N_3078);
and U5916 (N_5916,N_3374,N_2722);
xnor U5917 (N_5917,N_3620,N_2638);
nand U5918 (N_5918,N_4431,N_4413);
xor U5919 (N_5919,N_3714,N_3553);
xnor U5920 (N_5920,N_4716,N_2816);
nor U5921 (N_5921,N_4732,N_3217);
and U5922 (N_5922,N_2573,N_2773);
or U5923 (N_5923,N_4989,N_3304);
nand U5924 (N_5924,N_4802,N_2526);
and U5925 (N_5925,N_3396,N_4791);
nand U5926 (N_5926,N_4510,N_3860);
and U5927 (N_5927,N_3901,N_3106);
nand U5928 (N_5928,N_4121,N_4483);
nand U5929 (N_5929,N_3358,N_3587);
nand U5930 (N_5930,N_3055,N_3443);
or U5931 (N_5931,N_3393,N_3188);
and U5932 (N_5932,N_3723,N_2664);
nand U5933 (N_5933,N_3777,N_4488);
and U5934 (N_5934,N_4231,N_3914);
nand U5935 (N_5935,N_4608,N_3712);
nand U5936 (N_5936,N_3979,N_3168);
and U5937 (N_5937,N_2815,N_4159);
xnor U5938 (N_5938,N_4585,N_4215);
nand U5939 (N_5939,N_3002,N_4108);
and U5940 (N_5940,N_2881,N_2809);
or U5941 (N_5941,N_4265,N_3010);
or U5942 (N_5942,N_4805,N_4236);
xor U5943 (N_5943,N_4422,N_4702);
nand U5944 (N_5944,N_4543,N_2588);
nor U5945 (N_5945,N_2574,N_3354);
nand U5946 (N_5946,N_3243,N_4913);
and U5947 (N_5947,N_2915,N_4586);
nor U5948 (N_5948,N_4556,N_4862);
or U5949 (N_5949,N_2764,N_4856);
or U5950 (N_5950,N_3878,N_3748);
nor U5951 (N_5951,N_4136,N_4789);
or U5952 (N_5952,N_4260,N_3976);
xor U5953 (N_5953,N_3816,N_4986);
nand U5954 (N_5954,N_2735,N_2988);
xor U5955 (N_5955,N_3521,N_4210);
nand U5956 (N_5956,N_4191,N_3016);
and U5957 (N_5957,N_4320,N_4433);
and U5958 (N_5958,N_4641,N_3286);
nor U5959 (N_5959,N_3227,N_4685);
nand U5960 (N_5960,N_2714,N_4725);
or U5961 (N_5961,N_3957,N_4877);
or U5962 (N_5962,N_4346,N_3853);
or U5963 (N_5963,N_3695,N_2991);
xnor U5964 (N_5964,N_4695,N_2998);
xnor U5965 (N_5965,N_4227,N_3998);
nand U5966 (N_5966,N_3164,N_4269);
nor U5967 (N_5967,N_3366,N_3842);
and U5968 (N_5968,N_3423,N_3406);
xor U5969 (N_5969,N_3668,N_4751);
nor U5970 (N_5970,N_4906,N_2675);
and U5971 (N_5971,N_4444,N_3359);
and U5972 (N_5972,N_4924,N_3923);
and U5973 (N_5973,N_3506,N_2925);
nor U5974 (N_5974,N_3725,N_4632);
and U5975 (N_5975,N_3219,N_4955);
or U5976 (N_5976,N_3541,N_4252);
nand U5977 (N_5977,N_3427,N_4731);
nor U5978 (N_5978,N_4571,N_3280);
xor U5979 (N_5979,N_4857,N_2706);
and U5980 (N_5980,N_4312,N_3841);
and U5981 (N_5981,N_4206,N_4758);
nand U5982 (N_5982,N_4634,N_3113);
and U5983 (N_5983,N_4892,N_2678);
nand U5984 (N_5984,N_4761,N_4322);
and U5985 (N_5985,N_3646,N_2986);
xnor U5986 (N_5986,N_3592,N_4441);
xor U5987 (N_5987,N_4552,N_4943);
nand U5988 (N_5988,N_3263,N_2911);
and U5989 (N_5989,N_4077,N_4853);
nand U5990 (N_5990,N_4221,N_3469);
nand U5991 (N_5991,N_4553,N_4147);
or U5992 (N_5992,N_3481,N_2948);
or U5993 (N_5993,N_4278,N_4544);
xor U5994 (N_5994,N_3554,N_2727);
xnor U5995 (N_5995,N_4427,N_3886);
and U5996 (N_5996,N_2515,N_3057);
and U5997 (N_5997,N_4705,N_3925);
xnor U5998 (N_5998,N_3898,N_4667);
and U5999 (N_5999,N_2963,N_3404);
nor U6000 (N_6000,N_4698,N_3928);
xnor U6001 (N_6001,N_2791,N_2644);
or U6002 (N_6002,N_4949,N_2721);
nor U6003 (N_6003,N_4659,N_4551);
xor U6004 (N_6004,N_2970,N_3636);
and U6005 (N_6005,N_4601,N_4775);
nor U6006 (N_6006,N_3435,N_3522);
nand U6007 (N_6007,N_2704,N_2630);
xor U6008 (N_6008,N_2834,N_2872);
or U6009 (N_6009,N_3563,N_3633);
or U6010 (N_6010,N_3627,N_2851);
nor U6011 (N_6011,N_2616,N_4769);
xor U6012 (N_6012,N_2726,N_2622);
nand U6013 (N_6013,N_3283,N_2503);
nor U6014 (N_6014,N_2693,N_3176);
nor U6015 (N_6015,N_3798,N_4886);
xor U6016 (N_6016,N_3951,N_4350);
or U6017 (N_6017,N_3296,N_3231);
or U6018 (N_6018,N_2750,N_3962);
nand U6019 (N_6019,N_3742,N_4652);
xor U6020 (N_6020,N_3888,N_4056);
or U6021 (N_6021,N_4142,N_3083);
nand U6022 (N_6022,N_3102,N_4893);
or U6023 (N_6023,N_3819,N_3288);
and U6024 (N_6024,N_3383,N_3996);
or U6025 (N_6025,N_4851,N_3090);
nor U6026 (N_6026,N_4720,N_3145);
or U6027 (N_6027,N_4067,N_3347);
xor U6028 (N_6028,N_2682,N_4643);
xnor U6029 (N_6029,N_3341,N_2853);
or U6030 (N_6030,N_3751,N_3940);
nor U6031 (N_6031,N_4854,N_4219);
nor U6032 (N_6032,N_4449,N_3472);
nor U6033 (N_6033,N_2522,N_3077);
nor U6034 (N_6034,N_2821,N_3271);
and U6035 (N_6035,N_3701,N_4783);
and U6036 (N_6036,N_2793,N_4792);
and U6037 (N_6037,N_3602,N_3129);
and U6038 (N_6038,N_3667,N_2645);
nand U6039 (N_6039,N_3688,N_4232);
nand U6040 (N_6040,N_2829,N_3461);
or U6041 (N_6041,N_2555,N_3018);
xnor U6042 (N_6042,N_3956,N_4153);
nand U6043 (N_6043,N_3133,N_3737);
and U6044 (N_6044,N_4459,N_2846);
xor U6045 (N_6045,N_3025,N_2672);
nand U6046 (N_6046,N_3564,N_2592);
nor U6047 (N_6047,N_4214,N_3033);
nor U6048 (N_6048,N_2534,N_3464);
nor U6049 (N_6049,N_4654,N_4529);
nor U6050 (N_6050,N_4235,N_3407);
nand U6051 (N_6051,N_4297,N_4651);
or U6052 (N_6052,N_4247,N_3307);
nand U6053 (N_6053,N_3814,N_4606);
xor U6054 (N_6054,N_2501,N_4184);
nor U6055 (N_6055,N_4113,N_4790);
nand U6056 (N_6056,N_3682,N_3584);
or U6057 (N_6057,N_2624,N_2587);
nor U6058 (N_6058,N_3402,N_3111);
nand U6059 (N_6059,N_2819,N_3526);
nor U6060 (N_6060,N_4013,N_3637);
or U6061 (N_6061,N_4915,N_3117);
nor U6062 (N_6062,N_3954,N_4829);
and U6063 (N_6063,N_4845,N_4048);
nand U6064 (N_6064,N_2586,N_2966);
nand U6065 (N_6065,N_3605,N_4333);
nand U6066 (N_6066,N_4157,N_3754);
and U6067 (N_6067,N_2882,N_2896);
nand U6068 (N_6068,N_3557,N_4653);
or U6069 (N_6069,N_4841,N_3503);
xor U6070 (N_6070,N_4402,N_4085);
and U6071 (N_6071,N_3206,N_3038);
xnor U6072 (N_6072,N_4880,N_2658);
nand U6073 (N_6073,N_4978,N_3486);
xor U6074 (N_6074,N_2982,N_3317);
nor U6075 (N_6075,N_4125,N_3471);
and U6076 (N_6076,N_2833,N_4257);
nor U6077 (N_6077,N_2975,N_4119);
and U6078 (N_6078,N_4941,N_3719);
nor U6079 (N_6079,N_2771,N_4890);
and U6080 (N_6080,N_3586,N_3364);
nand U6081 (N_6081,N_4016,N_4340);
xor U6082 (N_6082,N_4672,N_4171);
nor U6083 (N_6083,N_3866,N_3495);
nand U6084 (N_6084,N_4909,N_3509);
or U6085 (N_6085,N_3309,N_3203);
and U6086 (N_6086,N_2744,N_2576);
or U6087 (N_6087,N_3096,N_4599);
or U6088 (N_6088,N_4660,N_2801);
or U6089 (N_6089,N_4554,N_2512);
nand U6090 (N_6090,N_3600,N_3749);
or U6091 (N_6091,N_3290,N_4001);
and U6092 (N_6092,N_3511,N_2891);
or U6093 (N_6093,N_4846,N_3815);
nand U6094 (N_6094,N_4994,N_4649);
and U6095 (N_6095,N_4120,N_3949);
or U6096 (N_6096,N_2837,N_2823);
xor U6097 (N_6097,N_3615,N_3915);
or U6098 (N_6098,N_3874,N_4006);
or U6099 (N_6099,N_4905,N_4041);
nor U6100 (N_6100,N_3027,N_2749);
nand U6101 (N_6101,N_4665,N_4051);
nand U6102 (N_6102,N_2608,N_4568);
or U6103 (N_6103,N_4212,N_2874);
nor U6104 (N_6104,N_3686,N_4678);
and U6105 (N_6105,N_4848,N_3174);
or U6106 (N_6106,N_4352,N_2657);
and U6107 (N_6107,N_3371,N_3428);
nor U6108 (N_6108,N_2762,N_4635);
nand U6109 (N_6109,N_3185,N_4781);
and U6110 (N_6110,N_2612,N_2546);
nor U6111 (N_6111,N_4421,N_4942);
nor U6112 (N_6112,N_4193,N_4456);
nor U6113 (N_6113,N_2886,N_4648);
xnor U6114 (N_6114,N_3045,N_3007);
nor U6115 (N_6115,N_4465,N_4202);
nor U6116 (N_6116,N_3377,N_3638);
or U6117 (N_6117,N_2892,N_2659);
xor U6118 (N_6118,N_3492,N_4849);
xnor U6119 (N_6119,N_4343,N_3569);
nor U6120 (N_6120,N_4364,N_4112);
nor U6121 (N_6121,N_4457,N_4011);
and U6122 (N_6122,N_4968,N_2995);
nor U6123 (N_6123,N_4096,N_3069);
nand U6124 (N_6124,N_3732,N_4603);
and U6125 (N_6125,N_4940,N_2932);
and U6126 (N_6126,N_2737,N_3042);
nor U6127 (N_6127,N_3381,N_3082);
nand U6128 (N_6128,N_2647,N_4823);
or U6129 (N_6129,N_3458,N_4390);
or U6130 (N_6130,N_3829,N_4254);
or U6131 (N_6131,N_2921,N_4873);
or U6132 (N_6132,N_4993,N_3105);
nor U6133 (N_6133,N_4296,N_4020);
nand U6134 (N_6134,N_2674,N_2619);
or U6135 (N_6135,N_4263,N_3207);
nor U6136 (N_6136,N_4241,N_4140);
nand U6137 (N_6137,N_4316,N_3310);
xor U6138 (N_6138,N_4303,N_3677);
nand U6139 (N_6139,N_4115,N_2609);
and U6140 (N_6140,N_4126,N_4436);
nand U6141 (N_6141,N_4738,N_3747);
xor U6142 (N_6142,N_2924,N_3987);
or U6143 (N_6143,N_2581,N_3693);
xor U6144 (N_6144,N_2884,N_3905);
nand U6145 (N_6145,N_2505,N_4187);
nor U6146 (N_6146,N_2778,N_3502);
xnor U6147 (N_6147,N_2745,N_3790);
nor U6148 (N_6148,N_4948,N_4624);
xor U6149 (N_6149,N_2504,N_2933);
nand U6150 (N_6150,N_4809,N_2792);
or U6151 (N_6151,N_4593,N_3520);
and U6152 (N_6152,N_4078,N_4897);
nand U6153 (N_6153,N_2552,N_4315);
and U6154 (N_6154,N_3361,N_2606);
nor U6155 (N_6155,N_3771,N_3342);
xor U6156 (N_6156,N_4884,N_3851);
xor U6157 (N_6157,N_4192,N_4690);
nor U6158 (N_6158,N_2757,N_4610);
or U6159 (N_6159,N_2796,N_4055);
and U6160 (N_6160,N_4984,N_3225);
or U6161 (N_6161,N_4273,N_4843);
nand U6162 (N_6162,N_3508,N_4946);
or U6163 (N_6163,N_3116,N_3632);
nor U6164 (N_6164,N_3218,N_2507);
nor U6165 (N_6165,N_2772,N_2780);
nand U6166 (N_6166,N_4062,N_4330);
or U6167 (N_6167,N_2528,N_4329);
and U6168 (N_6168,N_3946,N_4030);
xnor U6169 (N_6169,N_3856,N_3523);
and U6170 (N_6170,N_2519,N_2983);
or U6171 (N_6171,N_4583,N_3891);
xor U6172 (N_6172,N_2768,N_3200);
nor U6173 (N_6173,N_2985,N_3590);
xor U6174 (N_6174,N_3881,N_3000);
nor U6175 (N_6175,N_3023,N_4657);
nor U6176 (N_6176,N_4133,N_3351);
nand U6177 (N_6177,N_3978,N_3755);
xnor U6178 (N_6178,N_2521,N_3570);
or U6179 (N_6179,N_3131,N_3239);
xor U6180 (N_6180,N_4982,N_3059);
xnor U6181 (N_6181,N_2832,N_3068);
nand U6182 (N_6182,N_4793,N_3127);
and U6183 (N_6183,N_3548,N_3172);
nor U6184 (N_6184,N_4972,N_4976);
xnor U6185 (N_6185,N_4590,N_3711);
xor U6186 (N_6186,N_3356,N_3942);
nand U6187 (N_6187,N_4550,N_4392);
xnor U6188 (N_6188,N_3012,N_4696);
nand U6189 (N_6189,N_4458,N_4264);
xnor U6190 (N_6190,N_3598,N_4498);
nor U6191 (N_6191,N_4795,N_3229);
nor U6192 (N_6192,N_4177,N_3241);
xor U6193 (N_6193,N_4100,N_2575);
nor U6194 (N_6194,N_3854,N_4612);
xor U6195 (N_6195,N_3939,N_4847);
and U6196 (N_6196,N_3232,N_3659);
or U6197 (N_6197,N_4562,N_3299);
nor U6198 (N_6198,N_4484,N_3505);
and U6199 (N_6199,N_3882,N_2938);
and U6200 (N_6200,N_3828,N_3235);
nand U6201 (N_6201,N_4827,N_3379);
nand U6202 (N_6202,N_3525,N_4357);
nand U6203 (N_6203,N_4487,N_4916);
nor U6204 (N_6204,N_2804,N_3599);
nor U6205 (N_6205,N_3484,N_4726);
or U6206 (N_6206,N_3982,N_2956);
nor U6207 (N_6207,N_4124,N_4083);
nor U6208 (N_6208,N_4882,N_4114);
nor U6209 (N_6209,N_2688,N_3115);
nor U6210 (N_6210,N_3524,N_3652);
and U6211 (N_6211,N_3830,N_2946);
xor U6212 (N_6212,N_3301,N_4196);
and U6213 (N_6213,N_3644,N_2763);
xor U6214 (N_6214,N_2557,N_4706);
and U6215 (N_6215,N_4812,N_2669);
or U6216 (N_6216,N_3645,N_2739);
and U6217 (N_6217,N_3397,N_4704);
xor U6218 (N_6218,N_3034,N_2679);
or U6219 (N_6219,N_4628,N_2935);
nand U6220 (N_6220,N_4279,N_4128);
and U6221 (N_6221,N_4399,N_4010);
or U6222 (N_6222,N_3713,N_3741);
nand U6223 (N_6223,N_3617,N_4282);
nor U6224 (N_6224,N_3418,N_4037);
and U6225 (N_6225,N_2951,N_2705);
or U6226 (N_6226,N_3186,N_4973);
xnor U6227 (N_6227,N_3906,N_3974);
or U6228 (N_6228,N_2976,N_3970);
or U6229 (N_6229,N_3577,N_3234);
nor U6230 (N_6230,N_3967,N_4735);
nand U6231 (N_6231,N_3099,N_3772);
or U6232 (N_6232,N_3582,N_4058);
and U6233 (N_6233,N_3046,N_3700);
nor U6234 (N_6234,N_4198,N_4091);
nand U6235 (N_6235,N_3146,N_3415);
or U6236 (N_6236,N_3578,N_2684);
nor U6237 (N_6237,N_3324,N_3236);
nor U6238 (N_6238,N_4878,N_3156);
nand U6239 (N_6239,N_2807,N_3678);
and U6240 (N_6240,N_4885,N_4538);
or U6241 (N_6241,N_4931,N_2939);
nand U6242 (N_6242,N_4239,N_3480);
nand U6243 (N_6243,N_4446,N_2859);
and U6244 (N_6244,N_2718,N_4719);
nand U6245 (N_6245,N_3373,N_3022);
nand U6246 (N_6246,N_2533,N_4023);
xor U6247 (N_6247,N_3826,N_3368);
nor U6248 (N_6248,N_4460,N_4773);
and U6249 (N_6249,N_3917,N_4338);
nand U6250 (N_6250,N_3519,N_4658);
nand U6251 (N_6251,N_3153,N_3920);
xor U6252 (N_6252,N_3982,N_4675);
and U6253 (N_6253,N_2748,N_4392);
xnor U6254 (N_6254,N_4845,N_4343);
or U6255 (N_6255,N_3558,N_3962);
xnor U6256 (N_6256,N_3174,N_3460);
nor U6257 (N_6257,N_2594,N_4523);
or U6258 (N_6258,N_2543,N_3492);
nand U6259 (N_6259,N_4741,N_3176);
or U6260 (N_6260,N_2850,N_4164);
nor U6261 (N_6261,N_3081,N_4680);
xnor U6262 (N_6262,N_4976,N_3068);
xor U6263 (N_6263,N_3082,N_4875);
xnor U6264 (N_6264,N_3331,N_4068);
nand U6265 (N_6265,N_2846,N_3364);
nand U6266 (N_6266,N_2542,N_4748);
and U6267 (N_6267,N_3343,N_4867);
nand U6268 (N_6268,N_3955,N_4514);
and U6269 (N_6269,N_4965,N_2589);
xnor U6270 (N_6270,N_4329,N_2842);
and U6271 (N_6271,N_4914,N_4743);
and U6272 (N_6272,N_3410,N_4016);
and U6273 (N_6273,N_3844,N_3381);
and U6274 (N_6274,N_2523,N_3120);
or U6275 (N_6275,N_3169,N_4078);
nand U6276 (N_6276,N_3416,N_2892);
xor U6277 (N_6277,N_4109,N_2981);
xnor U6278 (N_6278,N_3363,N_4528);
and U6279 (N_6279,N_3461,N_4227);
and U6280 (N_6280,N_3096,N_3358);
nand U6281 (N_6281,N_3075,N_3742);
xnor U6282 (N_6282,N_3708,N_2896);
nand U6283 (N_6283,N_4689,N_4798);
xor U6284 (N_6284,N_4727,N_3021);
or U6285 (N_6285,N_2566,N_2626);
or U6286 (N_6286,N_4691,N_4831);
and U6287 (N_6287,N_4852,N_4333);
xor U6288 (N_6288,N_4195,N_4291);
xnor U6289 (N_6289,N_4250,N_4795);
nand U6290 (N_6290,N_3643,N_4182);
nand U6291 (N_6291,N_2925,N_4527);
or U6292 (N_6292,N_4534,N_3687);
nor U6293 (N_6293,N_4426,N_2905);
and U6294 (N_6294,N_4542,N_4392);
xnor U6295 (N_6295,N_3505,N_2661);
xnor U6296 (N_6296,N_4767,N_3388);
and U6297 (N_6297,N_4855,N_4518);
or U6298 (N_6298,N_3257,N_3013);
or U6299 (N_6299,N_4169,N_3237);
nand U6300 (N_6300,N_3704,N_4172);
or U6301 (N_6301,N_3544,N_4982);
nor U6302 (N_6302,N_3933,N_3960);
nand U6303 (N_6303,N_3550,N_3071);
or U6304 (N_6304,N_2963,N_4625);
and U6305 (N_6305,N_3114,N_3101);
and U6306 (N_6306,N_4770,N_4595);
or U6307 (N_6307,N_3167,N_3871);
and U6308 (N_6308,N_3668,N_3888);
nand U6309 (N_6309,N_3664,N_3201);
nand U6310 (N_6310,N_4740,N_3215);
xor U6311 (N_6311,N_4647,N_4735);
or U6312 (N_6312,N_4432,N_4103);
or U6313 (N_6313,N_3085,N_4095);
or U6314 (N_6314,N_4380,N_4314);
xor U6315 (N_6315,N_3797,N_4771);
and U6316 (N_6316,N_3192,N_4634);
and U6317 (N_6317,N_2860,N_4549);
or U6318 (N_6318,N_3501,N_2918);
or U6319 (N_6319,N_3430,N_4051);
xnor U6320 (N_6320,N_3028,N_3635);
nor U6321 (N_6321,N_3521,N_3981);
nor U6322 (N_6322,N_3521,N_4822);
or U6323 (N_6323,N_4830,N_3534);
and U6324 (N_6324,N_2813,N_2725);
and U6325 (N_6325,N_3700,N_4306);
nor U6326 (N_6326,N_2623,N_2507);
and U6327 (N_6327,N_2604,N_3391);
nor U6328 (N_6328,N_2926,N_4010);
and U6329 (N_6329,N_3001,N_3578);
and U6330 (N_6330,N_4695,N_4002);
or U6331 (N_6331,N_3868,N_3944);
nor U6332 (N_6332,N_4074,N_4857);
nor U6333 (N_6333,N_3370,N_2680);
and U6334 (N_6334,N_4013,N_4848);
nor U6335 (N_6335,N_3567,N_4155);
nor U6336 (N_6336,N_3452,N_2504);
nor U6337 (N_6337,N_4932,N_2510);
xor U6338 (N_6338,N_2712,N_3550);
xnor U6339 (N_6339,N_3620,N_3925);
xnor U6340 (N_6340,N_3564,N_3080);
nand U6341 (N_6341,N_2628,N_4479);
xnor U6342 (N_6342,N_2907,N_4855);
xor U6343 (N_6343,N_2774,N_2675);
or U6344 (N_6344,N_4792,N_4428);
or U6345 (N_6345,N_2657,N_4303);
or U6346 (N_6346,N_2835,N_4496);
xnor U6347 (N_6347,N_3881,N_2533);
or U6348 (N_6348,N_3179,N_3111);
nor U6349 (N_6349,N_4869,N_4189);
or U6350 (N_6350,N_2602,N_3608);
nor U6351 (N_6351,N_4857,N_3783);
xor U6352 (N_6352,N_3879,N_4436);
xnor U6353 (N_6353,N_4516,N_4654);
or U6354 (N_6354,N_4417,N_4526);
or U6355 (N_6355,N_3322,N_3124);
or U6356 (N_6356,N_2723,N_3834);
nor U6357 (N_6357,N_4303,N_4136);
xnor U6358 (N_6358,N_2660,N_4640);
nor U6359 (N_6359,N_3292,N_3795);
and U6360 (N_6360,N_3063,N_4284);
or U6361 (N_6361,N_3779,N_3818);
and U6362 (N_6362,N_4047,N_3529);
or U6363 (N_6363,N_3151,N_3910);
or U6364 (N_6364,N_4782,N_3407);
or U6365 (N_6365,N_4436,N_4613);
and U6366 (N_6366,N_3191,N_4627);
or U6367 (N_6367,N_4020,N_3468);
xnor U6368 (N_6368,N_4479,N_3964);
or U6369 (N_6369,N_4811,N_3945);
xnor U6370 (N_6370,N_3164,N_3020);
or U6371 (N_6371,N_4527,N_2822);
nand U6372 (N_6372,N_4095,N_4603);
and U6373 (N_6373,N_3471,N_4920);
or U6374 (N_6374,N_3705,N_4904);
nand U6375 (N_6375,N_4677,N_2923);
or U6376 (N_6376,N_3404,N_4889);
xor U6377 (N_6377,N_4977,N_3665);
xnor U6378 (N_6378,N_4307,N_4375);
nand U6379 (N_6379,N_4644,N_4403);
xor U6380 (N_6380,N_2963,N_3529);
nor U6381 (N_6381,N_3622,N_2693);
nand U6382 (N_6382,N_3084,N_3497);
nor U6383 (N_6383,N_3783,N_2829);
nand U6384 (N_6384,N_3776,N_2517);
and U6385 (N_6385,N_3961,N_3189);
and U6386 (N_6386,N_3519,N_4431);
nand U6387 (N_6387,N_4616,N_4685);
or U6388 (N_6388,N_2938,N_3926);
nor U6389 (N_6389,N_3516,N_4136);
and U6390 (N_6390,N_3046,N_4526);
or U6391 (N_6391,N_2913,N_3582);
nand U6392 (N_6392,N_4693,N_3339);
and U6393 (N_6393,N_4132,N_4516);
nand U6394 (N_6394,N_3806,N_3549);
and U6395 (N_6395,N_3079,N_3088);
and U6396 (N_6396,N_4786,N_2952);
nor U6397 (N_6397,N_3231,N_2807);
nand U6398 (N_6398,N_3488,N_3506);
nand U6399 (N_6399,N_4352,N_4739);
or U6400 (N_6400,N_3045,N_2803);
nand U6401 (N_6401,N_2657,N_4844);
or U6402 (N_6402,N_4762,N_4083);
and U6403 (N_6403,N_3189,N_3294);
or U6404 (N_6404,N_4810,N_3231);
and U6405 (N_6405,N_3439,N_4381);
xnor U6406 (N_6406,N_2649,N_3446);
xor U6407 (N_6407,N_3083,N_4075);
and U6408 (N_6408,N_4226,N_3835);
or U6409 (N_6409,N_3355,N_4464);
xnor U6410 (N_6410,N_4559,N_2725);
xnor U6411 (N_6411,N_2571,N_4700);
or U6412 (N_6412,N_4773,N_4079);
nand U6413 (N_6413,N_2675,N_3667);
nor U6414 (N_6414,N_2609,N_4991);
nand U6415 (N_6415,N_4988,N_4796);
nor U6416 (N_6416,N_4462,N_4786);
nand U6417 (N_6417,N_4119,N_4678);
or U6418 (N_6418,N_3929,N_4604);
or U6419 (N_6419,N_4143,N_3983);
nor U6420 (N_6420,N_4933,N_2651);
nand U6421 (N_6421,N_3411,N_2784);
or U6422 (N_6422,N_4869,N_3392);
nor U6423 (N_6423,N_3709,N_3599);
nand U6424 (N_6424,N_4575,N_3781);
xor U6425 (N_6425,N_4683,N_3939);
and U6426 (N_6426,N_4567,N_3300);
nor U6427 (N_6427,N_3103,N_3467);
or U6428 (N_6428,N_2573,N_3528);
or U6429 (N_6429,N_2768,N_3615);
and U6430 (N_6430,N_4577,N_2850);
and U6431 (N_6431,N_3775,N_2746);
nand U6432 (N_6432,N_3781,N_4340);
or U6433 (N_6433,N_2603,N_4500);
nor U6434 (N_6434,N_4169,N_3015);
xor U6435 (N_6435,N_2887,N_3693);
xor U6436 (N_6436,N_3733,N_3118);
xnor U6437 (N_6437,N_3130,N_2919);
nor U6438 (N_6438,N_3087,N_2875);
nor U6439 (N_6439,N_2667,N_4743);
nand U6440 (N_6440,N_2703,N_3379);
xor U6441 (N_6441,N_4327,N_3259);
nand U6442 (N_6442,N_4145,N_4770);
or U6443 (N_6443,N_3263,N_2552);
xor U6444 (N_6444,N_4670,N_3024);
nand U6445 (N_6445,N_4363,N_4932);
nor U6446 (N_6446,N_2664,N_2814);
and U6447 (N_6447,N_4025,N_3859);
nor U6448 (N_6448,N_2673,N_4048);
and U6449 (N_6449,N_4220,N_4913);
or U6450 (N_6450,N_3688,N_3655);
or U6451 (N_6451,N_4454,N_2643);
nand U6452 (N_6452,N_2539,N_3522);
xor U6453 (N_6453,N_4272,N_4034);
or U6454 (N_6454,N_3360,N_3257);
nor U6455 (N_6455,N_2656,N_3891);
or U6456 (N_6456,N_2527,N_4210);
xnor U6457 (N_6457,N_4976,N_4690);
xnor U6458 (N_6458,N_4238,N_4809);
or U6459 (N_6459,N_2754,N_2757);
or U6460 (N_6460,N_3498,N_4006);
nand U6461 (N_6461,N_2677,N_3910);
and U6462 (N_6462,N_3944,N_4890);
xnor U6463 (N_6463,N_4384,N_4443);
or U6464 (N_6464,N_3112,N_3674);
xnor U6465 (N_6465,N_2981,N_4124);
nand U6466 (N_6466,N_2800,N_3825);
and U6467 (N_6467,N_3356,N_3546);
nor U6468 (N_6468,N_3618,N_4895);
xnor U6469 (N_6469,N_4976,N_4688);
nor U6470 (N_6470,N_3816,N_4733);
xnor U6471 (N_6471,N_2635,N_4476);
and U6472 (N_6472,N_3108,N_4599);
nand U6473 (N_6473,N_3516,N_3249);
and U6474 (N_6474,N_4058,N_2543);
nor U6475 (N_6475,N_3579,N_3836);
xnor U6476 (N_6476,N_3493,N_4105);
nand U6477 (N_6477,N_2870,N_4900);
or U6478 (N_6478,N_3195,N_2645);
and U6479 (N_6479,N_3881,N_2681);
xor U6480 (N_6480,N_4963,N_2698);
nand U6481 (N_6481,N_4696,N_4484);
nor U6482 (N_6482,N_3011,N_3929);
and U6483 (N_6483,N_2560,N_3762);
nor U6484 (N_6484,N_4056,N_2789);
or U6485 (N_6485,N_4620,N_4628);
xnor U6486 (N_6486,N_4374,N_3491);
and U6487 (N_6487,N_4537,N_2803);
or U6488 (N_6488,N_2945,N_3510);
nor U6489 (N_6489,N_3236,N_3223);
or U6490 (N_6490,N_3063,N_3433);
xnor U6491 (N_6491,N_3203,N_4271);
nor U6492 (N_6492,N_3146,N_4538);
nand U6493 (N_6493,N_3106,N_4040);
nand U6494 (N_6494,N_3992,N_3576);
or U6495 (N_6495,N_3049,N_3814);
xnor U6496 (N_6496,N_4453,N_3141);
nand U6497 (N_6497,N_4669,N_2590);
nand U6498 (N_6498,N_3732,N_2933);
and U6499 (N_6499,N_3059,N_3037);
xor U6500 (N_6500,N_3018,N_4227);
and U6501 (N_6501,N_3544,N_3990);
xor U6502 (N_6502,N_4050,N_4556);
nor U6503 (N_6503,N_3967,N_3206);
and U6504 (N_6504,N_4481,N_3355);
and U6505 (N_6505,N_3060,N_3072);
and U6506 (N_6506,N_4264,N_2540);
or U6507 (N_6507,N_3336,N_4695);
nor U6508 (N_6508,N_4397,N_4314);
or U6509 (N_6509,N_2838,N_3036);
or U6510 (N_6510,N_2582,N_2771);
or U6511 (N_6511,N_3816,N_3067);
nor U6512 (N_6512,N_3863,N_2934);
nand U6513 (N_6513,N_4785,N_4858);
and U6514 (N_6514,N_4006,N_4506);
nor U6515 (N_6515,N_4138,N_3662);
and U6516 (N_6516,N_3216,N_3861);
or U6517 (N_6517,N_2932,N_3812);
or U6518 (N_6518,N_4461,N_3659);
nor U6519 (N_6519,N_4130,N_3347);
nand U6520 (N_6520,N_3915,N_3556);
and U6521 (N_6521,N_4712,N_3467);
nand U6522 (N_6522,N_2912,N_4470);
nand U6523 (N_6523,N_3254,N_3901);
nor U6524 (N_6524,N_4255,N_4901);
or U6525 (N_6525,N_2671,N_2921);
or U6526 (N_6526,N_3409,N_4503);
nand U6527 (N_6527,N_4948,N_4241);
xor U6528 (N_6528,N_2584,N_4325);
xnor U6529 (N_6529,N_4868,N_4691);
nor U6530 (N_6530,N_2535,N_4039);
or U6531 (N_6531,N_4312,N_3865);
xor U6532 (N_6532,N_4588,N_3517);
xor U6533 (N_6533,N_3760,N_3783);
nand U6534 (N_6534,N_4503,N_2570);
and U6535 (N_6535,N_2781,N_4912);
and U6536 (N_6536,N_4948,N_2571);
nand U6537 (N_6537,N_3276,N_3404);
xnor U6538 (N_6538,N_4391,N_4463);
nand U6539 (N_6539,N_3614,N_3040);
or U6540 (N_6540,N_4881,N_2817);
or U6541 (N_6541,N_2705,N_4896);
or U6542 (N_6542,N_3754,N_3405);
and U6543 (N_6543,N_4282,N_3678);
nand U6544 (N_6544,N_2515,N_4028);
nand U6545 (N_6545,N_4643,N_4071);
nand U6546 (N_6546,N_4643,N_4556);
nand U6547 (N_6547,N_4344,N_4424);
nand U6548 (N_6548,N_3337,N_4301);
or U6549 (N_6549,N_2680,N_4702);
and U6550 (N_6550,N_3784,N_4787);
nor U6551 (N_6551,N_3479,N_4779);
xor U6552 (N_6552,N_3616,N_4811);
or U6553 (N_6553,N_2587,N_2984);
or U6554 (N_6554,N_3797,N_2684);
or U6555 (N_6555,N_4035,N_3829);
nor U6556 (N_6556,N_4512,N_3691);
or U6557 (N_6557,N_4886,N_2514);
and U6558 (N_6558,N_2622,N_3174);
nand U6559 (N_6559,N_2734,N_3867);
or U6560 (N_6560,N_4638,N_3854);
and U6561 (N_6561,N_3527,N_4818);
nor U6562 (N_6562,N_2676,N_3980);
or U6563 (N_6563,N_3227,N_4376);
nor U6564 (N_6564,N_3536,N_2658);
and U6565 (N_6565,N_2951,N_3862);
nand U6566 (N_6566,N_3993,N_2916);
xor U6567 (N_6567,N_3241,N_4466);
or U6568 (N_6568,N_4223,N_3714);
and U6569 (N_6569,N_3708,N_2900);
xor U6570 (N_6570,N_4612,N_2860);
xor U6571 (N_6571,N_4760,N_4298);
xnor U6572 (N_6572,N_3654,N_4085);
nand U6573 (N_6573,N_2895,N_3940);
nand U6574 (N_6574,N_4343,N_3331);
and U6575 (N_6575,N_2815,N_3700);
nand U6576 (N_6576,N_4804,N_2716);
or U6577 (N_6577,N_2581,N_3391);
and U6578 (N_6578,N_2792,N_2539);
and U6579 (N_6579,N_3502,N_2694);
nand U6580 (N_6580,N_2590,N_2643);
nor U6581 (N_6581,N_3086,N_2810);
xor U6582 (N_6582,N_4002,N_3420);
nand U6583 (N_6583,N_2658,N_4142);
nor U6584 (N_6584,N_4155,N_4552);
nor U6585 (N_6585,N_4384,N_3587);
xor U6586 (N_6586,N_3753,N_4928);
nor U6587 (N_6587,N_3747,N_2528);
and U6588 (N_6588,N_4267,N_4800);
xnor U6589 (N_6589,N_2607,N_3809);
xor U6590 (N_6590,N_4730,N_2967);
xnor U6591 (N_6591,N_4453,N_3934);
or U6592 (N_6592,N_4878,N_4387);
nor U6593 (N_6593,N_3927,N_3883);
nor U6594 (N_6594,N_3174,N_3726);
or U6595 (N_6595,N_3671,N_2546);
xor U6596 (N_6596,N_3216,N_4347);
or U6597 (N_6597,N_2965,N_3019);
nor U6598 (N_6598,N_3258,N_3316);
and U6599 (N_6599,N_4769,N_2555);
or U6600 (N_6600,N_3568,N_3036);
or U6601 (N_6601,N_3764,N_3815);
xor U6602 (N_6602,N_4250,N_4438);
xor U6603 (N_6603,N_4223,N_3239);
and U6604 (N_6604,N_2610,N_4520);
nor U6605 (N_6605,N_4082,N_2721);
and U6606 (N_6606,N_4918,N_3853);
nor U6607 (N_6607,N_4016,N_3469);
xor U6608 (N_6608,N_2855,N_4488);
nand U6609 (N_6609,N_4774,N_3670);
nand U6610 (N_6610,N_3559,N_3871);
nor U6611 (N_6611,N_3538,N_3593);
xnor U6612 (N_6612,N_4822,N_2984);
nor U6613 (N_6613,N_3164,N_4942);
or U6614 (N_6614,N_3691,N_4730);
xnor U6615 (N_6615,N_3091,N_4824);
nand U6616 (N_6616,N_4301,N_4431);
xor U6617 (N_6617,N_2691,N_4480);
or U6618 (N_6618,N_4798,N_2775);
or U6619 (N_6619,N_4260,N_2720);
nand U6620 (N_6620,N_4001,N_4041);
xnor U6621 (N_6621,N_3341,N_4079);
and U6622 (N_6622,N_3958,N_4985);
nand U6623 (N_6623,N_3524,N_4374);
nand U6624 (N_6624,N_2943,N_3156);
nor U6625 (N_6625,N_4736,N_3846);
and U6626 (N_6626,N_4677,N_3783);
and U6627 (N_6627,N_3477,N_4750);
and U6628 (N_6628,N_2541,N_2984);
xnor U6629 (N_6629,N_4672,N_4099);
or U6630 (N_6630,N_4393,N_4907);
nor U6631 (N_6631,N_3930,N_4578);
nor U6632 (N_6632,N_2761,N_4789);
nor U6633 (N_6633,N_3353,N_2663);
nor U6634 (N_6634,N_4345,N_2810);
and U6635 (N_6635,N_4928,N_3672);
and U6636 (N_6636,N_3401,N_3711);
or U6637 (N_6637,N_4222,N_3314);
and U6638 (N_6638,N_2623,N_3794);
nor U6639 (N_6639,N_4270,N_3253);
nor U6640 (N_6640,N_3473,N_4098);
and U6641 (N_6641,N_3666,N_3787);
nand U6642 (N_6642,N_2874,N_2534);
and U6643 (N_6643,N_3856,N_4387);
or U6644 (N_6644,N_4613,N_4830);
xnor U6645 (N_6645,N_2968,N_3362);
nor U6646 (N_6646,N_4534,N_3456);
nand U6647 (N_6647,N_3373,N_4855);
xnor U6648 (N_6648,N_4402,N_3127);
xnor U6649 (N_6649,N_3449,N_3141);
nand U6650 (N_6650,N_4880,N_2795);
or U6651 (N_6651,N_2596,N_3299);
xor U6652 (N_6652,N_3764,N_4540);
xnor U6653 (N_6653,N_3324,N_3382);
nand U6654 (N_6654,N_3710,N_4478);
xor U6655 (N_6655,N_3828,N_3426);
nor U6656 (N_6656,N_3790,N_3860);
nand U6657 (N_6657,N_3079,N_3117);
or U6658 (N_6658,N_4227,N_4685);
xnor U6659 (N_6659,N_2708,N_3869);
and U6660 (N_6660,N_3342,N_3263);
nor U6661 (N_6661,N_4651,N_3393);
nand U6662 (N_6662,N_2955,N_4279);
nand U6663 (N_6663,N_3980,N_4618);
nand U6664 (N_6664,N_2640,N_4388);
nand U6665 (N_6665,N_4527,N_3152);
nand U6666 (N_6666,N_3283,N_4206);
nor U6667 (N_6667,N_3948,N_3445);
and U6668 (N_6668,N_3973,N_3838);
and U6669 (N_6669,N_4270,N_4243);
xor U6670 (N_6670,N_4755,N_3727);
nand U6671 (N_6671,N_2947,N_3805);
xor U6672 (N_6672,N_4247,N_4306);
and U6673 (N_6673,N_4343,N_2939);
or U6674 (N_6674,N_2869,N_3949);
and U6675 (N_6675,N_4229,N_3825);
nor U6676 (N_6676,N_4389,N_3218);
xor U6677 (N_6677,N_4505,N_3190);
or U6678 (N_6678,N_4318,N_3821);
and U6679 (N_6679,N_3760,N_3676);
nor U6680 (N_6680,N_2951,N_3667);
nor U6681 (N_6681,N_3533,N_3895);
nor U6682 (N_6682,N_4178,N_4381);
xor U6683 (N_6683,N_4323,N_3530);
or U6684 (N_6684,N_2576,N_4536);
nand U6685 (N_6685,N_4470,N_3256);
and U6686 (N_6686,N_2787,N_4565);
and U6687 (N_6687,N_4620,N_4821);
nor U6688 (N_6688,N_3791,N_4084);
nand U6689 (N_6689,N_4890,N_4887);
xor U6690 (N_6690,N_4806,N_3054);
and U6691 (N_6691,N_4407,N_3034);
and U6692 (N_6692,N_3601,N_2873);
and U6693 (N_6693,N_2887,N_3688);
nand U6694 (N_6694,N_4987,N_4034);
and U6695 (N_6695,N_4933,N_2754);
or U6696 (N_6696,N_3971,N_4421);
and U6697 (N_6697,N_4058,N_3118);
nor U6698 (N_6698,N_2965,N_4983);
and U6699 (N_6699,N_3231,N_2892);
nand U6700 (N_6700,N_3933,N_3893);
or U6701 (N_6701,N_4339,N_4144);
and U6702 (N_6702,N_2599,N_3636);
and U6703 (N_6703,N_3500,N_3387);
xnor U6704 (N_6704,N_4366,N_4471);
nand U6705 (N_6705,N_4518,N_2774);
xor U6706 (N_6706,N_4734,N_3211);
nor U6707 (N_6707,N_4479,N_4830);
nand U6708 (N_6708,N_3083,N_4581);
nand U6709 (N_6709,N_2646,N_4988);
or U6710 (N_6710,N_2737,N_4203);
and U6711 (N_6711,N_3070,N_3001);
nand U6712 (N_6712,N_4145,N_4098);
or U6713 (N_6713,N_4464,N_3322);
nand U6714 (N_6714,N_3029,N_3231);
nand U6715 (N_6715,N_4431,N_4475);
nor U6716 (N_6716,N_3067,N_4565);
or U6717 (N_6717,N_4561,N_3328);
and U6718 (N_6718,N_2996,N_3636);
or U6719 (N_6719,N_3122,N_4372);
nand U6720 (N_6720,N_4361,N_3897);
nor U6721 (N_6721,N_3616,N_3303);
or U6722 (N_6722,N_3397,N_3071);
nand U6723 (N_6723,N_4981,N_2573);
nor U6724 (N_6724,N_3832,N_4653);
nor U6725 (N_6725,N_3424,N_3274);
or U6726 (N_6726,N_3806,N_4448);
nor U6727 (N_6727,N_3972,N_2979);
nor U6728 (N_6728,N_4045,N_2890);
or U6729 (N_6729,N_4642,N_2988);
nand U6730 (N_6730,N_4582,N_4892);
or U6731 (N_6731,N_2736,N_3411);
and U6732 (N_6732,N_4105,N_3876);
nor U6733 (N_6733,N_4267,N_3442);
or U6734 (N_6734,N_4006,N_3310);
xor U6735 (N_6735,N_3139,N_4912);
xor U6736 (N_6736,N_4861,N_3776);
and U6737 (N_6737,N_3047,N_4499);
and U6738 (N_6738,N_4605,N_4975);
and U6739 (N_6739,N_3819,N_4753);
nor U6740 (N_6740,N_3217,N_4276);
nor U6741 (N_6741,N_4734,N_3962);
or U6742 (N_6742,N_4933,N_4651);
or U6743 (N_6743,N_4484,N_2827);
nand U6744 (N_6744,N_3551,N_4949);
and U6745 (N_6745,N_2527,N_2644);
nor U6746 (N_6746,N_4449,N_3890);
nand U6747 (N_6747,N_3256,N_3291);
nand U6748 (N_6748,N_4315,N_3211);
or U6749 (N_6749,N_2765,N_4062);
nand U6750 (N_6750,N_2949,N_4433);
and U6751 (N_6751,N_3316,N_3478);
nand U6752 (N_6752,N_2620,N_3343);
nand U6753 (N_6753,N_4762,N_3698);
and U6754 (N_6754,N_4793,N_3221);
nand U6755 (N_6755,N_2572,N_4968);
nand U6756 (N_6756,N_3518,N_2591);
and U6757 (N_6757,N_3415,N_3480);
nand U6758 (N_6758,N_2663,N_3437);
nor U6759 (N_6759,N_2951,N_3783);
xor U6760 (N_6760,N_2768,N_2549);
nor U6761 (N_6761,N_2954,N_3595);
nor U6762 (N_6762,N_4517,N_3623);
xor U6763 (N_6763,N_3715,N_4499);
nor U6764 (N_6764,N_2596,N_2513);
nor U6765 (N_6765,N_3777,N_4275);
nand U6766 (N_6766,N_3839,N_2518);
and U6767 (N_6767,N_4905,N_2508);
xor U6768 (N_6768,N_4953,N_3154);
nand U6769 (N_6769,N_2832,N_3579);
or U6770 (N_6770,N_4855,N_3730);
and U6771 (N_6771,N_3323,N_4317);
or U6772 (N_6772,N_3444,N_2987);
nand U6773 (N_6773,N_2962,N_3113);
nand U6774 (N_6774,N_4289,N_4927);
nor U6775 (N_6775,N_3974,N_2782);
xor U6776 (N_6776,N_3868,N_2769);
nand U6777 (N_6777,N_3531,N_2531);
nor U6778 (N_6778,N_3629,N_3071);
xnor U6779 (N_6779,N_2903,N_4998);
xor U6780 (N_6780,N_2841,N_4829);
or U6781 (N_6781,N_2585,N_4249);
xnor U6782 (N_6782,N_3516,N_4787);
nor U6783 (N_6783,N_4863,N_4109);
xor U6784 (N_6784,N_3653,N_4274);
or U6785 (N_6785,N_2586,N_3002);
and U6786 (N_6786,N_2787,N_3030);
nand U6787 (N_6787,N_4066,N_3861);
or U6788 (N_6788,N_4200,N_2865);
and U6789 (N_6789,N_3743,N_2586);
and U6790 (N_6790,N_2844,N_3671);
nand U6791 (N_6791,N_4233,N_4069);
and U6792 (N_6792,N_2619,N_3300);
nor U6793 (N_6793,N_3247,N_3527);
and U6794 (N_6794,N_4693,N_3328);
nand U6795 (N_6795,N_3357,N_4572);
nor U6796 (N_6796,N_3357,N_4467);
nand U6797 (N_6797,N_3446,N_3027);
xnor U6798 (N_6798,N_4468,N_4590);
and U6799 (N_6799,N_4015,N_4595);
or U6800 (N_6800,N_3030,N_2619);
and U6801 (N_6801,N_4658,N_4301);
nor U6802 (N_6802,N_4205,N_3084);
and U6803 (N_6803,N_2837,N_3412);
nand U6804 (N_6804,N_2594,N_2835);
nor U6805 (N_6805,N_3494,N_4639);
xor U6806 (N_6806,N_4500,N_4331);
nand U6807 (N_6807,N_4353,N_3468);
xor U6808 (N_6808,N_4377,N_4088);
nor U6809 (N_6809,N_2714,N_4245);
and U6810 (N_6810,N_3365,N_3675);
and U6811 (N_6811,N_3152,N_2906);
or U6812 (N_6812,N_3527,N_2545);
or U6813 (N_6813,N_3659,N_3464);
xor U6814 (N_6814,N_4713,N_4194);
nor U6815 (N_6815,N_3918,N_4027);
nor U6816 (N_6816,N_4537,N_4892);
or U6817 (N_6817,N_2670,N_3589);
nor U6818 (N_6818,N_4607,N_3520);
nor U6819 (N_6819,N_4433,N_4716);
xnor U6820 (N_6820,N_3789,N_3372);
nor U6821 (N_6821,N_3335,N_4594);
nand U6822 (N_6822,N_4722,N_3384);
or U6823 (N_6823,N_2661,N_3329);
xor U6824 (N_6824,N_3637,N_2787);
nand U6825 (N_6825,N_2783,N_3503);
and U6826 (N_6826,N_2526,N_2580);
nand U6827 (N_6827,N_3424,N_3912);
and U6828 (N_6828,N_3510,N_2900);
nor U6829 (N_6829,N_4471,N_3944);
or U6830 (N_6830,N_2805,N_4591);
nand U6831 (N_6831,N_4711,N_4390);
or U6832 (N_6832,N_3089,N_2903);
or U6833 (N_6833,N_3353,N_2988);
and U6834 (N_6834,N_3263,N_4319);
and U6835 (N_6835,N_3997,N_4873);
xor U6836 (N_6836,N_3981,N_4798);
and U6837 (N_6837,N_3133,N_4406);
xor U6838 (N_6838,N_3764,N_2771);
nor U6839 (N_6839,N_3138,N_4850);
or U6840 (N_6840,N_4152,N_4836);
or U6841 (N_6841,N_4933,N_4763);
and U6842 (N_6842,N_3886,N_3690);
xor U6843 (N_6843,N_3901,N_4118);
or U6844 (N_6844,N_4546,N_4930);
and U6845 (N_6845,N_3341,N_4426);
xor U6846 (N_6846,N_3215,N_3418);
nand U6847 (N_6847,N_3527,N_4175);
xor U6848 (N_6848,N_4421,N_3982);
or U6849 (N_6849,N_4365,N_3663);
nand U6850 (N_6850,N_3911,N_4112);
and U6851 (N_6851,N_2866,N_2859);
nor U6852 (N_6852,N_2745,N_3160);
and U6853 (N_6853,N_4304,N_4129);
nor U6854 (N_6854,N_4158,N_4085);
or U6855 (N_6855,N_3470,N_3716);
and U6856 (N_6856,N_2557,N_4386);
nand U6857 (N_6857,N_4526,N_4218);
and U6858 (N_6858,N_4388,N_4404);
nand U6859 (N_6859,N_2868,N_3624);
xor U6860 (N_6860,N_3340,N_3515);
xnor U6861 (N_6861,N_2832,N_2576);
xor U6862 (N_6862,N_2541,N_3800);
nor U6863 (N_6863,N_3301,N_4345);
and U6864 (N_6864,N_3292,N_3279);
or U6865 (N_6865,N_3807,N_4559);
nor U6866 (N_6866,N_2618,N_4754);
and U6867 (N_6867,N_3474,N_4287);
and U6868 (N_6868,N_2561,N_2879);
nor U6869 (N_6869,N_3433,N_3210);
and U6870 (N_6870,N_3545,N_2900);
nand U6871 (N_6871,N_3948,N_4677);
nor U6872 (N_6872,N_4374,N_3259);
xnor U6873 (N_6873,N_3262,N_4266);
and U6874 (N_6874,N_4779,N_4090);
or U6875 (N_6875,N_4267,N_4374);
or U6876 (N_6876,N_3202,N_4492);
nor U6877 (N_6877,N_4586,N_2701);
nand U6878 (N_6878,N_3724,N_2666);
or U6879 (N_6879,N_2977,N_4004);
or U6880 (N_6880,N_3592,N_3140);
xnor U6881 (N_6881,N_4835,N_4276);
or U6882 (N_6882,N_3934,N_4819);
nor U6883 (N_6883,N_3755,N_4209);
nor U6884 (N_6884,N_2876,N_4372);
and U6885 (N_6885,N_4542,N_4548);
and U6886 (N_6886,N_3982,N_4447);
and U6887 (N_6887,N_3133,N_3004);
and U6888 (N_6888,N_2998,N_3372);
nand U6889 (N_6889,N_4378,N_4789);
and U6890 (N_6890,N_4178,N_4351);
nor U6891 (N_6891,N_3839,N_2735);
xor U6892 (N_6892,N_4317,N_2723);
nand U6893 (N_6893,N_4398,N_3834);
nor U6894 (N_6894,N_4478,N_3885);
nand U6895 (N_6895,N_3167,N_4767);
nor U6896 (N_6896,N_3725,N_3456);
nor U6897 (N_6897,N_3243,N_3933);
xor U6898 (N_6898,N_4393,N_4611);
and U6899 (N_6899,N_3936,N_2632);
xor U6900 (N_6900,N_3532,N_2738);
nor U6901 (N_6901,N_4957,N_3198);
xnor U6902 (N_6902,N_2909,N_3360);
nor U6903 (N_6903,N_4094,N_4921);
or U6904 (N_6904,N_2958,N_3360);
nand U6905 (N_6905,N_3146,N_3929);
or U6906 (N_6906,N_4317,N_4291);
xor U6907 (N_6907,N_3940,N_3825);
nand U6908 (N_6908,N_3209,N_4611);
nor U6909 (N_6909,N_4740,N_3406);
nand U6910 (N_6910,N_2923,N_4128);
or U6911 (N_6911,N_3725,N_4013);
or U6912 (N_6912,N_2552,N_4312);
or U6913 (N_6913,N_3479,N_3422);
nor U6914 (N_6914,N_4413,N_2891);
nand U6915 (N_6915,N_3044,N_4187);
nand U6916 (N_6916,N_4845,N_4341);
nand U6917 (N_6917,N_4260,N_2569);
and U6918 (N_6918,N_3923,N_3862);
xnor U6919 (N_6919,N_4117,N_2881);
nor U6920 (N_6920,N_4157,N_3401);
nor U6921 (N_6921,N_4553,N_2562);
xnor U6922 (N_6922,N_4914,N_3964);
and U6923 (N_6923,N_3361,N_3024);
and U6924 (N_6924,N_3477,N_4864);
and U6925 (N_6925,N_4558,N_2602);
xnor U6926 (N_6926,N_4026,N_2969);
nand U6927 (N_6927,N_4384,N_3093);
nand U6928 (N_6928,N_3350,N_2542);
and U6929 (N_6929,N_4121,N_3373);
nand U6930 (N_6930,N_3968,N_4359);
xnor U6931 (N_6931,N_4799,N_4485);
and U6932 (N_6932,N_4828,N_3682);
xor U6933 (N_6933,N_3638,N_4507);
or U6934 (N_6934,N_2573,N_3796);
or U6935 (N_6935,N_3747,N_3065);
xnor U6936 (N_6936,N_3355,N_2825);
and U6937 (N_6937,N_3326,N_4477);
xor U6938 (N_6938,N_3374,N_4988);
or U6939 (N_6939,N_4342,N_4381);
and U6940 (N_6940,N_3363,N_2749);
or U6941 (N_6941,N_3431,N_4704);
nor U6942 (N_6942,N_2588,N_4171);
and U6943 (N_6943,N_3738,N_4316);
xnor U6944 (N_6944,N_3927,N_2539);
or U6945 (N_6945,N_2654,N_3818);
and U6946 (N_6946,N_4757,N_2595);
nand U6947 (N_6947,N_4723,N_4989);
nor U6948 (N_6948,N_3857,N_4016);
xnor U6949 (N_6949,N_3895,N_3511);
or U6950 (N_6950,N_4163,N_3287);
nor U6951 (N_6951,N_4591,N_3833);
nand U6952 (N_6952,N_3542,N_4138);
and U6953 (N_6953,N_4224,N_4075);
or U6954 (N_6954,N_4644,N_2870);
nor U6955 (N_6955,N_3165,N_4219);
nand U6956 (N_6956,N_4073,N_2776);
nor U6957 (N_6957,N_3556,N_4118);
or U6958 (N_6958,N_2855,N_3213);
or U6959 (N_6959,N_4827,N_3622);
nand U6960 (N_6960,N_3542,N_4867);
xnor U6961 (N_6961,N_3859,N_2878);
nor U6962 (N_6962,N_2569,N_4848);
xor U6963 (N_6963,N_4778,N_3525);
and U6964 (N_6964,N_2559,N_4555);
or U6965 (N_6965,N_2907,N_2708);
and U6966 (N_6966,N_4750,N_2957);
nor U6967 (N_6967,N_3840,N_3719);
or U6968 (N_6968,N_4900,N_4826);
and U6969 (N_6969,N_2922,N_2703);
xor U6970 (N_6970,N_4578,N_4061);
nor U6971 (N_6971,N_4758,N_3350);
or U6972 (N_6972,N_4821,N_4419);
nor U6973 (N_6973,N_4334,N_4452);
nor U6974 (N_6974,N_2717,N_4068);
and U6975 (N_6975,N_4086,N_2887);
or U6976 (N_6976,N_3078,N_3914);
nand U6977 (N_6977,N_3961,N_2726);
xor U6978 (N_6978,N_3272,N_3247);
or U6979 (N_6979,N_2763,N_4531);
nand U6980 (N_6980,N_4489,N_4931);
or U6981 (N_6981,N_2823,N_4161);
xor U6982 (N_6982,N_3923,N_3201);
xnor U6983 (N_6983,N_3500,N_3723);
xor U6984 (N_6984,N_3367,N_3068);
nand U6985 (N_6985,N_4914,N_4157);
xnor U6986 (N_6986,N_3669,N_3271);
and U6987 (N_6987,N_4689,N_3791);
nor U6988 (N_6988,N_4855,N_4093);
nor U6989 (N_6989,N_3386,N_4522);
or U6990 (N_6990,N_3258,N_4118);
nand U6991 (N_6991,N_4786,N_4783);
or U6992 (N_6992,N_4697,N_4269);
nand U6993 (N_6993,N_4653,N_3538);
and U6994 (N_6994,N_3775,N_4379);
and U6995 (N_6995,N_4069,N_4517);
nand U6996 (N_6996,N_3098,N_3742);
and U6997 (N_6997,N_4261,N_4249);
nand U6998 (N_6998,N_3742,N_4414);
and U6999 (N_6999,N_4413,N_4981);
nor U7000 (N_7000,N_4279,N_2852);
nand U7001 (N_7001,N_3340,N_3636);
nand U7002 (N_7002,N_4595,N_3509);
nor U7003 (N_7003,N_4064,N_4733);
and U7004 (N_7004,N_2947,N_3377);
nor U7005 (N_7005,N_4365,N_3248);
nor U7006 (N_7006,N_2562,N_2823);
xnor U7007 (N_7007,N_3066,N_2777);
nand U7008 (N_7008,N_4809,N_4340);
or U7009 (N_7009,N_4945,N_2969);
xor U7010 (N_7010,N_4654,N_3571);
xnor U7011 (N_7011,N_4563,N_3931);
and U7012 (N_7012,N_2538,N_3281);
or U7013 (N_7013,N_4620,N_4566);
nor U7014 (N_7014,N_3476,N_2796);
or U7015 (N_7015,N_3333,N_2866);
xnor U7016 (N_7016,N_3557,N_4855);
or U7017 (N_7017,N_3237,N_4502);
or U7018 (N_7018,N_4935,N_2939);
nand U7019 (N_7019,N_3962,N_3355);
nand U7020 (N_7020,N_3298,N_2655);
nand U7021 (N_7021,N_3077,N_3822);
nor U7022 (N_7022,N_3760,N_2689);
or U7023 (N_7023,N_3295,N_4757);
nor U7024 (N_7024,N_4587,N_4989);
xor U7025 (N_7025,N_4632,N_3319);
and U7026 (N_7026,N_4264,N_2752);
and U7027 (N_7027,N_4357,N_3117);
nand U7028 (N_7028,N_3568,N_3154);
nand U7029 (N_7029,N_3589,N_2628);
nand U7030 (N_7030,N_3988,N_3824);
nand U7031 (N_7031,N_4611,N_2566);
nor U7032 (N_7032,N_3484,N_4463);
nor U7033 (N_7033,N_3966,N_4469);
nor U7034 (N_7034,N_4287,N_4040);
nand U7035 (N_7035,N_2543,N_2856);
nor U7036 (N_7036,N_3868,N_4054);
or U7037 (N_7037,N_3277,N_4664);
xor U7038 (N_7038,N_2602,N_2840);
nor U7039 (N_7039,N_3148,N_3700);
nor U7040 (N_7040,N_3304,N_2782);
and U7041 (N_7041,N_3283,N_3993);
and U7042 (N_7042,N_2735,N_4510);
and U7043 (N_7043,N_2543,N_3002);
nor U7044 (N_7044,N_2514,N_4683);
nor U7045 (N_7045,N_4855,N_2871);
and U7046 (N_7046,N_4412,N_3765);
or U7047 (N_7047,N_4944,N_4838);
xnor U7048 (N_7048,N_3105,N_3437);
nand U7049 (N_7049,N_3579,N_4439);
nor U7050 (N_7050,N_3655,N_4154);
xnor U7051 (N_7051,N_3712,N_4038);
nand U7052 (N_7052,N_4507,N_3310);
xnor U7053 (N_7053,N_2577,N_2839);
nor U7054 (N_7054,N_3767,N_2836);
or U7055 (N_7055,N_4410,N_2802);
nor U7056 (N_7056,N_4040,N_4127);
nor U7057 (N_7057,N_3979,N_4439);
nand U7058 (N_7058,N_2639,N_2739);
and U7059 (N_7059,N_3156,N_3101);
nand U7060 (N_7060,N_4980,N_3233);
and U7061 (N_7061,N_3112,N_2872);
nor U7062 (N_7062,N_3721,N_4311);
nor U7063 (N_7063,N_4523,N_4395);
xnor U7064 (N_7064,N_2817,N_4562);
nand U7065 (N_7065,N_3819,N_4098);
nand U7066 (N_7066,N_3962,N_4207);
nor U7067 (N_7067,N_3407,N_3909);
and U7068 (N_7068,N_2640,N_2829);
nand U7069 (N_7069,N_4800,N_3860);
and U7070 (N_7070,N_3205,N_3152);
nor U7071 (N_7071,N_4949,N_3809);
xnor U7072 (N_7072,N_4619,N_4244);
and U7073 (N_7073,N_4528,N_3052);
or U7074 (N_7074,N_4413,N_4491);
and U7075 (N_7075,N_4291,N_2789);
or U7076 (N_7076,N_2546,N_2896);
nor U7077 (N_7077,N_3611,N_3563);
and U7078 (N_7078,N_2880,N_2988);
nor U7079 (N_7079,N_4476,N_3167);
nor U7080 (N_7080,N_2832,N_2735);
nand U7081 (N_7081,N_3594,N_2665);
and U7082 (N_7082,N_3223,N_3120);
or U7083 (N_7083,N_3951,N_4461);
xor U7084 (N_7084,N_2944,N_3085);
or U7085 (N_7085,N_4346,N_3572);
nand U7086 (N_7086,N_4428,N_4074);
nand U7087 (N_7087,N_3952,N_3881);
nor U7088 (N_7088,N_3561,N_4386);
or U7089 (N_7089,N_4816,N_2606);
xor U7090 (N_7090,N_2683,N_2685);
or U7091 (N_7091,N_4792,N_2830);
nand U7092 (N_7092,N_3825,N_4913);
or U7093 (N_7093,N_3446,N_2773);
and U7094 (N_7094,N_3662,N_4241);
nor U7095 (N_7095,N_3936,N_3044);
and U7096 (N_7096,N_4128,N_3663);
nand U7097 (N_7097,N_4059,N_4422);
or U7098 (N_7098,N_3364,N_4338);
nand U7099 (N_7099,N_3389,N_3638);
xor U7100 (N_7100,N_3116,N_4732);
nor U7101 (N_7101,N_2544,N_4697);
nor U7102 (N_7102,N_2587,N_2642);
nand U7103 (N_7103,N_3357,N_4543);
and U7104 (N_7104,N_4583,N_3215);
and U7105 (N_7105,N_4763,N_3586);
xnor U7106 (N_7106,N_4839,N_4820);
and U7107 (N_7107,N_3718,N_2536);
nor U7108 (N_7108,N_3260,N_2507);
nand U7109 (N_7109,N_3817,N_4480);
nand U7110 (N_7110,N_3342,N_2688);
or U7111 (N_7111,N_3945,N_4040);
nor U7112 (N_7112,N_3109,N_3166);
and U7113 (N_7113,N_3676,N_4163);
nand U7114 (N_7114,N_4395,N_2544);
nand U7115 (N_7115,N_2833,N_4546);
nor U7116 (N_7116,N_3470,N_3717);
nor U7117 (N_7117,N_3773,N_3741);
nor U7118 (N_7118,N_4068,N_3782);
xnor U7119 (N_7119,N_4265,N_4946);
and U7120 (N_7120,N_2973,N_4557);
or U7121 (N_7121,N_2687,N_3941);
xor U7122 (N_7122,N_4854,N_4451);
nand U7123 (N_7123,N_3473,N_3008);
or U7124 (N_7124,N_3950,N_4356);
xnor U7125 (N_7125,N_3355,N_2841);
nor U7126 (N_7126,N_3147,N_4045);
nand U7127 (N_7127,N_4682,N_4410);
and U7128 (N_7128,N_4284,N_4797);
nor U7129 (N_7129,N_3861,N_3007);
xor U7130 (N_7130,N_3207,N_4575);
xnor U7131 (N_7131,N_4173,N_2908);
or U7132 (N_7132,N_3689,N_3478);
and U7133 (N_7133,N_2813,N_4184);
xor U7134 (N_7134,N_3058,N_3470);
xnor U7135 (N_7135,N_2670,N_3872);
nand U7136 (N_7136,N_4760,N_3795);
xor U7137 (N_7137,N_2806,N_3828);
and U7138 (N_7138,N_4118,N_4514);
nand U7139 (N_7139,N_3725,N_4316);
nor U7140 (N_7140,N_3845,N_4996);
and U7141 (N_7141,N_3543,N_2981);
or U7142 (N_7142,N_3498,N_4928);
or U7143 (N_7143,N_3809,N_3975);
or U7144 (N_7144,N_2767,N_3577);
nor U7145 (N_7145,N_2909,N_3326);
xnor U7146 (N_7146,N_4722,N_3210);
nor U7147 (N_7147,N_4241,N_4881);
nand U7148 (N_7148,N_4970,N_3524);
nand U7149 (N_7149,N_4433,N_3992);
or U7150 (N_7150,N_4900,N_2874);
nor U7151 (N_7151,N_4309,N_3306);
nor U7152 (N_7152,N_4905,N_3538);
nor U7153 (N_7153,N_3711,N_4355);
xor U7154 (N_7154,N_4518,N_3141);
and U7155 (N_7155,N_2929,N_4355);
and U7156 (N_7156,N_2544,N_3525);
xor U7157 (N_7157,N_4179,N_4563);
xor U7158 (N_7158,N_4560,N_2781);
nor U7159 (N_7159,N_2564,N_4933);
nand U7160 (N_7160,N_3642,N_3787);
nor U7161 (N_7161,N_4466,N_4843);
nor U7162 (N_7162,N_4453,N_4915);
nor U7163 (N_7163,N_2725,N_3396);
nor U7164 (N_7164,N_3933,N_3966);
xnor U7165 (N_7165,N_3856,N_2515);
nand U7166 (N_7166,N_4955,N_2527);
nor U7167 (N_7167,N_3189,N_2503);
or U7168 (N_7168,N_2834,N_4479);
and U7169 (N_7169,N_3286,N_2759);
xor U7170 (N_7170,N_3969,N_3197);
or U7171 (N_7171,N_4585,N_3337);
or U7172 (N_7172,N_4259,N_4209);
and U7173 (N_7173,N_4984,N_4777);
nor U7174 (N_7174,N_2762,N_4220);
and U7175 (N_7175,N_3320,N_4248);
nand U7176 (N_7176,N_2762,N_3778);
or U7177 (N_7177,N_3984,N_4639);
and U7178 (N_7178,N_2917,N_3091);
xor U7179 (N_7179,N_4741,N_4867);
nand U7180 (N_7180,N_4963,N_2839);
and U7181 (N_7181,N_4794,N_3431);
nor U7182 (N_7182,N_3906,N_4387);
nor U7183 (N_7183,N_2573,N_3062);
xnor U7184 (N_7184,N_4188,N_4699);
xor U7185 (N_7185,N_3829,N_3026);
xor U7186 (N_7186,N_4798,N_4038);
or U7187 (N_7187,N_3209,N_3098);
nand U7188 (N_7188,N_2991,N_3858);
nand U7189 (N_7189,N_3446,N_2545);
xnor U7190 (N_7190,N_3760,N_3984);
nor U7191 (N_7191,N_2974,N_3997);
xor U7192 (N_7192,N_2995,N_3379);
and U7193 (N_7193,N_3817,N_4663);
and U7194 (N_7194,N_3092,N_3063);
and U7195 (N_7195,N_3047,N_3055);
nor U7196 (N_7196,N_3449,N_3158);
and U7197 (N_7197,N_3296,N_2618);
nand U7198 (N_7198,N_4159,N_4881);
or U7199 (N_7199,N_4251,N_4559);
xor U7200 (N_7200,N_2607,N_2582);
nor U7201 (N_7201,N_3977,N_4808);
nor U7202 (N_7202,N_3744,N_4850);
xor U7203 (N_7203,N_3162,N_3525);
and U7204 (N_7204,N_2811,N_4043);
nor U7205 (N_7205,N_3914,N_4694);
nor U7206 (N_7206,N_4292,N_2730);
nor U7207 (N_7207,N_2991,N_3656);
xnor U7208 (N_7208,N_3784,N_3840);
nor U7209 (N_7209,N_4228,N_4911);
nand U7210 (N_7210,N_3786,N_3531);
xnor U7211 (N_7211,N_4439,N_4793);
nand U7212 (N_7212,N_3835,N_3386);
and U7213 (N_7213,N_4031,N_2608);
xnor U7214 (N_7214,N_3100,N_4387);
xor U7215 (N_7215,N_2652,N_2843);
or U7216 (N_7216,N_2654,N_4562);
and U7217 (N_7217,N_3971,N_4610);
nand U7218 (N_7218,N_4858,N_3119);
and U7219 (N_7219,N_4262,N_3059);
xnor U7220 (N_7220,N_2980,N_2833);
nor U7221 (N_7221,N_3869,N_3914);
nand U7222 (N_7222,N_4061,N_2522);
or U7223 (N_7223,N_2813,N_4148);
or U7224 (N_7224,N_2697,N_2817);
nor U7225 (N_7225,N_4940,N_3132);
and U7226 (N_7226,N_2534,N_2759);
and U7227 (N_7227,N_3040,N_2502);
nand U7228 (N_7228,N_3626,N_3490);
xnor U7229 (N_7229,N_3951,N_4655);
nor U7230 (N_7230,N_3960,N_4774);
nor U7231 (N_7231,N_3674,N_3414);
and U7232 (N_7232,N_4788,N_2751);
nand U7233 (N_7233,N_4603,N_2522);
or U7234 (N_7234,N_4960,N_4050);
nor U7235 (N_7235,N_2701,N_4462);
or U7236 (N_7236,N_4895,N_3900);
xor U7237 (N_7237,N_2852,N_3376);
nand U7238 (N_7238,N_3940,N_4050);
nand U7239 (N_7239,N_4971,N_3579);
and U7240 (N_7240,N_3644,N_3655);
nor U7241 (N_7241,N_3914,N_3694);
nand U7242 (N_7242,N_4169,N_2962);
or U7243 (N_7243,N_3611,N_4743);
or U7244 (N_7244,N_3301,N_3934);
and U7245 (N_7245,N_3139,N_4520);
xor U7246 (N_7246,N_4726,N_4188);
nor U7247 (N_7247,N_2812,N_4053);
nor U7248 (N_7248,N_3265,N_4195);
nor U7249 (N_7249,N_3668,N_3903);
and U7250 (N_7250,N_3594,N_4755);
nand U7251 (N_7251,N_3386,N_4600);
and U7252 (N_7252,N_3548,N_4548);
and U7253 (N_7253,N_4804,N_2767);
nand U7254 (N_7254,N_4032,N_2663);
nand U7255 (N_7255,N_3212,N_2578);
nor U7256 (N_7256,N_3373,N_3455);
and U7257 (N_7257,N_2611,N_2756);
xnor U7258 (N_7258,N_4504,N_3481);
xnor U7259 (N_7259,N_3008,N_4556);
nor U7260 (N_7260,N_2552,N_4212);
xor U7261 (N_7261,N_4641,N_4189);
nand U7262 (N_7262,N_3179,N_3193);
nor U7263 (N_7263,N_3156,N_2820);
and U7264 (N_7264,N_4631,N_4439);
or U7265 (N_7265,N_3161,N_3343);
and U7266 (N_7266,N_3981,N_3749);
nor U7267 (N_7267,N_3134,N_3392);
xor U7268 (N_7268,N_4746,N_3728);
nor U7269 (N_7269,N_4209,N_4328);
or U7270 (N_7270,N_3128,N_4645);
nand U7271 (N_7271,N_4971,N_3192);
and U7272 (N_7272,N_4008,N_3509);
or U7273 (N_7273,N_2725,N_3436);
and U7274 (N_7274,N_4590,N_2812);
nand U7275 (N_7275,N_3111,N_4766);
xnor U7276 (N_7276,N_2590,N_2817);
nand U7277 (N_7277,N_4307,N_3183);
nor U7278 (N_7278,N_4831,N_3680);
nor U7279 (N_7279,N_3357,N_4606);
nand U7280 (N_7280,N_4334,N_4550);
xor U7281 (N_7281,N_2879,N_2824);
and U7282 (N_7282,N_3196,N_4672);
and U7283 (N_7283,N_3658,N_4390);
or U7284 (N_7284,N_2710,N_2839);
nand U7285 (N_7285,N_4494,N_3156);
or U7286 (N_7286,N_2682,N_4235);
nand U7287 (N_7287,N_3587,N_4174);
nor U7288 (N_7288,N_4683,N_4395);
nand U7289 (N_7289,N_2785,N_2841);
or U7290 (N_7290,N_4251,N_3568);
or U7291 (N_7291,N_4604,N_4008);
nor U7292 (N_7292,N_4441,N_2952);
nand U7293 (N_7293,N_3273,N_3249);
and U7294 (N_7294,N_3666,N_3539);
nor U7295 (N_7295,N_2890,N_3766);
or U7296 (N_7296,N_4262,N_4968);
or U7297 (N_7297,N_2890,N_4341);
or U7298 (N_7298,N_4447,N_3949);
or U7299 (N_7299,N_3429,N_3275);
xor U7300 (N_7300,N_3806,N_4396);
nor U7301 (N_7301,N_4665,N_4492);
nor U7302 (N_7302,N_3000,N_3320);
nor U7303 (N_7303,N_4869,N_2861);
nand U7304 (N_7304,N_3976,N_2575);
xor U7305 (N_7305,N_2999,N_4362);
xor U7306 (N_7306,N_4159,N_3358);
or U7307 (N_7307,N_3737,N_3180);
xor U7308 (N_7308,N_2928,N_3734);
nand U7309 (N_7309,N_3373,N_2899);
xnor U7310 (N_7310,N_4528,N_3196);
and U7311 (N_7311,N_2781,N_4106);
xnor U7312 (N_7312,N_2853,N_2709);
nand U7313 (N_7313,N_3101,N_4867);
xnor U7314 (N_7314,N_4734,N_4831);
nand U7315 (N_7315,N_2848,N_3838);
nor U7316 (N_7316,N_4587,N_3873);
xnor U7317 (N_7317,N_4700,N_3639);
or U7318 (N_7318,N_2889,N_4482);
or U7319 (N_7319,N_4459,N_2975);
nand U7320 (N_7320,N_4110,N_2927);
or U7321 (N_7321,N_2860,N_4459);
nor U7322 (N_7322,N_2697,N_2620);
or U7323 (N_7323,N_4368,N_3559);
nand U7324 (N_7324,N_3469,N_4161);
nand U7325 (N_7325,N_2563,N_2575);
nand U7326 (N_7326,N_3483,N_2585);
or U7327 (N_7327,N_3212,N_3269);
xnor U7328 (N_7328,N_4990,N_3453);
nor U7329 (N_7329,N_3991,N_2697);
nand U7330 (N_7330,N_3844,N_4984);
xor U7331 (N_7331,N_4521,N_2884);
xor U7332 (N_7332,N_3651,N_4315);
nand U7333 (N_7333,N_3118,N_3259);
nor U7334 (N_7334,N_3663,N_3799);
and U7335 (N_7335,N_4539,N_3393);
xnor U7336 (N_7336,N_4115,N_3327);
xor U7337 (N_7337,N_4614,N_3388);
nand U7338 (N_7338,N_2531,N_2635);
or U7339 (N_7339,N_3463,N_3283);
nor U7340 (N_7340,N_4368,N_2769);
or U7341 (N_7341,N_4523,N_3007);
and U7342 (N_7342,N_3444,N_4865);
xnor U7343 (N_7343,N_4181,N_2883);
xor U7344 (N_7344,N_3784,N_4188);
nand U7345 (N_7345,N_2698,N_4939);
xor U7346 (N_7346,N_2829,N_4287);
xor U7347 (N_7347,N_3320,N_4893);
and U7348 (N_7348,N_4393,N_3728);
or U7349 (N_7349,N_2835,N_4489);
nor U7350 (N_7350,N_4313,N_3288);
nand U7351 (N_7351,N_4391,N_3024);
nand U7352 (N_7352,N_4676,N_3565);
or U7353 (N_7353,N_3165,N_3716);
nand U7354 (N_7354,N_4247,N_3076);
nor U7355 (N_7355,N_3991,N_2969);
nand U7356 (N_7356,N_2535,N_3212);
nand U7357 (N_7357,N_4226,N_3831);
or U7358 (N_7358,N_4590,N_4863);
or U7359 (N_7359,N_4090,N_2516);
or U7360 (N_7360,N_3478,N_4854);
and U7361 (N_7361,N_4297,N_4312);
or U7362 (N_7362,N_2598,N_4108);
xor U7363 (N_7363,N_2897,N_3370);
xnor U7364 (N_7364,N_2834,N_4408);
nand U7365 (N_7365,N_3799,N_3153);
or U7366 (N_7366,N_4619,N_3795);
or U7367 (N_7367,N_3239,N_4667);
xor U7368 (N_7368,N_3638,N_3297);
or U7369 (N_7369,N_3435,N_4015);
or U7370 (N_7370,N_2863,N_2875);
xor U7371 (N_7371,N_3325,N_3668);
xor U7372 (N_7372,N_3736,N_4596);
nor U7373 (N_7373,N_4991,N_3238);
xor U7374 (N_7374,N_3705,N_3692);
nor U7375 (N_7375,N_4217,N_2937);
nand U7376 (N_7376,N_3245,N_3905);
or U7377 (N_7377,N_2851,N_4454);
nor U7378 (N_7378,N_2642,N_3506);
and U7379 (N_7379,N_3506,N_3496);
xor U7380 (N_7380,N_4790,N_3772);
xnor U7381 (N_7381,N_4352,N_4346);
xnor U7382 (N_7382,N_2516,N_4932);
nor U7383 (N_7383,N_3711,N_3347);
and U7384 (N_7384,N_3330,N_4306);
and U7385 (N_7385,N_4325,N_3467);
xor U7386 (N_7386,N_3526,N_3065);
xor U7387 (N_7387,N_3426,N_2607);
nor U7388 (N_7388,N_2700,N_3093);
nand U7389 (N_7389,N_2830,N_4027);
nor U7390 (N_7390,N_2996,N_3367);
nor U7391 (N_7391,N_4011,N_4423);
and U7392 (N_7392,N_3139,N_3563);
or U7393 (N_7393,N_4196,N_3682);
nor U7394 (N_7394,N_3378,N_4026);
nor U7395 (N_7395,N_3308,N_4112);
or U7396 (N_7396,N_4113,N_3388);
nor U7397 (N_7397,N_2536,N_3956);
and U7398 (N_7398,N_3829,N_4012);
and U7399 (N_7399,N_2988,N_3006);
or U7400 (N_7400,N_3480,N_3537);
xnor U7401 (N_7401,N_4750,N_4675);
and U7402 (N_7402,N_4607,N_3314);
and U7403 (N_7403,N_2821,N_4993);
or U7404 (N_7404,N_3313,N_3590);
xnor U7405 (N_7405,N_2655,N_4827);
nor U7406 (N_7406,N_3451,N_4460);
nand U7407 (N_7407,N_3837,N_4625);
nand U7408 (N_7408,N_4346,N_4689);
nand U7409 (N_7409,N_4114,N_4726);
or U7410 (N_7410,N_4267,N_2528);
nor U7411 (N_7411,N_3493,N_4050);
or U7412 (N_7412,N_4342,N_4822);
nor U7413 (N_7413,N_3744,N_4491);
nand U7414 (N_7414,N_4374,N_3482);
nand U7415 (N_7415,N_4844,N_3429);
nor U7416 (N_7416,N_2616,N_4252);
or U7417 (N_7417,N_2913,N_3496);
or U7418 (N_7418,N_2978,N_2839);
nor U7419 (N_7419,N_3517,N_3349);
xnor U7420 (N_7420,N_3400,N_3500);
xor U7421 (N_7421,N_4534,N_3186);
and U7422 (N_7422,N_3380,N_3213);
or U7423 (N_7423,N_4223,N_4460);
nand U7424 (N_7424,N_2582,N_4810);
and U7425 (N_7425,N_3063,N_4303);
nand U7426 (N_7426,N_3635,N_3985);
nor U7427 (N_7427,N_4455,N_3061);
or U7428 (N_7428,N_4219,N_3823);
xor U7429 (N_7429,N_3560,N_3609);
nor U7430 (N_7430,N_4797,N_2657);
and U7431 (N_7431,N_4337,N_2938);
nor U7432 (N_7432,N_3738,N_2882);
or U7433 (N_7433,N_4560,N_3125);
or U7434 (N_7434,N_3031,N_4516);
nor U7435 (N_7435,N_3725,N_2957);
nor U7436 (N_7436,N_3522,N_4679);
xnor U7437 (N_7437,N_3142,N_3421);
nor U7438 (N_7438,N_3474,N_2506);
and U7439 (N_7439,N_4878,N_4893);
xor U7440 (N_7440,N_3348,N_2940);
nand U7441 (N_7441,N_3268,N_2843);
nor U7442 (N_7442,N_4169,N_4868);
and U7443 (N_7443,N_2562,N_3558);
and U7444 (N_7444,N_2606,N_4329);
nand U7445 (N_7445,N_3319,N_4505);
nand U7446 (N_7446,N_2893,N_2771);
or U7447 (N_7447,N_4162,N_4955);
and U7448 (N_7448,N_4664,N_3958);
nor U7449 (N_7449,N_4644,N_4308);
nand U7450 (N_7450,N_4587,N_3713);
xor U7451 (N_7451,N_3307,N_4074);
xor U7452 (N_7452,N_3544,N_2790);
or U7453 (N_7453,N_3598,N_3544);
and U7454 (N_7454,N_2638,N_3496);
nand U7455 (N_7455,N_4298,N_2899);
nand U7456 (N_7456,N_4570,N_3853);
xnor U7457 (N_7457,N_3207,N_4982);
nor U7458 (N_7458,N_3033,N_4764);
nand U7459 (N_7459,N_3619,N_3618);
nor U7460 (N_7460,N_4811,N_2970);
and U7461 (N_7461,N_4106,N_3272);
xor U7462 (N_7462,N_4002,N_3353);
nand U7463 (N_7463,N_3210,N_2601);
nand U7464 (N_7464,N_3023,N_3707);
nand U7465 (N_7465,N_4885,N_4510);
nor U7466 (N_7466,N_3401,N_2949);
nor U7467 (N_7467,N_4108,N_4756);
xor U7468 (N_7468,N_3455,N_4658);
nand U7469 (N_7469,N_3607,N_4467);
nand U7470 (N_7470,N_3696,N_4023);
or U7471 (N_7471,N_3832,N_4595);
and U7472 (N_7472,N_3610,N_3873);
xnor U7473 (N_7473,N_4175,N_2556);
xnor U7474 (N_7474,N_4532,N_3724);
and U7475 (N_7475,N_3525,N_2960);
and U7476 (N_7476,N_4706,N_4605);
xor U7477 (N_7477,N_4486,N_4266);
nor U7478 (N_7478,N_3096,N_3044);
nand U7479 (N_7479,N_3889,N_4064);
or U7480 (N_7480,N_4160,N_2904);
nand U7481 (N_7481,N_3646,N_3872);
or U7482 (N_7482,N_4088,N_2942);
nor U7483 (N_7483,N_4090,N_3651);
and U7484 (N_7484,N_4771,N_4927);
or U7485 (N_7485,N_4207,N_2997);
or U7486 (N_7486,N_3794,N_3443);
nor U7487 (N_7487,N_3118,N_4406);
and U7488 (N_7488,N_2977,N_4387);
or U7489 (N_7489,N_4057,N_3681);
xor U7490 (N_7490,N_2564,N_4593);
or U7491 (N_7491,N_2673,N_4964);
and U7492 (N_7492,N_3281,N_3570);
and U7493 (N_7493,N_4427,N_3610);
nand U7494 (N_7494,N_3787,N_3972);
or U7495 (N_7495,N_4994,N_3024);
and U7496 (N_7496,N_4539,N_2546);
or U7497 (N_7497,N_2734,N_4631);
nand U7498 (N_7498,N_4683,N_3325);
xor U7499 (N_7499,N_2577,N_4183);
or U7500 (N_7500,N_5335,N_5407);
and U7501 (N_7501,N_6253,N_5664);
and U7502 (N_7502,N_5550,N_5008);
xnor U7503 (N_7503,N_7356,N_6861);
or U7504 (N_7504,N_5054,N_7439);
nor U7505 (N_7505,N_5044,N_6358);
nor U7506 (N_7506,N_5046,N_5962);
xor U7507 (N_7507,N_5721,N_5117);
nand U7508 (N_7508,N_5801,N_5539);
and U7509 (N_7509,N_6950,N_5441);
xnor U7510 (N_7510,N_7264,N_6022);
nor U7511 (N_7511,N_5951,N_6138);
xnor U7512 (N_7512,N_7149,N_6657);
nand U7513 (N_7513,N_6038,N_5241);
xor U7514 (N_7514,N_5723,N_5905);
xnor U7515 (N_7515,N_5496,N_6574);
xnor U7516 (N_7516,N_5031,N_7066);
nor U7517 (N_7517,N_6202,N_6801);
or U7518 (N_7518,N_6651,N_7312);
or U7519 (N_7519,N_6374,N_6229);
nand U7520 (N_7520,N_5236,N_6147);
xor U7521 (N_7521,N_6916,N_5870);
and U7522 (N_7522,N_5457,N_5213);
nor U7523 (N_7523,N_6378,N_7123);
nand U7524 (N_7524,N_5903,N_6522);
xnor U7525 (N_7525,N_6430,N_5231);
nand U7526 (N_7526,N_6132,N_5463);
or U7527 (N_7527,N_5183,N_5377);
and U7528 (N_7528,N_5641,N_5010);
xnor U7529 (N_7529,N_5192,N_6653);
or U7530 (N_7530,N_5502,N_7459);
nor U7531 (N_7531,N_5177,N_6943);
xor U7532 (N_7532,N_5286,N_6967);
or U7533 (N_7533,N_6620,N_5255);
and U7534 (N_7534,N_6420,N_7395);
nand U7535 (N_7535,N_7404,N_7362);
nand U7536 (N_7536,N_5531,N_7406);
nor U7537 (N_7537,N_7304,N_5529);
or U7538 (N_7538,N_7478,N_5625);
and U7539 (N_7539,N_6163,N_5928);
nor U7540 (N_7540,N_5712,N_6600);
xor U7541 (N_7541,N_6592,N_5420);
nand U7542 (N_7542,N_6211,N_5799);
xor U7543 (N_7543,N_6447,N_7462);
or U7544 (N_7544,N_7030,N_5590);
xnor U7545 (N_7545,N_6051,N_7436);
xor U7546 (N_7546,N_5789,N_5470);
nand U7547 (N_7547,N_6614,N_6937);
and U7548 (N_7548,N_7349,N_5105);
xor U7549 (N_7549,N_6213,N_6063);
nor U7550 (N_7550,N_7336,N_6333);
nor U7551 (N_7551,N_7485,N_5124);
nand U7552 (N_7552,N_7110,N_6047);
xor U7553 (N_7553,N_5796,N_6201);
xor U7554 (N_7554,N_6742,N_7164);
nand U7555 (N_7555,N_6429,N_6838);
or U7556 (N_7556,N_5964,N_5913);
and U7557 (N_7557,N_7449,N_5748);
xor U7558 (N_7558,N_5482,N_6035);
xor U7559 (N_7559,N_5917,N_6174);
and U7560 (N_7560,N_6509,N_5133);
and U7561 (N_7561,N_7230,N_6503);
xnor U7562 (N_7562,N_5922,N_5416);
xor U7563 (N_7563,N_6978,N_5452);
and U7564 (N_7564,N_6343,N_5070);
and U7565 (N_7565,N_5598,N_6575);
and U7566 (N_7566,N_5636,N_5665);
xor U7567 (N_7567,N_6621,N_7212);
xor U7568 (N_7568,N_5155,N_5994);
xor U7569 (N_7569,N_5719,N_7144);
or U7570 (N_7570,N_5972,N_6081);
and U7571 (N_7571,N_7352,N_6569);
xor U7572 (N_7572,N_6724,N_7060);
nor U7573 (N_7573,N_6252,N_5556);
or U7574 (N_7574,N_5528,N_6610);
nor U7575 (N_7575,N_5952,N_7393);
nand U7576 (N_7576,N_6307,N_6385);
xnor U7577 (N_7577,N_7488,N_6133);
or U7578 (N_7578,N_5029,N_6319);
nand U7579 (N_7579,N_5802,N_5708);
and U7580 (N_7580,N_6511,N_5426);
or U7581 (N_7581,N_5682,N_6406);
xor U7582 (N_7582,N_6564,N_5697);
xnor U7583 (N_7583,N_5091,N_6866);
and U7584 (N_7584,N_6197,N_6061);
nand U7585 (N_7585,N_6298,N_5674);
xor U7586 (N_7586,N_6074,N_6295);
or U7587 (N_7587,N_6984,N_6601);
nor U7588 (N_7588,N_6109,N_7106);
nor U7589 (N_7589,N_6495,N_5103);
or U7590 (N_7590,N_7423,N_6807);
nor U7591 (N_7591,N_5028,N_7027);
nand U7592 (N_7592,N_6561,N_6085);
and U7593 (N_7593,N_6888,N_6527);
xor U7594 (N_7594,N_6007,N_6744);
nand U7595 (N_7595,N_6203,N_6755);
nor U7596 (N_7596,N_7026,N_6587);
and U7597 (N_7597,N_6747,N_7112);
xor U7598 (N_7598,N_5466,N_5132);
nor U7599 (N_7599,N_5729,N_5626);
and U7600 (N_7600,N_7335,N_6011);
and U7601 (N_7601,N_7464,N_6686);
nor U7602 (N_7602,N_5373,N_6049);
nor U7603 (N_7603,N_7435,N_6336);
and U7604 (N_7604,N_5366,N_5861);
and U7605 (N_7605,N_5250,N_5309);
nor U7606 (N_7606,N_6894,N_6598);
and U7607 (N_7607,N_6041,N_7479);
and U7608 (N_7608,N_7351,N_7217);
nand U7609 (N_7609,N_6566,N_7353);
nor U7610 (N_7610,N_5546,N_7195);
nand U7611 (N_7611,N_6787,N_5246);
xor U7612 (N_7612,N_7205,N_6532);
and U7613 (N_7613,N_5396,N_6153);
or U7614 (N_7614,N_7199,N_6715);
and U7615 (N_7615,N_7220,N_5413);
nand U7616 (N_7616,N_5525,N_6478);
or U7617 (N_7617,N_5581,N_7460);
xor U7618 (N_7618,N_5143,N_6998);
and U7619 (N_7619,N_6642,N_5549);
or U7620 (N_7620,N_5524,N_6913);
xnor U7621 (N_7621,N_5532,N_6798);
or U7622 (N_7622,N_5571,N_7063);
and U7623 (N_7623,N_6139,N_5271);
xnor U7624 (N_7624,N_7113,N_7095);
and U7625 (N_7625,N_6393,N_6974);
nand U7626 (N_7626,N_5696,N_5785);
and U7627 (N_7627,N_5210,N_6518);
nor U7628 (N_7628,N_5382,N_6526);
and U7629 (N_7629,N_5656,N_6775);
nor U7630 (N_7630,N_6481,N_5062);
or U7631 (N_7631,N_6095,N_5737);
nand U7632 (N_7632,N_7234,N_5949);
nor U7633 (N_7633,N_6710,N_5148);
or U7634 (N_7634,N_7186,N_6398);
nand U7635 (N_7635,N_5631,N_6964);
nor U7636 (N_7636,N_5173,N_6331);
xor U7637 (N_7637,N_5400,N_5475);
and U7638 (N_7638,N_7021,N_7076);
nand U7639 (N_7639,N_7214,N_5042);
nor U7640 (N_7640,N_7366,N_6817);
nor U7641 (N_7641,N_6186,N_6157);
nand U7642 (N_7642,N_6165,N_7498);
nand U7643 (N_7643,N_5705,N_5527);
or U7644 (N_7644,N_5189,N_6870);
and U7645 (N_7645,N_6966,N_6571);
or U7646 (N_7646,N_6025,N_6730);
xnor U7647 (N_7647,N_6391,N_6367);
xor U7648 (N_7648,N_7469,N_6054);
and U7649 (N_7649,N_6951,N_6884);
and U7650 (N_7650,N_6005,N_5619);
xor U7651 (N_7651,N_5552,N_6176);
xnor U7652 (N_7652,N_5433,N_6542);
xor U7653 (N_7653,N_6226,N_6924);
or U7654 (N_7654,N_5436,N_6961);
xor U7655 (N_7655,N_6612,N_5965);
or U7656 (N_7656,N_5793,N_6364);
or U7657 (N_7657,N_6857,N_6265);
nor U7658 (N_7658,N_7370,N_6382);
nand U7659 (N_7659,N_6117,N_6264);
and U7660 (N_7660,N_5825,N_5120);
and U7661 (N_7661,N_6680,N_7048);
and U7662 (N_7662,N_5718,N_6324);
and U7663 (N_7663,N_6847,N_6193);
and U7664 (N_7664,N_7084,N_5021);
xor U7665 (N_7665,N_5545,N_5074);
and U7666 (N_7666,N_7382,N_5774);
or U7667 (N_7667,N_6591,N_5372);
or U7668 (N_7668,N_5242,N_6792);
nor U7669 (N_7669,N_7250,N_6434);
nand U7670 (N_7670,N_5461,N_6340);
nand U7671 (N_7671,N_6107,N_6917);
or U7672 (N_7672,N_7041,N_5112);
and U7673 (N_7673,N_5049,N_6028);
or U7674 (N_7674,N_7284,N_6065);
or U7675 (N_7675,N_7075,N_5230);
and U7676 (N_7676,N_5685,N_5940);
and U7677 (N_7677,N_5023,N_6266);
nor U7678 (N_7678,N_6623,N_5874);
xor U7679 (N_7679,N_5121,N_5043);
and U7680 (N_7680,N_6505,N_5228);
or U7681 (N_7681,N_7455,N_6781);
nor U7682 (N_7682,N_6523,N_6289);
nand U7683 (N_7683,N_6618,N_5934);
xor U7684 (N_7684,N_6513,N_7170);
nand U7685 (N_7685,N_6704,N_6414);
or U7686 (N_7686,N_6982,N_7394);
or U7687 (N_7687,N_7367,N_5069);
or U7688 (N_7688,N_6160,N_6667);
or U7689 (N_7689,N_6725,N_6108);
and U7690 (N_7690,N_5773,N_6239);
nor U7691 (N_7691,N_5232,N_6103);
xor U7692 (N_7692,N_7405,N_5788);
or U7693 (N_7693,N_5414,N_6013);
and U7694 (N_7694,N_6749,N_7252);
and U7695 (N_7695,N_7229,N_7444);
nand U7696 (N_7696,N_5841,N_6956);
xnor U7697 (N_7697,N_6624,N_6348);
or U7698 (N_7698,N_6057,N_7239);
or U7699 (N_7699,N_7391,N_6296);
or U7700 (N_7700,N_7289,N_5652);
nor U7701 (N_7701,N_7481,N_7174);
xnor U7702 (N_7702,N_6351,N_7342);
xor U7703 (N_7703,N_6825,N_5501);
nand U7704 (N_7704,N_6077,N_6435);
or U7705 (N_7705,N_6458,N_6622);
nand U7706 (N_7706,N_7099,N_7203);
xor U7707 (N_7707,N_5111,N_5185);
nor U7708 (N_7708,N_6630,N_6457);
nor U7709 (N_7709,N_6791,N_5826);
or U7710 (N_7710,N_7218,N_7417);
xnor U7711 (N_7711,N_7023,N_7355);
nor U7712 (N_7712,N_6327,N_5138);
or U7713 (N_7713,N_6795,N_6431);
or U7714 (N_7714,N_7088,N_6844);
xnor U7715 (N_7715,N_6415,N_6996);
or U7716 (N_7716,N_5688,N_6455);
nand U7717 (N_7717,N_5147,N_6119);
nor U7718 (N_7718,N_5569,N_7159);
xnor U7719 (N_7719,N_5852,N_7465);
or U7720 (N_7720,N_6145,N_5499);
nand U7721 (N_7721,N_5421,N_6088);
and U7722 (N_7722,N_5253,N_5090);
and U7723 (N_7723,N_5354,N_5566);
xor U7724 (N_7724,N_6948,N_5572);
nand U7725 (N_7725,N_5387,N_5710);
xnor U7726 (N_7726,N_6300,N_5776);
and U7727 (N_7727,N_6727,N_5711);
nand U7728 (N_7728,N_5163,N_7471);
nand U7729 (N_7729,N_6818,N_7116);
nor U7730 (N_7730,N_5097,N_7183);
or U7731 (N_7731,N_7412,N_5100);
or U7732 (N_7732,N_5498,N_5221);
nand U7733 (N_7733,N_6173,N_5586);
or U7734 (N_7734,N_6500,N_5215);
nand U7735 (N_7735,N_6131,N_5618);
nor U7736 (N_7736,N_7255,N_6446);
xnor U7737 (N_7737,N_7142,N_7044);
nand U7738 (N_7738,N_5842,N_7344);
nor U7739 (N_7739,N_6126,N_5259);
or U7740 (N_7740,N_6605,N_5967);
nand U7741 (N_7741,N_7376,N_6029);
xor U7742 (N_7742,N_5139,N_7420);
xnor U7743 (N_7743,N_5375,N_6552);
or U7744 (N_7744,N_6373,N_6177);
nand U7745 (N_7745,N_7003,N_6839);
xnor U7746 (N_7746,N_6106,N_5991);
nand U7747 (N_7747,N_7443,N_6769);
xnor U7748 (N_7748,N_5559,N_7249);
nand U7749 (N_7749,N_5521,N_5389);
nor U7750 (N_7750,N_6380,N_6835);
xor U7751 (N_7751,N_7499,N_6897);
xnor U7752 (N_7752,N_5386,N_6655);
nor U7753 (N_7753,N_7236,N_7381);
or U7754 (N_7754,N_6672,N_5233);
nor U7755 (N_7755,N_6314,N_6930);
or U7756 (N_7756,N_6635,N_6480);
nand U7757 (N_7757,N_6823,N_6467);
nand U7758 (N_7758,N_5122,N_7104);
xnor U7759 (N_7759,N_5486,N_5577);
xnor U7760 (N_7760,N_5272,N_5906);
and U7761 (N_7761,N_5827,N_6258);
xor U7762 (N_7762,N_6196,N_6171);
xor U7763 (N_7763,N_5180,N_7038);
nor U7764 (N_7764,N_5418,N_5076);
or U7765 (N_7765,N_6963,N_5495);
nand U7766 (N_7766,N_6159,N_6973);
or U7767 (N_7767,N_7163,N_7102);
or U7768 (N_7768,N_7422,N_5786);
nand U7769 (N_7769,N_6581,N_6277);
xnor U7770 (N_7770,N_6368,N_6304);
nor U7771 (N_7771,N_5654,N_5096);
xor U7772 (N_7772,N_5782,N_7225);
nand U7773 (N_7773,N_6826,N_6432);
xor U7774 (N_7774,N_5195,N_5284);
nand U7775 (N_7775,N_7155,N_7495);
and U7776 (N_7776,N_6908,N_6565);
and U7777 (N_7777,N_5219,N_6046);
nor U7778 (N_7778,N_5238,N_5815);
nand U7779 (N_7779,N_6899,N_7074);
nor U7780 (N_7780,N_5166,N_5283);
xor U7781 (N_7781,N_7338,N_6926);
nor U7782 (N_7782,N_5628,N_7117);
xnor U7783 (N_7783,N_7070,N_6115);
xor U7784 (N_7784,N_7094,N_7322);
and U7785 (N_7785,N_5035,N_6529);
nor U7786 (N_7786,N_6957,N_5114);
or U7787 (N_7787,N_6827,N_5522);
nand U7788 (N_7788,N_7019,N_5497);
or U7789 (N_7789,N_5607,N_5578);
nand U7790 (N_7790,N_6539,N_6925);
xor U7791 (N_7791,N_7055,N_5632);
or U7792 (N_7792,N_6733,N_6110);
xnor U7793 (N_7793,N_6362,N_6611);
or U7794 (N_7794,N_6221,N_5342);
and U7795 (N_7795,N_5363,N_6101);
nor U7796 (N_7796,N_7365,N_5585);
xor U7797 (N_7797,N_5536,N_5627);
or U7798 (N_7798,N_7384,N_6949);
xnor U7799 (N_7799,N_6472,N_6421);
and U7800 (N_7800,N_6248,N_5164);
nor U7801 (N_7801,N_6236,N_6355);
nand U7802 (N_7802,N_5307,N_6767);
nor U7803 (N_7803,N_5932,N_6369);
xor U7804 (N_7804,N_5968,N_7299);
nand U7805 (N_7805,N_6192,N_5199);
xor U7806 (N_7806,N_5084,N_6921);
or U7807 (N_7807,N_5423,N_5642);
nand U7808 (N_7808,N_6052,N_6498);
nor U7809 (N_7809,N_5863,N_7242);
and U7810 (N_7810,N_5813,N_5832);
and U7811 (N_7811,N_5287,N_6315);
nor U7812 (N_7812,N_6317,N_6875);
nor U7813 (N_7813,N_5385,N_5780);
nand U7814 (N_7814,N_7325,N_7161);
nand U7815 (N_7815,N_6896,N_6515);
xnor U7816 (N_7816,N_6709,N_6763);
nand U7817 (N_7817,N_7187,N_5371);
xnor U7818 (N_7818,N_5969,N_5986);
nand U7819 (N_7819,N_5762,N_7309);
or U7820 (N_7820,N_5993,N_6075);
nor U7821 (N_7821,N_6928,N_6089);
nor U7822 (N_7822,N_5765,N_6900);
nand U7823 (N_7823,N_7270,N_5515);
nand U7824 (N_7824,N_6227,N_7363);
xnor U7825 (N_7825,N_6806,N_5447);
nand U7826 (N_7826,N_6206,N_7022);
xnor U7827 (N_7827,N_7181,N_6312);
and U7828 (N_7828,N_5229,N_5595);
nand U7829 (N_7829,N_6599,N_5772);
and U7830 (N_7830,N_6705,N_6883);
xor U7831 (N_7831,N_5045,N_7379);
and U7832 (N_7832,N_6316,N_6768);
nor U7833 (N_7833,N_6701,N_5957);
and U7834 (N_7834,N_5643,N_5109);
xor U7835 (N_7835,N_6087,N_7167);
or U7836 (N_7836,N_5516,N_7191);
or U7837 (N_7837,N_7192,N_5388);
and U7838 (N_7838,N_5756,N_5188);
xnor U7839 (N_7839,N_5280,N_5040);
and U7840 (N_7840,N_6502,N_5145);
or U7841 (N_7841,N_5016,N_6869);
nor U7842 (N_7842,N_6673,N_6766);
nand U7843 (N_7843,N_6449,N_6790);
nand U7844 (N_7844,N_6661,N_5854);
nor U7845 (N_7845,N_5144,N_6760);
and U7846 (N_7846,N_6753,N_5432);
and U7847 (N_7847,N_7108,N_5974);
and U7848 (N_7848,N_6151,N_5411);
xor U7849 (N_7849,N_6335,N_7206);
and U7850 (N_7850,N_6627,N_7194);
nand U7851 (N_7851,N_5992,N_5247);
or U7852 (N_7852,N_7009,N_5623);
xnor U7853 (N_7853,N_6220,N_6568);
or U7854 (N_7854,N_5858,N_7141);
xor U7855 (N_7855,N_5835,N_6384);
or U7856 (N_7856,N_5582,N_5911);
nand U7857 (N_7857,N_5520,N_5768);
and U7858 (N_7858,N_7276,N_6032);
nor U7859 (N_7859,N_5583,N_7082);
xnor U7860 (N_7860,N_6815,N_6405);
nand U7861 (N_7861,N_5523,N_5009);
and U7862 (N_7862,N_6700,N_6895);
or U7863 (N_7863,N_7120,N_6423);
or U7864 (N_7864,N_7428,N_5184);
nor U7865 (N_7865,N_5669,N_5667);
or U7866 (N_7866,N_5065,N_6030);
nand U7867 (N_7867,N_5358,N_6987);
nand U7868 (N_7868,N_5961,N_6156);
nor U7869 (N_7869,N_5362,N_5990);
nor U7870 (N_7870,N_7091,N_7446);
or U7871 (N_7871,N_6267,N_7035);
nor U7872 (N_7872,N_5302,N_6158);
and U7873 (N_7873,N_5018,N_5717);
xor U7874 (N_7874,N_5314,N_7050);
and U7875 (N_7875,N_6656,N_5738);
nand U7876 (N_7876,N_6347,N_7399);
nand U7877 (N_7877,N_7244,N_5727);
nand U7878 (N_7878,N_5026,N_5837);
xor U7879 (N_7879,N_5931,N_5985);
xnor U7880 (N_7880,N_5442,N_6703);
nand U7881 (N_7881,N_7372,N_6958);
xnor U7882 (N_7882,N_6714,N_6770);
and U7883 (N_7883,N_5380,N_6489);
nand U7884 (N_7884,N_7392,N_7178);
xor U7885 (N_7885,N_6191,N_6015);
xnor U7886 (N_7886,N_7101,N_7388);
or U7887 (N_7887,N_5759,N_6450);
xnor U7888 (N_7888,N_6745,N_5912);
and U7889 (N_7889,N_6463,N_7288);
or U7890 (N_7890,N_7373,N_7346);
or U7891 (N_7891,N_5269,N_5439);
nand U7892 (N_7892,N_5194,N_5672);
xor U7893 (N_7893,N_5293,N_6994);
nand U7894 (N_7894,N_5172,N_6473);
xnor U7895 (N_7895,N_7315,N_6789);
nor U7896 (N_7896,N_6922,N_7345);
xor U7897 (N_7897,N_5419,N_5316);
xnor U7898 (N_7898,N_6273,N_6161);
and U7899 (N_7899,N_5805,N_5808);
or U7900 (N_7900,N_5935,N_7359);
xnor U7901 (N_7901,N_5322,N_6181);
nor U7902 (N_7902,N_7282,N_6969);
nand U7903 (N_7903,N_5429,N_6889);
xnor U7904 (N_7904,N_7177,N_6140);
xor U7905 (N_7905,N_5165,N_6127);
or U7906 (N_7906,N_7165,N_5666);
and U7907 (N_7907,N_5468,N_7450);
nand U7908 (N_7908,N_5547,N_5925);
or U7909 (N_7909,N_5104,N_7073);
xor U7910 (N_7910,N_6187,N_6175);
nor U7911 (N_7911,N_6501,N_6545);
or U7912 (N_7912,N_5510,N_5875);
or U7913 (N_7913,N_5170,N_5915);
and U7914 (N_7914,N_6858,N_5224);
nand U7915 (N_7915,N_5297,N_5146);
and U7916 (N_7916,N_6274,N_6892);
and U7917 (N_7917,N_6476,N_6471);
or U7918 (N_7918,N_7100,N_5136);
xor U7919 (N_7919,N_7259,N_6548);
xnor U7920 (N_7920,N_6649,N_6554);
and U7921 (N_7921,N_6965,N_5449);
nor U7922 (N_7922,N_5205,N_5127);
nor U7923 (N_7923,N_6379,N_7097);
xnor U7924 (N_7924,N_7251,N_7153);
or U7925 (N_7925,N_5966,N_6720);
and U7926 (N_7926,N_6019,N_6976);
nand U7927 (N_7927,N_6856,N_7330);
or U7928 (N_7928,N_7425,N_6230);
or U7929 (N_7929,N_7257,N_5014);
nor U7930 (N_7930,N_6448,N_6750);
and U7931 (N_7931,N_5067,N_7154);
or U7932 (N_7932,N_7016,N_5295);
and U7933 (N_7933,N_6233,N_6199);
and U7934 (N_7934,N_6474,N_5838);
nor U7935 (N_7935,N_7300,N_7087);
and U7936 (N_7936,N_5819,N_5655);
or U7937 (N_7937,N_7297,N_6756);
xor U7938 (N_7938,N_6843,N_5941);
nor U7939 (N_7939,N_5880,N_5490);
nor U7940 (N_7940,N_6282,N_7029);
and U7941 (N_7941,N_6339,N_7147);
xnor U7942 (N_7942,N_7246,N_6096);
xnor U7943 (N_7943,N_7248,N_6130);
nand U7944 (N_7944,N_7219,N_7197);
nor U7945 (N_7945,N_5364,N_5458);
xor U7946 (N_7946,N_6392,N_5444);
nand U7947 (N_7947,N_5999,N_6645);
nand U7948 (N_7948,N_6195,N_6670);
nor U7949 (N_7949,N_7010,N_6313);
nor U7950 (N_7950,N_5448,N_5594);
xnor U7951 (N_7951,N_6209,N_5503);
nand U7952 (N_7952,N_6692,N_6276);
nor U7953 (N_7953,N_7409,N_7015);
nand U7954 (N_7954,N_6440,N_6129);
nor U7955 (N_7955,N_5300,N_6521);
or U7956 (N_7956,N_5051,N_6208);
xor U7957 (N_7957,N_6902,N_7004);
xnor U7958 (N_7958,N_6939,N_6819);
nand U7959 (N_7959,N_7380,N_5956);
or U7960 (N_7960,N_5775,N_6759);
nand U7961 (N_7961,N_5267,N_6207);
xnor U7962 (N_7962,N_6915,N_5505);
nand U7963 (N_7963,N_6395,N_7032);
or U7964 (N_7964,N_7494,N_5828);
or U7965 (N_7965,N_6528,N_7081);
xor U7966 (N_7966,N_5193,N_6945);
or U7967 (N_7967,N_6142,N_5914);
nor U7968 (N_7968,N_6960,N_7343);
or U7969 (N_7969,N_6376,N_5794);
nand U7970 (N_7970,N_7017,N_7204);
and U7971 (N_7971,N_6488,N_5865);
xor U7972 (N_7972,N_5101,N_7286);
xor U7973 (N_7973,N_6562,N_5081);
or U7974 (N_7974,N_7115,N_6696);
xnor U7975 (N_7975,N_6255,N_6663);
xnor U7976 (N_7976,N_6991,N_6292);
nor U7977 (N_7977,N_6997,N_6425);
and U7978 (N_7978,N_5422,N_7296);
xnor U7979 (N_7979,N_6045,N_5512);
and U7980 (N_7980,N_6490,N_7316);
xor U7981 (N_7981,N_5116,N_5410);
xnor U7982 (N_7982,N_6270,N_7374);
nand U7983 (N_7983,N_5981,N_6836);
or U7984 (N_7984,N_5428,N_6416);
xor U7985 (N_7985,N_5003,N_5897);
or U7986 (N_7986,N_5893,N_6263);
nor U7987 (N_7987,N_7414,N_7331);
or U7988 (N_7988,N_5537,N_5102);
and U7989 (N_7989,N_5099,N_5971);
xor U7990 (N_7990,N_5020,N_5760);
nor U7991 (N_7991,N_5437,N_5401);
and U7992 (N_7992,N_6014,N_5381);
nand U7993 (N_7993,N_7262,N_5438);
nand U7994 (N_7994,N_6390,N_7285);
nor U7995 (N_7995,N_6690,N_6346);
and U7996 (N_7996,N_6018,N_7467);
and U7997 (N_7997,N_5824,N_7375);
nand U7998 (N_7998,N_5816,N_6402);
and U7999 (N_7999,N_5703,N_6762);
nand U8000 (N_8000,N_6086,N_7000);
nand U8001 (N_8001,N_5351,N_6178);
nand U8002 (N_8002,N_5644,N_6249);
and U8003 (N_8003,N_6050,N_5701);
xor U8004 (N_8004,N_5988,N_6732);
nor U8005 (N_8005,N_6520,N_6579);
and U8006 (N_8006,N_5326,N_5368);
xnor U8007 (N_8007,N_6810,N_5408);
or U8008 (N_8008,N_5534,N_6613);
or U8009 (N_8009,N_6071,N_5541);
and U8010 (N_8010,N_5034,N_7065);
xor U8011 (N_8011,N_5680,N_7416);
nand U8012 (N_8012,N_6034,N_5083);
and U8013 (N_8013,N_5763,N_6786);
and U8014 (N_8014,N_7169,N_5311);
nor U8015 (N_8015,N_6619,N_5171);
nor U8016 (N_8016,N_5347,N_6219);
and U8017 (N_8017,N_5191,N_5611);
or U8018 (N_8018,N_5621,N_5847);
and U8019 (N_8019,N_5662,N_5871);
xnor U8020 (N_8020,N_6040,N_5648);
and U8021 (N_8021,N_5698,N_5473);
xnor U8022 (N_8022,N_5263,N_7253);
and U8023 (N_8023,N_7275,N_7475);
xor U8024 (N_8024,N_6294,N_6179);
or U8025 (N_8025,N_6560,N_6682);
xnor U8026 (N_8026,N_5390,N_5454);
or U8027 (N_8027,N_7256,N_6944);
nand U8028 (N_8028,N_5947,N_5151);
xnor U8029 (N_8029,N_5857,N_5620);
nor U8030 (N_8030,N_7011,N_6694);
and U8031 (N_8031,N_5676,N_5591);
xnor U8032 (N_8032,N_5856,N_5910);
nand U8033 (N_8033,N_5299,N_7341);
or U8034 (N_8034,N_5739,N_6167);
and U8035 (N_8035,N_7271,N_6918);
or U8036 (N_8036,N_5519,N_5787);
and U8037 (N_8037,N_7001,N_5206);
and U8038 (N_8038,N_5465,N_7089);
or U8039 (N_8039,N_6111,N_6738);
or U8040 (N_8040,N_6090,N_7085);
nand U8041 (N_8041,N_6439,N_6719);
and U8042 (N_8042,N_7266,N_5208);
or U8043 (N_8043,N_6155,N_6217);
or U8044 (N_8044,N_7188,N_5251);
nor U8045 (N_8045,N_6009,N_5068);
nor U8046 (N_8046,N_5518,N_6322);
xor U8047 (N_8047,N_6754,N_7293);
nand U8048 (N_8048,N_6865,N_7317);
nand U8049 (N_8049,N_6468,N_5891);
or U8050 (N_8050,N_6607,N_5462);
nor U8051 (N_8051,N_6947,N_6357);
xor U8052 (N_8052,N_5288,N_6868);
xnor U8053 (N_8053,N_7339,N_7006);
nor U8054 (N_8054,N_5530,N_5235);
nand U8055 (N_8055,N_5995,N_5955);
and U8056 (N_8056,N_5349,N_7190);
or U8057 (N_8057,N_7442,N_7012);
xnor U8058 (N_8058,N_6855,N_6283);
nor U8059 (N_8059,N_5187,N_6125);
nor U8060 (N_8060,N_6625,N_6609);
nor U8061 (N_8061,N_6290,N_7007);
and U8062 (N_8062,N_5855,N_5025);
nand U8063 (N_8063,N_5728,N_7437);
nor U8064 (N_8064,N_6136,N_5430);
nor U8065 (N_8065,N_5744,N_7486);
or U8066 (N_8066,N_5334,N_7440);
and U8067 (N_8067,N_5777,N_5273);
xor U8068 (N_8068,N_5367,N_6002);
nor U8069 (N_8069,N_6793,N_6483);
nor U8070 (N_8070,N_6660,N_5359);
nand U8071 (N_8071,N_5344,N_7175);
nand U8072 (N_8072,N_7403,N_6721);
xor U8073 (N_8073,N_6235,N_6805);
or U8074 (N_8074,N_6780,N_5916);
nand U8075 (N_8075,N_5614,N_6647);
and U8076 (N_8076,N_5846,N_7456);
xnor U8077 (N_8077,N_6427,N_5060);
nand U8078 (N_8078,N_6496,N_6809);
xor U8079 (N_8079,N_7424,N_7137);
nor U8080 (N_8080,N_6058,N_6563);
nor U8081 (N_8081,N_6774,N_5707);
and U8082 (N_8082,N_6189,N_6350);
or U8083 (N_8083,N_7477,N_6540);
or U8084 (N_8084,N_7386,N_7148);
xor U8085 (N_8085,N_7311,N_5726);
or U8086 (N_8086,N_5810,N_7432);
and U8087 (N_8087,N_7415,N_7321);
nor U8088 (N_8088,N_6594,N_7245);
xnor U8089 (N_8089,N_6764,N_5252);
and U8090 (N_8090,N_5926,N_5226);
and U8091 (N_8091,N_5115,N_5989);
nor U8092 (N_8092,N_7451,N_7398);
or U8093 (N_8093,N_6757,N_5130);
nor U8094 (N_8094,N_5168,N_5562);
nor U8095 (N_8095,N_6699,N_7111);
and U8096 (N_8096,N_5544,N_7166);
nor U8097 (N_8097,N_6980,N_5218);
or U8098 (N_8098,N_5755,N_7083);
nand U8099 (N_8099,N_7086,N_6708);
nor U8100 (N_8100,N_5456,N_5217);
xnor U8101 (N_8101,N_7056,N_7396);
xnor U8102 (N_8102,N_6977,N_7463);
or U8103 (N_8103,N_6242,N_6979);
and U8104 (N_8104,N_7483,N_5107);
or U8105 (N_8105,N_5404,N_7461);
or U8106 (N_8106,N_5879,N_6586);
and U8107 (N_8107,N_7130,N_7361);
and U8108 (N_8108,N_6573,N_5730);
nor U8109 (N_8109,N_6275,N_5474);
xnor U8110 (N_8110,N_7310,N_5278);
or U8111 (N_8111,N_5092,N_5118);
or U8112 (N_8112,N_5002,N_7291);
and U8113 (N_8113,N_6940,N_5783);
or U8114 (N_8114,N_5973,N_5409);
nand U8115 (N_8115,N_5198,N_6010);
nand U8116 (N_8116,N_5024,N_7358);
or U8117 (N_8117,N_7371,N_6650);
xnor U8118 (N_8118,N_7068,N_7281);
nand U8119 (N_8119,N_5601,N_5223);
nand U8120 (N_8120,N_5001,N_7064);
xor U8121 (N_8121,N_5453,N_6589);
xnor U8122 (N_8122,N_6631,N_6422);
nor U8123 (N_8123,N_5262,N_6254);
or U8124 (N_8124,N_7221,N_6454);
or U8125 (N_8125,N_6269,N_5679);
nor U8126 (N_8126,N_5181,N_6079);
and U8127 (N_8127,N_6675,N_6531);
nand U8128 (N_8128,N_5766,N_5745);
nand U8129 (N_8129,N_6880,N_7079);
xnor U8130 (N_8130,N_5565,N_5997);
nand U8131 (N_8131,N_6517,N_5053);
nor U8132 (N_8132,N_6687,N_6626);
nand U8133 (N_8133,N_5681,N_6617);
and U8134 (N_8134,N_6683,N_5907);
or U8135 (N_8135,N_5807,N_5767);
nor U8136 (N_8136,N_6995,N_5869);
or U8137 (N_8137,N_5160,N_7334);
nand U8138 (N_8138,N_6008,N_6389);
nor U8139 (N_8139,N_6026,N_7493);
or U8140 (N_8140,N_5908,N_5743);
and U8141 (N_8141,N_6688,N_5950);
nor U8142 (N_8142,N_5277,N_7328);
nand U8143 (N_8143,N_6148,N_5939);
and U8144 (N_8144,N_7324,N_5153);
nor U8145 (N_8145,N_5976,N_6433);
nor U8146 (N_8146,N_7168,N_6638);
nor U8147 (N_8147,N_7237,N_6212);
nand U8148 (N_8148,N_6971,N_5784);
xor U8149 (N_8149,N_5650,N_7228);
xor U8150 (N_8150,N_7196,N_5919);
nor U8151 (N_8151,N_6365,N_6325);
or U8152 (N_8152,N_5174,N_7024);
nand U8153 (N_8153,N_6867,N_7295);
xor U8154 (N_8154,N_5303,N_7034);
or U8155 (N_8155,N_7261,N_6027);
or U8156 (N_8156,N_6437,N_6530);
xor U8157 (N_8157,N_5403,N_5379);
nand U8158 (N_8158,N_5629,N_6408);
or U8159 (N_8159,N_7265,N_6814);
and U8160 (N_8160,N_7233,N_7162);
nand U8161 (N_8161,N_6036,N_7119);
nor U8162 (N_8162,N_5369,N_6557);
and U8163 (N_8163,N_5849,N_5829);
nor U8164 (N_8164,N_6885,N_5616);
and U8165 (N_8165,N_6268,N_6043);
xnor U8166 (N_8166,N_6381,N_6419);
or U8167 (N_8167,N_6184,N_6832);
or U8168 (N_8168,N_6400,N_5812);
and U8169 (N_8169,N_7020,N_6905);
xor U8170 (N_8170,N_5348,N_5661);
nor U8171 (N_8171,N_5690,N_5019);
and U8172 (N_8172,N_6098,N_6305);
or U8173 (N_8173,N_5860,N_5047);
or U8174 (N_8174,N_6570,N_6407);
and U8175 (N_8175,N_6691,N_5050);
nand U8176 (N_8176,N_6772,N_6244);
or U8177 (N_8177,N_6652,N_6337);
xor U8178 (N_8178,N_6812,N_5467);
nand U8179 (N_8179,N_5352,N_6989);
or U8180 (N_8180,N_7263,N_6804);
nand U8181 (N_8181,N_7438,N_6603);
nor U8182 (N_8182,N_5647,N_6241);
and U8183 (N_8183,N_6225,N_5258);
xnor U8184 (N_8184,N_5814,N_6919);
nor U8185 (N_8185,N_7268,N_6550);
xor U8186 (N_8186,N_5699,N_6848);
nor U8187 (N_8187,N_5615,N_6674);
nor U8188 (N_8188,N_5085,N_6060);
and U8189 (N_8189,N_5695,N_5041);
or U8190 (N_8190,N_6716,N_5204);
xnor U8191 (N_8191,N_6999,N_6637);
nand U8192 (N_8192,N_5129,N_5378);
or U8193 (N_8193,N_5700,N_6728);
or U8194 (N_8194,N_5417,N_5017);
nand U8195 (N_8195,N_7054,N_7103);
nor U8196 (N_8196,N_6135,N_6188);
nand U8197 (N_8197,N_5469,N_6121);
or U8198 (N_8198,N_6286,N_5030);
xor U8199 (N_8199,N_6466,N_5579);
or U8200 (N_8200,N_5341,N_5182);
or U8201 (N_8201,N_5580,N_5340);
and U8202 (N_8202,N_5434,N_6628);
nand U8203 (N_8203,N_7061,N_5157);
nor U8204 (N_8204,N_5901,N_5249);
nor U8205 (N_8205,N_6361,N_6831);
nor U8206 (N_8206,N_6116,N_6146);
or U8207 (N_8207,N_6198,N_6851);
or U8208 (N_8208,N_5240,N_5472);
or U8209 (N_8209,N_5000,N_7152);
xor U8210 (N_8210,N_5716,N_7347);
and U8211 (N_8211,N_7418,N_7274);
nor U8212 (N_8212,N_5836,N_6931);
and U8213 (N_8213,N_6309,N_6771);
xnor U8214 (N_8214,N_6214,N_5658);
or U8215 (N_8215,N_7005,N_5178);
or U8216 (N_8216,N_6215,N_5007);
nand U8217 (N_8217,N_6070,N_5298);
nor U8218 (N_8218,N_6935,N_7198);
nor U8219 (N_8219,N_6354,N_5892);
nor U8220 (N_8220,N_6936,N_5878);
nor U8221 (N_8221,N_6706,N_5318);
and U8222 (N_8222,N_7458,N_5345);
nor U8223 (N_8223,N_7290,N_6853);
nand U8224 (N_8224,N_5909,N_6491);
nand U8225 (N_8225,N_5225,N_5924);
and U8226 (N_8226,N_7053,N_6684);
nand U8227 (N_8227,N_5850,N_7470);
nand U8228 (N_8228,N_5061,N_7320);
nand U8229 (N_8229,N_6954,N_6746);
or U8230 (N_8230,N_5004,N_5890);
and U8231 (N_8231,N_7185,N_6366);
and U8232 (N_8232,N_6693,N_5653);
xor U8233 (N_8233,N_7389,N_5504);
and U8234 (N_8234,N_7150,N_7071);
nand U8235 (N_8235,N_6210,N_6462);
and U8236 (N_8236,N_5290,N_6397);
and U8237 (N_8237,N_5011,N_6820);
and U8238 (N_8238,N_7340,N_5741);
or U8239 (N_8239,N_5058,N_5477);
nor U8240 (N_8240,N_5560,N_6172);
xor U8241 (N_8241,N_6363,N_6634);
or U8242 (N_8242,N_5677,N_6396);
xor U8243 (N_8243,N_6122,N_5125);
nand U8244 (N_8244,N_7385,N_6291);
or U8245 (N_8245,N_5075,N_5693);
nor U8246 (N_8246,N_6640,N_5613);
xor U8247 (N_8247,N_6953,N_7160);
nor U8248 (N_8248,N_6410,N_6606);
and U8249 (N_8249,N_5984,N_5570);
nand U8250 (N_8250,N_7377,N_7013);
xnor U8251 (N_8251,N_6261,N_6512);
nor U8252 (N_8252,N_7173,N_6580);
xor U8253 (N_8253,N_6303,N_7058);
xor U8254 (N_8254,N_5640,N_6487);
xnor U8255 (N_8255,N_7077,N_6118);
and U8256 (N_8256,N_5324,N_6084);
xor U8257 (N_8257,N_5450,N_5757);
nor U8258 (N_8258,N_6524,N_5149);
nor U8259 (N_8259,N_6204,N_7243);
and U8260 (N_8260,N_6062,N_6318);
nand U8261 (N_8261,N_5073,N_5315);
nor U8262 (N_8262,N_6927,N_6232);
or U8263 (N_8263,N_5207,N_6778);
nand U8264 (N_8264,N_5089,N_6829);
nor U8265 (N_8265,N_5894,N_5660);
nor U8266 (N_8266,N_6059,N_5946);
nand U8267 (N_8267,N_5978,N_6053);
and U8268 (N_8268,N_7468,N_6824);
or U8269 (N_8269,N_5360,N_7487);
nand U8270 (N_8270,N_6583,N_5921);
and U8271 (N_8271,N_5078,N_5087);
nand U8272 (N_8272,N_5402,N_5714);
or U8273 (N_8273,N_7387,N_6752);
nand U8274 (N_8274,N_5355,N_5574);
xor U8275 (N_8275,N_5753,N_5481);
nand U8276 (N_8276,N_6287,N_5724);
and U8277 (N_8277,N_5480,N_7182);
nor U8278 (N_8278,N_7292,N_5821);
nand U8279 (N_8279,N_6375,N_6681);
or U8280 (N_8280,N_7337,N_6162);
or U8281 (N_8281,N_7476,N_5176);
xnor U8282 (N_8282,N_5158,N_7109);
and U8283 (N_8283,N_5392,N_6907);
nor U8284 (N_8284,N_6537,N_5500);
or U8285 (N_8285,N_6461,N_6094);
nor U8286 (N_8286,N_5330,N_5605);
and U8287 (N_8287,N_6124,N_6541);
nand U8288 (N_8288,N_6394,N_7126);
nor U8289 (N_8289,N_7482,N_5764);
nand U8290 (N_8290,N_6278,N_6741);
or U8291 (N_8291,N_6597,N_5064);
and U8292 (N_8292,N_7305,N_7189);
nand U8293 (N_8293,N_7210,N_5088);
and U8294 (N_8294,N_5317,N_6881);
and U8295 (N_8295,N_5790,N_5602);
nand U8296 (N_8296,N_6559,N_5558);
nand U8297 (N_8297,N_6353,N_5624);
nor U8298 (N_8298,N_7400,N_5202);
or U8299 (N_8299,N_5175,N_6536);
or U8300 (N_8300,N_6726,N_5399);
or U8301 (N_8301,N_5929,N_6444);
and U8302 (N_8302,N_6852,N_5747);
and U8303 (N_8303,N_5960,N_6137);
and U8304 (N_8304,N_7057,N_6459);
nand U8305 (N_8305,N_5279,N_6845);
nor U8306 (N_8306,N_5131,N_5479);
nor U8307 (N_8307,N_6183,N_6854);
nor U8308 (N_8308,N_5154,N_6001);
and U8309 (N_8309,N_6923,N_5167);
nand U8310 (N_8310,N_6493,N_5142);
or U8311 (N_8311,N_6228,N_6359);
or U8312 (N_8312,N_6534,N_6942);
and U8313 (N_8313,N_5898,N_5374);
or U8314 (N_8314,N_7202,N_7090);
nand U8315 (N_8315,N_6073,N_5005);
xor U8316 (N_8316,N_7445,N_6371);
nor U8317 (N_8317,N_7235,N_7489);
and U8318 (N_8318,N_7302,N_5848);
or U8319 (N_8319,N_7121,N_6246);
nor U8320 (N_8320,N_6293,N_5365);
or U8321 (N_8321,N_5876,N_6797);
xor U8322 (N_8322,N_5758,N_6876);
xor U8323 (N_8323,N_6216,N_7046);
xor U8324 (N_8324,N_7039,N_6932);
or U8325 (N_8325,N_5156,N_5645);
xnor U8326 (N_8326,N_5904,N_6152);
nor U8327 (N_8327,N_5161,N_7298);
or U8328 (N_8328,N_5140,N_6662);
or U8329 (N_8329,N_5243,N_5622);
nor U8330 (N_8330,N_6068,N_6031);
and U8331 (N_8331,N_5670,N_5212);
xor U8332 (N_8332,N_6584,N_6535);
and U8333 (N_8333,N_5395,N_5673);
xor U8334 (N_8334,N_7454,N_7047);
and U8335 (N_8335,N_6372,N_6012);
nor U8336 (N_8336,N_6608,N_6508);
xnor U8337 (N_8337,N_5567,N_5119);
nor U8338 (N_8338,N_7283,N_7128);
xnor U8339 (N_8339,N_7172,N_7033);
or U8340 (N_8340,N_5840,N_5282);
nand U8341 (N_8341,N_7133,N_5274);
and U8342 (N_8342,N_6972,N_5668);
nand U8343 (N_8343,N_5489,N_6669);
nor U8344 (N_8344,N_6830,N_6840);
and U8345 (N_8345,N_5809,N_7411);
or U8346 (N_8346,N_6685,N_5948);
or U8347 (N_8347,N_6441,N_7105);
nand U8348 (N_8348,N_7413,N_5013);
xor U8349 (N_8349,N_7457,N_5639);
xor U8350 (N_8350,N_5464,N_6470);
or U8351 (N_8351,N_7145,N_6039);
nand U8352 (N_8352,N_6596,N_7211);
and U8353 (N_8353,N_6773,N_5584);
or U8354 (N_8354,N_6514,N_5321);
and U8355 (N_8355,N_7401,N_7143);
and U8356 (N_8356,N_6033,N_5883);
xor U8357 (N_8357,N_6100,N_7226);
nand U8358 (N_8358,N_6912,N_6914);
nor U8359 (N_8359,N_5977,N_5561);
and U8360 (N_8360,N_7433,N_5684);
or U8361 (N_8361,N_5511,N_7364);
nand U8362 (N_8362,N_6632,N_6578);
xnor U8363 (N_8363,N_5630,N_5460);
nor U8364 (N_8364,N_6668,N_5337);
nor U8365 (N_8365,N_6788,N_6658);
xor U8366 (N_8366,N_6409,N_6021);
or U8367 (N_8367,N_7231,N_6141);
nand U8368 (N_8368,N_5872,N_5435);
and U8369 (N_8369,N_6551,N_5294);
or U8370 (N_8370,N_6525,N_5289);
xor U8371 (N_8371,N_7480,N_6114);
nand U8372 (N_8372,N_5179,N_5292);
and U8373 (N_8373,N_6383,N_5227);
or U8374 (N_8374,N_5593,N_5998);
or U8375 (N_8375,N_6320,N_7434);
or U8376 (N_8376,N_6833,N_6123);
xnor U8377 (N_8377,N_7497,N_5963);
xnor U8378 (N_8378,N_7069,N_5750);
nand U8379 (N_8379,N_5459,N_6218);
and U8380 (N_8380,N_7028,N_6519);
nand U8381 (N_8381,N_7215,N_7043);
nand U8382 (N_8382,N_6418,N_5203);
xor U8383 (N_8383,N_7238,N_5725);
nor U8384 (N_8384,N_6445,N_5383);
nor U8385 (N_8385,N_5834,N_5339);
xnor U8386 (N_8386,N_6723,N_6872);
or U8387 (N_8387,N_5260,N_5671);
xnor U8388 (N_8388,N_5746,N_5350);
nor U8389 (N_8389,N_7157,N_7247);
nand U8390 (N_8390,N_6247,N_5811);
xor U8391 (N_8391,N_5778,N_5553);
nand U8392 (N_8392,N_5702,N_6507);
nand U8393 (N_8393,N_6332,N_5406);
and U8394 (N_8394,N_6898,N_6205);
and U8395 (N_8395,N_6689,N_5039);
nand U8396 (N_8396,N_5691,N_5356);
nand U8397 (N_8397,N_7368,N_5881);
nand U8398 (N_8398,N_6185,N_5169);
nand U8399 (N_8399,N_6841,N_6602);
or U8400 (N_8400,N_6166,N_5896);
or U8401 (N_8401,N_6654,N_5308);
nand U8402 (N_8402,N_5918,N_5599);
xor U8403 (N_8403,N_6739,N_5268);
or U8404 (N_8404,N_6479,N_6783);
nand U8405 (N_8405,N_7031,N_5657);
nand U8406 (N_8406,N_6516,N_6677);
xnor U8407 (N_8407,N_5048,N_6067);
nor U8408 (N_8408,N_6808,N_5333);
or U8409 (N_8409,N_5093,N_5927);
xnor U8410 (N_8410,N_5261,N_7326);
xnor U8411 (N_8411,N_6874,N_6482);
or U8412 (N_8412,N_6860,N_5804);
or U8413 (N_8413,N_6310,N_7350);
or U8414 (N_8414,N_5214,N_5305);
nand U8415 (N_8415,N_7306,N_5346);
nor U8416 (N_8416,N_6321,N_5740);
or U8417 (N_8417,N_7114,N_7240);
nor U8418 (N_8418,N_6262,N_7002);
nor U8419 (N_8419,N_6388,N_6992);
nor U8420 (N_8420,N_6751,N_5055);
xnor U8421 (N_8421,N_6465,N_5427);
nand U8422 (N_8422,N_6879,N_5633);
and U8423 (N_8423,N_6929,N_6890);
xor U8424 (N_8424,N_7452,N_5254);
nor U8425 (N_8425,N_7474,N_5692);
xnor U8426 (N_8426,N_5071,N_7158);
nor U8427 (N_8427,N_5270,N_6055);
nand U8428 (N_8428,N_5455,N_5720);
nand U8429 (N_8429,N_6938,N_5106);
nand U8430 (N_8430,N_6678,N_6451);
and U8431 (N_8431,N_6091,N_6492);
xnor U8432 (N_8432,N_6712,N_5683);
nand U8433 (N_8433,N_5851,N_5830);
or U8434 (N_8434,N_5754,N_5494);
or U8435 (N_8435,N_7036,N_6504);
or U8436 (N_8436,N_5376,N_5361);
nand U8437 (N_8437,N_5543,N_5186);
xor U8438 (N_8438,N_6475,N_7051);
xor U8439 (N_8439,N_6544,N_5770);
xor U8440 (N_8440,N_6665,N_6469);
nand U8441 (N_8441,N_7258,N_5323);
or U8442 (N_8442,N_6777,N_6636);
nand U8443 (N_8443,N_6401,N_5507);
nand U8444 (N_8444,N_6893,N_5587);
xnor U8445 (N_8445,N_5445,N_5032);
xnor U8446 (N_8446,N_7407,N_7303);
xnor U8447 (N_8447,N_5731,N_6962);
nor U8448 (N_8448,N_5742,N_5713);
and U8449 (N_8449,N_5319,N_5548);
nand U8450 (N_8450,N_5264,N_6911);
nor U8451 (N_8451,N_6311,N_6042);
xor U8452 (N_8452,N_6816,N_5134);
nand U8453 (N_8453,N_6105,N_6734);
xnor U8454 (N_8454,N_7049,N_6735);
or U8455 (N_8455,N_5080,N_7151);
xnor U8456 (N_8456,N_7078,N_5603);
and U8457 (N_8457,N_6194,N_5564);
xnor U8458 (N_8458,N_7383,N_5791);
nor U8459 (N_8459,N_6082,N_6859);
and U8460 (N_8460,N_5663,N_6803);
xnor U8461 (N_8461,N_5332,N_6386);
nand U8462 (N_8462,N_6387,N_7272);
or U8463 (N_8463,N_6076,N_5617);
xor U8464 (N_8464,N_5086,N_5492);
or U8465 (N_8465,N_5936,N_5150);
nor U8466 (N_8466,N_5575,N_7136);
nand U8467 (N_8467,N_6713,N_5689);
nand U8468 (N_8468,N_5281,N_5027);
or U8469 (N_8469,N_6765,N_6237);
nand U8470 (N_8470,N_7354,N_7184);
nor U8471 (N_8471,N_6485,N_5079);
nor U8472 (N_8472,N_6330,N_7140);
nand U8473 (N_8473,N_5296,N_6882);
and U8474 (N_8474,N_6679,N_6985);
xor U8475 (N_8475,N_7402,N_5197);
and U8476 (N_8476,N_6593,N_5820);
or U8477 (N_8477,N_5600,N_5135);
and U8478 (N_8478,N_5797,N_6442);
nand U8479 (N_8479,N_5216,N_6644);
or U8480 (N_8480,N_6328,N_5320);
and U8481 (N_8481,N_5845,N_6842);
or U8482 (N_8482,N_7447,N_5094);
nand U8483 (N_8483,N_7092,N_7059);
xor U8484 (N_8484,N_6112,N_6412);
xnor U8485 (N_8485,N_5864,N_6299);
xor U8486 (N_8486,N_5551,N_6871);
or U8487 (N_8487,N_6056,N_6048);
xnor U8488 (N_8488,N_6986,N_5588);
xnor U8489 (N_8489,N_5276,N_6302);
or U8490 (N_8490,N_5609,N_5722);
and U8491 (N_8491,N_7360,N_7132);
xnor U8492 (N_8492,N_6834,N_5887);
or U8493 (N_8493,N_5159,N_7301);
nor U8494 (N_8494,N_6629,N_6413);
nand U8495 (N_8495,N_6955,N_5391);
or U8496 (N_8496,N_6886,N_5798);
xnor U8497 (N_8497,N_5800,N_6256);
or U8498 (N_8498,N_6464,N_5678);
nor U8499 (N_8499,N_6301,N_7080);
or U8500 (N_8500,N_5930,N_5959);
or U8501 (N_8501,N_7357,N_5384);
nor U8502 (N_8502,N_7135,N_6595);
and U8503 (N_8503,N_6245,N_7269);
nand U8504 (N_8504,N_5113,N_5954);
or U8505 (N_8505,N_6604,N_6558);
or U8506 (N_8506,N_5209,N_5123);
xnor U8507 (N_8507,N_5394,N_6906);
xor U8508 (N_8508,N_5634,N_5888);
nand U8509 (N_8509,N_7213,N_7207);
nor U8510 (N_8510,N_6784,N_7332);
xnor U8511 (N_8511,N_6097,N_6983);
and U8512 (N_8512,N_6555,N_6164);
xor U8513 (N_8513,N_5508,N_6190);
and U8514 (N_8514,N_6411,N_6878);
and U8515 (N_8515,N_6981,N_6250);
or U8516 (N_8516,N_5222,N_5338);
xnor U8517 (N_8517,N_7260,N_7201);
xor U8518 (N_8518,N_6499,N_6284);
xor U8519 (N_8519,N_5884,N_6251);
or U8520 (N_8520,N_5608,N_6934);
or U8521 (N_8521,N_7319,N_7287);
and U8522 (N_8522,N_5706,N_6510);
or U8523 (N_8523,N_7138,N_5606);
nand U8524 (N_8524,N_5329,N_5899);
xnor U8525 (N_8525,N_7125,N_6648);
or U8526 (N_8526,N_7426,N_7294);
or U8527 (N_8527,N_5557,N_6664);
nor U8528 (N_8528,N_6240,N_6702);
and U8529 (N_8529,N_7193,N_5313);
nand U8530 (N_8530,N_6180,N_7176);
nor U8531 (N_8531,N_5237,N_5244);
or U8532 (N_8532,N_6484,N_7318);
xnor U8533 (N_8533,N_6811,N_7453);
xor U8534 (N_8534,N_5141,N_7067);
or U8535 (N_8535,N_6134,N_7040);
and U8536 (N_8536,N_6453,N_5190);
nor U8537 (N_8537,N_6323,N_7127);
or U8538 (N_8538,N_6092,N_5033);
xnor U8539 (N_8539,N_5735,N_6846);
xnor U8540 (N_8540,N_6901,N_5265);
and U8541 (N_8541,N_6443,N_6150);
nor U8542 (N_8542,N_5868,N_6993);
xnor U8543 (N_8543,N_5822,N_5491);
or U8544 (N_8544,N_5266,N_6403);
nor U8545 (N_8545,N_5895,N_5072);
xnor U8546 (N_8546,N_7216,N_6037);
xnor U8547 (N_8547,N_6828,N_6910);
and U8548 (N_8548,N_6356,N_6718);
and U8549 (N_8549,N_6120,N_7448);
or U8550 (N_8550,N_5514,N_7348);
nor U8551 (N_8551,N_6006,N_6200);
xnor U8552 (N_8552,N_6577,N_5592);
xnor U8553 (N_8553,N_6711,N_5542);
nand U8554 (N_8554,N_5331,N_5982);
nor U8555 (N_8555,N_7491,N_7267);
nand U8556 (N_8556,N_5877,N_7484);
or U8557 (N_8557,N_5555,N_5610);
xnor U8558 (N_8558,N_6946,N_6280);
nor U8559 (N_8559,N_5781,N_5443);
nand U8560 (N_8560,N_5245,N_5517);
nand U8561 (N_8561,N_5751,N_7466);
xnor U8562 (N_8562,N_5866,N_5077);
nand U8563 (N_8563,N_7427,N_6707);
nor U8564 (N_8564,N_5867,N_6020);
nand U8565 (N_8565,N_5471,N_5823);
and U8566 (N_8566,N_5357,N_5862);
nand U8567 (N_8567,N_7490,N_7171);
and U8568 (N_8568,N_6988,N_5006);
nand U8569 (N_8569,N_6740,N_5604);
nor U8570 (N_8570,N_6553,N_6281);
and U8571 (N_8571,N_6837,N_5256);
nor U8572 (N_8572,N_6850,N_5659);
and U8573 (N_8573,N_6231,N_5589);
nand U8574 (N_8574,N_7492,N_6802);
xor U8575 (N_8575,N_6909,N_5239);
nand U8576 (N_8576,N_6326,N_6024);
and U8577 (N_8577,N_5806,N_6891);
nand U8578 (N_8578,N_5709,N_6761);
and U8579 (N_8579,N_6486,N_5686);
nand U8580 (N_8580,N_6877,N_6671);
and U8581 (N_8581,N_6297,N_5843);
or U8582 (N_8582,N_7378,N_6069);
nand U8583 (N_8583,N_5882,N_6800);
nand U8584 (N_8584,N_5328,N_7208);
xor U8585 (N_8585,N_7232,N_5535);
xnor U8586 (N_8586,N_7397,N_5715);
xnor U8587 (N_8587,N_7139,N_5970);
nand U8588 (N_8588,N_6341,N_5902);
nand U8589 (N_8589,N_6813,N_5301);
nand U8590 (N_8590,N_6399,N_7018);
nand U8591 (N_8591,N_5052,N_7098);
or U8592 (N_8592,N_6873,N_5996);
nor U8593 (N_8593,N_5306,N_5487);
or U8594 (N_8594,N_6352,N_6863);
and U8595 (N_8595,N_6424,N_7093);
nand U8596 (N_8596,N_5980,N_5944);
nor U8597 (N_8597,N_7323,N_6970);
and U8598 (N_8598,N_7421,N_5485);
and U8599 (N_8599,N_7280,N_6168);
or U8600 (N_8600,N_7278,N_7227);
nor U8601 (N_8601,N_5736,N_5889);
nand U8602 (N_8602,N_5675,N_6543);
xor U8603 (N_8603,N_6224,N_6023);
nor U8604 (N_8604,N_5343,N_5012);
and U8605 (N_8605,N_6308,N_5370);
or U8606 (N_8606,N_5304,N_5853);
nand U8607 (N_8607,N_5063,N_5987);
xnor U8608 (N_8608,N_5873,N_5397);
nor U8609 (N_8609,N_5694,N_6072);
nor U8610 (N_8610,N_6952,N_7122);
and U8611 (N_8611,N_6695,N_6722);
nand U8612 (N_8612,N_6990,N_6779);
or U8613 (N_8613,N_5446,N_6776);
nor U8614 (N_8614,N_5152,N_7429);
nand U8615 (N_8615,N_6259,N_6576);
xnor U8616 (N_8616,N_6736,N_6567);
nor U8617 (N_8617,N_5234,N_5920);
nand U8618 (N_8618,N_5415,N_6547);
xor U8619 (N_8619,N_6641,N_5108);
xnor U8620 (N_8620,N_5937,N_6452);
and U8621 (N_8621,N_6104,N_5336);
xor U8622 (N_8622,N_6646,N_5425);
nor U8623 (N_8623,N_5540,N_5066);
nand U8624 (N_8624,N_6306,N_7200);
nor U8625 (N_8625,N_5015,N_5196);
or U8626 (N_8626,N_5831,N_6003);
and U8627 (N_8627,N_6582,N_5327);
xor U8628 (N_8628,N_6093,N_6549);
xor U8629 (N_8629,N_6864,N_5839);
nor U8630 (N_8630,N_6506,N_7045);
nand U8631 (N_8631,N_6698,N_5749);
or U8632 (N_8632,N_6968,N_6697);
nand U8633 (N_8633,N_6758,N_6064);
nor U8634 (N_8634,N_6279,N_6143);
or U8635 (N_8635,N_6080,N_6272);
xnor U8636 (N_8636,N_5488,N_7146);
nor U8637 (N_8637,N_6743,N_5953);
or U8638 (N_8638,N_7062,N_6428);
nor U8639 (N_8639,N_5200,N_6821);
and U8640 (N_8640,N_6271,N_6329);
or U8641 (N_8641,N_5211,N_6017);
xor U8642 (N_8642,N_6904,N_5818);
or U8643 (N_8643,N_7254,N_5036);
nor U8644 (N_8644,N_5022,N_5257);
and U8645 (N_8645,N_6616,N_6849);
xor U8646 (N_8646,N_6643,N_5325);
or U8647 (N_8647,N_6182,N_6349);
and U8648 (N_8648,N_6456,N_6113);
nor U8649 (N_8649,N_5038,N_6933);
xnor U8650 (N_8650,N_6257,N_6533);
and U8651 (N_8651,N_5597,N_6377);
and U8652 (N_8652,N_7134,N_6342);
nand U8653 (N_8653,N_5635,N_7307);
xnor U8654 (N_8654,N_7408,N_6223);
nor U8655 (N_8655,N_7496,N_5900);
xor U8656 (N_8656,N_5817,N_7279);
xnor U8657 (N_8657,N_5975,N_6862);
xor U8658 (N_8658,N_6785,N_6102);
xnor U8659 (N_8659,N_6572,N_6494);
or U8660 (N_8660,N_7313,N_6417);
xnor U8661 (N_8661,N_5859,N_5095);
xor U8662 (N_8662,N_5933,N_5612);
nand U8663 (N_8663,N_6676,N_5596);
nand U8664 (N_8664,N_7096,N_6234);
or U8665 (N_8665,N_5393,N_6546);
or U8666 (N_8666,N_7314,N_7333);
nor U8667 (N_8667,N_6260,N_7129);
and U8668 (N_8668,N_7430,N_5162);
nor U8669 (N_8669,N_5752,N_7124);
nor U8670 (N_8670,N_7222,N_7441);
xnor U8671 (N_8671,N_5424,N_5769);
nor U8672 (N_8672,N_7329,N_5576);
or U8673 (N_8673,N_6729,N_7273);
nand U8674 (N_8674,N_5886,N_5885);
or U8675 (N_8675,N_7209,N_5275);
or U8676 (N_8676,N_5943,N_5554);
or U8677 (N_8677,N_7042,N_5483);
nand U8678 (N_8678,N_6920,N_5923);
and U8679 (N_8679,N_5451,N_5938);
nand U8680 (N_8680,N_6222,N_5098);
or U8681 (N_8681,N_7052,N_7131);
nand U8682 (N_8682,N_6731,N_5732);
or U8683 (N_8683,N_6633,N_6585);
and U8684 (N_8684,N_5945,N_5440);
xor U8685 (N_8685,N_6334,N_5958);
nand U8686 (N_8686,N_7369,N_7118);
nor U8687 (N_8687,N_5637,N_5651);
or U8688 (N_8688,N_6078,N_6590);
and U8689 (N_8689,N_6799,N_6615);
xnor U8690 (N_8690,N_5478,N_7223);
nor U8691 (N_8691,N_5844,N_7156);
or U8692 (N_8692,N_6000,N_5646);
or U8693 (N_8693,N_5220,N_5059);
nand U8694 (N_8694,N_5979,N_5405);
or U8695 (N_8695,N_5687,N_7410);
and U8696 (N_8696,N_6099,N_6016);
and U8697 (N_8697,N_5310,N_5509);
xor U8698 (N_8698,N_5412,N_5779);
xnor U8699 (N_8699,N_5833,N_6796);
xnor U8700 (N_8700,N_6659,N_6639);
xor U8701 (N_8701,N_5312,N_5563);
nand U8702 (N_8702,N_6538,N_5533);
and U8703 (N_8703,N_5506,N_7224);
xor U8704 (N_8704,N_6243,N_6344);
or U8705 (N_8705,N_5761,N_5638);
xnor U8706 (N_8706,N_7473,N_6144);
xor U8707 (N_8707,N_7277,N_5568);
and U8708 (N_8708,N_7472,N_7037);
nor U8709 (N_8709,N_7308,N_6748);
nand U8710 (N_8710,N_6285,N_5056);
nor U8711 (N_8711,N_7072,N_5493);
xor U8712 (N_8712,N_5431,N_5128);
xor U8713 (N_8713,N_6238,N_7014);
nor U8714 (N_8714,N_5201,N_7431);
or U8715 (N_8715,N_6345,N_7241);
nand U8716 (N_8716,N_5398,N_6404);
xor U8717 (N_8717,N_5126,N_5484);
nor U8718 (N_8718,N_5353,N_5573);
xor U8719 (N_8719,N_6975,N_6717);
nor U8720 (N_8720,N_7327,N_5983);
nand U8721 (N_8721,N_5285,N_6903);
xnor U8722 (N_8722,N_7179,N_6044);
nor U8723 (N_8723,N_5733,N_6170);
and U8724 (N_8724,N_5771,N_6794);
nor U8725 (N_8725,N_5291,N_5037);
xor U8726 (N_8726,N_5110,N_5248);
nor U8727 (N_8727,N_6436,N_7025);
and U8728 (N_8728,N_6288,N_6588);
nand U8729 (N_8729,N_5792,N_6360);
and U8730 (N_8730,N_5803,N_5526);
nor U8731 (N_8731,N_6154,N_6004);
nor U8732 (N_8732,N_6782,N_6460);
xor U8733 (N_8733,N_5137,N_7107);
and U8734 (N_8734,N_6426,N_5538);
nand U8735 (N_8735,N_5734,N_6149);
nor U8736 (N_8736,N_5942,N_6497);
nand U8737 (N_8737,N_5795,N_7390);
nand U8738 (N_8738,N_6959,N_5704);
and U8739 (N_8739,N_6066,N_6370);
and U8740 (N_8740,N_6128,N_5057);
nand U8741 (N_8741,N_6666,N_5649);
or U8742 (N_8742,N_6941,N_6887);
xor U8743 (N_8743,N_6169,N_6438);
and U8744 (N_8744,N_6083,N_7008);
and U8745 (N_8745,N_5476,N_6338);
and U8746 (N_8746,N_6556,N_6822);
and U8747 (N_8747,N_5513,N_5082);
and U8748 (N_8748,N_7419,N_6737);
nor U8749 (N_8749,N_6477,N_7180);
and U8750 (N_8750,N_5642,N_7461);
xor U8751 (N_8751,N_6908,N_6209);
xnor U8752 (N_8752,N_6766,N_7391);
nand U8753 (N_8753,N_6314,N_6040);
xnor U8754 (N_8754,N_6900,N_5785);
xnor U8755 (N_8755,N_6123,N_6103);
xnor U8756 (N_8756,N_5833,N_5630);
xor U8757 (N_8757,N_6999,N_6084);
xnor U8758 (N_8758,N_6512,N_7481);
and U8759 (N_8759,N_6170,N_5494);
and U8760 (N_8760,N_6755,N_7169);
nor U8761 (N_8761,N_6894,N_6837);
nand U8762 (N_8762,N_5628,N_7024);
xnor U8763 (N_8763,N_5855,N_5207);
and U8764 (N_8764,N_6486,N_5639);
xor U8765 (N_8765,N_6831,N_7033);
and U8766 (N_8766,N_5125,N_7403);
xnor U8767 (N_8767,N_6561,N_6146);
and U8768 (N_8768,N_5626,N_5460);
nand U8769 (N_8769,N_6517,N_5048);
xnor U8770 (N_8770,N_6000,N_6045);
nand U8771 (N_8771,N_5889,N_5603);
and U8772 (N_8772,N_5874,N_5341);
and U8773 (N_8773,N_7108,N_5333);
nand U8774 (N_8774,N_6542,N_6633);
nor U8775 (N_8775,N_6466,N_5717);
nand U8776 (N_8776,N_5090,N_6214);
and U8777 (N_8777,N_7169,N_5196);
xor U8778 (N_8778,N_7256,N_5973);
and U8779 (N_8779,N_6395,N_5029);
nor U8780 (N_8780,N_5945,N_5924);
nand U8781 (N_8781,N_5696,N_6671);
xnor U8782 (N_8782,N_5363,N_7283);
and U8783 (N_8783,N_5409,N_7044);
nand U8784 (N_8784,N_5924,N_5518);
and U8785 (N_8785,N_6751,N_6797);
nor U8786 (N_8786,N_5872,N_7148);
nand U8787 (N_8787,N_6499,N_5122);
nor U8788 (N_8788,N_7101,N_6666);
xnor U8789 (N_8789,N_7447,N_5621);
and U8790 (N_8790,N_6678,N_5829);
nand U8791 (N_8791,N_5735,N_6214);
xnor U8792 (N_8792,N_6292,N_7318);
nand U8793 (N_8793,N_6837,N_6081);
and U8794 (N_8794,N_6866,N_5590);
nor U8795 (N_8795,N_6981,N_5078);
nand U8796 (N_8796,N_6108,N_6169);
xnor U8797 (N_8797,N_7321,N_6174);
and U8798 (N_8798,N_6938,N_6210);
xnor U8799 (N_8799,N_7473,N_5912);
nand U8800 (N_8800,N_5759,N_6811);
xnor U8801 (N_8801,N_7037,N_5970);
and U8802 (N_8802,N_6633,N_6928);
xnor U8803 (N_8803,N_5279,N_6402);
nand U8804 (N_8804,N_6049,N_5243);
and U8805 (N_8805,N_5523,N_6982);
or U8806 (N_8806,N_5613,N_5996);
or U8807 (N_8807,N_5800,N_7016);
xor U8808 (N_8808,N_6793,N_7430);
or U8809 (N_8809,N_7253,N_7350);
nor U8810 (N_8810,N_5662,N_6520);
and U8811 (N_8811,N_5123,N_6602);
nand U8812 (N_8812,N_5479,N_7165);
or U8813 (N_8813,N_7034,N_7319);
nand U8814 (N_8814,N_5698,N_6426);
and U8815 (N_8815,N_6016,N_6621);
nor U8816 (N_8816,N_6484,N_5982);
nand U8817 (N_8817,N_6423,N_6660);
xnor U8818 (N_8818,N_5969,N_6968);
nand U8819 (N_8819,N_5048,N_6122);
and U8820 (N_8820,N_5210,N_5632);
and U8821 (N_8821,N_6023,N_5691);
nand U8822 (N_8822,N_7419,N_6678);
and U8823 (N_8823,N_7211,N_6799);
xnor U8824 (N_8824,N_6602,N_5068);
or U8825 (N_8825,N_6754,N_6680);
and U8826 (N_8826,N_6459,N_7426);
and U8827 (N_8827,N_7260,N_5659);
and U8828 (N_8828,N_6934,N_7165);
xnor U8829 (N_8829,N_5078,N_6501);
or U8830 (N_8830,N_5150,N_7464);
nor U8831 (N_8831,N_7107,N_6324);
nand U8832 (N_8832,N_5106,N_5713);
xor U8833 (N_8833,N_7178,N_5049);
nand U8834 (N_8834,N_5081,N_6966);
and U8835 (N_8835,N_7111,N_5704);
and U8836 (N_8836,N_6117,N_6186);
nor U8837 (N_8837,N_6963,N_5996);
and U8838 (N_8838,N_6544,N_7364);
and U8839 (N_8839,N_5421,N_6986);
or U8840 (N_8840,N_6319,N_7328);
or U8841 (N_8841,N_6230,N_6021);
nor U8842 (N_8842,N_6296,N_7161);
or U8843 (N_8843,N_6147,N_5693);
nor U8844 (N_8844,N_5827,N_7017);
or U8845 (N_8845,N_5436,N_5692);
xnor U8846 (N_8846,N_7229,N_6304);
nand U8847 (N_8847,N_7116,N_6296);
nor U8848 (N_8848,N_5330,N_6930);
nand U8849 (N_8849,N_6102,N_5419);
nor U8850 (N_8850,N_5021,N_6736);
nand U8851 (N_8851,N_5446,N_6159);
or U8852 (N_8852,N_7455,N_5487);
nor U8853 (N_8853,N_6476,N_5658);
or U8854 (N_8854,N_5332,N_7064);
xnor U8855 (N_8855,N_5935,N_7267);
or U8856 (N_8856,N_5391,N_5183);
and U8857 (N_8857,N_5221,N_6449);
xnor U8858 (N_8858,N_7440,N_6451);
xor U8859 (N_8859,N_7403,N_5678);
or U8860 (N_8860,N_6813,N_7362);
nor U8861 (N_8861,N_5790,N_6621);
xor U8862 (N_8862,N_6287,N_7297);
and U8863 (N_8863,N_7276,N_7478);
and U8864 (N_8864,N_6581,N_5231);
or U8865 (N_8865,N_5169,N_6532);
or U8866 (N_8866,N_7236,N_7271);
and U8867 (N_8867,N_5764,N_6590);
nand U8868 (N_8868,N_6061,N_6798);
nand U8869 (N_8869,N_7023,N_6983);
nor U8870 (N_8870,N_6403,N_5289);
nand U8871 (N_8871,N_5018,N_5599);
or U8872 (N_8872,N_6959,N_7130);
or U8873 (N_8873,N_6956,N_5876);
and U8874 (N_8874,N_6243,N_7090);
nor U8875 (N_8875,N_6999,N_5548);
or U8876 (N_8876,N_5394,N_5743);
nor U8877 (N_8877,N_6673,N_5802);
nand U8878 (N_8878,N_7458,N_6907);
nor U8879 (N_8879,N_6128,N_7033);
nor U8880 (N_8880,N_6641,N_6601);
and U8881 (N_8881,N_5745,N_5785);
or U8882 (N_8882,N_6423,N_6865);
nor U8883 (N_8883,N_5540,N_6417);
xor U8884 (N_8884,N_5525,N_5251);
nand U8885 (N_8885,N_6520,N_5134);
xnor U8886 (N_8886,N_7314,N_6244);
xnor U8887 (N_8887,N_7242,N_6918);
nand U8888 (N_8888,N_5199,N_5763);
and U8889 (N_8889,N_6417,N_6989);
xor U8890 (N_8890,N_5823,N_6280);
nand U8891 (N_8891,N_6364,N_6328);
and U8892 (N_8892,N_6935,N_5826);
xor U8893 (N_8893,N_6212,N_7127);
nand U8894 (N_8894,N_6839,N_5243);
nor U8895 (N_8895,N_6412,N_6600);
xor U8896 (N_8896,N_5212,N_7373);
xnor U8897 (N_8897,N_6026,N_6408);
or U8898 (N_8898,N_6545,N_5654);
and U8899 (N_8899,N_5464,N_5051);
nand U8900 (N_8900,N_5927,N_5448);
or U8901 (N_8901,N_7148,N_5632);
nand U8902 (N_8902,N_6096,N_5685);
xor U8903 (N_8903,N_6660,N_6240);
xor U8904 (N_8904,N_5781,N_6927);
nand U8905 (N_8905,N_7473,N_5586);
and U8906 (N_8906,N_5586,N_5704);
nand U8907 (N_8907,N_6545,N_5967);
nand U8908 (N_8908,N_7135,N_5230);
or U8909 (N_8909,N_7457,N_5095);
nand U8910 (N_8910,N_5044,N_6933);
nor U8911 (N_8911,N_5507,N_5634);
nand U8912 (N_8912,N_6923,N_7188);
xnor U8913 (N_8913,N_5482,N_7092);
xor U8914 (N_8914,N_5989,N_5099);
and U8915 (N_8915,N_6956,N_5321);
nor U8916 (N_8916,N_6330,N_5812);
or U8917 (N_8917,N_5793,N_6101);
and U8918 (N_8918,N_7113,N_7224);
and U8919 (N_8919,N_6781,N_5506);
xor U8920 (N_8920,N_5022,N_5340);
xor U8921 (N_8921,N_5235,N_7079);
nor U8922 (N_8922,N_7341,N_5741);
xnor U8923 (N_8923,N_6844,N_6276);
and U8924 (N_8924,N_6625,N_5998);
and U8925 (N_8925,N_5390,N_6309);
xor U8926 (N_8926,N_7044,N_6424);
nand U8927 (N_8927,N_5368,N_5119);
nand U8928 (N_8928,N_6970,N_6085);
xnor U8929 (N_8929,N_6743,N_6239);
nor U8930 (N_8930,N_5246,N_5435);
nand U8931 (N_8931,N_6684,N_7219);
nand U8932 (N_8932,N_5044,N_6374);
xor U8933 (N_8933,N_6897,N_6014);
and U8934 (N_8934,N_6342,N_7379);
xnor U8935 (N_8935,N_7167,N_6502);
or U8936 (N_8936,N_5751,N_5919);
nand U8937 (N_8937,N_6013,N_7374);
and U8938 (N_8938,N_6396,N_6972);
nand U8939 (N_8939,N_5190,N_5951);
or U8940 (N_8940,N_5276,N_6681);
or U8941 (N_8941,N_6079,N_7400);
xor U8942 (N_8942,N_7106,N_6494);
xnor U8943 (N_8943,N_5549,N_5860);
and U8944 (N_8944,N_5837,N_6605);
nor U8945 (N_8945,N_5119,N_5797);
or U8946 (N_8946,N_6101,N_5973);
or U8947 (N_8947,N_6041,N_5501);
xnor U8948 (N_8948,N_6051,N_6131);
and U8949 (N_8949,N_6849,N_6520);
nor U8950 (N_8950,N_5260,N_7243);
nor U8951 (N_8951,N_7226,N_6229);
and U8952 (N_8952,N_7068,N_5873);
xnor U8953 (N_8953,N_5083,N_5592);
and U8954 (N_8954,N_6016,N_7058);
and U8955 (N_8955,N_6485,N_6327);
xor U8956 (N_8956,N_6968,N_6002);
nor U8957 (N_8957,N_5738,N_6474);
and U8958 (N_8958,N_6586,N_6827);
xor U8959 (N_8959,N_5616,N_7298);
nor U8960 (N_8960,N_6161,N_7428);
nor U8961 (N_8961,N_5089,N_7180);
nor U8962 (N_8962,N_6383,N_5610);
nand U8963 (N_8963,N_5868,N_5021);
xnor U8964 (N_8964,N_5510,N_6134);
and U8965 (N_8965,N_6347,N_7284);
nor U8966 (N_8966,N_6354,N_5929);
nor U8967 (N_8967,N_7269,N_5492);
and U8968 (N_8968,N_6335,N_6628);
nand U8969 (N_8969,N_6574,N_5329);
nor U8970 (N_8970,N_7187,N_5502);
nand U8971 (N_8971,N_6729,N_5138);
and U8972 (N_8972,N_6242,N_6094);
and U8973 (N_8973,N_6273,N_6525);
or U8974 (N_8974,N_6819,N_6195);
xor U8975 (N_8975,N_6143,N_6322);
nand U8976 (N_8976,N_6422,N_6801);
nor U8977 (N_8977,N_5844,N_6654);
and U8978 (N_8978,N_5704,N_5064);
and U8979 (N_8979,N_5178,N_6018);
nor U8980 (N_8980,N_5333,N_6801);
and U8981 (N_8981,N_5869,N_7371);
xnor U8982 (N_8982,N_5565,N_5894);
xnor U8983 (N_8983,N_6312,N_6609);
and U8984 (N_8984,N_7014,N_6825);
xor U8985 (N_8985,N_7223,N_5968);
and U8986 (N_8986,N_7191,N_5917);
nand U8987 (N_8987,N_6631,N_5674);
xnor U8988 (N_8988,N_6244,N_5818);
nand U8989 (N_8989,N_6863,N_7155);
nand U8990 (N_8990,N_7457,N_6800);
and U8991 (N_8991,N_5881,N_7134);
and U8992 (N_8992,N_6756,N_6512);
or U8993 (N_8993,N_6024,N_5811);
nand U8994 (N_8994,N_5165,N_6859);
or U8995 (N_8995,N_7464,N_6753);
nor U8996 (N_8996,N_5354,N_6946);
nand U8997 (N_8997,N_5887,N_5100);
and U8998 (N_8998,N_6180,N_5812);
nand U8999 (N_8999,N_6859,N_7292);
xor U9000 (N_9000,N_5681,N_6465);
or U9001 (N_9001,N_6380,N_6147);
xnor U9002 (N_9002,N_5800,N_7248);
or U9003 (N_9003,N_5496,N_6717);
nor U9004 (N_9004,N_6493,N_7179);
nand U9005 (N_9005,N_5138,N_5161);
nor U9006 (N_9006,N_6349,N_6036);
or U9007 (N_9007,N_6480,N_6349);
or U9008 (N_9008,N_5322,N_5076);
nand U9009 (N_9009,N_6542,N_6981);
or U9010 (N_9010,N_5248,N_6056);
nand U9011 (N_9011,N_7040,N_6095);
or U9012 (N_9012,N_7334,N_5190);
or U9013 (N_9013,N_5972,N_6316);
and U9014 (N_9014,N_5807,N_6665);
or U9015 (N_9015,N_5682,N_5513);
or U9016 (N_9016,N_6372,N_6826);
xnor U9017 (N_9017,N_5061,N_5156);
or U9018 (N_9018,N_6244,N_5164);
nor U9019 (N_9019,N_5888,N_6831);
nor U9020 (N_9020,N_6831,N_7261);
and U9021 (N_9021,N_6134,N_5878);
and U9022 (N_9022,N_5143,N_5728);
and U9023 (N_9023,N_7281,N_5058);
and U9024 (N_9024,N_7473,N_5768);
or U9025 (N_9025,N_6486,N_5183);
and U9026 (N_9026,N_5495,N_6402);
and U9027 (N_9027,N_6345,N_6834);
and U9028 (N_9028,N_5049,N_6244);
and U9029 (N_9029,N_5308,N_7083);
or U9030 (N_9030,N_7145,N_5601);
nor U9031 (N_9031,N_6140,N_5152);
xor U9032 (N_9032,N_6372,N_7372);
and U9033 (N_9033,N_5754,N_5604);
nand U9034 (N_9034,N_6525,N_6632);
and U9035 (N_9035,N_5192,N_7040);
nand U9036 (N_9036,N_7236,N_5315);
and U9037 (N_9037,N_7010,N_6037);
nand U9038 (N_9038,N_6575,N_5603);
or U9039 (N_9039,N_5184,N_5403);
xnor U9040 (N_9040,N_5379,N_6079);
and U9041 (N_9041,N_7408,N_6549);
nand U9042 (N_9042,N_5372,N_5280);
or U9043 (N_9043,N_5584,N_7058);
nor U9044 (N_9044,N_5087,N_5590);
nor U9045 (N_9045,N_6572,N_7419);
or U9046 (N_9046,N_7363,N_5892);
and U9047 (N_9047,N_5703,N_5949);
xor U9048 (N_9048,N_5619,N_6889);
nand U9049 (N_9049,N_6943,N_7164);
nor U9050 (N_9050,N_5273,N_7034);
xor U9051 (N_9051,N_7125,N_5307);
and U9052 (N_9052,N_7397,N_7367);
or U9053 (N_9053,N_5639,N_6821);
nand U9054 (N_9054,N_5746,N_5294);
nand U9055 (N_9055,N_5556,N_7469);
and U9056 (N_9056,N_6744,N_5340);
and U9057 (N_9057,N_5693,N_7462);
xnor U9058 (N_9058,N_6050,N_7291);
nor U9059 (N_9059,N_6893,N_6494);
or U9060 (N_9060,N_6305,N_7384);
and U9061 (N_9061,N_7471,N_7232);
nor U9062 (N_9062,N_6374,N_7290);
nor U9063 (N_9063,N_7046,N_7348);
xnor U9064 (N_9064,N_5346,N_7352);
nor U9065 (N_9065,N_5978,N_6502);
and U9066 (N_9066,N_5981,N_6342);
nor U9067 (N_9067,N_5815,N_7006);
or U9068 (N_9068,N_6175,N_7498);
nand U9069 (N_9069,N_5662,N_5433);
nor U9070 (N_9070,N_6874,N_5786);
xnor U9071 (N_9071,N_5608,N_6806);
xor U9072 (N_9072,N_5429,N_5464);
and U9073 (N_9073,N_5185,N_7277);
and U9074 (N_9074,N_6062,N_7329);
or U9075 (N_9075,N_5050,N_6441);
or U9076 (N_9076,N_6953,N_5078);
nor U9077 (N_9077,N_6427,N_6299);
nor U9078 (N_9078,N_7250,N_6250);
xnor U9079 (N_9079,N_7329,N_5691);
nor U9080 (N_9080,N_5823,N_5250);
and U9081 (N_9081,N_5418,N_7151);
and U9082 (N_9082,N_6292,N_6296);
or U9083 (N_9083,N_6519,N_6953);
nand U9084 (N_9084,N_6967,N_5416);
nand U9085 (N_9085,N_5515,N_5123);
and U9086 (N_9086,N_7363,N_6459);
and U9087 (N_9087,N_6801,N_5117);
nand U9088 (N_9088,N_6910,N_7002);
and U9089 (N_9089,N_5972,N_6598);
xor U9090 (N_9090,N_6509,N_7128);
and U9091 (N_9091,N_5159,N_6572);
or U9092 (N_9092,N_5573,N_6456);
xor U9093 (N_9093,N_6536,N_5418);
nor U9094 (N_9094,N_6517,N_6135);
nor U9095 (N_9095,N_7125,N_7430);
or U9096 (N_9096,N_5035,N_5710);
nor U9097 (N_9097,N_6047,N_5282);
or U9098 (N_9098,N_7300,N_5933);
nand U9099 (N_9099,N_6590,N_5554);
nor U9100 (N_9100,N_6717,N_5773);
nand U9101 (N_9101,N_5568,N_5869);
xnor U9102 (N_9102,N_7061,N_7158);
nand U9103 (N_9103,N_5109,N_5990);
nand U9104 (N_9104,N_7247,N_5460);
and U9105 (N_9105,N_5773,N_5671);
nor U9106 (N_9106,N_7369,N_6228);
or U9107 (N_9107,N_6780,N_6486);
or U9108 (N_9108,N_7117,N_7143);
xor U9109 (N_9109,N_7338,N_5780);
nor U9110 (N_9110,N_6730,N_6679);
nor U9111 (N_9111,N_7007,N_5400);
nor U9112 (N_9112,N_6616,N_6109);
or U9113 (N_9113,N_6272,N_6459);
nand U9114 (N_9114,N_5877,N_6136);
and U9115 (N_9115,N_7481,N_7411);
nor U9116 (N_9116,N_7453,N_7188);
and U9117 (N_9117,N_6622,N_5590);
or U9118 (N_9118,N_7148,N_6787);
and U9119 (N_9119,N_6924,N_5353);
nor U9120 (N_9120,N_7115,N_5309);
nor U9121 (N_9121,N_5786,N_7191);
xor U9122 (N_9122,N_7183,N_6092);
xnor U9123 (N_9123,N_6323,N_5285);
nor U9124 (N_9124,N_5496,N_6872);
nor U9125 (N_9125,N_7181,N_6200);
xor U9126 (N_9126,N_6572,N_7303);
or U9127 (N_9127,N_5184,N_5156);
and U9128 (N_9128,N_6402,N_7161);
or U9129 (N_9129,N_6392,N_6803);
nand U9130 (N_9130,N_7439,N_7077);
nor U9131 (N_9131,N_5687,N_5324);
xor U9132 (N_9132,N_5774,N_5627);
nor U9133 (N_9133,N_5162,N_5085);
xor U9134 (N_9134,N_5980,N_7260);
nand U9135 (N_9135,N_6967,N_6138);
nor U9136 (N_9136,N_5462,N_6928);
nor U9137 (N_9137,N_5626,N_7235);
nor U9138 (N_9138,N_5757,N_7438);
xor U9139 (N_9139,N_5443,N_6287);
nand U9140 (N_9140,N_7271,N_5793);
xor U9141 (N_9141,N_6677,N_7409);
or U9142 (N_9142,N_6339,N_5608);
nand U9143 (N_9143,N_5797,N_5692);
xor U9144 (N_9144,N_6264,N_7354);
nor U9145 (N_9145,N_5809,N_6759);
or U9146 (N_9146,N_6473,N_5539);
nand U9147 (N_9147,N_5835,N_5450);
nor U9148 (N_9148,N_6040,N_7490);
nor U9149 (N_9149,N_6265,N_6799);
nor U9150 (N_9150,N_5419,N_6341);
or U9151 (N_9151,N_5457,N_5432);
nand U9152 (N_9152,N_6045,N_6943);
and U9153 (N_9153,N_6836,N_6067);
xor U9154 (N_9154,N_6190,N_7060);
or U9155 (N_9155,N_6539,N_6929);
and U9156 (N_9156,N_7286,N_7443);
nor U9157 (N_9157,N_5105,N_5345);
xnor U9158 (N_9158,N_7017,N_5230);
nor U9159 (N_9159,N_6745,N_5394);
xor U9160 (N_9160,N_5736,N_6847);
nand U9161 (N_9161,N_6547,N_5017);
xnor U9162 (N_9162,N_6221,N_7081);
nor U9163 (N_9163,N_6334,N_5416);
xnor U9164 (N_9164,N_5206,N_5768);
xor U9165 (N_9165,N_6812,N_7157);
nand U9166 (N_9166,N_5345,N_5587);
xnor U9167 (N_9167,N_6034,N_6537);
xnor U9168 (N_9168,N_6836,N_6068);
xor U9169 (N_9169,N_6463,N_5325);
and U9170 (N_9170,N_6771,N_7208);
nor U9171 (N_9171,N_6885,N_5029);
xnor U9172 (N_9172,N_6343,N_5236);
xnor U9173 (N_9173,N_6260,N_5452);
xor U9174 (N_9174,N_5900,N_5214);
and U9175 (N_9175,N_5450,N_6002);
or U9176 (N_9176,N_5720,N_7033);
xor U9177 (N_9177,N_7403,N_6298);
xor U9178 (N_9178,N_6205,N_6097);
and U9179 (N_9179,N_5262,N_5079);
nor U9180 (N_9180,N_7272,N_6767);
nor U9181 (N_9181,N_5985,N_5749);
xor U9182 (N_9182,N_5240,N_5736);
xor U9183 (N_9183,N_5694,N_5578);
nand U9184 (N_9184,N_6486,N_6197);
and U9185 (N_9185,N_6991,N_6309);
or U9186 (N_9186,N_5066,N_5178);
or U9187 (N_9187,N_5201,N_5919);
xor U9188 (N_9188,N_7227,N_6275);
nor U9189 (N_9189,N_5776,N_5455);
xnor U9190 (N_9190,N_5843,N_5803);
nor U9191 (N_9191,N_6235,N_5387);
nand U9192 (N_9192,N_6754,N_5379);
or U9193 (N_9193,N_6721,N_6654);
nor U9194 (N_9194,N_6572,N_5215);
and U9195 (N_9195,N_7194,N_5398);
nand U9196 (N_9196,N_7234,N_5918);
xnor U9197 (N_9197,N_6936,N_7112);
or U9198 (N_9198,N_5086,N_5640);
or U9199 (N_9199,N_5438,N_7063);
nand U9200 (N_9200,N_7064,N_6646);
nor U9201 (N_9201,N_6725,N_6756);
xor U9202 (N_9202,N_7323,N_6418);
nor U9203 (N_9203,N_5154,N_5810);
and U9204 (N_9204,N_6157,N_5506);
and U9205 (N_9205,N_5695,N_6655);
and U9206 (N_9206,N_5361,N_5382);
or U9207 (N_9207,N_6189,N_5867);
xor U9208 (N_9208,N_6959,N_6110);
nor U9209 (N_9209,N_6361,N_6721);
or U9210 (N_9210,N_5095,N_5544);
or U9211 (N_9211,N_5204,N_5689);
nand U9212 (N_9212,N_5545,N_6475);
nor U9213 (N_9213,N_5281,N_5179);
xor U9214 (N_9214,N_6351,N_6784);
nand U9215 (N_9215,N_6734,N_7090);
or U9216 (N_9216,N_7454,N_7476);
and U9217 (N_9217,N_5748,N_5205);
and U9218 (N_9218,N_5492,N_6841);
or U9219 (N_9219,N_5081,N_7293);
xnor U9220 (N_9220,N_5554,N_7000);
nand U9221 (N_9221,N_7080,N_5822);
or U9222 (N_9222,N_5037,N_6644);
or U9223 (N_9223,N_7191,N_6767);
nand U9224 (N_9224,N_6488,N_5261);
or U9225 (N_9225,N_5494,N_7144);
xnor U9226 (N_9226,N_5467,N_7263);
xor U9227 (N_9227,N_7132,N_7173);
nor U9228 (N_9228,N_7311,N_7319);
xnor U9229 (N_9229,N_5803,N_5003);
and U9230 (N_9230,N_6963,N_5831);
nor U9231 (N_9231,N_6473,N_5955);
and U9232 (N_9232,N_6344,N_6509);
nand U9233 (N_9233,N_5717,N_6626);
and U9234 (N_9234,N_6522,N_6334);
nor U9235 (N_9235,N_5275,N_6996);
nor U9236 (N_9236,N_6016,N_6143);
xnor U9237 (N_9237,N_6872,N_5175);
nand U9238 (N_9238,N_5686,N_7065);
or U9239 (N_9239,N_5476,N_6583);
and U9240 (N_9240,N_7405,N_5310);
or U9241 (N_9241,N_7393,N_5051);
xnor U9242 (N_9242,N_6969,N_6202);
nand U9243 (N_9243,N_5764,N_6359);
or U9244 (N_9244,N_7245,N_6566);
nor U9245 (N_9245,N_5952,N_7245);
and U9246 (N_9246,N_5969,N_5344);
or U9247 (N_9247,N_6974,N_6583);
xnor U9248 (N_9248,N_6991,N_5343);
nor U9249 (N_9249,N_5836,N_6830);
or U9250 (N_9250,N_5341,N_5754);
nand U9251 (N_9251,N_6009,N_6586);
or U9252 (N_9252,N_5106,N_5703);
and U9253 (N_9253,N_7215,N_5519);
nand U9254 (N_9254,N_5185,N_5705);
and U9255 (N_9255,N_5704,N_6726);
or U9256 (N_9256,N_6423,N_6441);
and U9257 (N_9257,N_6520,N_5073);
xor U9258 (N_9258,N_6201,N_5450);
xor U9259 (N_9259,N_5456,N_5505);
nor U9260 (N_9260,N_6607,N_6420);
nand U9261 (N_9261,N_7431,N_6935);
xor U9262 (N_9262,N_7430,N_5018);
nor U9263 (N_9263,N_5431,N_5325);
nand U9264 (N_9264,N_7472,N_5106);
or U9265 (N_9265,N_5663,N_5685);
nand U9266 (N_9266,N_5845,N_6430);
or U9267 (N_9267,N_7126,N_5508);
and U9268 (N_9268,N_6670,N_6936);
nor U9269 (N_9269,N_5205,N_5823);
or U9270 (N_9270,N_7173,N_5930);
nand U9271 (N_9271,N_7431,N_6701);
nand U9272 (N_9272,N_6370,N_5366);
nand U9273 (N_9273,N_6630,N_6502);
xor U9274 (N_9274,N_6710,N_6309);
nand U9275 (N_9275,N_5575,N_7413);
nand U9276 (N_9276,N_5827,N_7097);
and U9277 (N_9277,N_5868,N_6154);
nor U9278 (N_9278,N_7202,N_7314);
and U9279 (N_9279,N_6827,N_6871);
and U9280 (N_9280,N_5623,N_6375);
nor U9281 (N_9281,N_5548,N_7119);
nor U9282 (N_9282,N_5745,N_5802);
nor U9283 (N_9283,N_6240,N_5888);
nor U9284 (N_9284,N_5573,N_5263);
xnor U9285 (N_9285,N_5764,N_7361);
nor U9286 (N_9286,N_5258,N_5675);
nand U9287 (N_9287,N_6283,N_6287);
or U9288 (N_9288,N_5159,N_6409);
nand U9289 (N_9289,N_5294,N_7368);
and U9290 (N_9290,N_6668,N_5322);
nor U9291 (N_9291,N_6101,N_7093);
and U9292 (N_9292,N_7069,N_7144);
and U9293 (N_9293,N_6470,N_6692);
and U9294 (N_9294,N_5543,N_7115);
nor U9295 (N_9295,N_6818,N_6422);
nor U9296 (N_9296,N_6910,N_7254);
nor U9297 (N_9297,N_6876,N_6120);
nor U9298 (N_9298,N_5566,N_6580);
and U9299 (N_9299,N_5197,N_5665);
and U9300 (N_9300,N_7139,N_7040);
nand U9301 (N_9301,N_6069,N_6649);
xnor U9302 (N_9302,N_5334,N_7356);
nand U9303 (N_9303,N_7326,N_7095);
and U9304 (N_9304,N_6337,N_6279);
nor U9305 (N_9305,N_5814,N_6479);
nand U9306 (N_9306,N_5079,N_6237);
or U9307 (N_9307,N_7207,N_6138);
xnor U9308 (N_9308,N_7158,N_7004);
or U9309 (N_9309,N_6545,N_7376);
nor U9310 (N_9310,N_5652,N_5845);
xor U9311 (N_9311,N_5455,N_5175);
nor U9312 (N_9312,N_5015,N_5665);
and U9313 (N_9313,N_6280,N_5719);
or U9314 (N_9314,N_6235,N_7326);
xor U9315 (N_9315,N_6902,N_6795);
and U9316 (N_9316,N_6592,N_5419);
xnor U9317 (N_9317,N_5114,N_6404);
and U9318 (N_9318,N_7075,N_6036);
or U9319 (N_9319,N_5319,N_5259);
nor U9320 (N_9320,N_6775,N_6326);
xnor U9321 (N_9321,N_5249,N_5545);
or U9322 (N_9322,N_5395,N_5477);
nand U9323 (N_9323,N_6331,N_6497);
and U9324 (N_9324,N_6984,N_7217);
nor U9325 (N_9325,N_7404,N_5754);
nand U9326 (N_9326,N_7013,N_5118);
nand U9327 (N_9327,N_6922,N_5358);
nand U9328 (N_9328,N_6957,N_6144);
nand U9329 (N_9329,N_7237,N_7106);
or U9330 (N_9330,N_5406,N_5094);
xor U9331 (N_9331,N_6834,N_5051);
nor U9332 (N_9332,N_6529,N_5453);
xor U9333 (N_9333,N_7495,N_5783);
nand U9334 (N_9334,N_7186,N_6626);
or U9335 (N_9335,N_5430,N_7316);
nand U9336 (N_9336,N_5828,N_5033);
nor U9337 (N_9337,N_5011,N_5061);
and U9338 (N_9338,N_6294,N_6084);
and U9339 (N_9339,N_5202,N_5824);
xnor U9340 (N_9340,N_5860,N_6057);
or U9341 (N_9341,N_6302,N_5751);
or U9342 (N_9342,N_6102,N_7497);
and U9343 (N_9343,N_6444,N_6709);
nand U9344 (N_9344,N_5584,N_5305);
and U9345 (N_9345,N_6971,N_6716);
nand U9346 (N_9346,N_7207,N_5011);
xor U9347 (N_9347,N_5523,N_5861);
and U9348 (N_9348,N_6968,N_7431);
xor U9349 (N_9349,N_6480,N_5428);
nor U9350 (N_9350,N_6746,N_5915);
nand U9351 (N_9351,N_5445,N_6647);
or U9352 (N_9352,N_5812,N_5556);
and U9353 (N_9353,N_7414,N_7089);
nand U9354 (N_9354,N_7054,N_6369);
or U9355 (N_9355,N_5695,N_6030);
and U9356 (N_9356,N_5933,N_7133);
xor U9357 (N_9357,N_6437,N_5453);
nand U9358 (N_9358,N_5129,N_6295);
xor U9359 (N_9359,N_7396,N_6971);
or U9360 (N_9360,N_5762,N_6467);
xor U9361 (N_9361,N_7179,N_5328);
or U9362 (N_9362,N_6561,N_5431);
or U9363 (N_9363,N_5110,N_5245);
xor U9364 (N_9364,N_7366,N_6064);
or U9365 (N_9365,N_7102,N_5114);
xnor U9366 (N_9366,N_6595,N_5476);
and U9367 (N_9367,N_7483,N_6913);
nand U9368 (N_9368,N_6832,N_6372);
xor U9369 (N_9369,N_7171,N_5811);
nor U9370 (N_9370,N_5888,N_5221);
nand U9371 (N_9371,N_6839,N_7355);
xnor U9372 (N_9372,N_7489,N_6948);
nor U9373 (N_9373,N_5110,N_5437);
and U9374 (N_9374,N_5103,N_6007);
and U9375 (N_9375,N_6813,N_5131);
nor U9376 (N_9376,N_5425,N_5211);
nor U9377 (N_9377,N_5831,N_6136);
xor U9378 (N_9378,N_6694,N_5163);
nand U9379 (N_9379,N_6881,N_6724);
xnor U9380 (N_9380,N_6668,N_7343);
xnor U9381 (N_9381,N_5530,N_5778);
and U9382 (N_9382,N_6510,N_5370);
nand U9383 (N_9383,N_6007,N_7348);
and U9384 (N_9384,N_7190,N_5680);
or U9385 (N_9385,N_7211,N_5027);
nor U9386 (N_9386,N_5371,N_6593);
nor U9387 (N_9387,N_6242,N_5487);
or U9388 (N_9388,N_7319,N_5875);
xnor U9389 (N_9389,N_6557,N_5267);
or U9390 (N_9390,N_6467,N_7217);
or U9391 (N_9391,N_5348,N_5475);
or U9392 (N_9392,N_7440,N_5314);
and U9393 (N_9393,N_7266,N_5639);
and U9394 (N_9394,N_5579,N_5235);
xor U9395 (N_9395,N_5224,N_6882);
and U9396 (N_9396,N_5404,N_6842);
or U9397 (N_9397,N_6613,N_6267);
nor U9398 (N_9398,N_7255,N_6765);
xnor U9399 (N_9399,N_5480,N_5308);
nand U9400 (N_9400,N_6407,N_6299);
and U9401 (N_9401,N_7401,N_5178);
nand U9402 (N_9402,N_5776,N_5708);
or U9403 (N_9403,N_6475,N_5330);
nand U9404 (N_9404,N_5339,N_5752);
nor U9405 (N_9405,N_5536,N_5321);
nor U9406 (N_9406,N_5407,N_5903);
and U9407 (N_9407,N_5025,N_5752);
nor U9408 (N_9408,N_5165,N_7321);
nand U9409 (N_9409,N_6926,N_7478);
and U9410 (N_9410,N_6005,N_5698);
nor U9411 (N_9411,N_6469,N_5583);
nand U9412 (N_9412,N_6692,N_5755);
or U9413 (N_9413,N_5330,N_6884);
and U9414 (N_9414,N_5809,N_5556);
nand U9415 (N_9415,N_6103,N_5017);
nand U9416 (N_9416,N_6767,N_6628);
xnor U9417 (N_9417,N_7087,N_5475);
xnor U9418 (N_9418,N_5915,N_6687);
and U9419 (N_9419,N_5566,N_7045);
xnor U9420 (N_9420,N_5043,N_6687);
and U9421 (N_9421,N_6986,N_6444);
nor U9422 (N_9422,N_6139,N_5953);
xor U9423 (N_9423,N_5711,N_5591);
or U9424 (N_9424,N_7152,N_5526);
nand U9425 (N_9425,N_7222,N_6297);
or U9426 (N_9426,N_7047,N_5916);
nand U9427 (N_9427,N_6876,N_6607);
xor U9428 (N_9428,N_7308,N_5947);
or U9429 (N_9429,N_5149,N_6430);
nand U9430 (N_9430,N_5169,N_5556);
xnor U9431 (N_9431,N_6657,N_5961);
nor U9432 (N_9432,N_6316,N_7492);
and U9433 (N_9433,N_6333,N_6474);
and U9434 (N_9434,N_7448,N_7344);
nor U9435 (N_9435,N_6858,N_6255);
xor U9436 (N_9436,N_6146,N_7221);
and U9437 (N_9437,N_6009,N_5523);
and U9438 (N_9438,N_5436,N_6902);
and U9439 (N_9439,N_6565,N_5341);
xor U9440 (N_9440,N_6643,N_6052);
and U9441 (N_9441,N_6481,N_5397);
nor U9442 (N_9442,N_7200,N_5802);
xor U9443 (N_9443,N_7298,N_6367);
and U9444 (N_9444,N_7175,N_5004);
xnor U9445 (N_9445,N_5495,N_7076);
xnor U9446 (N_9446,N_5408,N_7060);
nand U9447 (N_9447,N_5375,N_6548);
nor U9448 (N_9448,N_6371,N_5802);
xor U9449 (N_9449,N_5417,N_5280);
nand U9450 (N_9450,N_5925,N_6438);
or U9451 (N_9451,N_5942,N_7275);
nor U9452 (N_9452,N_6041,N_5661);
nand U9453 (N_9453,N_6351,N_6493);
or U9454 (N_9454,N_5918,N_6238);
or U9455 (N_9455,N_5123,N_5837);
and U9456 (N_9456,N_5240,N_6525);
and U9457 (N_9457,N_5662,N_5270);
or U9458 (N_9458,N_5439,N_6854);
or U9459 (N_9459,N_5959,N_5954);
or U9460 (N_9460,N_6870,N_5584);
nand U9461 (N_9461,N_6763,N_5576);
or U9462 (N_9462,N_6061,N_5159);
and U9463 (N_9463,N_7051,N_7338);
or U9464 (N_9464,N_5726,N_7231);
nand U9465 (N_9465,N_6062,N_6807);
or U9466 (N_9466,N_6407,N_5110);
nor U9467 (N_9467,N_5283,N_6413);
or U9468 (N_9468,N_5271,N_5177);
and U9469 (N_9469,N_6615,N_7315);
or U9470 (N_9470,N_6114,N_5457);
nand U9471 (N_9471,N_5381,N_6251);
xnor U9472 (N_9472,N_6154,N_5051);
nor U9473 (N_9473,N_6311,N_5303);
or U9474 (N_9474,N_5611,N_6636);
and U9475 (N_9475,N_6099,N_6454);
xor U9476 (N_9476,N_6938,N_6540);
or U9477 (N_9477,N_6065,N_5402);
and U9478 (N_9478,N_7494,N_5624);
xor U9479 (N_9479,N_5347,N_6435);
and U9480 (N_9480,N_5329,N_6391);
xnor U9481 (N_9481,N_5787,N_6726);
nor U9482 (N_9482,N_5323,N_6845);
and U9483 (N_9483,N_7024,N_6657);
and U9484 (N_9484,N_5210,N_5485);
and U9485 (N_9485,N_6216,N_7228);
and U9486 (N_9486,N_6913,N_5501);
nor U9487 (N_9487,N_5860,N_5473);
xnor U9488 (N_9488,N_6913,N_7100);
nand U9489 (N_9489,N_7457,N_7021);
or U9490 (N_9490,N_5023,N_6866);
and U9491 (N_9491,N_5575,N_5751);
or U9492 (N_9492,N_6180,N_5835);
xor U9493 (N_9493,N_5962,N_6890);
xnor U9494 (N_9494,N_5587,N_6072);
and U9495 (N_9495,N_6154,N_6056);
or U9496 (N_9496,N_5285,N_6066);
xnor U9497 (N_9497,N_7109,N_6541);
nor U9498 (N_9498,N_6309,N_7105);
or U9499 (N_9499,N_7080,N_6390);
or U9500 (N_9500,N_7201,N_5480);
nand U9501 (N_9501,N_5549,N_6053);
xor U9502 (N_9502,N_6869,N_5703);
nand U9503 (N_9503,N_6318,N_6024);
nor U9504 (N_9504,N_6906,N_5459);
and U9505 (N_9505,N_6681,N_5777);
nand U9506 (N_9506,N_5152,N_5109);
nand U9507 (N_9507,N_6467,N_6463);
nor U9508 (N_9508,N_5973,N_5625);
or U9509 (N_9509,N_5694,N_7495);
nor U9510 (N_9510,N_6985,N_6857);
and U9511 (N_9511,N_6901,N_7053);
xor U9512 (N_9512,N_6733,N_5405);
and U9513 (N_9513,N_6760,N_6127);
nand U9514 (N_9514,N_6136,N_6134);
xnor U9515 (N_9515,N_5291,N_7319);
or U9516 (N_9516,N_7112,N_6356);
and U9517 (N_9517,N_7164,N_5109);
or U9518 (N_9518,N_7318,N_7045);
xnor U9519 (N_9519,N_5801,N_5552);
xnor U9520 (N_9520,N_6330,N_5068);
nor U9521 (N_9521,N_7438,N_6960);
and U9522 (N_9522,N_6863,N_5762);
or U9523 (N_9523,N_6244,N_7279);
xor U9524 (N_9524,N_6160,N_6967);
nor U9525 (N_9525,N_5660,N_5307);
or U9526 (N_9526,N_5927,N_5045);
or U9527 (N_9527,N_5916,N_6521);
and U9528 (N_9528,N_7181,N_6385);
nand U9529 (N_9529,N_7123,N_6367);
and U9530 (N_9530,N_5398,N_7053);
nor U9531 (N_9531,N_5964,N_6561);
or U9532 (N_9532,N_6560,N_6000);
or U9533 (N_9533,N_6242,N_6059);
nor U9534 (N_9534,N_5006,N_7199);
and U9535 (N_9535,N_5068,N_6282);
nor U9536 (N_9536,N_6067,N_5128);
nand U9537 (N_9537,N_5016,N_5135);
xor U9538 (N_9538,N_6727,N_6122);
nor U9539 (N_9539,N_5655,N_7478);
and U9540 (N_9540,N_6520,N_6759);
and U9541 (N_9541,N_5168,N_5743);
xor U9542 (N_9542,N_6244,N_5082);
or U9543 (N_9543,N_6191,N_5164);
nand U9544 (N_9544,N_5169,N_7091);
xnor U9545 (N_9545,N_5969,N_6204);
nand U9546 (N_9546,N_6023,N_5180);
nand U9547 (N_9547,N_5836,N_6288);
or U9548 (N_9548,N_6689,N_6204);
nand U9549 (N_9549,N_7117,N_7147);
nor U9550 (N_9550,N_5179,N_5304);
xnor U9551 (N_9551,N_7440,N_5144);
and U9552 (N_9552,N_6476,N_5697);
xor U9553 (N_9553,N_6583,N_6945);
nor U9554 (N_9554,N_5988,N_5351);
xnor U9555 (N_9555,N_5244,N_5170);
nor U9556 (N_9556,N_5619,N_5268);
nor U9557 (N_9557,N_6766,N_5306);
and U9558 (N_9558,N_7240,N_6467);
nor U9559 (N_9559,N_5772,N_6905);
xnor U9560 (N_9560,N_5069,N_7330);
xnor U9561 (N_9561,N_6717,N_5744);
xor U9562 (N_9562,N_6329,N_7266);
and U9563 (N_9563,N_6376,N_6249);
xnor U9564 (N_9564,N_6103,N_6680);
nand U9565 (N_9565,N_5069,N_7035);
nand U9566 (N_9566,N_6185,N_7047);
and U9567 (N_9567,N_5424,N_5695);
or U9568 (N_9568,N_6144,N_6537);
nor U9569 (N_9569,N_6650,N_6283);
nor U9570 (N_9570,N_5469,N_7300);
nor U9571 (N_9571,N_6536,N_7075);
xor U9572 (N_9572,N_5083,N_6404);
or U9573 (N_9573,N_7172,N_5180);
or U9574 (N_9574,N_5789,N_7303);
nor U9575 (N_9575,N_6766,N_7274);
and U9576 (N_9576,N_7198,N_6546);
xor U9577 (N_9577,N_5740,N_5218);
nand U9578 (N_9578,N_7096,N_6852);
and U9579 (N_9579,N_6363,N_6114);
nand U9580 (N_9580,N_7147,N_6546);
nor U9581 (N_9581,N_5724,N_6202);
nand U9582 (N_9582,N_6547,N_7213);
nor U9583 (N_9583,N_6446,N_7379);
and U9584 (N_9584,N_6479,N_7258);
nor U9585 (N_9585,N_7012,N_6967);
and U9586 (N_9586,N_5773,N_7463);
xor U9587 (N_9587,N_5196,N_5446);
or U9588 (N_9588,N_7377,N_6927);
or U9589 (N_9589,N_6094,N_6447);
and U9590 (N_9590,N_5243,N_7305);
and U9591 (N_9591,N_6764,N_5598);
or U9592 (N_9592,N_6073,N_6414);
nand U9593 (N_9593,N_7276,N_5778);
or U9594 (N_9594,N_5049,N_5453);
and U9595 (N_9595,N_5362,N_7415);
or U9596 (N_9596,N_5315,N_7242);
nor U9597 (N_9597,N_6517,N_6389);
or U9598 (N_9598,N_6723,N_5446);
and U9599 (N_9599,N_5159,N_7329);
nand U9600 (N_9600,N_6865,N_7052);
and U9601 (N_9601,N_5806,N_5716);
nor U9602 (N_9602,N_5698,N_6887);
xnor U9603 (N_9603,N_7378,N_5003);
xor U9604 (N_9604,N_5962,N_5734);
xor U9605 (N_9605,N_6893,N_6527);
xnor U9606 (N_9606,N_5040,N_7258);
nand U9607 (N_9607,N_6097,N_5005);
xor U9608 (N_9608,N_7025,N_6715);
nor U9609 (N_9609,N_6945,N_5465);
nor U9610 (N_9610,N_5205,N_5469);
or U9611 (N_9611,N_6160,N_5412);
nor U9612 (N_9612,N_5258,N_6399);
xnor U9613 (N_9613,N_6305,N_6200);
nand U9614 (N_9614,N_6831,N_6032);
nand U9615 (N_9615,N_6119,N_5550);
xor U9616 (N_9616,N_6292,N_5593);
and U9617 (N_9617,N_7197,N_5052);
nand U9618 (N_9618,N_7054,N_5092);
nor U9619 (N_9619,N_5030,N_6367);
nor U9620 (N_9620,N_5823,N_5143);
and U9621 (N_9621,N_5265,N_6927);
and U9622 (N_9622,N_7452,N_5273);
nand U9623 (N_9623,N_7300,N_5957);
nor U9624 (N_9624,N_5189,N_5144);
and U9625 (N_9625,N_7175,N_5180);
nand U9626 (N_9626,N_6059,N_6901);
or U9627 (N_9627,N_5351,N_5872);
or U9628 (N_9628,N_6292,N_5451);
nand U9629 (N_9629,N_5273,N_6696);
nand U9630 (N_9630,N_7331,N_5853);
or U9631 (N_9631,N_6527,N_5647);
and U9632 (N_9632,N_5151,N_5982);
or U9633 (N_9633,N_7342,N_5835);
nand U9634 (N_9634,N_7410,N_5597);
and U9635 (N_9635,N_6007,N_6346);
nand U9636 (N_9636,N_5546,N_6344);
or U9637 (N_9637,N_5530,N_6303);
nor U9638 (N_9638,N_7465,N_6970);
nand U9639 (N_9639,N_5078,N_6370);
xnor U9640 (N_9640,N_7186,N_7328);
xnor U9641 (N_9641,N_6252,N_7374);
or U9642 (N_9642,N_5269,N_7335);
nand U9643 (N_9643,N_6661,N_6111);
nor U9644 (N_9644,N_5879,N_7115);
xnor U9645 (N_9645,N_7452,N_6454);
and U9646 (N_9646,N_7366,N_6512);
or U9647 (N_9647,N_6395,N_6800);
nor U9648 (N_9648,N_6177,N_5550);
nand U9649 (N_9649,N_6463,N_5312);
nand U9650 (N_9650,N_6499,N_6075);
or U9651 (N_9651,N_7116,N_7205);
xnor U9652 (N_9652,N_5829,N_5670);
nor U9653 (N_9653,N_5713,N_5446);
and U9654 (N_9654,N_6041,N_6329);
or U9655 (N_9655,N_7405,N_6156);
or U9656 (N_9656,N_5244,N_5229);
and U9657 (N_9657,N_5366,N_6170);
xnor U9658 (N_9658,N_5724,N_5745);
nand U9659 (N_9659,N_7393,N_6973);
or U9660 (N_9660,N_5702,N_7068);
and U9661 (N_9661,N_5527,N_6936);
xor U9662 (N_9662,N_6561,N_5057);
xor U9663 (N_9663,N_5010,N_5095);
nor U9664 (N_9664,N_5827,N_6499);
nor U9665 (N_9665,N_5667,N_5149);
and U9666 (N_9666,N_5356,N_5052);
nand U9667 (N_9667,N_5328,N_6118);
and U9668 (N_9668,N_6530,N_6073);
xor U9669 (N_9669,N_7090,N_6054);
nand U9670 (N_9670,N_5081,N_6542);
nor U9671 (N_9671,N_7007,N_6757);
or U9672 (N_9672,N_7463,N_6048);
or U9673 (N_9673,N_5266,N_6299);
nor U9674 (N_9674,N_5213,N_5722);
xnor U9675 (N_9675,N_5690,N_5047);
nand U9676 (N_9676,N_7265,N_5041);
nand U9677 (N_9677,N_6570,N_6336);
nor U9678 (N_9678,N_5367,N_7285);
xnor U9679 (N_9679,N_7149,N_6956);
nand U9680 (N_9680,N_6969,N_5342);
xnor U9681 (N_9681,N_6505,N_7371);
or U9682 (N_9682,N_6108,N_5351);
xor U9683 (N_9683,N_6844,N_5236);
and U9684 (N_9684,N_6156,N_6456);
nand U9685 (N_9685,N_6420,N_5564);
or U9686 (N_9686,N_6503,N_6245);
and U9687 (N_9687,N_5834,N_6921);
and U9688 (N_9688,N_7089,N_6319);
nor U9689 (N_9689,N_6917,N_7235);
or U9690 (N_9690,N_6090,N_5395);
nor U9691 (N_9691,N_5891,N_5986);
xnor U9692 (N_9692,N_7453,N_5745);
xor U9693 (N_9693,N_5418,N_7179);
nor U9694 (N_9694,N_5810,N_7149);
or U9695 (N_9695,N_6526,N_5113);
or U9696 (N_9696,N_6979,N_5319);
xor U9697 (N_9697,N_5519,N_6825);
or U9698 (N_9698,N_6529,N_5310);
nor U9699 (N_9699,N_6327,N_6813);
nor U9700 (N_9700,N_6176,N_6346);
or U9701 (N_9701,N_6461,N_6588);
nor U9702 (N_9702,N_6355,N_5565);
nor U9703 (N_9703,N_6017,N_5553);
xnor U9704 (N_9704,N_6850,N_6531);
or U9705 (N_9705,N_5526,N_5726);
nor U9706 (N_9706,N_6694,N_6527);
or U9707 (N_9707,N_7111,N_6662);
nand U9708 (N_9708,N_6096,N_6443);
xnor U9709 (N_9709,N_5877,N_6613);
nor U9710 (N_9710,N_6772,N_6466);
nor U9711 (N_9711,N_5051,N_7071);
xnor U9712 (N_9712,N_7404,N_5552);
nand U9713 (N_9713,N_7311,N_7089);
nor U9714 (N_9714,N_7242,N_6822);
and U9715 (N_9715,N_6935,N_7249);
nor U9716 (N_9716,N_5373,N_5652);
nand U9717 (N_9717,N_7302,N_6520);
nor U9718 (N_9718,N_6990,N_7387);
or U9719 (N_9719,N_5170,N_5878);
xor U9720 (N_9720,N_5235,N_6486);
or U9721 (N_9721,N_5655,N_6621);
xnor U9722 (N_9722,N_7400,N_7357);
nand U9723 (N_9723,N_5299,N_5393);
nor U9724 (N_9724,N_5691,N_6308);
nand U9725 (N_9725,N_5018,N_5508);
or U9726 (N_9726,N_6311,N_5076);
xnor U9727 (N_9727,N_6685,N_6211);
nor U9728 (N_9728,N_5941,N_7108);
nand U9729 (N_9729,N_5816,N_6430);
nand U9730 (N_9730,N_5662,N_7378);
xor U9731 (N_9731,N_7461,N_7197);
nor U9732 (N_9732,N_6750,N_7379);
xnor U9733 (N_9733,N_5922,N_5211);
nand U9734 (N_9734,N_6797,N_5742);
nand U9735 (N_9735,N_7216,N_6247);
nor U9736 (N_9736,N_6770,N_5686);
and U9737 (N_9737,N_6892,N_5013);
nor U9738 (N_9738,N_5358,N_5620);
and U9739 (N_9739,N_5323,N_6079);
xnor U9740 (N_9740,N_6455,N_6856);
nor U9741 (N_9741,N_5278,N_5093);
nor U9742 (N_9742,N_5520,N_6413);
nand U9743 (N_9743,N_5697,N_5403);
nor U9744 (N_9744,N_6172,N_6298);
and U9745 (N_9745,N_6679,N_7212);
nor U9746 (N_9746,N_6044,N_7412);
and U9747 (N_9747,N_5261,N_5097);
or U9748 (N_9748,N_6619,N_5159);
and U9749 (N_9749,N_7442,N_6962);
nor U9750 (N_9750,N_5423,N_5214);
nand U9751 (N_9751,N_6486,N_6860);
or U9752 (N_9752,N_5183,N_5825);
nand U9753 (N_9753,N_5374,N_6094);
nor U9754 (N_9754,N_6152,N_7159);
and U9755 (N_9755,N_6703,N_6361);
nand U9756 (N_9756,N_5635,N_5328);
nor U9757 (N_9757,N_5165,N_6707);
nor U9758 (N_9758,N_7041,N_5326);
nor U9759 (N_9759,N_5426,N_6949);
and U9760 (N_9760,N_6530,N_5350);
or U9761 (N_9761,N_6759,N_7219);
nor U9762 (N_9762,N_6641,N_6403);
nor U9763 (N_9763,N_5353,N_7155);
nand U9764 (N_9764,N_5770,N_5272);
xnor U9765 (N_9765,N_7325,N_6857);
and U9766 (N_9766,N_7316,N_6241);
nor U9767 (N_9767,N_6290,N_6254);
and U9768 (N_9768,N_5415,N_6718);
nor U9769 (N_9769,N_7084,N_5505);
nand U9770 (N_9770,N_6623,N_5413);
nand U9771 (N_9771,N_5748,N_5912);
xnor U9772 (N_9772,N_6600,N_6015);
xor U9773 (N_9773,N_5151,N_6548);
or U9774 (N_9774,N_6469,N_7360);
xnor U9775 (N_9775,N_5288,N_5268);
nand U9776 (N_9776,N_6641,N_5771);
and U9777 (N_9777,N_5230,N_5466);
nand U9778 (N_9778,N_6947,N_6757);
and U9779 (N_9779,N_5766,N_7182);
xnor U9780 (N_9780,N_5122,N_6787);
xor U9781 (N_9781,N_6804,N_5739);
nor U9782 (N_9782,N_5623,N_5735);
xor U9783 (N_9783,N_5115,N_7229);
nand U9784 (N_9784,N_6180,N_6834);
xor U9785 (N_9785,N_5176,N_7195);
nor U9786 (N_9786,N_6785,N_7323);
and U9787 (N_9787,N_7067,N_5101);
or U9788 (N_9788,N_5274,N_5023);
and U9789 (N_9789,N_7002,N_6045);
xnor U9790 (N_9790,N_7269,N_7326);
nand U9791 (N_9791,N_6105,N_5841);
xnor U9792 (N_9792,N_7114,N_6039);
and U9793 (N_9793,N_6555,N_6667);
and U9794 (N_9794,N_7110,N_6212);
and U9795 (N_9795,N_6227,N_6199);
nand U9796 (N_9796,N_6187,N_5490);
nand U9797 (N_9797,N_6390,N_6448);
nand U9798 (N_9798,N_5808,N_7166);
nand U9799 (N_9799,N_7130,N_7367);
nor U9800 (N_9800,N_5200,N_5610);
or U9801 (N_9801,N_7415,N_5644);
and U9802 (N_9802,N_6467,N_6802);
xor U9803 (N_9803,N_6784,N_5413);
nand U9804 (N_9804,N_6318,N_6924);
nor U9805 (N_9805,N_6538,N_6393);
and U9806 (N_9806,N_5731,N_5113);
xnor U9807 (N_9807,N_5792,N_5871);
or U9808 (N_9808,N_5925,N_7058);
and U9809 (N_9809,N_6604,N_7133);
nor U9810 (N_9810,N_6574,N_5642);
and U9811 (N_9811,N_5428,N_6407);
and U9812 (N_9812,N_5022,N_5262);
xor U9813 (N_9813,N_7193,N_6136);
nor U9814 (N_9814,N_5021,N_6885);
nor U9815 (N_9815,N_5230,N_5484);
nand U9816 (N_9816,N_5948,N_5739);
nor U9817 (N_9817,N_7312,N_5151);
and U9818 (N_9818,N_6500,N_7380);
or U9819 (N_9819,N_5088,N_5883);
nand U9820 (N_9820,N_5813,N_7185);
xor U9821 (N_9821,N_7210,N_5581);
nand U9822 (N_9822,N_5729,N_5743);
nand U9823 (N_9823,N_5508,N_5823);
xor U9824 (N_9824,N_6646,N_5423);
and U9825 (N_9825,N_5759,N_7311);
or U9826 (N_9826,N_5192,N_7211);
and U9827 (N_9827,N_6889,N_5362);
and U9828 (N_9828,N_6768,N_7090);
nand U9829 (N_9829,N_7002,N_5896);
and U9830 (N_9830,N_6980,N_6478);
xor U9831 (N_9831,N_6492,N_6342);
or U9832 (N_9832,N_5995,N_6084);
nor U9833 (N_9833,N_5162,N_6499);
or U9834 (N_9834,N_6244,N_7294);
and U9835 (N_9835,N_5330,N_5100);
nand U9836 (N_9836,N_7070,N_6675);
nand U9837 (N_9837,N_7072,N_5154);
and U9838 (N_9838,N_5231,N_7464);
xnor U9839 (N_9839,N_5361,N_5391);
nor U9840 (N_9840,N_6291,N_7160);
and U9841 (N_9841,N_7076,N_7007);
nor U9842 (N_9842,N_5594,N_7231);
nor U9843 (N_9843,N_5962,N_5105);
xnor U9844 (N_9844,N_6085,N_6835);
nor U9845 (N_9845,N_5263,N_7218);
nand U9846 (N_9846,N_5254,N_7121);
xnor U9847 (N_9847,N_5779,N_7072);
or U9848 (N_9848,N_7433,N_6529);
and U9849 (N_9849,N_7209,N_5404);
xor U9850 (N_9850,N_5031,N_7112);
nand U9851 (N_9851,N_6484,N_7398);
nand U9852 (N_9852,N_5102,N_7431);
or U9853 (N_9853,N_6705,N_5313);
and U9854 (N_9854,N_6402,N_5277);
or U9855 (N_9855,N_6759,N_7471);
xor U9856 (N_9856,N_5349,N_7413);
and U9857 (N_9857,N_5066,N_6175);
nor U9858 (N_9858,N_6540,N_6992);
nor U9859 (N_9859,N_5407,N_7167);
xnor U9860 (N_9860,N_5004,N_5181);
and U9861 (N_9861,N_7491,N_5979);
nand U9862 (N_9862,N_6506,N_6791);
and U9863 (N_9863,N_6736,N_6651);
or U9864 (N_9864,N_5476,N_5173);
nand U9865 (N_9865,N_7191,N_7357);
nor U9866 (N_9866,N_5931,N_6178);
nand U9867 (N_9867,N_5104,N_5335);
nor U9868 (N_9868,N_6760,N_5300);
nor U9869 (N_9869,N_6770,N_6229);
nor U9870 (N_9870,N_6925,N_6732);
and U9871 (N_9871,N_7032,N_5112);
xnor U9872 (N_9872,N_6378,N_6340);
or U9873 (N_9873,N_5658,N_6866);
nand U9874 (N_9874,N_7198,N_7494);
nor U9875 (N_9875,N_5494,N_5625);
nand U9876 (N_9876,N_5076,N_5580);
nor U9877 (N_9877,N_5656,N_7447);
nand U9878 (N_9878,N_5837,N_6802);
and U9879 (N_9879,N_6393,N_7154);
or U9880 (N_9880,N_6208,N_6760);
xnor U9881 (N_9881,N_5673,N_5022);
nand U9882 (N_9882,N_6177,N_6671);
and U9883 (N_9883,N_5148,N_7435);
or U9884 (N_9884,N_7485,N_7490);
xnor U9885 (N_9885,N_5390,N_6402);
or U9886 (N_9886,N_5815,N_7083);
and U9887 (N_9887,N_6305,N_7329);
nor U9888 (N_9888,N_5396,N_5491);
nor U9889 (N_9889,N_5163,N_5388);
or U9890 (N_9890,N_7207,N_5060);
or U9891 (N_9891,N_6158,N_7285);
and U9892 (N_9892,N_6715,N_6228);
xor U9893 (N_9893,N_5743,N_6821);
nor U9894 (N_9894,N_7340,N_5714);
xnor U9895 (N_9895,N_6346,N_7384);
or U9896 (N_9896,N_6483,N_5924);
and U9897 (N_9897,N_6128,N_6917);
xnor U9898 (N_9898,N_6708,N_6356);
nor U9899 (N_9899,N_6040,N_7102);
or U9900 (N_9900,N_6226,N_7443);
or U9901 (N_9901,N_6987,N_6602);
nor U9902 (N_9902,N_6662,N_7229);
or U9903 (N_9903,N_5239,N_7228);
or U9904 (N_9904,N_7036,N_5988);
or U9905 (N_9905,N_5716,N_7179);
xnor U9906 (N_9906,N_5780,N_7256);
and U9907 (N_9907,N_6186,N_5175);
xnor U9908 (N_9908,N_6648,N_5887);
nor U9909 (N_9909,N_7472,N_5887);
or U9910 (N_9910,N_6097,N_5639);
xnor U9911 (N_9911,N_7076,N_6487);
and U9912 (N_9912,N_6397,N_5123);
nor U9913 (N_9913,N_7245,N_6891);
xnor U9914 (N_9914,N_6890,N_6731);
or U9915 (N_9915,N_6058,N_7205);
or U9916 (N_9916,N_5885,N_5729);
and U9917 (N_9917,N_5849,N_5089);
nand U9918 (N_9918,N_5905,N_6512);
nand U9919 (N_9919,N_6873,N_5975);
nand U9920 (N_9920,N_5795,N_6131);
nor U9921 (N_9921,N_6258,N_6437);
nand U9922 (N_9922,N_6439,N_7434);
xnor U9923 (N_9923,N_6905,N_6000);
nand U9924 (N_9924,N_6591,N_5660);
xor U9925 (N_9925,N_6561,N_6012);
and U9926 (N_9926,N_7300,N_6053);
nand U9927 (N_9927,N_5224,N_6418);
nor U9928 (N_9928,N_7487,N_6417);
nor U9929 (N_9929,N_6360,N_7043);
and U9930 (N_9930,N_7265,N_6104);
nand U9931 (N_9931,N_5625,N_6137);
nand U9932 (N_9932,N_7412,N_6449);
or U9933 (N_9933,N_6646,N_6610);
or U9934 (N_9934,N_7197,N_7321);
and U9935 (N_9935,N_7309,N_5675);
nand U9936 (N_9936,N_6783,N_6301);
nand U9937 (N_9937,N_6799,N_6702);
xor U9938 (N_9938,N_7498,N_6316);
nor U9939 (N_9939,N_6310,N_5338);
and U9940 (N_9940,N_6910,N_7399);
xor U9941 (N_9941,N_6251,N_6796);
or U9942 (N_9942,N_7316,N_6932);
xor U9943 (N_9943,N_5935,N_5983);
and U9944 (N_9944,N_6497,N_6181);
nand U9945 (N_9945,N_5376,N_6930);
nand U9946 (N_9946,N_7275,N_7448);
nand U9947 (N_9947,N_6861,N_6332);
xnor U9948 (N_9948,N_6469,N_6572);
nor U9949 (N_9949,N_5289,N_5901);
xor U9950 (N_9950,N_5453,N_5820);
nor U9951 (N_9951,N_5764,N_7314);
or U9952 (N_9952,N_6485,N_6799);
nand U9953 (N_9953,N_5516,N_7067);
and U9954 (N_9954,N_6111,N_6560);
nor U9955 (N_9955,N_6146,N_6417);
and U9956 (N_9956,N_5930,N_5788);
and U9957 (N_9957,N_6703,N_5045);
or U9958 (N_9958,N_5572,N_5640);
nand U9959 (N_9959,N_7382,N_5851);
and U9960 (N_9960,N_6173,N_7315);
xnor U9961 (N_9961,N_7265,N_5839);
xnor U9962 (N_9962,N_5677,N_6031);
nand U9963 (N_9963,N_6226,N_7455);
nor U9964 (N_9964,N_7499,N_7229);
or U9965 (N_9965,N_6537,N_7147);
nor U9966 (N_9966,N_6097,N_5730);
xor U9967 (N_9967,N_7372,N_5575);
xor U9968 (N_9968,N_5396,N_5074);
xor U9969 (N_9969,N_6864,N_5229);
and U9970 (N_9970,N_6647,N_5357);
or U9971 (N_9971,N_5771,N_5694);
or U9972 (N_9972,N_5309,N_5331);
nor U9973 (N_9973,N_5468,N_7298);
nor U9974 (N_9974,N_6123,N_6750);
or U9975 (N_9975,N_5100,N_5291);
and U9976 (N_9976,N_6285,N_7478);
or U9977 (N_9977,N_7295,N_6516);
nor U9978 (N_9978,N_6276,N_6002);
or U9979 (N_9979,N_7052,N_6286);
or U9980 (N_9980,N_5323,N_5442);
nand U9981 (N_9981,N_5349,N_6852);
nand U9982 (N_9982,N_6450,N_5200);
nor U9983 (N_9983,N_7151,N_5535);
and U9984 (N_9984,N_7111,N_7053);
and U9985 (N_9985,N_5226,N_5663);
xor U9986 (N_9986,N_6785,N_5995);
nand U9987 (N_9987,N_5349,N_5167);
nand U9988 (N_9988,N_5707,N_7399);
xnor U9989 (N_9989,N_6076,N_5717);
or U9990 (N_9990,N_6221,N_5067);
or U9991 (N_9991,N_5217,N_5927);
or U9992 (N_9992,N_5957,N_6676);
nand U9993 (N_9993,N_7446,N_7120);
or U9994 (N_9994,N_7232,N_7053);
nand U9995 (N_9995,N_6008,N_7064);
nor U9996 (N_9996,N_5740,N_7053);
xnor U9997 (N_9997,N_6789,N_5284);
xnor U9998 (N_9998,N_5453,N_5067);
and U9999 (N_9999,N_7292,N_5331);
xor U10000 (N_10000,N_8617,N_7834);
and U10001 (N_10001,N_9606,N_9691);
nor U10002 (N_10002,N_9459,N_8292);
and U10003 (N_10003,N_9794,N_9620);
nand U10004 (N_10004,N_8507,N_7808);
or U10005 (N_10005,N_8179,N_8470);
nor U10006 (N_10006,N_8294,N_9415);
and U10007 (N_10007,N_7591,N_8106);
nor U10008 (N_10008,N_8895,N_9372);
nand U10009 (N_10009,N_8672,N_9856);
nand U10010 (N_10010,N_8373,N_8473);
or U10011 (N_10011,N_8398,N_8392);
or U10012 (N_10012,N_9171,N_9199);
and U10013 (N_10013,N_7904,N_8939);
nand U10014 (N_10014,N_7606,N_8879);
and U10015 (N_10015,N_9401,N_8213);
or U10016 (N_10016,N_8546,N_9407);
and U10017 (N_10017,N_8386,N_7599);
and U10018 (N_10018,N_7940,N_7567);
nor U10019 (N_10019,N_9833,N_9524);
and U10020 (N_10020,N_8836,N_8323);
xnor U10021 (N_10021,N_8839,N_7915);
or U10022 (N_10022,N_8030,N_8985);
nor U10023 (N_10023,N_9374,N_8361);
xnor U10024 (N_10024,N_8013,N_9671);
and U10025 (N_10025,N_7559,N_9702);
nand U10026 (N_10026,N_8930,N_9067);
and U10027 (N_10027,N_7903,N_9250);
xnor U10028 (N_10028,N_9118,N_7548);
nor U10029 (N_10029,N_9168,N_9533);
nand U10030 (N_10030,N_7635,N_9701);
or U10031 (N_10031,N_9455,N_9882);
or U10032 (N_10032,N_8845,N_7821);
xnor U10033 (N_10033,N_9737,N_9529);
nor U10034 (N_10034,N_8891,N_9842);
nor U10035 (N_10035,N_9886,N_8431);
xor U10036 (N_10036,N_8677,N_8664);
nor U10037 (N_10037,N_8814,N_7889);
nor U10038 (N_10038,N_9971,N_9380);
and U10039 (N_10039,N_8926,N_9367);
nor U10040 (N_10040,N_8936,N_9958);
and U10041 (N_10041,N_8194,N_9177);
and U10042 (N_10042,N_8422,N_8667);
xor U10043 (N_10043,N_9190,N_8940);
nand U10044 (N_10044,N_9685,N_9617);
xor U10045 (N_10045,N_9313,N_8548);
xor U10046 (N_10046,N_8807,N_8728);
or U10047 (N_10047,N_9488,N_8056);
xor U10048 (N_10048,N_8004,N_9229);
and U10049 (N_10049,N_8295,N_8559);
or U10050 (N_10050,N_8161,N_9649);
nor U10051 (N_10051,N_8883,N_8584);
and U10052 (N_10052,N_9591,N_9608);
or U10053 (N_10053,N_9818,N_9065);
and U10054 (N_10054,N_9351,N_9744);
xor U10055 (N_10055,N_8107,N_8867);
nor U10056 (N_10056,N_9628,N_9343);
or U10057 (N_10057,N_8994,N_8627);
and U10058 (N_10058,N_9817,N_8254);
xor U10059 (N_10059,N_7870,N_8819);
nand U10060 (N_10060,N_8840,N_8597);
nor U10061 (N_10061,N_8674,N_8172);
or U10062 (N_10062,N_9275,N_8525);
nand U10063 (N_10063,N_7705,N_7984);
nand U10064 (N_10064,N_8729,N_7879);
nor U10065 (N_10065,N_8218,N_9866);
or U10066 (N_10066,N_9003,N_8259);
xnor U10067 (N_10067,N_8448,N_7780);
nand U10068 (N_10068,N_9472,N_9422);
or U10069 (N_10069,N_9449,N_8698);
nor U10070 (N_10070,N_8544,N_8184);
xnor U10071 (N_10071,N_9453,N_7899);
xnor U10072 (N_10072,N_7817,N_7779);
xnor U10073 (N_10073,N_9166,N_8281);
nand U10074 (N_10074,N_8964,N_8658);
xor U10075 (N_10075,N_7991,N_8562);
nor U10076 (N_10076,N_9396,N_7596);
nand U10077 (N_10077,N_8193,N_7977);
or U10078 (N_10078,N_8601,N_8374);
or U10079 (N_10079,N_9032,N_8523);
nor U10080 (N_10080,N_9498,N_8219);
and U10081 (N_10081,N_8810,N_8125);
and U10082 (N_10082,N_9743,N_9814);
nor U10083 (N_10083,N_8183,N_7850);
nor U10084 (N_10084,N_9518,N_8232);
xnor U10085 (N_10085,N_8874,N_9384);
nor U10086 (N_10086,N_9115,N_9854);
or U10087 (N_10087,N_9345,N_9651);
xor U10088 (N_10088,N_9815,N_9385);
and U10089 (N_10089,N_7981,N_7842);
or U10090 (N_10090,N_9318,N_9416);
nand U10091 (N_10091,N_8980,N_8445);
and U10092 (N_10092,N_9182,N_9820);
or U10093 (N_10093,N_9145,N_9360);
xnor U10094 (N_10094,N_9536,N_9424);
nand U10095 (N_10095,N_8931,N_8089);
and U10096 (N_10096,N_9219,N_9892);
nor U10097 (N_10097,N_9107,N_9297);
or U10098 (N_10098,N_8649,N_9478);
xor U10099 (N_10099,N_9515,N_8261);
or U10100 (N_10100,N_9873,N_9953);
xor U10101 (N_10101,N_8616,N_8847);
and U10102 (N_10102,N_8241,N_9633);
xnor U10103 (N_10103,N_9878,N_9226);
nand U10104 (N_10104,N_9995,N_7974);
nor U10105 (N_10105,N_9456,N_8607);
or U10106 (N_10106,N_8449,N_8778);
and U10107 (N_10107,N_8159,N_8384);
xor U10108 (N_10108,N_8045,N_8954);
or U10109 (N_10109,N_8355,N_8497);
nand U10110 (N_10110,N_7883,N_9317);
nand U10111 (N_10111,N_7593,N_9753);
nand U10112 (N_10112,N_7936,N_8304);
and U10113 (N_10113,N_7756,N_8419);
nor U10114 (N_10114,N_9266,N_9054);
or U10115 (N_10115,N_8668,N_9733);
or U10116 (N_10116,N_8971,N_9026);
or U10117 (N_10117,N_7960,N_8909);
nand U10118 (N_10118,N_8841,N_9872);
or U10119 (N_10119,N_9444,N_8828);
nand U10120 (N_10120,N_9011,N_8215);
xor U10121 (N_10121,N_9732,N_8972);
nand U10122 (N_10122,N_9601,N_7733);
nor U10123 (N_10123,N_8765,N_7822);
nor U10124 (N_10124,N_8220,N_9289);
and U10125 (N_10125,N_8624,N_7696);
nor U10126 (N_10126,N_8310,N_9029);
xnor U10127 (N_10127,N_8965,N_9073);
nand U10128 (N_10128,N_9272,N_7659);
and U10129 (N_10129,N_9208,N_7546);
and U10130 (N_10130,N_9548,N_8663);
and U10131 (N_10131,N_9673,N_8790);
nand U10132 (N_10132,N_7776,N_7755);
xnor U10133 (N_10133,N_7877,N_9001);
xor U10134 (N_10134,N_8103,N_8817);
xor U10135 (N_10135,N_8858,N_9043);
nand U10136 (N_10136,N_9954,N_9224);
and U10137 (N_10137,N_9722,N_8015);
and U10138 (N_10138,N_9710,N_9550);
xor U10139 (N_10139,N_7540,N_8735);
nor U10140 (N_10140,N_8691,N_8651);
nor U10141 (N_10141,N_9883,N_7841);
and U10142 (N_10142,N_8852,N_8461);
xnor U10143 (N_10143,N_9085,N_9075);
or U10144 (N_10144,N_7708,N_7661);
and U10145 (N_10145,N_8214,N_8745);
xnor U10146 (N_10146,N_9699,N_7771);
or U10147 (N_10147,N_9920,N_8039);
or U10148 (N_10148,N_7939,N_8586);
and U10149 (N_10149,N_8212,N_8471);
and U10150 (N_10150,N_9981,N_9486);
and U10151 (N_10151,N_7930,N_9526);
nand U10152 (N_10152,N_8750,N_8889);
xor U10153 (N_10153,N_9139,N_9725);
nand U10154 (N_10154,N_9062,N_8661);
nor U10155 (N_10155,N_8288,N_9688);
nor U10156 (N_10156,N_9364,N_9893);
xnor U10157 (N_10157,N_8365,N_8353);
nor U10158 (N_10158,N_9778,N_8849);
and U10159 (N_10159,N_8657,N_7713);
or U10160 (N_10160,N_7990,N_9235);
nand U10161 (N_10161,N_8088,N_9996);
or U10162 (N_10162,N_8427,N_8185);
nor U10163 (N_10163,N_8370,N_9090);
or U10164 (N_10164,N_7504,N_9175);
or U10165 (N_10165,N_8153,N_9331);
nor U10166 (N_10166,N_9354,N_7876);
and U10167 (N_10167,N_9353,N_8394);
and U10168 (N_10168,N_9220,N_9309);
and U10169 (N_10169,N_9863,N_9096);
nand U10170 (N_10170,N_7742,N_7524);
and U10171 (N_10171,N_8912,N_8770);
or U10172 (N_10172,N_8812,N_8527);
nor U10173 (N_10173,N_7740,N_9538);
xor U10174 (N_10174,N_9112,N_8513);
xnor U10175 (N_10175,N_9657,N_8169);
nand U10176 (N_10176,N_8751,N_8341);
and U10177 (N_10177,N_8446,N_9823);
nand U10178 (N_10178,N_7793,N_8113);
nand U10179 (N_10179,N_8011,N_7999);
or U10180 (N_10180,N_9582,N_7769);
xor U10181 (N_10181,N_9489,N_7773);
or U10182 (N_10182,N_8332,N_8065);
nand U10183 (N_10183,N_8522,N_9980);
and U10184 (N_10184,N_8614,N_7777);
xnor U10185 (N_10185,N_7586,N_8000);
and U10186 (N_10186,N_8280,N_8073);
and U10187 (N_10187,N_9805,N_9947);
and U10188 (N_10188,N_8942,N_9709);
nor U10189 (N_10189,N_8742,N_9781);
nand U10190 (N_10190,N_8483,N_9927);
nor U10191 (N_10191,N_7820,N_8626);
nor U10192 (N_10192,N_8076,N_9173);
xnor U10193 (N_10193,N_7588,N_8404);
and U10194 (N_10194,N_9638,N_9670);
or U10195 (N_10195,N_7537,N_9680);
and U10196 (N_10196,N_9358,N_8192);
or U10197 (N_10197,N_7997,N_8864);
or U10198 (N_10198,N_9894,N_7768);
xnor U10199 (N_10199,N_8884,N_8300);
nand U10200 (N_10200,N_8561,N_9776);
xnor U10201 (N_10201,N_9361,N_8162);
and U10202 (N_10202,N_8020,N_9986);
xnor U10203 (N_10203,N_9768,N_8547);
or U10204 (N_10204,N_9740,N_9267);
xnor U10205 (N_10205,N_9296,N_8347);
or U10206 (N_10206,N_9643,N_8919);
xnor U10207 (N_10207,N_8612,N_9060);
nand U10208 (N_10208,N_9473,N_8808);
nor U10209 (N_10209,N_8163,N_8393);
nand U10210 (N_10210,N_7642,N_8476);
nor U10211 (N_10211,N_7953,N_8025);
or U10212 (N_10212,N_8204,N_8943);
or U10213 (N_10213,N_8075,N_8488);
xor U10214 (N_10214,N_8682,N_9004);
nand U10215 (N_10215,N_7772,N_8780);
and U10216 (N_10216,N_9223,N_9884);
nor U10217 (N_10217,N_8631,N_9809);
xor U10218 (N_10218,N_8805,N_9084);
and U10219 (N_10219,N_8899,N_9625);
nor U10220 (N_10220,N_9482,N_9905);
nor U10221 (N_10221,N_9637,N_9503);
and U10222 (N_10222,N_8689,N_8575);
or U10223 (N_10223,N_9057,N_9254);
nand U10224 (N_10224,N_7574,N_8222);
nor U10225 (N_10225,N_8415,N_7547);
or U10226 (N_10226,N_7600,N_8813);
and U10227 (N_10227,N_8190,N_7946);
and U10228 (N_10228,N_7668,N_7554);
xor U10229 (N_10229,N_9058,N_9588);
nand U10230 (N_10230,N_9316,N_8591);
nand U10231 (N_10231,N_9544,N_8122);
nor U10232 (N_10232,N_9227,N_7503);
and U10233 (N_10233,N_8989,N_9280);
or U10234 (N_10234,N_8210,N_7767);
xnor U10235 (N_10235,N_8003,N_7792);
nor U10236 (N_10236,N_9613,N_9329);
nor U10237 (N_10237,N_8043,N_8900);
nor U10238 (N_10238,N_9150,N_8733);
or U10239 (N_10239,N_7597,N_8352);
and U10240 (N_10240,N_8779,N_8769);
and U10241 (N_10241,N_8540,N_9707);
and U10242 (N_10242,N_8702,N_8203);
nand U10243 (N_10243,N_8560,N_9988);
and U10244 (N_10244,N_9914,N_8875);
or U10245 (N_10245,N_9770,N_7592);
xnor U10246 (N_10246,N_9308,N_7602);
nand U10247 (N_10247,N_7750,N_8727);
nand U10248 (N_10248,N_9501,N_9630);
nor U10249 (N_10249,N_7803,N_8499);
nor U10250 (N_10250,N_9851,N_9417);
nand U10251 (N_10251,N_9747,N_8549);
or U10252 (N_10252,N_8619,N_8152);
or U10253 (N_10253,N_7992,N_8094);
or U10254 (N_10254,N_7695,N_8274);
nand U10255 (N_10255,N_9349,N_9957);
and U10256 (N_10256,N_9587,N_9039);
and U10257 (N_10257,N_8823,N_9757);
xor U10258 (N_10258,N_9287,N_9471);
nand U10259 (N_10259,N_8558,N_8041);
nor U10260 (N_10260,N_9721,N_7715);
nor U10261 (N_10261,N_8681,N_9255);
and U10262 (N_10262,N_9595,N_8506);
nand U10263 (N_10263,N_8485,N_8240);
and U10264 (N_10264,N_8257,N_9889);
or U10265 (N_10265,N_8686,N_9285);
nor U10266 (N_10266,N_7565,N_8798);
or U10267 (N_10267,N_8615,N_9769);
xnor U10268 (N_10268,N_9154,N_7672);
or U10269 (N_10269,N_9551,N_9406);
and U10270 (N_10270,N_9252,N_9298);
or U10271 (N_10271,N_8662,N_9355);
xor U10272 (N_10272,N_9100,N_9314);
and U10273 (N_10273,N_9136,N_9627);
or U10274 (N_10274,N_8425,N_8604);
or U10275 (N_10275,N_9454,N_9196);
nor U10276 (N_10276,N_7631,N_8364);
and U10277 (N_10277,N_9063,N_7798);
nor U10278 (N_10278,N_8277,N_8478);
nand U10279 (N_10279,N_7854,N_7910);
and U10280 (N_10280,N_8412,N_9910);
and U10281 (N_10281,N_8818,N_9605);
nor U10282 (N_10282,N_7994,N_9428);
nor U10283 (N_10283,N_9214,N_7667);
nor U10284 (N_10284,N_7749,N_9047);
and U10285 (N_10285,N_8695,N_7675);
nor U10286 (N_10286,N_8827,N_7542);
xor U10287 (N_10287,N_8298,N_7920);
nand U10288 (N_10288,N_9751,N_7951);
xnor U10289 (N_10289,N_8786,N_8986);
and U10290 (N_10290,N_8990,N_9007);
xor U10291 (N_10291,N_8960,N_9938);
and U10292 (N_10292,N_9077,N_8583);
nor U10293 (N_10293,N_7860,N_8367);
nor U10294 (N_10294,N_7555,N_8670);
nor U10295 (N_10295,N_8938,N_7685);
nor U10296 (N_10296,N_9506,N_9881);
and U10297 (N_10297,N_7641,N_8719);
and U10298 (N_10298,N_9644,N_8628);
and U10299 (N_10299,N_9681,N_8570);
or U10300 (N_10300,N_9813,N_8378);
and U10301 (N_10301,N_9928,N_8230);
xnor U10302 (N_10302,N_8967,N_7684);
nor U10303 (N_10303,N_8166,N_8486);
xor U10304 (N_10304,N_9338,N_9600);
and U10305 (N_10305,N_8582,N_8890);
or U10306 (N_10306,N_9779,N_7968);
or U10307 (N_10307,N_7500,N_8198);
or U10308 (N_10308,N_9051,N_8878);
and U10309 (N_10309,N_9727,N_7979);
xnor U10310 (N_10310,N_9592,N_8359);
xor U10311 (N_10311,N_9865,N_7736);
xnor U10312 (N_10312,N_9697,N_9155);
nand U10313 (N_10313,N_9824,N_8197);
nor U10314 (N_10314,N_9717,N_9931);
nor U10315 (N_10315,N_9645,N_9762);
nor U10316 (N_10316,N_8968,N_8437);
and U10317 (N_10317,N_9724,N_9556);
nor U10318 (N_10318,N_7637,N_7628);
nor U10319 (N_10319,N_7948,N_8579);
xnor U10320 (N_10320,N_9241,N_8340);
or U10321 (N_10321,N_8226,N_9410);
nor U10322 (N_10322,N_8072,N_8642);
xnor U10323 (N_10323,N_9438,N_9803);
xnor U10324 (N_10324,N_9540,N_9729);
or U10325 (N_10325,N_9991,N_9450);
and U10326 (N_10326,N_8555,N_9868);
or U10327 (N_10327,N_9165,N_8757);
nand U10328 (N_10328,N_9408,N_8620);
xor U10329 (N_10329,N_9333,N_8687);
and U10330 (N_10330,N_9485,N_7702);
or U10331 (N_10331,N_9277,N_8268);
or U10332 (N_10332,N_9774,N_9507);
nand U10333 (N_10333,N_9151,N_8600);
xnor U10334 (N_10334,N_7678,N_7783);
nor U10335 (N_10335,N_8587,N_7873);
or U10336 (N_10336,N_9461,N_9496);
nor U10337 (N_10337,N_8498,N_7896);
nor U10338 (N_10338,N_9098,N_8363);
nand U10339 (N_10339,N_8068,N_8708);
nor U10340 (N_10340,N_9426,N_7624);
or U10341 (N_10341,N_8503,N_9016);
nand U10342 (N_10342,N_8234,N_9200);
nand U10343 (N_10343,N_7723,N_9977);
nand U10344 (N_10344,N_8955,N_9499);
or U10345 (N_10345,N_7691,N_8296);
nand U10346 (N_10346,N_7827,N_7687);
or U10347 (N_10347,N_7816,N_9906);
nand U10348 (N_10348,N_7794,N_8436);
nand U10349 (N_10349,N_8060,N_9270);
and U10350 (N_10350,N_9201,N_8469);
or U10351 (N_10351,N_7673,N_8126);
or U10352 (N_10352,N_8801,N_8851);
nor U10353 (N_10353,N_9755,N_8286);
nand U10354 (N_10354,N_7603,N_9926);
nand U10355 (N_10355,N_9127,N_9913);
nor U10356 (N_10356,N_9631,N_8988);
or U10357 (N_10357,N_8763,N_8822);
nand U10358 (N_10358,N_9716,N_8181);
xnor U10359 (N_10359,N_8428,N_9346);
xnor U10360 (N_10360,N_9879,N_9373);
or U10361 (N_10361,N_8608,N_7644);
xnor U10362 (N_10362,N_9457,N_9326);
and U10363 (N_10363,N_8846,N_8520);
nor U10364 (N_10364,N_9647,N_8264);
or U10365 (N_10365,N_8462,N_9321);
and U10366 (N_10366,N_8111,N_8784);
xnor U10367 (N_10367,N_9447,N_7698);
nor U10368 (N_10368,N_9341,N_8731);
nor U10369 (N_10369,N_9965,N_9974);
and U10370 (N_10370,N_8921,N_8863);
or U10371 (N_10371,N_7502,N_8475);
nor U10372 (N_10372,N_9782,N_9393);
or U10373 (N_10373,N_7797,N_9650);
nor U10374 (N_10374,N_8052,N_7710);
or U10375 (N_10375,N_8444,N_8741);
nand U10376 (N_10376,N_8652,N_7781);
nor U10377 (N_10377,N_7786,N_7814);
xor U10378 (N_10378,N_8149,N_7895);
and U10379 (N_10379,N_9930,N_8081);
or U10380 (N_10380,N_7533,N_9804);
nand U10381 (N_10381,N_9398,N_8792);
or U10382 (N_10382,N_8115,N_9106);
and U10383 (N_10383,N_9369,N_9147);
nor U10384 (N_10384,N_9849,N_9514);
nand U10385 (N_10385,N_8411,N_9248);
and U10386 (N_10386,N_9885,N_7614);
nand U10387 (N_10387,N_7844,N_8070);
and U10388 (N_10388,N_8932,N_8079);
nand U10389 (N_10389,N_8429,N_7971);
nand U10390 (N_10390,N_8518,N_9000);
nand U10391 (N_10391,N_8743,N_8935);
or U10392 (N_10392,N_9121,N_9108);
nor U10393 (N_10393,N_9510,N_8135);
or U10394 (N_10394,N_9901,N_9086);
nor U10395 (N_10395,N_7847,N_9246);
xnor U10396 (N_10396,N_9972,N_8399);
and U10397 (N_10397,N_8430,N_7833);
and U10398 (N_10398,N_7619,N_9783);
nand U10399 (N_10399,N_9480,N_7681);
or U10400 (N_10400,N_9463,N_9114);
or U10401 (N_10401,N_7837,N_9193);
xnor U10402 (N_10402,N_7583,N_8040);
nand U10403 (N_10403,N_7944,N_8371);
nand U10404 (N_10404,N_9713,N_8262);
or U10405 (N_10405,N_7615,N_8235);
nor U10406 (N_10406,N_8904,N_9436);
or U10407 (N_10407,N_9520,N_8694);
xnor U10408 (N_10408,N_9832,N_7505);
or U10409 (N_10409,N_9403,N_9135);
or U10410 (N_10410,N_8973,N_9312);
and U10411 (N_10411,N_8588,N_7795);
and U10412 (N_10412,N_8958,N_8305);
or U10413 (N_10413,N_8250,N_9042);
nor U10414 (N_10414,N_9511,N_8956);
and U10415 (N_10415,N_8716,N_7728);
nor U10416 (N_10416,N_9213,N_8961);
nor U10417 (N_10417,N_8996,N_7601);
nand U10418 (N_10418,N_8188,N_8306);
xnor U10419 (N_10419,N_8703,N_8740);
xor U10420 (N_10420,N_8258,N_9677);
nand U10421 (N_10421,N_7526,N_9577);
nand U10422 (N_10422,N_9443,N_8815);
or U10423 (N_10423,N_8233,N_7987);
nand U10424 (N_10424,N_7993,N_9089);
and U10425 (N_10425,N_7976,N_9619);
nor U10426 (N_10426,N_9950,N_8354);
xnor U10427 (N_10427,N_9074,N_8944);
nand U10428 (N_10428,N_8142,N_8118);
xnor U10429 (N_10429,N_8002,N_9294);
or U10430 (N_10430,N_8151,N_8150);
or U10431 (N_10431,N_8881,N_9432);
and U10432 (N_10432,N_7894,N_7626);
nor U10433 (N_10433,N_9187,N_9648);
xnor U10434 (N_10434,N_8322,N_8334);
or U10435 (N_10435,N_9476,N_8265);
nand U10436 (N_10436,N_7513,N_9907);
nand U10437 (N_10437,N_9458,N_8069);
and U10438 (N_10438,N_9575,N_7518);
xor U10439 (N_10439,N_9186,N_8046);
and U10440 (N_10440,N_9574,N_9976);
nand U10441 (N_10441,N_9006,N_7892);
or U10442 (N_10442,N_7867,N_7802);
xnor U10443 (N_10443,N_9900,N_8267);
xor U10444 (N_10444,N_9464,N_8100);
or U10445 (N_10445,N_8237,N_8330);
xor U10446 (N_10446,N_8344,N_9189);
and U10447 (N_10447,N_8328,N_8123);
or U10448 (N_10448,N_8247,N_7874);
nor U10449 (N_10449,N_9033,N_8857);
or U10450 (N_10450,N_9500,N_9133);
and U10451 (N_10451,N_9912,N_9584);
and U10452 (N_10452,N_9315,N_8574);
and U10453 (N_10453,N_9908,N_7907);
and U10454 (N_10454,N_8385,N_9875);
xnor U10455 (N_10455,N_8725,N_8933);
nand U10456 (N_10456,N_9799,N_9470);
nor U10457 (N_10457,N_9259,N_9903);
and U10458 (N_10458,N_8414,N_7764);
and U10459 (N_10459,N_7552,N_8684);
and U10460 (N_10460,N_7564,N_9069);
nor U10461 (N_10461,N_9793,N_8707);
and U10462 (N_10462,N_9348,N_9162);
nand U10463 (N_10463,N_7884,N_9128);
and U10464 (N_10464,N_9841,N_9839);
and U10465 (N_10465,N_8886,N_8132);
and U10466 (N_10466,N_9429,N_9983);
xnor U10467 (N_10467,N_7612,N_9734);
and U10468 (N_10468,N_9561,N_9853);
or U10469 (N_10469,N_8675,N_9292);
or U10470 (N_10470,N_7525,N_9466);
nor U10471 (N_10471,N_8400,N_9874);
nor U10472 (N_10472,N_9547,N_9120);
nand U10473 (N_10473,N_9435,N_7535);
xnor U10474 (N_10474,N_9379,N_7625);
and U10475 (N_10475,N_9093,N_9391);
or U10476 (N_10476,N_9565,N_7534);
xnor U10477 (N_10477,N_8335,N_9508);
and U10478 (N_10478,N_9792,N_8572);
and U10479 (N_10479,N_8033,N_9634);
nand U10480 (N_10480,N_7763,N_9568);
xor U10481 (N_10481,N_7664,N_8569);
or U10482 (N_10482,N_8730,N_7627);
nand U10483 (N_10483,N_9694,N_8880);
nor U10484 (N_10484,N_9594,N_7881);
or U10485 (N_10485,N_7765,N_8129);
nand U10486 (N_10486,N_9347,N_9687);
and U10487 (N_10487,N_9798,N_8737);
nor U10488 (N_10488,N_9421,N_9388);
xnor U10489 (N_10489,N_7954,N_7871);
nand U10490 (N_10490,N_8744,N_9390);
nand U10491 (N_10491,N_8245,N_7510);
nor U10492 (N_10492,N_7509,N_8829);
and U10493 (N_10493,N_7726,N_9442);
and U10494 (N_10494,N_7665,N_8034);
or U10495 (N_10495,N_7862,N_7530);
or U10496 (N_10496,N_9366,N_9119);
nor U10497 (N_10497,N_7682,N_7645);
nand U10498 (N_10498,N_8516,N_8061);
nand U10499 (N_10499,N_9052,N_8001);
xor U10500 (N_10500,N_9545,N_8551);
xnor U10501 (N_10501,N_8911,N_9256);
xnor U10502 (N_10502,N_9357,N_8905);
nor U10503 (N_10503,N_8282,N_9225);
or U10504 (N_10504,N_9935,N_9959);
nand U10505 (N_10505,N_9251,N_7507);
nor U10506 (N_10506,N_9174,N_8249);
nor U10507 (N_10507,N_7980,N_9376);
nor U10508 (N_10508,N_9936,N_7891);
nor U10509 (N_10509,N_9835,N_9966);
nor U10510 (N_10510,N_9258,N_8545);
and U10511 (N_10511,N_7928,N_8995);
or U10512 (N_10512,N_9754,N_8242);
or U10513 (N_10513,N_7810,N_7790);
and U10514 (N_10514,N_9159,N_9413);
nor U10515 (N_10515,N_7815,N_9371);
nor U10516 (N_10516,N_8148,N_8833);
nand U10517 (N_10517,N_7970,N_8552);
and U10518 (N_10518,N_7737,N_7739);
xnor U10519 (N_10519,N_8934,N_7751);
or U10520 (N_10520,N_8390,N_8317);
or U10521 (N_10521,N_7935,N_9233);
nand U10522 (N_10522,N_7670,N_9116);
xnor U10523 (N_10523,N_7701,N_9205);
and U10524 (N_10524,N_8848,N_8538);
and U10525 (N_10525,N_8372,N_8057);
nor U10526 (N_10526,N_8244,N_8855);
or U10527 (N_10527,N_7924,N_9730);
and U10528 (N_10528,N_9736,N_7880);
nand U10529 (N_10529,N_8508,N_8105);
or U10530 (N_10530,N_9869,N_9284);
or U10531 (N_10531,N_9602,N_9640);
nand U10532 (N_10532,N_8278,N_8055);
nand U10533 (N_10533,N_8640,N_9216);
nor U10534 (N_10534,N_7523,N_9149);
and U10535 (N_10535,N_8860,N_8914);
and U10536 (N_10536,N_8023,N_8309);
or U10537 (N_10537,N_8632,N_8256);
or U10538 (N_10538,N_7585,N_9325);
xnor U10539 (N_10539,N_9335,N_8736);
xor U10540 (N_10540,N_8993,N_9780);
or U10541 (N_10541,N_9802,N_9240);
nor U10542 (N_10542,N_8221,N_7529);
nor U10543 (N_10543,N_9700,N_9024);
and U10544 (N_10544,N_9666,N_9243);
xnor U10545 (N_10545,N_9599,N_9639);
xnor U10546 (N_10546,N_8625,N_8468);
nor U10547 (N_10547,N_7720,N_9609);
xor U10548 (N_10548,N_9720,N_9646);
xnor U10549 (N_10549,N_7866,N_7758);
nor U10550 (N_10550,N_7836,N_9773);
and U10551 (N_10551,N_9117,N_9260);
nand U10552 (N_10552,N_8690,N_9847);
xnor U10553 (N_10553,N_8866,N_8481);
and U10554 (N_10554,N_9791,N_7828);
nor U10555 (N_10555,N_9377,N_9955);
nand U10556 (N_10556,N_7578,N_8648);
nand U10557 (N_10557,N_9020,N_9969);
nand U10558 (N_10558,N_8199,N_8269);
nand U10559 (N_10559,N_8952,N_8139);
or U10560 (N_10560,N_9273,N_9923);
nand U10561 (N_10561,N_9484,N_8077);
nand U10562 (N_10562,N_7890,N_8673);
or U10563 (N_10563,N_8724,N_9553);
nand U10564 (N_10564,N_7840,N_8382);
and U10565 (N_10565,N_9542,N_7731);
xnor U10566 (N_10566,N_7556,N_8850);
nor U10567 (N_10567,N_7909,N_9295);
or U10568 (N_10568,N_8116,N_9961);
and U10569 (N_10569,N_8165,N_8660);
xnor U10570 (N_10570,N_9035,N_7658);
nand U10571 (N_10571,N_8284,N_9549);
nand U10572 (N_10572,N_9967,N_8715);
nor U10573 (N_10573,N_7782,N_8659);
nor U10574 (N_10574,N_9855,N_9897);
and U10575 (N_10575,N_7683,N_7888);
or U10576 (N_10576,N_9477,N_9846);
nor U10577 (N_10577,N_9693,N_9728);
nand U10578 (N_10578,N_7914,N_8010);
xor U10579 (N_10579,N_8346,N_9336);
nand U10580 (N_10580,N_8091,N_9714);
nor U10581 (N_10581,N_8653,N_9990);
nor U10582 (N_10582,N_8528,N_9812);
xor U10583 (N_10583,N_9559,N_9045);
nor U10584 (N_10584,N_9386,N_8945);
or U10585 (N_10585,N_8031,N_7738);
nor U10586 (N_10586,N_7825,N_8869);
nand U10587 (N_10587,N_9641,N_9245);
xnor U10588 (N_10588,N_7959,N_9777);
nor U10589 (N_10589,N_7865,N_9286);
xnor U10590 (N_10590,N_8195,N_7522);
xnor U10591 (N_10591,N_9467,N_9365);
nand U10592 (N_10592,N_8327,N_8922);
nand U10593 (N_10593,N_7789,N_9053);
nand U10594 (N_10594,N_9370,N_7653);
nor U10595 (N_10595,N_8903,N_8289);
and U10596 (N_10596,N_7945,N_8474);
or U10597 (N_10597,N_7694,N_8760);
nor U10598 (N_10598,N_9180,N_8457);
nand U10599 (N_10599,N_9002,N_8466);
nor U10600 (N_10600,N_8458,N_8882);
nor U10601 (N_10601,N_8820,N_9183);
nor U10602 (N_10602,N_8293,N_8440);
nand U10603 (N_10603,N_8090,N_9621);
nor U10604 (N_10604,N_7573,N_8164);
or U10605 (N_10605,N_9682,N_9404);
and U10606 (N_10606,N_9179,N_9099);
xnor U10607 (N_10607,N_7813,N_8791);
or U10608 (N_10608,N_8112,N_8680);
nand U10609 (N_10609,N_9402,N_9445);
or U10610 (N_10610,N_8999,N_9263);
nand U10611 (N_10611,N_9409,N_8178);
and U10612 (N_10612,N_9434,N_8979);
nor U10613 (N_10613,N_7632,N_8861);
nand U10614 (N_10614,N_8134,N_8239);
nor U10615 (N_10615,N_8700,N_8026);
and U10616 (N_10616,N_8360,N_8155);
nor U10617 (N_10617,N_8732,N_9899);
nor U10618 (N_10618,N_8208,N_9695);
xor U10619 (N_10619,N_8211,N_9993);
and U10620 (N_10620,N_8051,N_9130);
nand U10621 (N_10621,N_9786,N_8832);
nor U10622 (N_10622,N_8379,N_7549);
nand U10623 (N_10623,N_8785,N_8279);
nand U10624 (N_10624,N_8270,N_8493);
nand U10625 (N_10625,N_9539,N_9519);
nand U10626 (N_10626,N_7610,N_9198);
xnor U10627 (N_10627,N_9212,N_7925);
or U10628 (N_10628,N_8592,N_8156);
and U10629 (N_10629,N_8017,N_9537);
xor U10630 (N_10630,N_7575,N_8124);
or U10631 (N_10631,N_9939,N_9672);
nand U10632 (N_10632,N_7746,N_7856);
or U10633 (N_10633,N_8225,N_7989);
nor U10634 (N_10634,N_8984,N_9218);
nand U10635 (N_10635,N_9337,N_8666);
and U10636 (N_10636,N_8018,N_9230);
and U10637 (N_10637,N_9411,N_8974);
xnor U10638 (N_10638,N_8871,N_9902);
nor U10639 (N_10639,N_8170,N_8826);
nor U10640 (N_10640,N_8263,N_9399);
or U10641 (N_10641,N_8550,N_8217);
nand U10642 (N_10642,N_8062,N_9163);
and U10643 (N_10643,N_8892,N_7900);
nand U10644 (N_10644,N_8243,N_9414);
nand U10645 (N_10645,N_9745,N_7973);
xor U10646 (N_10646,N_7778,N_9146);
or U10647 (N_10647,N_9142,N_9945);
or U10648 (N_10648,N_8227,N_8835);
and U10649 (N_10649,N_8618,N_7514);
or U10650 (N_10650,N_8492,N_7829);
and U10651 (N_10651,N_9037,N_8494);
or U10652 (N_10652,N_8676,N_8231);
and U10653 (N_10653,N_8087,N_9554);
xnor U10654 (N_10654,N_9615,N_7893);
nor U10655 (N_10655,N_8410,N_8865);
nand U10656 (N_10656,N_7543,N_8568);
nand U10657 (N_10657,N_7811,N_9304);
nand U10658 (N_10658,N_9843,N_8782);
nand U10659 (N_10659,N_7947,N_9784);
and U10660 (N_10660,N_8885,N_8610);
and U10661 (N_10661,N_9038,N_9741);
xnor U10662 (N_10662,N_8910,N_8187);
and U10663 (N_10663,N_8870,N_8064);
xnor U10664 (N_10664,N_8201,N_9509);
nand U10665 (N_10665,N_9686,N_8888);
and U10666 (N_10666,N_8924,N_7655);
and U10667 (N_10667,N_9632,N_9068);
nor U10668 (N_10668,N_8276,N_7747);
and U10669 (N_10669,N_8928,N_7957);
nor U10670 (N_10670,N_7952,N_8012);
xnor U10671 (N_10671,N_7908,N_7704);
nor U10672 (N_10672,N_8417,N_8248);
and U10673 (N_10673,N_7923,N_9940);
or U10674 (N_10674,N_8356,N_9921);
nand U10675 (N_10675,N_7921,N_7809);
nand U10676 (N_10676,N_9027,N_7966);
xnor U10677 (N_10677,N_8722,N_7916);
or U10678 (N_10678,N_7689,N_9663);
or U10679 (N_10679,N_9876,N_9097);
or U10680 (N_10680,N_9748,N_9659);
and U10681 (N_10681,N_9059,N_7544);
nand U10682 (N_10682,N_9522,N_8074);
nor U10683 (N_10683,N_9567,N_9276);
or U10684 (N_10684,N_7897,N_9491);
nand U10685 (N_10685,N_8772,N_9046);
nand U10686 (N_10686,N_9028,N_8158);
or U10687 (N_10687,N_8781,N_7982);
and U10688 (N_10688,N_7853,N_9564);
nor U10689 (N_10689,N_7787,N_7577);
xnor U10690 (N_10690,N_9852,N_9465);
xnor U10691 (N_10691,N_8567,N_7757);
and U10692 (N_10692,N_7680,N_8128);
and U10693 (N_10693,N_8788,N_7905);
or U10694 (N_10694,N_8349,N_7650);
nor U10695 (N_10695,N_9094,N_9998);
and U10696 (N_10696,N_9319,N_8898);
nand U10697 (N_10697,N_8207,N_7654);
and U10698 (N_10698,N_9572,N_7519);
nand U10699 (N_10699,N_9137,N_8809);
nor U10700 (N_10700,N_8571,N_8711);
and U10701 (N_10701,N_9160,N_7831);
nand U10702 (N_10702,N_8271,N_7796);
and U10703 (N_10703,N_7734,N_7697);
or U10704 (N_10704,N_9756,N_8173);
nand U10705 (N_10705,N_9712,N_8389);
and U10706 (N_10706,N_8441,N_8997);
nor U10707 (N_10707,N_8451,N_8811);
or U10708 (N_10708,N_8176,N_7933);
nor U10709 (N_10709,N_9342,N_9845);
nor U10710 (N_10710,N_8721,N_8524);
or U10711 (N_10711,N_8771,N_9204);
nand U10712 (N_10712,N_7978,N_7770);
nand U10713 (N_10713,N_9040,N_9664);
nand U10714 (N_10714,N_7652,N_8606);
xnor U10715 (N_10715,N_9916,N_9871);
nand U10716 (N_10716,N_9268,N_9624);
nand U10717 (N_10717,N_7609,N_9530);
nand U10718 (N_10718,N_9126,N_7721);
or U10719 (N_10719,N_8180,N_9661);
or U10720 (N_10720,N_8917,N_9512);
nor U10721 (N_10721,N_9767,N_8748);
nand U10722 (N_10722,N_7613,N_7640);
xnor U10723 (N_10723,N_7748,N_9018);
or U10724 (N_10724,N_9382,N_7775);
nand U10725 (N_10725,N_9560,N_7707);
or U10726 (N_10726,N_7963,N_7699);
nand U10727 (N_10727,N_7617,N_8800);
nand U10728 (N_10728,N_7969,N_9956);
and U10729 (N_10729,N_7571,N_9178);
or U10730 (N_10730,N_8369,N_7528);
xnor U10731 (N_10731,N_7986,N_7643);
nor U10732 (N_10732,N_8251,N_8959);
nor U10733 (N_10733,N_7872,N_8998);
or U10734 (N_10734,N_8216,N_7804);
nand U10735 (N_10735,N_8634,N_8893);
xnor U10736 (N_10736,N_8581,N_9985);
xor U10737 (N_10737,N_9080,N_7633);
nor U10738 (N_10738,N_8957,N_8854);
nor U10739 (N_10739,N_9420,N_9997);
nor U10740 (N_10740,N_8720,N_8168);
and U10741 (N_10741,N_9339,N_9877);
nor U10742 (N_10742,N_8450,N_9237);
nand U10743 (N_10743,N_9994,N_8140);
xnor U10744 (N_10744,N_7594,N_9164);
nor U10745 (N_10745,N_8275,N_9618);
or U10746 (N_10746,N_8726,N_9264);
xor U10747 (N_10747,N_9231,N_7716);
or U10748 (N_10748,N_9806,N_9676);
nand U10749 (N_10749,N_9704,N_9202);
nor U10750 (N_10750,N_8147,N_9775);
nand U10751 (N_10751,N_9257,N_9895);
nor U10752 (N_10752,N_7590,N_8024);
or U10753 (N_10753,N_8053,N_8443);
or U10754 (N_10754,N_9660,N_7972);
or U10755 (N_10755,N_9143,N_9968);
nand U10756 (N_10756,N_7516,N_9066);
and U10757 (N_10757,N_9984,N_8747);
xnor U10758 (N_10758,N_9169,N_9124);
or U10759 (N_10759,N_9103,N_8141);
xor U10760 (N_10760,N_9944,N_9848);
and U10761 (N_10761,N_9941,N_9495);
or U10762 (N_10762,N_7735,N_9274);
and U10763 (N_10763,N_7807,N_7561);
and U10764 (N_10764,N_9683,N_7819);
and U10765 (N_10765,N_9772,N_9962);
xnor U10766 (N_10766,N_8764,N_9684);
xor U10767 (N_10767,N_7622,N_8144);
nor U10768 (N_10768,N_8542,N_8102);
nand U10769 (N_10769,N_9808,N_8793);
or U10770 (N_10770,N_9829,N_7692);
nor U10771 (N_10771,N_8491,N_7589);
nand U10772 (N_10772,N_7913,N_9917);
nor U10773 (N_10773,N_7832,N_9323);
and U10774 (N_10774,N_7902,N_9827);
nor U10775 (N_10775,N_9596,N_8343);
and U10776 (N_10776,N_8096,N_9576);
xnor U10777 (N_10777,N_7709,N_8585);
nor U10778 (N_10778,N_7955,N_7927);
nand U10779 (N_10779,N_8517,N_8976);
and U10780 (N_10780,N_9049,N_7669);
or U10781 (N_10781,N_8655,N_9764);
and U10782 (N_10782,N_8044,N_9111);
xor U10783 (N_10783,N_8795,N_8117);
nand U10784 (N_10784,N_9723,N_9742);
nand U10785 (N_10785,N_9232,N_8638);
nand U10786 (N_10786,N_8391,N_9924);
or U10787 (N_10787,N_8902,N_8643);
nand U10788 (N_10788,N_9738,N_8629);
and U10789 (N_10789,N_9711,N_8641);
nand U10790 (N_10790,N_9134,N_9350);
nor U10791 (N_10791,N_9104,N_7634);
nor U10792 (N_10792,N_8983,N_8929);
nor U10793 (N_10793,N_9788,N_9221);
and U10794 (N_10794,N_8776,N_8032);
and U10795 (N_10795,N_8167,N_9138);
nand U10796 (N_10796,N_7620,N_9228);
and U10797 (N_10797,N_9061,N_8734);
and U10798 (N_10798,N_9705,N_9766);
or U10799 (N_10799,N_9299,N_7570);
xor U10800 (N_10800,N_7929,N_8202);
xor U10801 (N_10801,N_9055,N_9381);
nand U10802 (N_10802,N_8472,N_7677);
xnor U10803 (N_10803,N_9013,N_8067);
xnor U10804 (N_10804,N_7774,N_8531);
xor U10805 (N_10805,N_8027,N_7646);
and U10806 (N_10806,N_8283,N_7838);
nand U10807 (N_10807,N_9933,N_9973);
and U10808 (N_10808,N_7674,N_8273);
or U10809 (N_10809,N_9439,N_8099);
nor U10810 (N_10810,N_9718,N_8223);
and U10811 (N_10811,N_9440,N_9759);
nand U10812 (N_10812,N_7511,N_9992);
xor U10813 (N_10813,N_8477,N_8992);
or U10814 (N_10814,N_9611,N_9181);
nand U10815 (N_10815,N_9209,N_8796);
xor U10816 (N_10816,N_7917,N_8821);
and U10817 (N_10817,N_8981,N_8894);
nand U10818 (N_10818,N_7639,N_8953);
xor U10819 (N_10819,N_9761,N_8453);
nand U10820 (N_10820,N_8182,N_8238);
nor U10821 (N_10821,N_9161,N_9964);
and U10822 (N_10822,N_7688,N_8773);
xnor U10823 (N_10823,N_8537,N_7722);
nor U10824 (N_10824,N_8844,N_9831);
or U10825 (N_10825,N_7846,N_7712);
nand U10826 (N_10826,N_8948,N_7501);
nor U10827 (N_10827,N_8291,N_8563);
and U10828 (N_10828,N_8401,N_8329);
xor U10829 (N_10829,N_9392,N_9328);
nand U10830 (N_10830,N_7569,N_8837);
and U10831 (N_10831,N_9948,N_8704);
nand U10832 (N_10832,N_9834,N_8541);
or U10833 (N_10833,N_7693,N_9698);
and U10834 (N_10834,N_9573,N_9431);
and U10835 (N_10835,N_8028,N_9517);
or U10836 (N_10836,N_9989,N_9904);
and U10837 (N_10837,N_8396,N_9056);
or U10838 (N_10838,N_8048,N_9504);
or U10839 (N_10839,N_9585,N_7800);
and U10840 (N_10840,N_7730,N_8502);
xnor U10841 (N_10841,N_9244,N_8482);
or U10842 (N_10842,N_7849,N_8054);
or U10843 (N_10843,N_8873,N_7806);
or U10844 (N_10844,N_9469,N_8253);
and U10845 (N_10845,N_9678,N_9765);
nor U10846 (N_10846,N_8036,N_7882);
and U10847 (N_10847,N_8311,N_8637);
xnor U10848 (N_10848,N_7868,N_9746);
and U10849 (N_10849,N_8205,N_8504);
or U10850 (N_10850,N_8029,N_7579);
nor U10851 (N_10851,N_7662,N_8007);
or U10852 (N_10852,N_8375,N_9125);
or U10853 (N_10853,N_8767,N_9265);
nor U10854 (N_10854,N_9934,N_9797);
xor U10855 (N_10855,N_8157,N_8557);
or U10856 (N_10856,N_8577,N_9356);
or U10857 (N_10857,N_7686,N_9460);
or U10858 (N_10858,N_9800,N_8092);
nand U10859 (N_10859,N_8019,N_8014);
nand U10860 (N_10860,N_8008,N_7938);
or U10861 (N_10861,N_9022,N_9552);
and U10862 (N_10862,N_8138,N_9087);
nand U10863 (N_10863,N_7759,N_9234);
nand U10864 (N_10864,N_9320,N_9857);
xor U10865 (N_10865,N_8876,N_9222);
nor U10866 (N_10866,N_9975,N_8709);
xnor U10867 (N_10867,N_8665,N_8339);
nand U10868 (N_10868,N_8505,N_8130);
xor U10869 (N_10869,N_9692,N_8966);
nand U10870 (N_10870,N_9375,N_7531);
and U10871 (N_10871,N_8119,N_8526);
or U10872 (N_10872,N_8521,N_8095);
or U10873 (N_10873,N_8383,N_9195);
xor U10874 (N_10874,N_7717,N_8906);
nand U10875 (N_10875,N_9044,N_8977);
xnor U10876 (N_10876,N_7732,N_8080);
nor U10877 (N_10877,N_7937,N_9064);
nand U10878 (N_10878,N_9113,N_9896);
xnor U10879 (N_10879,N_8171,N_8975);
and U10880 (N_10880,N_9423,N_9490);
nor U10881 (N_10881,N_7863,N_9562);
nand U10882 (N_10882,N_9288,N_8775);
nor U10883 (N_10883,N_8137,N_7538);
and U10884 (N_10884,N_9952,N_9690);
nor U10885 (N_10885,N_9311,N_9612);
or U10886 (N_10886,N_9674,N_9534);
nor U10887 (N_10887,N_8059,N_8143);
and U10888 (N_10888,N_8645,N_8447);
and U10889 (N_10889,N_9468,N_9194);
nand U10890 (N_10890,N_9891,N_9656);
xor U10891 (N_10891,N_9132,N_7855);
xor U10892 (N_10892,N_8316,N_9942);
or U10893 (N_10893,N_9604,N_9122);
or U10894 (N_10894,N_8022,N_7762);
nand U10895 (N_10895,N_8397,N_8951);
or U10896 (N_10896,N_7942,N_9750);
nand U10897 (N_10897,N_8037,N_9807);
nor U10898 (N_10898,N_7918,N_9437);
nand U10899 (N_10899,N_9271,N_8464);
nand U10900 (N_10900,N_9071,N_8434);
nand U10901 (N_10901,N_9050,N_9590);
nor U10902 (N_10902,N_9362,N_8463);
nor U10903 (N_10903,N_7830,N_9383);
nor U10904 (N_10904,N_8416,N_7851);
xor U10905 (N_10905,N_9979,N_9025);
xnor U10906 (N_10906,N_9703,N_8500);
nand U10907 (N_10907,N_7962,N_7941);
nand U10908 (N_10908,N_7563,N_9844);
or U10909 (N_10909,N_9334,N_9479);
and U10910 (N_10910,N_9951,N_8564);
nor U10911 (N_10911,N_8459,N_9448);
or U10912 (N_10912,N_7912,N_9811);
or U10913 (N_10913,N_7580,N_9005);
and U10914 (N_10914,N_7657,N_9279);
nand U10915 (N_10915,N_8084,N_9034);
or U10916 (N_10916,N_8066,N_7604);
and U10917 (N_10917,N_7727,N_9278);
nor U10918 (N_10918,N_9653,N_8696);
and U10919 (N_10919,N_9502,N_8947);
nor U10920 (N_10920,N_8533,N_8312);
nor U10921 (N_10921,N_8535,N_9655);
nand U10922 (N_10922,N_9191,N_8603);
and U10923 (N_10923,N_9726,N_8362);
xor U10924 (N_10924,N_9521,N_7875);
and U10925 (N_10925,N_7761,N_8406);
and U10926 (N_10926,N_8565,N_9301);
nand U10927 (N_10927,N_8692,N_9669);
and U10928 (N_10928,N_7651,N_7517);
nand U10929 (N_10929,N_9419,N_9352);
and U10930 (N_10930,N_8916,N_9172);
or U10931 (N_10931,N_8738,N_7965);
or U10932 (N_10932,N_9079,N_7852);
nor U10933 (N_10933,N_9523,N_7988);
nor U10934 (N_10934,N_8101,N_8712);
and U10935 (N_10935,N_8897,N_9283);
or U10936 (N_10936,N_8816,N_7898);
xnor U10937 (N_10937,N_9433,N_8435);
nor U10938 (N_10938,N_9825,N_8654);
and U10939 (N_10939,N_8512,N_9394);
nor U10940 (N_10940,N_9197,N_7520);
nor U10941 (N_10941,N_8196,N_8758);
xor U10942 (N_10942,N_8887,N_7906);
nand U10943 (N_10943,N_8611,N_8623);
nor U10944 (N_10944,N_9689,N_8553);
xnor U10945 (N_10945,N_9253,N_8006);
xnor U10946 (N_10946,N_8460,N_9752);
and U10947 (N_10947,N_7605,N_8644);
nand U10948 (N_10948,N_7824,N_9282);
and U10949 (N_10949,N_7512,N_8646);
nand U10950 (N_10950,N_7719,N_8287);
xor U10951 (N_10951,N_9579,N_7859);
or U10952 (N_10952,N_9015,N_9070);
nor U10953 (N_10953,N_9867,N_7656);
and U10954 (N_10954,N_9012,N_9887);
or U10955 (N_10955,N_7711,N_9675);
or U10956 (N_10956,N_9929,N_9262);
xnor U10957 (N_10957,N_8962,N_9494);
nor U10958 (N_10958,N_8331,N_7964);
or U10959 (N_10959,N_7956,N_9790);
nand U10960 (N_10960,N_8907,N_8578);
nand U10961 (N_10961,N_7961,N_8418);
xor U10962 (N_10962,N_9581,N_8266);
and U10963 (N_10963,N_8872,N_8756);
and U10964 (N_10964,N_8083,N_7725);
nor U10965 (N_10965,N_9010,N_9614);
and U10966 (N_10966,N_8405,N_9247);
nand U10967 (N_10967,N_8345,N_9749);
xnor U10968 (N_10968,N_9236,N_9571);
or U10969 (N_10969,N_8376,N_9558);
nor U10970 (N_10970,N_7508,N_8590);
and U10971 (N_10971,N_8209,N_9091);
or U10972 (N_10972,N_8787,N_9801);
or U10973 (N_10973,N_7598,N_8206);
nand U10974 (N_10974,N_8131,N_8774);
nand U10975 (N_10975,N_8908,N_7551);
nor U10976 (N_10976,N_9300,N_9513);
nand U10977 (N_10977,N_8487,N_8490);
nor U10978 (N_10978,N_9840,N_9101);
xnor U10979 (N_10979,N_8302,N_8543);
xor U10980 (N_10980,N_8050,N_9837);
or U10981 (N_10981,N_7648,N_8589);
and U10982 (N_10982,N_9610,N_8701);
xnor U10983 (N_10983,N_9217,N_8501);
and U10984 (N_10984,N_9543,N_8136);
and U10985 (N_10985,N_9451,N_8970);
nor U10986 (N_10986,N_9528,N_7539);
or U10987 (N_10987,N_9327,N_9462);
xnor U10988 (N_10988,N_7967,N_9888);
or U10989 (N_10989,N_9144,N_9636);
nand U10990 (N_10990,N_9535,N_7724);
nor U10991 (N_10991,N_9566,N_8368);
xnor U10992 (N_10992,N_8042,N_9302);
or U10993 (N_10993,N_9999,N_8154);
and U10994 (N_10994,N_8868,N_7532);
nand U10995 (N_10995,N_9131,N_8093);
xor U10996 (N_10996,N_8452,N_8315);
nand U10997 (N_10997,N_7784,N_8937);
xor U10998 (N_10998,N_8656,N_8358);
and U10999 (N_10999,N_7788,N_8484);
nand U11000 (N_11000,N_9525,N_9859);
xor U11001 (N_11001,N_7861,N_9915);
nand U11002 (N_11002,N_8324,N_8946);
or U11003 (N_11003,N_9185,N_8454);
nand U11004 (N_11004,N_9023,N_9861);
or U11005 (N_11005,N_8366,N_8380);
nand U11006 (N_11006,N_9405,N_8489);
and U11007 (N_11007,N_9763,N_9668);
and U11008 (N_11008,N_8357,N_7636);
nand U11009 (N_11009,N_8016,N_9557);
xnor U11010 (N_11010,N_7703,N_7995);
nand U11011 (N_11011,N_9153,N_7690);
or U11012 (N_11012,N_8301,N_9188);
or U11013 (N_11013,N_8071,N_8723);
nand U11014 (N_11014,N_9425,N_8260);
or U11015 (N_11015,N_7845,N_9036);
nand U11016 (N_11016,N_9963,N_9821);
xnor U11017 (N_11017,N_8950,N_9397);
nand U11018 (N_11018,N_9332,N_9937);
and U11019 (N_11019,N_9481,N_9076);
or U11020 (N_11020,N_9911,N_9307);
nor U11021 (N_11021,N_8432,N_7679);
nor U11022 (N_11022,N_8599,N_7560);
xnor U11023 (N_11023,N_9589,N_7541);
nand U11024 (N_11024,N_7506,N_9427);
nand U11025 (N_11025,N_9836,N_7676);
or U11026 (N_11026,N_9215,N_9946);
or U11027 (N_11027,N_7623,N_9021);
and U11028 (N_11028,N_9658,N_8337);
nor U11029 (N_11029,N_8797,N_9586);
nor U11030 (N_11030,N_9890,N_8104);
and U11031 (N_11031,N_9157,N_8514);
or U11032 (N_11032,N_8318,N_9909);
or U11033 (N_11033,N_7671,N_8825);
and U11034 (N_11034,N_8063,N_9210);
or U11035 (N_11035,N_9970,N_9483);
or U11036 (N_11036,N_7587,N_9789);
nand U11037 (N_11037,N_8755,N_7848);
nor U11038 (N_11038,N_9828,N_8927);
nand U11039 (N_11039,N_8480,N_8442);
xor U11040 (N_11040,N_8699,N_9344);
nand U11041 (N_11041,N_8336,N_9092);
nand U11042 (N_11042,N_7843,N_7752);
or U11043 (N_11043,N_9810,N_9982);
xor U11044 (N_11044,N_8186,N_9662);
and U11045 (N_11045,N_9919,N_8925);
or U11046 (N_11046,N_7886,N_8114);
nand U11047 (N_11047,N_8987,N_8308);
or U11048 (N_11048,N_7536,N_7663);
xnor U11049 (N_11049,N_7595,N_9838);
nor U11050 (N_11050,N_7607,N_8455);
nor U11051 (N_11051,N_8843,N_7812);
nand U11052 (N_11052,N_9078,N_7885);
nand U11053 (N_11053,N_9816,N_8630);
xnor U11054 (N_11054,N_8566,N_8789);
and U11055 (N_11055,N_7718,N_8108);
xor U11056 (N_11056,N_8613,N_9322);
or U11057 (N_11057,N_9603,N_7932);
nand U11058 (N_11058,N_7878,N_8439);
xor U11059 (N_11059,N_8175,N_8338);
xnor U11060 (N_11060,N_8802,N_9368);
or U11061 (N_11061,N_9925,N_8918);
and U11062 (N_11062,N_8465,N_8313);
and U11063 (N_11063,N_7839,N_7566);
and U11064 (N_11064,N_8536,N_8669);
nor U11065 (N_11065,N_9148,N_9041);
or U11066 (N_11066,N_7584,N_8714);
nor U11067 (N_11067,N_8529,N_9580);
nor U11068 (N_11068,N_7649,N_9898);
nand U11069 (N_11069,N_8749,N_8949);
xor U11070 (N_11070,N_8333,N_7608);
nor U11071 (N_11071,N_9819,N_8824);
and U11072 (N_11072,N_7527,N_9167);
or U11073 (N_11073,N_9441,N_9546);
nand U11074 (N_11074,N_8146,N_7630);
xnor U11075 (N_11075,N_7582,N_9031);
nor U11076 (N_11076,N_8718,N_9158);
xor U11077 (N_11077,N_9239,N_8838);
xor U11078 (N_11078,N_7581,N_7743);
nor U11079 (N_11079,N_8433,N_8963);
xnor U11080 (N_11080,N_8806,N_9527);
and U11081 (N_11081,N_8576,N_8255);
and U11082 (N_11082,N_9306,N_8408);
nand U11083 (N_11083,N_9583,N_8650);
xor U11084 (N_11084,N_7706,N_8556);
or U11085 (N_11085,N_7801,N_8539);
nand U11086 (N_11086,N_8423,N_8706);
and U11087 (N_11087,N_8321,N_8596);
xnor U11088 (N_11088,N_7943,N_9665);
nand U11089 (N_11089,N_9019,N_8272);
nor U11090 (N_11090,N_9497,N_8325);
xnor U11091 (N_11091,N_8697,N_8622);
nor U11092 (N_11092,N_9696,N_8754);
nor U11093 (N_11093,N_9735,N_9009);
xor U11094 (N_11094,N_7618,N_9184);
or U11095 (N_11095,N_7835,N_8058);
nand U11096 (N_11096,N_7998,N_9771);
nand U11097 (N_11097,N_9269,N_8685);
or U11098 (N_11098,N_8739,N_9922);
and U11099 (N_11099,N_8804,N_8252);
nand U11100 (N_11100,N_9830,N_7823);
nand U11101 (N_11101,N_8799,N_9412);
nand U11102 (N_11102,N_7521,N_8761);
or U11103 (N_11103,N_8783,N_7621);
and U11104 (N_11104,N_8923,N_8683);
nand U11105 (N_11105,N_8830,N_7858);
nor U11106 (N_11106,N_8766,N_8595);
and U11107 (N_11107,N_8762,N_9593);
or U11108 (N_11108,N_9826,N_7745);
nor U11109 (N_11109,N_7901,N_7949);
and U11110 (N_11110,N_9170,N_9758);
nor U11111 (N_11111,N_9796,N_7568);
nand U11112 (N_11112,N_9152,N_8009);
nand U11113 (N_11113,N_8246,N_9418);
or U11114 (N_11114,N_9487,N_8978);
xnor U11115 (N_11115,N_8110,N_9017);
xor U11116 (N_11116,N_8969,N_9474);
nand U11117 (N_11117,N_8424,N_8420);
or U11118 (N_11118,N_8285,N_9987);
and U11119 (N_11119,N_7753,N_9708);
and U11120 (N_11120,N_9140,N_8290);
xnor U11121 (N_11121,N_8145,N_7791);
xor U11122 (N_11122,N_7616,N_8746);
or U11123 (N_11123,N_9395,N_8307);
nand U11124 (N_11124,N_8515,N_7926);
or U11125 (N_11125,N_9008,N_8350);
or U11126 (N_11126,N_9141,N_9563);
nor U11127 (N_11127,N_8082,N_8049);
nand U11128 (N_11128,N_7700,N_7996);
nand U11129 (N_11129,N_9156,N_8859);
xor U11130 (N_11130,N_8342,N_8413);
or U11131 (N_11131,N_9293,N_8456);
nand U11132 (N_11132,N_9679,N_9932);
nand U11133 (N_11133,N_8636,N_9960);
nor U11134 (N_11134,N_8047,N_8915);
or U11135 (N_11135,N_8403,N_7558);
or U11136 (N_11136,N_9850,N_8639);
xnor U11137 (N_11137,N_8421,N_8035);
nand U11138 (N_11138,N_7818,N_8794);
or U11139 (N_11139,N_7864,N_7799);
or U11140 (N_11140,N_9739,N_8753);
nor U11141 (N_11141,N_8679,N_9864);
xnor U11142 (N_11142,N_8532,N_8509);
nor U11143 (N_11143,N_9531,N_8303);
xor U11144 (N_11144,N_8678,N_9597);
or U11145 (N_11145,N_9072,N_8621);
nor U11146 (N_11146,N_9475,N_8991);
xor U11147 (N_11147,N_7557,N_8097);
nor U11148 (N_11148,N_8299,N_8593);
xnor U11149 (N_11149,N_9446,N_9715);
or U11150 (N_11150,N_8877,N_7629);
nor U11151 (N_11151,N_8853,N_8693);
nor U11152 (N_11152,N_9206,N_9014);
xnor U11153 (N_11153,N_8038,N_9860);
and U11154 (N_11154,N_8913,N_8387);
and U11155 (N_11155,N_7934,N_9629);
xor U11156 (N_11156,N_8598,N_9795);
and U11157 (N_11157,N_9541,N_8120);
nand U11158 (N_11158,N_8467,N_8496);
or U11159 (N_11159,N_8127,N_8348);
or U11160 (N_11160,N_9760,N_9870);
or U11161 (N_11161,N_9787,N_7958);
nor U11162 (N_11162,N_7869,N_8160);
nand U11163 (N_11163,N_9493,N_9110);
xnor U11164 (N_11164,N_8402,N_8409);
nand U11165 (N_11165,N_9261,N_7975);
xnor U11166 (N_11166,N_8580,N_8377);
nand U11167 (N_11167,N_8633,N_9203);
or U11168 (N_11168,N_9378,N_9555);
or U11169 (N_11169,N_9635,N_9281);
xor U11170 (N_11170,N_8752,N_9731);
or U11171 (N_11171,N_9642,N_8842);
nor U11172 (N_11172,N_8896,N_7545);
or U11173 (N_11173,N_8982,N_8479);
xnor U11174 (N_11174,N_7572,N_8710);
xor U11175 (N_11175,N_9822,N_8189);
xor U11176 (N_11176,N_9340,N_9949);
or U11177 (N_11177,N_7754,N_7766);
and U11178 (N_11178,N_8717,N_8297);
or U11179 (N_11179,N_9862,N_9291);
nand U11180 (N_11180,N_9290,N_9129);
and U11181 (N_11181,N_8021,N_7550);
xnor U11182 (N_11182,N_8228,N_9607);
or U11183 (N_11183,N_8573,N_9452);
nand U11184 (N_11184,N_9310,N_8086);
xor U11185 (N_11185,N_9123,N_9858);
nor U11186 (N_11186,N_9785,N_8901);
and U11187 (N_11187,N_8109,N_9192);
xor U11188 (N_11188,N_7887,N_8759);
nand U11189 (N_11189,N_7805,N_8229);
xor U11190 (N_11190,N_8941,N_7647);
xor U11191 (N_11191,N_9430,N_9505);
or U11192 (N_11192,N_9622,N_9324);
nor U11193 (N_11193,N_7515,N_8534);
or U11194 (N_11194,N_8635,N_7666);
or U11195 (N_11195,N_8834,N_8609);
nand U11196 (N_11196,N_9626,N_8647);
or U11197 (N_11197,N_8121,N_9532);
or U11198 (N_11198,N_9083,N_9359);
nand U11199 (N_11199,N_8200,N_8388);
or U11200 (N_11200,N_8510,N_9918);
nor U11201 (N_11201,N_8856,N_8326);
and U11202 (N_11202,N_9048,N_7983);
and U11203 (N_11203,N_9095,N_7611);
and U11204 (N_11204,N_9330,N_9305);
xor U11205 (N_11205,N_8688,N_9207);
or U11206 (N_11206,N_9082,N_9654);
and U11207 (N_11207,N_9578,N_8314);
nand U11208 (N_11208,N_8495,N_8426);
nand U11209 (N_11209,N_7985,N_8438);
nand U11210 (N_11210,N_9667,N_9569);
xor U11211 (N_11211,N_7714,N_9363);
and U11212 (N_11212,N_7562,N_9978);
nor U11213 (N_11213,N_8519,N_9616);
nand U11214 (N_11214,N_8381,N_8803);
nand U11215 (N_11215,N_8530,N_7660);
nand U11216 (N_11216,N_8671,N_8078);
xnor U11217 (N_11217,N_8177,N_8133);
and U11218 (N_11218,N_7785,N_8554);
and U11219 (N_11219,N_9623,N_8605);
or U11220 (N_11220,N_9176,N_9387);
xor U11221 (N_11221,N_7911,N_9598);
and U11222 (N_11222,N_7576,N_8236);
nand U11223 (N_11223,N_9088,N_7922);
or U11224 (N_11224,N_9880,N_8713);
or U11225 (N_11225,N_9706,N_8174);
and U11226 (N_11226,N_7744,N_9249);
nor U11227 (N_11227,N_9105,N_8191);
xnor U11228 (N_11228,N_7729,N_8705);
and U11229 (N_11229,N_9081,N_9516);
and U11230 (N_11230,N_9652,N_8862);
xnor U11231 (N_11231,N_8594,N_8320);
or U11232 (N_11232,N_7931,N_9400);
nand U11233 (N_11233,N_8224,N_7826);
and U11234 (N_11234,N_7950,N_8005);
nand U11235 (N_11235,N_8920,N_9492);
nor U11236 (N_11236,N_8085,N_9238);
nand U11237 (N_11237,N_9303,N_9389);
and U11238 (N_11238,N_7741,N_8777);
nand U11239 (N_11239,N_8768,N_8511);
xnor U11240 (N_11240,N_9242,N_9211);
nor U11241 (N_11241,N_7857,N_8098);
and U11242 (N_11242,N_9109,N_9943);
nand U11243 (N_11243,N_8351,N_9570);
nand U11244 (N_11244,N_8395,N_7760);
or U11245 (N_11245,N_8407,N_7638);
nor U11246 (N_11246,N_9719,N_7919);
and U11247 (N_11247,N_8602,N_7553);
xor U11248 (N_11248,N_9030,N_8319);
nand U11249 (N_11249,N_8831,N_9102);
xnor U11250 (N_11250,N_9795,N_8387);
and U11251 (N_11251,N_9014,N_8065);
or U11252 (N_11252,N_9031,N_7671);
and U11253 (N_11253,N_7695,N_7960);
and U11254 (N_11254,N_9716,N_9496);
xnor U11255 (N_11255,N_7565,N_7623);
and U11256 (N_11256,N_8001,N_9615);
nor U11257 (N_11257,N_9351,N_8973);
xor U11258 (N_11258,N_8446,N_8841);
xor U11259 (N_11259,N_9408,N_7679);
nand U11260 (N_11260,N_9741,N_7867);
xor U11261 (N_11261,N_8186,N_8685);
and U11262 (N_11262,N_8652,N_8577);
nand U11263 (N_11263,N_9626,N_8355);
nor U11264 (N_11264,N_9575,N_9027);
nand U11265 (N_11265,N_8666,N_7773);
or U11266 (N_11266,N_8513,N_9398);
nand U11267 (N_11267,N_7761,N_9937);
nand U11268 (N_11268,N_8978,N_8640);
and U11269 (N_11269,N_7830,N_7639);
nor U11270 (N_11270,N_9208,N_8093);
and U11271 (N_11271,N_8458,N_8767);
or U11272 (N_11272,N_7837,N_9198);
or U11273 (N_11273,N_8120,N_8332);
and U11274 (N_11274,N_8990,N_7675);
nand U11275 (N_11275,N_9258,N_9494);
xor U11276 (N_11276,N_9942,N_8870);
nand U11277 (N_11277,N_9224,N_8471);
nand U11278 (N_11278,N_8780,N_9731);
nor U11279 (N_11279,N_8055,N_8214);
or U11280 (N_11280,N_7691,N_9902);
nand U11281 (N_11281,N_9404,N_9527);
nand U11282 (N_11282,N_8160,N_9413);
or U11283 (N_11283,N_8079,N_8154);
nor U11284 (N_11284,N_9076,N_9996);
or U11285 (N_11285,N_9547,N_9461);
and U11286 (N_11286,N_8051,N_7558);
and U11287 (N_11287,N_9073,N_9542);
xnor U11288 (N_11288,N_9716,N_7618);
xnor U11289 (N_11289,N_8072,N_8877);
nor U11290 (N_11290,N_8987,N_9610);
and U11291 (N_11291,N_8570,N_7873);
nand U11292 (N_11292,N_8788,N_8875);
nand U11293 (N_11293,N_8632,N_8391);
nor U11294 (N_11294,N_8021,N_8017);
nand U11295 (N_11295,N_9354,N_8084);
xor U11296 (N_11296,N_9637,N_7879);
nor U11297 (N_11297,N_7632,N_8005);
and U11298 (N_11298,N_8864,N_8872);
or U11299 (N_11299,N_9429,N_7576);
nor U11300 (N_11300,N_9181,N_8362);
nor U11301 (N_11301,N_9478,N_8417);
or U11302 (N_11302,N_9344,N_7954);
nor U11303 (N_11303,N_9626,N_9172);
xnor U11304 (N_11304,N_8061,N_8172);
and U11305 (N_11305,N_7547,N_8235);
and U11306 (N_11306,N_8766,N_9276);
nand U11307 (N_11307,N_9871,N_8610);
and U11308 (N_11308,N_8977,N_8677);
and U11309 (N_11309,N_8386,N_7831);
nand U11310 (N_11310,N_9755,N_9013);
xnor U11311 (N_11311,N_8084,N_9138);
nor U11312 (N_11312,N_9264,N_9656);
xnor U11313 (N_11313,N_8652,N_8683);
xnor U11314 (N_11314,N_7510,N_8782);
and U11315 (N_11315,N_7736,N_9174);
xor U11316 (N_11316,N_8353,N_9707);
or U11317 (N_11317,N_8191,N_7745);
nor U11318 (N_11318,N_9450,N_9826);
nand U11319 (N_11319,N_8081,N_9450);
nand U11320 (N_11320,N_7552,N_8366);
or U11321 (N_11321,N_8066,N_9388);
nand U11322 (N_11322,N_8463,N_9509);
xnor U11323 (N_11323,N_8465,N_8598);
and U11324 (N_11324,N_9780,N_8424);
nor U11325 (N_11325,N_8248,N_9942);
xnor U11326 (N_11326,N_9532,N_9952);
and U11327 (N_11327,N_8475,N_7549);
nand U11328 (N_11328,N_7531,N_8992);
or U11329 (N_11329,N_9865,N_9884);
and U11330 (N_11330,N_8998,N_7699);
nor U11331 (N_11331,N_8924,N_9055);
nor U11332 (N_11332,N_8750,N_9908);
and U11333 (N_11333,N_7774,N_8398);
xor U11334 (N_11334,N_9716,N_9808);
nand U11335 (N_11335,N_9618,N_8467);
xor U11336 (N_11336,N_7914,N_9043);
or U11337 (N_11337,N_8410,N_8025);
xnor U11338 (N_11338,N_7614,N_7584);
nand U11339 (N_11339,N_9195,N_8938);
nand U11340 (N_11340,N_7886,N_8010);
and U11341 (N_11341,N_8637,N_9608);
xor U11342 (N_11342,N_8675,N_8275);
xor U11343 (N_11343,N_9731,N_9835);
xnor U11344 (N_11344,N_8910,N_9329);
nor U11345 (N_11345,N_8179,N_8541);
nand U11346 (N_11346,N_9404,N_8919);
or U11347 (N_11347,N_9496,N_9900);
nor U11348 (N_11348,N_9481,N_9623);
xor U11349 (N_11349,N_9649,N_9713);
and U11350 (N_11350,N_8245,N_7674);
xor U11351 (N_11351,N_8810,N_9445);
nor U11352 (N_11352,N_9272,N_8299);
nand U11353 (N_11353,N_9673,N_7587);
nand U11354 (N_11354,N_8957,N_9503);
or U11355 (N_11355,N_7823,N_7837);
xnor U11356 (N_11356,N_8837,N_7941);
nand U11357 (N_11357,N_8346,N_9989);
xnor U11358 (N_11358,N_9889,N_9302);
or U11359 (N_11359,N_8885,N_8368);
and U11360 (N_11360,N_8739,N_8850);
nand U11361 (N_11361,N_8283,N_8366);
and U11362 (N_11362,N_7608,N_9232);
nand U11363 (N_11363,N_8123,N_8331);
nor U11364 (N_11364,N_8801,N_8398);
nor U11365 (N_11365,N_8348,N_9360);
nor U11366 (N_11366,N_8702,N_7669);
nand U11367 (N_11367,N_9558,N_9749);
xnor U11368 (N_11368,N_7881,N_8609);
or U11369 (N_11369,N_8752,N_7548);
nor U11370 (N_11370,N_8881,N_7508);
and U11371 (N_11371,N_8258,N_9834);
xor U11372 (N_11372,N_8280,N_9299);
and U11373 (N_11373,N_9520,N_7610);
or U11374 (N_11374,N_8082,N_9206);
or U11375 (N_11375,N_9085,N_8833);
xnor U11376 (N_11376,N_9369,N_8251);
nand U11377 (N_11377,N_8164,N_9548);
nand U11378 (N_11378,N_9361,N_8672);
and U11379 (N_11379,N_9964,N_8172);
nand U11380 (N_11380,N_8227,N_9326);
or U11381 (N_11381,N_8936,N_9394);
nor U11382 (N_11382,N_8519,N_8150);
nor U11383 (N_11383,N_8639,N_7825);
or U11384 (N_11384,N_8055,N_7553);
nor U11385 (N_11385,N_7660,N_8007);
and U11386 (N_11386,N_8538,N_9545);
and U11387 (N_11387,N_9469,N_8795);
nand U11388 (N_11388,N_8313,N_9144);
xor U11389 (N_11389,N_8122,N_8408);
or U11390 (N_11390,N_9814,N_9587);
and U11391 (N_11391,N_9209,N_8121);
xor U11392 (N_11392,N_7781,N_8958);
or U11393 (N_11393,N_9115,N_8004);
nor U11394 (N_11394,N_9262,N_8470);
nand U11395 (N_11395,N_8286,N_8651);
xor U11396 (N_11396,N_8677,N_9053);
and U11397 (N_11397,N_9784,N_9066);
xnor U11398 (N_11398,N_8730,N_7536);
or U11399 (N_11399,N_8384,N_8535);
or U11400 (N_11400,N_9237,N_9633);
xnor U11401 (N_11401,N_8339,N_7750);
nor U11402 (N_11402,N_9995,N_8233);
nand U11403 (N_11403,N_9719,N_8875);
nand U11404 (N_11404,N_8516,N_8079);
nor U11405 (N_11405,N_9848,N_8603);
and U11406 (N_11406,N_7831,N_9981);
nand U11407 (N_11407,N_7979,N_9340);
nand U11408 (N_11408,N_8718,N_7581);
nand U11409 (N_11409,N_9720,N_7783);
nand U11410 (N_11410,N_9423,N_8557);
xor U11411 (N_11411,N_8903,N_9839);
and U11412 (N_11412,N_9168,N_9117);
nand U11413 (N_11413,N_8790,N_9793);
xnor U11414 (N_11414,N_9151,N_7836);
nand U11415 (N_11415,N_9583,N_9156);
nor U11416 (N_11416,N_7899,N_9549);
nand U11417 (N_11417,N_7806,N_9133);
or U11418 (N_11418,N_9829,N_9923);
xor U11419 (N_11419,N_7913,N_8835);
nand U11420 (N_11420,N_9766,N_9578);
xor U11421 (N_11421,N_9786,N_9116);
or U11422 (N_11422,N_7928,N_8204);
nand U11423 (N_11423,N_8027,N_9285);
nor U11424 (N_11424,N_7971,N_7545);
and U11425 (N_11425,N_8159,N_8188);
or U11426 (N_11426,N_7842,N_8478);
nand U11427 (N_11427,N_9706,N_8226);
or U11428 (N_11428,N_7757,N_8762);
or U11429 (N_11429,N_8109,N_9222);
xor U11430 (N_11430,N_9703,N_9228);
xor U11431 (N_11431,N_9461,N_8535);
nand U11432 (N_11432,N_7902,N_8676);
and U11433 (N_11433,N_8392,N_8327);
and U11434 (N_11434,N_9602,N_7750);
and U11435 (N_11435,N_9932,N_8319);
nand U11436 (N_11436,N_9687,N_9229);
xnor U11437 (N_11437,N_8644,N_9736);
and U11438 (N_11438,N_9387,N_9567);
or U11439 (N_11439,N_9293,N_9449);
nor U11440 (N_11440,N_9870,N_8439);
xnor U11441 (N_11441,N_8515,N_9319);
nor U11442 (N_11442,N_9247,N_7507);
and U11443 (N_11443,N_8284,N_7610);
or U11444 (N_11444,N_9184,N_9705);
xnor U11445 (N_11445,N_7869,N_8181);
or U11446 (N_11446,N_8462,N_8375);
nor U11447 (N_11447,N_8447,N_9095);
nor U11448 (N_11448,N_9122,N_9156);
and U11449 (N_11449,N_9089,N_9747);
or U11450 (N_11450,N_7987,N_9277);
and U11451 (N_11451,N_7662,N_9982);
nor U11452 (N_11452,N_9899,N_8951);
or U11453 (N_11453,N_8048,N_7560);
and U11454 (N_11454,N_7886,N_9003);
nand U11455 (N_11455,N_9507,N_8558);
nand U11456 (N_11456,N_8934,N_7705);
nand U11457 (N_11457,N_9416,N_7953);
nor U11458 (N_11458,N_9152,N_9585);
and U11459 (N_11459,N_9998,N_9119);
nor U11460 (N_11460,N_8344,N_9631);
nand U11461 (N_11461,N_7924,N_9432);
and U11462 (N_11462,N_9957,N_9375);
and U11463 (N_11463,N_8546,N_7841);
xor U11464 (N_11464,N_8609,N_9419);
nor U11465 (N_11465,N_7757,N_9693);
nor U11466 (N_11466,N_8833,N_9862);
and U11467 (N_11467,N_9638,N_9239);
or U11468 (N_11468,N_7875,N_8690);
nand U11469 (N_11469,N_8504,N_8320);
nand U11470 (N_11470,N_9487,N_8051);
and U11471 (N_11471,N_9630,N_8565);
nand U11472 (N_11472,N_7921,N_8683);
nand U11473 (N_11473,N_8315,N_8051);
or U11474 (N_11474,N_8971,N_9191);
and U11475 (N_11475,N_9389,N_8275);
and U11476 (N_11476,N_9949,N_7778);
nor U11477 (N_11477,N_7876,N_9471);
or U11478 (N_11478,N_9041,N_9014);
nand U11479 (N_11479,N_8075,N_7643);
nand U11480 (N_11480,N_7653,N_9684);
or U11481 (N_11481,N_7636,N_8001);
nor U11482 (N_11482,N_9580,N_9091);
nor U11483 (N_11483,N_7897,N_8618);
xor U11484 (N_11484,N_8009,N_8929);
nand U11485 (N_11485,N_9142,N_8983);
nand U11486 (N_11486,N_8656,N_9311);
nand U11487 (N_11487,N_9474,N_7529);
and U11488 (N_11488,N_7812,N_9795);
or U11489 (N_11489,N_8616,N_9828);
nand U11490 (N_11490,N_8812,N_9934);
or U11491 (N_11491,N_8134,N_9777);
and U11492 (N_11492,N_9711,N_9128);
xnor U11493 (N_11493,N_8160,N_9520);
xnor U11494 (N_11494,N_9899,N_7968);
nor U11495 (N_11495,N_8127,N_9452);
xnor U11496 (N_11496,N_9557,N_9239);
xor U11497 (N_11497,N_9179,N_9797);
nand U11498 (N_11498,N_9690,N_9514);
or U11499 (N_11499,N_8547,N_8112);
xnor U11500 (N_11500,N_7824,N_9715);
nand U11501 (N_11501,N_9299,N_8987);
nor U11502 (N_11502,N_8608,N_8563);
or U11503 (N_11503,N_7903,N_7688);
and U11504 (N_11504,N_8705,N_7631);
nor U11505 (N_11505,N_7547,N_8316);
and U11506 (N_11506,N_7987,N_9140);
or U11507 (N_11507,N_8271,N_7725);
xor U11508 (N_11508,N_8156,N_9287);
and U11509 (N_11509,N_8611,N_8600);
nand U11510 (N_11510,N_9829,N_8227);
nand U11511 (N_11511,N_9527,N_9604);
nor U11512 (N_11512,N_9382,N_8097);
nor U11513 (N_11513,N_9599,N_9841);
and U11514 (N_11514,N_8959,N_7650);
or U11515 (N_11515,N_9961,N_9691);
or U11516 (N_11516,N_8235,N_8341);
nor U11517 (N_11517,N_8874,N_9901);
and U11518 (N_11518,N_8180,N_8102);
nand U11519 (N_11519,N_9727,N_9739);
xor U11520 (N_11520,N_9065,N_8866);
xor U11521 (N_11521,N_8643,N_9914);
nor U11522 (N_11522,N_9020,N_9916);
nor U11523 (N_11523,N_8430,N_9704);
nor U11524 (N_11524,N_9357,N_8515);
and U11525 (N_11525,N_9232,N_8822);
or U11526 (N_11526,N_9750,N_8633);
nand U11527 (N_11527,N_9256,N_8094);
nor U11528 (N_11528,N_8760,N_7638);
and U11529 (N_11529,N_8901,N_8173);
or U11530 (N_11530,N_9791,N_8672);
nand U11531 (N_11531,N_9883,N_8042);
and U11532 (N_11532,N_8988,N_8698);
nor U11533 (N_11533,N_9308,N_7519);
and U11534 (N_11534,N_8742,N_9218);
nor U11535 (N_11535,N_7664,N_8999);
nor U11536 (N_11536,N_8789,N_9706);
xor U11537 (N_11537,N_8434,N_8389);
xor U11538 (N_11538,N_9511,N_9013);
and U11539 (N_11539,N_9018,N_8656);
or U11540 (N_11540,N_9722,N_9860);
xor U11541 (N_11541,N_8761,N_7542);
and U11542 (N_11542,N_8347,N_9401);
xor U11543 (N_11543,N_7998,N_9472);
xnor U11544 (N_11544,N_8688,N_9086);
nand U11545 (N_11545,N_8516,N_8181);
nor U11546 (N_11546,N_7834,N_8462);
nor U11547 (N_11547,N_8471,N_7823);
or U11548 (N_11548,N_9693,N_7530);
nor U11549 (N_11549,N_8481,N_9361);
nand U11550 (N_11550,N_8648,N_9702);
and U11551 (N_11551,N_8935,N_8736);
and U11552 (N_11552,N_7935,N_9208);
nor U11553 (N_11553,N_7998,N_7647);
and U11554 (N_11554,N_9092,N_8591);
and U11555 (N_11555,N_8732,N_9275);
nand U11556 (N_11556,N_9524,N_9839);
nand U11557 (N_11557,N_7815,N_8354);
nor U11558 (N_11558,N_8122,N_7960);
nand U11559 (N_11559,N_7650,N_8357);
nand U11560 (N_11560,N_8969,N_8879);
nand U11561 (N_11561,N_9454,N_8733);
or U11562 (N_11562,N_7616,N_9903);
nand U11563 (N_11563,N_8712,N_8292);
nand U11564 (N_11564,N_9342,N_9963);
nand U11565 (N_11565,N_8591,N_9701);
or U11566 (N_11566,N_9619,N_9547);
nor U11567 (N_11567,N_7914,N_7735);
nor U11568 (N_11568,N_7776,N_8163);
and U11569 (N_11569,N_8440,N_8513);
nor U11570 (N_11570,N_8883,N_9455);
nor U11571 (N_11571,N_8533,N_8670);
xor U11572 (N_11572,N_9927,N_7844);
xor U11573 (N_11573,N_8316,N_8381);
or U11574 (N_11574,N_7895,N_7968);
xor U11575 (N_11575,N_8958,N_8028);
and U11576 (N_11576,N_7733,N_8926);
and U11577 (N_11577,N_8910,N_7527);
nand U11578 (N_11578,N_9626,N_9086);
or U11579 (N_11579,N_9356,N_8768);
nor U11580 (N_11580,N_8092,N_8228);
xnor U11581 (N_11581,N_9230,N_8843);
nand U11582 (N_11582,N_9178,N_8864);
and U11583 (N_11583,N_7946,N_9906);
nand U11584 (N_11584,N_8181,N_8565);
xnor U11585 (N_11585,N_8966,N_8722);
nor U11586 (N_11586,N_9079,N_8680);
nand U11587 (N_11587,N_9384,N_8943);
or U11588 (N_11588,N_8479,N_8078);
or U11589 (N_11589,N_9175,N_9614);
nand U11590 (N_11590,N_9694,N_8158);
or U11591 (N_11591,N_9626,N_8754);
nand U11592 (N_11592,N_8409,N_8030);
or U11593 (N_11593,N_7954,N_8361);
or U11594 (N_11594,N_7891,N_9826);
or U11595 (N_11595,N_8352,N_7665);
nand U11596 (N_11596,N_7608,N_8448);
and U11597 (N_11597,N_8518,N_9130);
xor U11598 (N_11598,N_9852,N_8700);
nand U11599 (N_11599,N_9672,N_8352);
nand U11600 (N_11600,N_8466,N_9221);
and U11601 (N_11601,N_7762,N_7552);
xor U11602 (N_11602,N_9006,N_8470);
or U11603 (N_11603,N_9089,N_9134);
and U11604 (N_11604,N_9661,N_8518);
nor U11605 (N_11605,N_9847,N_9768);
nor U11606 (N_11606,N_8006,N_9191);
nor U11607 (N_11607,N_9788,N_8687);
xor U11608 (N_11608,N_9359,N_8036);
nand U11609 (N_11609,N_7694,N_7994);
and U11610 (N_11610,N_9506,N_9409);
nor U11611 (N_11611,N_8006,N_7620);
nor U11612 (N_11612,N_7599,N_9429);
xnor U11613 (N_11613,N_7970,N_8367);
or U11614 (N_11614,N_8864,N_8416);
or U11615 (N_11615,N_9121,N_9941);
nor U11616 (N_11616,N_9291,N_9648);
or U11617 (N_11617,N_9617,N_7540);
and U11618 (N_11618,N_9708,N_9802);
nor U11619 (N_11619,N_9250,N_9153);
nor U11620 (N_11620,N_7542,N_8866);
nand U11621 (N_11621,N_7567,N_8739);
nand U11622 (N_11622,N_9944,N_9245);
or U11623 (N_11623,N_8412,N_8477);
nand U11624 (N_11624,N_9412,N_8779);
xor U11625 (N_11625,N_8894,N_8383);
and U11626 (N_11626,N_9585,N_9053);
nand U11627 (N_11627,N_9725,N_8464);
or U11628 (N_11628,N_8491,N_9488);
nor U11629 (N_11629,N_8711,N_8853);
nor U11630 (N_11630,N_8415,N_7552);
or U11631 (N_11631,N_7531,N_8436);
nor U11632 (N_11632,N_8900,N_9193);
xor U11633 (N_11633,N_7826,N_8584);
and U11634 (N_11634,N_8618,N_8336);
nor U11635 (N_11635,N_7653,N_7828);
nor U11636 (N_11636,N_8541,N_9659);
nand U11637 (N_11637,N_7883,N_9303);
nand U11638 (N_11638,N_8140,N_7566);
nor U11639 (N_11639,N_8658,N_7529);
xor U11640 (N_11640,N_7883,N_9733);
and U11641 (N_11641,N_8020,N_7634);
and U11642 (N_11642,N_9265,N_9173);
or U11643 (N_11643,N_7549,N_9570);
or U11644 (N_11644,N_8600,N_9662);
xnor U11645 (N_11645,N_7736,N_8177);
xor U11646 (N_11646,N_8048,N_9743);
nor U11647 (N_11647,N_9045,N_9948);
and U11648 (N_11648,N_9890,N_8072);
or U11649 (N_11649,N_8395,N_8380);
nand U11650 (N_11650,N_8906,N_8813);
nand U11651 (N_11651,N_9086,N_8840);
xnor U11652 (N_11652,N_9648,N_8455);
and U11653 (N_11653,N_7725,N_8415);
nor U11654 (N_11654,N_8586,N_8394);
nand U11655 (N_11655,N_9622,N_8497);
and U11656 (N_11656,N_9326,N_9471);
or U11657 (N_11657,N_8753,N_8060);
nand U11658 (N_11658,N_7547,N_8425);
xnor U11659 (N_11659,N_9315,N_9820);
xnor U11660 (N_11660,N_8177,N_7584);
xor U11661 (N_11661,N_9299,N_8638);
or U11662 (N_11662,N_8943,N_9554);
and U11663 (N_11663,N_8309,N_8409);
and U11664 (N_11664,N_8337,N_9376);
xnor U11665 (N_11665,N_9654,N_8489);
xor U11666 (N_11666,N_7803,N_8884);
nor U11667 (N_11667,N_7660,N_9376);
nand U11668 (N_11668,N_7747,N_8421);
nor U11669 (N_11669,N_8987,N_8309);
nor U11670 (N_11670,N_8895,N_8509);
nand U11671 (N_11671,N_9286,N_8718);
nor U11672 (N_11672,N_8155,N_9203);
and U11673 (N_11673,N_7899,N_9570);
or U11674 (N_11674,N_8565,N_8683);
nand U11675 (N_11675,N_8022,N_8164);
or U11676 (N_11676,N_9244,N_9827);
or U11677 (N_11677,N_8619,N_7611);
and U11678 (N_11678,N_9274,N_8413);
and U11679 (N_11679,N_7858,N_9507);
xnor U11680 (N_11680,N_8825,N_9175);
xor U11681 (N_11681,N_9904,N_7715);
and U11682 (N_11682,N_9694,N_9761);
nand U11683 (N_11683,N_7646,N_9881);
and U11684 (N_11684,N_8095,N_9189);
and U11685 (N_11685,N_9606,N_7793);
or U11686 (N_11686,N_7653,N_8646);
and U11687 (N_11687,N_9237,N_8250);
nand U11688 (N_11688,N_9437,N_7853);
xnor U11689 (N_11689,N_9647,N_9681);
nand U11690 (N_11690,N_8245,N_8410);
nand U11691 (N_11691,N_8230,N_9161);
nor U11692 (N_11692,N_9370,N_8260);
nand U11693 (N_11693,N_7893,N_7708);
xor U11694 (N_11694,N_8710,N_8526);
and U11695 (N_11695,N_9674,N_8041);
and U11696 (N_11696,N_9368,N_8171);
nor U11697 (N_11697,N_7972,N_9721);
xor U11698 (N_11698,N_9524,N_8449);
and U11699 (N_11699,N_7951,N_8910);
xor U11700 (N_11700,N_9704,N_8456);
xnor U11701 (N_11701,N_9894,N_7710);
and U11702 (N_11702,N_8927,N_9093);
and U11703 (N_11703,N_7819,N_7587);
and U11704 (N_11704,N_8445,N_9158);
nor U11705 (N_11705,N_8213,N_9165);
nor U11706 (N_11706,N_7902,N_8768);
or U11707 (N_11707,N_9557,N_8910);
and U11708 (N_11708,N_8668,N_8388);
nand U11709 (N_11709,N_8752,N_9541);
nor U11710 (N_11710,N_8613,N_8675);
and U11711 (N_11711,N_7936,N_8589);
or U11712 (N_11712,N_8088,N_8831);
and U11713 (N_11713,N_8482,N_9836);
nand U11714 (N_11714,N_8672,N_7947);
and U11715 (N_11715,N_9015,N_9354);
xnor U11716 (N_11716,N_9527,N_8376);
nand U11717 (N_11717,N_8309,N_7574);
and U11718 (N_11718,N_8418,N_9874);
and U11719 (N_11719,N_8407,N_9789);
xnor U11720 (N_11720,N_9654,N_7501);
xor U11721 (N_11721,N_9885,N_7815);
and U11722 (N_11722,N_9408,N_8126);
nand U11723 (N_11723,N_9102,N_8265);
nor U11724 (N_11724,N_8506,N_8684);
nand U11725 (N_11725,N_9537,N_9171);
nand U11726 (N_11726,N_8593,N_8394);
and U11727 (N_11727,N_7963,N_9624);
nand U11728 (N_11728,N_9489,N_8277);
nand U11729 (N_11729,N_7887,N_7675);
nand U11730 (N_11730,N_7775,N_7750);
nand U11731 (N_11731,N_9327,N_7768);
nor U11732 (N_11732,N_9758,N_8805);
or U11733 (N_11733,N_8894,N_8235);
or U11734 (N_11734,N_9034,N_8162);
or U11735 (N_11735,N_8057,N_7854);
nor U11736 (N_11736,N_9440,N_9083);
nor U11737 (N_11737,N_8491,N_9076);
and U11738 (N_11738,N_9937,N_7656);
xnor U11739 (N_11739,N_8517,N_8427);
nand U11740 (N_11740,N_9793,N_9398);
nand U11741 (N_11741,N_7769,N_8291);
and U11742 (N_11742,N_8463,N_9393);
or U11743 (N_11743,N_8133,N_8198);
and U11744 (N_11744,N_9322,N_7908);
nand U11745 (N_11745,N_9051,N_8305);
nor U11746 (N_11746,N_9559,N_9501);
or U11747 (N_11747,N_9746,N_8317);
nor U11748 (N_11748,N_7690,N_9372);
or U11749 (N_11749,N_8513,N_9239);
nor U11750 (N_11750,N_9152,N_8392);
nor U11751 (N_11751,N_9491,N_8746);
nor U11752 (N_11752,N_8541,N_9513);
nor U11753 (N_11753,N_8857,N_9433);
xor U11754 (N_11754,N_8578,N_7676);
and U11755 (N_11755,N_7705,N_8872);
and U11756 (N_11756,N_7666,N_7917);
nand U11757 (N_11757,N_9704,N_7515);
or U11758 (N_11758,N_7970,N_7874);
and U11759 (N_11759,N_8432,N_8775);
nand U11760 (N_11760,N_9704,N_7765);
and U11761 (N_11761,N_8971,N_7938);
xor U11762 (N_11762,N_8165,N_8320);
and U11763 (N_11763,N_8201,N_9690);
nor U11764 (N_11764,N_7552,N_8897);
nor U11765 (N_11765,N_9992,N_8021);
xor U11766 (N_11766,N_8684,N_8554);
and U11767 (N_11767,N_9884,N_9778);
xor U11768 (N_11768,N_9095,N_9864);
and U11769 (N_11769,N_9518,N_7951);
or U11770 (N_11770,N_9973,N_8750);
or U11771 (N_11771,N_8966,N_8380);
and U11772 (N_11772,N_8110,N_7714);
nand U11773 (N_11773,N_9498,N_9380);
or U11774 (N_11774,N_9950,N_8319);
or U11775 (N_11775,N_8429,N_9874);
and U11776 (N_11776,N_7757,N_9778);
nand U11777 (N_11777,N_7756,N_7775);
and U11778 (N_11778,N_8894,N_8367);
xor U11779 (N_11779,N_8234,N_9943);
or U11780 (N_11780,N_8948,N_8191);
xnor U11781 (N_11781,N_9439,N_8596);
or U11782 (N_11782,N_9894,N_9902);
nor U11783 (N_11783,N_9749,N_7889);
or U11784 (N_11784,N_7810,N_9621);
nand U11785 (N_11785,N_9803,N_9176);
nand U11786 (N_11786,N_8341,N_8759);
and U11787 (N_11787,N_8585,N_7543);
nor U11788 (N_11788,N_7577,N_9410);
xor U11789 (N_11789,N_7591,N_9703);
nand U11790 (N_11790,N_9187,N_8101);
xor U11791 (N_11791,N_9198,N_9316);
or U11792 (N_11792,N_9957,N_8463);
and U11793 (N_11793,N_9605,N_8035);
nand U11794 (N_11794,N_9596,N_8972);
nand U11795 (N_11795,N_7645,N_9944);
xnor U11796 (N_11796,N_9096,N_8119);
nand U11797 (N_11797,N_8410,N_9706);
or U11798 (N_11798,N_8785,N_7639);
nand U11799 (N_11799,N_7990,N_7626);
and U11800 (N_11800,N_7760,N_9461);
xor U11801 (N_11801,N_8761,N_9438);
or U11802 (N_11802,N_8144,N_7964);
or U11803 (N_11803,N_9668,N_8741);
and U11804 (N_11804,N_9511,N_8816);
xor U11805 (N_11805,N_8168,N_7899);
nor U11806 (N_11806,N_9631,N_7836);
xnor U11807 (N_11807,N_9056,N_8351);
nand U11808 (N_11808,N_9276,N_9772);
nand U11809 (N_11809,N_7813,N_9897);
or U11810 (N_11810,N_8152,N_9577);
nand U11811 (N_11811,N_7927,N_7637);
nand U11812 (N_11812,N_9164,N_8827);
and U11813 (N_11813,N_7939,N_8492);
or U11814 (N_11814,N_7969,N_7875);
nor U11815 (N_11815,N_8333,N_8464);
nor U11816 (N_11816,N_8656,N_7743);
or U11817 (N_11817,N_9089,N_9236);
nand U11818 (N_11818,N_7708,N_7901);
nor U11819 (N_11819,N_7610,N_7823);
xor U11820 (N_11820,N_8005,N_9503);
nand U11821 (N_11821,N_9650,N_8285);
nor U11822 (N_11822,N_7569,N_9312);
xnor U11823 (N_11823,N_9727,N_8601);
nor U11824 (N_11824,N_9922,N_8062);
xnor U11825 (N_11825,N_9945,N_9951);
nand U11826 (N_11826,N_9126,N_9574);
xnor U11827 (N_11827,N_8663,N_8082);
nor U11828 (N_11828,N_7574,N_9822);
and U11829 (N_11829,N_7886,N_7785);
or U11830 (N_11830,N_9195,N_9763);
and U11831 (N_11831,N_7946,N_7827);
xor U11832 (N_11832,N_8364,N_7936);
xor U11833 (N_11833,N_8069,N_9300);
xor U11834 (N_11834,N_9819,N_9748);
nand U11835 (N_11835,N_7670,N_9678);
and U11836 (N_11836,N_7648,N_8376);
xor U11837 (N_11837,N_9825,N_8511);
and U11838 (N_11838,N_8889,N_7701);
and U11839 (N_11839,N_8315,N_9675);
and U11840 (N_11840,N_7914,N_8909);
nand U11841 (N_11841,N_8860,N_8207);
nand U11842 (N_11842,N_7614,N_8127);
xnor U11843 (N_11843,N_9298,N_9396);
nand U11844 (N_11844,N_8833,N_8476);
or U11845 (N_11845,N_8324,N_9725);
nor U11846 (N_11846,N_9371,N_7728);
or U11847 (N_11847,N_9044,N_7700);
and U11848 (N_11848,N_9900,N_9204);
nor U11849 (N_11849,N_7697,N_7924);
and U11850 (N_11850,N_8977,N_9914);
nand U11851 (N_11851,N_7628,N_9781);
and U11852 (N_11852,N_8224,N_8821);
and U11853 (N_11853,N_9309,N_9065);
and U11854 (N_11854,N_8370,N_8504);
xnor U11855 (N_11855,N_9774,N_9081);
and U11856 (N_11856,N_8467,N_9666);
xnor U11857 (N_11857,N_9874,N_8391);
xor U11858 (N_11858,N_8991,N_9403);
and U11859 (N_11859,N_9309,N_7545);
or U11860 (N_11860,N_8498,N_9157);
and U11861 (N_11861,N_7834,N_9782);
nor U11862 (N_11862,N_7674,N_9619);
and U11863 (N_11863,N_9114,N_8382);
or U11864 (N_11864,N_9665,N_8026);
nand U11865 (N_11865,N_9672,N_8966);
and U11866 (N_11866,N_8748,N_9928);
or U11867 (N_11867,N_7650,N_8623);
and U11868 (N_11868,N_8065,N_8165);
xor U11869 (N_11869,N_8645,N_8753);
xor U11870 (N_11870,N_9866,N_7851);
nand U11871 (N_11871,N_9041,N_8611);
xor U11872 (N_11872,N_7915,N_9294);
nand U11873 (N_11873,N_7899,N_9744);
nor U11874 (N_11874,N_8613,N_8223);
or U11875 (N_11875,N_8939,N_9994);
nor U11876 (N_11876,N_9679,N_9859);
or U11877 (N_11877,N_8432,N_7750);
or U11878 (N_11878,N_8156,N_9626);
or U11879 (N_11879,N_9758,N_8600);
xnor U11880 (N_11880,N_7905,N_9515);
xnor U11881 (N_11881,N_9822,N_7978);
nor U11882 (N_11882,N_7698,N_7738);
nand U11883 (N_11883,N_9282,N_9324);
xnor U11884 (N_11884,N_7920,N_9028);
nand U11885 (N_11885,N_9221,N_8559);
nand U11886 (N_11886,N_7898,N_9985);
xnor U11887 (N_11887,N_8449,N_9865);
nor U11888 (N_11888,N_7916,N_8112);
and U11889 (N_11889,N_8770,N_9924);
nand U11890 (N_11890,N_8500,N_8174);
nand U11891 (N_11891,N_8513,N_8312);
xor U11892 (N_11892,N_9697,N_9836);
nand U11893 (N_11893,N_8478,N_7780);
nor U11894 (N_11894,N_9507,N_9538);
nand U11895 (N_11895,N_7828,N_8765);
nand U11896 (N_11896,N_9537,N_8591);
nand U11897 (N_11897,N_8502,N_7804);
nor U11898 (N_11898,N_7991,N_7968);
or U11899 (N_11899,N_9310,N_8089);
and U11900 (N_11900,N_8183,N_9477);
and U11901 (N_11901,N_8691,N_7651);
or U11902 (N_11902,N_7915,N_9129);
and U11903 (N_11903,N_9684,N_9770);
xnor U11904 (N_11904,N_9019,N_8079);
nor U11905 (N_11905,N_8455,N_9676);
or U11906 (N_11906,N_7610,N_8371);
nand U11907 (N_11907,N_8146,N_8331);
and U11908 (N_11908,N_8813,N_8287);
xnor U11909 (N_11909,N_7886,N_7892);
or U11910 (N_11910,N_8166,N_9236);
nor U11911 (N_11911,N_9279,N_9740);
or U11912 (N_11912,N_8636,N_8254);
xor U11913 (N_11913,N_9265,N_9664);
xor U11914 (N_11914,N_7907,N_8392);
or U11915 (N_11915,N_7597,N_7905);
nor U11916 (N_11916,N_7844,N_8770);
xnor U11917 (N_11917,N_9133,N_9466);
nor U11918 (N_11918,N_8906,N_8525);
or U11919 (N_11919,N_8537,N_8928);
or U11920 (N_11920,N_7627,N_7930);
and U11921 (N_11921,N_8627,N_9983);
nor U11922 (N_11922,N_9832,N_8769);
nor U11923 (N_11923,N_8419,N_8607);
nor U11924 (N_11924,N_7859,N_9154);
nand U11925 (N_11925,N_9223,N_9429);
xnor U11926 (N_11926,N_9995,N_7863);
or U11927 (N_11927,N_9595,N_9709);
nor U11928 (N_11928,N_9704,N_8030);
nor U11929 (N_11929,N_9743,N_9787);
xor U11930 (N_11930,N_9185,N_9731);
and U11931 (N_11931,N_8222,N_9076);
nor U11932 (N_11932,N_7578,N_8945);
xor U11933 (N_11933,N_8883,N_8179);
and U11934 (N_11934,N_8546,N_8972);
nand U11935 (N_11935,N_9368,N_9641);
xnor U11936 (N_11936,N_9565,N_9904);
nand U11937 (N_11937,N_9907,N_7931);
and U11938 (N_11938,N_8670,N_8036);
nand U11939 (N_11939,N_9232,N_8908);
nand U11940 (N_11940,N_7943,N_9109);
nor U11941 (N_11941,N_8211,N_8352);
xor U11942 (N_11942,N_8963,N_8521);
xnor U11943 (N_11943,N_8922,N_7938);
nand U11944 (N_11944,N_8384,N_8913);
and U11945 (N_11945,N_7513,N_8008);
and U11946 (N_11946,N_9916,N_9370);
nand U11947 (N_11947,N_9447,N_8655);
nand U11948 (N_11948,N_8050,N_9544);
and U11949 (N_11949,N_7859,N_8688);
xor U11950 (N_11950,N_9591,N_7583);
or U11951 (N_11951,N_9187,N_9639);
nor U11952 (N_11952,N_8484,N_7979);
nor U11953 (N_11953,N_7741,N_8179);
or U11954 (N_11954,N_7876,N_8696);
and U11955 (N_11955,N_8231,N_9272);
and U11956 (N_11956,N_9066,N_7695);
or U11957 (N_11957,N_7556,N_9310);
and U11958 (N_11958,N_8570,N_8510);
nor U11959 (N_11959,N_8394,N_8902);
xor U11960 (N_11960,N_9476,N_9399);
and U11961 (N_11961,N_7921,N_7731);
xnor U11962 (N_11962,N_8501,N_7843);
nand U11963 (N_11963,N_8022,N_8270);
or U11964 (N_11964,N_7904,N_8055);
nor U11965 (N_11965,N_9223,N_7550);
and U11966 (N_11966,N_9421,N_9299);
nand U11967 (N_11967,N_9512,N_8550);
or U11968 (N_11968,N_9750,N_9700);
nor U11969 (N_11969,N_9451,N_8099);
and U11970 (N_11970,N_7764,N_9426);
or U11971 (N_11971,N_9179,N_8285);
nand U11972 (N_11972,N_8597,N_9446);
nor U11973 (N_11973,N_7764,N_8845);
and U11974 (N_11974,N_9444,N_7712);
nor U11975 (N_11975,N_9617,N_7635);
or U11976 (N_11976,N_9131,N_8229);
nand U11977 (N_11977,N_9728,N_7664);
xor U11978 (N_11978,N_7623,N_9600);
nor U11979 (N_11979,N_7547,N_9725);
or U11980 (N_11980,N_8632,N_7875);
and U11981 (N_11981,N_9270,N_8774);
and U11982 (N_11982,N_9007,N_9602);
xor U11983 (N_11983,N_8616,N_9857);
xor U11984 (N_11984,N_9782,N_7530);
xnor U11985 (N_11985,N_7953,N_9089);
nand U11986 (N_11986,N_8611,N_8787);
nor U11987 (N_11987,N_8427,N_9947);
nor U11988 (N_11988,N_8339,N_9696);
xnor U11989 (N_11989,N_9821,N_8384);
xor U11990 (N_11990,N_7858,N_9076);
and U11991 (N_11991,N_8540,N_7575);
nand U11992 (N_11992,N_9708,N_8403);
and U11993 (N_11993,N_8226,N_9273);
or U11994 (N_11994,N_9106,N_9539);
and U11995 (N_11995,N_8646,N_7746);
xnor U11996 (N_11996,N_7960,N_8947);
or U11997 (N_11997,N_9134,N_9460);
xnor U11998 (N_11998,N_8113,N_8371);
nor U11999 (N_11999,N_8508,N_9577);
or U12000 (N_12000,N_7508,N_9749);
and U12001 (N_12001,N_9316,N_9536);
xor U12002 (N_12002,N_8379,N_9498);
nand U12003 (N_12003,N_8005,N_9449);
nor U12004 (N_12004,N_7854,N_8740);
and U12005 (N_12005,N_8395,N_8489);
nor U12006 (N_12006,N_9349,N_9492);
or U12007 (N_12007,N_8034,N_9894);
nor U12008 (N_12008,N_8472,N_9092);
and U12009 (N_12009,N_9358,N_7508);
nand U12010 (N_12010,N_7820,N_9835);
nand U12011 (N_12011,N_7753,N_9362);
nor U12012 (N_12012,N_8100,N_7933);
nor U12013 (N_12013,N_7631,N_9122);
nor U12014 (N_12014,N_9880,N_9656);
xor U12015 (N_12015,N_9520,N_7937);
nand U12016 (N_12016,N_9258,N_8066);
nor U12017 (N_12017,N_7888,N_9644);
nand U12018 (N_12018,N_9587,N_9532);
nand U12019 (N_12019,N_7761,N_9342);
nand U12020 (N_12020,N_9479,N_9657);
nand U12021 (N_12021,N_8340,N_8495);
xnor U12022 (N_12022,N_9258,N_9199);
nor U12023 (N_12023,N_9098,N_7543);
or U12024 (N_12024,N_9736,N_9236);
nor U12025 (N_12025,N_7541,N_8875);
nor U12026 (N_12026,N_9171,N_7634);
and U12027 (N_12027,N_9167,N_8093);
and U12028 (N_12028,N_7932,N_7953);
nor U12029 (N_12029,N_8288,N_8615);
xnor U12030 (N_12030,N_9128,N_8334);
or U12031 (N_12031,N_9098,N_8124);
nand U12032 (N_12032,N_8924,N_9379);
xor U12033 (N_12033,N_9194,N_7786);
nor U12034 (N_12034,N_8034,N_8732);
or U12035 (N_12035,N_7955,N_8900);
and U12036 (N_12036,N_9772,N_8874);
nor U12037 (N_12037,N_9846,N_7948);
or U12038 (N_12038,N_8757,N_8908);
and U12039 (N_12039,N_9034,N_8477);
nor U12040 (N_12040,N_9079,N_8336);
nand U12041 (N_12041,N_8356,N_7899);
or U12042 (N_12042,N_9010,N_8374);
nor U12043 (N_12043,N_9489,N_9412);
and U12044 (N_12044,N_8510,N_7902);
and U12045 (N_12045,N_7683,N_7594);
xor U12046 (N_12046,N_9322,N_7951);
nand U12047 (N_12047,N_9609,N_7550);
nand U12048 (N_12048,N_9301,N_9886);
nand U12049 (N_12049,N_9936,N_7888);
nand U12050 (N_12050,N_7868,N_8578);
xor U12051 (N_12051,N_8695,N_8941);
nand U12052 (N_12052,N_9030,N_9833);
nor U12053 (N_12053,N_7560,N_8235);
and U12054 (N_12054,N_8971,N_7886);
and U12055 (N_12055,N_9780,N_9674);
and U12056 (N_12056,N_9822,N_9914);
nand U12057 (N_12057,N_8250,N_9971);
nand U12058 (N_12058,N_7952,N_9203);
nor U12059 (N_12059,N_9390,N_9665);
xor U12060 (N_12060,N_8625,N_9409);
or U12061 (N_12061,N_9491,N_8225);
or U12062 (N_12062,N_9348,N_8709);
nor U12063 (N_12063,N_8007,N_7673);
nor U12064 (N_12064,N_9478,N_9992);
xor U12065 (N_12065,N_9874,N_9090);
and U12066 (N_12066,N_8491,N_8612);
and U12067 (N_12067,N_9662,N_7775);
nor U12068 (N_12068,N_8639,N_8191);
nand U12069 (N_12069,N_9000,N_8258);
nand U12070 (N_12070,N_8777,N_7615);
xor U12071 (N_12071,N_8182,N_8866);
nand U12072 (N_12072,N_9361,N_8777);
and U12073 (N_12073,N_8204,N_9308);
nor U12074 (N_12074,N_8029,N_8922);
nor U12075 (N_12075,N_9106,N_8084);
xnor U12076 (N_12076,N_7694,N_8901);
and U12077 (N_12077,N_7596,N_8801);
nand U12078 (N_12078,N_8403,N_9395);
and U12079 (N_12079,N_9974,N_8758);
xnor U12080 (N_12080,N_8141,N_9233);
nor U12081 (N_12081,N_8866,N_8183);
nand U12082 (N_12082,N_8648,N_9653);
and U12083 (N_12083,N_9934,N_7971);
or U12084 (N_12084,N_7806,N_7527);
xor U12085 (N_12085,N_8758,N_9437);
nand U12086 (N_12086,N_9130,N_9590);
xor U12087 (N_12087,N_7703,N_7555);
xnor U12088 (N_12088,N_9605,N_9235);
nand U12089 (N_12089,N_8637,N_9911);
nor U12090 (N_12090,N_8779,N_7981);
or U12091 (N_12091,N_9202,N_9206);
or U12092 (N_12092,N_9409,N_9430);
xor U12093 (N_12093,N_8407,N_7730);
xor U12094 (N_12094,N_8049,N_9611);
and U12095 (N_12095,N_9562,N_8803);
or U12096 (N_12096,N_8150,N_8778);
and U12097 (N_12097,N_9155,N_8783);
nor U12098 (N_12098,N_9709,N_7967);
and U12099 (N_12099,N_8535,N_8740);
and U12100 (N_12100,N_8674,N_9565);
nand U12101 (N_12101,N_7698,N_9132);
and U12102 (N_12102,N_9401,N_8189);
nand U12103 (N_12103,N_9794,N_8629);
xnor U12104 (N_12104,N_9746,N_7907);
xnor U12105 (N_12105,N_8078,N_8804);
and U12106 (N_12106,N_9721,N_9863);
nand U12107 (N_12107,N_9201,N_9381);
or U12108 (N_12108,N_8847,N_8945);
and U12109 (N_12109,N_7750,N_9383);
and U12110 (N_12110,N_8393,N_7520);
and U12111 (N_12111,N_9595,N_9137);
xor U12112 (N_12112,N_9947,N_7759);
and U12113 (N_12113,N_8233,N_8278);
nor U12114 (N_12114,N_8359,N_8907);
nand U12115 (N_12115,N_8823,N_7881);
nor U12116 (N_12116,N_9352,N_8376);
xor U12117 (N_12117,N_8115,N_7581);
xor U12118 (N_12118,N_9628,N_9323);
nand U12119 (N_12119,N_8054,N_9222);
nor U12120 (N_12120,N_7923,N_8446);
and U12121 (N_12121,N_7702,N_8932);
nand U12122 (N_12122,N_7937,N_8996);
nand U12123 (N_12123,N_9035,N_8701);
xnor U12124 (N_12124,N_9923,N_8659);
nor U12125 (N_12125,N_7543,N_9560);
and U12126 (N_12126,N_8547,N_8610);
and U12127 (N_12127,N_9173,N_9361);
nor U12128 (N_12128,N_7570,N_9711);
xor U12129 (N_12129,N_9724,N_8972);
and U12130 (N_12130,N_7888,N_7997);
nor U12131 (N_12131,N_7610,N_8236);
and U12132 (N_12132,N_9451,N_7650);
or U12133 (N_12133,N_9847,N_9422);
xor U12134 (N_12134,N_8033,N_9766);
nand U12135 (N_12135,N_7825,N_8771);
nor U12136 (N_12136,N_9167,N_9615);
and U12137 (N_12137,N_8411,N_7595);
nor U12138 (N_12138,N_9036,N_8723);
and U12139 (N_12139,N_9772,N_8851);
nand U12140 (N_12140,N_9355,N_9626);
nor U12141 (N_12141,N_7833,N_9306);
nor U12142 (N_12142,N_8915,N_9946);
nor U12143 (N_12143,N_9638,N_9992);
and U12144 (N_12144,N_8204,N_7676);
and U12145 (N_12145,N_8284,N_8980);
xor U12146 (N_12146,N_8972,N_9095);
xnor U12147 (N_12147,N_8941,N_8936);
nand U12148 (N_12148,N_9069,N_9579);
xnor U12149 (N_12149,N_8898,N_7944);
or U12150 (N_12150,N_8029,N_9248);
nand U12151 (N_12151,N_8821,N_9788);
xnor U12152 (N_12152,N_8293,N_8646);
nor U12153 (N_12153,N_9200,N_9539);
xnor U12154 (N_12154,N_7780,N_9273);
nor U12155 (N_12155,N_9752,N_9849);
or U12156 (N_12156,N_9452,N_7717);
nor U12157 (N_12157,N_9586,N_8435);
xnor U12158 (N_12158,N_9110,N_9426);
nand U12159 (N_12159,N_8253,N_8121);
nand U12160 (N_12160,N_9537,N_9959);
nand U12161 (N_12161,N_7725,N_9656);
or U12162 (N_12162,N_7795,N_8187);
nand U12163 (N_12163,N_9729,N_8555);
nor U12164 (N_12164,N_8905,N_8303);
nor U12165 (N_12165,N_8511,N_8842);
nand U12166 (N_12166,N_9038,N_7907);
nand U12167 (N_12167,N_9912,N_8166);
and U12168 (N_12168,N_8239,N_8028);
nand U12169 (N_12169,N_9831,N_8753);
nor U12170 (N_12170,N_8346,N_7732);
nand U12171 (N_12171,N_8703,N_9410);
xnor U12172 (N_12172,N_8337,N_7845);
nor U12173 (N_12173,N_8033,N_8743);
nand U12174 (N_12174,N_9161,N_8465);
xor U12175 (N_12175,N_9333,N_8108);
or U12176 (N_12176,N_8572,N_7743);
nor U12177 (N_12177,N_9396,N_8224);
and U12178 (N_12178,N_7830,N_9535);
nand U12179 (N_12179,N_9448,N_8162);
or U12180 (N_12180,N_9320,N_8841);
or U12181 (N_12181,N_8624,N_8332);
or U12182 (N_12182,N_8366,N_9097);
or U12183 (N_12183,N_9541,N_8183);
and U12184 (N_12184,N_8790,N_9421);
and U12185 (N_12185,N_9070,N_7981);
nor U12186 (N_12186,N_8870,N_9394);
nor U12187 (N_12187,N_9996,N_7585);
and U12188 (N_12188,N_8468,N_7828);
xnor U12189 (N_12189,N_9685,N_9402);
nor U12190 (N_12190,N_9648,N_9667);
xor U12191 (N_12191,N_9573,N_9893);
nor U12192 (N_12192,N_9947,N_9339);
nor U12193 (N_12193,N_9157,N_7616);
xnor U12194 (N_12194,N_7536,N_8215);
xnor U12195 (N_12195,N_8778,N_9461);
nand U12196 (N_12196,N_8317,N_7819);
xnor U12197 (N_12197,N_8126,N_9264);
nor U12198 (N_12198,N_8766,N_9602);
or U12199 (N_12199,N_9648,N_8125);
nand U12200 (N_12200,N_8946,N_9938);
or U12201 (N_12201,N_8002,N_9553);
and U12202 (N_12202,N_8802,N_8879);
and U12203 (N_12203,N_9753,N_9433);
nand U12204 (N_12204,N_9738,N_8206);
nor U12205 (N_12205,N_9771,N_9921);
xnor U12206 (N_12206,N_8651,N_9989);
or U12207 (N_12207,N_9582,N_9136);
xor U12208 (N_12208,N_7942,N_9490);
nor U12209 (N_12209,N_9003,N_9232);
and U12210 (N_12210,N_8120,N_7930);
or U12211 (N_12211,N_8350,N_8720);
nand U12212 (N_12212,N_7542,N_9167);
and U12213 (N_12213,N_9201,N_7617);
and U12214 (N_12214,N_8800,N_8041);
or U12215 (N_12215,N_9508,N_9216);
nand U12216 (N_12216,N_9906,N_8723);
nor U12217 (N_12217,N_8756,N_8572);
xnor U12218 (N_12218,N_8656,N_9947);
nand U12219 (N_12219,N_9984,N_9278);
nand U12220 (N_12220,N_8673,N_8554);
and U12221 (N_12221,N_8470,N_9333);
and U12222 (N_12222,N_9147,N_7845);
nor U12223 (N_12223,N_8159,N_8584);
xnor U12224 (N_12224,N_7765,N_7742);
or U12225 (N_12225,N_8619,N_9165);
or U12226 (N_12226,N_8450,N_8039);
xnor U12227 (N_12227,N_9389,N_8730);
or U12228 (N_12228,N_8290,N_9354);
and U12229 (N_12229,N_8290,N_8704);
nand U12230 (N_12230,N_9133,N_9955);
nor U12231 (N_12231,N_9584,N_7998);
xor U12232 (N_12232,N_8679,N_8355);
and U12233 (N_12233,N_9766,N_8754);
nor U12234 (N_12234,N_8152,N_9153);
or U12235 (N_12235,N_9203,N_9394);
xnor U12236 (N_12236,N_8601,N_9990);
nand U12237 (N_12237,N_8172,N_9897);
nor U12238 (N_12238,N_9699,N_9907);
nand U12239 (N_12239,N_9293,N_9027);
or U12240 (N_12240,N_8595,N_8574);
xnor U12241 (N_12241,N_9558,N_9382);
nor U12242 (N_12242,N_7527,N_8726);
nor U12243 (N_12243,N_9801,N_7858);
or U12244 (N_12244,N_8064,N_9418);
nor U12245 (N_12245,N_8092,N_8627);
and U12246 (N_12246,N_8151,N_7899);
or U12247 (N_12247,N_7796,N_9670);
nand U12248 (N_12248,N_7936,N_9162);
or U12249 (N_12249,N_7827,N_7828);
nor U12250 (N_12250,N_8891,N_9222);
nor U12251 (N_12251,N_9962,N_7521);
or U12252 (N_12252,N_8900,N_8752);
and U12253 (N_12253,N_9612,N_9036);
xnor U12254 (N_12254,N_8097,N_9022);
nand U12255 (N_12255,N_9855,N_7943);
or U12256 (N_12256,N_9889,N_9291);
xor U12257 (N_12257,N_7799,N_9653);
xnor U12258 (N_12258,N_7808,N_9380);
and U12259 (N_12259,N_8650,N_9861);
nor U12260 (N_12260,N_8901,N_9095);
and U12261 (N_12261,N_7748,N_9466);
xor U12262 (N_12262,N_8948,N_9115);
nor U12263 (N_12263,N_9651,N_9013);
nand U12264 (N_12264,N_8974,N_8688);
and U12265 (N_12265,N_7792,N_9084);
or U12266 (N_12266,N_8737,N_9894);
xnor U12267 (N_12267,N_9962,N_8071);
nor U12268 (N_12268,N_8831,N_9325);
or U12269 (N_12269,N_9757,N_8991);
nand U12270 (N_12270,N_9998,N_9121);
and U12271 (N_12271,N_8633,N_8847);
and U12272 (N_12272,N_8716,N_8618);
nor U12273 (N_12273,N_8574,N_8166);
xor U12274 (N_12274,N_8874,N_7573);
nor U12275 (N_12275,N_8920,N_8832);
nand U12276 (N_12276,N_9179,N_9518);
xor U12277 (N_12277,N_8928,N_8790);
nand U12278 (N_12278,N_8573,N_8683);
nor U12279 (N_12279,N_9928,N_9264);
xor U12280 (N_12280,N_9603,N_9707);
or U12281 (N_12281,N_9984,N_9220);
xnor U12282 (N_12282,N_7840,N_8219);
and U12283 (N_12283,N_9409,N_9939);
and U12284 (N_12284,N_7662,N_7816);
nand U12285 (N_12285,N_9755,N_9176);
or U12286 (N_12286,N_7566,N_7855);
xor U12287 (N_12287,N_8592,N_9571);
xnor U12288 (N_12288,N_9324,N_9920);
nand U12289 (N_12289,N_8008,N_9730);
nand U12290 (N_12290,N_8881,N_9977);
nor U12291 (N_12291,N_8250,N_7912);
and U12292 (N_12292,N_8919,N_9871);
or U12293 (N_12293,N_7806,N_9383);
xnor U12294 (N_12294,N_7707,N_9444);
and U12295 (N_12295,N_9192,N_9324);
or U12296 (N_12296,N_8179,N_9824);
and U12297 (N_12297,N_8633,N_7650);
and U12298 (N_12298,N_7634,N_9479);
or U12299 (N_12299,N_8473,N_8463);
nand U12300 (N_12300,N_9970,N_9340);
xor U12301 (N_12301,N_9186,N_8722);
xnor U12302 (N_12302,N_8100,N_8746);
nand U12303 (N_12303,N_9646,N_9791);
nand U12304 (N_12304,N_8695,N_8789);
and U12305 (N_12305,N_8789,N_8757);
or U12306 (N_12306,N_8534,N_9174);
xnor U12307 (N_12307,N_9624,N_8513);
nand U12308 (N_12308,N_8926,N_8858);
xor U12309 (N_12309,N_9214,N_8914);
nor U12310 (N_12310,N_8410,N_8723);
and U12311 (N_12311,N_9159,N_9262);
nor U12312 (N_12312,N_9730,N_7576);
nand U12313 (N_12313,N_7664,N_9444);
and U12314 (N_12314,N_9526,N_8207);
and U12315 (N_12315,N_9527,N_7805);
or U12316 (N_12316,N_9391,N_8619);
nor U12317 (N_12317,N_8963,N_8934);
nor U12318 (N_12318,N_7820,N_8170);
xnor U12319 (N_12319,N_8614,N_8770);
nand U12320 (N_12320,N_7592,N_8984);
or U12321 (N_12321,N_8105,N_9840);
nor U12322 (N_12322,N_8363,N_9370);
or U12323 (N_12323,N_8000,N_7682);
xor U12324 (N_12324,N_7583,N_8657);
nor U12325 (N_12325,N_9357,N_8972);
xor U12326 (N_12326,N_9793,N_9896);
and U12327 (N_12327,N_8868,N_9649);
and U12328 (N_12328,N_9655,N_8893);
xnor U12329 (N_12329,N_9605,N_7962);
nor U12330 (N_12330,N_9486,N_7990);
nand U12331 (N_12331,N_7725,N_9775);
and U12332 (N_12332,N_9998,N_8943);
xor U12333 (N_12333,N_8185,N_8297);
xor U12334 (N_12334,N_9231,N_9328);
nand U12335 (N_12335,N_9412,N_8343);
nand U12336 (N_12336,N_9167,N_9135);
nand U12337 (N_12337,N_7682,N_9883);
xor U12338 (N_12338,N_9301,N_8487);
xor U12339 (N_12339,N_9150,N_9925);
xnor U12340 (N_12340,N_8088,N_8089);
nand U12341 (N_12341,N_8687,N_9650);
xor U12342 (N_12342,N_8979,N_7855);
xnor U12343 (N_12343,N_9425,N_8374);
xor U12344 (N_12344,N_8354,N_7689);
or U12345 (N_12345,N_7552,N_8106);
nand U12346 (N_12346,N_8212,N_9256);
and U12347 (N_12347,N_8331,N_8501);
or U12348 (N_12348,N_8269,N_8150);
or U12349 (N_12349,N_9275,N_7593);
nor U12350 (N_12350,N_9813,N_8290);
and U12351 (N_12351,N_7563,N_9322);
nor U12352 (N_12352,N_8457,N_9292);
nand U12353 (N_12353,N_7897,N_9449);
and U12354 (N_12354,N_9207,N_8419);
xnor U12355 (N_12355,N_7811,N_7854);
nand U12356 (N_12356,N_9486,N_8800);
nand U12357 (N_12357,N_9389,N_9550);
and U12358 (N_12358,N_7854,N_7655);
nand U12359 (N_12359,N_8207,N_8518);
nand U12360 (N_12360,N_7998,N_8353);
nor U12361 (N_12361,N_8915,N_8404);
nor U12362 (N_12362,N_9351,N_9276);
nor U12363 (N_12363,N_7606,N_9662);
nor U12364 (N_12364,N_7723,N_7681);
nand U12365 (N_12365,N_7781,N_9604);
xor U12366 (N_12366,N_9721,N_8471);
and U12367 (N_12367,N_7841,N_9201);
nand U12368 (N_12368,N_9257,N_9772);
xor U12369 (N_12369,N_8405,N_9199);
and U12370 (N_12370,N_8688,N_9677);
or U12371 (N_12371,N_9563,N_8905);
xnor U12372 (N_12372,N_9922,N_9576);
nor U12373 (N_12373,N_8564,N_9539);
or U12374 (N_12374,N_8037,N_8184);
nor U12375 (N_12375,N_8134,N_9869);
xor U12376 (N_12376,N_9413,N_7701);
xnor U12377 (N_12377,N_7929,N_8017);
nand U12378 (N_12378,N_8926,N_8918);
and U12379 (N_12379,N_7882,N_9817);
nor U12380 (N_12380,N_9096,N_7525);
nor U12381 (N_12381,N_7619,N_8511);
nand U12382 (N_12382,N_8227,N_8921);
or U12383 (N_12383,N_8777,N_8005);
and U12384 (N_12384,N_7577,N_8918);
or U12385 (N_12385,N_7705,N_8360);
nand U12386 (N_12386,N_8200,N_8263);
nand U12387 (N_12387,N_7579,N_9593);
or U12388 (N_12388,N_8781,N_9844);
or U12389 (N_12389,N_9144,N_8195);
or U12390 (N_12390,N_7953,N_9471);
xor U12391 (N_12391,N_7902,N_8723);
nor U12392 (N_12392,N_9800,N_7858);
and U12393 (N_12393,N_8501,N_9569);
nor U12394 (N_12394,N_9530,N_9844);
or U12395 (N_12395,N_9383,N_8192);
xor U12396 (N_12396,N_8532,N_9974);
xnor U12397 (N_12397,N_8474,N_8969);
nor U12398 (N_12398,N_8782,N_8667);
nand U12399 (N_12399,N_9781,N_9381);
xor U12400 (N_12400,N_8353,N_8652);
nand U12401 (N_12401,N_9059,N_8058);
xnor U12402 (N_12402,N_8154,N_9026);
and U12403 (N_12403,N_9430,N_7730);
or U12404 (N_12404,N_8570,N_8602);
nor U12405 (N_12405,N_9037,N_9659);
nor U12406 (N_12406,N_7964,N_8813);
xnor U12407 (N_12407,N_8957,N_9699);
nor U12408 (N_12408,N_8326,N_9426);
xnor U12409 (N_12409,N_9874,N_9994);
nand U12410 (N_12410,N_9127,N_9253);
nor U12411 (N_12411,N_7531,N_7826);
nand U12412 (N_12412,N_7695,N_9243);
or U12413 (N_12413,N_9592,N_8494);
xnor U12414 (N_12414,N_8592,N_9768);
nand U12415 (N_12415,N_7823,N_8949);
nor U12416 (N_12416,N_8201,N_8222);
nand U12417 (N_12417,N_9420,N_8942);
xor U12418 (N_12418,N_7869,N_9000);
or U12419 (N_12419,N_8972,N_9796);
xor U12420 (N_12420,N_7838,N_9639);
nor U12421 (N_12421,N_9661,N_9604);
and U12422 (N_12422,N_9359,N_7835);
xor U12423 (N_12423,N_9585,N_9403);
or U12424 (N_12424,N_9107,N_7944);
or U12425 (N_12425,N_9284,N_9442);
nand U12426 (N_12426,N_8323,N_8278);
and U12427 (N_12427,N_8974,N_9300);
and U12428 (N_12428,N_9875,N_7917);
and U12429 (N_12429,N_7666,N_9527);
nand U12430 (N_12430,N_7666,N_7576);
nand U12431 (N_12431,N_9934,N_8254);
or U12432 (N_12432,N_8973,N_9555);
or U12433 (N_12433,N_7818,N_9025);
nor U12434 (N_12434,N_9078,N_8383);
or U12435 (N_12435,N_7788,N_7940);
nor U12436 (N_12436,N_9357,N_8348);
xnor U12437 (N_12437,N_8126,N_9706);
nor U12438 (N_12438,N_9561,N_8294);
and U12439 (N_12439,N_9486,N_8947);
and U12440 (N_12440,N_9039,N_8995);
nor U12441 (N_12441,N_8840,N_9964);
nor U12442 (N_12442,N_9973,N_8330);
and U12443 (N_12443,N_7678,N_9945);
nand U12444 (N_12444,N_9998,N_7805);
nor U12445 (N_12445,N_9494,N_9875);
xnor U12446 (N_12446,N_7976,N_8576);
nand U12447 (N_12447,N_7599,N_9554);
nand U12448 (N_12448,N_8306,N_9422);
or U12449 (N_12449,N_8637,N_7759);
nor U12450 (N_12450,N_9915,N_8893);
xnor U12451 (N_12451,N_7993,N_8684);
or U12452 (N_12452,N_9831,N_7668);
xnor U12453 (N_12453,N_8789,N_9309);
nand U12454 (N_12454,N_8474,N_9180);
xor U12455 (N_12455,N_8259,N_7646);
nor U12456 (N_12456,N_7763,N_7878);
xnor U12457 (N_12457,N_7815,N_8107);
or U12458 (N_12458,N_8667,N_8899);
nand U12459 (N_12459,N_8697,N_9568);
and U12460 (N_12460,N_8862,N_9524);
nor U12461 (N_12461,N_9581,N_8942);
nor U12462 (N_12462,N_9896,N_8842);
xor U12463 (N_12463,N_9821,N_9834);
xnor U12464 (N_12464,N_8820,N_8866);
nand U12465 (N_12465,N_7621,N_7863);
nand U12466 (N_12466,N_9608,N_9703);
nand U12467 (N_12467,N_9337,N_8481);
and U12468 (N_12468,N_9268,N_9075);
and U12469 (N_12469,N_7934,N_9071);
and U12470 (N_12470,N_8025,N_7943);
xnor U12471 (N_12471,N_8666,N_9961);
nand U12472 (N_12472,N_8027,N_9831);
or U12473 (N_12473,N_8860,N_9030);
nor U12474 (N_12474,N_9203,N_8498);
xnor U12475 (N_12475,N_7912,N_8195);
or U12476 (N_12476,N_8745,N_7802);
or U12477 (N_12477,N_9462,N_8942);
nor U12478 (N_12478,N_8252,N_9809);
nor U12479 (N_12479,N_7864,N_9922);
xor U12480 (N_12480,N_8754,N_7849);
and U12481 (N_12481,N_9743,N_9661);
nor U12482 (N_12482,N_7767,N_9737);
nand U12483 (N_12483,N_9747,N_9662);
nand U12484 (N_12484,N_9384,N_9338);
and U12485 (N_12485,N_9300,N_9210);
and U12486 (N_12486,N_7994,N_8855);
or U12487 (N_12487,N_9000,N_8385);
or U12488 (N_12488,N_9141,N_9477);
or U12489 (N_12489,N_7822,N_8299);
and U12490 (N_12490,N_9586,N_8218);
nor U12491 (N_12491,N_9161,N_8633);
nor U12492 (N_12492,N_7725,N_8774);
nand U12493 (N_12493,N_9590,N_7538);
or U12494 (N_12494,N_8130,N_9123);
nand U12495 (N_12495,N_7629,N_9593);
xor U12496 (N_12496,N_8290,N_9614);
xnor U12497 (N_12497,N_8929,N_8595);
nand U12498 (N_12498,N_9395,N_7657);
xnor U12499 (N_12499,N_7895,N_8673);
xnor U12500 (N_12500,N_11431,N_10915);
xor U12501 (N_12501,N_11882,N_11938);
xnor U12502 (N_12502,N_12368,N_11883);
and U12503 (N_12503,N_11174,N_12111);
or U12504 (N_12504,N_10427,N_11454);
or U12505 (N_12505,N_11961,N_12133);
nand U12506 (N_12506,N_12106,N_11237);
nor U12507 (N_12507,N_12374,N_11985);
xor U12508 (N_12508,N_10560,N_10203);
or U12509 (N_12509,N_11274,N_10200);
or U12510 (N_12510,N_12156,N_10658);
nor U12511 (N_12511,N_10565,N_10387);
nand U12512 (N_12512,N_11689,N_10342);
or U12513 (N_12513,N_12383,N_12105);
nor U12514 (N_12514,N_10063,N_12011);
nand U12515 (N_12515,N_10976,N_12141);
and U12516 (N_12516,N_12357,N_12277);
xnor U12517 (N_12517,N_10491,N_10157);
nor U12518 (N_12518,N_10390,N_12012);
nor U12519 (N_12519,N_10174,N_11583);
xor U12520 (N_12520,N_12470,N_11624);
nand U12521 (N_12521,N_10636,N_11255);
nand U12522 (N_12522,N_11111,N_11369);
and U12523 (N_12523,N_12196,N_11975);
xor U12524 (N_12524,N_10949,N_11780);
nand U12525 (N_12525,N_10146,N_12436);
xor U12526 (N_12526,N_10569,N_11004);
or U12527 (N_12527,N_10627,N_11208);
and U12528 (N_12528,N_10317,N_10988);
nand U12529 (N_12529,N_10444,N_12082);
and U12530 (N_12530,N_10014,N_12272);
and U12531 (N_12531,N_10013,N_11435);
xor U12532 (N_12532,N_11867,N_11118);
or U12533 (N_12533,N_10113,N_11341);
and U12534 (N_12534,N_10354,N_10183);
and U12535 (N_12535,N_12055,N_11771);
nor U12536 (N_12536,N_10034,N_11407);
nor U12537 (N_12537,N_12227,N_11535);
and U12538 (N_12538,N_10641,N_12154);
nor U12539 (N_12539,N_10248,N_10144);
and U12540 (N_12540,N_10796,N_12188);
and U12541 (N_12541,N_10494,N_12481);
or U12542 (N_12542,N_10101,N_12119);
and U12543 (N_12543,N_12038,N_11748);
nand U12544 (N_12544,N_11877,N_11155);
nor U12545 (N_12545,N_11272,N_11443);
nor U12546 (N_12546,N_11198,N_12139);
and U12547 (N_12547,N_11891,N_10746);
nor U12548 (N_12548,N_11516,N_10417);
xor U12549 (N_12549,N_10630,N_11502);
or U12550 (N_12550,N_10587,N_11756);
nand U12551 (N_12551,N_10980,N_10100);
and U12552 (N_12552,N_10679,N_10234);
and U12553 (N_12553,N_11219,N_12427);
nand U12554 (N_12554,N_10622,N_11621);
and U12555 (N_12555,N_11599,N_10716);
nor U12556 (N_12556,N_11787,N_11165);
and U12557 (N_12557,N_10628,N_11334);
nand U12558 (N_12558,N_12483,N_11193);
xnor U12559 (N_12559,N_11013,N_10530);
nor U12560 (N_12560,N_10793,N_12214);
or U12561 (N_12561,N_12009,N_11082);
and U12562 (N_12562,N_12278,N_11500);
and U12563 (N_12563,N_12376,N_12144);
or U12564 (N_12564,N_10030,N_11721);
or U12565 (N_12565,N_12304,N_12155);
or U12566 (N_12566,N_10833,N_11186);
or U12567 (N_12567,N_10676,N_11570);
nor U12568 (N_12568,N_11293,N_10597);
and U12569 (N_12569,N_11052,N_10753);
or U12570 (N_12570,N_11055,N_11762);
nor U12571 (N_12571,N_11180,N_11349);
xor U12572 (N_12572,N_11241,N_11470);
nand U12573 (N_12573,N_11826,N_11916);
nor U12574 (N_12574,N_12322,N_11409);
or U12575 (N_12575,N_11283,N_11618);
and U12576 (N_12576,N_11852,N_12053);
xnor U12577 (N_12577,N_11727,N_11973);
nand U12578 (N_12578,N_11853,N_10149);
or U12579 (N_12579,N_10650,N_11758);
and U12580 (N_12580,N_10859,N_11956);
nor U12581 (N_12581,N_11113,N_11396);
or U12582 (N_12582,N_10791,N_10270);
xnor U12583 (N_12583,N_11368,N_10255);
nand U12584 (N_12584,N_11311,N_12181);
and U12585 (N_12585,N_12403,N_11009);
xnor U12586 (N_12586,N_11143,N_11517);
or U12587 (N_12587,N_11838,N_10640);
nand U12588 (N_12588,N_10700,N_11147);
nor U12589 (N_12589,N_10900,N_10201);
nor U12590 (N_12590,N_10111,N_10947);
nand U12591 (N_12591,N_12281,N_12245);
or U12592 (N_12592,N_11121,N_10575);
or U12593 (N_12593,N_11954,N_10328);
nand U12594 (N_12594,N_10286,N_10067);
nand U12595 (N_12595,N_11706,N_12173);
or U12596 (N_12596,N_10142,N_10792);
or U12597 (N_12597,N_11753,N_12107);
xor U12598 (N_12598,N_11430,N_12120);
xor U12599 (N_12599,N_10849,N_10618);
nand U12600 (N_12600,N_10367,N_10432);
and U12601 (N_12601,N_10683,N_11587);
xor U12602 (N_12602,N_10840,N_11868);
xor U12603 (N_12603,N_10845,N_10141);
or U12604 (N_12604,N_10528,N_10508);
and U12605 (N_12605,N_11832,N_10023);
or U12606 (N_12606,N_11148,N_11209);
and U12607 (N_12607,N_11402,N_12222);
xor U12608 (N_12608,N_12033,N_10841);
or U12609 (N_12609,N_10937,N_11002);
or U12610 (N_12610,N_10971,N_11432);
and U12611 (N_12611,N_11476,N_10264);
nor U12612 (N_12612,N_11589,N_10969);
nor U12613 (N_12613,N_12429,N_10300);
xor U12614 (N_12614,N_10288,N_11811);
xnor U12615 (N_12615,N_12242,N_10522);
or U12616 (N_12616,N_10254,N_12293);
nor U12617 (N_12617,N_11153,N_10842);
nor U12618 (N_12618,N_10661,N_12152);
nand U12619 (N_12619,N_11722,N_10684);
nand U12620 (N_12620,N_11647,N_11588);
nor U12621 (N_12621,N_10393,N_10523);
xnor U12622 (N_12622,N_12412,N_11046);
xnor U12623 (N_12623,N_11640,N_12269);
xor U12624 (N_12624,N_10357,N_12497);
and U12625 (N_12625,N_10327,N_11295);
nand U12626 (N_12626,N_10245,N_11804);
xnor U12627 (N_12627,N_10782,N_11623);
and U12628 (N_12628,N_12330,N_11875);
xor U12629 (N_12629,N_10031,N_10130);
nand U12630 (N_12630,N_10340,N_10785);
or U12631 (N_12631,N_10088,N_11923);
and U12632 (N_12632,N_10828,N_10046);
and U12633 (N_12633,N_11404,N_12070);
and U12634 (N_12634,N_11918,N_11459);
nor U12635 (N_12635,N_10957,N_11253);
xnor U12636 (N_12636,N_12402,N_11466);
and U12637 (N_12637,N_11783,N_10419);
or U12638 (N_12638,N_10017,N_12075);
xnor U12639 (N_12639,N_11936,N_11854);
xnor U12640 (N_12640,N_12236,N_10206);
and U12641 (N_12641,N_11890,N_12093);
and U12642 (N_12642,N_10158,N_10552);
or U12643 (N_12643,N_12375,N_11702);
xnor U12644 (N_12644,N_11742,N_11665);
xnor U12645 (N_12645,N_11486,N_10148);
nor U12646 (N_12646,N_10981,N_10706);
nand U12647 (N_12647,N_11108,N_10389);
nand U12648 (N_12648,N_11651,N_10495);
nor U12649 (N_12649,N_12489,N_11371);
nor U12650 (N_12650,N_10068,N_10790);
and U12651 (N_12651,N_10663,N_11426);
or U12652 (N_12652,N_12089,N_11061);
and U12653 (N_12653,N_10098,N_11413);
or U12654 (N_12654,N_11805,N_10708);
and U12655 (N_12655,N_12298,N_12165);
and U12656 (N_12656,N_11455,N_11541);
nor U12657 (N_12657,N_12232,N_10576);
and U12658 (N_12658,N_12319,N_10179);
nand U12659 (N_12659,N_11419,N_10103);
nand U12660 (N_12660,N_10305,N_10194);
or U12661 (N_12661,N_12449,N_11635);
and U12662 (N_12662,N_12078,N_12099);
or U12663 (N_12663,N_11841,N_10431);
nor U12664 (N_12664,N_10167,N_11513);
xor U12665 (N_12665,N_10208,N_11194);
nand U12666 (N_12666,N_10211,N_11851);
or U12667 (N_12667,N_12389,N_11417);
and U12668 (N_12668,N_10446,N_11090);
xnor U12669 (N_12669,N_10048,N_10757);
xor U12670 (N_12670,N_10341,N_10225);
xor U12671 (N_12671,N_12345,N_12225);
nand U12672 (N_12672,N_12036,N_10540);
or U12673 (N_12673,N_11515,N_10818);
nor U12674 (N_12674,N_11873,N_10909);
or U12675 (N_12675,N_11896,N_10052);
nand U12676 (N_12676,N_11187,N_10513);
or U12677 (N_12677,N_10449,N_12294);
nand U12678 (N_12678,N_12025,N_12018);
or U12679 (N_12679,N_10244,N_12359);
or U12680 (N_12680,N_11031,N_11083);
nand U12681 (N_12681,N_10262,N_10302);
nor U12682 (N_12682,N_12360,N_12339);
nor U12683 (N_12683,N_10715,N_11669);
or U12684 (N_12684,N_11150,N_11590);
xnor U12685 (N_12685,N_11709,N_12349);
and U12686 (N_12686,N_10370,N_11385);
or U12687 (N_12687,N_11955,N_12194);
and U12688 (N_12688,N_10418,N_11595);
and U12689 (N_12689,N_11444,N_11892);
xnor U12690 (N_12690,N_12302,N_12076);
and U12691 (N_12691,N_11097,N_11633);
or U12692 (N_12692,N_11981,N_11792);
or U12693 (N_12693,N_10107,N_12109);
xor U12694 (N_12694,N_11585,N_10453);
nand U12695 (N_12695,N_12179,N_11644);
nor U12696 (N_12696,N_10611,N_10751);
nor U12697 (N_12697,N_12084,N_11858);
xor U12698 (N_12698,N_12217,N_10811);
nand U12699 (N_12699,N_10074,N_10136);
or U12700 (N_12700,N_12145,N_11586);
and U12701 (N_12701,N_10821,N_10968);
xor U12702 (N_12702,N_12421,N_11415);
nand U12703 (N_12703,N_10222,N_11078);
xor U12704 (N_12704,N_10917,N_11324);
or U12705 (N_12705,N_10786,N_10664);
nor U12706 (N_12706,N_10693,N_10723);
or U12707 (N_12707,N_12324,N_10524);
xnor U12708 (N_12708,N_11682,N_10333);
and U12709 (N_12709,N_11440,N_10325);
or U12710 (N_12710,N_12467,N_11372);
or U12711 (N_12711,N_10826,N_11309);
nor U12712 (N_12712,N_11262,N_10187);
nor U12713 (N_12713,N_10344,N_11196);
and U12714 (N_12714,N_11197,N_11549);
or U12715 (N_12715,N_10816,N_11625);
and U12716 (N_12716,N_10586,N_11740);
nand U12717 (N_12717,N_10865,N_12477);
xnor U12718 (N_12718,N_10794,N_11354);
xnor U12719 (N_12719,N_10115,N_11845);
or U12720 (N_12720,N_12183,N_12388);
nand U12721 (N_12721,N_10941,N_11144);
and U12722 (N_12722,N_12333,N_10623);
or U12723 (N_12723,N_10078,N_11183);
and U12724 (N_12724,N_10454,N_10110);
xor U12725 (N_12725,N_11604,N_10766);
and U12726 (N_12726,N_10061,N_12387);
and U12727 (N_12727,N_10553,N_12118);
nand U12728 (N_12728,N_12142,N_12331);
and U12729 (N_12729,N_10780,N_12444);
or U12730 (N_12730,N_11442,N_10091);
xor U12731 (N_12731,N_11478,N_10185);
nor U12732 (N_12732,N_10551,N_10882);
xnor U12733 (N_12733,N_12343,N_11266);
xor U12734 (N_12734,N_11984,N_10891);
and U12735 (N_12735,N_11017,N_11356);
xnor U12736 (N_12736,N_11021,N_10484);
and U12737 (N_12737,N_11375,N_11622);
xor U12738 (N_12738,N_11364,N_12317);
nand U12739 (N_12739,N_11317,N_10682);
xor U12740 (N_12740,N_10666,N_12068);
xnor U12741 (N_12741,N_10516,N_10671);
and U12742 (N_12742,N_11037,N_10955);
and U12743 (N_12743,N_12060,N_11462);
nor U12744 (N_12744,N_11292,N_12346);
nand U12745 (N_12745,N_11914,N_12447);
or U12746 (N_12746,N_10163,N_10173);
and U12747 (N_12747,N_11434,N_11260);
xnor U12748 (N_12748,N_10363,N_11377);
and U12749 (N_12749,N_12042,N_10927);
xor U12750 (N_12750,N_11510,N_11678);
nand U12751 (N_12751,N_10614,N_11384);
nand U12752 (N_12752,N_11089,N_10235);
or U12753 (N_12753,N_10388,N_12377);
nand U12754 (N_12754,N_10733,N_10594);
nor U12755 (N_12755,N_10625,N_11073);
xnor U12756 (N_12756,N_10020,N_11287);
or U12757 (N_12757,N_11149,N_12046);
or U12758 (N_12758,N_11632,N_12426);
and U12759 (N_12759,N_10297,N_11701);
nor U12760 (N_12760,N_11910,N_10874);
nor U12761 (N_12761,N_11879,N_11636);
nor U12762 (N_12762,N_11860,N_10605);
and U12763 (N_12763,N_10436,N_12441);
and U12764 (N_12764,N_11857,N_11726);
or U12765 (N_12765,N_11014,N_11765);
nand U12766 (N_12766,N_10543,N_12460);
nand U12767 (N_12767,N_11942,N_11104);
nor U12768 (N_12768,N_10692,N_12292);
and U12769 (N_12769,N_10515,N_12406);
and U12770 (N_12770,N_11573,N_10120);
nand U12771 (N_12771,N_11393,N_10642);
nor U12772 (N_12772,N_10485,N_11359);
or U12773 (N_12773,N_11849,N_10750);
xnor U12774 (N_12774,N_11100,N_12271);
nor U12775 (N_12775,N_10080,N_10345);
nand U12776 (N_12776,N_12126,N_11238);
nor U12777 (N_12777,N_12000,N_11081);
nor U12778 (N_12778,N_10801,N_10273);
nor U12779 (N_12779,N_10137,N_10272);
nand U12780 (N_12780,N_11107,N_11968);
nor U12781 (N_12781,N_10462,N_10466);
nor U12782 (N_12782,N_12007,N_10942);
nor U12783 (N_12783,N_10198,N_10744);
nand U12784 (N_12784,N_11642,N_12401);
xor U12785 (N_12785,N_11784,N_11836);
xor U12786 (N_12786,N_11294,N_10645);
or U12787 (N_12787,N_12233,N_10878);
nor U12788 (N_12788,N_11302,N_12239);
and U12789 (N_12789,N_11313,N_10867);
xor U12790 (N_12790,N_11339,N_12305);
xnor U12791 (N_12791,N_10775,N_10373);
and U12792 (N_12792,N_11029,N_12466);
nand U12793 (N_12793,N_10404,N_11778);
or U12794 (N_12794,N_11130,N_10348);
and U12795 (N_12795,N_11720,N_11275);
and U12796 (N_12796,N_11249,N_11994);
nor U12797 (N_12797,N_12422,N_12158);
nand U12798 (N_12798,N_12417,N_11305);
or U12799 (N_12799,N_12351,N_12485);
nand U12800 (N_12800,N_12226,N_11504);
nand U12801 (N_12801,N_10531,N_10987);
xnor U12802 (N_12802,N_12344,N_10369);
xor U12803 (N_12803,N_11831,N_10691);
xor U12804 (N_12804,N_10820,N_12229);
nor U12805 (N_12805,N_11752,N_10555);
nor U12806 (N_12806,N_10298,N_10675);
nor U12807 (N_12807,N_11609,N_12086);
nor U12808 (N_12808,N_10226,N_11764);
or U12809 (N_12809,N_12061,N_11978);
nor U12810 (N_12810,N_10376,N_10637);
or U12811 (N_12811,N_12031,N_11050);
nand U12812 (N_12812,N_12315,N_10643);
xnor U12813 (N_12813,N_11527,N_10282);
nand U12814 (N_12814,N_10392,N_12313);
nand U12815 (N_12815,N_12321,N_10456);
or U12816 (N_12816,N_10126,N_11724);
nand U12817 (N_12817,N_10481,N_11245);
nand U12818 (N_12818,N_12207,N_12097);
and U12819 (N_12819,N_12049,N_11710);
xnor U12820 (N_12820,N_11472,N_11657);
nand U12821 (N_12821,N_12172,N_10619);
xor U12822 (N_12822,N_10506,N_10151);
xnor U12823 (N_12823,N_10318,N_11593);
nand U12824 (N_12824,N_10421,N_11801);
nand U12825 (N_12825,N_11566,N_10534);
or U12826 (N_12826,N_11224,N_11986);
nor U12827 (N_12827,N_10773,N_10724);
nor U12828 (N_12828,N_12342,N_11864);
nand U12829 (N_12829,N_10680,N_11946);
or U12830 (N_12830,N_10043,N_11025);
nand U12831 (N_12831,N_12115,N_10138);
or U12832 (N_12832,N_12301,N_11005);
or U12833 (N_12833,N_10940,N_12017);
and U12834 (N_12834,N_11420,N_11673);
nand U12835 (N_12835,N_12438,N_12205);
nor U12836 (N_12836,N_12320,N_10958);
or U12837 (N_12837,N_11766,N_10905);
nand U12838 (N_12838,N_11565,N_10592);
and U12839 (N_12839,N_11285,N_10056);
xnor U12840 (N_12840,N_11373,N_10218);
nand U12841 (N_12841,N_10104,N_10799);
nor U12842 (N_12842,N_10055,N_11102);
and U12843 (N_12843,N_12473,N_11592);
nor U12844 (N_12844,N_10191,N_10321);
nand U12845 (N_12845,N_10492,N_11919);
nand U12846 (N_12846,N_10735,N_11460);
xor U12847 (N_12847,N_12113,N_12102);
or U12848 (N_12848,N_11229,N_12202);
or U12849 (N_12849,N_12323,N_11821);
xor U12850 (N_12850,N_11553,N_11619);
nor U12851 (N_12851,N_10422,N_10946);
xnor U12852 (N_12852,N_11427,N_11788);
xnor U12853 (N_12853,N_11785,N_11508);
or U12854 (N_12854,N_11559,N_10756);
or U12855 (N_12855,N_11878,N_12486);
xnor U12856 (N_12856,N_11908,N_10155);
and U12857 (N_12857,N_10379,N_10351);
xor U12858 (N_12858,N_12187,N_10921);
nor U12859 (N_12859,N_10258,N_12338);
nor U12860 (N_12860,N_11607,N_11181);
or U12861 (N_12861,N_10525,N_10916);
nand U12862 (N_12862,N_11794,N_12288);
nand U12863 (N_12863,N_10159,N_10143);
and U12864 (N_12864,N_10924,N_11700);
xor U12865 (N_12865,N_11615,N_10761);
and U12866 (N_12866,N_10223,N_10129);
nand U12867 (N_12867,N_12191,N_10536);
or U12868 (N_12868,N_12475,N_11828);
and U12869 (N_12869,N_11132,N_10895);
xor U12870 (N_12870,N_10097,N_11536);
and U12871 (N_12871,N_11070,N_10696);
and U12872 (N_12872,N_12094,N_11518);
and U12873 (N_12873,N_11812,N_10268);
nand U12874 (N_12874,N_11716,N_12228);
xnor U12875 (N_12875,N_11707,N_11033);
or U12876 (N_12876,N_10337,N_11893);
xor U12877 (N_12877,N_12458,N_10251);
nand U12878 (N_12878,N_10171,N_11803);
and U12879 (N_12879,N_11221,N_11388);
or U12880 (N_12880,N_12405,N_10378);
xor U12881 (N_12881,N_12221,N_11163);
or U12882 (N_12882,N_10058,N_10974);
xor U12883 (N_12883,N_11989,N_10669);
xor U12884 (N_12884,N_10220,N_11468);
or U12885 (N_12885,N_11256,N_12353);
and U12886 (N_12886,N_10473,N_10105);
nor U12887 (N_12887,N_10985,N_11581);
nor U12888 (N_12888,N_12445,N_11905);
xnor U12889 (N_12889,N_11705,N_11880);
or U12890 (N_12890,N_11112,N_10975);
or U12891 (N_12891,N_11370,N_12079);
nand U12892 (N_12892,N_10871,N_10612);
xnor U12893 (N_12893,N_11129,N_12128);
and U12894 (N_12894,N_10320,N_12480);
xnor U12895 (N_12895,N_10809,N_11280);
xor U12896 (N_12896,N_10938,N_12066);
and U12897 (N_12897,N_11212,N_10764);
xnor U12898 (N_12898,N_10933,N_10434);
or U12899 (N_12899,N_10907,N_12051);
or U12900 (N_12900,N_11361,N_12056);
xor U12901 (N_12901,N_10073,N_10480);
xnor U12902 (N_12902,N_11790,N_10463);
nor U12903 (N_12903,N_12280,N_10464);
xnor U12904 (N_12904,N_10616,N_11703);
nand U12905 (N_12905,N_10638,N_10287);
xnor U12906 (N_12906,N_11259,N_11983);
or U12907 (N_12907,N_10918,N_12425);
nor U12908 (N_12908,N_10595,N_12235);
nand U12909 (N_12909,N_12492,N_11437);
or U12910 (N_12910,N_11079,N_11063);
nor U12911 (N_12911,N_10131,N_12266);
and U12912 (N_12912,N_12310,N_11917);
nor U12913 (N_12913,N_11667,N_11929);
xor U12914 (N_12914,N_10970,N_10016);
and U12915 (N_12915,N_10677,N_10960);
xnor U12916 (N_12916,N_11164,N_11243);
and U12917 (N_12917,N_10134,N_12147);
xor U12918 (N_12918,N_11213,N_11216);
and U12919 (N_12919,N_11582,N_12208);
or U12920 (N_12920,N_11234,N_10065);
and U12921 (N_12921,N_11833,N_10240);
nor U12922 (N_12922,N_11214,N_12326);
nor U12923 (N_12923,N_12148,N_12185);
xor U12924 (N_12924,N_11494,N_10800);
and U12925 (N_12925,N_10028,N_10010);
or U12926 (N_12926,N_12382,N_11060);
nor U12927 (N_12927,N_10311,N_12169);
and U12928 (N_12928,N_11085,N_10497);
or U12929 (N_12929,N_10936,N_11066);
xor U12930 (N_12930,N_11357,N_11547);
and U12931 (N_12931,N_12220,N_10527);
or U12932 (N_12932,N_11556,N_11117);
nor U12933 (N_12933,N_10346,N_11834);
nand U12934 (N_12934,N_11477,N_10116);
nand U12935 (N_12935,N_12204,N_10224);
nand U12936 (N_12936,N_12498,N_11023);
or U12937 (N_12937,N_10019,N_11326);
or U12938 (N_12938,N_11552,N_10656);
nor U12939 (N_12939,N_10604,N_11137);
nand U12940 (N_12940,N_11827,N_11489);
or U12941 (N_12941,N_10922,N_11408);
or U12942 (N_12942,N_12309,N_10573);
nand U12943 (N_12943,N_11136,N_12409);
and U12944 (N_12944,N_12218,N_10275);
xor U12945 (N_12945,N_11053,N_11554);
nor U12946 (N_12946,N_11521,N_10205);
xnor U12947 (N_12947,N_10386,N_11899);
xor U12948 (N_12948,N_10364,N_11416);
xor U12949 (N_12949,N_10591,N_10526);
xnor U12950 (N_12950,N_11217,N_10885);
or U12951 (N_12951,N_10039,N_10606);
nor U12952 (N_12952,N_10577,N_11944);
nor U12953 (N_12953,N_12080,N_12354);
xnor U12954 (N_12954,N_11146,N_11514);
nand U12955 (N_12955,N_11533,N_10954);
and U12956 (N_12956,N_10152,N_10465);
nand U12957 (N_12957,N_10053,N_11846);
and U12958 (N_12958,N_10868,N_11410);
or U12959 (N_12959,N_11131,N_12484);
and U12960 (N_12960,N_11015,N_10263);
nor U12961 (N_12961,N_12246,N_11022);
nand U12962 (N_12962,N_12307,N_12316);
xnor U12963 (N_12963,N_11451,N_11481);
nand U12964 (N_12964,N_10475,N_11051);
or U12965 (N_12965,N_10079,N_10247);
or U12966 (N_12966,N_10762,N_12295);
nand U12967 (N_12967,N_10440,N_11943);
and U12968 (N_12968,N_11822,N_12058);
or U12969 (N_12969,N_10292,N_11628);
and U12970 (N_12970,N_11076,N_12267);
nor U12971 (N_12971,N_10660,N_10556);
nand U12972 (N_12972,N_11800,N_10580);
nor U12973 (N_12973,N_10760,N_11452);
nand U12974 (N_12974,N_10003,N_12199);
nand U12975 (N_12975,N_10479,N_11679);
nor U12976 (N_12976,N_12090,N_10549);
nand U12977 (N_12977,N_11158,N_10380);
and U12978 (N_12978,N_11348,N_11273);
nand U12979 (N_12979,N_11597,N_11523);
or U12980 (N_12980,N_12397,N_12190);
xnor U12981 (N_12981,N_10332,N_11603);
or U12982 (N_12982,N_10807,N_11134);
and U12983 (N_12983,N_10309,N_10951);
and U12984 (N_12984,N_10740,N_10928);
xor U12985 (N_12985,N_10992,N_12478);
nor U12986 (N_12986,N_10424,N_11674);
nor U12987 (N_12987,N_10629,N_10731);
nor U12988 (N_12988,N_11677,N_10662);
nor U12989 (N_12989,N_10903,N_11874);
nand U12990 (N_12990,N_11738,N_12071);
or U12991 (N_12991,N_11340,N_11650);
nor U12992 (N_12992,N_10932,N_10261);
or U12993 (N_12993,N_10728,N_11096);
xor U12994 (N_12994,N_12136,N_10727);
nor U12995 (N_12995,N_12116,N_11218);
or U12996 (N_12996,N_12092,N_11842);
or U12997 (N_12997,N_10400,N_10216);
xnor U12998 (N_12998,N_10186,N_12216);
nand U12999 (N_12999,N_12462,N_10215);
nand U13000 (N_13000,N_10803,N_10172);
and U13001 (N_13001,N_11865,N_11655);
nand U13002 (N_13002,N_10391,N_12312);
xnor U13003 (N_13003,N_10445,N_11161);
nand U13004 (N_13004,N_12015,N_12340);
nand U13005 (N_13005,N_12201,N_10950);
xnor U13006 (N_13006,N_12437,N_12325);
and U13007 (N_13007,N_11390,N_10714);
xnor U13008 (N_13008,N_11047,N_11350);
or U13009 (N_13009,N_11652,N_10655);
or U13010 (N_13010,N_11360,N_11059);
and U13011 (N_13011,N_10861,N_10886);
and U13012 (N_13012,N_12180,N_11139);
or U13013 (N_13013,N_10857,N_10926);
or U13014 (N_13014,N_12495,N_11663);
xnor U13015 (N_13015,N_12265,N_10721);
xor U13016 (N_13016,N_10360,N_10024);
and U13017 (N_13017,N_10181,N_11457);
and U13018 (N_13018,N_12479,N_12399);
nand U13019 (N_13019,N_11088,N_10274);
and U13020 (N_13020,N_12446,N_12423);
and U13021 (N_13021,N_10064,N_11571);
or U13022 (N_13022,N_12127,N_12121);
or U13023 (N_13023,N_11438,N_10720);
xnor U13024 (N_13024,N_10877,N_10477);
nor U13025 (N_13025,N_10169,N_10122);
and U13026 (N_13026,N_10678,N_10574);
nor U13027 (N_13027,N_10123,N_10368);
nor U13028 (N_13028,N_10511,N_11101);
xor U13029 (N_13029,N_10631,N_11115);
or U13030 (N_13030,N_11534,N_10410);
nand U13031 (N_13031,N_12013,N_10836);
nor U13032 (N_13032,N_10711,N_10382);
or U13033 (N_13033,N_11487,N_11791);
xnor U13034 (N_13034,N_10910,N_10168);
nor U13035 (N_13035,N_10140,N_11122);
nor U13036 (N_13036,N_11840,N_11316);
and U13037 (N_13037,N_11931,N_11352);
or U13038 (N_13038,N_10219,N_10366);
or U13039 (N_13039,N_11501,N_10355);
nand U13040 (N_13040,N_11577,N_10310);
or U13041 (N_13041,N_11484,N_11694);
xor U13042 (N_13042,N_12366,N_11227);
nor U13043 (N_13043,N_10117,N_12253);
xor U13044 (N_13044,N_10253,N_10266);
nor U13045 (N_13045,N_10579,N_12420);
xor U13046 (N_13046,N_10075,N_11866);
nor U13047 (N_13047,N_10967,N_10241);
nor U13048 (N_13048,N_11483,N_10672);
and U13049 (N_13049,N_11028,N_10461);
and U13050 (N_13050,N_10822,N_10002);
or U13051 (N_13051,N_12219,N_11793);
nor U13052 (N_13052,N_10827,N_12254);
and U13053 (N_13053,N_12224,N_12371);
nand U13054 (N_13054,N_10889,N_10929);
xor U13055 (N_13055,N_12122,N_10635);
nor U13056 (N_13056,N_10986,N_11531);
or U13057 (N_13057,N_11296,N_10593);
nand U13058 (N_13058,N_12268,N_10407);
xor U13059 (N_13059,N_10385,N_10006);
and U13060 (N_13060,N_11817,N_11332);
and U13061 (N_13061,N_11068,N_11969);
or U13062 (N_13062,N_11524,N_11176);
and U13063 (N_13063,N_11167,N_10093);
nand U13064 (N_13064,N_12175,N_11123);
xnor U13065 (N_13065,N_11400,N_12240);
and U13066 (N_13066,N_10228,N_11401);
nand U13067 (N_13067,N_11889,N_10854);
nor U13068 (N_13068,N_11799,N_12212);
nor U13069 (N_13069,N_10601,N_10265);
nand U13070 (N_13070,N_10923,N_11290);
nand U13071 (N_13071,N_12211,N_10999);
xor U13072 (N_13072,N_11639,N_10397);
xnor U13073 (N_13073,N_11634,N_11230);
and U13074 (N_13074,N_10314,N_10457);
nor U13075 (N_13075,N_10808,N_11611);
or U13076 (N_13076,N_12407,N_11380);
nand U13077 (N_13077,N_10331,N_11715);
xnor U13078 (N_13078,N_11281,N_10529);
nor U13079 (N_13079,N_10581,N_11646);
nor U13080 (N_13080,N_10798,N_12282);
xnor U13081 (N_13081,N_11220,N_11550);
and U13082 (N_13082,N_10202,N_10209);
nor U13083 (N_13083,N_10428,N_11211);
nand U13084 (N_13084,N_10359,N_12398);
and U13085 (N_13085,N_11049,N_11103);
or U13086 (N_13086,N_12419,N_11203);
nor U13087 (N_13087,N_12250,N_11269);
xnor U13088 (N_13088,N_10548,N_11928);
nor U13089 (N_13089,N_11843,N_10162);
or U13090 (N_13090,N_11786,N_11848);
xor U13091 (N_13091,N_11567,N_12104);
xnor U13092 (N_13092,N_10467,N_11095);
or U13093 (N_13093,N_11043,N_12231);
or U13094 (N_13094,N_10694,N_11303);
xnor U13095 (N_13095,N_12384,N_11449);
and U13096 (N_13096,N_11987,N_10831);
and U13097 (N_13097,N_10358,N_11080);
nand U13098 (N_13098,N_11901,N_11925);
nand U13099 (N_13099,N_12361,N_11769);
and U13100 (N_13100,N_12408,N_10983);
xor U13101 (N_13101,N_10705,N_10356);
and U13102 (N_13102,N_10725,N_11363);
nor U13103 (N_13103,N_11177,N_10229);
and U13104 (N_13104,N_10184,N_11116);
or U13105 (N_13105,N_11945,N_11353);
nand U13106 (N_13106,N_11268,N_10127);
and U13107 (N_13107,N_10564,N_10726);
or U13108 (N_13108,N_10787,N_11045);
and U13109 (N_13109,N_10788,N_10870);
xor U13110 (N_13110,N_10306,N_10853);
nand U13111 (N_13111,N_11630,N_11206);
xor U13112 (N_13112,N_11251,N_11734);
nand U13113 (N_13113,N_10990,N_10227);
nor U13114 (N_13114,N_10177,N_10486);
and U13115 (N_13115,N_12260,N_11745);
nand U13116 (N_13116,N_10626,N_12257);
nor U13117 (N_13117,N_12095,N_11959);
nor U13118 (N_13118,N_10283,N_11027);
xor U13119 (N_13119,N_11491,N_11808);
or U13120 (N_13120,N_10763,N_10182);
nor U13121 (N_13121,N_11411,N_10180);
or U13122 (N_13122,N_10860,N_11145);
xor U13123 (N_13123,N_10718,N_11030);
nand U13124 (N_13124,N_10277,N_10584);
xor U13125 (N_13125,N_11271,N_10866);
nor U13126 (N_13126,N_10313,N_12482);
nand U13127 (N_13127,N_12270,N_10897);
or U13128 (N_13128,N_11320,N_10135);
xnor U13129 (N_13129,N_10469,N_10027);
xor U13130 (N_13130,N_12037,N_11937);
nand U13131 (N_13131,N_11512,N_10839);
and U13132 (N_13132,N_11962,N_10654);
and U13133 (N_13133,N_10051,N_10076);
and U13134 (N_13134,N_10646,N_12140);
xnor U13135 (N_13135,N_10559,N_10546);
and U13136 (N_13136,N_12215,N_10402);
xnor U13137 (N_13137,N_12442,N_11934);
and U13138 (N_13138,N_11572,N_10879);
and U13139 (N_13139,N_11328,N_10966);
or U13140 (N_13140,N_12451,N_11242);
nor U13141 (N_13141,N_12362,N_12069);
or U13142 (N_13142,N_11421,N_11939);
nor U13143 (N_13143,N_10192,N_11178);
nand U13144 (N_13144,N_11254,N_11200);
or U13145 (N_13145,N_11574,N_10069);
and U13146 (N_13146,N_11346,N_11963);
and U13147 (N_13147,N_11894,N_12456);
and U13148 (N_13148,N_12448,N_11725);
and U13149 (N_13149,N_11869,N_11915);
and U13150 (N_13150,N_11754,N_12378);
nand U13151 (N_13151,N_11856,N_10883);
or U13152 (N_13152,N_10197,N_12369);
or U13153 (N_13153,N_11614,N_11069);
nor U13154 (N_13154,N_10176,N_12162);
or U13155 (N_13155,N_11497,N_12044);
nor U13156 (N_13156,N_12276,N_10004);
xor U13157 (N_13157,N_10041,N_11496);
and U13158 (N_13158,N_11714,N_11662);
nor U13159 (N_13159,N_11003,N_11712);
and U13160 (N_13160,N_10517,N_10349);
nand U13161 (N_13161,N_11568,N_12248);
nor U13162 (N_13162,N_11898,N_10108);
xor U13163 (N_13163,N_10022,N_12110);
and U13164 (N_13164,N_11751,N_11162);
nor U13165 (N_13165,N_11498,N_12299);
nand U13166 (N_13166,N_11862,N_11056);
nand U13167 (N_13167,N_11172,N_11995);
nor U13168 (N_13168,N_10539,N_12415);
xor U13169 (N_13169,N_10651,N_11094);
or U13170 (N_13170,N_11258,N_11016);
or U13171 (N_13171,N_12189,N_10301);
nand U13172 (N_13172,N_12153,N_11830);
or U13173 (N_13173,N_11333,N_11345);
nand U13174 (N_13174,N_11998,N_11114);
nor U13175 (N_13175,N_12264,N_11605);
nor U13176 (N_13176,N_11479,N_11680);
or U13177 (N_13177,N_10814,N_10709);
nand U13178 (N_13178,N_10872,N_10070);
or U13179 (N_13179,N_11074,N_10621);
and U13180 (N_13180,N_11106,N_11695);
nand U13181 (N_13181,N_12455,N_11367);
and U13182 (N_13182,N_12249,N_10686);
and U13183 (N_13183,N_10906,N_11071);
or U13184 (N_13184,N_11850,N_12289);
nand U13185 (N_13185,N_11598,N_12290);
nand U13186 (N_13186,N_10189,N_11819);
xor U13187 (N_13187,N_11040,N_12040);
or U13188 (N_13188,N_10600,N_12108);
xnor U13189 (N_13189,N_11668,N_10893);
xor U13190 (N_13190,N_10246,N_10930);
nand U13191 (N_13191,N_11814,N_11596);
xor U13192 (N_13192,N_11761,N_10784);
or U13193 (N_13193,N_10478,N_11949);
and U13194 (N_13194,N_11519,N_11990);
and U13195 (N_13195,N_10869,N_11579);
xnor U13196 (N_13196,N_10280,N_10498);
nand U13197 (N_13197,N_10741,N_11569);
xnor U13198 (N_13198,N_12143,N_10094);
nor U13199 (N_13199,N_11641,N_12063);
nand U13200 (N_13200,N_11506,N_11418);
or U13201 (N_13201,N_10011,N_11188);
or U13202 (N_13202,N_11397,N_10894);
or U13203 (N_13203,N_10077,N_11156);
xnor U13204 (N_13204,N_12432,N_10541);
xnor U13205 (N_13205,N_10112,N_11561);
nor U13206 (N_13206,N_12129,N_10758);
and U13207 (N_13207,N_10817,N_10460);
xnor U13208 (N_13208,N_10249,N_12352);
and U13209 (N_13209,N_11087,N_12135);
nand U13210 (N_13210,N_12251,N_10106);
xnor U13211 (N_13211,N_11192,N_10420);
and U13212 (N_13212,N_12255,N_11157);
nand U13213 (N_13213,N_10729,N_11347);
or U13214 (N_13214,N_11717,N_12252);
or U13215 (N_13215,N_11691,N_11291);
nand U13216 (N_13216,N_11480,N_11903);
and U13217 (N_13217,N_10087,N_12192);
and U13218 (N_13218,N_12150,N_10468);
nor U13219 (N_13219,N_10778,N_10852);
xor U13220 (N_13220,N_10804,N_11729);
nand U13221 (N_13221,N_11412,N_10912);
nand U13222 (N_13222,N_10008,N_10326);
nand U13223 (N_13223,N_11135,N_11863);
or U13224 (N_13224,N_11120,N_11463);
or U13225 (N_13225,N_11337,N_11676);
xor U13226 (N_13226,N_11277,N_11528);
nand U13227 (N_13227,N_10873,N_11127);
or U13228 (N_13228,N_10532,N_11979);
and U13229 (N_13229,N_10082,N_11697);
nor U13230 (N_13230,N_12032,N_10304);
nand U13231 (N_13231,N_12072,N_11201);
nand U13232 (N_13232,N_11439,N_12167);
nor U13233 (N_13233,N_10090,N_10697);
and U13234 (N_13234,N_12379,N_11323);
nor U13235 (N_13235,N_10114,N_10147);
or U13236 (N_13236,N_11325,N_11687);
xor U13237 (N_13237,N_10953,N_11887);
and U13238 (N_13238,N_11637,N_12035);
nor U13239 (N_13239,N_11119,N_10510);
and U13240 (N_13240,N_12464,N_10490);
nand U13241 (N_13241,N_11374,N_12138);
nand U13242 (N_13242,N_11952,N_10435);
or U13243 (N_13243,N_11058,N_11760);
and U13244 (N_13244,N_10118,N_10059);
nor U13245 (N_13245,N_11141,N_11093);
and U13246 (N_13246,N_10307,N_12300);
nor U13247 (N_13247,N_11286,N_10805);
or U13248 (N_13248,N_10335,N_10608);
and U13249 (N_13249,N_12241,N_11684);
xnor U13250 (N_13250,N_10685,N_11759);
or U13251 (N_13251,N_10047,N_11429);
and U13252 (N_13252,N_11926,N_12160);
and U13253 (N_13253,N_12465,N_11299);
nand U13254 (N_13254,N_12230,N_11236);
or U13255 (N_13255,N_11927,N_10441);
xnor U13256 (N_13256,N_10670,N_11823);
or U13257 (N_13257,N_10243,N_11876);
nand U13258 (N_13258,N_10768,N_11247);
or U13259 (N_13259,N_11704,N_11215);
nor U13260 (N_13260,N_11578,N_11991);
or U13261 (N_13261,N_12453,N_12314);
or U13262 (N_13262,N_10881,N_10170);
xor U13263 (N_13263,N_12367,N_10846);
nand U13264 (N_13264,N_12452,N_12306);
and U13265 (N_13265,N_12329,N_10150);
nand U13266 (N_13266,N_11276,N_11798);
and U13267 (N_13267,N_12177,N_11772);
and U13268 (N_13268,N_11656,N_10851);
and U13269 (N_13269,N_12430,N_11376);
xor U13270 (N_13270,N_12026,N_11777);
nand U13271 (N_13271,N_12393,N_10823);
xor U13272 (N_13272,N_11034,N_11310);
and U13273 (N_13273,N_12024,N_11490);
nor U13274 (N_13274,N_11315,N_12001);
or U13275 (N_13275,N_11816,N_10858);
xnor U13276 (N_13276,N_11661,N_10767);
or U13277 (N_13277,N_11226,N_11246);
nand U13278 (N_13278,N_10312,N_11072);
nor U13279 (N_13279,N_11601,N_10290);
and U13280 (N_13280,N_12182,N_10085);
xnor U13281 (N_13281,N_11110,N_10835);
nand U13282 (N_13282,N_11750,N_10099);
nand U13283 (N_13283,N_10789,N_11499);
xor U13284 (N_13284,N_11733,N_10021);
nand U13285 (N_13285,N_11026,N_10813);
xor U13286 (N_13286,N_10558,N_12087);
or U13287 (N_13287,N_11306,N_10972);
nor U13288 (N_13288,N_11160,N_11681);
or U13289 (N_13289,N_10610,N_10084);
nor U13290 (N_13290,N_12117,N_10092);
nor U13291 (N_13291,N_10702,N_10588);
nand U13292 (N_13292,N_12385,N_10336);
and U13293 (N_13293,N_10769,N_12130);
nand U13294 (N_13294,N_12380,N_11781);
nand U13295 (N_13295,N_11996,N_11041);
or U13296 (N_13296,N_10520,N_11543);
xnor U13297 (N_13297,N_10830,N_11529);
or U13298 (N_13298,N_11244,N_11683);
and U13299 (N_13299,N_10001,N_11235);
nand U13300 (N_13300,N_12041,N_10514);
or U13301 (N_13301,N_11739,N_10772);
nor U13302 (N_13302,N_10408,N_11594);
and U13303 (N_13303,N_10834,N_11105);
or U13304 (N_13304,N_12176,N_10864);
or U13305 (N_13305,N_10876,N_11820);
and U13306 (N_13306,N_10956,N_10880);
and U13307 (N_13307,N_11768,N_11839);
xnor U13308 (N_13308,N_11403,N_10395);
nand U13309 (N_13309,N_10199,N_10613);
nand U13310 (N_13310,N_10755,N_12067);
nor U13311 (N_13311,N_11307,N_11548);
nand U13312 (N_13312,N_10590,N_11062);
xnor U13313 (N_13313,N_12125,N_10779);
nor U13314 (N_13314,N_12435,N_10856);
nor U13315 (N_13315,N_10012,N_12029);
nand U13316 (N_13316,N_11974,N_10737);
xnor U13317 (N_13317,N_11648,N_11329);
and U13318 (N_13318,N_10000,N_10607);
or U13319 (N_13319,N_11728,N_11600);
and U13320 (N_13320,N_10736,N_11692);
nand U13321 (N_13321,N_11278,N_10742);
xnor U13322 (N_13322,N_10620,N_11343);
xor U13323 (N_13323,N_11921,N_11126);
and U13324 (N_13324,N_11392,N_11741);
nand U13325 (N_13325,N_10850,N_10086);
xnor U13326 (N_13326,N_11252,N_10699);
nor U13327 (N_13327,N_11447,N_12391);
nand U13328 (N_13328,N_12350,N_12200);
or U13329 (N_13329,N_10125,N_12499);
and U13330 (N_13330,N_11128,N_10236);
or U13331 (N_13331,N_10781,N_10452);
nand U13332 (N_13332,N_10566,N_10096);
and U13333 (N_13333,N_10221,N_11185);
nand U13334 (N_13334,N_10993,N_11179);
or U13335 (N_13335,N_10233,N_10770);
and U13336 (N_13336,N_10945,N_11124);
and U13337 (N_13337,N_11744,N_11084);
nor U13338 (N_13338,N_11965,N_11233);
or U13339 (N_13339,N_11737,N_10542);
or U13340 (N_13340,N_11099,N_11327);
nor U13341 (N_13341,N_10384,N_10322);
and U13342 (N_13342,N_10703,N_11670);
xnor U13343 (N_13343,N_11012,N_11428);
xor U13344 (N_13344,N_12198,N_11972);
nor U13345 (N_13345,N_11608,N_10704);
nor U13346 (N_13346,N_10267,N_10284);
or U13347 (N_13347,N_12131,N_10752);
nor U13348 (N_13348,N_10681,N_10164);
nor U13349 (N_13349,N_10698,N_10832);
nor U13350 (N_13350,N_11471,N_11967);
nor U13351 (N_13351,N_10081,N_11446);
nand U13352 (N_13352,N_10375,N_11482);
and U13353 (N_13353,N_10128,N_11532);
xnor U13354 (N_13354,N_12085,N_10824);
nand U13355 (N_13355,N_10257,N_12287);
nor U13356 (N_13356,N_10231,N_11749);
nand U13357 (N_13357,N_11885,N_11011);
or U13358 (N_13358,N_11736,N_10687);
and U13359 (N_13359,N_11199,N_10035);
xnor U13360 (N_13360,N_12184,N_11763);
nor U13361 (N_13361,N_12163,N_12414);
nand U13362 (N_13362,N_11638,N_10501);
nor U13363 (N_13363,N_11152,N_10214);
nor U13364 (N_13364,N_10353,N_10371);
and U13365 (N_13365,N_10291,N_10863);
nor U13366 (N_13366,N_10888,N_10913);
nand U13367 (N_13367,N_10557,N_11999);
nand U13368 (N_13368,N_11191,N_11539);
or U13369 (N_13369,N_11966,N_11284);
xnor U13370 (N_13370,N_10734,N_12416);
or U13371 (N_13371,N_10279,N_10190);
xor U13372 (N_13372,N_10278,N_11331);
nor U13373 (N_13373,N_10213,N_11282);
or U13374 (N_13374,N_10509,N_12256);
or U13375 (N_13375,N_11886,N_12490);
nor U13376 (N_13376,N_11988,N_11629);
nand U13377 (N_13377,N_10260,N_12157);
nand U13378 (N_13378,N_10488,N_11488);
nor U13379 (N_13379,N_10451,N_10196);
and U13380 (N_13380,N_11643,N_11168);
xor U13381 (N_13381,N_12439,N_10754);
nand U13382 (N_13382,N_12210,N_11560);
or U13383 (N_13383,N_10896,N_12091);
and U13384 (N_13384,N_10657,N_12274);
xnor U13385 (N_13385,N_11461,N_10049);
nand U13386 (N_13386,N_11660,N_12159);
or U13387 (N_13387,N_12258,N_12468);
and U13388 (N_13388,N_10009,N_12064);
and U13389 (N_13389,N_10589,N_10503);
xor U13390 (N_13390,N_11904,N_10747);
or U13391 (N_13391,N_10961,N_11048);
xnor U13392 (N_13392,N_10673,N_11602);
nor U13393 (N_13393,N_11950,N_12004);
nor U13394 (N_13394,N_11270,N_12263);
nand U13395 (N_13395,N_11649,N_10296);
nor U13396 (N_13396,N_10365,N_11982);
and U13397 (N_13397,N_10450,N_11351);
nand U13398 (N_13398,N_10230,N_12146);
xnor U13399 (N_13399,N_11300,N_11086);
and U13400 (N_13400,N_11653,N_11475);
xnor U13401 (N_13401,N_12433,N_11835);
nor U13402 (N_13402,N_12059,N_10898);
or U13403 (N_13403,N_11797,N_11210);
nand U13404 (N_13404,N_11010,N_12411);
nor U13405 (N_13405,N_11755,N_10083);
and U13406 (N_13406,N_11774,N_11493);
nor U13407 (N_13407,N_10507,N_10437);
xor U13408 (N_13408,N_10242,N_10695);
xor U13409 (N_13409,N_10901,N_11563);
and U13410 (N_13410,N_10330,N_11690);
xor U13411 (N_13411,N_12062,N_11039);
or U13412 (N_13412,N_10890,N_11064);
nand U13413 (N_13413,N_10795,N_11054);
xor U13414 (N_13414,N_10471,N_12463);
or U13415 (N_13415,N_10276,N_10771);
or U13416 (N_13416,N_11239,N_12030);
nor U13417 (N_13417,N_11024,N_12297);
nand U13418 (N_13418,N_11228,N_11202);
or U13419 (N_13419,N_10374,N_11902);
and U13420 (N_13420,N_12461,N_10535);
nor U13421 (N_13421,N_11708,N_11773);
nor U13422 (N_13422,N_10025,N_10425);
and U13423 (N_13423,N_11441,N_11922);
xor U13424 (N_13424,N_11473,N_10959);
or U13425 (N_13425,N_12100,N_10533);
or U13426 (N_13426,N_12336,N_10738);
and U13427 (N_13427,N_12123,N_12347);
and U13428 (N_13428,N_11795,N_11008);
and U13429 (N_13429,N_11077,N_10944);
xor U13430 (N_13430,N_12178,N_10537);
nor U13431 (N_13431,N_11394,N_11019);
nor U13432 (N_13432,N_10405,N_11240);
or U13433 (N_13433,N_10295,N_11562);
and U13434 (N_13434,N_12431,N_10571);
and U13435 (N_13435,N_11338,N_11723);
or U13436 (N_13436,N_11613,N_10745);
xnor U13437 (N_13437,N_10193,N_10633);
nor U13438 (N_13438,N_10701,N_11279);
or U13439 (N_13439,N_10188,N_11318);
nand U13440 (N_13440,N_11503,N_11906);
nand U13441 (N_13441,N_11020,N_12386);
or U13442 (N_13442,N_12174,N_12050);
or U13443 (N_13443,N_11696,N_10978);
nor U13444 (N_13444,N_10582,N_12124);
nor U13445 (N_13445,N_12054,N_10352);
nand U13446 (N_13446,N_11542,N_11231);
or U13447 (N_13447,N_12450,N_10665);
nand U13448 (N_13448,N_11386,N_12213);
and U13449 (N_13449,N_11829,N_11151);
xnor U13450 (N_13450,N_10415,N_12243);
nor U13451 (N_13451,N_12151,N_11289);
xnor U13452 (N_13452,N_12373,N_12014);
nand U13453 (N_13453,N_11511,N_12372);
and U13454 (N_13454,N_10977,N_11698);
nand U13455 (N_13455,N_10299,N_10829);
xor U13456 (N_13456,N_10394,N_10042);
xnor U13457 (N_13457,N_10712,N_11399);
nor U13458 (N_13458,N_10991,N_11824);
nand U13459 (N_13459,N_11558,N_10518);
xor U13460 (N_13460,N_11620,N_10521);
nand U13461 (N_13461,N_10647,N_11564);
nor U13462 (N_13462,N_10476,N_11948);
nand U13463 (N_13463,N_10139,N_11414);
xnor U13464 (N_13464,N_11626,N_10343);
xnor U13465 (N_13465,N_10914,N_10920);
or U13466 (N_13466,N_10545,N_10339);
nand U13467 (N_13467,N_10217,N_11545);
or U13468 (N_13468,N_11855,N_10195);
nor U13469 (N_13469,N_12028,N_11171);
nand U13470 (N_13470,N_12392,N_10578);
nor U13471 (N_13471,N_11433,N_11450);
and U13472 (N_13472,N_10281,N_12098);
and U13473 (N_13473,N_12022,N_12283);
xnor U13474 (N_13474,N_11810,N_11335);
or U13475 (N_13475,N_10562,N_12003);
xnor U13476 (N_13476,N_10207,N_11718);
nand U13477 (N_13477,N_12327,N_12261);
nand U13478 (N_13478,N_11610,N_10238);
nand U13479 (N_13479,N_11312,N_11342);
nand U13480 (N_13480,N_11007,N_11525);
and U13481 (N_13481,N_12496,N_12356);
xnor U13482 (N_13482,N_11993,N_10033);
nand U13483 (N_13483,N_11977,N_10609);
and U13484 (N_13484,N_11314,N_11184);
xor U13485 (N_13485,N_11322,N_10430);
nand U13486 (N_13486,N_12019,N_12363);
xnor U13487 (N_13487,N_12348,N_10572);
and U13488 (N_13488,N_10668,N_12404);
xnor U13489 (N_13489,N_10018,N_12285);
or U13490 (N_13490,N_11207,N_10563);
or U13491 (N_13491,N_10487,N_11142);
nand U13492 (N_13492,N_11960,N_10285);
nor U13493 (N_13493,N_12074,N_10057);
xor U13494 (N_13494,N_11067,N_10347);
nand U13495 (N_13495,N_10413,N_10998);
nor U13496 (N_13496,N_11870,N_10965);
nor U13497 (N_13497,N_11591,N_11884);
and U13498 (N_13498,N_10997,N_11847);
or U13499 (N_13499,N_11182,N_12171);
nor U13500 (N_13500,N_11319,N_12039);
xnor U13501 (N_13501,N_10815,N_12203);
xor U13502 (N_13502,N_10443,N_12457);
nor U13503 (N_13503,N_10710,N_11770);
xor U13504 (N_13504,N_11422,N_11909);
nand U13505 (N_13505,N_11664,N_11757);
nor U13506 (N_13506,N_10232,N_11711);
nor U13507 (N_13507,N_12381,N_11298);
nor U13508 (N_13508,N_10943,N_10689);
nand U13509 (N_13509,N_10567,N_10416);
nor U13510 (N_13510,N_11170,N_10429);
xor U13511 (N_13511,N_11900,N_11920);
nand U13512 (N_13512,N_10596,N_10838);
nand U13513 (N_13513,N_10362,N_10806);
nand U13514 (N_13514,N_10294,N_12234);
or U13515 (N_13515,N_11895,N_12308);
or U13516 (N_13516,N_12493,N_10496);
or U13517 (N_13517,N_10289,N_10050);
nand U13518 (N_13518,N_11796,N_12088);
nor U13519 (N_13519,N_10145,N_11509);
and U13520 (N_13520,N_11065,N_11992);
or U13521 (N_13521,N_11474,N_11631);
or U13522 (N_13522,N_10783,N_11837);
nor U13523 (N_13523,N_10777,N_12020);
or U13524 (N_13524,N_11001,N_11775);
and U13525 (N_13525,N_10095,N_10156);
and U13526 (N_13526,N_12443,N_10812);
or U13527 (N_13527,N_10825,N_11456);
nor U13528 (N_13528,N_11546,N_11297);
or U13529 (N_13529,N_10963,N_11584);
xor U13530 (N_13530,N_12279,N_11495);
nand U13531 (N_13531,N_11807,N_11267);
xnor U13532 (N_13532,N_11913,N_10269);
or U13533 (N_13533,N_10398,N_10717);
nor U13534 (N_13534,N_10996,N_10743);
and U13535 (N_13535,N_12469,N_10066);
xor U13536 (N_13536,N_12149,N_12043);
and U13537 (N_13537,N_12394,N_10401);
or U13538 (N_13538,N_10765,N_12355);
or U13539 (N_13539,N_10252,N_11406);
xnor U13540 (N_13540,N_10502,N_10438);
nand U13541 (N_13541,N_11580,N_11304);
xnor U13542 (N_13542,N_10153,N_10102);
xor U13543 (N_13543,N_11735,N_11924);
xor U13544 (N_13544,N_11000,N_10015);
or U13545 (N_13545,N_10411,N_11381);
or U13546 (N_13546,N_12396,N_11997);
and U13547 (N_13547,N_12341,N_12337);
xor U13548 (N_13548,N_12476,N_12023);
nand U13549 (N_13549,N_10038,N_10489);
and U13550 (N_13550,N_11405,N_10624);
and U13551 (N_13551,N_10414,N_11505);
nand U13552 (N_13552,N_11485,N_10154);
nor U13553 (N_13553,N_10649,N_10204);
nand U13554 (N_13554,N_12491,N_12016);
or U13555 (N_13555,N_11248,N_10583);
and U13556 (N_13556,N_11190,N_11861);
or U13557 (N_13557,N_11222,N_10644);
or U13558 (N_13558,N_10964,N_10455);
nand U13559 (N_13559,N_10166,N_12335);
and U13560 (N_13560,N_12114,N_11379);
xnor U13561 (N_13561,N_11540,N_10160);
or U13562 (N_13562,N_12244,N_12318);
xor U13563 (N_13563,N_12413,N_10931);
nand U13564 (N_13564,N_12073,N_10603);
nor U13565 (N_13565,N_10919,N_10119);
and U13566 (N_13566,N_11091,N_11693);
nand U13567 (N_13567,N_11940,N_11688);
and U13568 (N_13568,N_10739,N_11719);
and U13569 (N_13569,N_10409,N_11806);
or U13570 (N_13570,N_10005,N_11225);
xnor U13571 (N_13571,N_10653,N_10617);
or U13572 (N_13572,N_12083,N_10599);
or U13573 (N_13573,N_10474,N_12365);
nor U13574 (N_13574,N_11957,N_11301);
nor U13575 (N_13575,N_11057,N_11458);
or U13576 (N_13576,N_12077,N_11453);
and U13577 (N_13577,N_12206,N_11844);
nand U13578 (N_13578,N_11365,N_11154);
and U13579 (N_13579,N_12223,N_10381);
xor U13580 (N_13580,N_10615,N_10632);
xor U13581 (N_13581,N_12132,N_12209);
or U13582 (N_13582,N_11645,N_12296);
xnor U13583 (N_13583,N_10544,N_12390);
and U13584 (N_13584,N_10377,N_11813);
nor U13585 (N_13585,N_10029,N_10902);
nand U13586 (N_13586,N_10259,N_11424);
nand U13587 (N_13587,N_11958,N_10036);
xnor U13588 (N_13588,N_11907,N_12057);
nand U13589 (N_13589,N_11933,N_10482);
or U13590 (N_13590,N_11036,N_10044);
nand U13591 (N_13591,N_11098,N_11038);
and U13592 (N_13592,N_10448,N_10032);
or U13593 (N_13593,N_10802,N_11606);
nor U13594 (N_13594,N_12103,N_10948);
or U13595 (N_13595,N_11330,N_12008);
nand U13596 (N_13596,N_10007,N_10722);
or U13597 (N_13597,N_10538,N_10212);
or U13598 (N_13598,N_10887,N_12161);
and U13599 (N_13599,N_12034,N_10423);
nor U13600 (N_13600,N_12021,N_12328);
xnor U13601 (N_13601,N_11362,N_10433);
xnor U13602 (N_13602,N_10271,N_11378);
and U13603 (N_13603,N_11767,N_10323);
nor U13604 (N_13604,N_11469,N_12006);
nor U13605 (N_13605,N_10989,N_10334);
and U13606 (N_13606,N_10504,N_11616);
nand U13607 (N_13607,N_10383,N_10713);
or U13608 (N_13608,N_12027,N_11818);
xor U13609 (N_13609,N_12052,N_12164);
xor U13610 (N_13610,N_12487,N_12311);
nand U13611 (N_13611,N_10892,N_11018);
and U13612 (N_13612,N_10659,N_11109);
xnor U13613 (N_13613,N_11951,N_10554);
nand U13614 (N_13614,N_12291,N_10447);
nor U13615 (N_13615,N_10748,N_10648);
and U13616 (N_13616,N_10568,N_12262);
nor U13617 (N_13617,N_11932,N_11445);
xor U13618 (N_13618,N_11205,N_11809);
and U13619 (N_13619,N_10875,N_11888);
nor U13620 (N_13620,N_11859,N_10667);
or U13621 (N_13621,N_11526,N_11658);
nor U13622 (N_13622,N_10072,N_10994);
nor U13623 (N_13623,N_12259,N_11815);
nand U13624 (N_13624,N_11173,N_10519);
nand U13625 (N_13625,N_10324,N_11617);
xnor U13626 (N_13626,N_10934,N_10984);
and U13627 (N_13627,N_10315,N_10837);
or U13628 (N_13628,N_12334,N_10848);
nor U13629 (N_13629,N_11263,N_12112);
xnor U13630 (N_13630,N_11897,N_11355);
xnor U13631 (N_13631,N_10303,N_11935);
or U13632 (N_13632,N_11336,N_10759);
nand U13633 (N_13633,N_11175,N_11947);
nand U13634 (N_13634,N_11344,N_11971);
nand U13635 (N_13635,N_11075,N_10719);
or U13636 (N_13636,N_11159,N_12237);
xnor U13637 (N_13637,N_10973,N_11257);
and U13638 (N_13638,N_11612,N_11389);
nand U13639 (N_13639,N_11507,N_11464);
nor U13640 (N_13640,N_12370,N_11467);
nor U13641 (N_13641,N_10962,N_10045);
or U13642 (N_13642,N_10338,N_10570);
and U13643 (N_13643,N_11032,N_12002);
nor U13644 (N_13644,N_10512,N_10939);
nor U13645 (N_13645,N_10884,N_12494);
nor U13646 (N_13646,N_10855,N_10797);
and U13647 (N_13647,N_11537,N_10040);
xnor U13648 (N_13648,N_10844,N_11802);
or U13649 (N_13649,N_12424,N_11189);
xnor U13650 (N_13650,N_10372,N_12081);
or U13651 (N_13651,N_11544,N_10732);
nor U13652 (N_13652,N_12286,N_11125);
nor U13653 (N_13653,N_10210,N_10256);
xnor U13654 (N_13654,N_10935,N_12137);
nand U13655 (N_13655,N_10062,N_12166);
or U13656 (N_13656,N_11980,N_10674);
nand U13657 (N_13657,N_12238,N_10361);
or U13658 (N_13658,N_10547,N_11398);
and U13659 (N_13659,N_10350,N_10749);
nand U13660 (N_13660,N_11250,N_10121);
nand U13661 (N_13661,N_11911,N_10911);
and U13662 (N_13662,N_11204,N_10071);
nand U13663 (N_13663,N_12488,N_10979);
nor U13664 (N_13664,N_11042,N_11672);
xor U13665 (N_13665,N_12273,N_11423);
xor U13666 (N_13666,N_10403,N_10329);
and U13667 (N_13667,N_11261,N_11522);
nor U13668 (N_13668,N_10505,N_12065);
xnor U13669 (N_13669,N_11358,N_11465);
or U13670 (N_13670,N_10634,N_10925);
xnor U13671 (N_13671,N_12474,N_10843);
nand U13672 (N_13672,N_10237,N_10037);
xnor U13673 (N_13673,N_10585,N_11223);
or U13674 (N_13674,N_10308,N_10293);
xnor U13675 (N_13675,N_10862,N_11881);
xor U13676 (N_13676,N_12364,N_10847);
nor U13677 (N_13677,N_10178,N_11195);
nor U13678 (N_13678,N_10819,N_11383);
nand U13679 (N_13679,N_12168,N_11551);
nor U13680 (N_13680,N_10165,N_11659);
xnor U13681 (N_13681,N_10952,N_12410);
and U13682 (N_13682,N_10442,N_10239);
or U13683 (N_13683,N_11425,N_12358);
and U13684 (N_13684,N_10060,N_11743);
nor U13685 (N_13685,N_10026,N_11686);
xor U13686 (N_13686,N_10652,N_10133);
nor U13687 (N_13687,N_11520,N_11970);
nand U13688 (N_13688,N_10124,N_10399);
xor U13689 (N_13689,N_10904,N_10550);
or U13690 (N_13690,N_11575,N_11006);
or U13691 (N_13691,N_10483,N_10499);
nand U13692 (N_13692,N_12247,N_11133);
nor U13693 (N_13693,N_12440,N_12418);
nor U13694 (N_13694,N_11538,N_12005);
and U13695 (N_13695,N_11654,N_10459);
nand U13696 (N_13696,N_11746,N_11092);
or U13697 (N_13697,N_12275,N_11789);
nor U13698 (N_13698,N_10132,N_12400);
nor U13699 (N_13699,N_10458,N_10175);
or U13700 (N_13700,N_11395,N_11492);
or U13701 (N_13701,N_11675,N_10406);
or U13702 (N_13702,N_12010,N_12472);
nand U13703 (N_13703,N_12195,N_10089);
and U13704 (N_13704,N_12134,N_11140);
nand U13705 (N_13705,N_11391,N_12471);
nand U13706 (N_13706,N_10109,N_12096);
nand U13707 (N_13707,N_11035,N_11265);
or U13708 (N_13708,N_12303,N_11941);
or U13709 (N_13709,N_12434,N_11872);
or U13710 (N_13710,N_11953,N_11699);
nand U13711 (N_13711,N_12101,N_11871);
and U13712 (N_13712,N_11731,N_10396);
nand U13713 (N_13713,N_12332,N_10690);
or U13714 (N_13714,N_10899,N_10412);
and U13715 (N_13715,N_12186,N_11232);
nor U13716 (N_13716,N_11308,N_11264);
or U13717 (N_13717,N_12284,N_10774);
nand U13718 (N_13718,N_12170,N_11166);
xnor U13719 (N_13719,N_10688,N_12047);
nor U13720 (N_13720,N_11366,N_11530);
and U13721 (N_13721,N_11964,N_11825);
nor U13722 (N_13722,N_11666,N_11576);
and U13723 (N_13723,N_11912,N_10250);
nand U13724 (N_13724,N_10602,N_10316);
nand U13725 (N_13725,N_11671,N_11782);
nand U13726 (N_13726,N_10707,N_11930);
and U13727 (N_13727,N_10472,N_11713);
and U13728 (N_13728,N_12395,N_12459);
nor U13729 (N_13729,N_11382,N_11776);
or U13730 (N_13730,N_10730,N_11321);
nor U13731 (N_13731,N_11732,N_10319);
nand U13732 (N_13732,N_11976,N_11555);
and U13733 (N_13733,N_10598,N_10639);
nor U13734 (N_13734,N_10493,N_11044);
nor U13735 (N_13735,N_10995,N_10500);
or U13736 (N_13736,N_10161,N_11169);
nand U13737 (N_13737,N_12193,N_10439);
nor U13738 (N_13738,N_11557,N_11288);
nand U13739 (N_13739,N_11138,N_12045);
nor U13740 (N_13740,N_10982,N_11747);
nand U13741 (N_13741,N_11436,N_11448);
or U13742 (N_13742,N_11627,N_10810);
and U13743 (N_13743,N_10908,N_11387);
or U13744 (N_13744,N_10776,N_12428);
and U13745 (N_13745,N_12048,N_11685);
or U13746 (N_13746,N_10561,N_10054);
and U13747 (N_13747,N_12197,N_11730);
xor U13748 (N_13748,N_10470,N_11779);
nor U13749 (N_13749,N_12454,N_10426);
nor U13750 (N_13750,N_10048,N_11504);
and U13751 (N_13751,N_11134,N_10929);
or U13752 (N_13752,N_11121,N_10383);
or U13753 (N_13753,N_12132,N_12038);
and U13754 (N_13754,N_11995,N_10566);
xnor U13755 (N_13755,N_11895,N_10635);
nor U13756 (N_13756,N_11188,N_10318);
xnor U13757 (N_13757,N_10363,N_11554);
or U13758 (N_13758,N_10391,N_10760);
nand U13759 (N_13759,N_10122,N_11709);
nor U13760 (N_13760,N_11503,N_10763);
nor U13761 (N_13761,N_10995,N_11975);
nand U13762 (N_13762,N_10969,N_11312);
and U13763 (N_13763,N_12385,N_10786);
nor U13764 (N_13764,N_10971,N_11151);
xor U13765 (N_13765,N_10911,N_11878);
nand U13766 (N_13766,N_12036,N_12254);
nand U13767 (N_13767,N_11724,N_11864);
xnor U13768 (N_13768,N_12379,N_11027);
nor U13769 (N_13769,N_11322,N_12011);
xor U13770 (N_13770,N_12359,N_11847);
xnor U13771 (N_13771,N_10657,N_10718);
and U13772 (N_13772,N_11513,N_12440);
and U13773 (N_13773,N_10932,N_11721);
or U13774 (N_13774,N_10713,N_11337);
and U13775 (N_13775,N_12109,N_11757);
or U13776 (N_13776,N_10813,N_11876);
and U13777 (N_13777,N_10922,N_12051);
or U13778 (N_13778,N_10114,N_10427);
and U13779 (N_13779,N_10231,N_10080);
and U13780 (N_13780,N_11037,N_10256);
and U13781 (N_13781,N_10509,N_10974);
and U13782 (N_13782,N_10188,N_10941);
and U13783 (N_13783,N_12456,N_12113);
nand U13784 (N_13784,N_10033,N_10991);
or U13785 (N_13785,N_11408,N_11868);
and U13786 (N_13786,N_10810,N_10742);
and U13787 (N_13787,N_11090,N_12108);
nor U13788 (N_13788,N_11868,N_11005);
nand U13789 (N_13789,N_11205,N_11984);
nand U13790 (N_13790,N_10396,N_12278);
nand U13791 (N_13791,N_11628,N_10950);
and U13792 (N_13792,N_11903,N_12472);
and U13793 (N_13793,N_10700,N_12004);
nand U13794 (N_13794,N_11060,N_10815);
or U13795 (N_13795,N_10402,N_12284);
xor U13796 (N_13796,N_12151,N_10084);
and U13797 (N_13797,N_11847,N_10696);
or U13798 (N_13798,N_12495,N_10548);
nand U13799 (N_13799,N_10128,N_11654);
xnor U13800 (N_13800,N_10485,N_11030);
and U13801 (N_13801,N_10773,N_11356);
or U13802 (N_13802,N_10680,N_11076);
xnor U13803 (N_13803,N_11114,N_10743);
nand U13804 (N_13804,N_12366,N_11100);
nand U13805 (N_13805,N_10039,N_10356);
or U13806 (N_13806,N_10747,N_11003);
and U13807 (N_13807,N_10776,N_11606);
nor U13808 (N_13808,N_11220,N_10171);
or U13809 (N_13809,N_12499,N_11733);
and U13810 (N_13810,N_11385,N_10729);
nor U13811 (N_13811,N_11296,N_11854);
or U13812 (N_13812,N_10881,N_12085);
nand U13813 (N_13813,N_10305,N_12295);
xnor U13814 (N_13814,N_10846,N_11849);
xor U13815 (N_13815,N_11187,N_10124);
nor U13816 (N_13816,N_10873,N_10897);
nand U13817 (N_13817,N_11524,N_11882);
and U13818 (N_13818,N_10614,N_11205);
nor U13819 (N_13819,N_10943,N_10480);
and U13820 (N_13820,N_12009,N_11492);
xor U13821 (N_13821,N_10684,N_12057);
or U13822 (N_13822,N_10787,N_11942);
nor U13823 (N_13823,N_10123,N_11448);
xnor U13824 (N_13824,N_12145,N_10085);
xnor U13825 (N_13825,N_10287,N_10522);
and U13826 (N_13826,N_11416,N_10672);
nor U13827 (N_13827,N_12400,N_11588);
xor U13828 (N_13828,N_11369,N_10721);
nand U13829 (N_13829,N_11821,N_11736);
nor U13830 (N_13830,N_10482,N_11843);
xnor U13831 (N_13831,N_10108,N_12143);
and U13832 (N_13832,N_12118,N_11729);
nand U13833 (N_13833,N_12485,N_11163);
nand U13834 (N_13834,N_11609,N_10658);
or U13835 (N_13835,N_11728,N_11855);
nor U13836 (N_13836,N_12495,N_10509);
xor U13837 (N_13837,N_11446,N_10608);
or U13838 (N_13838,N_10492,N_12077);
nor U13839 (N_13839,N_11328,N_11685);
nor U13840 (N_13840,N_10420,N_11980);
nor U13841 (N_13841,N_11916,N_10449);
nor U13842 (N_13842,N_12224,N_11209);
and U13843 (N_13843,N_11948,N_10017);
nand U13844 (N_13844,N_10598,N_11292);
nor U13845 (N_13845,N_12033,N_12292);
nand U13846 (N_13846,N_11933,N_12492);
or U13847 (N_13847,N_10277,N_11512);
xnor U13848 (N_13848,N_12227,N_12063);
and U13849 (N_13849,N_11539,N_12058);
nand U13850 (N_13850,N_10328,N_10703);
and U13851 (N_13851,N_12051,N_12080);
or U13852 (N_13852,N_11949,N_11164);
and U13853 (N_13853,N_12245,N_10072);
nor U13854 (N_13854,N_10847,N_10999);
nand U13855 (N_13855,N_11863,N_10450);
or U13856 (N_13856,N_12183,N_12206);
and U13857 (N_13857,N_11362,N_11105);
nor U13858 (N_13858,N_10342,N_11749);
or U13859 (N_13859,N_12014,N_10650);
xnor U13860 (N_13860,N_10351,N_10759);
nand U13861 (N_13861,N_10212,N_11028);
nor U13862 (N_13862,N_12144,N_10287);
nor U13863 (N_13863,N_10920,N_10693);
xnor U13864 (N_13864,N_11090,N_11283);
nand U13865 (N_13865,N_10492,N_12106);
xnor U13866 (N_13866,N_11026,N_12190);
xor U13867 (N_13867,N_11307,N_10673);
nor U13868 (N_13868,N_12250,N_12216);
nor U13869 (N_13869,N_12347,N_11715);
nor U13870 (N_13870,N_10961,N_11277);
and U13871 (N_13871,N_10805,N_10872);
or U13872 (N_13872,N_12193,N_10184);
xnor U13873 (N_13873,N_11008,N_11946);
nand U13874 (N_13874,N_10513,N_10776);
nor U13875 (N_13875,N_11731,N_11318);
nor U13876 (N_13876,N_10143,N_11246);
xor U13877 (N_13877,N_11122,N_10953);
xor U13878 (N_13878,N_12235,N_11984);
nand U13879 (N_13879,N_11142,N_11616);
nand U13880 (N_13880,N_12258,N_11070);
and U13881 (N_13881,N_10016,N_12027);
and U13882 (N_13882,N_11337,N_11745);
nor U13883 (N_13883,N_10470,N_12265);
or U13884 (N_13884,N_12278,N_10909);
nor U13885 (N_13885,N_12217,N_10607);
xor U13886 (N_13886,N_10118,N_11812);
and U13887 (N_13887,N_11228,N_11882);
nor U13888 (N_13888,N_11746,N_10759);
nand U13889 (N_13889,N_12239,N_10661);
xor U13890 (N_13890,N_10506,N_10750);
or U13891 (N_13891,N_10234,N_11071);
and U13892 (N_13892,N_12001,N_10265);
or U13893 (N_13893,N_10890,N_12254);
nand U13894 (N_13894,N_10703,N_11579);
nor U13895 (N_13895,N_11490,N_12136);
or U13896 (N_13896,N_12224,N_10159);
xor U13897 (N_13897,N_11681,N_11906);
xor U13898 (N_13898,N_11590,N_11061);
nand U13899 (N_13899,N_12190,N_10989);
nand U13900 (N_13900,N_11895,N_10876);
or U13901 (N_13901,N_10130,N_11812);
and U13902 (N_13902,N_11779,N_11214);
and U13903 (N_13903,N_10298,N_10895);
and U13904 (N_13904,N_12163,N_10311);
nor U13905 (N_13905,N_12275,N_10185);
nand U13906 (N_13906,N_11551,N_12406);
nor U13907 (N_13907,N_11776,N_12195);
and U13908 (N_13908,N_12230,N_12358);
nand U13909 (N_13909,N_11692,N_11615);
nand U13910 (N_13910,N_11884,N_12362);
and U13911 (N_13911,N_12449,N_10779);
or U13912 (N_13912,N_11841,N_10021);
nand U13913 (N_13913,N_10655,N_11053);
and U13914 (N_13914,N_12076,N_11507);
xor U13915 (N_13915,N_11360,N_10997);
xor U13916 (N_13916,N_11511,N_10161);
nor U13917 (N_13917,N_11278,N_12048);
nor U13918 (N_13918,N_10772,N_11045);
xor U13919 (N_13919,N_11990,N_12003);
xnor U13920 (N_13920,N_11278,N_12447);
xnor U13921 (N_13921,N_10169,N_11765);
nand U13922 (N_13922,N_11895,N_10873);
or U13923 (N_13923,N_11301,N_11311);
nand U13924 (N_13924,N_12469,N_11381);
and U13925 (N_13925,N_11763,N_11429);
and U13926 (N_13926,N_10652,N_12069);
and U13927 (N_13927,N_10870,N_10439);
and U13928 (N_13928,N_10446,N_10709);
nand U13929 (N_13929,N_11264,N_11651);
or U13930 (N_13930,N_11560,N_11280);
nand U13931 (N_13931,N_11269,N_12172);
or U13932 (N_13932,N_11413,N_10671);
nor U13933 (N_13933,N_11357,N_12229);
nor U13934 (N_13934,N_11898,N_12479);
or U13935 (N_13935,N_12059,N_10266);
nand U13936 (N_13936,N_11890,N_11406);
xor U13937 (N_13937,N_11706,N_10098);
or U13938 (N_13938,N_10154,N_10315);
or U13939 (N_13939,N_10729,N_11645);
nor U13940 (N_13940,N_10062,N_11832);
xnor U13941 (N_13941,N_11602,N_10709);
and U13942 (N_13942,N_10200,N_11828);
or U13943 (N_13943,N_12238,N_10283);
xnor U13944 (N_13944,N_10674,N_12039);
xnor U13945 (N_13945,N_11810,N_11012);
nand U13946 (N_13946,N_11044,N_12350);
nor U13947 (N_13947,N_10538,N_10755);
xnor U13948 (N_13948,N_11387,N_11621);
xor U13949 (N_13949,N_10954,N_10320);
nand U13950 (N_13950,N_11379,N_11505);
nor U13951 (N_13951,N_10770,N_10585);
nand U13952 (N_13952,N_10865,N_11959);
nand U13953 (N_13953,N_11094,N_10899);
nor U13954 (N_13954,N_10143,N_11749);
and U13955 (N_13955,N_11246,N_11383);
and U13956 (N_13956,N_10161,N_11879);
nor U13957 (N_13957,N_10815,N_10343);
and U13958 (N_13958,N_11752,N_10125);
nand U13959 (N_13959,N_12034,N_11023);
nor U13960 (N_13960,N_12491,N_11367);
or U13961 (N_13961,N_10788,N_11541);
or U13962 (N_13962,N_11168,N_10868);
nor U13963 (N_13963,N_11479,N_11917);
or U13964 (N_13964,N_11015,N_10811);
and U13965 (N_13965,N_11533,N_10908);
and U13966 (N_13966,N_11766,N_12391);
nor U13967 (N_13967,N_12418,N_12112);
nand U13968 (N_13968,N_11706,N_10266);
nand U13969 (N_13969,N_10807,N_11181);
or U13970 (N_13970,N_10513,N_11478);
nand U13971 (N_13971,N_10428,N_10197);
xnor U13972 (N_13972,N_11079,N_10938);
or U13973 (N_13973,N_10935,N_10283);
or U13974 (N_13974,N_12389,N_12044);
or U13975 (N_13975,N_10018,N_10232);
nor U13976 (N_13976,N_10641,N_10411);
or U13977 (N_13977,N_12458,N_10859);
nor U13978 (N_13978,N_10953,N_11995);
nor U13979 (N_13979,N_12424,N_12112);
or U13980 (N_13980,N_10623,N_10628);
nand U13981 (N_13981,N_10583,N_10766);
or U13982 (N_13982,N_11546,N_11613);
nand U13983 (N_13983,N_11376,N_10947);
or U13984 (N_13984,N_10941,N_10628);
and U13985 (N_13985,N_11289,N_10777);
nand U13986 (N_13986,N_10857,N_12002);
nor U13987 (N_13987,N_11729,N_12063);
and U13988 (N_13988,N_11450,N_11121);
nand U13989 (N_13989,N_10539,N_12347);
nand U13990 (N_13990,N_12158,N_10007);
xnor U13991 (N_13991,N_11109,N_11739);
nand U13992 (N_13992,N_11110,N_11260);
or U13993 (N_13993,N_12128,N_11886);
nor U13994 (N_13994,N_10210,N_12049);
nand U13995 (N_13995,N_10966,N_10967);
nand U13996 (N_13996,N_10924,N_11137);
nand U13997 (N_13997,N_12089,N_12294);
nor U13998 (N_13998,N_12117,N_10523);
or U13999 (N_13999,N_10278,N_10527);
nor U14000 (N_14000,N_10906,N_10728);
xor U14001 (N_14001,N_10167,N_10755);
nand U14002 (N_14002,N_10625,N_10964);
or U14003 (N_14003,N_11311,N_11676);
xor U14004 (N_14004,N_10368,N_11250);
xnor U14005 (N_14005,N_11473,N_11543);
nand U14006 (N_14006,N_11184,N_12446);
and U14007 (N_14007,N_10078,N_10234);
nor U14008 (N_14008,N_10241,N_12490);
or U14009 (N_14009,N_11508,N_11595);
xnor U14010 (N_14010,N_11614,N_10118);
and U14011 (N_14011,N_11486,N_11820);
xnor U14012 (N_14012,N_10463,N_11667);
nor U14013 (N_14013,N_11776,N_12261);
xor U14014 (N_14014,N_12484,N_10127);
or U14015 (N_14015,N_12386,N_11574);
or U14016 (N_14016,N_10014,N_11996);
nor U14017 (N_14017,N_10225,N_11216);
xor U14018 (N_14018,N_10510,N_11308);
xnor U14019 (N_14019,N_10555,N_11120);
and U14020 (N_14020,N_11467,N_11982);
and U14021 (N_14021,N_10828,N_10393);
xnor U14022 (N_14022,N_10520,N_10949);
xnor U14023 (N_14023,N_11060,N_10558);
nor U14024 (N_14024,N_10177,N_11811);
or U14025 (N_14025,N_11478,N_11780);
nor U14026 (N_14026,N_12464,N_10930);
and U14027 (N_14027,N_10807,N_10757);
or U14028 (N_14028,N_10771,N_11934);
nor U14029 (N_14029,N_10599,N_11843);
nand U14030 (N_14030,N_12106,N_10584);
or U14031 (N_14031,N_11402,N_10892);
or U14032 (N_14032,N_10990,N_11426);
and U14033 (N_14033,N_11644,N_12366);
or U14034 (N_14034,N_11307,N_11602);
nor U14035 (N_14035,N_11939,N_11378);
nand U14036 (N_14036,N_11619,N_11002);
or U14037 (N_14037,N_10391,N_12122);
nand U14038 (N_14038,N_12441,N_10871);
nor U14039 (N_14039,N_10060,N_11873);
or U14040 (N_14040,N_11171,N_11387);
and U14041 (N_14041,N_11008,N_11523);
nor U14042 (N_14042,N_12473,N_10315);
and U14043 (N_14043,N_12315,N_10525);
xor U14044 (N_14044,N_11770,N_10988);
xnor U14045 (N_14045,N_11992,N_10642);
nor U14046 (N_14046,N_10380,N_10008);
or U14047 (N_14047,N_12437,N_10921);
nand U14048 (N_14048,N_10440,N_12392);
and U14049 (N_14049,N_10161,N_12360);
and U14050 (N_14050,N_10700,N_10860);
nor U14051 (N_14051,N_11959,N_12074);
and U14052 (N_14052,N_10896,N_11591);
xor U14053 (N_14053,N_11862,N_10325);
xor U14054 (N_14054,N_11899,N_11819);
nand U14055 (N_14055,N_10819,N_11434);
nor U14056 (N_14056,N_11185,N_12142);
and U14057 (N_14057,N_10856,N_10000);
nand U14058 (N_14058,N_11323,N_12105);
and U14059 (N_14059,N_11316,N_11925);
nand U14060 (N_14060,N_12426,N_12098);
xnor U14061 (N_14061,N_12308,N_12300);
or U14062 (N_14062,N_11477,N_11227);
xnor U14063 (N_14063,N_12232,N_10940);
or U14064 (N_14064,N_10243,N_10761);
nor U14065 (N_14065,N_11481,N_11932);
nand U14066 (N_14066,N_11444,N_11653);
and U14067 (N_14067,N_10085,N_11647);
or U14068 (N_14068,N_11214,N_11116);
or U14069 (N_14069,N_10612,N_10467);
nand U14070 (N_14070,N_10581,N_11921);
nand U14071 (N_14071,N_10311,N_12419);
nor U14072 (N_14072,N_10430,N_12166);
or U14073 (N_14073,N_11483,N_11222);
and U14074 (N_14074,N_11442,N_10272);
and U14075 (N_14075,N_11182,N_10035);
and U14076 (N_14076,N_12288,N_12227);
nand U14077 (N_14077,N_10692,N_10552);
xor U14078 (N_14078,N_11179,N_11770);
nand U14079 (N_14079,N_11843,N_10289);
or U14080 (N_14080,N_12205,N_11048);
xnor U14081 (N_14081,N_12396,N_11819);
and U14082 (N_14082,N_11151,N_11444);
nor U14083 (N_14083,N_12071,N_10572);
nor U14084 (N_14084,N_12108,N_12497);
xor U14085 (N_14085,N_10702,N_10357);
or U14086 (N_14086,N_10759,N_11520);
nor U14087 (N_14087,N_12037,N_11955);
nor U14088 (N_14088,N_10796,N_11598);
nor U14089 (N_14089,N_12154,N_11210);
and U14090 (N_14090,N_10747,N_12083);
nor U14091 (N_14091,N_10104,N_10311);
xor U14092 (N_14092,N_11543,N_11479);
nor U14093 (N_14093,N_10764,N_11764);
and U14094 (N_14094,N_12061,N_11723);
nor U14095 (N_14095,N_10747,N_10544);
and U14096 (N_14096,N_12484,N_10456);
xor U14097 (N_14097,N_10670,N_10876);
nor U14098 (N_14098,N_10558,N_10776);
and U14099 (N_14099,N_11698,N_12329);
nor U14100 (N_14100,N_11800,N_11344);
or U14101 (N_14101,N_12120,N_11324);
or U14102 (N_14102,N_11444,N_12088);
or U14103 (N_14103,N_11197,N_11316);
nand U14104 (N_14104,N_12164,N_11552);
or U14105 (N_14105,N_10330,N_11499);
nor U14106 (N_14106,N_10691,N_10622);
xnor U14107 (N_14107,N_10231,N_10932);
nand U14108 (N_14108,N_10299,N_11071);
xor U14109 (N_14109,N_12053,N_11737);
nor U14110 (N_14110,N_11175,N_11542);
xnor U14111 (N_14111,N_11181,N_11163);
nand U14112 (N_14112,N_11062,N_10441);
xnor U14113 (N_14113,N_11797,N_10722);
or U14114 (N_14114,N_11222,N_12038);
nand U14115 (N_14115,N_12236,N_10687);
or U14116 (N_14116,N_11347,N_10462);
nor U14117 (N_14117,N_12424,N_12186);
nand U14118 (N_14118,N_10757,N_11705);
and U14119 (N_14119,N_10493,N_11242);
and U14120 (N_14120,N_10236,N_10914);
or U14121 (N_14121,N_12404,N_11632);
xnor U14122 (N_14122,N_11951,N_11425);
or U14123 (N_14123,N_11719,N_12012);
and U14124 (N_14124,N_11173,N_11747);
nor U14125 (N_14125,N_11967,N_11842);
nor U14126 (N_14126,N_11237,N_10590);
xor U14127 (N_14127,N_12077,N_10101);
nand U14128 (N_14128,N_11796,N_10382);
xor U14129 (N_14129,N_10782,N_10536);
xnor U14130 (N_14130,N_11209,N_11876);
nor U14131 (N_14131,N_10890,N_11815);
nor U14132 (N_14132,N_10999,N_10050);
nor U14133 (N_14133,N_12287,N_12345);
xor U14134 (N_14134,N_12490,N_10126);
and U14135 (N_14135,N_12191,N_10458);
nand U14136 (N_14136,N_10257,N_10756);
and U14137 (N_14137,N_11675,N_12183);
nand U14138 (N_14138,N_10586,N_10641);
and U14139 (N_14139,N_12358,N_10065);
or U14140 (N_14140,N_12182,N_12439);
nor U14141 (N_14141,N_10569,N_10478);
or U14142 (N_14142,N_11383,N_10262);
or U14143 (N_14143,N_10042,N_10352);
or U14144 (N_14144,N_11151,N_11636);
xor U14145 (N_14145,N_12213,N_12177);
nor U14146 (N_14146,N_11923,N_11611);
nor U14147 (N_14147,N_10394,N_12317);
xor U14148 (N_14148,N_10821,N_10035);
nand U14149 (N_14149,N_12142,N_11253);
nand U14150 (N_14150,N_11927,N_11903);
nor U14151 (N_14151,N_11976,N_10092);
or U14152 (N_14152,N_10462,N_11568);
xnor U14153 (N_14153,N_11390,N_11465);
xnor U14154 (N_14154,N_10233,N_11995);
or U14155 (N_14155,N_11055,N_12366);
xnor U14156 (N_14156,N_11182,N_11407);
nor U14157 (N_14157,N_12054,N_10924);
and U14158 (N_14158,N_10504,N_10435);
nand U14159 (N_14159,N_12414,N_12110);
xor U14160 (N_14160,N_11794,N_11991);
or U14161 (N_14161,N_11380,N_12142);
nand U14162 (N_14162,N_10100,N_10106);
xnor U14163 (N_14163,N_11591,N_12202);
or U14164 (N_14164,N_11005,N_10712);
nand U14165 (N_14165,N_11605,N_10506);
or U14166 (N_14166,N_10830,N_11792);
xnor U14167 (N_14167,N_12222,N_10548);
nand U14168 (N_14168,N_10374,N_10717);
or U14169 (N_14169,N_10953,N_11359);
or U14170 (N_14170,N_11008,N_11308);
xnor U14171 (N_14171,N_12168,N_10793);
nor U14172 (N_14172,N_11040,N_12127);
nand U14173 (N_14173,N_11545,N_12361);
and U14174 (N_14174,N_10534,N_10915);
nor U14175 (N_14175,N_12066,N_11044);
and U14176 (N_14176,N_11166,N_12158);
and U14177 (N_14177,N_11595,N_11429);
nor U14178 (N_14178,N_11905,N_11893);
nor U14179 (N_14179,N_10173,N_10763);
and U14180 (N_14180,N_11826,N_10825);
and U14181 (N_14181,N_11507,N_12492);
nor U14182 (N_14182,N_10456,N_12165);
nand U14183 (N_14183,N_12092,N_10184);
xnor U14184 (N_14184,N_11967,N_10167);
nand U14185 (N_14185,N_10814,N_10416);
and U14186 (N_14186,N_11222,N_11679);
nor U14187 (N_14187,N_11066,N_10520);
xor U14188 (N_14188,N_10339,N_11256);
nand U14189 (N_14189,N_10303,N_10774);
xnor U14190 (N_14190,N_11952,N_10923);
or U14191 (N_14191,N_10811,N_10548);
nand U14192 (N_14192,N_10338,N_10291);
xnor U14193 (N_14193,N_11425,N_11840);
nand U14194 (N_14194,N_11602,N_11055);
xor U14195 (N_14195,N_12298,N_11854);
nor U14196 (N_14196,N_11019,N_11105);
xnor U14197 (N_14197,N_10274,N_11479);
and U14198 (N_14198,N_11872,N_12033);
and U14199 (N_14199,N_12207,N_10641);
xnor U14200 (N_14200,N_10729,N_12118);
nand U14201 (N_14201,N_10116,N_12340);
nand U14202 (N_14202,N_10312,N_10160);
nand U14203 (N_14203,N_10731,N_10724);
nor U14204 (N_14204,N_10667,N_11423);
xor U14205 (N_14205,N_11361,N_11727);
xnor U14206 (N_14206,N_10660,N_12318);
nand U14207 (N_14207,N_11107,N_10612);
or U14208 (N_14208,N_11595,N_12311);
or U14209 (N_14209,N_10945,N_12491);
and U14210 (N_14210,N_11401,N_12483);
nor U14211 (N_14211,N_11549,N_11442);
nor U14212 (N_14212,N_12458,N_11318);
xnor U14213 (N_14213,N_10918,N_11064);
and U14214 (N_14214,N_11823,N_11469);
xor U14215 (N_14215,N_12365,N_10990);
nand U14216 (N_14216,N_11879,N_12107);
nor U14217 (N_14217,N_10086,N_10378);
or U14218 (N_14218,N_11138,N_10249);
nor U14219 (N_14219,N_12179,N_10377);
or U14220 (N_14220,N_10594,N_10656);
and U14221 (N_14221,N_10422,N_11177);
nand U14222 (N_14222,N_11382,N_12453);
nand U14223 (N_14223,N_11177,N_12407);
or U14224 (N_14224,N_11739,N_11639);
and U14225 (N_14225,N_10505,N_11907);
and U14226 (N_14226,N_10755,N_10444);
nand U14227 (N_14227,N_11151,N_11327);
xor U14228 (N_14228,N_11950,N_10044);
nor U14229 (N_14229,N_11137,N_11776);
nor U14230 (N_14230,N_11442,N_12272);
nor U14231 (N_14231,N_12022,N_12413);
nand U14232 (N_14232,N_10381,N_12096);
xnor U14233 (N_14233,N_12070,N_11179);
and U14234 (N_14234,N_10590,N_12292);
nand U14235 (N_14235,N_11725,N_12391);
and U14236 (N_14236,N_10428,N_11693);
nor U14237 (N_14237,N_10817,N_10026);
or U14238 (N_14238,N_10151,N_11850);
or U14239 (N_14239,N_10337,N_11065);
xnor U14240 (N_14240,N_11946,N_10398);
nand U14241 (N_14241,N_10800,N_10329);
or U14242 (N_14242,N_11468,N_10270);
and U14243 (N_14243,N_10437,N_10008);
or U14244 (N_14244,N_11174,N_10330);
and U14245 (N_14245,N_10905,N_10112);
nor U14246 (N_14246,N_12018,N_12128);
nor U14247 (N_14247,N_10457,N_12177);
nor U14248 (N_14248,N_11338,N_12173);
or U14249 (N_14249,N_12290,N_12284);
nor U14250 (N_14250,N_11471,N_10311);
or U14251 (N_14251,N_10517,N_11798);
nor U14252 (N_14252,N_12379,N_10273);
xnor U14253 (N_14253,N_10130,N_10054);
xor U14254 (N_14254,N_10404,N_10984);
nor U14255 (N_14255,N_11827,N_10236);
and U14256 (N_14256,N_11984,N_11977);
or U14257 (N_14257,N_12487,N_11866);
nand U14258 (N_14258,N_10683,N_11863);
and U14259 (N_14259,N_10945,N_10767);
and U14260 (N_14260,N_10959,N_10561);
or U14261 (N_14261,N_12418,N_12153);
nand U14262 (N_14262,N_10458,N_10981);
or U14263 (N_14263,N_10372,N_11995);
or U14264 (N_14264,N_12425,N_11015);
and U14265 (N_14265,N_10911,N_11750);
nor U14266 (N_14266,N_10934,N_11760);
nor U14267 (N_14267,N_11008,N_10569);
and U14268 (N_14268,N_12342,N_11713);
xnor U14269 (N_14269,N_11609,N_10267);
and U14270 (N_14270,N_10858,N_12092);
or U14271 (N_14271,N_11193,N_10279);
xor U14272 (N_14272,N_11482,N_10607);
and U14273 (N_14273,N_10810,N_10489);
nand U14274 (N_14274,N_12229,N_11013);
nor U14275 (N_14275,N_11609,N_10939);
xnor U14276 (N_14276,N_10353,N_11651);
or U14277 (N_14277,N_11147,N_10309);
or U14278 (N_14278,N_12335,N_12447);
nand U14279 (N_14279,N_11560,N_12030);
nand U14280 (N_14280,N_12194,N_10554);
nor U14281 (N_14281,N_10932,N_11659);
xor U14282 (N_14282,N_12123,N_11111);
xor U14283 (N_14283,N_12392,N_11803);
xor U14284 (N_14284,N_11172,N_10733);
or U14285 (N_14285,N_11203,N_12042);
nor U14286 (N_14286,N_11136,N_11405);
xnor U14287 (N_14287,N_12211,N_10123);
or U14288 (N_14288,N_11597,N_10196);
xnor U14289 (N_14289,N_10120,N_10106);
or U14290 (N_14290,N_10255,N_11308);
nor U14291 (N_14291,N_10067,N_12063);
or U14292 (N_14292,N_12199,N_11373);
nand U14293 (N_14293,N_12331,N_12484);
nor U14294 (N_14294,N_11438,N_11222);
xnor U14295 (N_14295,N_11021,N_10320);
nor U14296 (N_14296,N_11178,N_11904);
nand U14297 (N_14297,N_11795,N_11319);
nand U14298 (N_14298,N_10977,N_10228);
and U14299 (N_14299,N_10571,N_11374);
nand U14300 (N_14300,N_11636,N_11565);
and U14301 (N_14301,N_11475,N_10955);
and U14302 (N_14302,N_11171,N_12434);
and U14303 (N_14303,N_12106,N_11789);
xor U14304 (N_14304,N_12233,N_11443);
xor U14305 (N_14305,N_11681,N_10307);
and U14306 (N_14306,N_10326,N_12306);
nor U14307 (N_14307,N_11206,N_11938);
and U14308 (N_14308,N_11516,N_11787);
nor U14309 (N_14309,N_12408,N_10312);
and U14310 (N_14310,N_11094,N_11682);
nand U14311 (N_14311,N_12195,N_11684);
or U14312 (N_14312,N_11662,N_11423);
nand U14313 (N_14313,N_11802,N_11888);
nor U14314 (N_14314,N_10145,N_11245);
nor U14315 (N_14315,N_11120,N_11833);
and U14316 (N_14316,N_10140,N_11627);
nand U14317 (N_14317,N_10831,N_10900);
or U14318 (N_14318,N_10050,N_11146);
xnor U14319 (N_14319,N_12049,N_11654);
xnor U14320 (N_14320,N_10486,N_11587);
xnor U14321 (N_14321,N_10939,N_12248);
and U14322 (N_14322,N_10877,N_11429);
and U14323 (N_14323,N_10669,N_11532);
nand U14324 (N_14324,N_10081,N_10636);
nor U14325 (N_14325,N_10256,N_10965);
and U14326 (N_14326,N_12232,N_10912);
or U14327 (N_14327,N_10694,N_11825);
xor U14328 (N_14328,N_10088,N_12219);
xnor U14329 (N_14329,N_12339,N_11257);
xor U14330 (N_14330,N_11022,N_10010);
or U14331 (N_14331,N_12052,N_10420);
or U14332 (N_14332,N_10917,N_10447);
or U14333 (N_14333,N_10569,N_11231);
nor U14334 (N_14334,N_11641,N_11819);
nand U14335 (N_14335,N_12052,N_10274);
and U14336 (N_14336,N_12109,N_10051);
xor U14337 (N_14337,N_10375,N_12130);
and U14338 (N_14338,N_12364,N_11483);
nor U14339 (N_14339,N_11446,N_10956);
nor U14340 (N_14340,N_12233,N_10828);
and U14341 (N_14341,N_10339,N_11201);
and U14342 (N_14342,N_12272,N_11144);
and U14343 (N_14343,N_10390,N_12309);
and U14344 (N_14344,N_11370,N_10447);
xor U14345 (N_14345,N_12280,N_11813);
and U14346 (N_14346,N_11843,N_12215);
and U14347 (N_14347,N_12192,N_11300);
and U14348 (N_14348,N_10274,N_11911);
xnor U14349 (N_14349,N_11897,N_12456);
nor U14350 (N_14350,N_10822,N_10343);
or U14351 (N_14351,N_11829,N_11978);
and U14352 (N_14352,N_10715,N_11092);
and U14353 (N_14353,N_11381,N_11735);
or U14354 (N_14354,N_12257,N_10010);
xnor U14355 (N_14355,N_11989,N_11480);
and U14356 (N_14356,N_12179,N_10956);
nand U14357 (N_14357,N_10790,N_12319);
or U14358 (N_14358,N_12400,N_11770);
or U14359 (N_14359,N_10186,N_11346);
nor U14360 (N_14360,N_11255,N_10063);
xnor U14361 (N_14361,N_10127,N_12046);
or U14362 (N_14362,N_11058,N_11763);
or U14363 (N_14363,N_12058,N_11740);
or U14364 (N_14364,N_11370,N_10535);
or U14365 (N_14365,N_12132,N_10537);
xnor U14366 (N_14366,N_10657,N_11101);
nand U14367 (N_14367,N_10949,N_12288);
or U14368 (N_14368,N_10253,N_12344);
nor U14369 (N_14369,N_11401,N_10422);
or U14370 (N_14370,N_12272,N_10506);
or U14371 (N_14371,N_12063,N_10357);
and U14372 (N_14372,N_10615,N_10919);
xor U14373 (N_14373,N_10072,N_12281);
or U14374 (N_14374,N_10843,N_10184);
or U14375 (N_14375,N_11212,N_11163);
or U14376 (N_14376,N_11952,N_11129);
nand U14377 (N_14377,N_10495,N_10492);
nor U14378 (N_14378,N_11236,N_11803);
nand U14379 (N_14379,N_12131,N_11371);
and U14380 (N_14380,N_10116,N_10866);
nor U14381 (N_14381,N_10353,N_11159);
nand U14382 (N_14382,N_10861,N_11938);
and U14383 (N_14383,N_10808,N_10385);
and U14384 (N_14384,N_12061,N_12060);
and U14385 (N_14385,N_10434,N_12489);
or U14386 (N_14386,N_10215,N_12248);
xor U14387 (N_14387,N_11100,N_10926);
nand U14388 (N_14388,N_10081,N_11082);
or U14389 (N_14389,N_12286,N_10840);
xor U14390 (N_14390,N_11655,N_12126);
nand U14391 (N_14391,N_11955,N_10160);
nor U14392 (N_14392,N_12093,N_10094);
and U14393 (N_14393,N_12155,N_12016);
or U14394 (N_14394,N_10230,N_11215);
or U14395 (N_14395,N_10400,N_12330);
or U14396 (N_14396,N_12136,N_10110);
and U14397 (N_14397,N_11391,N_11344);
or U14398 (N_14398,N_11161,N_11750);
nand U14399 (N_14399,N_12361,N_10161);
nor U14400 (N_14400,N_10691,N_11971);
nor U14401 (N_14401,N_11684,N_12309);
or U14402 (N_14402,N_11544,N_10757);
or U14403 (N_14403,N_11270,N_11843);
and U14404 (N_14404,N_12319,N_10886);
and U14405 (N_14405,N_10267,N_11300);
or U14406 (N_14406,N_10956,N_10738);
or U14407 (N_14407,N_11679,N_10607);
or U14408 (N_14408,N_10280,N_11576);
nand U14409 (N_14409,N_11226,N_12477);
nor U14410 (N_14410,N_11881,N_12081);
xnor U14411 (N_14411,N_11762,N_11924);
nor U14412 (N_14412,N_10606,N_12362);
or U14413 (N_14413,N_11274,N_10385);
and U14414 (N_14414,N_10025,N_10531);
xor U14415 (N_14415,N_11276,N_12381);
nor U14416 (N_14416,N_12398,N_11142);
or U14417 (N_14417,N_11581,N_10066);
nor U14418 (N_14418,N_11728,N_10515);
or U14419 (N_14419,N_11764,N_12406);
nor U14420 (N_14420,N_11228,N_12355);
xnor U14421 (N_14421,N_10575,N_10921);
nand U14422 (N_14422,N_10979,N_10642);
nand U14423 (N_14423,N_12252,N_10321);
nand U14424 (N_14424,N_10055,N_11779);
nand U14425 (N_14425,N_10487,N_10467);
nand U14426 (N_14426,N_10355,N_10461);
and U14427 (N_14427,N_10943,N_11361);
xnor U14428 (N_14428,N_10229,N_11606);
xnor U14429 (N_14429,N_11974,N_10367);
xnor U14430 (N_14430,N_11224,N_10316);
and U14431 (N_14431,N_11599,N_12270);
nand U14432 (N_14432,N_11677,N_11553);
and U14433 (N_14433,N_10414,N_10768);
nor U14434 (N_14434,N_11759,N_10989);
nand U14435 (N_14435,N_10950,N_12172);
nor U14436 (N_14436,N_11390,N_11328);
nor U14437 (N_14437,N_10540,N_10811);
and U14438 (N_14438,N_11431,N_10352);
nand U14439 (N_14439,N_10362,N_11690);
nand U14440 (N_14440,N_12146,N_11722);
nor U14441 (N_14441,N_10040,N_10966);
and U14442 (N_14442,N_11433,N_11223);
and U14443 (N_14443,N_11997,N_10888);
xor U14444 (N_14444,N_12022,N_12248);
and U14445 (N_14445,N_11744,N_12032);
xnor U14446 (N_14446,N_11634,N_12395);
and U14447 (N_14447,N_10592,N_10723);
or U14448 (N_14448,N_10051,N_12323);
xor U14449 (N_14449,N_11532,N_11341);
or U14450 (N_14450,N_11745,N_10531);
and U14451 (N_14451,N_10020,N_12245);
or U14452 (N_14452,N_11392,N_10506);
nand U14453 (N_14453,N_10341,N_10967);
nand U14454 (N_14454,N_12058,N_10348);
xnor U14455 (N_14455,N_12371,N_10528);
and U14456 (N_14456,N_11651,N_10587);
nor U14457 (N_14457,N_10766,N_11265);
and U14458 (N_14458,N_11048,N_11167);
and U14459 (N_14459,N_11517,N_11729);
or U14460 (N_14460,N_10173,N_11709);
or U14461 (N_14461,N_12322,N_10211);
nor U14462 (N_14462,N_12476,N_10631);
nand U14463 (N_14463,N_10927,N_10965);
xnor U14464 (N_14464,N_12080,N_10844);
or U14465 (N_14465,N_11803,N_11624);
nand U14466 (N_14466,N_11141,N_11024);
or U14467 (N_14467,N_12239,N_10304);
nor U14468 (N_14468,N_12427,N_11261);
xor U14469 (N_14469,N_10133,N_11432);
or U14470 (N_14470,N_12091,N_10592);
and U14471 (N_14471,N_10988,N_11169);
and U14472 (N_14472,N_11177,N_11395);
and U14473 (N_14473,N_10651,N_10575);
or U14474 (N_14474,N_12050,N_12332);
nand U14475 (N_14475,N_11570,N_10899);
or U14476 (N_14476,N_11349,N_10001);
xnor U14477 (N_14477,N_11060,N_11615);
or U14478 (N_14478,N_10966,N_11748);
nor U14479 (N_14479,N_10550,N_11668);
and U14480 (N_14480,N_10933,N_11662);
or U14481 (N_14481,N_11226,N_10587);
and U14482 (N_14482,N_10390,N_10129);
or U14483 (N_14483,N_10664,N_12419);
and U14484 (N_14484,N_10677,N_10483);
or U14485 (N_14485,N_12348,N_11956);
xor U14486 (N_14486,N_11635,N_11790);
or U14487 (N_14487,N_11095,N_11745);
and U14488 (N_14488,N_11622,N_10751);
xor U14489 (N_14489,N_11851,N_11681);
or U14490 (N_14490,N_12155,N_10124);
xnor U14491 (N_14491,N_10736,N_12472);
and U14492 (N_14492,N_10990,N_12161);
nor U14493 (N_14493,N_11996,N_10152);
or U14494 (N_14494,N_11216,N_10653);
nand U14495 (N_14495,N_11828,N_11361);
xnor U14496 (N_14496,N_11246,N_11855);
or U14497 (N_14497,N_12044,N_10743);
or U14498 (N_14498,N_11009,N_11478);
nor U14499 (N_14499,N_10850,N_12306);
xor U14500 (N_14500,N_11209,N_11249);
or U14501 (N_14501,N_12172,N_10348);
nor U14502 (N_14502,N_10729,N_12332);
xor U14503 (N_14503,N_11016,N_12330);
nand U14504 (N_14504,N_10109,N_12136);
and U14505 (N_14505,N_12003,N_10184);
or U14506 (N_14506,N_11656,N_10669);
nor U14507 (N_14507,N_10188,N_11124);
nor U14508 (N_14508,N_11030,N_11431);
xnor U14509 (N_14509,N_11738,N_10976);
and U14510 (N_14510,N_10594,N_10190);
or U14511 (N_14511,N_12158,N_10731);
xor U14512 (N_14512,N_10293,N_11106);
or U14513 (N_14513,N_11011,N_10693);
and U14514 (N_14514,N_10868,N_12374);
nand U14515 (N_14515,N_11065,N_11776);
xnor U14516 (N_14516,N_12396,N_10090);
or U14517 (N_14517,N_11040,N_11987);
nor U14518 (N_14518,N_10412,N_10878);
or U14519 (N_14519,N_10310,N_11815);
xor U14520 (N_14520,N_10848,N_10129);
and U14521 (N_14521,N_10263,N_11732);
and U14522 (N_14522,N_10576,N_10772);
nor U14523 (N_14523,N_12480,N_10509);
nor U14524 (N_14524,N_12460,N_10397);
nand U14525 (N_14525,N_10482,N_12377);
or U14526 (N_14526,N_11171,N_11834);
and U14527 (N_14527,N_10372,N_10260);
or U14528 (N_14528,N_11990,N_10345);
and U14529 (N_14529,N_10077,N_12147);
or U14530 (N_14530,N_10216,N_11653);
xnor U14531 (N_14531,N_11048,N_11494);
nand U14532 (N_14532,N_11346,N_12412);
xnor U14533 (N_14533,N_11805,N_11940);
or U14534 (N_14534,N_10822,N_12025);
or U14535 (N_14535,N_10632,N_11793);
nor U14536 (N_14536,N_11729,N_11286);
nand U14537 (N_14537,N_11755,N_11695);
xor U14538 (N_14538,N_10702,N_10945);
or U14539 (N_14539,N_11752,N_10003);
and U14540 (N_14540,N_12371,N_11309);
or U14541 (N_14541,N_12382,N_12358);
nor U14542 (N_14542,N_10715,N_12079);
xor U14543 (N_14543,N_10628,N_10540);
nand U14544 (N_14544,N_11343,N_11256);
and U14545 (N_14545,N_11354,N_10063);
or U14546 (N_14546,N_11506,N_12401);
nand U14547 (N_14547,N_10933,N_11489);
nand U14548 (N_14548,N_11596,N_10256);
or U14549 (N_14549,N_11034,N_10803);
nand U14550 (N_14550,N_11849,N_10769);
or U14551 (N_14551,N_11465,N_12405);
nor U14552 (N_14552,N_10151,N_11384);
or U14553 (N_14553,N_11799,N_10278);
nand U14554 (N_14554,N_12329,N_10126);
or U14555 (N_14555,N_10358,N_10965);
xnor U14556 (N_14556,N_11447,N_12003);
and U14557 (N_14557,N_10599,N_12081);
and U14558 (N_14558,N_10248,N_12341);
xor U14559 (N_14559,N_11047,N_11733);
nand U14560 (N_14560,N_11423,N_10566);
nor U14561 (N_14561,N_12277,N_12139);
nor U14562 (N_14562,N_10010,N_10497);
and U14563 (N_14563,N_10363,N_10755);
and U14564 (N_14564,N_11799,N_10452);
nor U14565 (N_14565,N_10369,N_11472);
nor U14566 (N_14566,N_11488,N_12285);
nand U14567 (N_14567,N_10419,N_10891);
or U14568 (N_14568,N_10344,N_12409);
nor U14569 (N_14569,N_11097,N_10792);
and U14570 (N_14570,N_10720,N_10661);
nand U14571 (N_14571,N_11826,N_11056);
or U14572 (N_14572,N_10359,N_11444);
nand U14573 (N_14573,N_10618,N_11102);
nand U14574 (N_14574,N_10592,N_11485);
nand U14575 (N_14575,N_12407,N_12456);
and U14576 (N_14576,N_11247,N_11180);
nor U14577 (N_14577,N_11443,N_12338);
nand U14578 (N_14578,N_10207,N_11983);
and U14579 (N_14579,N_11017,N_11634);
and U14580 (N_14580,N_10353,N_12100);
and U14581 (N_14581,N_10127,N_12395);
nand U14582 (N_14582,N_11079,N_11429);
xor U14583 (N_14583,N_12057,N_12370);
nand U14584 (N_14584,N_11094,N_11727);
nor U14585 (N_14585,N_10741,N_12348);
xor U14586 (N_14586,N_10745,N_10329);
xor U14587 (N_14587,N_11288,N_11265);
nor U14588 (N_14588,N_11654,N_12092);
or U14589 (N_14589,N_12221,N_11583);
and U14590 (N_14590,N_11653,N_10028);
and U14591 (N_14591,N_10005,N_12368);
and U14592 (N_14592,N_10808,N_11266);
and U14593 (N_14593,N_11170,N_11406);
nand U14594 (N_14594,N_10899,N_11425);
and U14595 (N_14595,N_11712,N_10447);
or U14596 (N_14596,N_11816,N_11702);
xor U14597 (N_14597,N_11079,N_11936);
nand U14598 (N_14598,N_10424,N_12092);
xnor U14599 (N_14599,N_10154,N_10598);
or U14600 (N_14600,N_10314,N_12065);
nand U14601 (N_14601,N_10679,N_10369);
xor U14602 (N_14602,N_12496,N_10394);
nor U14603 (N_14603,N_10358,N_11802);
or U14604 (N_14604,N_10196,N_11728);
nor U14605 (N_14605,N_11357,N_10209);
or U14606 (N_14606,N_11663,N_11930);
nor U14607 (N_14607,N_12365,N_10285);
nand U14608 (N_14608,N_10576,N_12404);
nand U14609 (N_14609,N_10440,N_11379);
xor U14610 (N_14610,N_11375,N_12489);
or U14611 (N_14611,N_12283,N_11494);
or U14612 (N_14612,N_11177,N_11202);
or U14613 (N_14613,N_11409,N_12463);
xnor U14614 (N_14614,N_10313,N_10673);
nor U14615 (N_14615,N_10285,N_11627);
and U14616 (N_14616,N_12457,N_10292);
nor U14617 (N_14617,N_11573,N_11589);
or U14618 (N_14618,N_11123,N_10762);
nor U14619 (N_14619,N_11101,N_12209);
xor U14620 (N_14620,N_11999,N_12296);
nand U14621 (N_14621,N_10691,N_12081);
nor U14622 (N_14622,N_12059,N_11944);
nand U14623 (N_14623,N_12268,N_10633);
xnor U14624 (N_14624,N_11705,N_11019);
nand U14625 (N_14625,N_10919,N_12498);
nor U14626 (N_14626,N_11354,N_10948);
xor U14627 (N_14627,N_10268,N_11852);
and U14628 (N_14628,N_11848,N_10026);
or U14629 (N_14629,N_11973,N_12066);
or U14630 (N_14630,N_10678,N_12496);
nor U14631 (N_14631,N_10077,N_12031);
xor U14632 (N_14632,N_10161,N_10527);
nor U14633 (N_14633,N_10341,N_12087);
nand U14634 (N_14634,N_10814,N_11733);
nor U14635 (N_14635,N_11049,N_11564);
or U14636 (N_14636,N_10230,N_12064);
xor U14637 (N_14637,N_12112,N_10132);
nand U14638 (N_14638,N_11899,N_10624);
nor U14639 (N_14639,N_10372,N_10093);
nor U14640 (N_14640,N_11233,N_11580);
nand U14641 (N_14641,N_10329,N_12455);
xor U14642 (N_14642,N_11681,N_12220);
xnor U14643 (N_14643,N_11084,N_10079);
or U14644 (N_14644,N_11486,N_10437);
and U14645 (N_14645,N_10781,N_10954);
xor U14646 (N_14646,N_11448,N_10656);
and U14647 (N_14647,N_10015,N_11081);
or U14648 (N_14648,N_11260,N_11122);
and U14649 (N_14649,N_12086,N_11273);
and U14650 (N_14650,N_10407,N_11183);
or U14651 (N_14651,N_11364,N_11104);
or U14652 (N_14652,N_12432,N_10242);
nand U14653 (N_14653,N_11785,N_10657);
nor U14654 (N_14654,N_11347,N_11073);
or U14655 (N_14655,N_11516,N_12061);
xnor U14656 (N_14656,N_10765,N_11075);
nand U14657 (N_14657,N_12232,N_12416);
and U14658 (N_14658,N_11704,N_10845);
and U14659 (N_14659,N_11221,N_10800);
or U14660 (N_14660,N_11440,N_10871);
nor U14661 (N_14661,N_12460,N_12473);
and U14662 (N_14662,N_10201,N_10835);
or U14663 (N_14663,N_11595,N_10525);
nor U14664 (N_14664,N_12165,N_12447);
nor U14665 (N_14665,N_11948,N_12431);
and U14666 (N_14666,N_12195,N_11380);
nor U14667 (N_14667,N_11075,N_12013);
nor U14668 (N_14668,N_11060,N_10299);
nor U14669 (N_14669,N_11121,N_11898);
nand U14670 (N_14670,N_11343,N_11651);
and U14671 (N_14671,N_12499,N_10070);
xnor U14672 (N_14672,N_12078,N_11693);
and U14673 (N_14673,N_11953,N_10982);
nand U14674 (N_14674,N_10558,N_12078);
xnor U14675 (N_14675,N_11001,N_10265);
nor U14676 (N_14676,N_10574,N_11187);
and U14677 (N_14677,N_11633,N_10634);
nand U14678 (N_14678,N_11411,N_10690);
and U14679 (N_14679,N_11640,N_11969);
and U14680 (N_14680,N_12413,N_10517);
xnor U14681 (N_14681,N_12037,N_12345);
xnor U14682 (N_14682,N_10165,N_11953);
nor U14683 (N_14683,N_10107,N_12241);
nor U14684 (N_14684,N_11464,N_10248);
nor U14685 (N_14685,N_10984,N_12424);
xor U14686 (N_14686,N_12148,N_11511);
or U14687 (N_14687,N_11096,N_11869);
or U14688 (N_14688,N_12022,N_12416);
nor U14689 (N_14689,N_10296,N_10349);
nand U14690 (N_14690,N_12458,N_10628);
and U14691 (N_14691,N_11051,N_10362);
or U14692 (N_14692,N_10857,N_11640);
nand U14693 (N_14693,N_11173,N_11861);
and U14694 (N_14694,N_12025,N_10043);
xor U14695 (N_14695,N_12056,N_11160);
nand U14696 (N_14696,N_10765,N_12300);
nand U14697 (N_14697,N_11380,N_11279);
nand U14698 (N_14698,N_11931,N_10977);
nor U14699 (N_14699,N_11951,N_11385);
nor U14700 (N_14700,N_10269,N_11768);
or U14701 (N_14701,N_11938,N_10468);
nor U14702 (N_14702,N_12023,N_11047);
nand U14703 (N_14703,N_10962,N_12326);
and U14704 (N_14704,N_12419,N_11217);
nor U14705 (N_14705,N_11042,N_12424);
nand U14706 (N_14706,N_11407,N_12206);
xnor U14707 (N_14707,N_12024,N_10805);
and U14708 (N_14708,N_10230,N_12391);
nand U14709 (N_14709,N_12337,N_10714);
and U14710 (N_14710,N_12009,N_11706);
xnor U14711 (N_14711,N_10942,N_11803);
nand U14712 (N_14712,N_12298,N_12491);
nor U14713 (N_14713,N_11125,N_11012);
nor U14714 (N_14714,N_11307,N_11560);
xor U14715 (N_14715,N_12199,N_10518);
and U14716 (N_14716,N_10365,N_10695);
and U14717 (N_14717,N_10523,N_10052);
and U14718 (N_14718,N_11535,N_11646);
nor U14719 (N_14719,N_10107,N_12398);
xnor U14720 (N_14720,N_12026,N_10654);
or U14721 (N_14721,N_12402,N_11812);
xnor U14722 (N_14722,N_11484,N_12222);
or U14723 (N_14723,N_11957,N_10469);
or U14724 (N_14724,N_10815,N_10738);
or U14725 (N_14725,N_11970,N_10581);
nand U14726 (N_14726,N_10881,N_11107);
nand U14727 (N_14727,N_10202,N_12429);
nand U14728 (N_14728,N_11847,N_12165);
nor U14729 (N_14729,N_10163,N_11322);
and U14730 (N_14730,N_12169,N_12407);
nand U14731 (N_14731,N_12069,N_10955);
xor U14732 (N_14732,N_10332,N_10833);
nand U14733 (N_14733,N_12053,N_10822);
and U14734 (N_14734,N_11519,N_11538);
or U14735 (N_14735,N_11998,N_11609);
or U14736 (N_14736,N_11965,N_12418);
nor U14737 (N_14737,N_12299,N_11219);
xor U14738 (N_14738,N_10034,N_12174);
or U14739 (N_14739,N_10239,N_10520);
or U14740 (N_14740,N_12458,N_11906);
and U14741 (N_14741,N_11622,N_11789);
or U14742 (N_14742,N_10486,N_11180);
nor U14743 (N_14743,N_11846,N_10062);
xnor U14744 (N_14744,N_12276,N_12112);
nand U14745 (N_14745,N_11203,N_12460);
or U14746 (N_14746,N_11631,N_11156);
or U14747 (N_14747,N_10613,N_11931);
nand U14748 (N_14748,N_12270,N_12122);
nor U14749 (N_14749,N_12258,N_10093);
and U14750 (N_14750,N_11919,N_11669);
and U14751 (N_14751,N_11469,N_12138);
or U14752 (N_14752,N_10117,N_11332);
nand U14753 (N_14753,N_10055,N_10592);
and U14754 (N_14754,N_10088,N_11969);
nor U14755 (N_14755,N_11110,N_12011);
xor U14756 (N_14756,N_11445,N_10909);
and U14757 (N_14757,N_12425,N_11157);
nor U14758 (N_14758,N_10468,N_10919);
or U14759 (N_14759,N_12198,N_11121);
xnor U14760 (N_14760,N_11796,N_10777);
nor U14761 (N_14761,N_11034,N_10995);
or U14762 (N_14762,N_12441,N_10451);
and U14763 (N_14763,N_12181,N_11972);
and U14764 (N_14764,N_12112,N_11289);
and U14765 (N_14765,N_11331,N_10329);
and U14766 (N_14766,N_11164,N_11504);
or U14767 (N_14767,N_12484,N_11547);
or U14768 (N_14768,N_10170,N_11678);
xnor U14769 (N_14769,N_11302,N_11910);
nand U14770 (N_14770,N_10929,N_12198);
or U14771 (N_14771,N_10464,N_11306);
nor U14772 (N_14772,N_10440,N_12376);
nor U14773 (N_14773,N_10245,N_10699);
and U14774 (N_14774,N_10183,N_10237);
nand U14775 (N_14775,N_12184,N_11037);
xor U14776 (N_14776,N_11631,N_12459);
or U14777 (N_14777,N_10099,N_10455);
and U14778 (N_14778,N_11129,N_11205);
or U14779 (N_14779,N_10043,N_11298);
xor U14780 (N_14780,N_11905,N_12383);
nor U14781 (N_14781,N_11241,N_11078);
or U14782 (N_14782,N_11038,N_11635);
nor U14783 (N_14783,N_10778,N_10759);
nand U14784 (N_14784,N_11200,N_11564);
and U14785 (N_14785,N_11883,N_11202);
nand U14786 (N_14786,N_12484,N_11573);
and U14787 (N_14787,N_12215,N_12197);
or U14788 (N_14788,N_11236,N_10775);
nand U14789 (N_14789,N_10192,N_11933);
nor U14790 (N_14790,N_10061,N_11440);
or U14791 (N_14791,N_10561,N_11761);
nor U14792 (N_14792,N_12430,N_10295);
or U14793 (N_14793,N_10063,N_11028);
xnor U14794 (N_14794,N_12402,N_10738);
nand U14795 (N_14795,N_11991,N_11129);
or U14796 (N_14796,N_11392,N_10940);
or U14797 (N_14797,N_11658,N_10046);
nor U14798 (N_14798,N_12182,N_11673);
or U14799 (N_14799,N_12075,N_11023);
or U14800 (N_14800,N_11618,N_10471);
nand U14801 (N_14801,N_12253,N_11366);
nor U14802 (N_14802,N_10682,N_12261);
xor U14803 (N_14803,N_10654,N_10448);
nor U14804 (N_14804,N_12028,N_10869);
nand U14805 (N_14805,N_11214,N_11243);
nand U14806 (N_14806,N_10416,N_10165);
xnor U14807 (N_14807,N_10283,N_11097);
nor U14808 (N_14808,N_10842,N_12407);
or U14809 (N_14809,N_11348,N_10926);
nand U14810 (N_14810,N_11831,N_11603);
nor U14811 (N_14811,N_11463,N_11065);
xnor U14812 (N_14812,N_10642,N_10375);
and U14813 (N_14813,N_11868,N_11977);
nand U14814 (N_14814,N_11275,N_11231);
or U14815 (N_14815,N_12079,N_10998);
xnor U14816 (N_14816,N_11269,N_10569);
nor U14817 (N_14817,N_12348,N_11630);
and U14818 (N_14818,N_11896,N_10166);
xnor U14819 (N_14819,N_12488,N_11657);
or U14820 (N_14820,N_11515,N_12426);
nand U14821 (N_14821,N_10710,N_10885);
nand U14822 (N_14822,N_11331,N_11480);
nand U14823 (N_14823,N_10584,N_11259);
or U14824 (N_14824,N_10209,N_10653);
nor U14825 (N_14825,N_12081,N_12174);
and U14826 (N_14826,N_12455,N_10459);
nor U14827 (N_14827,N_11536,N_11734);
or U14828 (N_14828,N_11410,N_12496);
nor U14829 (N_14829,N_12015,N_12476);
nand U14830 (N_14830,N_10256,N_11760);
or U14831 (N_14831,N_10769,N_11771);
or U14832 (N_14832,N_12270,N_10432);
or U14833 (N_14833,N_11491,N_12119);
nor U14834 (N_14834,N_12134,N_11553);
nor U14835 (N_14835,N_11594,N_10045);
or U14836 (N_14836,N_11654,N_12205);
xnor U14837 (N_14837,N_11033,N_10319);
xor U14838 (N_14838,N_10905,N_11198);
nor U14839 (N_14839,N_11198,N_10347);
or U14840 (N_14840,N_11896,N_11793);
or U14841 (N_14841,N_12357,N_12172);
xor U14842 (N_14842,N_10210,N_11998);
or U14843 (N_14843,N_11511,N_12445);
nand U14844 (N_14844,N_10271,N_10656);
nor U14845 (N_14845,N_11971,N_12421);
nor U14846 (N_14846,N_11784,N_11579);
or U14847 (N_14847,N_10108,N_10315);
xnor U14848 (N_14848,N_10808,N_10766);
and U14849 (N_14849,N_11405,N_12492);
nand U14850 (N_14850,N_12314,N_11019);
nor U14851 (N_14851,N_10258,N_10798);
xor U14852 (N_14852,N_10963,N_10168);
or U14853 (N_14853,N_12290,N_11312);
nor U14854 (N_14854,N_11392,N_11724);
nor U14855 (N_14855,N_11762,N_10795);
and U14856 (N_14856,N_11007,N_10036);
or U14857 (N_14857,N_10228,N_10971);
xnor U14858 (N_14858,N_12287,N_12410);
and U14859 (N_14859,N_10853,N_12398);
or U14860 (N_14860,N_10056,N_11853);
nand U14861 (N_14861,N_12133,N_11998);
nor U14862 (N_14862,N_10518,N_11951);
or U14863 (N_14863,N_10788,N_11204);
or U14864 (N_14864,N_11470,N_11618);
nor U14865 (N_14865,N_10663,N_11295);
and U14866 (N_14866,N_10405,N_11370);
nor U14867 (N_14867,N_10254,N_10929);
nand U14868 (N_14868,N_10866,N_11116);
xor U14869 (N_14869,N_10288,N_10169);
nor U14870 (N_14870,N_10000,N_11594);
nor U14871 (N_14871,N_11034,N_10012);
nand U14872 (N_14872,N_10055,N_11378);
nor U14873 (N_14873,N_11936,N_11397);
xnor U14874 (N_14874,N_10195,N_10541);
nor U14875 (N_14875,N_11984,N_10958);
nand U14876 (N_14876,N_10638,N_10106);
and U14877 (N_14877,N_11604,N_11017);
xor U14878 (N_14878,N_11009,N_10074);
nand U14879 (N_14879,N_11796,N_12042);
nor U14880 (N_14880,N_11694,N_12187);
xnor U14881 (N_14881,N_10520,N_10607);
or U14882 (N_14882,N_10301,N_12334);
or U14883 (N_14883,N_11562,N_12312);
xor U14884 (N_14884,N_11650,N_10768);
or U14885 (N_14885,N_10949,N_10604);
and U14886 (N_14886,N_11259,N_12040);
nand U14887 (N_14887,N_11744,N_12211);
or U14888 (N_14888,N_11742,N_12195);
or U14889 (N_14889,N_10626,N_12477);
xor U14890 (N_14890,N_11639,N_10222);
nand U14891 (N_14891,N_12341,N_10394);
nand U14892 (N_14892,N_10288,N_12013);
or U14893 (N_14893,N_10104,N_12112);
or U14894 (N_14894,N_10044,N_12392);
nor U14895 (N_14895,N_10796,N_12193);
nor U14896 (N_14896,N_10974,N_10038);
xnor U14897 (N_14897,N_10892,N_10555);
or U14898 (N_14898,N_12086,N_11837);
xor U14899 (N_14899,N_11531,N_11462);
nand U14900 (N_14900,N_10616,N_11544);
nand U14901 (N_14901,N_10050,N_10523);
or U14902 (N_14902,N_12125,N_11334);
nor U14903 (N_14903,N_11027,N_11643);
nor U14904 (N_14904,N_11021,N_10134);
nor U14905 (N_14905,N_11996,N_10111);
and U14906 (N_14906,N_10331,N_12146);
xnor U14907 (N_14907,N_10666,N_10178);
or U14908 (N_14908,N_11226,N_11477);
and U14909 (N_14909,N_10001,N_11974);
xnor U14910 (N_14910,N_11610,N_10825);
nand U14911 (N_14911,N_11732,N_10166);
and U14912 (N_14912,N_11164,N_10165);
xor U14913 (N_14913,N_12387,N_11190);
nand U14914 (N_14914,N_10543,N_11239);
or U14915 (N_14915,N_10158,N_11156);
or U14916 (N_14916,N_10329,N_11492);
xor U14917 (N_14917,N_12056,N_10363);
or U14918 (N_14918,N_11023,N_12024);
nor U14919 (N_14919,N_11353,N_11649);
xnor U14920 (N_14920,N_12149,N_11951);
nand U14921 (N_14921,N_10298,N_10440);
nand U14922 (N_14922,N_11906,N_10874);
nand U14923 (N_14923,N_10659,N_11830);
nor U14924 (N_14924,N_11739,N_10058);
nor U14925 (N_14925,N_11729,N_10487);
and U14926 (N_14926,N_12480,N_11379);
and U14927 (N_14927,N_11816,N_12459);
or U14928 (N_14928,N_10868,N_10840);
nand U14929 (N_14929,N_10918,N_11166);
xnor U14930 (N_14930,N_10761,N_11878);
nor U14931 (N_14931,N_11863,N_10306);
nor U14932 (N_14932,N_11357,N_11244);
or U14933 (N_14933,N_10134,N_10692);
xnor U14934 (N_14934,N_11941,N_11272);
and U14935 (N_14935,N_11217,N_11415);
and U14936 (N_14936,N_11282,N_12104);
xnor U14937 (N_14937,N_10241,N_12438);
nand U14938 (N_14938,N_12068,N_12174);
and U14939 (N_14939,N_10929,N_11910);
xor U14940 (N_14940,N_10288,N_11589);
nand U14941 (N_14941,N_10009,N_11761);
or U14942 (N_14942,N_12210,N_10102);
and U14943 (N_14943,N_11297,N_12024);
nor U14944 (N_14944,N_10123,N_12006);
and U14945 (N_14945,N_11550,N_12141);
xnor U14946 (N_14946,N_11131,N_11063);
xor U14947 (N_14947,N_10933,N_11570);
xnor U14948 (N_14948,N_10828,N_12421);
or U14949 (N_14949,N_11186,N_12180);
nor U14950 (N_14950,N_10796,N_10909);
or U14951 (N_14951,N_11257,N_11614);
and U14952 (N_14952,N_12157,N_11685);
xnor U14953 (N_14953,N_11801,N_10397);
nor U14954 (N_14954,N_11905,N_12377);
or U14955 (N_14955,N_12107,N_10918);
xnor U14956 (N_14956,N_11998,N_10608);
nor U14957 (N_14957,N_10583,N_11768);
nand U14958 (N_14958,N_11112,N_10969);
nor U14959 (N_14959,N_10391,N_10863);
and U14960 (N_14960,N_10426,N_10777);
xnor U14961 (N_14961,N_11093,N_11818);
and U14962 (N_14962,N_11000,N_12393);
nor U14963 (N_14963,N_12176,N_10478);
nor U14964 (N_14964,N_12453,N_10606);
xnor U14965 (N_14965,N_10097,N_10713);
or U14966 (N_14966,N_12319,N_11999);
or U14967 (N_14967,N_11687,N_11849);
nand U14968 (N_14968,N_11177,N_10057);
xnor U14969 (N_14969,N_11267,N_12390);
or U14970 (N_14970,N_11699,N_10973);
nor U14971 (N_14971,N_11998,N_11249);
nand U14972 (N_14972,N_12215,N_11384);
nand U14973 (N_14973,N_12117,N_11314);
nor U14974 (N_14974,N_11889,N_12256);
and U14975 (N_14975,N_10709,N_11250);
nor U14976 (N_14976,N_10910,N_11708);
nand U14977 (N_14977,N_10265,N_11683);
and U14978 (N_14978,N_12413,N_12142);
or U14979 (N_14979,N_10497,N_10766);
nand U14980 (N_14980,N_10688,N_10484);
and U14981 (N_14981,N_12343,N_11969);
nand U14982 (N_14982,N_11309,N_11895);
nand U14983 (N_14983,N_11294,N_11735);
nand U14984 (N_14984,N_12170,N_11217);
nor U14985 (N_14985,N_11892,N_10454);
and U14986 (N_14986,N_10556,N_10892);
nor U14987 (N_14987,N_10636,N_11702);
xor U14988 (N_14988,N_11674,N_11934);
nor U14989 (N_14989,N_12281,N_12194);
nor U14990 (N_14990,N_11895,N_12448);
nor U14991 (N_14991,N_10510,N_10048);
nor U14992 (N_14992,N_11099,N_12050);
or U14993 (N_14993,N_11295,N_10705);
nand U14994 (N_14994,N_10050,N_10659);
and U14995 (N_14995,N_11704,N_10332);
and U14996 (N_14996,N_11540,N_11653);
nand U14997 (N_14997,N_10290,N_11772);
xnor U14998 (N_14998,N_10974,N_10321);
or U14999 (N_14999,N_11437,N_12092);
or U15000 (N_15000,N_13186,N_13110);
and U15001 (N_15001,N_14266,N_13322);
nor U15002 (N_15002,N_12778,N_14500);
and U15003 (N_15003,N_13154,N_13805);
and U15004 (N_15004,N_12743,N_13395);
nor U15005 (N_15005,N_14768,N_13712);
nor U15006 (N_15006,N_12735,N_13949);
nand U15007 (N_15007,N_14193,N_12903);
nor U15008 (N_15008,N_12622,N_14561);
or U15009 (N_15009,N_13878,N_12900);
and U15010 (N_15010,N_12727,N_13102);
nand U15011 (N_15011,N_14424,N_13737);
and U15012 (N_15012,N_14603,N_12546);
nand U15013 (N_15013,N_14051,N_13830);
xor U15014 (N_15014,N_14939,N_13937);
and U15015 (N_15015,N_14822,N_13926);
xor U15016 (N_15016,N_14435,N_12698);
xnor U15017 (N_15017,N_14735,N_13918);
xnor U15018 (N_15018,N_14781,N_12607);
nor U15019 (N_15019,N_14619,N_14226);
nand U15020 (N_15020,N_12838,N_14810);
or U15021 (N_15021,N_14366,N_14802);
and U15022 (N_15022,N_14682,N_13515);
nor U15023 (N_15023,N_14380,N_13270);
or U15024 (N_15024,N_14972,N_13351);
nand U15025 (N_15025,N_13132,N_14031);
xor U15026 (N_15026,N_13907,N_13657);
nor U15027 (N_15027,N_14512,N_14940);
xor U15028 (N_15028,N_12979,N_13751);
xnor U15029 (N_15029,N_14566,N_14182);
and U15030 (N_15030,N_12664,N_14184);
nor U15031 (N_15031,N_14362,N_13084);
xor U15032 (N_15032,N_12609,N_14992);
nor U15033 (N_15033,N_13250,N_14683);
and U15034 (N_15034,N_13734,N_14626);
nand U15035 (N_15035,N_14263,N_13310);
and U15036 (N_15036,N_14705,N_14841);
nor U15037 (N_15037,N_12887,N_14149);
xor U15038 (N_15038,N_13095,N_14658);
xor U15039 (N_15039,N_14976,N_13984);
or U15040 (N_15040,N_14487,N_13879);
nor U15041 (N_15041,N_13632,N_12804);
nand U15042 (N_15042,N_13890,N_12644);
nand U15043 (N_15043,N_14472,N_14058);
and U15044 (N_15044,N_14563,N_14886);
nor U15045 (N_15045,N_13855,N_12898);
nand U15046 (N_15046,N_12686,N_12848);
nor U15047 (N_15047,N_13847,N_13628);
and U15048 (N_15048,N_14686,N_14309);
and U15049 (N_15049,N_13498,N_13278);
xor U15050 (N_15050,N_13073,N_13086);
and U15051 (N_15051,N_14722,N_13802);
nand U15052 (N_15052,N_14891,N_13258);
nor U15053 (N_15053,N_14475,N_14406);
and U15054 (N_15054,N_14013,N_13414);
and U15055 (N_15055,N_14957,N_14291);
xnor U15056 (N_15056,N_14392,N_13396);
xor U15057 (N_15057,N_13425,N_12982);
or U15058 (N_15058,N_14355,N_12562);
and U15059 (N_15059,N_13538,N_14079);
and U15060 (N_15060,N_14648,N_14896);
nor U15061 (N_15061,N_14174,N_12542);
and U15062 (N_15062,N_14229,N_13156);
nand U15063 (N_15063,N_14697,N_13402);
or U15064 (N_15064,N_12933,N_14926);
nand U15065 (N_15065,N_14847,N_14173);
or U15066 (N_15066,N_14457,N_14659);
nor U15067 (N_15067,N_14170,N_14937);
xor U15068 (N_15068,N_13493,N_13374);
xnor U15069 (N_15069,N_12864,N_13481);
xor U15070 (N_15070,N_12641,N_14812);
and U15071 (N_15071,N_13016,N_14503);
xnor U15072 (N_15072,N_14534,N_12591);
nand U15073 (N_15073,N_14752,N_14430);
nand U15074 (N_15074,N_13832,N_14140);
nor U15075 (N_15075,N_12732,N_12714);
and U15076 (N_15076,N_12565,N_12932);
nor U15077 (N_15077,N_12974,N_13764);
xor U15078 (N_15078,N_14642,N_13383);
nor U15079 (N_15079,N_14879,N_13698);
or U15080 (N_15080,N_13298,N_12695);
and U15081 (N_15081,N_14832,N_14462);
xor U15082 (N_15082,N_12750,N_12598);
or U15083 (N_15083,N_13811,N_14662);
xor U15084 (N_15084,N_14025,N_13637);
or U15085 (N_15085,N_14459,N_14617);
and U15086 (N_15086,N_14265,N_12703);
or U15087 (N_15087,N_14733,N_13381);
nand U15088 (N_15088,N_14687,N_13329);
or U15089 (N_15089,N_13333,N_13041);
and U15090 (N_15090,N_14456,N_13638);
and U15091 (N_15091,N_14502,N_12883);
and U15092 (N_15092,N_13806,N_13605);
nand U15093 (N_15093,N_14077,N_13813);
nand U15094 (N_15094,N_14283,N_12919);
and U15095 (N_15095,N_13226,N_14298);
xor U15096 (N_15096,N_14168,N_12529);
nand U15097 (N_15097,N_14312,N_13865);
or U15098 (N_15098,N_14023,N_14734);
xor U15099 (N_15099,N_14531,N_14273);
nand U15100 (N_15100,N_14093,N_13793);
and U15101 (N_15101,N_12999,N_13417);
or U15102 (N_15102,N_13145,N_14047);
nor U15103 (N_15103,N_14147,N_13025);
or U15104 (N_15104,N_14506,N_13265);
nor U15105 (N_15105,N_12771,N_13319);
nand U15106 (N_15106,N_13761,N_12923);
nand U15107 (N_15107,N_13560,N_14954);
xor U15108 (N_15108,N_14723,N_13662);
or U15109 (N_15109,N_13267,N_14056);
xor U15110 (N_15110,N_14755,N_13977);
nand U15111 (N_15111,N_14836,N_14578);
nor U15112 (N_15112,N_13910,N_14152);
or U15113 (N_15113,N_14910,N_12726);
and U15114 (N_15114,N_14460,N_14809);
nor U15115 (N_15115,N_13990,N_12926);
xnor U15116 (N_15116,N_12780,N_13993);
nor U15117 (N_15117,N_13519,N_14767);
nor U15118 (N_15118,N_12696,N_14119);
and U15119 (N_15119,N_12573,N_14092);
and U15120 (N_15120,N_13624,N_14553);
and U15121 (N_15121,N_13777,N_14053);
and U15122 (N_15122,N_14924,N_14772);
and U15123 (N_15123,N_14632,N_12613);
nand U15124 (N_15124,N_12527,N_14038);
and U15125 (N_15125,N_12840,N_14613);
nand U15126 (N_15126,N_14669,N_12540);
or U15127 (N_15127,N_13211,N_14412);
or U15128 (N_15128,N_14465,N_14318);
or U15129 (N_15129,N_14766,N_13924);
xnor U15130 (N_15130,N_14749,N_12803);
nor U15131 (N_15131,N_12504,N_13405);
nand U15132 (N_15132,N_13376,N_12774);
nor U15133 (N_15133,N_12597,N_14702);
xor U15134 (N_15134,N_14605,N_12998);
nor U15135 (N_15135,N_12841,N_14679);
or U15136 (N_15136,N_14271,N_13053);
or U15137 (N_15137,N_14095,N_13429);
nand U15138 (N_15138,N_14712,N_13610);
nand U15139 (N_15139,N_13261,N_13942);
and U15140 (N_15140,N_12619,N_14858);
nor U15141 (N_15141,N_14145,N_13994);
and U15142 (N_15142,N_13339,N_12751);
and U15143 (N_15143,N_14082,N_13645);
or U15144 (N_15144,N_13786,N_12501);
nor U15145 (N_15145,N_12618,N_14912);
or U15146 (N_15146,N_13072,N_13240);
nand U15147 (N_15147,N_13553,N_13001);
nor U15148 (N_15148,N_12967,N_13394);
xnor U15149 (N_15149,N_13227,N_14064);
nand U15150 (N_15150,N_14208,N_14970);
and U15151 (N_15151,N_13520,N_14109);
nor U15152 (N_15152,N_14484,N_13087);
or U15153 (N_15153,N_13308,N_13044);
xor U15154 (N_15154,N_14138,N_12801);
nand U15155 (N_15155,N_12675,N_14695);
and U15156 (N_15156,N_12904,N_14044);
and U15157 (N_15157,N_13778,N_13646);
nor U15158 (N_15158,N_12694,N_14532);
and U15159 (N_15159,N_13375,N_14934);
and U15160 (N_15160,N_13530,N_14980);
xor U15161 (N_15161,N_12748,N_14009);
nor U15162 (N_15162,N_13077,N_14432);
and U15163 (N_15163,N_13201,N_14139);
and U15164 (N_15164,N_14215,N_13356);
and U15165 (N_15165,N_14798,N_13100);
or U15166 (N_15166,N_14815,N_14122);
xor U15167 (N_15167,N_14586,N_12506);
xnor U15168 (N_15168,N_13238,N_13194);
or U15169 (N_15169,N_13433,N_13792);
or U15170 (N_15170,N_12868,N_14654);
and U15171 (N_15171,N_13074,N_14762);
and U15172 (N_15172,N_13998,N_12709);
or U15173 (N_15173,N_13683,N_14335);
or U15174 (N_15174,N_13219,N_13244);
nand U15175 (N_15175,N_13281,N_14745);
nor U15176 (N_15176,N_14133,N_14728);
xor U15177 (N_15177,N_14811,N_13930);
nor U15178 (N_15178,N_13835,N_14350);
and U15179 (N_15179,N_13393,N_14482);
or U15180 (N_15180,N_14527,N_13817);
and U15181 (N_15181,N_12781,N_13453);
nor U15182 (N_15182,N_14395,N_12907);
or U15183 (N_15183,N_13531,N_13153);
nand U15184 (N_15184,N_13502,N_13739);
and U15185 (N_15185,N_14376,N_13325);
nand U15186 (N_15186,N_14065,N_14385);
nor U15187 (N_15187,N_12997,N_13328);
or U15188 (N_15188,N_13920,N_14628);
or U15189 (N_15189,N_12881,N_12867);
nor U15190 (N_15190,N_12634,N_13913);
nor U15191 (N_15191,N_14343,N_14630);
or U15192 (N_15192,N_14699,N_14547);
and U15193 (N_15193,N_12543,N_14638);
nor U15194 (N_15194,N_13863,N_14998);
nand U15195 (N_15195,N_12639,N_14657);
nor U15196 (N_15196,N_14339,N_12722);
xnor U15197 (N_15197,N_14540,N_13678);
nor U15198 (N_15198,N_14983,N_13633);
nor U15199 (N_15199,N_14151,N_14245);
nor U15200 (N_15200,N_13845,N_14943);
and U15201 (N_15201,N_12901,N_13972);
xor U15202 (N_15202,N_13247,N_14369);
or U15203 (N_15203,N_13639,N_13691);
nor U15204 (N_15204,N_13634,N_12761);
or U15205 (N_15205,N_14242,N_12912);
nand U15206 (N_15206,N_13583,N_13821);
nor U15207 (N_15207,N_13163,N_14351);
and U15208 (N_15208,N_13602,N_13717);
xor U15209 (N_15209,N_14277,N_13934);
nand U15210 (N_15210,N_13180,N_14279);
and U15211 (N_15211,N_14169,N_13217);
nor U15212 (N_15212,N_13936,N_12582);
nor U15213 (N_15213,N_14608,N_14902);
or U15214 (N_15214,N_13781,N_14663);
or U15215 (N_15215,N_12844,N_14743);
xnor U15216 (N_15216,N_13135,N_14227);
or U15217 (N_15217,N_13164,N_14288);
xor U15218 (N_15218,N_14377,N_14548);
xnor U15219 (N_15219,N_13331,N_13545);
nor U15220 (N_15220,N_12990,N_12757);
xnor U15221 (N_15221,N_14769,N_13853);
nand U15222 (N_15222,N_14904,N_14823);
nor U15223 (N_15223,N_13916,N_14741);
or U15224 (N_15224,N_14621,N_14523);
and U15225 (N_15225,N_12853,N_14602);
nand U15226 (N_15226,N_13588,N_13723);
and U15227 (N_15227,N_14337,N_13800);
or U15228 (N_15228,N_13663,N_14916);
or U15229 (N_15229,N_13134,N_14796);
nor U15230 (N_15230,N_14320,N_13214);
and U15231 (N_15231,N_14834,N_14496);
or U15232 (N_15232,N_14282,N_14570);
nor U15233 (N_15233,N_12986,N_13293);
nand U15234 (N_15234,N_14718,N_13000);
nand U15235 (N_15235,N_12627,N_13886);
and U15236 (N_15236,N_14311,N_14901);
nor U15237 (N_15237,N_13565,N_12966);
and U15238 (N_15238,N_14596,N_14678);
or U15239 (N_15239,N_13479,N_12895);
nand U15240 (N_15240,N_14756,N_14293);
or U15241 (N_15241,N_13911,N_14454);
and U15242 (N_15242,N_12524,N_14297);
xor U15243 (N_15243,N_14782,N_14421);
nor U15244 (N_15244,N_13722,N_13148);
nand U15245 (N_15245,N_14765,N_13131);
nor U15246 (N_15246,N_13980,N_12776);
and U15247 (N_15247,N_14923,N_12813);
nor U15248 (N_15248,N_14063,N_12739);
nor U15249 (N_15249,N_13507,N_14685);
nand U15250 (N_15250,N_14330,N_13345);
or U15251 (N_15251,N_13669,N_14719);
and U15252 (N_15252,N_13872,N_14061);
xnor U15253 (N_15253,N_13208,N_12585);
and U15254 (N_15254,N_12855,N_14116);
or U15255 (N_15255,N_14352,N_14439);
xnor U15256 (N_15256,N_12516,N_14994);
xnor U15257 (N_15257,N_13141,N_13031);
and U15258 (N_15258,N_13048,N_12560);
nand U15259 (N_15259,N_14759,N_14449);
nand U15260 (N_15260,N_13590,N_14448);
nor U15261 (N_15261,N_13315,N_14130);
xor U15262 (N_15262,N_12687,N_14990);
xor U15263 (N_15263,N_14304,N_12545);
and U15264 (N_15264,N_12947,N_13917);
nand U15265 (N_15265,N_14565,N_13754);
or U15266 (N_15266,N_14470,N_13415);
nand U15267 (N_15267,N_13313,N_14520);
and U15268 (N_15268,N_14709,N_13796);
nor U15269 (N_15269,N_12720,N_14526);
and U15270 (N_15270,N_14591,N_14236);
xnor U15271 (N_15271,N_14046,N_13651);
or U15272 (N_15272,N_13528,N_13978);
and U15273 (N_15273,N_12580,N_13051);
nand U15274 (N_15274,N_13883,N_13659);
nor U15275 (N_15275,N_14224,N_14387);
nor U15276 (N_15276,N_14495,N_13787);
nand U15277 (N_15277,N_13511,N_13670);
nor U15278 (N_15278,N_14711,N_13416);
and U15279 (N_15279,N_14597,N_13488);
xor U15280 (N_15280,N_14689,N_14622);
nor U15281 (N_15281,N_13501,N_14577);
nor U15282 (N_15282,N_13504,N_14704);
nand U15283 (N_15283,N_14404,N_14529);
and U15284 (N_15284,N_13860,N_12921);
nor U15285 (N_15285,N_12817,N_13795);
nand U15286 (N_15286,N_13305,N_13005);
or U15287 (N_15287,N_14217,N_14600);
nand U15288 (N_15288,N_13704,N_13594);
and U15289 (N_15289,N_14251,N_12526);
nand U15290 (N_15290,N_13388,N_13815);
xor U15291 (N_15291,N_14838,N_12793);
nor U15292 (N_15292,N_13411,N_13367);
or U15293 (N_15293,N_13940,N_14157);
nand U15294 (N_15294,N_14096,N_13181);
nand U15295 (N_15295,N_14108,N_14931);
or U15296 (N_15296,N_14447,N_14115);
xnor U15297 (N_15297,N_13775,N_13713);
nor U15298 (N_15298,N_13970,N_13486);
or U15299 (N_15299,N_14442,N_13126);
nand U15300 (N_15300,N_12831,N_13033);
nor U15301 (N_15301,N_14588,N_13640);
xor U15302 (N_15302,N_13973,N_13446);
nor U15303 (N_15303,N_13252,N_13757);
and U15304 (N_15304,N_14515,N_12617);
xor U15305 (N_15305,N_14666,N_14325);
xor U15306 (N_15306,N_14007,N_14285);
xor U15307 (N_15307,N_14249,N_12699);
and U15308 (N_15308,N_12683,N_13695);
nor U15309 (N_15309,N_13080,N_14198);
or U15310 (N_15310,N_14250,N_13321);
nand U15311 (N_15311,N_14189,N_13312);
or U15312 (N_15312,N_13516,N_13706);
or U15313 (N_15313,N_12507,N_14473);
nand U15314 (N_15314,N_13123,N_14346);
xnor U15315 (N_15315,N_13062,N_12615);
nand U15316 (N_15316,N_14885,N_13473);
or U15317 (N_15317,N_14476,N_13716);
and U15318 (N_15318,N_14107,N_13071);
or U15319 (N_15319,N_12837,N_13841);
or U15320 (N_15320,N_12691,N_12632);
nand U15321 (N_15321,N_12711,N_14211);
nand U15322 (N_15322,N_14196,N_13901);
nand U15323 (N_15323,N_13412,N_12812);
and U15324 (N_15324,N_13850,N_12861);
xor U15325 (N_15325,N_14358,N_14589);
or U15326 (N_15326,N_12595,N_14892);
or U15327 (N_15327,N_13579,N_14490);
nand U15328 (N_15328,N_14505,N_12769);
or U15329 (N_15329,N_12706,N_13589);
nor U15330 (N_15330,N_13692,N_14895);
and U15331 (N_15331,N_13159,N_14787);
or U15332 (N_15332,N_12672,N_13810);
nand U15333 (N_15333,N_13665,N_14431);
or U15334 (N_15334,N_13463,N_12559);
nand U15335 (N_15335,N_14579,N_14386);
or U15336 (N_15336,N_14461,N_13643);
nand U15337 (N_15337,N_14156,N_12952);
xor U15338 (N_15338,N_13253,N_14212);
nand U15339 (N_15339,N_13581,N_12969);
nor U15340 (N_15340,N_14870,N_12878);
and U15341 (N_15341,N_14111,N_13089);
and U15342 (N_15342,N_13785,N_14536);
nand U15343 (N_15343,N_14960,N_12563);
nand U15344 (N_15344,N_13763,N_14706);
and U15345 (N_15345,N_12625,N_13045);
or U15346 (N_15346,N_12719,N_14786);
or U15347 (N_15347,N_13797,N_14422);
or U15348 (N_15348,N_13999,N_14326);
or U15349 (N_15349,N_13184,N_14135);
or U15350 (N_15350,N_14067,N_14004);
nand U15351 (N_15351,N_14598,N_13218);
nor U15352 (N_15352,N_14855,N_13812);
and U15353 (N_15353,N_14868,N_13272);
or U15354 (N_15354,N_13648,N_13483);
nand U15355 (N_15355,N_13569,N_14090);
xor U15356 (N_15356,N_14464,N_13894);
or U15357 (N_15357,N_12610,N_13213);
xnor U15358 (N_15358,N_14006,N_12800);
nand U15359 (N_15359,N_12535,N_13022);
or U15360 (N_15360,N_13036,N_13465);
or U15361 (N_15361,N_14480,N_14037);
nor U15362 (N_15362,N_14732,N_14202);
or U15363 (N_15363,N_12785,N_14367);
nor U15364 (N_15364,N_13303,N_14969);
and U15365 (N_15365,N_14729,N_14036);
nand U15366 (N_15366,N_12522,N_14877);
nor U15367 (N_15367,N_13058,N_13011);
nand U15368 (N_15368,N_12816,N_14979);
and U15369 (N_15369,N_13040,N_12910);
nand U15370 (N_15370,N_13615,N_14019);
xnor U15371 (N_15371,N_14008,N_12980);
or U15372 (N_15372,N_14074,N_14143);
and U15373 (N_15373,N_12984,N_14308);
or U15374 (N_15374,N_12658,N_12541);
nand U15375 (N_15375,N_14106,N_12624);
nand U15376 (N_15376,N_12949,N_14200);
xnor U15377 (N_15377,N_12572,N_13391);
and U15378 (N_15378,N_12890,N_14268);
and U15379 (N_15379,N_13431,N_13686);
nor U15380 (N_15380,N_12889,N_13408);
nand U15381 (N_15381,N_14821,N_13275);
or U15382 (N_15382,N_13870,N_13378);
and U15383 (N_15383,N_14649,N_14777);
and U15384 (N_15384,N_13401,N_12943);
xnor U15385 (N_15385,N_14947,N_13578);
nand U15386 (N_15386,N_13893,N_14113);
and U15387 (N_15387,N_14725,N_14022);
nand U15388 (N_15388,N_14651,N_12608);
nand U15389 (N_15389,N_13818,N_12849);
nor U15390 (N_15390,N_13789,N_12832);
nand U15391 (N_15391,N_13028,N_14477);
nand U15392 (N_15392,N_13107,N_13057);
nor U15393 (N_15393,N_12987,N_13149);
xor U15394 (N_15394,N_14830,N_12682);
or U15395 (N_15395,N_13838,N_14129);
nand U15396 (N_15396,N_14562,N_12937);
or U15397 (N_15397,N_14382,N_12941);
or U15398 (N_15398,N_13491,N_14825);
nor U15399 (N_15399,N_14999,N_14295);
xnor U15400 (N_15400,N_12668,N_13361);
nand U15401 (N_15401,N_13963,N_13434);
xnor U15402 (N_15402,N_13284,N_13108);
and U15403 (N_15403,N_14073,N_14889);
or U15404 (N_15404,N_13768,N_13803);
and U15405 (N_15405,N_13353,N_13948);
nand U15406 (N_15406,N_14123,N_14427);
nand U15407 (N_15407,N_12620,N_12554);
or U15408 (N_15408,N_14555,N_14329);
or U15409 (N_15409,N_14340,N_13851);
nor U15410 (N_15410,N_14039,N_13944);
nand U15411 (N_15411,N_13038,N_13241);
nand U15412 (N_15412,N_14347,N_14650);
nor U15413 (N_15413,N_13008,N_13599);
and U15414 (N_15414,N_12946,N_13547);
nor U15415 (N_15415,N_14593,N_13466);
and U15416 (N_15416,N_13666,N_12708);
or U15417 (N_15417,N_13889,N_14917);
nor U15418 (N_15418,N_13960,N_13840);
nand U15419 (N_15419,N_14055,N_13617);
xnor U15420 (N_15420,N_13199,N_12570);
xnor U15421 (N_15421,N_12825,N_14606);
nor U15422 (N_15422,N_14091,N_13982);
and U15423 (N_15423,N_13891,N_12530);
and U15424 (N_15424,N_13532,N_13232);
and U15425 (N_15425,N_12718,N_14963);
or U15426 (N_15426,N_13454,N_13090);
nor U15427 (N_15427,N_14042,N_12762);
nand U15428 (N_15428,N_14903,N_14919);
nand U15429 (N_15429,N_13623,N_14209);
nor U15430 (N_15430,N_13554,N_14195);
xnor U15431 (N_15431,N_14610,N_14966);
or U15432 (N_15432,N_14882,N_14296);
and U15433 (N_15433,N_14574,N_14788);
or U15434 (N_15434,N_14513,N_13189);
xnor U15435 (N_15435,N_12942,N_12772);
and U15436 (N_15436,N_13826,N_14831);
nand U15437 (N_15437,N_13603,N_14290);
nand U15438 (N_15438,N_14636,N_13575);
nand U15439 (N_15439,N_13869,N_14255);
xnor U15440 (N_15440,N_12577,N_12944);
nor U15441 (N_15441,N_13492,N_14517);
nor U15442 (N_15442,N_14178,N_12725);
nand U15443 (N_15443,N_13458,N_13816);
nor U15444 (N_15444,N_13738,N_12651);
and U15445 (N_15445,N_13043,N_13030);
nor U15446 (N_15446,N_13721,N_14700);
nand U15447 (N_15447,N_14911,N_13567);
and U15448 (N_15448,N_13544,N_12665);
xor U15449 (N_15449,N_14974,N_14398);
nor U15450 (N_15450,N_14664,N_13675);
nor U15451 (N_15451,N_14890,N_12792);
or U15452 (N_15452,N_14428,N_14192);
xor U15453 (N_15453,N_12767,N_13297);
nand U15454 (N_15454,N_12697,N_12886);
nor U15455 (N_15455,N_14244,N_14501);
nand U15456 (N_15456,N_12531,N_14444);
nor U15457 (N_15457,N_14614,N_14371);
and U15458 (N_15458,N_12700,N_12827);
nor U15459 (N_15459,N_13462,N_13898);
or U15460 (N_15460,N_13302,N_13526);
nand U15461 (N_15461,N_13047,N_14419);
nand U15462 (N_15462,N_14389,N_13584);
xor U15463 (N_15463,N_13067,N_13234);
or U15464 (N_15464,N_12971,N_13546);
nand U15465 (N_15465,N_14751,N_12938);
xor U15466 (N_15466,N_14001,N_13694);
nand U15467 (N_15467,N_12517,N_13200);
and U15468 (N_15468,N_13887,N_14417);
xor U15469 (N_15469,N_14854,N_14467);
nand U15470 (N_15470,N_14322,N_13941);
nor U15471 (N_15471,N_13061,N_13447);
or U15472 (N_15472,N_13981,N_12502);
nand U15473 (N_15473,N_14564,N_13834);
or U15474 (N_15474,N_14101,N_13206);
or U15475 (N_15475,N_12790,N_13193);
nor U15476 (N_15476,N_13996,N_14537);
and U15477 (N_15477,N_14824,N_12765);
xnor U15478 (N_15478,N_14552,N_14443);
or U15479 (N_15479,N_14445,N_13573);
nand U15480 (N_15480,N_14738,N_14846);
nor U15481 (N_15481,N_13566,N_13334);
and U15482 (N_15482,N_14860,N_13032);
and U15483 (N_15483,N_14909,N_13014);
and U15484 (N_15484,N_14887,N_13956);
nand U15485 (N_15485,N_12862,N_12896);
and U15486 (N_15486,N_14763,N_12809);
xnor U15487 (N_15487,N_14356,N_13731);
nor U15488 (N_15488,N_13188,N_12603);
or U15489 (N_15489,N_12555,N_14844);
xor U15490 (N_15490,N_14900,N_13460);
nor U15491 (N_15491,N_14437,N_14070);
xnor U15492 (N_15492,N_13760,N_13056);
and U15493 (N_15493,N_14744,N_14011);
nor U15494 (N_15494,N_14816,N_12972);
xor U15495 (N_15495,N_13083,N_13562);
nand U15496 (N_15496,N_13324,N_13748);
nand U15497 (N_15497,N_14511,N_12717);
xnor U15498 (N_15498,N_12532,N_12660);
or U15499 (N_15499,N_13745,N_13006);
nand U15500 (N_15500,N_13668,N_13702);
and U15501 (N_15501,N_14270,N_14615);
and U15502 (N_15502,N_13260,N_13660);
or U15503 (N_15503,N_14086,N_13344);
and U15504 (N_15504,N_14066,N_13158);
xor U15505 (N_15505,N_14235,N_12604);
xnor U15506 (N_15506,N_14803,N_13825);
or U15507 (N_15507,N_12839,N_13958);
xor U15508 (N_15508,N_14967,N_14584);
and U15509 (N_15509,N_14665,N_13866);
or U15510 (N_15510,N_12593,N_13882);
and U15511 (N_15511,N_14724,N_12742);
nand U15512 (N_15512,N_12806,N_13457);
nand U15513 (N_15513,N_13952,N_13557);
or U15514 (N_15514,N_13836,N_13183);
nand U15515 (N_15515,N_13833,N_14188);
nor U15516 (N_15516,N_14869,N_13468);
and U15517 (N_15517,N_13551,N_13535);
xnor U15518 (N_15518,N_14713,N_14201);
or U15519 (N_15519,N_14349,N_13065);
or U15520 (N_15520,N_14897,N_12755);
xor U15521 (N_15521,N_12643,N_13221);
nand U15522 (N_15522,N_14862,N_12842);
or U15523 (N_15523,N_14426,N_13561);
nand U15524 (N_15524,N_14021,N_14571);
nor U15525 (N_15525,N_12836,N_14819);
or U15526 (N_15526,N_12959,N_13185);
xor U15527 (N_15527,N_13861,N_12847);
nor U15528 (N_15528,N_13403,N_14493);
and U15529 (N_15529,N_13814,N_13349);
or U15530 (N_15530,N_13112,N_13309);
nand U15531 (N_15531,N_14372,N_14218);
nand U15532 (N_15532,N_13727,N_12548);
nand U15533 (N_15533,N_13155,N_14690);
or U15534 (N_15534,N_13330,N_13983);
nor U15535 (N_15535,N_14549,N_12770);
and U15536 (N_15536,N_14252,N_14867);
nor U15537 (N_15537,N_13782,N_14098);
nor U15538 (N_15538,N_13513,N_14027);
xnor U15539 (N_15539,N_13004,N_14436);
xor U15540 (N_15540,N_12656,N_13327);
and U15541 (N_15541,N_14453,N_14225);
nor U15542 (N_15542,N_13875,N_14094);
or U15543 (N_15543,N_12623,N_14985);
or U15544 (N_15544,N_14012,N_13974);
and U15545 (N_15545,N_14797,N_13222);
or U15546 (N_15546,N_14975,N_14083);
or U15547 (N_15547,N_13390,N_12807);
or U15548 (N_15548,N_13233,N_14345);
and U15549 (N_15549,N_13224,N_14300);
xnor U15550 (N_15550,N_13109,N_14546);
nand U15551 (N_15551,N_14582,N_13054);
xor U15552 (N_15552,N_12536,N_14873);
xnor U15553 (N_15553,N_14522,N_13740);
xnor U15554 (N_15554,N_14175,N_12551);
xnor U15555 (N_15555,N_14671,N_13759);
or U15556 (N_15556,N_14441,N_14374);
or U15557 (N_15557,N_13558,N_12876);
nor U15558 (N_15558,N_14378,N_12666);
or U15559 (N_15559,N_13791,N_13876);
nor U15560 (N_15560,N_13762,N_12915);
nor U15561 (N_15561,N_13550,N_13017);
xnor U15562 (N_15562,N_14936,N_13859);
nor U15563 (N_15563,N_13995,N_12788);
xor U15564 (N_15564,N_14524,N_12519);
nor U15565 (N_15565,N_13652,N_12823);
nand U15566 (N_15566,N_13497,N_12830);
xor U15567 (N_15567,N_13644,N_14866);
xnor U15568 (N_15568,N_13771,N_14692);
or U15569 (N_15569,N_14958,N_14826);
nor U15570 (N_15570,N_13225,N_14396);
nor U15571 (N_15571,N_14757,N_13746);
or U15572 (N_15572,N_13294,N_13326);
nand U15573 (N_15573,N_12583,N_12851);
xor U15574 (N_15574,N_14315,N_14518);
nor U15575 (N_15575,N_13961,N_14469);
nor U15576 (N_15576,N_14360,N_13173);
nand U15577 (N_15577,N_14416,N_13207);
nor U15578 (N_15578,N_13755,N_14136);
xor U15579 (N_15579,N_14907,N_13205);
xor U15580 (N_15580,N_13162,N_13177);
nand U15581 (N_15581,N_14206,N_12843);
or U15582 (N_15582,N_13824,N_14760);
and U15583 (N_15583,N_13563,N_12596);
nand U15584 (N_15584,N_12779,N_13059);
and U15585 (N_15585,N_12983,N_12599);
and U15586 (N_15586,N_13667,N_12721);
and U15587 (N_15587,N_13255,N_14394);
nor U15588 (N_15588,N_13939,N_12549);
nand U15589 (N_15589,N_14035,N_12701);
or U15590 (N_15590,N_14057,N_13042);
xnor U15591 (N_15591,N_12865,N_13280);
nand U15592 (N_15592,N_12539,N_14590);
xnor U15593 (N_15593,N_13574,N_13518);
or U15594 (N_15594,N_14471,N_13867);
xor U15595 (N_15595,N_13626,N_13864);
and U15596 (N_15596,N_13398,N_13690);
nor U15597 (N_15597,N_13279,N_13441);
nand U15598 (N_15598,N_13407,N_14986);
nand U15599 (N_15599,N_13078,N_13400);
xnor U15600 (N_15600,N_13092,N_13827);
xor U15601 (N_15601,N_13175,N_12601);
nand U15602 (N_15602,N_14514,N_13066);
nor U15603 (N_15603,N_13957,N_14307);
or U15604 (N_15604,N_14951,N_13929);
and U15605 (N_15605,N_12574,N_14468);
or U15606 (N_15606,N_13317,N_14219);
nor U15607 (N_15607,N_14029,N_13242);
or U15608 (N_15608,N_13655,N_13992);
xnor U15609 (N_15609,N_13075,N_14328);
nand U15610 (N_15610,N_13783,N_12693);
nor U15611 (N_15611,N_14808,N_12951);
nor U15612 (N_15612,N_14996,N_13621);
nand U15613 (N_15613,N_13277,N_13210);
or U15614 (N_15614,N_13262,N_12586);
nand U15615 (N_15615,N_14016,N_14408);
nor U15616 (N_15616,N_12612,N_13069);
nand U15617 (N_15617,N_14783,N_12931);
and U15618 (N_15618,N_14914,N_12892);
xor U15619 (N_15619,N_14117,N_13572);
or U15620 (N_15620,N_14932,N_14921);
or U15621 (N_15621,N_14631,N_14569);
nand U15622 (N_15622,N_13003,N_13534);
or U15623 (N_15623,N_12602,N_12970);
nor U15624 (N_15624,N_13172,N_13650);
nand U15625 (N_15625,N_12616,N_14587);
xnor U15626 (N_15626,N_14258,N_13854);
nand U15627 (N_15627,N_14388,N_13050);
nand U15628 (N_15628,N_13143,N_14221);
nand U15629 (N_15629,N_13971,N_14278);
nand U15630 (N_15630,N_13595,N_12799);
and U15631 (N_15631,N_13256,N_14871);
xor U15632 (N_15632,N_14827,N_13475);
nor U15633 (N_15633,N_12828,N_12927);
nor U15634 (N_15634,N_13953,N_13012);
nor U15635 (N_15635,N_13469,N_14373);
xor U15636 (N_15636,N_13082,N_14941);
nand U15637 (N_15637,N_14521,N_13076);
nor U15638 (N_15638,N_12653,N_13607);
nand U15639 (N_15639,N_14248,N_12909);
nor U15640 (N_15640,N_13904,N_13888);
and U15641 (N_15641,N_13604,N_13340);
nand U15642 (N_15642,N_12654,N_14771);
and U15643 (N_15643,N_12723,N_13756);
nor U15644 (N_15644,N_14795,N_14440);
nand U15645 (N_15645,N_14045,N_12858);
xor U15646 (N_15646,N_13780,N_13248);
or U15647 (N_15647,N_14478,N_12661);
nor U15648 (N_15648,N_14127,N_12537);
and U15649 (N_15649,N_14674,N_13007);
xor U15650 (N_15650,N_13341,N_14576);
and U15651 (N_15651,N_14059,N_14888);
or U15652 (N_15652,N_12523,N_12760);
or U15653 (N_15653,N_14479,N_12674);
nand U15654 (N_15654,N_14102,N_12796);
and U15655 (N_15655,N_14601,N_13673);
and U15656 (N_15656,N_13426,N_14141);
xnor U15657 (N_15657,N_14163,N_14232);
or U15658 (N_15658,N_14334,N_13616);
nand U15659 (N_15659,N_14599,N_13899);
nor U15660 (N_15660,N_13151,N_14884);
and U15661 (N_15661,N_14281,N_13478);
nor U15662 (N_15662,N_13807,N_13915);
and U15663 (N_15663,N_13286,N_14483);
nand U15664 (N_15664,N_14410,N_13360);
nand U15665 (N_15665,N_14499,N_12670);
xor U15666 (N_15666,N_12592,N_14927);
and U15667 (N_15667,N_12764,N_14099);
or U15668 (N_15668,N_13570,N_14541);
xor U15669 (N_15669,N_13943,N_14289);
nand U15670 (N_15670,N_14929,N_13707);
xnor U15671 (N_15671,N_13456,N_12925);
or U15672 (N_15672,N_14993,N_13674);
and U15673 (N_15673,N_13452,N_12885);
nor U15674 (N_15674,N_13438,N_13608);
nand U15675 (N_15675,N_12635,N_13338);
or U15676 (N_15676,N_14731,N_14354);
xor U15677 (N_15677,N_13052,N_13413);
nor U15678 (N_15678,N_14616,N_14321);
xor U15679 (N_15679,N_13139,N_13099);
nor U15680 (N_15680,N_13711,N_13965);
or U15681 (N_15681,N_13552,N_14627);
or U15682 (N_15682,N_14861,N_14407);
and U15683 (N_15683,N_14736,N_14162);
nor U15684 (N_15684,N_14849,N_14859);
and U15685 (N_15685,N_14661,N_12628);
or U15686 (N_15686,N_13938,N_13529);
or U15687 (N_15687,N_13348,N_14714);
nor U15688 (N_15688,N_14655,N_12880);
or U15689 (N_15689,N_13923,N_14420);
nand U15690 (N_15690,N_13630,N_13564);
nand U15691 (N_15691,N_13122,N_14609);
and U15692 (N_15692,N_13203,N_13753);
xor U15693 (N_15693,N_14383,N_12505);
nand U15694 (N_15694,N_14949,N_13880);
nand U15695 (N_15695,N_13366,N_13510);
xnor U15696 (N_15696,N_14612,N_13013);
nand U15697 (N_15697,N_12857,N_14539);
nand U15698 (N_15698,N_14332,N_14171);
nor U15699 (N_15699,N_12513,N_14804);
and U15700 (N_15700,N_14852,N_13735);
nand U15701 (N_15701,N_13820,N_13091);
xnor U15702 (N_15702,N_13140,N_13912);
nand U15703 (N_15703,N_12514,N_14839);
nand U15704 (N_15704,N_13450,N_12647);
or U15705 (N_15705,N_13470,N_13455);
or U15706 (N_15706,N_14556,N_13467);
or U15707 (N_15707,N_14186,N_12977);
xnor U15708 (N_15708,N_14458,N_12600);
or U15709 (N_15709,N_13612,N_13724);
and U15710 (N_15710,N_13397,N_13658);
nand U15711 (N_15711,N_13664,N_14843);
xor U15712 (N_15712,N_13976,N_13598);
xor U15713 (N_15713,N_13523,N_13461);
nor U15714 (N_15714,N_14306,N_13142);
nand U15715 (N_15715,N_13766,N_13779);
and U15716 (N_15716,N_14629,N_13424);
and U15717 (N_15717,N_13220,N_14179);
nand U15718 (N_15718,N_14327,N_12914);
or U15719 (N_15719,N_13732,N_14833);
or U15720 (N_15720,N_14237,N_14853);
nand U15721 (N_15721,N_13176,N_14401);
or U15722 (N_15722,N_12707,N_13606);
nand U15723 (N_15723,N_12820,N_12854);
nand U15724 (N_15724,N_12655,N_14348);
nor U15725 (N_15725,N_14260,N_12978);
nor U15726 (N_15726,N_14807,N_12834);
xor U15727 (N_15727,N_12588,N_13451);
xor U15728 (N_15728,N_13582,N_13288);
xnor U15729 (N_15729,N_13254,N_14172);
and U15730 (N_15730,N_13150,N_12775);
and U15731 (N_15731,N_12510,N_14411);
or U15732 (N_15732,N_14688,N_13198);
and U15733 (N_15733,N_13986,N_13121);
and U15734 (N_15734,N_13116,N_13427);
xor U15735 (N_15735,N_13494,N_13037);
nand U15736 (N_15736,N_12684,N_14088);
or U15737 (N_15737,N_13962,N_13120);
xor U15738 (N_15738,N_12567,N_14062);
nand U15739 (N_15739,N_12652,N_14041);
xor U15740 (N_15740,N_13620,N_14933);
nand U15741 (N_15741,N_14210,N_13024);
xor U15742 (N_15742,N_13568,N_14492);
nand U15743 (N_15743,N_14778,N_13178);
nand U15744 (N_15744,N_12512,N_14640);
or U15745 (N_15745,N_13527,N_14050);
and U15746 (N_15746,N_13885,N_12960);
or U15747 (N_15747,N_13104,N_14944);
nor U15748 (N_15748,N_12648,N_12879);
xor U15749 (N_15749,N_13117,N_14753);
or U15750 (N_15750,N_13715,N_13306);
xnor U15751 (N_15751,N_13165,N_14187);
nor U15752 (N_15752,N_14125,N_13487);
xor U15753 (N_15753,N_14525,N_14028);
nor U15754 (N_15754,N_12594,N_12621);
xnor U15755 (N_15755,N_13541,N_14384);
nand U15756 (N_15756,N_14359,N_14399);
nand U15757 (N_15757,N_13619,N_13829);
nand U15758 (N_15758,N_13743,N_13436);
and U15759 (N_15759,N_12918,N_14848);
or U15760 (N_15760,N_12902,N_14883);
xnor U15761 (N_15761,N_13389,N_13231);
xor U15762 (N_15762,N_13118,N_12754);
xnor U15763 (N_15763,N_12657,N_13896);
xor U15764 (N_15764,N_13365,N_12752);
and U15765 (N_15765,N_13914,N_14364);
nor U15766 (N_15766,N_12746,N_13799);
and U15767 (N_15767,N_12955,N_12503);
nand U15768 (N_15768,N_14559,N_14754);
nand U15769 (N_15769,N_12869,N_13085);
and U15770 (N_15770,N_13576,N_14105);
xor U15771 (N_15771,N_12822,N_12753);
xor U15772 (N_15772,N_13020,N_14997);
nand U15773 (N_15773,N_13774,N_14267);
nor U15774 (N_15774,N_13215,N_13409);
and U15775 (N_15775,N_13874,N_14652);
nand U15776 (N_15776,N_12797,N_13699);
xnor U15777 (N_15777,N_12899,N_13496);
nor U15778 (N_15778,N_14672,N_12590);
xor U15779 (N_15779,N_13649,N_14681);
nand U15780 (N_15780,N_14390,N_13548);
nor U15781 (N_15781,N_12629,N_12587);
or U15782 (N_15782,N_14434,N_13223);
nor U15783 (N_15783,N_12508,N_13169);
nand U15784 (N_15784,N_14573,N_13432);
nand U15785 (N_15785,N_13370,N_14403);
or U15786 (N_15786,N_14955,N_12908);
nand U15787 (N_15787,N_14842,N_12863);
xor U15788 (N_15788,N_14850,N_14946);
xnor U15789 (N_15789,N_14930,N_14204);
nand U15790 (N_15790,N_14747,N_12534);
or U15791 (N_15791,N_13283,N_14799);
xor U15792 (N_15792,N_13129,N_14393);
or U15793 (N_15793,N_12729,N_13684);
or U15794 (N_15794,N_13296,N_14764);
or U15795 (N_15795,N_13273,N_13063);
nor U15796 (N_15796,N_13420,N_14049);
or U15797 (N_15797,N_14299,N_13537);
nor U15798 (N_15798,N_14792,N_14104);
nand U15799 (N_15799,N_14637,N_13804);
and U15800 (N_15800,N_12936,N_13928);
xor U15801 (N_15801,N_12731,N_13877);
xnor U15802 (N_15802,N_12961,N_13418);
and U15803 (N_15803,N_12733,N_14773);
xor U15804 (N_15804,N_13900,N_14677);
or U15805 (N_15805,N_14301,N_14120);
nor U15806 (N_15806,N_12741,N_13170);
nor U15807 (N_15807,N_13274,N_14857);
xnor U15808 (N_15808,N_14793,N_13146);
xnor U15809 (N_15809,N_13848,N_14342);
or U15810 (N_15810,N_13591,N_14987);
nor U15811 (N_15811,N_12663,N_12710);
nor U15812 (N_15812,N_13357,N_14872);
xnor U15813 (N_15813,N_14071,N_14126);
and U15814 (N_15814,N_14222,N_12811);
and U15815 (N_15815,N_13015,N_13354);
and U15816 (N_15816,N_14150,N_13167);
nand U15817 (N_15817,N_13839,N_12747);
nor U15818 (N_15818,N_14452,N_13239);
or U15819 (N_15819,N_14761,N_12515);
or U15820 (N_15820,N_12758,N_14575);
xnor U15821 (N_15821,N_12829,N_13627);
or U15822 (N_15822,N_13857,N_13776);
xnor U15823 (N_15823,N_14368,N_14875);
nand U15824 (N_15824,N_12988,N_14317);
and U15825 (N_15825,N_14269,N_14784);
or U15826 (N_15826,N_14581,N_14906);
xor U15827 (N_15827,N_13430,N_14474);
nand U15828 (N_15828,N_12728,N_12884);
and U15829 (N_15829,N_13744,N_13701);
and U15830 (N_15830,N_13105,N_12784);
and U15831 (N_15831,N_13975,N_14341);
or U15832 (N_15832,N_14451,N_12680);
nor U15833 (N_15833,N_14361,N_12667);
xnor U15834 (N_15834,N_12662,N_12552);
xor U15835 (N_15835,N_12875,N_12805);
nand U15836 (N_15836,N_13881,N_13229);
xor U15837 (N_15837,N_13742,N_14696);
nor U15838 (N_15838,N_12859,N_14568);
nor U15839 (N_15839,N_13794,N_14670);
nor U15840 (N_15840,N_12940,N_13119);
and U15841 (N_15841,N_14010,N_13714);
nand U15842 (N_15842,N_13685,N_13399);
and U15843 (N_15843,N_14942,N_13517);
nor U15844 (N_15844,N_12561,N_12678);
nor U15845 (N_15845,N_13323,N_13216);
and U15846 (N_15846,N_13259,N_13935);
nand U15847 (N_15847,N_14148,N_13823);
and U15848 (N_15848,N_14002,N_14623);
xnor U15849 (N_15849,N_14925,N_12749);
and U15850 (N_15850,N_14450,N_14893);
xor U15851 (N_15851,N_13113,N_12985);
xnor U15852 (N_15852,N_14336,N_13472);
nand U15853 (N_15853,N_12745,N_12738);
xor U15854 (N_15854,N_14611,N_13856);
nor U15855 (N_15855,N_12579,N_14054);
nand U15856 (N_15856,N_12794,N_13307);
and U15857 (N_15857,N_14257,N_13289);
xor U15858 (N_15858,N_14205,N_13749);
nand U15859 (N_15859,N_14305,N_14913);
nor U15860 (N_15860,N_13873,N_12950);
nand U15861 (N_15861,N_12673,N_13243);
xnor U15862 (N_15862,N_14624,N_14243);
nor U15863 (N_15863,N_14164,N_13371);
nand U15864 (N_15864,N_13555,N_13439);
or U15865 (N_15865,N_13046,N_13202);
nor U15866 (N_15866,N_14805,N_14018);
and U15867 (N_15867,N_12782,N_14239);
nand U15868 (N_15868,N_12789,N_14253);
nor U15869 (N_15869,N_13251,N_13837);
nor U15870 (N_15870,N_14280,N_14716);
and U15871 (N_15871,N_14197,N_13257);
nor U15872 (N_15872,N_14668,N_13521);
or U15873 (N_15873,N_14405,N_12928);
or U15874 (N_15874,N_13474,N_12872);
xnor U15875 (N_15875,N_14415,N_12996);
or U15876 (N_15876,N_13618,N_12773);
or U15877 (N_15877,N_14118,N_12704);
or U15878 (N_15878,N_14181,N_14533);
xor U15879 (N_15879,N_13919,N_12500);
xnor U15880 (N_15880,N_12702,N_13729);
xor U15881 (N_15881,N_14989,N_13765);
nand U15882 (N_15882,N_13710,N_13508);
and U15883 (N_15883,N_13115,N_12556);
or U15884 (N_15884,N_13613,N_13809);
and U15885 (N_15885,N_14707,N_13314);
and U15886 (N_15886,N_12906,N_12677);
nand U15887 (N_15887,N_12581,N_14114);
nor U15888 (N_15888,N_13505,N_13355);
nor U15889 (N_15889,N_13946,N_13539);
and U15890 (N_15890,N_14656,N_13679);
xor U15891 (N_15891,N_14968,N_14894);
xnor U15892 (N_15892,N_13895,N_12642);
nand U15893 (N_15893,N_13846,N_12873);
nand U15894 (N_15894,N_12891,N_13369);
nor U15895 (N_15895,N_14995,N_12689);
nor U15896 (N_15896,N_14489,N_13191);
and U15897 (N_15897,N_12783,N_14880);
and U15898 (N_15898,N_14691,N_14247);
or U15899 (N_15899,N_14413,N_12511);
nor U15900 (N_15900,N_14213,N_14020);
xnor U15901 (N_15901,N_12578,N_12845);
or U15902 (N_15902,N_14837,N_13300);
nand U15903 (N_15903,N_14048,N_12713);
and U15904 (N_15904,N_13377,N_13945);
or U15905 (N_15905,N_12538,N_14604);
and U15906 (N_15906,N_13094,N_13922);
or U15907 (N_15907,N_13587,N_14780);
nor U15908 (N_15908,N_13585,N_13464);
nand U15909 (N_15909,N_13021,N_14177);
or U15910 (N_15910,N_14375,N_13160);
nor U15911 (N_15911,N_14899,N_13019);
nand U15912 (N_15912,N_13533,N_13964);
nor U15913 (N_15913,N_14567,N_14455);
xor U15914 (N_15914,N_12860,N_13106);
and U15915 (N_15915,N_14953,N_14530);
nor U15916 (N_15916,N_13332,N_12948);
nand U15917 (N_15917,N_12525,N_14190);
nor U15918 (N_15918,N_14775,N_12520);
xnor U15919 (N_15919,N_13098,N_12965);
nand U15920 (N_15920,N_14742,N_14863);
xor U15921 (N_15921,N_14081,N_14504);
nor U15922 (N_15922,N_14234,N_13490);
nor U15923 (N_15923,N_14915,N_13600);
nand U15924 (N_15924,N_12866,N_13858);
and U15925 (N_15925,N_12584,N_13212);
and U15926 (N_15926,N_14155,N_14737);
nand U15927 (N_15927,N_13653,N_13733);
nor U15928 (N_15928,N_12736,N_13725);
or U15929 (N_15929,N_14545,N_12833);
nor U15930 (N_15930,N_14425,N_12815);
nor U15931 (N_15931,N_13230,N_12856);
nor U15932 (N_15932,N_12649,N_13884);
or U15933 (N_15933,N_13392,N_13902);
and U15934 (N_15934,N_14864,N_13525);
nor U15935 (N_15935,N_14015,N_14800);
xnor U15936 (N_15936,N_14161,N_14121);
and U15937 (N_15937,N_14103,N_12976);
xor U15938 (N_15938,N_13625,N_13197);
nand U15939 (N_15939,N_13897,N_13741);
nand U15940 (N_15940,N_12991,N_14856);
xor U15941 (N_15941,N_13245,N_13192);
nand U15942 (N_15942,N_14851,N_13459);
and U15943 (N_15943,N_12650,N_14558);
xor U15944 (N_15944,N_14717,N_14779);
xnor U15945 (N_15945,N_14646,N_14580);
and U15946 (N_15946,N_12564,N_14144);
and U15947 (N_15947,N_13635,N_14446);
or U15948 (N_15948,N_13784,N_14262);
or U15949 (N_15949,N_13337,N_14167);
xnor U15950 (N_15950,N_14758,N_13577);
and U15951 (N_15951,N_14216,N_14381);
xor U15952 (N_15952,N_14684,N_14026);
or U15953 (N_15953,N_12993,N_14494);
xnor U15954 (N_15954,N_14550,N_13693);
or U15955 (N_15955,N_12737,N_14344);
and U15956 (N_15956,N_13849,N_12802);
or U15957 (N_15957,N_13967,N_13147);
or U15958 (N_15958,N_14794,N_13304);
and U15959 (N_15959,N_13124,N_12894);
xnor U15960 (N_15960,N_13654,N_14076);
or U15961 (N_15961,N_14363,N_14040);
and U15962 (N_15962,N_14409,N_14982);
nor U15963 (N_15963,N_12716,N_13026);
and U15964 (N_15964,N_14820,N_14097);
and U15965 (N_15965,N_14003,N_13503);
and U15966 (N_15966,N_14981,N_12905);
nor U15967 (N_15967,N_13027,N_14176);
nor U15968 (N_15968,N_13384,N_13422);
and U15969 (N_15969,N_14594,N_13536);
nor U15970 (N_15970,N_14698,N_13363);
and U15971 (N_15971,N_13512,N_13689);
or U15972 (N_15972,N_14554,N_13404);
or U15973 (N_15973,N_14231,N_13647);
and U15974 (N_15974,N_14720,N_14710);
or U15975 (N_15975,N_13237,N_14774);
nand U15976 (N_15976,N_14653,N_14261);
nor U15977 (N_15977,N_13018,N_14284);
and U15978 (N_15978,N_14191,N_14400);
and U15979 (N_15979,N_14078,N_14303);
or U15980 (N_15980,N_13372,N_14959);
or U15981 (N_15981,N_14032,N_12558);
nand U15982 (N_15982,N_13593,N_13444);
nor U15983 (N_15983,N_14633,N_14331);
nor U15984 (N_15984,N_12712,N_13482);
or U15985 (N_15985,N_13509,N_13359);
or U15986 (N_15986,N_12930,N_13580);
nand U15987 (N_15987,N_12945,N_14313);
and U15988 (N_15988,N_13979,N_13892);
and U15989 (N_15989,N_12766,N_12671);
nand U15990 (N_15990,N_13364,N_13114);
nor U15991 (N_15991,N_13540,N_14034);
and U15992 (N_15992,N_13622,N_13111);
nand U15993 (N_15993,N_13991,N_14543);
nand U15994 (N_15994,N_13808,N_14486);
and U15995 (N_15995,N_12724,N_12888);
nand U15996 (N_15996,N_13346,N_12973);
and U15997 (N_15997,N_13290,N_12808);
xor U15998 (N_15998,N_13336,N_13264);
xnor U15999 (N_15999,N_12640,N_13969);
nand U16000 (N_16000,N_14033,N_12631);
nand U16001 (N_16001,N_12688,N_13773);
and U16002 (N_16002,N_14314,N_12669);
nand U16003 (N_16003,N_12550,N_14159);
or U16004 (N_16004,N_13932,N_13386);
or U16005 (N_16005,N_14323,N_14324);
nand U16006 (N_16006,N_14874,N_13471);
nor U16007 (N_16007,N_13697,N_14230);
or U16008 (N_16008,N_13428,N_14418);
nand U16009 (N_16009,N_13641,N_14302);
xor U16010 (N_16010,N_14272,N_13362);
nand U16011 (N_16011,N_13614,N_13718);
and U16012 (N_16012,N_12835,N_14881);
nand U16013 (N_16013,N_13423,N_14072);
nor U16014 (N_16014,N_12756,N_12759);
xnor U16015 (N_16015,N_14319,N_12575);
or U16016 (N_16016,N_13843,N_14703);
nor U16017 (N_16017,N_12533,N_14708);
or U16018 (N_16018,N_14789,N_14551);
xnor U16019 (N_16019,N_13174,N_14014);
and U16020 (N_16020,N_13676,N_12981);
or U16021 (N_16021,N_12553,N_13903);
nor U16022 (N_16022,N_14918,N_13750);
nand U16023 (N_16023,N_14645,N_13182);
xor U16024 (N_16024,N_14806,N_13842);
nor U16025 (N_16025,N_14160,N_13068);
nor U16026 (N_16026,N_12685,N_13291);
or U16027 (N_16027,N_14538,N_12557);
xor U16028 (N_16028,N_14214,N_12681);
and U16029 (N_16029,N_12850,N_13152);
xnor U16030 (N_16030,N_12913,N_14813);
nand U16031 (N_16031,N_12611,N_13542);
xnor U16032 (N_16032,N_14727,N_13959);
or U16033 (N_16033,N_12989,N_12826);
xnor U16034 (N_16034,N_14908,N_14560);
and U16035 (N_16035,N_12734,N_12626);
and U16036 (N_16036,N_13730,N_13772);
xor U16037 (N_16037,N_14770,N_13703);
or U16038 (N_16038,N_14370,N_13009);
xnor U16039 (N_16039,N_13088,N_14516);
nor U16040 (N_16040,N_13133,N_14365);
and U16041 (N_16041,N_13137,N_14085);
nand U16042 (N_16042,N_13263,N_13950);
nand U16043 (N_16043,N_13988,N_13187);
nand U16044 (N_16044,N_14185,N_12962);
xor U16045 (N_16045,N_14276,N_13276);
xor U16046 (N_16046,N_14146,N_12975);
and U16047 (N_16047,N_14693,N_14952);
and U16048 (N_16048,N_12571,N_14510);
or U16049 (N_16049,N_14264,N_14124);
xnor U16050 (N_16050,N_14316,N_14154);
xor U16051 (N_16051,N_14402,N_13292);
nor U16052 (N_16052,N_14286,N_13136);
nand U16053 (N_16053,N_14984,N_12920);
xor U16054 (N_16054,N_13954,N_13769);
xnor U16055 (N_16055,N_13266,N_14748);
nand U16056 (N_16056,N_12939,N_13445);
nor U16057 (N_16057,N_12768,N_13586);
nand U16058 (N_16058,N_13543,N_12568);
nor U16059 (N_16059,N_13705,N_14973);
and U16060 (N_16060,N_12786,N_13822);
nand U16061 (N_16061,N_14991,N_14508);
xor U16062 (N_16062,N_13559,N_14180);
or U16063 (N_16063,N_13514,N_14275);
xor U16064 (N_16064,N_14087,N_14238);
xnor U16065 (N_16065,N_14715,N_14945);
xnor U16066 (N_16066,N_12547,N_13343);
nand U16067 (N_16067,N_12968,N_14100);
or U16068 (N_16068,N_12871,N_13125);
nor U16069 (N_16069,N_14519,N_12814);
nand U16070 (N_16070,N_13299,N_14817);
nand U16071 (N_16071,N_13249,N_14660);
or U16072 (N_16072,N_14978,N_14259);
xor U16073 (N_16073,N_13549,N_14294);
and U16074 (N_16074,N_12715,N_13097);
or U16075 (N_16075,N_12798,N_13629);
xor U16076 (N_16076,N_13927,N_14845);
xnor U16077 (N_16077,N_14739,N_13687);
and U16078 (N_16078,N_13485,N_13871);
xnor U16079 (N_16079,N_12569,N_14840);
nand U16080 (N_16080,N_14287,N_13350);
or U16081 (N_16081,N_14528,N_14542);
xnor U16082 (N_16082,N_14950,N_14043);
nor U16083 (N_16083,N_13320,N_13556);
nor U16084 (N_16084,N_12630,N_12763);
nor U16085 (N_16085,N_13335,N_12544);
or U16086 (N_16086,N_14791,N_13010);
nand U16087 (N_16087,N_12791,N_14680);
and U16088 (N_16088,N_14466,N_14488);
nor U16089 (N_16089,N_13448,N_14052);
nor U16090 (N_16090,N_14491,N_13443);
nand U16091 (N_16091,N_14644,N_13921);
and U16092 (N_16092,N_13495,N_13947);
and U16093 (N_16093,N_14814,N_13642);
nand U16094 (N_16094,N_12882,N_13318);
nor U16095 (N_16095,N_14634,N_14746);
or U16096 (N_16096,N_14977,N_13597);
nand U16097 (N_16097,N_13039,N_14357);
nand U16098 (N_16098,N_14639,N_14507);
xnor U16099 (N_16099,N_14620,N_12637);
and U16100 (N_16100,N_13168,N_14089);
or U16101 (N_16101,N_13301,N_14618);
nor U16102 (N_16102,N_12659,N_14740);
or U16103 (N_16103,N_13034,N_14338);
nand U16104 (N_16104,N_13406,N_13421);
or U16105 (N_16105,N_13093,N_13190);
and U16106 (N_16106,N_14750,N_12992);
nand U16107 (N_16107,N_14835,N_14776);
xnor U16108 (N_16108,N_13908,N_13295);
nor U16109 (N_16109,N_14397,N_13196);
nor U16110 (N_16110,N_14607,N_12528);
nor U16111 (N_16111,N_13596,N_13788);
and U16112 (N_16112,N_13228,N_14132);
or U16113 (N_16113,N_14865,N_13747);
nor U16114 (N_16114,N_14433,N_13440);
xor U16115 (N_16115,N_13798,N_14585);
nor U16116 (N_16116,N_12929,N_14438);
nand U16117 (N_16117,N_13285,N_14905);
or U16118 (N_16118,N_12917,N_13925);
nor U16119 (N_16119,N_14110,N_12645);
xnor U16120 (N_16120,N_12994,N_14165);
xor U16121 (N_16121,N_12576,N_13352);
and U16122 (N_16122,N_14030,N_12810);
and U16123 (N_16123,N_13868,N_13688);
nor U16124 (N_16124,N_14142,N_12818);
or U16125 (N_16125,N_14485,N_13656);
xnor U16126 (N_16126,N_14721,N_12954);
or U16127 (N_16127,N_13955,N_12870);
nand U16128 (N_16128,N_14068,N_14557);
and U16129 (N_16129,N_13671,N_13437);
xor U16130 (N_16130,N_14498,N_14935);
nand U16131 (N_16131,N_13682,N_13101);
and U16132 (N_16132,N_12934,N_13358);
and U16133 (N_16133,N_13592,N_12636);
nor U16134 (N_16134,N_13235,N_14131);
nor U16135 (N_16135,N_13631,N_13828);
and U16136 (N_16136,N_12958,N_13728);
or U16137 (N_16137,N_13720,N_12744);
xor U16138 (N_16138,N_14158,N_14207);
and U16139 (N_16139,N_13752,N_12935);
nor U16140 (N_16140,N_13246,N_14497);
nor U16141 (N_16141,N_14667,N_14228);
nor U16142 (N_16142,N_14965,N_12819);
and U16143 (N_16143,N_13342,N_13103);
nor U16144 (N_16144,N_13571,N_13379);
or U16145 (N_16145,N_13661,N_12787);
or U16146 (N_16146,N_14948,N_13700);
xnor U16147 (N_16147,N_12509,N_13128);
nand U16148 (N_16148,N_14274,N_13029);
and U16149 (N_16149,N_13387,N_13373);
xnor U16150 (N_16150,N_12777,N_14084);
nand U16151 (N_16151,N_14790,N_14509);
or U16152 (N_16152,N_13968,N_12924);
nor U16153 (N_16153,N_12614,N_13906);
xor U16154 (N_16154,N_14818,N_12995);
nand U16155 (N_16155,N_13282,N_12705);
or U16156 (N_16156,N_14194,N_12893);
nor U16157 (N_16157,N_14956,N_13987);
xnor U16158 (N_16158,N_13506,N_14183);
xor U16159 (N_16159,N_13801,N_13382);
or U16160 (N_16160,N_13611,N_13966);
nor U16161 (N_16161,N_12690,N_13144);
and U16162 (N_16162,N_14069,N_13055);
and U16163 (N_16163,N_13997,N_12740);
or U16164 (N_16164,N_14246,N_13347);
nor U16165 (N_16165,N_12605,N_14220);
and U16166 (N_16166,N_14694,N_13166);
nand U16167 (N_16167,N_14635,N_14310);
xnor U16168 (N_16168,N_13677,N_12964);
xor U16169 (N_16169,N_13770,N_14878);
xnor U16170 (N_16170,N_13951,N_14673);
xor U16171 (N_16171,N_13157,N_13524);
xor U16172 (N_16172,N_12679,N_13931);
nand U16173 (N_16173,N_14675,N_12852);
nand U16174 (N_16174,N_14137,N_14641);
nand U16175 (N_16175,N_13171,N_13002);
nand U16176 (N_16176,N_13410,N_14625);
and U16177 (N_16177,N_14333,N_13130);
xor U16178 (N_16178,N_14535,N_12606);
nand U16179 (N_16179,N_12676,N_14876);
nand U16180 (N_16180,N_13905,N_14701);
nand U16181 (N_16181,N_14128,N_14828);
or U16182 (N_16182,N_13268,N_13380);
nor U16183 (N_16183,N_12916,N_14379);
or U16184 (N_16184,N_13909,N_13680);
nand U16185 (N_16185,N_13209,N_13844);
nand U16186 (N_16186,N_13758,N_14233);
and U16187 (N_16187,N_13609,N_14595);
or U16188 (N_16188,N_14254,N_13435);
and U16189 (N_16189,N_14017,N_14112);
nand U16190 (N_16190,N_12566,N_13096);
nor U16191 (N_16191,N_14060,N_13933);
nand U16192 (N_16192,N_13023,N_14647);
or U16193 (N_16193,N_14240,N_12518);
and U16194 (N_16194,N_12821,N_13060);
and U16195 (N_16195,N_13419,N_14643);
nand U16196 (N_16196,N_14592,N_12877);
and U16197 (N_16197,N_13852,N_14971);
and U16198 (N_16198,N_14583,N_12521);
or U16199 (N_16199,N_14391,N_14964);
or U16200 (N_16200,N_13709,N_13790);
xor U16201 (N_16201,N_13049,N_13636);
xnor U16202 (N_16202,N_13204,N_14024);
or U16203 (N_16203,N_14481,N_12897);
nor U16204 (N_16204,N_13271,N_13681);
xnor U16205 (N_16205,N_13862,N_12953);
nor U16206 (N_16206,N_13480,N_14256);
nand U16207 (N_16207,N_14203,N_12638);
nand U16208 (N_16208,N_14080,N_14223);
nand U16209 (N_16209,N_14134,N_13079);
nand U16210 (N_16210,N_13070,N_13127);
nand U16211 (N_16211,N_14785,N_13269);
nor U16212 (N_16212,N_13719,N_12846);
nor U16213 (N_16213,N_14544,N_13989);
nor U16214 (N_16214,N_14730,N_14801);
nor U16215 (N_16215,N_14676,N_14726);
nand U16216 (N_16216,N_13476,N_14829);
xor U16217 (N_16217,N_13449,N_14166);
and U16218 (N_16218,N_14353,N_14988);
nand U16219 (N_16219,N_13708,N_12646);
nand U16220 (N_16220,N_13368,N_13819);
nand U16221 (N_16221,N_12956,N_13179);
and U16222 (N_16222,N_14005,N_13161);
and U16223 (N_16223,N_13035,N_14423);
or U16224 (N_16224,N_12911,N_13385);
xnor U16225 (N_16225,N_14241,N_12922);
nor U16226 (N_16226,N_13311,N_14199);
xnor U16227 (N_16227,N_14429,N_14920);
nor U16228 (N_16228,N_12957,N_13726);
nor U16229 (N_16229,N_13736,N_14928);
nand U16230 (N_16230,N_14000,N_13064);
and U16231 (N_16231,N_12795,N_13442);
xor U16232 (N_16232,N_14153,N_13499);
and U16233 (N_16233,N_12730,N_12824);
xor U16234 (N_16234,N_14898,N_14922);
nor U16235 (N_16235,N_13287,N_13985);
nor U16236 (N_16236,N_13767,N_12874);
or U16237 (N_16237,N_13672,N_13081);
nand U16238 (N_16238,N_13500,N_14938);
or U16239 (N_16239,N_13831,N_12589);
nand U16240 (N_16240,N_13316,N_12692);
xor U16241 (N_16241,N_13477,N_14075);
or U16242 (N_16242,N_14463,N_13522);
xor U16243 (N_16243,N_13195,N_14572);
nor U16244 (N_16244,N_13236,N_14292);
nand U16245 (N_16245,N_13484,N_14414);
and U16246 (N_16246,N_13601,N_12633);
nor U16247 (N_16247,N_13489,N_13696);
xnor U16248 (N_16248,N_14962,N_13138);
and U16249 (N_16249,N_12963,N_14961);
nor U16250 (N_16250,N_12891,N_13707);
or U16251 (N_16251,N_14099,N_13444);
nand U16252 (N_16252,N_14936,N_13607);
nand U16253 (N_16253,N_14052,N_13493);
nand U16254 (N_16254,N_13207,N_14678);
nand U16255 (N_16255,N_12809,N_14365);
and U16256 (N_16256,N_14998,N_14811);
or U16257 (N_16257,N_13853,N_13612);
and U16258 (N_16258,N_14198,N_14454);
and U16259 (N_16259,N_13143,N_13860);
xor U16260 (N_16260,N_12724,N_12974);
and U16261 (N_16261,N_13208,N_12730);
xor U16262 (N_16262,N_12797,N_13531);
and U16263 (N_16263,N_14874,N_13552);
nor U16264 (N_16264,N_13848,N_14359);
xor U16265 (N_16265,N_13560,N_14644);
and U16266 (N_16266,N_14959,N_13190);
or U16267 (N_16267,N_12530,N_14813);
xnor U16268 (N_16268,N_13047,N_12933);
nor U16269 (N_16269,N_13816,N_13976);
nand U16270 (N_16270,N_13570,N_14329);
or U16271 (N_16271,N_12870,N_14297);
nor U16272 (N_16272,N_13639,N_13211);
xnor U16273 (N_16273,N_14153,N_14555);
or U16274 (N_16274,N_13360,N_13845);
nor U16275 (N_16275,N_14410,N_12847);
nor U16276 (N_16276,N_14501,N_13971);
xor U16277 (N_16277,N_14187,N_14979);
nor U16278 (N_16278,N_13168,N_14039);
and U16279 (N_16279,N_12511,N_14051);
xor U16280 (N_16280,N_14575,N_14823);
nand U16281 (N_16281,N_12754,N_13646);
nand U16282 (N_16282,N_12961,N_14086);
nor U16283 (N_16283,N_14565,N_13295);
nor U16284 (N_16284,N_12907,N_13631);
nand U16285 (N_16285,N_13187,N_12579);
xor U16286 (N_16286,N_12587,N_14524);
nand U16287 (N_16287,N_13553,N_12892);
xor U16288 (N_16288,N_13513,N_13427);
xor U16289 (N_16289,N_12995,N_12895);
and U16290 (N_16290,N_13417,N_14323);
and U16291 (N_16291,N_14663,N_12643);
or U16292 (N_16292,N_13756,N_13150);
xnor U16293 (N_16293,N_12637,N_13573);
and U16294 (N_16294,N_12860,N_13177);
nor U16295 (N_16295,N_13719,N_14525);
nor U16296 (N_16296,N_13490,N_14971);
nand U16297 (N_16297,N_14637,N_13786);
nor U16298 (N_16298,N_14355,N_12592);
and U16299 (N_16299,N_12753,N_14074);
nand U16300 (N_16300,N_14251,N_13884);
xnor U16301 (N_16301,N_14595,N_12639);
nand U16302 (N_16302,N_13147,N_12902);
or U16303 (N_16303,N_13310,N_12847);
xnor U16304 (N_16304,N_13575,N_14904);
and U16305 (N_16305,N_13508,N_13937);
and U16306 (N_16306,N_12669,N_13566);
nor U16307 (N_16307,N_14669,N_14861);
or U16308 (N_16308,N_12877,N_13219);
xor U16309 (N_16309,N_13643,N_14538);
nor U16310 (N_16310,N_12536,N_12939);
nand U16311 (N_16311,N_14268,N_14839);
nand U16312 (N_16312,N_14307,N_12839);
nor U16313 (N_16313,N_13142,N_14777);
nor U16314 (N_16314,N_14649,N_14906);
or U16315 (N_16315,N_14560,N_14988);
nor U16316 (N_16316,N_13844,N_14465);
and U16317 (N_16317,N_14813,N_12772);
nand U16318 (N_16318,N_13038,N_14553);
and U16319 (N_16319,N_14433,N_14879);
nand U16320 (N_16320,N_14411,N_13101);
or U16321 (N_16321,N_12716,N_12985);
or U16322 (N_16322,N_14141,N_12924);
and U16323 (N_16323,N_14147,N_14897);
and U16324 (N_16324,N_14399,N_13713);
xnor U16325 (N_16325,N_13632,N_13951);
nor U16326 (N_16326,N_13001,N_14979);
xnor U16327 (N_16327,N_12770,N_13663);
and U16328 (N_16328,N_14236,N_13477);
nand U16329 (N_16329,N_12961,N_14133);
xor U16330 (N_16330,N_14057,N_14088);
xor U16331 (N_16331,N_14238,N_14320);
xor U16332 (N_16332,N_13989,N_12503);
or U16333 (N_16333,N_13666,N_14875);
and U16334 (N_16334,N_12812,N_14398);
and U16335 (N_16335,N_14679,N_13035);
and U16336 (N_16336,N_14297,N_14579);
or U16337 (N_16337,N_13888,N_12735);
xor U16338 (N_16338,N_12751,N_14773);
xor U16339 (N_16339,N_14127,N_13104);
xnor U16340 (N_16340,N_12733,N_13456);
or U16341 (N_16341,N_14918,N_14859);
nor U16342 (N_16342,N_12534,N_13829);
xnor U16343 (N_16343,N_14579,N_12839);
or U16344 (N_16344,N_13211,N_13335);
or U16345 (N_16345,N_13418,N_14497);
nor U16346 (N_16346,N_13175,N_14858);
and U16347 (N_16347,N_14366,N_12647);
nand U16348 (N_16348,N_13468,N_14560);
and U16349 (N_16349,N_13148,N_13952);
nand U16350 (N_16350,N_12773,N_14751);
or U16351 (N_16351,N_13564,N_13274);
nor U16352 (N_16352,N_14234,N_14747);
and U16353 (N_16353,N_14791,N_14625);
or U16354 (N_16354,N_14798,N_14532);
nand U16355 (N_16355,N_12611,N_13001);
or U16356 (N_16356,N_13899,N_12768);
nand U16357 (N_16357,N_14746,N_13791);
or U16358 (N_16358,N_13318,N_14885);
xor U16359 (N_16359,N_14481,N_12861);
nand U16360 (N_16360,N_13792,N_12827);
xnor U16361 (N_16361,N_14308,N_12908);
nand U16362 (N_16362,N_14535,N_14282);
xor U16363 (N_16363,N_13023,N_13218);
or U16364 (N_16364,N_14226,N_12818);
nor U16365 (N_16365,N_12741,N_13864);
nand U16366 (N_16366,N_12912,N_14783);
nor U16367 (N_16367,N_14477,N_14668);
nand U16368 (N_16368,N_13473,N_14966);
nand U16369 (N_16369,N_13107,N_14186);
and U16370 (N_16370,N_13892,N_13289);
xor U16371 (N_16371,N_14212,N_13466);
nor U16372 (N_16372,N_14335,N_13120);
nor U16373 (N_16373,N_12808,N_14520);
nand U16374 (N_16374,N_14299,N_14450);
and U16375 (N_16375,N_12568,N_14399);
xor U16376 (N_16376,N_13212,N_14021);
and U16377 (N_16377,N_12979,N_14697);
or U16378 (N_16378,N_13539,N_13807);
and U16379 (N_16379,N_13053,N_13183);
nand U16380 (N_16380,N_14622,N_14458);
and U16381 (N_16381,N_13613,N_14827);
and U16382 (N_16382,N_14216,N_14337);
or U16383 (N_16383,N_13394,N_14679);
nand U16384 (N_16384,N_13583,N_13731);
or U16385 (N_16385,N_14390,N_12558);
xnor U16386 (N_16386,N_14163,N_13951);
or U16387 (N_16387,N_13714,N_12942);
or U16388 (N_16388,N_14174,N_13607);
or U16389 (N_16389,N_14140,N_13297);
nor U16390 (N_16390,N_13443,N_13228);
or U16391 (N_16391,N_14690,N_12680);
xor U16392 (N_16392,N_12982,N_13516);
xnor U16393 (N_16393,N_13225,N_13338);
nor U16394 (N_16394,N_14437,N_12690);
and U16395 (N_16395,N_12804,N_14154);
and U16396 (N_16396,N_13483,N_12628);
nor U16397 (N_16397,N_13700,N_13225);
nor U16398 (N_16398,N_13286,N_13375);
nor U16399 (N_16399,N_12952,N_14783);
nor U16400 (N_16400,N_14026,N_13916);
xor U16401 (N_16401,N_14661,N_12734);
or U16402 (N_16402,N_12788,N_14651);
and U16403 (N_16403,N_12926,N_12932);
nand U16404 (N_16404,N_12853,N_13990);
or U16405 (N_16405,N_14137,N_14128);
xnor U16406 (N_16406,N_13597,N_13277);
and U16407 (N_16407,N_13897,N_14887);
and U16408 (N_16408,N_12639,N_12705);
and U16409 (N_16409,N_14040,N_14149);
or U16410 (N_16410,N_14752,N_12892);
nor U16411 (N_16411,N_14863,N_14987);
and U16412 (N_16412,N_12997,N_14791);
xnor U16413 (N_16413,N_13440,N_14931);
xor U16414 (N_16414,N_13788,N_14288);
and U16415 (N_16415,N_14594,N_12768);
xor U16416 (N_16416,N_13229,N_14062);
and U16417 (N_16417,N_14086,N_13945);
or U16418 (N_16418,N_12538,N_13542);
xnor U16419 (N_16419,N_14745,N_14770);
xnor U16420 (N_16420,N_14978,N_14835);
xnor U16421 (N_16421,N_13792,N_13585);
or U16422 (N_16422,N_12628,N_13548);
or U16423 (N_16423,N_13716,N_14205);
or U16424 (N_16424,N_14498,N_13366);
nor U16425 (N_16425,N_12713,N_13304);
and U16426 (N_16426,N_14742,N_13400);
nor U16427 (N_16427,N_13648,N_13176);
nor U16428 (N_16428,N_14140,N_13121);
nand U16429 (N_16429,N_14276,N_13401);
or U16430 (N_16430,N_14697,N_14831);
nor U16431 (N_16431,N_13762,N_14469);
and U16432 (N_16432,N_13394,N_12691);
nand U16433 (N_16433,N_12860,N_14054);
and U16434 (N_16434,N_14002,N_13038);
xor U16435 (N_16435,N_14978,N_13109);
nor U16436 (N_16436,N_12698,N_13858);
or U16437 (N_16437,N_12866,N_14755);
nand U16438 (N_16438,N_13842,N_14826);
or U16439 (N_16439,N_14110,N_12653);
nand U16440 (N_16440,N_14225,N_13845);
xor U16441 (N_16441,N_14314,N_12696);
nand U16442 (N_16442,N_14712,N_12752);
nor U16443 (N_16443,N_13781,N_14251);
or U16444 (N_16444,N_14408,N_12542);
and U16445 (N_16445,N_14187,N_13613);
and U16446 (N_16446,N_14471,N_14635);
xor U16447 (N_16447,N_14196,N_13649);
nand U16448 (N_16448,N_14834,N_12965);
nor U16449 (N_16449,N_14002,N_14048);
xnor U16450 (N_16450,N_13334,N_12594);
nand U16451 (N_16451,N_12527,N_12687);
xor U16452 (N_16452,N_13453,N_14594);
xnor U16453 (N_16453,N_12894,N_13712);
and U16454 (N_16454,N_12532,N_12515);
or U16455 (N_16455,N_14632,N_14443);
nor U16456 (N_16456,N_14605,N_14648);
and U16457 (N_16457,N_14306,N_13208);
nand U16458 (N_16458,N_13225,N_13801);
nand U16459 (N_16459,N_13357,N_14509);
xnor U16460 (N_16460,N_14967,N_12792);
xnor U16461 (N_16461,N_12873,N_13070);
xnor U16462 (N_16462,N_14491,N_13616);
or U16463 (N_16463,N_13266,N_14371);
nor U16464 (N_16464,N_14112,N_13707);
xnor U16465 (N_16465,N_13951,N_14969);
nor U16466 (N_16466,N_12879,N_14008);
or U16467 (N_16467,N_14693,N_14861);
nand U16468 (N_16468,N_14433,N_13343);
and U16469 (N_16469,N_13140,N_12799);
nand U16470 (N_16470,N_12539,N_14749);
nand U16471 (N_16471,N_12662,N_14120);
xnor U16472 (N_16472,N_13734,N_14698);
or U16473 (N_16473,N_14584,N_14849);
or U16474 (N_16474,N_13339,N_14243);
nor U16475 (N_16475,N_13372,N_13126);
and U16476 (N_16476,N_14252,N_13486);
and U16477 (N_16477,N_13736,N_14353);
nor U16478 (N_16478,N_13088,N_14284);
nor U16479 (N_16479,N_14230,N_13078);
nand U16480 (N_16480,N_13321,N_12756);
nand U16481 (N_16481,N_13983,N_13424);
nor U16482 (N_16482,N_14742,N_14419);
and U16483 (N_16483,N_14219,N_13042);
nor U16484 (N_16484,N_14639,N_14752);
nand U16485 (N_16485,N_14925,N_14860);
nand U16486 (N_16486,N_14344,N_14305);
nor U16487 (N_16487,N_14706,N_13194);
nand U16488 (N_16488,N_14301,N_12870);
xor U16489 (N_16489,N_12614,N_12670);
and U16490 (N_16490,N_14542,N_14259);
nor U16491 (N_16491,N_12801,N_13124);
or U16492 (N_16492,N_12894,N_14766);
nor U16493 (N_16493,N_13305,N_13964);
nor U16494 (N_16494,N_13064,N_13271);
nor U16495 (N_16495,N_13452,N_12628);
xnor U16496 (N_16496,N_13137,N_12813);
and U16497 (N_16497,N_13259,N_14196);
or U16498 (N_16498,N_12999,N_14136);
or U16499 (N_16499,N_14998,N_14288);
nor U16500 (N_16500,N_14837,N_12502);
nand U16501 (N_16501,N_14135,N_14844);
and U16502 (N_16502,N_14840,N_13760);
nor U16503 (N_16503,N_13669,N_13633);
or U16504 (N_16504,N_13174,N_14236);
or U16505 (N_16505,N_13825,N_12734);
nand U16506 (N_16506,N_14440,N_14997);
or U16507 (N_16507,N_13557,N_14894);
xor U16508 (N_16508,N_13093,N_12640);
nand U16509 (N_16509,N_14407,N_13898);
or U16510 (N_16510,N_14504,N_12783);
or U16511 (N_16511,N_14795,N_12874);
xor U16512 (N_16512,N_12608,N_14576);
and U16513 (N_16513,N_14018,N_13334);
xnor U16514 (N_16514,N_12509,N_12763);
nor U16515 (N_16515,N_12540,N_14314);
nor U16516 (N_16516,N_13074,N_12830);
or U16517 (N_16517,N_14610,N_13792);
xor U16518 (N_16518,N_12949,N_14630);
and U16519 (N_16519,N_14961,N_13903);
xor U16520 (N_16520,N_12628,N_13759);
nand U16521 (N_16521,N_13661,N_12530);
nor U16522 (N_16522,N_14069,N_13195);
or U16523 (N_16523,N_14441,N_14608);
nor U16524 (N_16524,N_13598,N_12987);
and U16525 (N_16525,N_13537,N_14316);
or U16526 (N_16526,N_14082,N_14351);
or U16527 (N_16527,N_14860,N_13563);
and U16528 (N_16528,N_12993,N_12674);
nand U16529 (N_16529,N_13482,N_13705);
or U16530 (N_16530,N_12814,N_14212);
xnor U16531 (N_16531,N_14591,N_14090);
or U16532 (N_16532,N_14525,N_14103);
and U16533 (N_16533,N_13169,N_12639);
nand U16534 (N_16534,N_13398,N_14006);
or U16535 (N_16535,N_14756,N_13544);
xnor U16536 (N_16536,N_14743,N_13923);
and U16537 (N_16537,N_13011,N_14063);
nand U16538 (N_16538,N_14714,N_12534);
and U16539 (N_16539,N_13901,N_13812);
nor U16540 (N_16540,N_14343,N_14998);
nor U16541 (N_16541,N_13123,N_14035);
xor U16542 (N_16542,N_14869,N_14529);
nor U16543 (N_16543,N_14097,N_14859);
nand U16544 (N_16544,N_14440,N_14057);
or U16545 (N_16545,N_14850,N_13426);
nor U16546 (N_16546,N_12622,N_14974);
nand U16547 (N_16547,N_13791,N_13982);
and U16548 (N_16548,N_12583,N_13245);
nor U16549 (N_16549,N_13232,N_13099);
nor U16550 (N_16550,N_13429,N_14411);
nand U16551 (N_16551,N_12782,N_14935);
xor U16552 (N_16552,N_12662,N_12605);
xnor U16553 (N_16553,N_14733,N_14703);
nand U16554 (N_16554,N_12805,N_13121);
nand U16555 (N_16555,N_14848,N_13374);
nor U16556 (N_16556,N_13672,N_14499);
xor U16557 (N_16557,N_14044,N_12598);
nand U16558 (N_16558,N_14112,N_12615);
and U16559 (N_16559,N_13603,N_13105);
or U16560 (N_16560,N_12506,N_12582);
nand U16561 (N_16561,N_14751,N_14340);
xor U16562 (N_16562,N_13319,N_14525);
and U16563 (N_16563,N_13329,N_12708);
or U16564 (N_16564,N_12563,N_13263);
and U16565 (N_16565,N_14689,N_14129);
or U16566 (N_16566,N_12850,N_14977);
or U16567 (N_16567,N_12854,N_13323);
nor U16568 (N_16568,N_14758,N_12744);
nor U16569 (N_16569,N_14822,N_12513);
and U16570 (N_16570,N_12837,N_14049);
and U16571 (N_16571,N_14456,N_13698);
nor U16572 (N_16572,N_14720,N_14167);
or U16573 (N_16573,N_12939,N_12671);
nor U16574 (N_16574,N_13747,N_13605);
or U16575 (N_16575,N_12634,N_12864);
xor U16576 (N_16576,N_14868,N_14554);
nand U16577 (N_16577,N_13506,N_14342);
xor U16578 (N_16578,N_13775,N_13910);
xor U16579 (N_16579,N_13259,N_13273);
and U16580 (N_16580,N_14259,N_14695);
nand U16581 (N_16581,N_12956,N_13233);
and U16582 (N_16582,N_14088,N_13918);
xor U16583 (N_16583,N_13626,N_13907);
or U16584 (N_16584,N_13004,N_14602);
xor U16585 (N_16585,N_14687,N_14062);
nor U16586 (N_16586,N_13221,N_12503);
nand U16587 (N_16587,N_14248,N_13849);
and U16588 (N_16588,N_13899,N_13479);
and U16589 (N_16589,N_13669,N_14081);
and U16590 (N_16590,N_12699,N_13769);
nor U16591 (N_16591,N_13983,N_13423);
nand U16592 (N_16592,N_14279,N_12780);
nand U16593 (N_16593,N_14926,N_14556);
xor U16594 (N_16594,N_14060,N_13190);
and U16595 (N_16595,N_12830,N_13239);
and U16596 (N_16596,N_12536,N_14396);
or U16597 (N_16597,N_14801,N_13991);
nor U16598 (N_16598,N_14334,N_12812);
or U16599 (N_16599,N_12952,N_13201);
nand U16600 (N_16600,N_13605,N_12886);
and U16601 (N_16601,N_13540,N_13440);
nand U16602 (N_16602,N_14469,N_12645);
nand U16603 (N_16603,N_12886,N_12770);
and U16604 (N_16604,N_13335,N_14904);
xor U16605 (N_16605,N_14088,N_14315);
or U16606 (N_16606,N_13634,N_13501);
and U16607 (N_16607,N_12529,N_13021);
and U16608 (N_16608,N_13143,N_12669);
nor U16609 (N_16609,N_12771,N_13713);
nor U16610 (N_16610,N_13713,N_14798);
nand U16611 (N_16611,N_13623,N_12652);
or U16612 (N_16612,N_12893,N_13527);
or U16613 (N_16613,N_14173,N_12700);
and U16614 (N_16614,N_12771,N_14654);
xnor U16615 (N_16615,N_13794,N_13622);
and U16616 (N_16616,N_13996,N_12786);
and U16617 (N_16617,N_14645,N_14010);
or U16618 (N_16618,N_12844,N_14905);
or U16619 (N_16619,N_14294,N_14325);
nand U16620 (N_16620,N_13457,N_14797);
nand U16621 (N_16621,N_14254,N_13883);
nor U16622 (N_16622,N_14383,N_13252);
nand U16623 (N_16623,N_13252,N_14361);
xnor U16624 (N_16624,N_12587,N_13947);
nor U16625 (N_16625,N_14060,N_14380);
or U16626 (N_16626,N_12844,N_13179);
or U16627 (N_16627,N_13692,N_12953);
and U16628 (N_16628,N_13924,N_14064);
nor U16629 (N_16629,N_12882,N_12876);
xor U16630 (N_16630,N_13532,N_14897);
or U16631 (N_16631,N_14795,N_13258);
xnor U16632 (N_16632,N_14734,N_13683);
nand U16633 (N_16633,N_13578,N_12715);
xor U16634 (N_16634,N_14576,N_14402);
or U16635 (N_16635,N_14832,N_12695);
nand U16636 (N_16636,N_14734,N_12657);
and U16637 (N_16637,N_13027,N_14011);
nand U16638 (N_16638,N_14263,N_12979);
nand U16639 (N_16639,N_13520,N_13387);
and U16640 (N_16640,N_14072,N_14337);
nand U16641 (N_16641,N_14108,N_12889);
nand U16642 (N_16642,N_12514,N_13833);
nor U16643 (N_16643,N_12910,N_13151);
nor U16644 (N_16644,N_13401,N_14887);
or U16645 (N_16645,N_14655,N_14647);
nand U16646 (N_16646,N_12592,N_13832);
or U16647 (N_16647,N_12849,N_13940);
or U16648 (N_16648,N_13587,N_14636);
or U16649 (N_16649,N_13641,N_14895);
or U16650 (N_16650,N_13898,N_14142);
xnor U16651 (N_16651,N_14712,N_14315);
nor U16652 (N_16652,N_14596,N_12749);
and U16653 (N_16653,N_14968,N_13253);
nand U16654 (N_16654,N_14218,N_14142);
xnor U16655 (N_16655,N_13805,N_12642);
or U16656 (N_16656,N_13477,N_13376);
xor U16657 (N_16657,N_12926,N_13213);
nor U16658 (N_16658,N_13197,N_12722);
and U16659 (N_16659,N_14646,N_13880);
nor U16660 (N_16660,N_12935,N_13469);
xor U16661 (N_16661,N_13124,N_12993);
or U16662 (N_16662,N_13279,N_13158);
nor U16663 (N_16663,N_13810,N_13317);
nand U16664 (N_16664,N_14864,N_14147);
nor U16665 (N_16665,N_14535,N_13366);
or U16666 (N_16666,N_14589,N_14785);
nand U16667 (N_16667,N_14447,N_13201);
nand U16668 (N_16668,N_14659,N_14483);
xor U16669 (N_16669,N_13352,N_14505);
and U16670 (N_16670,N_14224,N_12881);
nand U16671 (N_16671,N_14463,N_13942);
xor U16672 (N_16672,N_14066,N_13919);
nor U16673 (N_16673,N_14522,N_13802);
nor U16674 (N_16674,N_13798,N_13511);
xnor U16675 (N_16675,N_13591,N_13459);
nand U16676 (N_16676,N_12921,N_14139);
nor U16677 (N_16677,N_13501,N_13358);
xor U16678 (N_16678,N_14098,N_14629);
xnor U16679 (N_16679,N_13072,N_12751);
or U16680 (N_16680,N_13467,N_13273);
nor U16681 (N_16681,N_13489,N_14824);
and U16682 (N_16682,N_14054,N_13372);
nand U16683 (N_16683,N_13499,N_13501);
and U16684 (N_16684,N_12636,N_14110);
and U16685 (N_16685,N_13438,N_14783);
or U16686 (N_16686,N_14165,N_13201);
and U16687 (N_16687,N_12565,N_13134);
nand U16688 (N_16688,N_14035,N_14923);
xor U16689 (N_16689,N_13707,N_12996);
nor U16690 (N_16690,N_13065,N_14685);
nor U16691 (N_16691,N_12718,N_14325);
nor U16692 (N_16692,N_14585,N_13427);
nand U16693 (N_16693,N_14195,N_13241);
nor U16694 (N_16694,N_14647,N_14125);
xnor U16695 (N_16695,N_14145,N_12967);
nand U16696 (N_16696,N_14007,N_14338);
or U16697 (N_16697,N_12580,N_13799);
xor U16698 (N_16698,N_14989,N_14205);
nor U16699 (N_16699,N_14955,N_14917);
nor U16700 (N_16700,N_14528,N_12572);
xnor U16701 (N_16701,N_12686,N_12697);
or U16702 (N_16702,N_13351,N_13997);
nor U16703 (N_16703,N_12704,N_13248);
or U16704 (N_16704,N_12535,N_13840);
and U16705 (N_16705,N_12941,N_12812);
nand U16706 (N_16706,N_14008,N_12554);
and U16707 (N_16707,N_14762,N_13565);
xor U16708 (N_16708,N_12725,N_13412);
nand U16709 (N_16709,N_14892,N_13146);
nand U16710 (N_16710,N_14985,N_13069);
nand U16711 (N_16711,N_14045,N_12697);
or U16712 (N_16712,N_14959,N_13314);
nand U16713 (N_16713,N_14434,N_13732);
xor U16714 (N_16714,N_14587,N_14105);
nand U16715 (N_16715,N_12824,N_14036);
or U16716 (N_16716,N_13642,N_12527);
nor U16717 (N_16717,N_13476,N_14599);
xnor U16718 (N_16718,N_14388,N_14819);
xnor U16719 (N_16719,N_13960,N_13365);
nor U16720 (N_16720,N_13927,N_14748);
nor U16721 (N_16721,N_13149,N_13990);
nand U16722 (N_16722,N_12570,N_13171);
nor U16723 (N_16723,N_12777,N_13580);
and U16724 (N_16724,N_13805,N_13871);
or U16725 (N_16725,N_14744,N_14027);
and U16726 (N_16726,N_13111,N_12933);
xor U16727 (N_16727,N_13337,N_14256);
and U16728 (N_16728,N_13257,N_14265);
or U16729 (N_16729,N_12913,N_14861);
nand U16730 (N_16730,N_14737,N_14844);
and U16731 (N_16731,N_14825,N_14832);
nor U16732 (N_16732,N_12608,N_14204);
nor U16733 (N_16733,N_12887,N_14724);
nand U16734 (N_16734,N_13808,N_13195);
xor U16735 (N_16735,N_14479,N_14006);
or U16736 (N_16736,N_14202,N_13118);
nor U16737 (N_16737,N_12689,N_14655);
nand U16738 (N_16738,N_14208,N_14089);
and U16739 (N_16739,N_14151,N_14481);
nor U16740 (N_16740,N_14395,N_12709);
or U16741 (N_16741,N_12951,N_13765);
and U16742 (N_16742,N_14645,N_13537);
and U16743 (N_16743,N_12696,N_12934);
or U16744 (N_16744,N_12993,N_13163);
nor U16745 (N_16745,N_13861,N_14063);
or U16746 (N_16746,N_14080,N_14448);
and U16747 (N_16747,N_14064,N_14870);
nor U16748 (N_16748,N_13929,N_14027);
xor U16749 (N_16749,N_12929,N_14369);
nor U16750 (N_16750,N_13829,N_13728);
and U16751 (N_16751,N_14369,N_13272);
xor U16752 (N_16752,N_13992,N_13878);
or U16753 (N_16753,N_14430,N_14877);
nand U16754 (N_16754,N_14152,N_13650);
nor U16755 (N_16755,N_12926,N_14464);
or U16756 (N_16756,N_14602,N_13135);
nand U16757 (N_16757,N_13466,N_13506);
nand U16758 (N_16758,N_12667,N_14341);
xnor U16759 (N_16759,N_13888,N_12628);
nor U16760 (N_16760,N_14191,N_14606);
and U16761 (N_16761,N_14647,N_13958);
xnor U16762 (N_16762,N_12722,N_14031);
nand U16763 (N_16763,N_13194,N_14788);
and U16764 (N_16764,N_13671,N_14886);
or U16765 (N_16765,N_13847,N_14466);
xnor U16766 (N_16766,N_12798,N_13923);
and U16767 (N_16767,N_12983,N_12700);
nor U16768 (N_16768,N_13420,N_13995);
and U16769 (N_16769,N_14310,N_14428);
nor U16770 (N_16770,N_13711,N_13301);
or U16771 (N_16771,N_13718,N_12911);
xor U16772 (N_16772,N_13510,N_14939);
nand U16773 (N_16773,N_13930,N_14306);
and U16774 (N_16774,N_13687,N_13274);
or U16775 (N_16775,N_14537,N_12530);
or U16776 (N_16776,N_14346,N_14619);
nor U16777 (N_16777,N_14048,N_12849);
nand U16778 (N_16778,N_13907,N_13901);
nand U16779 (N_16779,N_13750,N_13109);
or U16780 (N_16780,N_13953,N_14509);
or U16781 (N_16781,N_13948,N_14852);
or U16782 (N_16782,N_14132,N_13655);
and U16783 (N_16783,N_14849,N_14210);
nand U16784 (N_16784,N_13617,N_13776);
nand U16785 (N_16785,N_14257,N_12896);
or U16786 (N_16786,N_14181,N_14561);
xor U16787 (N_16787,N_14629,N_12941);
nor U16788 (N_16788,N_13782,N_13747);
or U16789 (N_16789,N_13384,N_13171);
nand U16790 (N_16790,N_12559,N_14256);
xor U16791 (N_16791,N_14863,N_12578);
xnor U16792 (N_16792,N_14501,N_13837);
nor U16793 (N_16793,N_14460,N_14094);
nor U16794 (N_16794,N_13430,N_13955);
nand U16795 (N_16795,N_14392,N_13982);
xor U16796 (N_16796,N_14086,N_12816);
nand U16797 (N_16797,N_14620,N_13234);
nor U16798 (N_16798,N_13402,N_14441);
nand U16799 (N_16799,N_13576,N_14548);
and U16800 (N_16800,N_14843,N_14547);
nor U16801 (N_16801,N_12888,N_12717);
nand U16802 (N_16802,N_13243,N_12573);
xor U16803 (N_16803,N_13979,N_13756);
nor U16804 (N_16804,N_13493,N_14043);
xor U16805 (N_16805,N_13765,N_14693);
and U16806 (N_16806,N_12739,N_14027);
or U16807 (N_16807,N_13056,N_13595);
nor U16808 (N_16808,N_13189,N_12800);
or U16809 (N_16809,N_14396,N_13723);
nor U16810 (N_16810,N_14865,N_14882);
or U16811 (N_16811,N_12981,N_13530);
nand U16812 (N_16812,N_14497,N_12549);
and U16813 (N_16813,N_13107,N_13510);
nor U16814 (N_16814,N_14773,N_12952);
xnor U16815 (N_16815,N_13014,N_14549);
xor U16816 (N_16816,N_14245,N_14789);
xnor U16817 (N_16817,N_13481,N_14583);
and U16818 (N_16818,N_14141,N_14467);
or U16819 (N_16819,N_13998,N_13033);
or U16820 (N_16820,N_14201,N_14263);
and U16821 (N_16821,N_14988,N_14672);
xor U16822 (N_16822,N_13527,N_14278);
nand U16823 (N_16823,N_13242,N_12660);
xor U16824 (N_16824,N_14255,N_13281);
xnor U16825 (N_16825,N_13118,N_14055);
nand U16826 (N_16826,N_12670,N_12787);
xnor U16827 (N_16827,N_14602,N_12571);
nand U16828 (N_16828,N_12808,N_13591);
or U16829 (N_16829,N_13270,N_13613);
nor U16830 (N_16830,N_14792,N_14694);
nor U16831 (N_16831,N_13466,N_13416);
xnor U16832 (N_16832,N_13134,N_13508);
and U16833 (N_16833,N_14997,N_13241);
nand U16834 (N_16834,N_12849,N_14075);
nand U16835 (N_16835,N_14309,N_14723);
or U16836 (N_16836,N_12978,N_13567);
nor U16837 (N_16837,N_14408,N_13111);
xor U16838 (N_16838,N_13324,N_14609);
or U16839 (N_16839,N_13415,N_13316);
and U16840 (N_16840,N_12600,N_14107);
nor U16841 (N_16841,N_12747,N_13277);
or U16842 (N_16842,N_13866,N_14609);
and U16843 (N_16843,N_13219,N_13844);
nand U16844 (N_16844,N_14774,N_13058);
nand U16845 (N_16845,N_12703,N_13113);
and U16846 (N_16846,N_13137,N_12574);
and U16847 (N_16847,N_14037,N_14391);
or U16848 (N_16848,N_13440,N_13284);
nand U16849 (N_16849,N_12512,N_14579);
or U16850 (N_16850,N_14843,N_14404);
or U16851 (N_16851,N_13210,N_14568);
nand U16852 (N_16852,N_13622,N_13493);
nor U16853 (N_16853,N_14503,N_14765);
and U16854 (N_16854,N_14082,N_13366);
nor U16855 (N_16855,N_14869,N_12945);
nand U16856 (N_16856,N_13287,N_13692);
nand U16857 (N_16857,N_13193,N_13623);
nand U16858 (N_16858,N_14212,N_13397);
and U16859 (N_16859,N_13784,N_14329);
or U16860 (N_16860,N_13374,N_14517);
or U16861 (N_16861,N_14039,N_14596);
nor U16862 (N_16862,N_14518,N_13327);
or U16863 (N_16863,N_13955,N_12749);
or U16864 (N_16864,N_13908,N_13096);
nor U16865 (N_16865,N_14321,N_13142);
nor U16866 (N_16866,N_13354,N_14866);
nand U16867 (N_16867,N_13116,N_13844);
or U16868 (N_16868,N_13966,N_14759);
nand U16869 (N_16869,N_13964,N_13722);
xnor U16870 (N_16870,N_14151,N_13265);
or U16871 (N_16871,N_13835,N_14892);
nor U16872 (N_16872,N_14119,N_12893);
nand U16873 (N_16873,N_13036,N_14090);
nand U16874 (N_16874,N_14785,N_13445);
nor U16875 (N_16875,N_13495,N_14927);
nor U16876 (N_16876,N_12860,N_12722);
nor U16877 (N_16877,N_14827,N_13403);
nor U16878 (N_16878,N_12676,N_14795);
nand U16879 (N_16879,N_14034,N_13517);
and U16880 (N_16880,N_13929,N_12650);
xor U16881 (N_16881,N_14416,N_14402);
xnor U16882 (N_16882,N_13273,N_12849);
nand U16883 (N_16883,N_14501,N_13545);
nor U16884 (N_16884,N_12852,N_13838);
or U16885 (N_16885,N_12667,N_14794);
nand U16886 (N_16886,N_13482,N_14035);
and U16887 (N_16887,N_13301,N_12528);
or U16888 (N_16888,N_13708,N_13780);
and U16889 (N_16889,N_13914,N_12814);
or U16890 (N_16890,N_14013,N_14237);
or U16891 (N_16891,N_12778,N_14755);
nor U16892 (N_16892,N_13822,N_13729);
nand U16893 (N_16893,N_13366,N_13820);
xnor U16894 (N_16894,N_12575,N_14579);
or U16895 (N_16895,N_14547,N_13949);
nand U16896 (N_16896,N_13707,N_14043);
or U16897 (N_16897,N_13081,N_13126);
nand U16898 (N_16898,N_12896,N_14716);
nor U16899 (N_16899,N_13531,N_13745);
xnor U16900 (N_16900,N_14036,N_13393);
nand U16901 (N_16901,N_14862,N_13591);
nand U16902 (N_16902,N_12832,N_13316);
or U16903 (N_16903,N_12930,N_14665);
and U16904 (N_16904,N_14636,N_13151);
and U16905 (N_16905,N_14870,N_13197);
nor U16906 (N_16906,N_14027,N_13285);
nor U16907 (N_16907,N_14670,N_12938);
xor U16908 (N_16908,N_14308,N_13866);
or U16909 (N_16909,N_14475,N_13984);
nand U16910 (N_16910,N_12731,N_12826);
nand U16911 (N_16911,N_14355,N_14269);
and U16912 (N_16912,N_13528,N_13788);
xnor U16913 (N_16913,N_12873,N_13411);
nor U16914 (N_16914,N_12776,N_13866);
or U16915 (N_16915,N_14867,N_13123);
nand U16916 (N_16916,N_13326,N_14370);
or U16917 (N_16917,N_14526,N_13832);
nand U16918 (N_16918,N_14378,N_12741);
nor U16919 (N_16919,N_14712,N_13689);
nand U16920 (N_16920,N_13425,N_14185);
nor U16921 (N_16921,N_13886,N_13492);
and U16922 (N_16922,N_13242,N_14166);
xor U16923 (N_16923,N_13136,N_13377);
and U16924 (N_16924,N_13331,N_13522);
xnor U16925 (N_16925,N_14503,N_13196);
and U16926 (N_16926,N_13255,N_14590);
and U16927 (N_16927,N_12697,N_14704);
nand U16928 (N_16928,N_12924,N_14166);
xor U16929 (N_16929,N_12503,N_14059);
nor U16930 (N_16930,N_14800,N_12970);
nor U16931 (N_16931,N_12556,N_14596);
nand U16932 (N_16932,N_12840,N_12696);
xnor U16933 (N_16933,N_12977,N_14089);
xor U16934 (N_16934,N_14613,N_14684);
and U16935 (N_16935,N_13893,N_13107);
and U16936 (N_16936,N_13074,N_12960);
or U16937 (N_16937,N_14324,N_13774);
or U16938 (N_16938,N_13697,N_13000);
nand U16939 (N_16939,N_12766,N_12579);
nand U16940 (N_16940,N_12523,N_13019);
nand U16941 (N_16941,N_14526,N_13694);
or U16942 (N_16942,N_12541,N_13430);
and U16943 (N_16943,N_13380,N_14248);
or U16944 (N_16944,N_13181,N_14787);
or U16945 (N_16945,N_14799,N_14183);
xnor U16946 (N_16946,N_13301,N_14780);
and U16947 (N_16947,N_13325,N_13487);
nor U16948 (N_16948,N_13386,N_13837);
and U16949 (N_16949,N_14587,N_14487);
xor U16950 (N_16950,N_14317,N_13749);
nand U16951 (N_16951,N_14110,N_14340);
and U16952 (N_16952,N_13057,N_12829);
nand U16953 (N_16953,N_12816,N_13089);
xnor U16954 (N_16954,N_14534,N_14378);
and U16955 (N_16955,N_14296,N_14026);
nand U16956 (N_16956,N_12689,N_13745);
xnor U16957 (N_16957,N_13244,N_13652);
xor U16958 (N_16958,N_14249,N_13645);
nand U16959 (N_16959,N_14435,N_14218);
xor U16960 (N_16960,N_14687,N_14403);
xor U16961 (N_16961,N_14606,N_14046);
xor U16962 (N_16962,N_12695,N_13413);
or U16963 (N_16963,N_13931,N_13677);
nor U16964 (N_16964,N_13666,N_14849);
nand U16965 (N_16965,N_13100,N_12775);
and U16966 (N_16966,N_13603,N_14245);
xor U16967 (N_16967,N_13300,N_14410);
and U16968 (N_16968,N_12780,N_14897);
or U16969 (N_16969,N_14771,N_13847);
and U16970 (N_16970,N_13946,N_13414);
or U16971 (N_16971,N_13578,N_12844);
and U16972 (N_16972,N_14289,N_14962);
xor U16973 (N_16973,N_13527,N_12653);
and U16974 (N_16974,N_14936,N_12746);
and U16975 (N_16975,N_13059,N_14094);
nor U16976 (N_16976,N_14078,N_13799);
or U16977 (N_16977,N_14273,N_14225);
xor U16978 (N_16978,N_13711,N_14103);
nor U16979 (N_16979,N_14070,N_14513);
xnor U16980 (N_16980,N_12811,N_14817);
or U16981 (N_16981,N_14327,N_13386);
nor U16982 (N_16982,N_13051,N_13297);
xnor U16983 (N_16983,N_14437,N_14369);
or U16984 (N_16984,N_13339,N_13073);
and U16985 (N_16985,N_14845,N_12916);
xnor U16986 (N_16986,N_14569,N_14673);
or U16987 (N_16987,N_12556,N_14726);
nand U16988 (N_16988,N_13534,N_14684);
xnor U16989 (N_16989,N_14962,N_13541);
nor U16990 (N_16990,N_13130,N_13068);
nor U16991 (N_16991,N_13729,N_14679);
xor U16992 (N_16992,N_13606,N_13183);
nand U16993 (N_16993,N_13443,N_14908);
or U16994 (N_16994,N_13682,N_13422);
and U16995 (N_16995,N_13629,N_13464);
nand U16996 (N_16996,N_14600,N_13326);
and U16997 (N_16997,N_14122,N_14778);
and U16998 (N_16998,N_12864,N_12899);
nor U16999 (N_16999,N_13296,N_12749);
or U17000 (N_17000,N_14054,N_13847);
nand U17001 (N_17001,N_14903,N_12735);
nor U17002 (N_17002,N_14275,N_13971);
xor U17003 (N_17003,N_13743,N_13562);
and U17004 (N_17004,N_14016,N_12813);
and U17005 (N_17005,N_14552,N_13451);
nand U17006 (N_17006,N_13949,N_13202);
nor U17007 (N_17007,N_13737,N_13636);
and U17008 (N_17008,N_13360,N_14045);
and U17009 (N_17009,N_14013,N_13510);
or U17010 (N_17010,N_14963,N_14726);
nor U17011 (N_17011,N_13379,N_12859);
and U17012 (N_17012,N_12504,N_14311);
or U17013 (N_17013,N_14966,N_14063);
or U17014 (N_17014,N_13788,N_12572);
and U17015 (N_17015,N_14123,N_12984);
nand U17016 (N_17016,N_12565,N_13692);
nand U17017 (N_17017,N_13293,N_12528);
nand U17018 (N_17018,N_13312,N_12529);
and U17019 (N_17019,N_14763,N_13674);
and U17020 (N_17020,N_13033,N_13494);
or U17021 (N_17021,N_14387,N_14496);
and U17022 (N_17022,N_12579,N_13264);
nor U17023 (N_17023,N_13950,N_13136);
and U17024 (N_17024,N_14522,N_14400);
nand U17025 (N_17025,N_13005,N_14357);
nor U17026 (N_17026,N_14341,N_13737);
nand U17027 (N_17027,N_14848,N_14044);
nand U17028 (N_17028,N_13484,N_12950);
nand U17029 (N_17029,N_14826,N_13439);
nor U17030 (N_17030,N_12625,N_13532);
xor U17031 (N_17031,N_14124,N_12586);
and U17032 (N_17032,N_14157,N_13673);
xnor U17033 (N_17033,N_14976,N_14305);
nand U17034 (N_17034,N_12949,N_12899);
nor U17035 (N_17035,N_14566,N_14759);
nand U17036 (N_17036,N_12549,N_13002);
nor U17037 (N_17037,N_12849,N_12732);
xnor U17038 (N_17038,N_13629,N_13864);
nor U17039 (N_17039,N_13368,N_13268);
nand U17040 (N_17040,N_13853,N_13449);
or U17041 (N_17041,N_12510,N_14739);
or U17042 (N_17042,N_14831,N_13704);
or U17043 (N_17043,N_13598,N_12722);
nor U17044 (N_17044,N_14640,N_13964);
or U17045 (N_17045,N_13510,N_14827);
nor U17046 (N_17046,N_13761,N_13212);
and U17047 (N_17047,N_12771,N_14341);
nor U17048 (N_17048,N_12694,N_12704);
and U17049 (N_17049,N_13647,N_14897);
and U17050 (N_17050,N_13201,N_14309);
xor U17051 (N_17051,N_13666,N_13386);
or U17052 (N_17052,N_13900,N_13624);
nand U17053 (N_17053,N_14664,N_12680);
nor U17054 (N_17054,N_13269,N_13107);
xor U17055 (N_17055,N_14353,N_12958);
xnor U17056 (N_17056,N_13514,N_14572);
nor U17057 (N_17057,N_13546,N_12980);
and U17058 (N_17058,N_12970,N_13585);
nand U17059 (N_17059,N_13503,N_13469);
nor U17060 (N_17060,N_14646,N_14181);
nand U17061 (N_17061,N_14298,N_12562);
nand U17062 (N_17062,N_14975,N_14213);
and U17063 (N_17063,N_12747,N_13458);
xnor U17064 (N_17064,N_13082,N_13216);
and U17065 (N_17065,N_13827,N_13633);
nor U17066 (N_17066,N_12688,N_12676);
xor U17067 (N_17067,N_13971,N_13845);
xnor U17068 (N_17068,N_14465,N_14472);
nand U17069 (N_17069,N_14853,N_13577);
xnor U17070 (N_17070,N_14529,N_13486);
nand U17071 (N_17071,N_14702,N_14742);
and U17072 (N_17072,N_14951,N_13973);
and U17073 (N_17073,N_12848,N_12786);
or U17074 (N_17074,N_13013,N_13121);
nor U17075 (N_17075,N_14701,N_13299);
and U17076 (N_17076,N_14755,N_13349);
and U17077 (N_17077,N_13179,N_12662);
xnor U17078 (N_17078,N_13460,N_13701);
xor U17079 (N_17079,N_14621,N_14506);
nor U17080 (N_17080,N_12504,N_13890);
or U17081 (N_17081,N_14217,N_12808);
xor U17082 (N_17082,N_14593,N_13724);
or U17083 (N_17083,N_12572,N_13355);
and U17084 (N_17084,N_13415,N_13629);
or U17085 (N_17085,N_13563,N_13900);
xnor U17086 (N_17086,N_13763,N_13490);
xor U17087 (N_17087,N_13882,N_13793);
nor U17088 (N_17088,N_14828,N_12658);
nor U17089 (N_17089,N_14076,N_13574);
or U17090 (N_17090,N_14730,N_14495);
nor U17091 (N_17091,N_14659,N_13592);
nor U17092 (N_17092,N_14588,N_12953);
nor U17093 (N_17093,N_14916,N_13951);
nor U17094 (N_17094,N_14784,N_12765);
nand U17095 (N_17095,N_12930,N_14738);
or U17096 (N_17096,N_13355,N_12995);
nor U17097 (N_17097,N_12644,N_14495);
and U17098 (N_17098,N_12799,N_14218);
and U17099 (N_17099,N_14277,N_14110);
nand U17100 (N_17100,N_14538,N_14063);
and U17101 (N_17101,N_13826,N_14862);
xor U17102 (N_17102,N_14532,N_12702);
and U17103 (N_17103,N_14404,N_13199);
xor U17104 (N_17104,N_14866,N_13007);
nand U17105 (N_17105,N_13752,N_14642);
xor U17106 (N_17106,N_14547,N_13910);
nor U17107 (N_17107,N_14778,N_13875);
and U17108 (N_17108,N_13664,N_14324);
nand U17109 (N_17109,N_13195,N_14970);
or U17110 (N_17110,N_14760,N_14722);
and U17111 (N_17111,N_13997,N_14645);
and U17112 (N_17112,N_13376,N_12624);
nand U17113 (N_17113,N_12993,N_14676);
nor U17114 (N_17114,N_12906,N_12661);
nor U17115 (N_17115,N_13596,N_14156);
xnor U17116 (N_17116,N_13072,N_13597);
and U17117 (N_17117,N_13720,N_14657);
xor U17118 (N_17118,N_14756,N_14462);
xor U17119 (N_17119,N_14044,N_13276);
nor U17120 (N_17120,N_12803,N_13941);
nor U17121 (N_17121,N_12689,N_14906);
or U17122 (N_17122,N_14888,N_14567);
or U17123 (N_17123,N_14440,N_13840);
and U17124 (N_17124,N_12741,N_14618);
nor U17125 (N_17125,N_12990,N_13588);
xor U17126 (N_17126,N_13526,N_12663);
and U17127 (N_17127,N_13264,N_12938);
nand U17128 (N_17128,N_12640,N_12538);
nor U17129 (N_17129,N_13767,N_13821);
nor U17130 (N_17130,N_14464,N_14565);
xnor U17131 (N_17131,N_14644,N_14171);
nand U17132 (N_17132,N_12678,N_13375);
nand U17133 (N_17133,N_12552,N_14744);
xnor U17134 (N_17134,N_14378,N_12788);
or U17135 (N_17135,N_13240,N_13642);
or U17136 (N_17136,N_14617,N_13132);
xor U17137 (N_17137,N_14097,N_14439);
xnor U17138 (N_17138,N_12738,N_13727);
nand U17139 (N_17139,N_12506,N_13718);
or U17140 (N_17140,N_14119,N_14546);
or U17141 (N_17141,N_13323,N_12984);
or U17142 (N_17142,N_12776,N_14443);
and U17143 (N_17143,N_14231,N_14128);
nor U17144 (N_17144,N_14021,N_13304);
nand U17145 (N_17145,N_14647,N_14861);
xnor U17146 (N_17146,N_13612,N_13062);
xor U17147 (N_17147,N_13906,N_14655);
nor U17148 (N_17148,N_12821,N_13928);
nor U17149 (N_17149,N_14764,N_13487);
or U17150 (N_17150,N_12502,N_13204);
and U17151 (N_17151,N_12614,N_14645);
and U17152 (N_17152,N_12705,N_12527);
or U17153 (N_17153,N_12543,N_13527);
nor U17154 (N_17154,N_14717,N_12807);
xor U17155 (N_17155,N_14328,N_13166);
xor U17156 (N_17156,N_14460,N_14262);
xnor U17157 (N_17157,N_13097,N_14600);
nand U17158 (N_17158,N_13392,N_12742);
and U17159 (N_17159,N_14692,N_14849);
nor U17160 (N_17160,N_14167,N_12999);
and U17161 (N_17161,N_13900,N_12741);
and U17162 (N_17162,N_13669,N_12621);
nand U17163 (N_17163,N_14585,N_12808);
nor U17164 (N_17164,N_13995,N_14580);
nor U17165 (N_17165,N_12988,N_14342);
xnor U17166 (N_17166,N_14328,N_14439);
or U17167 (N_17167,N_13484,N_13878);
nor U17168 (N_17168,N_14102,N_14478);
xnor U17169 (N_17169,N_14231,N_12714);
nand U17170 (N_17170,N_14010,N_14793);
nor U17171 (N_17171,N_13018,N_13354);
or U17172 (N_17172,N_14149,N_13275);
or U17173 (N_17173,N_14264,N_14655);
xnor U17174 (N_17174,N_12527,N_12896);
nand U17175 (N_17175,N_14490,N_13109);
xnor U17176 (N_17176,N_13674,N_12877);
nand U17177 (N_17177,N_13624,N_14649);
nor U17178 (N_17178,N_12789,N_13344);
xor U17179 (N_17179,N_14736,N_14434);
and U17180 (N_17180,N_12988,N_14529);
or U17181 (N_17181,N_12668,N_14696);
nor U17182 (N_17182,N_14247,N_14898);
nand U17183 (N_17183,N_13529,N_13437);
nand U17184 (N_17184,N_13616,N_13513);
nand U17185 (N_17185,N_13424,N_13639);
xor U17186 (N_17186,N_14470,N_13359);
and U17187 (N_17187,N_14215,N_12793);
nand U17188 (N_17188,N_14458,N_14736);
xnor U17189 (N_17189,N_13837,N_13333);
or U17190 (N_17190,N_13963,N_13888);
and U17191 (N_17191,N_14530,N_14954);
and U17192 (N_17192,N_14737,N_14772);
xor U17193 (N_17193,N_14468,N_13091);
nor U17194 (N_17194,N_14356,N_14345);
nand U17195 (N_17195,N_13153,N_13498);
or U17196 (N_17196,N_14520,N_13060);
and U17197 (N_17197,N_13366,N_12869);
nand U17198 (N_17198,N_14106,N_14184);
nand U17199 (N_17199,N_14040,N_12960);
or U17200 (N_17200,N_14666,N_13367);
xor U17201 (N_17201,N_14793,N_13054);
xnor U17202 (N_17202,N_13885,N_13866);
nand U17203 (N_17203,N_12957,N_12784);
nand U17204 (N_17204,N_13039,N_13666);
nand U17205 (N_17205,N_13718,N_13728);
nor U17206 (N_17206,N_13161,N_14198);
xor U17207 (N_17207,N_14912,N_14930);
and U17208 (N_17208,N_12832,N_14955);
or U17209 (N_17209,N_12544,N_14368);
nor U17210 (N_17210,N_14727,N_12572);
nor U17211 (N_17211,N_12527,N_12977);
and U17212 (N_17212,N_13074,N_13383);
xnor U17213 (N_17213,N_13487,N_13013);
nor U17214 (N_17214,N_14396,N_13051);
and U17215 (N_17215,N_14750,N_14163);
and U17216 (N_17216,N_13811,N_12937);
or U17217 (N_17217,N_12759,N_12608);
or U17218 (N_17218,N_13491,N_12854);
nand U17219 (N_17219,N_12831,N_13628);
nor U17220 (N_17220,N_14992,N_13998);
nand U17221 (N_17221,N_13330,N_12804);
and U17222 (N_17222,N_14205,N_14325);
nor U17223 (N_17223,N_14119,N_12678);
nor U17224 (N_17224,N_14487,N_14827);
xor U17225 (N_17225,N_13640,N_12524);
nor U17226 (N_17226,N_13311,N_14692);
or U17227 (N_17227,N_14862,N_13447);
or U17228 (N_17228,N_14786,N_13106);
nor U17229 (N_17229,N_14771,N_13394);
nor U17230 (N_17230,N_13948,N_13182);
xor U17231 (N_17231,N_13786,N_13401);
xnor U17232 (N_17232,N_14468,N_14402);
or U17233 (N_17233,N_13538,N_13980);
nor U17234 (N_17234,N_13367,N_14520);
or U17235 (N_17235,N_13475,N_13730);
or U17236 (N_17236,N_12701,N_14642);
or U17237 (N_17237,N_12827,N_12829);
and U17238 (N_17238,N_14033,N_12997);
nor U17239 (N_17239,N_14843,N_14378);
and U17240 (N_17240,N_13730,N_14853);
nor U17241 (N_17241,N_13893,N_12562);
nor U17242 (N_17242,N_14173,N_13467);
nor U17243 (N_17243,N_12827,N_12739);
or U17244 (N_17244,N_14177,N_14398);
xor U17245 (N_17245,N_13859,N_12580);
nand U17246 (N_17246,N_13640,N_12870);
xnor U17247 (N_17247,N_14336,N_14499);
nand U17248 (N_17248,N_14248,N_13412);
or U17249 (N_17249,N_14447,N_13219);
xor U17250 (N_17250,N_12899,N_14718);
and U17251 (N_17251,N_14841,N_14586);
xnor U17252 (N_17252,N_14643,N_14104);
nor U17253 (N_17253,N_14100,N_13006);
or U17254 (N_17254,N_13400,N_14741);
nor U17255 (N_17255,N_14173,N_13045);
nand U17256 (N_17256,N_12749,N_14374);
or U17257 (N_17257,N_14941,N_14047);
or U17258 (N_17258,N_14234,N_13175);
xor U17259 (N_17259,N_13586,N_13215);
and U17260 (N_17260,N_14148,N_13748);
nand U17261 (N_17261,N_14713,N_12963);
or U17262 (N_17262,N_13293,N_13333);
or U17263 (N_17263,N_13962,N_14504);
nor U17264 (N_17264,N_14520,N_14020);
nor U17265 (N_17265,N_14095,N_14121);
nor U17266 (N_17266,N_14254,N_13050);
nand U17267 (N_17267,N_13500,N_12825);
or U17268 (N_17268,N_13109,N_14631);
nor U17269 (N_17269,N_14271,N_13525);
and U17270 (N_17270,N_14354,N_13726);
nor U17271 (N_17271,N_14419,N_12816);
or U17272 (N_17272,N_14383,N_12917);
or U17273 (N_17273,N_13222,N_14514);
or U17274 (N_17274,N_14864,N_14626);
and U17275 (N_17275,N_13052,N_12883);
nor U17276 (N_17276,N_13864,N_14990);
or U17277 (N_17277,N_13555,N_14716);
xor U17278 (N_17278,N_13022,N_13301);
xnor U17279 (N_17279,N_14341,N_14707);
or U17280 (N_17280,N_13688,N_13135);
nand U17281 (N_17281,N_13769,N_12627);
and U17282 (N_17282,N_13606,N_13774);
nor U17283 (N_17283,N_13650,N_13945);
nor U17284 (N_17284,N_14933,N_13632);
nor U17285 (N_17285,N_14794,N_14325);
xnor U17286 (N_17286,N_14476,N_14663);
or U17287 (N_17287,N_13123,N_13402);
xor U17288 (N_17288,N_14917,N_13836);
nor U17289 (N_17289,N_12577,N_13917);
or U17290 (N_17290,N_12586,N_13137);
nand U17291 (N_17291,N_14673,N_14882);
nor U17292 (N_17292,N_12668,N_13351);
or U17293 (N_17293,N_14527,N_13063);
or U17294 (N_17294,N_13577,N_14735);
and U17295 (N_17295,N_14010,N_14942);
and U17296 (N_17296,N_13255,N_14100);
and U17297 (N_17297,N_12818,N_13130);
nand U17298 (N_17298,N_13402,N_14751);
xnor U17299 (N_17299,N_13180,N_14405);
or U17300 (N_17300,N_13910,N_13925);
nand U17301 (N_17301,N_14444,N_12855);
nand U17302 (N_17302,N_12741,N_14542);
or U17303 (N_17303,N_13356,N_13290);
nor U17304 (N_17304,N_14823,N_14300);
xnor U17305 (N_17305,N_12662,N_14706);
nor U17306 (N_17306,N_14758,N_13439);
and U17307 (N_17307,N_14593,N_12799);
xnor U17308 (N_17308,N_13450,N_13618);
nor U17309 (N_17309,N_14145,N_14161);
xnor U17310 (N_17310,N_14200,N_13348);
nand U17311 (N_17311,N_14584,N_13601);
nand U17312 (N_17312,N_13818,N_14645);
nand U17313 (N_17313,N_13390,N_12779);
or U17314 (N_17314,N_14020,N_14185);
or U17315 (N_17315,N_13667,N_14111);
or U17316 (N_17316,N_14896,N_13234);
xnor U17317 (N_17317,N_13661,N_13446);
or U17318 (N_17318,N_14926,N_14016);
nand U17319 (N_17319,N_13992,N_14264);
nor U17320 (N_17320,N_13633,N_14684);
or U17321 (N_17321,N_13748,N_13813);
and U17322 (N_17322,N_13557,N_13581);
and U17323 (N_17323,N_13974,N_13448);
and U17324 (N_17324,N_13434,N_14161);
nand U17325 (N_17325,N_14400,N_13428);
or U17326 (N_17326,N_13773,N_14559);
nor U17327 (N_17327,N_12810,N_14721);
nor U17328 (N_17328,N_14020,N_13823);
and U17329 (N_17329,N_13748,N_14205);
and U17330 (N_17330,N_13631,N_14916);
nand U17331 (N_17331,N_13756,N_12735);
nand U17332 (N_17332,N_14150,N_12636);
or U17333 (N_17333,N_14405,N_13355);
nand U17334 (N_17334,N_13150,N_12866);
xor U17335 (N_17335,N_14510,N_14975);
nand U17336 (N_17336,N_13331,N_14273);
nor U17337 (N_17337,N_14352,N_12872);
or U17338 (N_17338,N_12870,N_14116);
and U17339 (N_17339,N_14998,N_14130);
xnor U17340 (N_17340,N_12724,N_13706);
nor U17341 (N_17341,N_14718,N_13852);
nor U17342 (N_17342,N_13481,N_14653);
or U17343 (N_17343,N_14638,N_13354);
and U17344 (N_17344,N_13074,N_14069);
xor U17345 (N_17345,N_13962,N_14694);
and U17346 (N_17346,N_14304,N_14936);
or U17347 (N_17347,N_14443,N_12835);
nor U17348 (N_17348,N_13085,N_12814);
nand U17349 (N_17349,N_13272,N_14922);
nand U17350 (N_17350,N_14788,N_13004);
xnor U17351 (N_17351,N_13481,N_14679);
and U17352 (N_17352,N_13058,N_14323);
or U17353 (N_17353,N_14827,N_13868);
xor U17354 (N_17354,N_13111,N_13970);
nand U17355 (N_17355,N_13105,N_12681);
nor U17356 (N_17356,N_14540,N_14593);
nand U17357 (N_17357,N_13251,N_14788);
nand U17358 (N_17358,N_13013,N_13770);
nand U17359 (N_17359,N_12904,N_13062);
xor U17360 (N_17360,N_14639,N_12721);
nor U17361 (N_17361,N_12849,N_12674);
or U17362 (N_17362,N_14860,N_13888);
or U17363 (N_17363,N_13341,N_14295);
or U17364 (N_17364,N_14088,N_13113);
xor U17365 (N_17365,N_14274,N_14504);
nand U17366 (N_17366,N_13647,N_14048);
nand U17367 (N_17367,N_14283,N_13463);
or U17368 (N_17368,N_12840,N_13490);
and U17369 (N_17369,N_14704,N_14529);
nand U17370 (N_17370,N_13462,N_12746);
and U17371 (N_17371,N_14865,N_13546);
nand U17372 (N_17372,N_13758,N_14955);
nand U17373 (N_17373,N_12648,N_13902);
nor U17374 (N_17374,N_14878,N_14051);
or U17375 (N_17375,N_12803,N_14554);
nand U17376 (N_17376,N_14308,N_14197);
and U17377 (N_17377,N_13797,N_12939);
or U17378 (N_17378,N_12764,N_13584);
xnor U17379 (N_17379,N_14728,N_13457);
nand U17380 (N_17380,N_14776,N_12641);
nor U17381 (N_17381,N_13256,N_13240);
nor U17382 (N_17382,N_13658,N_12990);
xor U17383 (N_17383,N_13430,N_14909);
nand U17384 (N_17384,N_14380,N_14419);
nor U17385 (N_17385,N_13632,N_14436);
or U17386 (N_17386,N_13956,N_13221);
and U17387 (N_17387,N_12860,N_13071);
nor U17388 (N_17388,N_14083,N_13931);
and U17389 (N_17389,N_14689,N_13506);
xnor U17390 (N_17390,N_13633,N_14294);
or U17391 (N_17391,N_14808,N_14269);
or U17392 (N_17392,N_13137,N_14826);
xnor U17393 (N_17393,N_12785,N_13395);
and U17394 (N_17394,N_14670,N_13808);
nand U17395 (N_17395,N_13141,N_14508);
and U17396 (N_17396,N_13924,N_13191);
nor U17397 (N_17397,N_14594,N_14179);
and U17398 (N_17398,N_14281,N_12881);
or U17399 (N_17399,N_14169,N_14814);
or U17400 (N_17400,N_13824,N_14253);
xnor U17401 (N_17401,N_13420,N_14659);
and U17402 (N_17402,N_13159,N_13361);
or U17403 (N_17403,N_14263,N_14253);
or U17404 (N_17404,N_13832,N_14904);
nand U17405 (N_17405,N_13542,N_13356);
nor U17406 (N_17406,N_12920,N_14527);
xor U17407 (N_17407,N_14701,N_12533);
and U17408 (N_17408,N_14537,N_12505);
nor U17409 (N_17409,N_13176,N_13766);
nor U17410 (N_17410,N_13845,N_13057);
nor U17411 (N_17411,N_12513,N_14831);
nor U17412 (N_17412,N_14580,N_14511);
nand U17413 (N_17413,N_13899,N_12688);
xnor U17414 (N_17414,N_14434,N_13569);
xnor U17415 (N_17415,N_13799,N_13864);
nand U17416 (N_17416,N_14881,N_12598);
or U17417 (N_17417,N_14555,N_13602);
or U17418 (N_17418,N_13370,N_12976);
and U17419 (N_17419,N_14178,N_14750);
or U17420 (N_17420,N_14223,N_12781);
nand U17421 (N_17421,N_14860,N_14192);
or U17422 (N_17422,N_14800,N_13951);
and U17423 (N_17423,N_14591,N_14463);
and U17424 (N_17424,N_14679,N_13786);
or U17425 (N_17425,N_13938,N_12957);
xnor U17426 (N_17426,N_13757,N_13933);
or U17427 (N_17427,N_13394,N_14686);
xnor U17428 (N_17428,N_14216,N_12919);
nor U17429 (N_17429,N_14718,N_13408);
nor U17430 (N_17430,N_12708,N_14855);
xnor U17431 (N_17431,N_14067,N_14889);
nand U17432 (N_17432,N_13068,N_13968);
nand U17433 (N_17433,N_12748,N_14279);
and U17434 (N_17434,N_14645,N_12987);
nand U17435 (N_17435,N_14225,N_12538);
nand U17436 (N_17436,N_12510,N_12874);
or U17437 (N_17437,N_13537,N_13805);
xor U17438 (N_17438,N_13199,N_13236);
nor U17439 (N_17439,N_14234,N_13675);
nand U17440 (N_17440,N_12736,N_12913);
or U17441 (N_17441,N_13520,N_14874);
nor U17442 (N_17442,N_13221,N_14269);
nor U17443 (N_17443,N_12880,N_13659);
or U17444 (N_17444,N_14124,N_14543);
and U17445 (N_17445,N_14079,N_13982);
and U17446 (N_17446,N_13789,N_14013);
nor U17447 (N_17447,N_14051,N_14993);
nand U17448 (N_17448,N_14870,N_12540);
nand U17449 (N_17449,N_13393,N_13725);
nand U17450 (N_17450,N_14924,N_12666);
nand U17451 (N_17451,N_14791,N_14201);
or U17452 (N_17452,N_13869,N_13974);
nand U17453 (N_17453,N_12817,N_13845);
nand U17454 (N_17454,N_14102,N_14076);
or U17455 (N_17455,N_13776,N_14595);
or U17456 (N_17456,N_13042,N_13210);
or U17457 (N_17457,N_13099,N_14944);
or U17458 (N_17458,N_14768,N_14509);
nand U17459 (N_17459,N_14385,N_12822);
nor U17460 (N_17460,N_14709,N_14797);
or U17461 (N_17461,N_13610,N_12755);
nand U17462 (N_17462,N_14839,N_14278);
xnor U17463 (N_17463,N_14014,N_12754);
or U17464 (N_17464,N_12804,N_14428);
nand U17465 (N_17465,N_13185,N_14153);
and U17466 (N_17466,N_14391,N_14285);
xor U17467 (N_17467,N_13270,N_13475);
nand U17468 (N_17468,N_13905,N_13096);
and U17469 (N_17469,N_14641,N_13873);
xor U17470 (N_17470,N_13398,N_12652);
and U17471 (N_17471,N_13033,N_14073);
nor U17472 (N_17472,N_14970,N_13111);
nor U17473 (N_17473,N_13071,N_13782);
nand U17474 (N_17474,N_14251,N_14129);
or U17475 (N_17475,N_13513,N_14851);
xnor U17476 (N_17476,N_13950,N_14951);
or U17477 (N_17477,N_14440,N_12895);
and U17478 (N_17478,N_12513,N_13419);
or U17479 (N_17479,N_13981,N_13518);
or U17480 (N_17480,N_14333,N_12844);
xnor U17481 (N_17481,N_13839,N_13263);
nand U17482 (N_17482,N_14501,N_13439);
nor U17483 (N_17483,N_14975,N_12937);
nand U17484 (N_17484,N_13653,N_13450);
or U17485 (N_17485,N_12776,N_13596);
nand U17486 (N_17486,N_14162,N_13523);
nand U17487 (N_17487,N_12959,N_13190);
or U17488 (N_17488,N_14592,N_14254);
nand U17489 (N_17489,N_12867,N_13224);
and U17490 (N_17490,N_13035,N_12535);
nor U17491 (N_17491,N_14565,N_14653);
xor U17492 (N_17492,N_13519,N_12809);
nand U17493 (N_17493,N_13078,N_12921);
nor U17494 (N_17494,N_14161,N_12687);
nand U17495 (N_17495,N_13410,N_14825);
nand U17496 (N_17496,N_13130,N_12886);
or U17497 (N_17497,N_14541,N_13385);
and U17498 (N_17498,N_14881,N_14837);
and U17499 (N_17499,N_12612,N_13408);
or U17500 (N_17500,N_17448,N_16377);
or U17501 (N_17501,N_15025,N_16132);
xor U17502 (N_17502,N_16606,N_15766);
or U17503 (N_17503,N_16928,N_17468);
and U17504 (N_17504,N_15224,N_15537);
nor U17505 (N_17505,N_15395,N_16618);
xor U17506 (N_17506,N_15273,N_16477);
nand U17507 (N_17507,N_16411,N_16648);
or U17508 (N_17508,N_15062,N_16898);
nor U17509 (N_17509,N_15606,N_15105);
or U17510 (N_17510,N_17376,N_17357);
or U17511 (N_17511,N_15049,N_16322);
or U17512 (N_17512,N_17186,N_15467);
xnor U17513 (N_17513,N_16050,N_15861);
nand U17514 (N_17514,N_16067,N_16309);
xor U17515 (N_17515,N_15250,N_15800);
nand U17516 (N_17516,N_16273,N_17205);
xor U17517 (N_17517,N_15389,N_16524);
xor U17518 (N_17518,N_16634,N_15318);
and U17519 (N_17519,N_16848,N_17447);
nor U17520 (N_17520,N_15840,N_17259);
or U17521 (N_17521,N_16741,N_15540);
nor U17522 (N_17522,N_16931,N_16297);
or U17523 (N_17523,N_15297,N_16265);
nand U17524 (N_17524,N_15447,N_16123);
and U17525 (N_17525,N_15039,N_15289);
and U17526 (N_17526,N_17358,N_15698);
nand U17527 (N_17527,N_15979,N_16417);
or U17528 (N_17528,N_15917,N_15108);
nor U17529 (N_17529,N_16504,N_15975);
or U17530 (N_17530,N_16399,N_17207);
xor U17531 (N_17531,N_17200,N_15076);
and U17532 (N_17532,N_16646,N_16983);
xnor U17533 (N_17533,N_17002,N_16760);
nand U17534 (N_17534,N_15130,N_15786);
nor U17535 (N_17535,N_15860,N_17393);
nor U17536 (N_17536,N_16320,N_15689);
and U17537 (N_17537,N_16497,N_16304);
and U17538 (N_17538,N_16246,N_15521);
and U17539 (N_17539,N_17096,N_16144);
xor U17540 (N_17540,N_16193,N_16012);
xor U17541 (N_17541,N_15134,N_16861);
and U17542 (N_17542,N_17389,N_15003);
xnor U17543 (N_17543,N_15191,N_16856);
nor U17544 (N_17544,N_15822,N_16323);
and U17545 (N_17545,N_15737,N_17435);
xnor U17546 (N_17546,N_16083,N_16074);
and U17547 (N_17547,N_15077,N_15805);
or U17548 (N_17548,N_16667,N_15534);
and U17549 (N_17549,N_15332,N_15645);
nand U17550 (N_17550,N_15608,N_15502);
nand U17551 (N_17551,N_15122,N_16576);
nand U17552 (N_17552,N_16212,N_15754);
nand U17553 (N_17553,N_16626,N_16813);
or U17554 (N_17554,N_16156,N_17400);
and U17555 (N_17555,N_16680,N_16272);
xnor U17556 (N_17556,N_15053,N_16047);
nor U17557 (N_17557,N_16126,N_15022);
nand U17558 (N_17558,N_17165,N_17007);
nor U17559 (N_17559,N_15565,N_16247);
and U17560 (N_17560,N_16435,N_16048);
nand U17561 (N_17561,N_16698,N_15222);
and U17562 (N_17562,N_16799,N_17113);
or U17563 (N_17563,N_17278,N_16117);
xor U17564 (N_17564,N_15402,N_15387);
and U17565 (N_17565,N_16260,N_15765);
xnor U17566 (N_17566,N_15489,N_17341);
nor U17567 (N_17567,N_17420,N_15528);
nor U17568 (N_17568,N_15089,N_16054);
or U17569 (N_17569,N_15519,N_15581);
or U17570 (N_17570,N_16287,N_16657);
nand U17571 (N_17571,N_16881,N_17204);
and U17572 (N_17572,N_15662,N_15201);
nor U17573 (N_17573,N_17212,N_17285);
or U17574 (N_17574,N_16505,N_16714);
xnor U17575 (N_17575,N_17330,N_16089);
or U17576 (N_17576,N_15738,N_16575);
or U17577 (N_17577,N_15789,N_16990);
xor U17578 (N_17578,N_15441,N_15562);
nor U17579 (N_17579,N_15398,N_16356);
nand U17580 (N_17580,N_15729,N_17059);
and U17581 (N_17581,N_15769,N_15004);
and U17582 (N_17582,N_15679,N_15094);
and U17583 (N_17583,N_15506,N_16883);
and U17584 (N_17584,N_16864,N_15811);
nand U17585 (N_17585,N_15329,N_17168);
nand U17586 (N_17586,N_15381,N_15020);
nand U17587 (N_17587,N_15604,N_15874);
nor U17588 (N_17588,N_16368,N_16347);
or U17589 (N_17589,N_16224,N_16199);
nor U17590 (N_17590,N_16364,N_17099);
and U17591 (N_17591,N_16758,N_15964);
or U17592 (N_17592,N_17078,N_16652);
nand U17593 (N_17593,N_17225,N_17156);
and U17594 (N_17594,N_15196,N_17060);
and U17595 (N_17595,N_16059,N_15579);
nor U17596 (N_17596,N_16078,N_16527);
and U17597 (N_17597,N_16404,N_15223);
or U17598 (N_17598,N_17344,N_16509);
nor U17599 (N_17599,N_15696,N_16939);
or U17600 (N_17600,N_16984,N_16540);
and U17601 (N_17601,N_15166,N_16027);
nand U17602 (N_17602,N_17157,N_15192);
nand U17603 (N_17603,N_17049,N_15001);
nor U17604 (N_17604,N_15051,N_16807);
or U17605 (N_17605,N_16378,N_15624);
and U17606 (N_17606,N_16619,N_16585);
nand U17607 (N_17607,N_17419,N_17459);
and U17608 (N_17608,N_16623,N_17476);
and U17609 (N_17609,N_15055,N_16985);
nand U17610 (N_17610,N_16582,N_16907);
or U17611 (N_17611,N_16070,N_17114);
or U17612 (N_17612,N_17401,N_16029);
xnor U17613 (N_17613,N_17016,N_17137);
and U17614 (N_17614,N_16017,N_17479);
xnor U17615 (N_17615,N_15732,N_15850);
or U17616 (N_17616,N_15072,N_17245);
xor U17617 (N_17617,N_16361,N_15725);
and U17618 (N_17618,N_16837,N_16946);
and U17619 (N_17619,N_16024,N_15873);
and U17620 (N_17620,N_16607,N_16281);
xor U17621 (N_17621,N_16266,N_16267);
and U17622 (N_17622,N_15995,N_15203);
and U17623 (N_17623,N_17219,N_16337);
nand U17624 (N_17624,N_16009,N_15199);
nand U17625 (N_17625,N_15948,N_15981);
nand U17626 (N_17626,N_15317,N_17230);
nor U17627 (N_17627,N_17035,N_16120);
nand U17628 (N_17628,N_17295,N_15205);
nand U17629 (N_17629,N_15002,N_17170);
and U17630 (N_17630,N_16348,N_15755);
nor U17631 (N_17631,N_16778,N_16472);
nand U17632 (N_17632,N_16002,N_16092);
or U17633 (N_17633,N_15690,N_16581);
and U17634 (N_17634,N_16484,N_15971);
nand U17635 (N_17635,N_16995,N_16787);
nand U17636 (N_17636,N_15556,N_15287);
nor U17637 (N_17637,N_16410,N_16063);
nor U17638 (N_17638,N_15504,N_15063);
nor U17639 (N_17639,N_17257,N_15328);
nand U17640 (N_17640,N_17343,N_16234);
or U17641 (N_17641,N_17196,N_15268);
or U17642 (N_17642,N_15272,N_16970);
nor U17643 (N_17643,N_15911,N_15079);
nand U17644 (N_17644,N_15631,N_16537);
nand U17645 (N_17645,N_15210,N_15548);
xor U17646 (N_17646,N_15838,N_15292);
nand U17647 (N_17647,N_16904,N_15591);
nor U17648 (N_17648,N_15980,N_15070);
nand U17649 (N_17649,N_17377,N_16616);
nand U17650 (N_17650,N_16510,N_17471);
nor U17651 (N_17651,N_16767,N_16419);
or U17652 (N_17652,N_15507,N_17098);
xnor U17653 (N_17653,N_15152,N_17406);
and U17654 (N_17654,N_16747,N_17014);
xor U17655 (N_17655,N_15773,N_17409);
and U17656 (N_17656,N_15875,N_15877);
nor U17657 (N_17657,N_16157,N_16955);
xor U17658 (N_17658,N_16906,N_15054);
nor U17659 (N_17659,N_16519,N_15969);
nor U17660 (N_17660,N_16525,N_15307);
xor U17661 (N_17661,N_16206,N_16895);
xnor U17662 (N_17662,N_15028,N_16943);
nor U17663 (N_17663,N_16911,N_16423);
nand U17664 (N_17664,N_17314,N_17130);
nand U17665 (N_17665,N_16232,N_15753);
nand U17666 (N_17666,N_16683,N_15081);
nand U17667 (N_17667,N_15139,N_17206);
nor U17668 (N_17668,N_15177,N_15869);
nor U17669 (N_17669,N_15988,N_17457);
and U17670 (N_17670,N_15767,N_15339);
nand U17671 (N_17671,N_17227,N_16549);
xnor U17672 (N_17672,N_16069,N_16737);
and U17673 (N_17673,N_15867,N_15804);
or U17674 (N_17674,N_15904,N_15090);
xor U17675 (N_17675,N_17005,N_16820);
nor U17676 (N_17676,N_15570,N_15693);
xnor U17677 (N_17677,N_16960,N_15324);
xor U17678 (N_17678,N_15728,N_17260);
nor U17679 (N_17679,N_17316,N_15095);
xnor U17680 (N_17680,N_17410,N_17361);
nand U17681 (N_17681,N_16730,N_16553);
and U17682 (N_17682,N_15891,N_17199);
nor U17683 (N_17683,N_16969,N_15116);
and U17684 (N_17684,N_17485,N_15849);
nor U17685 (N_17685,N_15087,N_16044);
xor U17686 (N_17686,N_17082,N_15279);
and U17687 (N_17687,N_17001,N_15516);
xnor U17688 (N_17688,N_16244,N_15684);
nand U17689 (N_17689,N_16803,N_16629);
nor U17690 (N_17690,N_15270,N_15644);
or U17691 (N_17691,N_15910,N_16798);
xor U17692 (N_17692,N_17434,N_16682);
and U17693 (N_17693,N_16631,N_16200);
xor U17694 (N_17694,N_16021,N_16049);
nor U17695 (N_17695,N_15385,N_17027);
xnor U17696 (N_17696,N_15791,N_16727);
nand U17697 (N_17697,N_15675,N_16738);
or U17698 (N_17698,N_16420,N_15221);
nand U17699 (N_17699,N_17415,N_15851);
or U17700 (N_17700,N_17104,N_15623);
and U17701 (N_17701,N_15550,N_16494);
and U17702 (N_17702,N_16734,N_17238);
and U17703 (N_17703,N_16408,N_17412);
nand U17704 (N_17704,N_15554,N_15155);
or U17705 (N_17705,N_17092,N_16324);
nand U17706 (N_17706,N_16192,N_16489);
nor U17707 (N_17707,N_15060,N_16233);
and U17708 (N_17708,N_16498,N_15425);
nor U17709 (N_17709,N_16901,N_15702);
nor U17710 (N_17710,N_17369,N_17497);
xor U17711 (N_17711,N_17375,N_16174);
nand U17712 (N_17712,N_15123,N_15240);
nand U17713 (N_17713,N_16994,N_15058);
and U17714 (N_17714,N_15341,N_15311);
nor U17715 (N_17715,N_16301,N_15494);
xor U17716 (N_17716,N_17045,N_15371);
nand U17717 (N_17717,N_15589,N_15496);
xor U17718 (N_17718,N_15430,N_15140);
xnor U17719 (N_17719,N_16896,N_16215);
nor U17720 (N_17720,N_17129,N_16674);
or U17721 (N_17721,N_15300,N_16934);
and U17722 (N_17722,N_17193,N_16467);
nand U17723 (N_17723,N_17475,N_15573);
and U17724 (N_17724,N_16830,N_16314);
nor U17725 (N_17725,N_16141,N_17011);
nor U17726 (N_17726,N_17179,N_16339);
nand U17727 (N_17727,N_16045,N_16219);
or U17728 (N_17728,N_16022,N_15484);
xnor U17729 (N_17729,N_15687,N_15056);
nand U17730 (N_17730,N_15012,N_15626);
nor U17731 (N_17731,N_17181,N_17152);
and U17732 (N_17732,N_16902,N_16279);
and U17733 (N_17733,N_16713,N_15437);
xnor U17734 (N_17734,N_15609,N_16603);
and U17735 (N_17735,N_16086,N_15463);
xor U17736 (N_17736,N_16468,N_16428);
xor U17737 (N_17737,N_15460,N_15774);
nand U17738 (N_17738,N_15383,N_16940);
nand U17739 (N_17739,N_16613,N_16333);
or U17740 (N_17740,N_15067,N_16298);
nand U17741 (N_17741,N_15149,N_15432);
or U17742 (N_17742,N_16222,N_16715);
xnor U17743 (N_17743,N_15816,N_16046);
or U17744 (N_17744,N_16572,N_15459);
nor U17745 (N_17745,N_16143,N_16185);
nor U17746 (N_17746,N_16521,N_17110);
nand U17747 (N_17747,N_16796,N_16443);
nand U17748 (N_17748,N_15741,N_17301);
nand U17749 (N_17749,N_17483,N_17440);
nor U17750 (N_17750,N_15065,N_16513);
or U17751 (N_17751,N_16614,N_17154);
nor U17752 (N_17752,N_16753,N_16073);
xor U17753 (N_17753,N_16422,N_17058);
nand U17754 (N_17754,N_16407,N_15600);
and U17755 (N_17755,N_16186,N_16914);
nand U17756 (N_17756,N_16462,N_15450);
nand U17757 (N_17757,N_15832,N_16668);
or U17758 (N_17758,N_15170,N_16128);
nor U17759 (N_17759,N_16599,N_15319);
nand U17760 (N_17760,N_15595,N_15135);
and U17761 (N_17761,N_16712,N_17489);
or U17762 (N_17762,N_16094,N_16036);
xor U17763 (N_17763,N_16366,N_16355);
or U17764 (N_17764,N_15726,N_16650);
and U17765 (N_17765,N_17438,N_17499);
nor U17766 (N_17766,N_16016,N_17022);
xnor U17767 (N_17767,N_15985,N_15704);
xor U17768 (N_17768,N_17090,N_17074);
nand U17769 (N_17769,N_16863,N_16884);
nand U17770 (N_17770,N_17167,N_15209);
nor U17771 (N_17771,N_15742,N_15491);
nand U17772 (N_17772,N_15949,N_15409);
or U17773 (N_17773,N_16000,N_15603);
xnor U17774 (N_17774,N_15808,N_15173);
xor U17775 (N_17775,N_15740,N_15810);
nand U17776 (N_17776,N_16845,N_16439);
xor U17777 (N_17777,N_16085,N_15715);
and U17778 (N_17778,N_16485,N_15705);
xor U17779 (N_17779,N_16291,N_16033);
nor U17780 (N_17780,N_16925,N_16312);
nand U17781 (N_17781,N_15040,N_15453);
or U17782 (N_17782,N_15627,N_17124);
nand U17783 (N_17783,N_15780,N_16349);
xor U17784 (N_17784,N_16950,N_15700);
or U17785 (N_17785,N_17408,N_17055);
xnor U17786 (N_17786,N_15817,N_16146);
xor U17787 (N_17787,N_15227,N_15326);
or U17788 (N_17788,N_17398,N_15636);
or U17789 (N_17789,N_16963,N_15617);
and U17790 (N_17790,N_16604,N_15331);
or U17791 (N_17791,N_15370,N_16814);
nand U17792 (N_17792,N_17122,N_15819);
xor U17793 (N_17793,N_16353,N_16104);
xor U17794 (N_17794,N_17056,N_16373);
xnor U17795 (N_17795,N_16892,N_15593);
and U17796 (N_17796,N_16724,N_15306);
xnor U17797 (N_17797,N_15871,N_17378);
nand U17798 (N_17798,N_17033,N_17272);
nor U17799 (N_17799,N_15634,N_16563);
or U17800 (N_17800,N_16098,N_15750);
nand U17801 (N_17801,N_17454,N_17392);
or U17802 (N_17802,N_15778,N_16557);
or U17803 (N_17803,N_17224,N_15336);
xor U17804 (N_17804,N_17148,N_15366);
xnor U17805 (N_17805,N_17150,N_16989);
or U17806 (N_17806,N_16437,N_15722);
nor U17807 (N_17807,N_15234,N_16460);
xnor U17808 (N_17808,N_15934,N_15179);
nand U17809 (N_17809,N_16728,N_15423);
nand U17810 (N_17810,N_16037,N_15872);
nand U17811 (N_17811,N_15796,N_15085);
xor U17812 (N_17812,N_16153,N_17450);
or U17813 (N_17813,N_16122,N_17388);
nand U17814 (N_17814,N_16823,N_16427);
nand U17815 (N_17815,N_16384,N_15847);
and U17816 (N_17816,N_15416,N_16426);
nor U17817 (N_17817,N_17387,N_17268);
nor U17818 (N_17818,N_17243,N_15375);
nand U17819 (N_17819,N_15782,N_16538);
nor U17820 (N_17820,N_15165,N_16360);
xnor U17821 (N_17821,N_16751,N_15878);
nand U17822 (N_17822,N_17432,N_15345);
xnor U17823 (N_17823,N_17477,N_16996);
nand U17824 (N_17824,N_15731,N_15527);
and U17825 (N_17825,N_16262,N_15577);
or U17826 (N_17826,N_16066,N_15592);
nor U17827 (N_17827,N_15440,N_17337);
or U17828 (N_17828,N_17094,N_15315);
nor U17829 (N_17829,N_16729,N_15661);
xor U17830 (N_17830,N_15957,N_16237);
and U17831 (N_17831,N_16469,N_17403);
or U17832 (N_17832,N_15610,N_16697);
nand U17833 (N_17833,N_16953,N_15515);
nor U17834 (N_17834,N_16295,N_15490);
nand U17835 (N_17835,N_17293,N_15566);
nand U17836 (N_17836,N_16238,N_16545);
xnor U17837 (N_17837,N_15812,N_17372);
xor U17838 (N_17838,N_16843,N_17057);
and U17839 (N_17839,N_15935,N_15378);
and U17840 (N_17840,N_15730,N_15718);
xnor U17841 (N_17841,N_16303,N_15543);
or U17842 (N_17842,N_16555,N_15455);
xnor U17843 (N_17843,N_15555,N_16152);
xnor U17844 (N_17844,N_16177,N_15266);
or U17845 (N_17845,N_15772,N_17313);
and U17846 (N_17846,N_16535,N_15184);
xnor U17847 (N_17847,N_15427,N_17211);
xnor U17848 (N_17848,N_16750,N_16182);
nor U17849 (N_17849,N_16035,N_15466);
or U17850 (N_17850,N_15893,N_15043);
nand U17851 (N_17851,N_15733,N_16025);
nor U17852 (N_17852,N_15285,N_15362);
and U17853 (N_17853,N_16701,N_15924);
xor U17854 (N_17854,N_16775,N_15674);
and U17855 (N_17855,N_16254,N_16255);
nand U17856 (N_17856,N_16721,N_16743);
and U17857 (N_17857,N_17445,N_15508);
nor U17858 (N_17858,N_15676,N_15866);
nand U17859 (N_17859,N_15121,N_15312);
nand U17860 (N_17860,N_15202,N_15106);
nor U17861 (N_17861,N_17010,N_16972);
nand U17862 (N_17862,N_16844,N_15158);
nand U17863 (N_17863,N_16197,N_15894);
or U17864 (N_17864,N_15410,N_15906);
nor U17865 (N_17865,N_15656,N_17487);
and U17866 (N_17866,N_17048,N_16442);
or U17867 (N_17867,N_16586,N_15172);
and U17868 (N_17868,N_15779,N_17101);
and U17869 (N_17869,N_16294,N_16293);
nor U17870 (N_17870,N_16615,N_16717);
nand U17871 (N_17871,N_16057,N_17021);
xnor U17872 (N_17872,N_17315,N_15044);
or U17873 (N_17873,N_15241,N_15369);
xnor U17874 (N_17874,N_15833,N_15628);
xnor U17875 (N_17875,N_15294,N_17080);
nor U17876 (N_17876,N_15288,N_16894);
or U17877 (N_17877,N_15278,N_16154);
nand U17878 (N_17878,N_15218,N_16877);
nand U17879 (N_17879,N_15783,N_15193);
nand U17880 (N_17880,N_16371,N_15686);
or U17881 (N_17881,N_16159,N_17063);
or U17882 (N_17882,N_16833,N_16080);
nand U17883 (N_17883,N_16811,N_16447);
nand U17884 (N_17884,N_15436,N_16097);
and U17885 (N_17885,N_15126,N_15763);
and U17886 (N_17886,N_17362,N_16374);
nor U17887 (N_17887,N_15228,N_16998);
nor U17888 (N_17888,N_16478,N_16782);
xor U17889 (N_17889,N_16250,N_17198);
xnor U17890 (N_17890,N_15485,N_16138);
xor U17891 (N_17891,N_15807,N_16913);
and U17892 (N_17892,N_15298,N_17202);
nand U17893 (N_17893,N_17395,N_15276);
nand U17894 (N_17894,N_15259,N_17474);
nor U17895 (N_17895,N_16957,N_17303);
nand U17896 (N_17896,N_15439,N_15185);
and U17897 (N_17897,N_16779,N_15394);
nor U17898 (N_17898,N_17026,N_17134);
and U17899 (N_17899,N_16058,N_15344);
xor U17900 (N_17900,N_15762,N_15029);
xor U17901 (N_17901,N_17418,N_15182);
and U17902 (N_17902,N_17064,N_16413);
nor U17903 (N_17903,N_17201,N_16474);
nor U17904 (N_17904,N_16819,N_15413);
or U17905 (N_17905,N_16841,N_15225);
nor U17906 (N_17906,N_16882,N_16274);
nor U17907 (N_17907,N_15136,N_17384);
xor U17908 (N_17908,N_16261,N_16305);
xor U17909 (N_17909,N_16018,N_16430);
nand U17910 (N_17910,N_15846,N_17276);
and U17911 (N_17911,N_15982,N_15658);
nor U17912 (N_17912,N_15163,N_16429);
or U17913 (N_17913,N_16772,N_16038);
xor U17914 (N_17914,N_17332,N_15734);
nand U17915 (N_17915,N_17373,N_15015);
nand U17916 (N_17916,N_16597,N_16825);
nand U17917 (N_17917,N_15009,N_16006);
or U17918 (N_17918,N_15560,N_16977);
nor U17919 (N_17919,N_16664,N_15213);
or U17920 (N_17920,N_16554,N_17484);
xor U17921 (N_17921,N_15882,N_16321);
and U17922 (N_17922,N_17486,N_15751);
and U17923 (N_17923,N_16511,N_16973);
or U17924 (N_17924,N_16687,N_15187);
nor U17925 (N_17925,N_16948,N_15613);
xnor U17926 (N_17926,N_16887,N_16308);
xnor U17927 (N_17927,N_16167,N_16662);
nor U17928 (N_17928,N_16005,N_17283);
xor U17929 (N_17929,N_16195,N_16096);
or U17930 (N_17930,N_15921,N_16180);
or U17931 (N_17931,N_17149,N_15124);
nor U17932 (N_17932,N_17284,N_15803);
nand U17933 (N_17933,N_16139,N_16201);
or U17934 (N_17934,N_16531,N_15073);
or U17935 (N_17935,N_16490,N_15137);
or U17936 (N_17936,N_15444,N_16453);
nor U17937 (N_17937,N_17191,N_15501);
nand U17938 (N_17938,N_15446,N_17436);
xor U17939 (N_17939,N_16380,N_16552);
nor U17940 (N_17940,N_16952,N_15238);
nor U17941 (N_17941,N_15792,N_16720);
nor U17942 (N_17942,N_16269,N_16259);
and U17943 (N_17943,N_16726,N_16190);
nor U17944 (N_17944,N_17494,N_16745);
nor U17945 (N_17945,N_17430,N_15093);
and U17946 (N_17946,N_15113,N_16396);
nand U17947 (N_17947,N_16971,N_17309);
nand U17948 (N_17948,N_17009,N_17032);
nor U17949 (N_17949,N_16391,N_15518);
nand U17950 (N_17950,N_17209,N_15230);
nor U17951 (N_17951,N_15468,N_15414);
nor U17952 (N_17952,N_15876,N_17119);
or U17953 (N_17953,N_16444,N_17380);
nand U17954 (N_17954,N_16529,N_16740);
and U17955 (N_17955,N_17465,N_15434);
nor U17956 (N_17956,N_16935,N_15724);
nand U17957 (N_17957,N_15900,N_15034);
xnor U17958 (N_17958,N_15487,N_17472);
nor U17959 (N_17959,N_15342,N_15277);
nor U17960 (N_17960,N_16785,N_16622);
xor U17961 (N_17961,N_15488,N_15647);
and U17962 (N_17962,N_16431,N_17121);
and U17963 (N_17963,N_15781,N_15057);
nand U17964 (N_17964,N_17139,N_15069);
nand U17965 (N_17965,N_17405,N_15244);
and U17966 (N_17966,N_16533,N_16452);
or U17967 (N_17967,N_16240,N_15358);
xor U17968 (N_17968,N_17107,N_15157);
nor U17969 (N_17969,N_15016,N_15933);
or U17970 (N_17970,N_15403,N_15156);
or U17971 (N_17971,N_17287,N_15181);
and U17972 (N_17972,N_16210,N_16547);
xnor U17973 (N_17973,N_15974,N_16241);
nor U17974 (N_17974,N_16860,N_16577);
or U17975 (N_17975,N_15707,N_16317);
or U17976 (N_17976,N_15685,N_15760);
and U17977 (N_17977,N_15408,N_15212);
nor U17978 (N_17978,N_16363,N_16627);
or U17979 (N_17979,N_16824,N_15945);
xor U17980 (N_17980,N_16327,N_16661);
nand U17981 (N_17981,N_15902,N_15844);
xnor U17982 (N_17982,N_16561,N_15236);
xor U17983 (N_17983,N_16655,N_16810);
or U17984 (N_17984,N_15598,N_16299);
nand U17985 (N_17985,N_16885,N_17299);
and U17986 (N_17986,N_17034,N_16217);
and U17987 (N_17987,N_15552,N_15839);
and U17988 (N_17988,N_17173,N_15481);
and U17989 (N_17989,N_17282,N_16744);
nand U17990 (N_17990,N_15913,N_17239);
nand U17991 (N_17991,N_16169,N_15574);
xnor U17992 (N_17992,N_15880,N_16409);
and U17993 (N_17993,N_15611,N_15190);
nor U17994 (N_17994,N_16358,N_15952);
or U17995 (N_17995,N_16220,N_15903);
or U17996 (N_17996,N_16328,N_16506);
nand U17997 (N_17997,N_15084,N_15918);
xnor U17998 (N_17998,N_15007,N_15545);
nor U17999 (N_17999,N_17345,N_15367);
nor U18000 (N_18000,N_15111,N_16475);
or U18001 (N_18001,N_15042,N_16838);
and U18002 (N_18002,N_17294,N_17297);
nand U18003 (N_18003,N_16993,N_15448);
nor U18004 (N_18004,N_15264,N_16013);
nor U18005 (N_18005,N_17370,N_17146);
and U18006 (N_18006,N_15271,N_16578);
xnor U18007 (N_18007,N_15989,N_16258);
or U18008 (N_18008,N_16216,N_17300);
or U18009 (N_18009,N_15586,N_17462);
nand U18010 (N_18010,N_15727,N_16644);
or U18011 (N_18011,N_15118,N_15396);
xnor U18012 (N_18012,N_17103,N_15529);
nand U18013 (N_18013,N_16082,N_17320);
nor U18014 (N_18014,N_16056,N_17171);
or U18015 (N_18015,N_17237,N_15691);
xor U18016 (N_18016,N_16277,N_15777);
nand U18017 (N_18017,N_16592,N_16161);
xnor U18018 (N_18018,N_15976,N_15021);
nor U18019 (N_18019,N_15997,N_17258);
and U18020 (N_18020,N_16875,N_16310);
nor U18021 (N_18021,N_16670,N_16111);
nor U18022 (N_18022,N_16672,N_17052);
nand U18023 (N_18023,N_17267,N_15119);
xor U18024 (N_18024,N_17087,N_15712);
and U18025 (N_18025,N_17086,N_16988);
or U18026 (N_18026,N_16776,N_16570);
xor U18027 (N_18027,N_16099,N_15401);
nor U18028 (N_18028,N_16568,N_16754);
and U18029 (N_18029,N_15831,N_16736);
and U18030 (N_18030,N_17469,N_17428);
and U18031 (N_18031,N_16105,N_15257);
nor U18032 (N_18032,N_17286,N_16802);
nor U18033 (N_18033,N_16286,N_16677);
xor U18034 (N_18034,N_16397,N_16432);
and U18035 (N_18035,N_17414,N_17037);
or U18036 (N_18036,N_16815,N_16797);
and U18037 (N_18037,N_15036,N_16765);
and U18038 (N_18038,N_15665,N_15511);
xnor U18039 (N_18039,N_15245,N_15513);
or U18040 (N_18040,N_16264,N_15252);
nand U18041 (N_18041,N_16756,N_16981);
nor U18042 (N_18042,N_15884,N_16365);
nor U18043 (N_18043,N_15648,N_16958);
nand U18044 (N_18044,N_15098,N_15078);
nor U18045 (N_18045,N_16704,N_15443);
nand U18046 (N_18046,N_17091,N_15642);
nor U18047 (N_18047,N_15219,N_16956);
nor U18048 (N_18048,N_15350,N_16019);
nor U18049 (N_18049,N_16415,N_16938);
nand U18050 (N_18050,N_15823,N_17263);
or U18051 (N_18051,N_16868,N_16486);
nand U18052 (N_18052,N_17453,N_15886);
nand U18053 (N_18053,N_15670,N_16163);
xor U18054 (N_18054,N_16421,N_16878);
nand U18055 (N_18055,N_16112,N_15563);
xor U18056 (N_18056,N_16857,N_16596);
or U18057 (N_18057,N_15602,N_16296);
xnor U18058 (N_18058,N_16659,N_16214);
and U18059 (N_18059,N_16658,N_15097);
nand U18060 (N_18060,N_16318,N_16449);
or U18061 (N_18061,N_17456,N_17366);
xnor U18062 (N_18062,N_15357,N_16542);
xnor U18063 (N_18063,N_15770,N_15462);
nand U18064 (N_18064,N_15638,N_15164);
xnor U18065 (N_18065,N_16976,N_17070);
nand U18066 (N_18066,N_16155,N_16283);
nor U18067 (N_18067,N_15061,N_16937);
and U18068 (N_18068,N_15499,N_15129);
and U18069 (N_18069,N_16909,N_16459);
and U18070 (N_18070,N_17273,N_17163);
nand U18071 (N_18071,N_15825,N_15154);
xnor U18072 (N_18072,N_15692,N_15486);
nor U18073 (N_18073,N_16307,N_16425);
xor U18074 (N_18074,N_15435,N_17394);
xnor U18075 (N_18075,N_16218,N_17397);
or U18076 (N_18076,N_16921,N_16381);
and U18077 (N_18077,N_15605,N_15709);
xnor U18078 (N_18078,N_15887,N_16891);
xor U18079 (N_18079,N_15359,N_15597);
nand U18080 (N_18080,N_17252,N_15338);
nand U18081 (N_18081,N_17274,N_16718);
nor U18082 (N_18082,N_16788,N_16929);
nor U18083 (N_18083,N_17416,N_15785);
xnor U18084 (N_18084,N_16330,N_16870);
or U18085 (N_18085,N_16383,N_15788);
xnor U18086 (N_18086,N_16762,N_16242);
nand U18087 (N_18087,N_16023,N_17463);
nor U18088 (N_18088,N_15747,N_16665);
nand U18089 (N_18089,N_16532,N_16918);
and U18090 (N_18090,N_17351,N_15281);
and U18091 (N_18091,N_17160,N_16580);
xnor U18092 (N_18092,N_15551,N_15682);
and U18093 (N_18093,N_16978,N_17017);
xnor U18094 (N_18094,N_15046,N_15719);
xor U18095 (N_18095,N_16367,N_15008);
and U18096 (N_18096,N_17144,N_17019);
nor U18097 (N_18097,N_16862,N_16703);
xor U18098 (N_18098,N_15461,N_15207);
or U18099 (N_18099,N_15784,N_15445);
xnor U18100 (N_18100,N_16424,N_16418);
or U18101 (N_18101,N_17085,N_16800);
nor U18102 (N_18102,N_15759,N_16731);
and U18103 (N_18103,N_15428,N_15038);
nor U18104 (N_18104,N_16643,N_17155);
xor U18105 (N_18105,N_16487,N_17190);
and U18106 (N_18106,N_16926,N_16357);
nor U18107 (N_18107,N_16786,N_16847);
nand U18108 (N_18108,N_17417,N_16528);
or U18109 (N_18109,N_17251,N_16839);
nor U18110 (N_18110,N_15836,N_17495);
and U18111 (N_18111,N_15128,N_15286);
xor U18112 (N_18112,N_15100,N_17184);
and U18113 (N_18113,N_15478,N_17030);
nand U18114 (N_18114,N_15930,N_15291);
nand U18115 (N_18115,N_17047,N_16759);
or U18116 (N_18116,N_16932,N_16346);
or U18117 (N_18117,N_16865,N_15701);
or U18118 (N_18118,N_15965,N_16311);
and U18119 (N_18119,N_15535,N_17340);
xnor U18120 (N_18120,N_16684,N_15858);
nand U18121 (N_18121,N_16198,N_16051);
and U18122 (N_18122,N_16840,N_15475);
nand U18123 (N_18123,N_15041,N_15932);
nor U18124 (N_18124,N_16959,N_15809);
and U18125 (N_18125,N_17253,N_17277);
or U18126 (N_18126,N_16239,N_15594);
xor U18127 (N_18127,N_15806,N_16434);
and U18128 (N_18128,N_16852,N_17248);
nand U18129 (N_18129,N_15418,N_16223);
nor U18130 (N_18130,N_16379,N_17215);
and U18131 (N_18131,N_16917,N_16835);
and U18132 (N_18132,N_17280,N_15265);
or U18133 (N_18133,N_16465,N_15746);
nor U18134 (N_18134,N_15267,N_15295);
nor U18135 (N_18135,N_16292,N_16628);
xnor U18136 (N_18136,N_15643,N_16821);
nand U18137 (N_18137,N_17138,N_15852);
xnor U18138 (N_18138,N_17359,N_15799);
and U18139 (N_18139,N_16842,N_16075);
nor U18140 (N_18140,N_16947,N_15464);
xnor U18141 (N_18141,N_15080,N_17319);
nor U18142 (N_18142,N_15923,N_16951);
or U18143 (N_18143,N_15633,N_15005);
nand U18144 (N_18144,N_17342,N_15253);
nand U18145 (N_18145,N_15862,N_16793);
and U18146 (N_18146,N_15818,N_16871);
or U18147 (N_18147,N_15429,N_17203);
nor U18148 (N_18148,N_16390,N_16567);
nand U18149 (N_18149,N_17467,N_17000);
and U18150 (N_18150,N_16590,N_16617);
nand U18151 (N_18151,N_16028,N_16007);
and U18152 (N_18152,N_16534,N_15584);
nand U18153 (N_18153,N_16202,N_17466);
or U18154 (N_18154,N_17443,N_15492);
or U18155 (N_18155,N_17363,N_15568);
nand U18156 (N_18156,N_16794,N_16846);
nand U18157 (N_18157,N_15006,N_15651);
nand U18158 (N_18158,N_16113,N_16343);
or U18159 (N_18159,N_15301,N_15826);
nor U18160 (N_18160,N_16031,N_17004);
nand U18161 (N_18161,N_15354,N_16780);
nand U18162 (N_18162,N_16053,N_16671);
xor U18163 (N_18163,N_15400,N_16256);
xnor U18164 (N_18164,N_16725,N_15373);
xnor U18165 (N_18165,N_15120,N_17141);
or U18166 (N_18166,N_17236,N_15269);
nor U18167 (N_18167,N_15939,N_15530);
nor U18168 (N_18168,N_16688,N_15333);
nand U18169 (N_18169,N_15960,N_15208);
or U18170 (N_18170,N_16573,N_15639);
nor U18171 (N_18171,N_17310,N_17413);
and U18172 (N_18172,N_16602,N_15901);
nor U18173 (N_18173,N_16691,N_15787);
nand U18174 (N_18174,N_17246,N_15950);
nor U18175 (N_18175,N_15102,N_17374);
nand U18176 (N_18176,N_15083,N_17386);
xnor U18177 (N_18177,N_16685,N_15681);
nor U18178 (N_18178,N_15013,N_16101);
nor U18179 (N_18179,N_17053,N_15853);
nand U18180 (N_18180,N_15915,N_16784);
nor U18181 (N_18181,N_15708,N_15379);
nor U18182 (N_18182,N_15204,N_16503);
nand U18183 (N_18183,N_15842,N_17195);
or U18184 (N_18184,N_17188,N_17326);
xor U18185 (N_18185,N_15558,N_15293);
nor U18186 (N_18186,N_16257,N_17136);
nand U18187 (N_18187,N_15983,N_15262);
xnor U18188 (N_18188,N_16587,N_15929);
and U18189 (N_18189,N_15959,N_16342);
nand U18190 (N_18190,N_16121,N_15951);
nor U18191 (N_18191,N_16205,N_17089);
or U18192 (N_18192,N_17135,N_15316);
nand U18193 (N_18193,N_17242,N_15797);
and U18194 (N_18194,N_17335,N_16352);
nor U18195 (N_18195,N_15532,N_16369);
nor U18196 (N_18196,N_15571,N_16072);
or U18197 (N_18197,N_16880,N_17426);
or U18198 (N_18198,N_15421,N_16032);
and U18199 (N_18199,N_17185,N_16874);
nor U18200 (N_18200,N_15397,N_15365);
or U18201 (N_18201,N_17062,N_16151);
nor U18202 (N_18202,N_16136,N_16278);
xor U18203 (N_18203,N_17231,N_15171);
nor U18204 (N_18204,N_16967,N_15133);
or U18205 (N_18205,N_16817,N_15821);
xnor U18206 (N_18206,N_15247,N_16213);
or U18207 (N_18207,N_15168,N_15998);
nor U18208 (N_18208,N_15382,N_15465);
nand U18209 (N_18209,N_17365,N_15473);
nand U18210 (N_18210,N_17083,N_16689);
nor U18211 (N_18211,N_16869,N_16855);
xnor U18212 (N_18212,N_16093,N_16412);
xnor U18213 (N_18213,N_15739,N_16920);
xnor U18214 (N_18214,N_15019,N_16134);
xor U18215 (N_18215,N_15538,N_16338);
and U18216 (N_18216,N_16605,N_15567);
nand U18217 (N_18217,N_16164,N_17452);
and U18218 (N_18218,N_17348,N_15321);
xor U18219 (N_18219,N_15612,N_15148);
nand U18220 (N_18220,N_16571,N_17312);
or U18221 (N_18221,N_15677,N_15000);
xnor U18222 (N_18222,N_17125,N_15757);
and U18223 (N_18223,N_17161,N_15848);
nor U18224 (N_18224,N_15183,N_16483);
nand U18225 (N_18225,N_17329,N_16905);
nand U18226 (N_18226,N_17429,N_15688);
nor U18227 (N_18227,N_17226,N_15296);
nand U18228 (N_18228,N_17222,N_17304);
nand U18229 (N_18229,N_16207,N_16476);
or U18230 (N_18230,N_16135,N_16965);
or U18231 (N_18231,N_16081,N_15601);
and U18232 (N_18232,N_16872,N_15899);
nor U18233 (N_18233,N_16345,N_16001);
nor U18234 (N_18234,N_17311,N_15066);
xor U18235 (N_18235,N_16226,N_16229);
nor U18236 (N_18236,N_15417,N_17317);
nand U18237 (N_18237,N_15533,N_15620);
or U18238 (N_18238,N_15260,N_16897);
nand U18239 (N_18239,N_17355,N_15327);
nor U18240 (N_18240,N_15314,N_16451);
or U18241 (N_18241,N_15374,N_15030);
xnor U18242 (N_18242,N_15865,N_17288);
and U18243 (N_18243,N_16763,N_15578);
or U18244 (N_18244,N_15994,N_15977);
or U18245 (N_18245,N_16129,N_15109);
xor U18246 (N_18246,N_15820,N_17336);
nor U18247 (N_18247,N_15010,N_16560);
and U18248 (N_18248,N_17324,N_16647);
and U18249 (N_18249,N_17159,N_15984);
and U18250 (N_18250,N_15576,N_15426);
nor U18251 (N_18251,N_15101,N_15059);
nand U18252 (N_18252,N_17264,N_16319);
xor U18253 (N_18253,N_15180,N_16591);
and U18254 (N_18254,N_16491,N_16656);
xor U18255 (N_18255,N_16912,N_16398);
or U18256 (N_18256,N_15232,N_15655);
or U18257 (N_18257,N_16933,N_15657);
and U18258 (N_18258,N_16043,N_17289);
and U18259 (N_18259,N_17120,N_16441);
or U18260 (N_18260,N_16621,N_16010);
xnor U18261 (N_18261,N_16204,N_16389);
nand U18262 (N_18262,N_15735,N_16103);
nand U18263 (N_18263,N_15305,N_16927);
nor U18264 (N_18264,N_16574,N_16666);
xor U18265 (N_18265,N_16109,N_15625);
nand U18266 (N_18266,N_16004,N_16732);
nor U18267 (N_18267,N_15561,N_17162);
nand U18268 (N_18268,N_15795,N_16187);
nand U18269 (N_18269,N_17402,N_16107);
nand U18270 (N_18270,N_16777,N_15999);
or U18271 (N_18271,N_16088,N_16673);
nor U18272 (N_18272,N_15239,N_17368);
and U18273 (N_18273,N_17234,N_16165);
or U18274 (N_18274,N_17220,N_17182);
or U18275 (N_18275,N_16499,N_15667);
and U18276 (N_18276,N_16761,N_15368);
xnor U18277 (N_18277,N_16593,N_16079);
xor U18278 (N_18278,N_17076,N_17192);
xnor U18279 (N_18279,N_16235,N_16400);
nand U18280 (N_18280,N_16523,N_15304);
or U18281 (N_18281,N_16370,N_15653);
and U18282 (N_18282,N_16055,N_17275);
nand U18283 (N_18283,N_15536,N_16236);
xnor U18284 (N_18284,N_17292,N_16100);
nor U18285 (N_18285,N_17423,N_15035);
and U18286 (N_18286,N_15883,N_15514);
nand U18287 (N_18287,N_16620,N_17088);
nand U18288 (N_18288,N_16694,N_15474);
nor U18289 (N_18289,N_16642,N_15162);
or U18290 (N_18290,N_15678,N_15249);
xnor U18291 (N_18291,N_15226,N_16166);
nor U18292 (N_18292,N_17197,N_15828);
or U18293 (N_18293,N_16061,N_17491);
or U18294 (N_18294,N_16457,N_15088);
and U18295 (N_18295,N_15052,N_15553);
nand U18296 (N_18296,N_16610,N_17131);
or U18297 (N_18297,N_16790,N_15151);
nand U18298 (N_18298,N_16888,N_16653);
and U18299 (N_18299,N_15458,N_15220);
nand U18300 (N_18300,N_16276,N_15159);
and U18301 (N_18301,N_16150,N_15334);
xnor U18302 (N_18302,N_16243,N_17084);
nand U18303 (N_18303,N_16284,N_16375);
or U18304 (N_18304,N_15011,N_17018);
and U18305 (N_18305,N_15050,N_16579);
nor U18306 (N_18306,N_17111,N_16065);
or U18307 (N_18307,N_16340,N_15827);
or U18308 (N_18308,N_16014,N_15255);
or U18309 (N_18309,N_16288,N_17247);
or U18310 (N_18310,N_16518,N_15346);
or U18311 (N_18311,N_15697,N_15967);
or U18312 (N_18312,N_16764,N_17223);
and U18313 (N_18313,N_15254,N_17240);
and U18314 (N_18314,N_17302,N_17265);
nor U18315 (N_18315,N_15033,N_15195);
xnor U18316 (N_18316,N_15864,N_16401);
nor U18317 (N_18317,N_15907,N_16832);
nand U18318 (N_18318,N_15233,N_17360);
or U18319 (N_18319,N_17051,N_16332);
nor U18320 (N_18320,N_17003,N_17425);
or U18321 (N_18321,N_16102,N_17254);
or U18322 (N_18322,N_15668,N_16601);
xnor U18323 (N_18323,N_16849,N_15717);
nand U18324 (N_18324,N_16645,N_16313);
nor U18325 (N_18325,N_16137,N_15587);
nor U18326 (N_18326,N_17178,N_16916);
and U18327 (N_18327,N_16804,N_16149);
nor U18328 (N_18328,N_15824,N_15031);
nand U18329 (N_18329,N_16336,N_15830);
nand U18330 (N_18330,N_17281,N_15635);
nand U18331 (N_18331,N_16612,N_16071);
nand U18332 (N_18332,N_16248,N_16270);
or U18333 (N_18333,N_16030,N_16635);
xor U18334 (N_18334,N_15074,N_15023);
xor U18335 (N_18335,N_16702,N_17024);
nand U18336 (N_18336,N_15348,N_15096);
or U18337 (N_18337,N_17334,N_17318);
or U18338 (N_18338,N_16382,N_16915);
xor U18339 (N_18339,N_16188,N_15559);
nand U18340 (N_18340,N_15752,N_15813);
and U18341 (N_18341,N_17189,N_15946);
or U18342 (N_18342,N_16600,N_15973);
or U18343 (N_18343,N_15954,N_16968);
and U18344 (N_18344,N_17028,N_15340);
and U18345 (N_18345,N_15673,N_16003);
nor U18346 (N_18346,N_17071,N_15176);
xor U18347 (N_18347,N_15482,N_16696);
xor U18348 (N_18348,N_17346,N_16020);
nand U18349 (N_18349,N_15420,N_17183);
xnor U18350 (N_18350,N_15086,N_15026);
or U18351 (N_18351,N_15380,N_16565);
nand U18352 (N_18352,N_16556,N_16191);
nor U18353 (N_18353,N_16015,N_16060);
xnor U18354 (N_18354,N_16245,N_17147);
nor U18355 (N_18355,N_16160,N_15798);
and U18356 (N_18356,N_15457,N_17492);
nand U18357 (N_18357,N_16791,N_16394);
or U18358 (N_18358,N_16748,N_15743);
xnor U18359 (N_18359,N_17323,N_15928);
xor U18360 (N_18360,N_15986,N_15663);
xnor U18361 (N_18361,N_16249,N_15914);
xnor U18362 (N_18362,N_16454,N_16651);
and U18363 (N_18363,N_15582,N_17347);
or U18364 (N_18364,N_16630,N_16624);
and U18365 (N_18365,N_16710,N_16041);
nand U18366 (N_18366,N_15776,N_16639);
xor U18367 (N_18367,N_16326,N_16773);
and U18368 (N_18368,N_16470,N_15198);
nor U18369 (N_18369,N_16583,N_16039);
or U18370 (N_18370,N_15363,N_15407);
xor U18371 (N_18371,N_16699,N_15211);
or U18372 (N_18372,N_16828,N_15117);
nor U18373 (N_18373,N_15472,N_15308);
and U18374 (N_18374,N_17404,N_17354);
nor U18375 (N_18375,N_15027,N_16302);
xnor U18376 (N_18376,N_15547,N_17279);
xor U18377 (N_18377,N_15520,N_17322);
nor U18378 (N_18378,N_16675,N_15991);
and U18379 (N_18379,N_15433,N_16178);
and U18380 (N_18380,N_15360,N_16633);
and U18381 (N_18381,N_17164,N_15768);
and U18382 (N_18382,N_17441,N_15870);
or U18383 (N_18383,N_15146,N_16118);
nand U18384 (N_18384,N_16508,N_16227);
and U18385 (N_18385,N_15857,N_16042);
nand U18386 (N_18386,N_17249,N_16436);
nor U18387 (N_18387,N_15958,N_16280);
nand U18388 (N_18388,N_15284,N_15131);
and U18389 (N_18389,N_16867,N_17490);
xnor U18390 (N_18390,N_17488,N_15541);
nor U18391 (N_18391,N_17338,N_17081);
and U18392 (N_18392,N_15153,N_16733);
or U18393 (N_18393,N_16488,N_15082);
or U18394 (N_18394,N_16595,N_17133);
and U18395 (N_18395,N_17214,N_17123);
and U18396 (N_18396,N_15896,N_15493);
nor U18397 (N_18397,N_16125,N_17232);
xor U18398 (N_18398,N_15721,N_15024);
and U18399 (N_18399,N_16516,N_16514);
or U18400 (N_18400,N_16809,N_15160);
xor U18401 (N_18401,N_16769,N_17306);
xnor U18402 (N_18402,N_15672,N_15442);
or U18403 (N_18403,N_16087,N_17473);
nor U18404 (N_18404,N_16812,N_16709);
xor U18405 (N_18405,N_17172,N_16632);
nor U18406 (N_18406,N_16640,N_17493);
nand U18407 (N_18407,N_16446,N_15364);
nor U18408 (N_18408,N_16681,N_17116);
xnor U18409 (N_18409,N_16350,N_16091);
nand U18410 (N_18410,N_15542,N_16594);
nor U18411 (N_18411,N_16859,N_16908);
xor U18412 (N_18412,N_16637,N_16403);
and U18413 (N_18413,N_16466,N_15356);
nand U18414 (N_18414,N_15863,N_15925);
nand U18415 (N_18415,N_15909,N_16517);
xor U18416 (N_18416,N_15926,N_15916);
xnor U18417 (N_18417,N_16695,N_15214);
and U18418 (N_18418,N_17327,N_15075);
or U18419 (N_18419,N_17068,N_16372);
or U18420 (N_18420,N_17025,N_17180);
or U18421 (N_18421,N_15669,N_15942);
and U18422 (N_18422,N_16886,N_15912);
xor U18423 (N_18423,N_17013,N_17325);
and U18424 (N_18424,N_16676,N_17461);
nor U18425 (N_18425,N_16792,N_17383);
and U18426 (N_18426,N_16746,N_15337);
or U18427 (N_18427,N_17271,N_17097);
nor U18428 (N_18428,N_16546,N_17108);
and U18429 (N_18429,N_15399,N_16473);
or U18430 (N_18430,N_16705,N_17241);
xnor U18431 (N_18431,N_17075,N_15290);
or U18432 (N_18432,N_17385,N_17458);
or U18433 (N_18433,N_17115,N_16290);
nor U18434 (N_18434,N_15216,N_16090);
or U18435 (N_18435,N_16271,N_17498);
nor U18436 (N_18436,N_16636,N_15169);
nor U18437 (N_18437,N_15694,N_16130);
nor U18438 (N_18438,N_17093,N_17433);
or U18439 (N_18439,N_15699,N_16530);
nor U18440 (N_18440,N_17127,N_16716);
xor U18441 (N_18441,N_15652,N_17140);
nor U18442 (N_18442,N_15922,N_16196);
or U18443 (N_18443,N_16289,N_15110);
nand U18444 (N_18444,N_17221,N_16611);
and U18445 (N_18445,N_17128,N_16980);
and U18446 (N_18446,N_16551,N_15422);
or U18447 (N_18447,N_17261,N_15972);
and U18448 (N_18448,N_15549,N_16783);
xor U18449 (N_18449,N_15411,N_17470);
or U18450 (N_18450,N_15720,N_16801);
xor U18451 (N_18451,N_17118,N_17339);
or U18452 (N_18452,N_15944,N_16795);
nand U18453 (N_18453,N_17379,N_16145);
and U18454 (N_18454,N_15174,N_16742);
and U18455 (N_18455,N_17029,N_15320);
and U18456 (N_18456,N_15415,N_15431);
xnor U18457 (N_18457,N_17041,N_17106);
xnor U18458 (N_18458,N_16184,N_16522);
xnor U18459 (N_18459,N_15353,N_16062);
xor U18460 (N_18460,N_17153,N_16438);
nor U18461 (N_18461,N_15758,N_15531);
nor U18462 (N_18462,N_16826,N_15895);
nand U18463 (N_18463,N_15114,N_15941);
nor U18464 (N_18464,N_15525,N_17216);
nor U18465 (N_18465,N_15351,N_16387);
or U18466 (N_18466,N_15412,N_16209);
or U18467 (N_18467,N_15659,N_16974);
or U18468 (N_18468,N_15217,N_15037);
or U18469 (N_18469,N_17437,N_15947);
nor U18470 (N_18470,N_15881,N_15517);
nor U18471 (N_18471,N_15064,N_15641);
and U18472 (N_18472,N_15127,N_16520);
and U18473 (N_18473,N_15014,N_15920);
nand U18474 (N_18474,N_16584,N_15744);
nor U18475 (N_18475,N_16942,N_16334);
and U18476 (N_18476,N_16722,N_15186);
xnor U18477 (N_18477,N_15775,N_16335);
and U18478 (N_18478,N_17194,N_16515);
or U18479 (N_18479,N_15256,N_16341);
nand U18480 (N_18480,N_15953,N_16966);
xnor U18481 (N_18481,N_16781,N_15588);
xnor U18482 (N_18482,N_15963,N_16922);
xnor U18483 (N_18483,N_16116,N_17290);
xor U18484 (N_18484,N_16189,N_16512);
or U18485 (N_18485,N_16115,N_15143);
and U18486 (N_18486,N_15283,N_16464);
xor U18487 (N_18487,N_16316,N_16818);
nor U18488 (N_18488,N_15615,N_17250);
nand U18489 (N_18489,N_15452,N_16654);
or U18490 (N_18490,N_16690,N_16331);
nand U18491 (N_18491,N_15405,N_17174);
nor U18492 (N_18492,N_17069,N_15424);
and U18493 (N_18493,N_17356,N_16944);
nand U18494 (N_18494,N_16405,N_17175);
nand U18495 (N_18495,N_15897,N_17095);
xnor U18496 (N_18496,N_16982,N_16147);
nand U18497 (N_18497,N_15544,N_16416);
nor U18498 (N_18498,N_15261,N_16376);
nor U18499 (N_18499,N_15711,N_17480);
or U18500 (N_18500,N_15931,N_15616);
and U18501 (N_18501,N_15714,N_16501);
or U18502 (N_18502,N_17352,N_15274);
nor U18503 (N_18503,N_16766,N_15384);
nor U18504 (N_18504,N_15138,N_15905);
nor U18505 (N_18505,N_16836,N_16124);
or U18506 (N_18506,N_15583,N_15618);
nor U18507 (N_18507,N_15480,N_17073);
nand U18508 (N_18508,N_15680,N_15145);
or U18509 (N_18509,N_16068,N_15936);
nor U18510 (N_18510,N_17399,N_17008);
and U18511 (N_18511,N_17210,N_16999);
and U18512 (N_18512,N_16084,N_17439);
nor U18513 (N_18513,N_16693,N_16850);
nand U18514 (N_18514,N_17187,N_17166);
nor U18515 (N_18515,N_17213,N_15637);
xnor U18516 (N_18516,N_17455,N_17350);
nor U18517 (N_18517,N_15325,N_15451);
or U18518 (N_18518,N_16388,N_16221);
nand U18519 (N_18519,N_17023,N_16344);
nand U18520 (N_18520,N_16406,N_16749);
and U18521 (N_18521,N_15355,N_15068);
nand U18522 (N_18522,N_15966,N_16181);
xnor U18523 (N_18523,N_17061,N_15585);
and U18524 (N_18524,N_17331,N_17460);
or U18525 (N_18525,N_15017,N_16541);
nand U18526 (N_18526,N_16158,N_17396);
nor U18527 (N_18527,N_15630,N_16739);
and U18528 (N_18528,N_15723,N_15352);
nand U18529 (N_18529,N_15671,N_17067);
nor U18530 (N_18530,N_15569,N_16834);
xnor U18531 (N_18531,N_15323,N_15683);
and U18532 (N_18532,N_17482,N_15859);
nand U18533 (N_18533,N_15303,N_16445);
nand U18534 (N_18534,N_17046,N_17256);
nand U18535 (N_18535,N_15189,N_15032);
and U18536 (N_18536,N_16052,N_17367);
and U18537 (N_18537,N_17444,N_15018);
nor U18538 (N_18538,N_16026,N_16495);
or U18539 (N_18539,N_16194,N_16502);
and U18540 (N_18540,N_17321,N_17478);
nand U18541 (N_18541,N_16707,N_16679);
or U18542 (N_18542,N_16543,N_15495);
nand U18543 (N_18543,N_15470,N_17065);
or U18544 (N_18544,N_15716,N_16179);
and U18545 (N_18545,N_15392,N_15500);
nor U18546 (N_18546,N_15251,N_15469);
xor U18547 (N_18547,N_17132,N_15524);
or U18548 (N_18548,N_16641,N_17427);
and U18549 (N_18549,N_17169,N_16076);
or U18550 (N_18550,N_15045,N_15390);
nor U18551 (N_18551,N_17038,N_16133);
xor U18552 (N_18552,N_15814,N_15388);
and U18553 (N_18553,N_15282,N_15841);
nand U18554 (N_18554,N_16458,N_15391);
and U18555 (N_18555,N_16771,N_15654);
xnor U18556 (N_18556,N_16127,N_15629);
nor U18557 (N_18557,N_16162,N_15483);
xor U18558 (N_18558,N_15793,N_17044);
and U18559 (N_18559,N_16106,N_16481);
and U18560 (N_18560,N_16986,N_15361);
nor U18561 (N_18561,N_15996,N_16708);
nand U18562 (N_18562,N_16669,N_16251);
xnor U18563 (N_18563,N_15961,N_15161);
and U18564 (N_18564,N_15393,N_15302);
or U18565 (N_18565,N_16228,N_16649);
and U18566 (N_18566,N_16325,N_16831);
or U18567 (N_18567,N_15992,N_17496);
nand U18568 (N_18568,N_15649,N_16987);
nor U18569 (N_18569,N_16354,N_15575);
nand U18570 (N_18570,N_16598,N_15099);
nand U18571 (N_18571,N_16402,N_16285);
xor U18572 (N_18572,N_15509,N_15835);
nor U18573 (N_18573,N_16479,N_15048);
xnor U18574 (N_18574,N_15736,N_17109);
xor U18575 (N_18575,N_17307,N_17054);
xnor U18576 (N_18576,N_15313,N_16816);
and U18577 (N_18577,N_15275,N_16455);
or U18578 (N_18578,N_15322,N_16829);
xnor U18579 (N_18579,N_15476,N_15978);
and U18580 (N_18580,N_15215,N_15557);
and U18581 (N_18581,N_17451,N_15112);
xnor U18582 (N_18582,N_15640,N_15854);
xnor U18583 (N_18583,N_16482,N_15477);
nor U18584 (N_18584,N_15646,N_17333);
nor U18585 (N_18585,N_17050,N_17382);
or U18586 (N_18586,N_15107,N_17020);
nor U18587 (N_18587,N_16608,N_15280);
xnor U18588 (N_18588,N_17112,N_16609);
nor U18589 (N_18589,N_15175,N_17411);
and U18590 (N_18590,N_16997,N_16700);
nor U18591 (N_18591,N_16385,N_16889);
nand U18592 (N_18592,N_15419,N_15596);
and U18593 (N_18593,N_15614,N_15347);
nor U18594 (N_18594,N_17031,N_16774);
and U18595 (N_18595,N_16735,N_16903);
xnor U18596 (N_18596,N_15607,N_15330);
nand U18597 (N_18597,N_15406,N_16208);
nor U18598 (N_18598,N_15632,N_17143);
or U18599 (N_18599,N_15539,N_17270);
or U18600 (N_18600,N_16924,N_16808);
xor U18601 (N_18601,N_15456,N_15523);
nor U18602 (N_18602,N_16131,N_16034);
xor U18603 (N_18603,N_17177,N_16962);
nor U18604 (N_18604,N_16806,N_16108);
and U18605 (N_18605,N_16558,N_16176);
or U18606 (N_18606,N_15206,N_15970);
nor U18607 (N_18607,N_16851,N_16077);
and U18608 (N_18608,N_15147,N_17105);
nand U18609 (N_18609,N_15856,N_15248);
nand U18610 (N_18610,N_16119,N_17100);
xnor U18611 (N_18611,N_17218,N_16919);
or U18612 (N_18612,N_17176,N_16930);
nand U18613 (N_18613,N_15512,N_15713);
nor U18614 (N_18614,N_17235,N_16110);
xnor U18615 (N_18615,N_16386,N_17349);
xnor U18616 (N_18616,N_15888,N_17079);
and U18617 (N_18617,N_15955,N_17364);
and U18618 (N_18618,N_16496,N_16770);
nor U18619 (N_18619,N_17464,N_16203);
or U18620 (N_18620,N_16064,N_16678);
nor U18621 (N_18621,N_15309,N_15815);
or U18622 (N_18622,N_15622,N_16300);
nor U18623 (N_18623,N_15372,N_17043);
nand U18624 (N_18624,N_15510,N_16638);
nor U18625 (N_18625,N_15993,N_16853);
nor U18626 (N_18626,N_17442,N_16275);
nor U18627 (N_18627,N_15115,N_15829);
or U18628 (N_18628,N_16230,N_15505);
xor U18629 (N_18629,N_15103,N_15938);
and U18630 (N_18630,N_15599,N_15890);
nand U18631 (N_18631,N_16253,N_16625);
nor U18632 (N_18632,N_16991,N_17308);
nand U18633 (N_18633,N_16566,N_15650);
and U18634 (N_18634,N_15943,N_16550);
nor U18635 (N_18635,N_15235,N_17217);
and U18636 (N_18636,N_15197,N_16359);
nor U18637 (N_18637,N_16140,N_15837);
and U18638 (N_18638,N_16755,N_15968);
nor U18639 (N_18639,N_16456,N_15335);
and U18640 (N_18640,N_16114,N_16493);
and U18641 (N_18641,N_16719,N_17126);
nand U18642 (N_18642,N_17381,N_16329);
nor U18643 (N_18643,N_16263,N_15522);
or U18644 (N_18644,N_15845,N_17421);
xnor U18645 (N_18645,N_16992,N_17072);
nand U18646 (N_18646,N_16559,N_15167);
xnor U18647 (N_18647,N_15092,N_17012);
nor U18648 (N_18648,N_15619,N_16392);
or U18649 (N_18649,N_16876,N_16768);
xor U18650 (N_18650,N_16362,N_17228);
or U18651 (N_18651,N_15749,N_17036);
xor U18652 (N_18652,N_16564,N_16526);
and U18653 (N_18653,N_15229,N_16536);
and U18654 (N_18654,N_16548,N_17353);
nand U18655 (N_18655,N_16822,N_17390);
nand U18656 (N_18656,N_15386,N_16945);
nor U18657 (N_18657,N_16282,N_17269);
nor U18658 (N_18658,N_16142,N_16827);
or U18659 (N_18659,N_15343,N_15263);
xnor U18660 (N_18660,N_17066,N_16008);
nand U18661 (N_18661,N_15889,N_17151);
nand U18662 (N_18662,N_17446,N_17291);
xor U18663 (N_18663,N_16393,N_17117);
and U18664 (N_18664,N_15310,N_15141);
or U18665 (N_18665,N_17298,N_15243);
and U18666 (N_18666,N_15194,N_16706);
and U18667 (N_18667,N_15231,N_16171);
nand U18668 (N_18668,N_15471,N_16663);
and U18669 (N_18669,N_17424,N_15142);
and U18670 (N_18670,N_17244,N_17145);
xnor U18671 (N_18671,N_16268,N_17006);
xor U18672 (N_18672,N_15756,N_16395);
nand U18673 (N_18673,N_16414,N_15178);
nor U18674 (N_18674,N_16231,N_15104);
nor U18675 (N_18675,N_15299,N_16854);
xnor U18676 (N_18676,N_15377,N_16306);
nor U18677 (N_18677,N_16440,N_15666);
and U18678 (N_18678,N_16941,N_16893);
or U18679 (N_18679,N_15144,N_17481);
and U18680 (N_18680,N_15834,N_16975);
xnor U18681 (N_18681,N_15376,N_15710);
xnor U18682 (N_18682,N_16757,N_16723);
xor U18683 (N_18683,N_17042,N_15919);
or U18684 (N_18684,N_16461,N_17431);
xor U18685 (N_18685,N_16789,N_16899);
xnor U18686 (N_18686,N_17039,N_15242);
or U18687 (N_18687,N_15962,N_16183);
and U18688 (N_18688,N_16588,N_17255);
xnor U18689 (N_18689,N_15790,N_16964);
and U18690 (N_18690,N_15927,N_15660);
nor U18691 (N_18691,N_16539,N_15843);
or U18692 (N_18692,N_15454,N_15479);
and U18693 (N_18693,N_15246,N_15071);
and U18694 (N_18694,N_16752,N_16858);
and U18695 (N_18695,N_16890,N_15908);
or U18696 (N_18696,N_15892,N_16463);
xnor U18697 (N_18697,N_17040,N_17305);
and U18698 (N_18698,N_15200,N_15580);
and U18699 (N_18699,N_16315,N_15748);
xnor U18700 (N_18700,N_16544,N_16095);
nor U18701 (N_18701,N_16711,N_15125);
nor U18702 (N_18702,N_16866,N_15940);
xnor U18703 (N_18703,N_16507,N_17208);
or U18704 (N_18704,N_17449,N_15237);
xor U18705 (N_18705,N_16910,N_15047);
and U18706 (N_18706,N_16954,N_16900);
nand U18707 (N_18707,N_16351,N_16225);
nand U18708 (N_18708,N_16011,N_15794);
and U18709 (N_18709,N_16168,N_16949);
nand U18710 (N_18710,N_16936,N_15802);
or U18711 (N_18711,N_15621,N_15590);
xnor U18712 (N_18712,N_15546,N_16805);
and U18713 (N_18713,N_15526,N_16173);
xor U18714 (N_18714,N_17328,N_15188);
xnor U18715 (N_18715,N_17262,N_15937);
xor U18716 (N_18716,N_16480,N_15503);
and U18717 (N_18717,N_16040,N_15258);
xor U18718 (N_18718,N_17102,N_15885);
and U18719 (N_18719,N_16589,N_17158);
or U18720 (N_18720,N_15761,N_16923);
nor U18721 (N_18721,N_15349,N_15855);
or U18722 (N_18722,N_16450,N_16873);
or U18723 (N_18723,N_15879,N_15498);
and U18724 (N_18724,N_15745,N_15091);
nor U18725 (N_18725,N_16692,N_15764);
or U18726 (N_18726,N_16961,N_17015);
nand U18727 (N_18727,N_16148,N_17422);
and U18728 (N_18728,N_17229,N_17077);
nor U18729 (N_18729,N_15703,N_15898);
nor U18730 (N_18730,N_16979,N_16448);
nor U18731 (N_18731,N_15664,N_16562);
xnor U18732 (N_18732,N_15706,N_16252);
nand U18733 (N_18733,N_17371,N_15497);
or U18734 (N_18734,N_16500,N_17142);
nand U18735 (N_18735,N_16569,N_15404);
nand U18736 (N_18736,N_15572,N_16492);
nor U18737 (N_18737,N_16172,N_17296);
and U18738 (N_18738,N_15801,N_15695);
or U18739 (N_18739,N_15132,N_15564);
nand U18740 (N_18740,N_17266,N_16170);
and U18741 (N_18741,N_15771,N_16175);
xor U18742 (N_18742,N_16660,N_15990);
xnor U18743 (N_18743,N_17407,N_16433);
or U18744 (N_18744,N_16471,N_15987);
or U18745 (N_18745,N_15956,N_17233);
and U18746 (N_18746,N_15868,N_16686);
or U18747 (N_18747,N_17391,N_15150);
xnor U18748 (N_18748,N_16879,N_15449);
and U18749 (N_18749,N_15438,N_16211);
nand U18750 (N_18750,N_17265,N_16482);
xor U18751 (N_18751,N_16916,N_17102);
nand U18752 (N_18752,N_17308,N_15933);
and U18753 (N_18753,N_15633,N_16760);
or U18754 (N_18754,N_15770,N_16774);
xnor U18755 (N_18755,N_16171,N_16101);
xnor U18756 (N_18756,N_16871,N_17213);
xor U18757 (N_18757,N_17169,N_15885);
and U18758 (N_18758,N_16172,N_15021);
xnor U18759 (N_18759,N_16642,N_15205);
and U18760 (N_18760,N_15035,N_15712);
nor U18761 (N_18761,N_17056,N_16918);
nor U18762 (N_18762,N_17205,N_16740);
nand U18763 (N_18763,N_15365,N_17492);
and U18764 (N_18764,N_15593,N_16819);
and U18765 (N_18765,N_15217,N_16546);
nor U18766 (N_18766,N_17176,N_17428);
nor U18767 (N_18767,N_16127,N_16088);
xnor U18768 (N_18768,N_16097,N_16909);
and U18769 (N_18769,N_17196,N_15368);
xnor U18770 (N_18770,N_16982,N_16997);
or U18771 (N_18771,N_15698,N_16358);
nor U18772 (N_18772,N_15916,N_16781);
xnor U18773 (N_18773,N_16294,N_16899);
nand U18774 (N_18774,N_16987,N_17481);
or U18775 (N_18775,N_16306,N_16126);
xor U18776 (N_18776,N_15256,N_15729);
nor U18777 (N_18777,N_15101,N_15933);
and U18778 (N_18778,N_17274,N_17242);
xor U18779 (N_18779,N_16070,N_16020);
nand U18780 (N_18780,N_17221,N_15897);
nor U18781 (N_18781,N_17009,N_15953);
nor U18782 (N_18782,N_15610,N_16836);
or U18783 (N_18783,N_16306,N_15137);
or U18784 (N_18784,N_16654,N_15200);
or U18785 (N_18785,N_16349,N_15645);
or U18786 (N_18786,N_15155,N_16451);
and U18787 (N_18787,N_16293,N_16276);
nor U18788 (N_18788,N_15400,N_16371);
xor U18789 (N_18789,N_16274,N_15813);
xor U18790 (N_18790,N_16945,N_16110);
nand U18791 (N_18791,N_16274,N_16185);
nand U18792 (N_18792,N_16511,N_15144);
xnor U18793 (N_18793,N_17064,N_17028);
and U18794 (N_18794,N_16908,N_16391);
nand U18795 (N_18795,N_17125,N_16748);
nor U18796 (N_18796,N_15261,N_16765);
nor U18797 (N_18797,N_15687,N_17278);
xnor U18798 (N_18798,N_15100,N_16578);
or U18799 (N_18799,N_17006,N_16559);
and U18800 (N_18800,N_15518,N_15211);
xnor U18801 (N_18801,N_15048,N_16272);
nor U18802 (N_18802,N_15911,N_15692);
xor U18803 (N_18803,N_17338,N_15162);
or U18804 (N_18804,N_15290,N_16688);
or U18805 (N_18805,N_15294,N_15501);
nor U18806 (N_18806,N_16462,N_15658);
nor U18807 (N_18807,N_15571,N_16958);
xnor U18808 (N_18808,N_16312,N_15069);
or U18809 (N_18809,N_15733,N_15550);
xnor U18810 (N_18810,N_17256,N_17306);
xnor U18811 (N_18811,N_15099,N_15831);
nor U18812 (N_18812,N_16864,N_15074);
nand U18813 (N_18813,N_16844,N_16239);
nand U18814 (N_18814,N_15302,N_17465);
nor U18815 (N_18815,N_16956,N_15117);
nor U18816 (N_18816,N_15790,N_15823);
nor U18817 (N_18817,N_16633,N_16257);
nand U18818 (N_18818,N_15540,N_16421);
nand U18819 (N_18819,N_16704,N_15234);
nand U18820 (N_18820,N_17383,N_15145);
xnor U18821 (N_18821,N_16174,N_16439);
xor U18822 (N_18822,N_16766,N_15529);
nand U18823 (N_18823,N_16021,N_16184);
or U18824 (N_18824,N_15196,N_16417);
nor U18825 (N_18825,N_16496,N_16731);
nand U18826 (N_18826,N_16486,N_16859);
nand U18827 (N_18827,N_15298,N_16932);
xor U18828 (N_18828,N_15426,N_16665);
or U18829 (N_18829,N_17419,N_15203);
and U18830 (N_18830,N_16533,N_15095);
nor U18831 (N_18831,N_15632,N_17439);
xnor U18832 (N_18832,N_17421,N_16711);
nand U18833 (N_18833,N_17209,N_15081);
nor U18834 (N_18834,N_16170,N_16226);
nand U18835 (N_18835,N_16761,N_15400);
or U18836 (N_18836,N_16731,N_17418);
and U18837 (N_18837,N_15454,N_16051);
and U18838 (N_18838,N_15935,N_15617);
nor U18839 (N_18839,N_16395,N_15036);
nand U18840 (N_18840,N_17498,N_15340);
xor U18841 (N_18841,N_16877,N_16851);
nor U18842 (N_18842,N_15329,N_15304);
nand U18843 (N_18843,N_15814,N_16930);
or U18844 (N_18844,N_15630,N_16827);
xor U18845 (N_18845,N_15235,N_16429);
nor U18846 (N_18846,N_16796,N_17269);
nor U18847 (N_18847,N_16533,N_16432);
xnor U18848 (N_18848,N_15239,N_15552);
nor U18849 (N_18849,N_15124,N_17248);
and U18850 (N_18850,N_16314,N_15142);
nor U18851 (N_18851,N_17319,N_17094);
nand U18852 (N_18852,N_16695,N_15709);
nor U18853 (N_18853,N_17171,N_15645);
nand U18854 (N_18854,N_16372,N_16983);
and U18855 (N_18855,N_15775,N_15207);
nor U18856 (N_18856,N_15285,N_16231);
or U18857 (N_18857,N_15902,N_16725);
or U18858 (N_18858,N_17274,N_16143);
and U18859 (N_18859,N_15925,N_17024);
xor U18860 (N_18860,N_17406,N_16842);
xnor U18861 (N_18861,N_15142,N_15516);
and U18862 (N_18862,N_16039,N_17381);
or U18863 (N_18863,N_15221,N_16896);
xnor U18864 (N_18864,N_16074,N_16984);
xnor U18865 (N_18865,N_15822,N_16931);
nand U18866 (N_18866,N_15609,N_15991);
and U18867 (N_18867,N_16797,N_15099);
and U18868 (N_18868,N_15508,N_16244);
nand U18869 (N_18869,N_16474,N_17476);
and U18870 (N_18870,N_15604,N_16916);
nor U18871 (N_18871,N_16010,N_17085);
xnor U18872 (N_18872,N_15545,N_17097);
xor U18873 (N_18873,N_15333,N_16261);
or U18874 (N_18874,N_16680,N_16181);
and U18875 (N_18875,N_17001,N_15524);
xnor U18876 (N_18876,N_17450,N_15224);
or U18877 (N_18877,N_15129,N_15647);
nand U18878 (N_18878,N_17391,N_16012);
nor U18879 (N_18879,N_15935,N_15905);
or U18880 (N_18880,N_17026,N_15783);
xnor U18881 (N_18881,N_16793,N_16895);
nor U18882 (N_18882,N_16463,N_16979);
xnor U18883 (N_18883,N_15502,N_15215);
or U18884 (N_18884,N_17424,N_15145);
nor U18885 (N_18885,N_16537,N_16016);
xor U18886 (N_18886,N_16534,N_16264);
xor U18887 (N_18887,N_16691,N_17173);
or U18888 (N_18888,N_15014,N_16538);
and U18889 (N_18889,N_15792,N_16960);
or U18890 (N_18890,N_15111,N_16721);
and U18891 (N_18891,N_15160,N_17288);
xor U18892 (N_18892,N_16406,N_15000);
or U18893 (N_18893,N_17169,N_16902);
or U18894 (N_18894,N_16508,N_17249);
or U18895 (N_18895,N_16043,N_15069);
nand U18896 (N_18896,N_15358,N_16293);
nor U18897 (N_18897,N_16103,N_17164);
nand U18898 (N_18898,N_17096,N_17194);
or U18899 (N_18899,N_15514,N_16015);
xnor U18900 (N_18900,N_16985,N_15937);
xnor U18901 (N_18901,N_17303,N_15279);
and U18902 (N_18902,N_17305,N_15978);
and U18903 (N_18903,N_17429,N_16421);
nand U18904 (N_18904,N_16679,N_16464);
nand U18905 (N_18905,N_16239,N_15897);
xor U18906 (N_18906,N_17293,N_15884);
xnor U18907 (N_18907,N_16962,N_15019);
nor U18908 (N_18908,N_15672,N_16211);
or U18909 (N_18909,N_16570,N_17160);
nand U18910 (N_18910,N_15211,N_16604);
and U18911 (N_18911,N_15685,N_15425);
nor U18912 (N_18912,N_17349,N_17000);
or U18913 (N_18913,N_16503,N_16662);
nor U18914 (N_18914,N_15418,N_16031);
nor U18915 (N_18915,N_16937,N_15245);
or U18916 (N_18916,N_15274,N_15844);
nand U18917 (N_18917,N_15912,N_15975);
and U18918 (N_18918,N_15303,N_17283);
or U18919 (N_18919,N_15155,N_17112);
xnor U18920 (N_18920,N_15943,N_16913);
xnor U18921 (N_18921,N_15238,N_17279);
nand U18922 (N_18922,N_15762,N_17250);
and U18923 (N_18923,N_17016,N_16203);
and U18924 (N_18924,N_15602,N_17351);
nor U18925 (N_18925,N_15823,N_15462);
or U18926 (N_18926,N_16675,N_16851);
xor U18927 (N_18927,N_15515,N_15476);
or U18928 (N_18928,N_15262,N_16226);
or U18929 (N_18929,N_16324,N_16887);
or U18930 (N_18930,N_17433,N_15473);
nor U18931 (N_18931,N_15555,N_16041);
nor U18932 (N_18932,N_16328,N_15523);
xnor U18933 (N_18933,N_15346,N_15369);
xnor U18934 (N_18934,N_16830,N_17249);
xnor U18935 (N_18935,N_15043,N_15083);
and U18936 (N_18936,N_15237,N_16159);
and U18937 (N_18937,N_16788,N_15252);
nor U18938 (N_18938,N_15467,N_16340);
nand U18939 (N_18939,N_16991,N_15513);
or U18940 (N_18940,N_15096,N_16854);
and U18941 (N_18941,N_16348,N_15504);
nand U18942 (N_18942,N_16924,N_17479);
nand U18943 (N_18943,N_15932,N_17113);
nand U18944 (N_18944,N_15529,N_15924);
or U18945 (N_18945,N_17373,N_15773);
nand U18946 (N_18946,N_16403,N_16736);
and U18947 (N_18947,N_16787,N_16969);
or U18948 (N_18948,N_15859,N_15966);
or U18949 (N_18949,N_15253,N_17012);
or U18950 (N_18950,N_15010,N_15286);
xor U18951 (N_18951,N_16394,N_15683);
nor U18952 (N_18952,N_16050,N_15303);
nor U18953 (N_18953,N_16110,N_15200);
or U18954 (N_18954,N_16911,N_15311);
nand U18955 (N_18955,N_16919,N_17058);
and U18956 (N_18956,N_15918,N_16017);
xor U18957 (N_18957,N_16545,N_15716);
and U18958 (N_18958,N_16617,N_17318);
xnor U18959 (N_18959,N_15822,N_15862);
nor U18960 (N_18960,N_16864,N_17183);
nand U18961 (N_18961,N_16089,N_16516);
nor U18962 (N_18962,N_16459,N_15073);
and U18963 (N_18963,N_15823,N_16198);
or U18964 (N_18964,N_15697,N_15454);
and U18965 (N_18965,N_15616,N_16459);
nand U18966 (N_18966,N_16341,N_16912);
nand U18967 (N_18967,N_16041,N_16030);
and U18968 (N_18968,N_16880,N_15818);
xor U18969 (N_18969,N_17164,N_16628);
xnor U18970 (N_18970,N_15429,N_15991);
xor U18971 (N_18971,N_15260,N_15448);
nand U18972 (N_18972,N_16662,N_17071);
xor U18973 (N_18973,N_17052,N_17407);
nor U18974 (N_18974,N_16072,N_15595);
or U18975 (N_18975,N_16407,N_15220);
and U18976 (N_18976,N_17318,N_15213);
or U18977 (N_18977,N_16595,N_15453);
nand U18978 (N_18978,N_16073,N_16776);
and U18979 (N_18979,N_15422,N_15620);
and U18980 (N_18980,N_17485,N_15562);
or U18981 (N_18981,N_16821,N_15800);
nand U18982 (N_18982,N_16127,N_16214);
xnor U18983 (N_18983,N_15500,N_16810);
nand U18984 (N_18984,N_17229,N_16222);
nand U18985 (N_18985,N_16828,N_15547);
xnor U18986 (N_18986,N_16263,N_17057);
or U18987 (N_18987,N_17371,N_15959);
or U18988 (N_18988,N_15827,N_17319);
xnor U18989 (N_18989,N_15610,N_15158);
nor U18990 (N_18990,N_16137,N_15395);
or U18991 (N_18991,N_16823,N_15379);
or U18992 (N_18992,N_15267,N_16969);
and U18993 (N_18993,N_16907,N_16371);
and U18994 (N_18994,N_15746,N_15910);
nor U18995 (N_18995,N_15829,N_16905);
xnor U18996 (N_18996,N_15975,N_15951);
xnor U18997 (N_18997,N_16516,N_16785);
xor U18998 (N_18998,N_15878,N_16560);
nor U18999 (N_18999,N_15562,N_15030);
or U19000 (N_19000,N_16728,N_16644);
or U19001 (N_19001,N_16808,N_15796);
or U19002 (N_19002,N_17303,N_16137);
nand U19003 (N_19003,N_16003,N_15830);
nand U19004 (N_19004,N_15134,N_17431);
or U19005 (N_19005,N_15662,N_15350);
nor U19006 (N_19006,N_15370,N_16563);
and U19007 (N_19007,N_15610,N_16797);
and U19008 (N_19008,N_15975,N_17019);
nor U19009 (N_19009,N_16247,N_15562);
nor U19010 (N_19010,N_17228,N_16561);
or U19011 (N_19011,N_17245,N_16091);
nand U19012 (N_19012,N_15918,N_16923);
or U19013 (N_19013,N_15351,N_15922);
nor U19014 (N_19014,N_15881,N_15257);
xnor U19015 (N_19015,N_15625,N_16641);
nor U19016 (N_19016,N_17123,N_17300);
and U19017 (N_19017,N_16336,N_15329);
or U19018 (N_19018,N_15251,N_15065);
xnor U19019 (N_19019,N_16149,N_16268);
or U19020 (N_19020,N_16548,N_15374);
xnor U19021 (N_19021,N_15952,N_17092);
nand U19022 (N_19022,N_15793,N_17185);
and U19023 (N_19023,N_16518,N_16155);
or U19024 (N_19024,N_16697,N_17252);
or U19025 (N_19025,N_16426,N_16393);
or U19026 (N_19026,N_15020,N_15521);
or U19027 (N_19027,N_15462,N_17443);
nand U19028 (N_19028,N_15057,N_16602);
or U19029 (N_19029,N_15551,N_17259);
or U19030 (N_19030,N_16039,N_16675);
or U19031 (N_19031,N_15564,N_15100);
or U19032 (N_19032,N_17319,N_17438);
nand U19033 (N_19033,N_16386,N_15383);
nand U19034 (N_19034,N_16203,N_16095);
nor U19035 (N_19035,N_15337,N_15056);
or U19036 (N_19036,N_15455,N_16406);
and U19037 (N_19037,N_15410,N_17238);
nor U19038 (N_19038,N_15177,N_15626);
and U19039 (N_19039,N_17475,N_17133);
nor U19040 (N_19040,N_16250,N_16118);
or U19041 (N_19041,N_16244,N_17098);
xnor U19042 (N_19042,N_16084,N_17462);
nand U19043 (N_19043,N_16781,N_15070);
nor U19044 (N_19044,N_16760,N_17132);
xor U19045 (N_19045,N_17083,N_15845);
or U19046 (N_19046,N_16806,N_17237);
xor U19047 (N_19047,N_16578,N_16942);
nor U19048 (N_19048,N_15008,N_17457);
xnor U19049 (N_19049,N_17315,N_15380);
xnor U19050 (N_19050,N_17246,N_15294);
xor U19051 (N_19051,N_15565,N_16203);
nand U19052 (N_19052,N_16822,N_15955);
nor U19053 (N_19053,N_15117,N_16214);
nand U19054 (N_19054,N_16556,N_16287);
nor U19055 (N_19055,N_15604,N_15935);
nand U19056 (N_19056,N_15236,N_16282);
or U19057 (N_19057,N_15577,N_17261);
nor U19058 (N_19058,N_17105,N_15402);
and U19059 (N_19059,N_15141,N_16356);
nor U19060 (N_19060,N_15980,N_15333);
xor U19061 (N_19061,N_16426,N_17013);
and U19062 (N_19062,N_16796,N_17160);
nor U19063 (N_19063,N_15874,N_16376);
and U19064 (N_19064,N_15515,N_15159);
and U19065 (N_19065,N_16275,N_16079);
nand U19066 (N_19066,N_15507,N_16269);
nor U19067 (N_19067,N_16942,N_15159);
xnor U19068 (N_19068,N_16187,N_16704);
nand U19069 (N_19069,N_15798,N_16877);
nand U19070 (N_19070,N_17464,N_15356);
xnor U19071 (N_19071,N_16365,N_16111);
nor U19072 (N_19072,N_15956,N_15233);
xor U19073 (N_19073,N_17432,N_17414);
nor U19074 (N_19074,N_17468,N_16558);
and U19075 (N_19075,N_16662,N_17093);
or U19076 (N_19076,N_15940,N_15078);
and U19077 (N_19077,N_16213,N_16650);
xnor U19078 (N_19078,N_17282,N_17020);
nor U19079 (N_19079,N_17406,N_15286);
xnor U19080 (N_19080,N_16030,N_17074);
nor U19081 (N_19081,N_15227,N_16813);
or U19082 (N_19082,N_17096,N_15753);
and U19083 (N_19083,N_16089,N_15465);
or U19084 (N_19084,N_17014,N_17388);
xor U19085 (N_19085,N_16871,N_17304);
nand U19086 (N_19086,N_15186,N_17328);
and U19087 (N_19087,N_15028,N_16651);
xnor U19088 (N_19088,N_15870,N_16369);
nand U19089 (N_19089,N_17134,N_15962);
xnor U19090 (N_19090,N_16056,N_15402);
xor U19091 (N_19091,N_16108,N_15426);
and U19092 (N_19092,N_17370,N_17091);
or U19093 (N_19093,N_15656,N_16687);
nor U19094 (N_19094,N_15644,N_16952);
or U19095 (N_19095,N_16806,N_15020);
or U19096 (N_19096,N_16572,N_17151);
nor U19097 (N_19097,N_16993,N_16534);
nand U19098 (N_19098,N_16128,N_15993);
or U19099 (N_19099,N_16722,N_15005);
and U19100 (N_19100,N_15852,N_16782);
nor U19101 (N_19101,N_15821,N_16287);
and U19102 (N_19102,N_17223,N_16407);
or U19103 (N_19103,N_16708,N_16782);
nand U19104 (N_19104,N_15947,N_16350);
nor U19105 (N_19105,N_15588,N_17051);
xor U19106 (N_19106,N_16389,N_17381);
or U19107 (N_19107,N_15555,N_16419);
nor U19108 (N_19108,N_15905,N_15321);
nor U19109 (N_19109,N_17213,N_17426);
nand U19110 (N_19110,N_16925,N_15657);
xnor U19111 (N_19111,N_17420,N_17373);
or U19112 (N_19112,N_16736,N_16874);
xor U19113 (N_19113,N_17123,N_15064);
and U19114 (N_19114,N_17431,N_15796);
and U19115 (N_19115,N_16033,N_17361);
or U19116 (N_19116,N_16076,N_15229);
or U19117 (N_19117,N_17111,N_17329);
xnor U19118 (N_19118,N_16642,N_17301);
nor U19119 (N_19119,N_16371,N_16104);
or U19120 (N_19120,N_15979,N_17144);
and U19121 (N_19121,N_15748,N_16343);
nand U19122 (N_19122,N_16664,N_17449);
nor U19123 (N_19123,N_17002,N_16131);
nand U19124 (N_19124,N_17106,N_15312);
and U19125 (N_19125,N_17110,N_16370);
nor U19126 (N_19126,N_17030,N_16080);
and U19127 (N_19127,N_15864,N_15342);
nor U19128 (N_19128,N_17481,N_17330);
and U19129 (N_19129,N_15846,N_15826);
or U19130 (N_19130,N_15562,N_15379);
or U19131 (N_19131,N_15301,N_15302);
nor U19132 (N_19132,N_16065,N_15376);
nor U19133 (N_19133,N_16018,N_16971);
and U19134 (N_19134,N_16590,N_15913);
xnor U19135 (N_19135,N_15004,N_16930);
nor U19136 (N_19136,N_16458,N_17244);
nor U19137 (N_19137,N_16147,N_17452);
xor U19138 (N_19138,N_15947,N_15463);
nand U19139 (N_19139,N_16240,N_15865);
and U19140 (N_19140,N_16327,N_17485);
or U19141 (N_19141,N_16672,N_16060);
or U19142 (N_19142,N_16793,N_15634);
nand U19143 (N_19143,N_17103,N_16918);
or U19144 (N_19144,N_15657,N_16056);
or U19145 (N_19145,N_16505,N_16223);
nor U19146 (N_19146,N_15005,N_15384);
nor U19147 (N_19147,N_15252,N_17185);
or U19148 (N_19148,N_16430,N_17110);
and U19149 (N_19149,N_16264,N_16093);
or U19150 (N_19150,N_17383,N_15308);
and U19151 (N_19151,N_17059,N_17424);
nor U19152 (N_19152,N_16615,N_16186);
nand U19153 (N_19153,N_15289,N_15699);
or U19154 (N_19154,N_16209,N_15281);
nor U19155 (N_19155,N_16555,N_17388);
nor U19156 (N_19156,N_17237,N_15924);
xor U19157 (N_19157,N_15706,N_15996);
and U19158 (N_19158,N_16486,N_15960);
or U19159 (N_19159,N_17029,N_16164);
or U19160 (N_19160,N_16596,N_16359);
and U19161 (N_19161,N_15984,N_17336);
and U19162 (N_19162,N_15619,N_16575);
xor U19163 (N_19163,N_16799,N_16147);
xor U19164 (N_19164,N_16772,N_17483);
nand U19165 (N_19165,N_17034,N_16228);
nor U19166 (N_19166,N_16167,N_15704);
or U19167 (N_19167,N_15678,N_16601);
or U19168 (N_19168,N_15516,N_16957);
nand U19169 (N_19169,N_17221,N_16915);
or U19170 (N_19170,N_15182,N_15755);
or U19171 (N_19171,N_17030,N_15249);
nor U19172 (N_19172,N_15357,N_16681);
or U19173 (N_19173,N_17201,N_17428);
and U19174 (N_19174,N_15699,N_16058);
and U19175 (N_19175,N_15870,N_16032);
and U19176 (N_19176,N_15705,N_15610);
nor U19177 (N_19177,N_16024,N_17177);
nand U19178 (N_19178,N_17054,N_17206);
nand U19179 (N_19179,N_16947,N_16177);
nand U19180 (N_19180,N_16700,N_15587);
and U19181 (N_19181,N_16738,N_16085);
xnor U19182 (N_19182,N_16911,N_15881);
nand U19183 (N_19183,N_17338,N_15890);
nor U19184 (N_19184,N_15360,N_16152);
and U19185 (N_19185,N_15589,N_16765);
or U19186 (N_19186,N_15177,N_16512);
and U19187 (N_19187,N_16541,N_15817);
nor U19188 (N_19188,N_15098,N_16165);
nand U19189 (N_19189,N_16804,N_16239);
and U19190 (N_19190,N_16084,N_16213);
xnor U19191 (N_19191,N_15196,N_15464);
nand U19192 (N_19192,N_16301,N_17196);
nand U19193 (N_19193,N_16614,N_15884);
nor U19194 (N_19194,N_17098,N_15764);
nand U19195 (N_19195,N_15609,N_17046);
nor U19196 (N_19196,N_16944,N_16114);
or U19197 (N_19197,N_17242,N_17272);
nand U19198 (N_19198,N_15795,N_15889);
nor U19199 (N_19199,N_16419,N_15590);
nand U19200 (N_19200,N_15310,N_16934);
or U19201 (N_19201,N_17387,N_17212);
or U19202 (N_19202,N_15345,N_15673);
xor U19203 (N_19203,N_15402,N_15919);
xor U19204 (N_19204,N_16640,N_15882);
or U19205 (N_19205,N_16156,N_15467);
or U19206 (N_19206,N_17391,N_15770);
nor U19207 (N_19207,N_16330,N_17059);
nor U19208 (N_19208,N_15974,N_15075);
nand U19209 (N_19209,N_15807,N_17180);
nand U19210 (N_19210,N_16101,N_15747);
or U19211 (N_19211,N_17106,N_16403);
or U19212 (N_19212,N_17003,N_17291);
nand U19213 (N_19213,N_15402,N_15716);
xor U19214 (N_19214,N_16403,N_17076);
nand U19215 (N_19215,N_16024,N_16508);
xnor U19216 (N_19216,N_15668,N_17381);
xnor U19217 (N_19217,N_17433,N_17079);
nor U19218 (N_19218,N_15259,N_15738);
nand U19219 (N_19219,N_16020,N_17005);
nand U19220 (N_19220,N_15005,N_15797);
nand U19221 (N_19221,N_15638,N_15361);
or U19222 (N_19222,N_15804,N_16687);
xor U19223 (N_19223,N_15146,N_16961);
and U19224 (N_19224,N_15546,N_17067);
or U19225 (N_19225,N_16381,N_15495);
xor U19226 (N_19226,N_17323,N_15819);
and U19227 (N_19227,N_15924,N_16439);
nand U19228 (N_19228,N_15490,N_17014);
nor U19229 (N_19229,N_15014,N_17189);
or U19230 (N_19230,N_17226,N_17313);
or U19231 (N_19231,N_15653,N_15737);
xor U19232 (N_19232,N_17283,N_16944);
and U19233 (N_19233,N_15873,N_15962);
and U19234 (N_19234,N_17321,N_15247);
xnor U19235 (N_19235,N_15634,N_17194);
or U19236 (N_19236,N_15072,N_16837);
and U19237 (N_19237,N_16945,N_15811);
or U19238 (N_19238,N_15346,N_16291);
or U19239 (N_19239,N_15306,N_16651);
xnor U19240 (N_19240,N_16753,N_15955);
xor U19241 (N_19241,N_17128,N_15973);
nor U19242 (N_19242,N_16497,N_15266);
nor U19243 (N_19243,N_15634,N_17236);
nand U19244 (N_19244,N_16112,N_16212);
nand U19245 (N_19245,N_15757,N_15347);
nand U19246 (N_19246,N_15066,N_15536);
or U19247 (N_19247,N_16224,N_15917);
or U19248 (N_19248,N_16665,N_15256);
and U19249 (N_19249,N_16586,N_15662);
and U19250 (N_19250,N_16740,N_17497);
nor U19251 (N_19251,N_15524,N_15496);
or U19252 (N_19252,N_15860,N_17270);
xor U19253 (N_19253,N_15554,N_16420);
and U19254 (N_19254,N_16439,N_15964);
and U19255 (N_19255,N_15611,N_15770);
nor U19256 (N_19256,N_15309,N_15569);
or U19257 (N_19257,N_17408,N_16303);
nand U19258 (N_19258,N_16447,N_17289);
nand U19259 (N_19259,N_17296,N_16860);
nor U19260 (N_19260,N_15350,N_17020);
xor U19261 (N_19261,N_16045,N_16007);
nor U19262 (N_19262,N_15026,N_16545);
nand U19263 (N_19263,N_16149,N_17497);
xor U19264 (N_19264,N_15164,N_16875);
and U19265 (N_19265,N_16860,N_16392);
xor U19266 (N_19266,N_15375,N_17417);
nor U19267 (N_19267,N_15001,N_16248);
nor U19268 (N_19268,N_15091,N_17168);
or U19269 (N_19269,N_16018,N_17082);
nor U19270 (N_19270,N_15085,N_17279);
or U19271 (N_19271,N_16270,N_16347);
or U19272 (N_19272,N_15957,N_15060);
nor U19273 (N_19273,N_17050,N_16777);
nor U19274 (N_19274,N_15256,N_17154);
or U19275 (N_19275,N_16323,N_16567);
nand U19276 (N_19276,N_17220,N_17354);
and U19277 (N_19277,N_15288,N_17256);
nand U19278 (N_19278,N_15510,N_16267);
and U19279 (N_19279,N_17385,N_16300);
nor U19280 (N_19280,N_16818,N_16514);
nand U19281 (N_19281,N_15454,N_17197);
and U19282 (N_19282,N_15011,N_15599);
or U19283 (N_19283,N_15157,N_16081);
nor U19284 (N_19284,N_16640,N_15788);
xnor U19285 (N_19285,N_15701,N_15822);
or U19286 (N_19286,N_16866,N_16623);
xor U19287 (N_19287,N_15464,N_15023);
xnor U19288 (N_19288,N_15623,N_16715);
xor U19289 (N_19289,N_16102,N_16263);
xor U19290 (N_19290,N_16785,N_15926);
or U19291 (N_19291,N_16183,N_16342);
and U19292 (N_19292,N_16285,N_15708);
nor U19293 (N_19293,N_16179,N_15567);
or U19294 (N_19294,N_17205,N_15856);
nand U19295 (N_19295,N_17414,N_17111);
xnor U19296 (N_19296,N_17131,N_16476);
nor U19297 (N_19297,N_15863,N_15762);
or U19298 (N_19298,N_16431,N_17131);
and U19299 (N_19299,N_16175,N_16542);
xor U19300 (N_19300,N_15252,N_15417);
xor U19301 (N_19301,N_16446,N_17054);
or U19302 (N_19302,N_15427,N_15113);
or U19303 (N_19303,N_15375,N_17010);
and U19304 (N_19304,N_17469,N_16264);
or U19305 (N_19305,N_16863,N_15442);
and U19306 (N_19306,N_15839,N_15312);
nand U19307 (N_19307,N_16780,N_17390);
nand U19308 (N_19308,N_16063,N_15428);
xnor U19309 (N_19309,N_15347,N_16664);
and U19310 (N_19310,N_16854,N_17403);
xnor U19311 (N_19311,N_17072,N_17212);
and U19312 (N_19312,N_17276,N_15314);
nand U19313 (N_19313,N_15591,N_15847);
and U19314 (N_19314,N_16730,N_16523);
nor U19315 (N_19315,N_17143,N_16582);
and U19316 (N_19316,N_17329,N_17212);
nand U19317 (N_19317,N_16051,N_16707);
nor U19318 (N_19318,N_16184,N_16257);
nand U19319 (N_19319,N_17042,N_16344);
nor U19320 (N_19320,N_16273,N_17338);
or U19321 (N_19321,N_16751,N_16075);
xnor U19322 (N_19322,N_17277,N_16212);
nand U19323 (N_19323,N_17147,N_15723);
nand U19324 (N_19324,N_15435,N_15829);
nor U19325 (N_19325,N_15857,N_15750);
nand U19326 (N_19326,N_15729,N_15686);
and U19327 (N_19327,N_15557,N_15297);
xor U19328 (N_19328,N_16554,N_15639);
xnor U19329 (N_19329,N_16541,N_15996);
and U19330 (N_19330,N_15250,N_16457);
nand U19331 (N_19331,N_15272,N_16897);
and U19332 (N_19332,N_15493,N_16592);
xnor U19333 (N_19333,N_15502,N_16102);
or U19334 (N_19334,N_17105,N_15937);
nor U19335 (N_19335,N_15582,N_16820);
nand U19336 (N_19336,N_15315,N_15159);
xor U19337 (N_19337,N_15706,N_15955);
or U19338 (N_19338,N_16641,N_16021);
xnor U19339 (N_19339,N_17141,N_16416);
nand U19340 (N_19340,N_15561,N_15109);
and U19341 (N_19341,N_16363,N_16130);
xor U19342 (N_19342,N_15839,N_15040);
nand U19343 (N_19343,N_15495,N_16637);
or U19344 (N_19344,N_16112,N_15456);
or U19345 (N_19345,N_15239,N_16899);
xnor U19346 (N_19346,N_16346,N_17008);
nand U19347 (N_19347,N_15054,N_15797);
nor U19348 (N_19348,N_16836,N_15506);
nand U19349 (N_19349,N_16169,N_16662);
nor U19350 (N_19350,N_15017,N_16685);
nand U19351 (N_19351,N_16994,N_17337);
nand U19352 (N_19352,N_17224,N_15752);
xnor U19353 (N_19353,N_16779,N_16377);
nand U19354 (N_19354,N_15302,N_15431);
or U19355 (N_19355,N_17107,N_17439);
nor U19356 (N_19356,N_17040,N_16809);
or U19357 (N_19357,N_15977,N_15723);
and U19358 (N_19358,N_15482,N_16003);
nor U19359 (N_19359,N_15019,N_15987);
and U19360 (N_19360,N_17488,N_15791);
nor U19361 (N_19361,N_15914,N_16191);
nand U19362 (N_19362,N_16145,N_16758);
nor U19363 (N_19363,N_17470,N_16673);
nor U19364 (N_19364,N_17188,N_17269);
or U19365 (N_19365,N_15529,N_17225);
nor U19366 (N_19366,N_17320,N_15660);
xor U19367 (N_19367,N_17272,N_16000);
or U19368 (N_19368,N_16914,N_16510);
and U19369 (N_19369,N_16507,N_17116);
xnor U19370 (N_19370,N_15530,N_15740);
or U19371 (N_19371,N_15132,N_16122);
nor U19372 (N_19372,N_17199,N_15582);
and U19373 (N_19373,N_15208,N_15682);
xor U19374 (N_19374,N_16256,N_17119);
nand U19375 (N_19375,N_15064,N_15303);
nor U19376 (N_19376,N_17311,N_15169);
and U19377 (N_19377,N_16175,N_17361);
and U19378 (N_19378,N_16425,N_17337);
nand U19379 (N_19379,N_17227,N_16714);
xor U19380 (N_19380,N_15990,N_16470);
nor U19381 (N_19381,N_15221,N_17009);
nor U19382 (N_19382,N_16583,N_17107);
nand U19383 (N_19383,N_15376,N_16377);
nor U19384 (N_19384,N_15433,N_15472);
nand U19385 (N_19385,N_16225,N_17032);
or U19386 (N_19386,N_16752,N_16677);
nor U19387 (N_19387,N_16046,N_16289);
nor U19388 (N_19388,N_16901,N_17107);
xnor U19389 (N_19389,N_15843,N_15689);
and U19390 (N_19390,N_15692,N_17114);
and U19391 (N_19391,N_15534,N_16481);
nand U19392 (N_19392,N_15444,N_17284);
xor U19393 (N_19393,N_16818,N_16383);
xor U19394 (N_19394,N_15818,N_16148);
or U19395 (N_19395,N_17186,N_15353);
and U19396 (N_19396,N_15930,N_15574);
nor U19397 (N_19397,N_16439,N_16729);
and U19398 (N_19398,N_15652,N_15552);
nand U19399 (N_19399,N_15427,N_16010);
or U19400 (N_19400,N_15080,N_17092);
or U19401 (N_19401,N_15934,N_16130);
and U19402 (N_19402,N_16192,N_15922);
xnor U19403 (N_19403,N_15195,N_15505);
or U19404 (N_19404,N_15203,N_15110);
nor U19405 (N_19405,N_15699,N_16302);
xor U19406 (N_19406,N_17215,N_16755);
or U19407 (N_19407,N_15068,N_16553);
and U19408 (N_19408,N_16477,N_16414);
nand U19409 (N_19409,N_15127,N_15723);
and U19410 (N_19410,N_15328,N_16703);
and U19411 (N_19411,N_16452,N_17167);
nor U19412 (N_19412,N_15788,N_17298);
xnor U19413 (N_19413,N_16089,N_17448);
or U19414 (N_19414,N_15201,N_15917);
and U19415 (N_19415,N_15631,N_16215);
xor U19416 (N_19416,N_15222,N_15592);
and U19417 (N_19417,N_15297,N_16159);
or U19418 (N_19418,N_16013,N_17403);
or U19419 (N_19419,N_17186,N_16571);
nand U19420 (N_19420,N_15869,N_17429);
nand U19421 (N_19421,N_15466,N_17440);
and U19422 (N_19422,N_16233,N_17071);
nor U19423 (N_19423,N_16284,N_17055);
nand U19424 (N_19424,N_17440,N_16627);
and U19425 (N_19425,N_15391,N_17434);
nor U19426 (N_19426,N_17380,N_16883);
or U19427 (N_19427,N_17170,N_16912);
nand U19428 (N_19428,N_15666,N_17048);
nor U19429 (N_19429,N_17041,N_15715);
or U19430 (N_19430,N_16682,N_15762);
and U19431 (N_19431,N_16425,N_15651);
or U19432 (N_19432,N_15303,N_16484);
nor U19433 (N_19433,N_15872,N_15384);
nor U19434 (N_19434,N_15757,N_17409);
nor U19435 (N_19435,N_15531,N_15056);
nor U19436 (N_19436,N_16302,N_15455);
nand U19437 (N_19437,N_15013,N_15030);
or U19438 (N_19438,N_16967,N_16355);
nor U19439 (N_19439,N_15072,N_16966);
nand U19440 (N_19440,N_16758,N_15566);
nor U19441 (N_19441,N_16092,N_16882);
or U19442 (N_19442,N_16180,N_15110);
or U19443 (N_19443,N_16743,N_15402);
nor U19444 (N_19444,N_15047,N_16232);
or U19445 (N_19445,N_15384,N_16236);
and U19446 (N_19446,N_16975,N_15743);
nor U19447 (N_19447,N_17228,N_16184);
xnor U19448 (N_19448,N_16245,N_16501);
nor U19449 (N_19449,N_17051,N_16431);
xnor U19450 (N_19450,N_17333,N_15027);
nand U19451 (N_19451,N_17456,N_15610);
nor U19452 (N_19452,N_17313,N_17456);
nor U19453 (N_19453,N_16488,N_16707);
or U19454 (N_19454,N_15562,N_17420);
and U19455 (N_19455,N_15080,N_17193);
nor U19456 (N_19456,N_17134,N_16747);
xor U19457 (N_19457,N_16714,N_15220);
and U19458 (N_19458,N_17054,N_16417);
or U19459 (N_19459,N_17251,N_17353);
or U19460 (N_19460,N_17377,N_15135);
xor U19461 (N_19461,N_16545,N_16657);
or U19462 (N_19462,N_16564,N_16901);
nand U19463 (N_19463,N_16784,N_15334);
xnor U19464 (N_19464,N_15084,N_16722);
nor U19465 (N_19465,N_16164,N_17304);
or U19466 (N_19466,N_15667,N_16138);
xor U19467 (N_19467,N_17028,N_15349);
nor U19468 (N_19468,N_15404,N_16290);
and U19469 (N_19469,N_17443,N_15124);
nor U19470 (N_19470,N_16955,N_16104);
or U19471 (N_19471,N_16140,N_16408);
nand U19472 (N_19472,N_15801,N_15450);
and U19473 (N_19473,N_15211,N_16471);
nand U19474 (N_19474,N_15310,N_16671);
xnor U19475 (N_19475,N_16159,N_15904);
and U19476 (N_19476,N_16439,N_16636);
nor U19477 (N_19477,N_16330,N_15023);
nor U19478 (N_19478,N_15323,N_17015);
and U19479 (N_19479,N_15163,N_16267);
nand U19480 (N_19480,N_16881,N_15603);
or U19481 (N_19481,N_16130,N_16649);
xnor U19482 (N_19482,N_15341,N_16687);
or U19483 (N_19483,N_16375,N_16415);
and U19484 (N_19484,N_15892,N_16508);
nand U19485 (N_19485,N_16175,N_16605);
nand U19486 (N_19486,N_17373,N_17150);
nand U19487 (N_19487,N_17139,N_15118);
or U19488 (N_19488,N_16168,N_16229);
and U19489 (N_19489,N_15094,N_16971);
and U19490 (N_19490,N_17436,N_15824);
and U19491 (N_19491,N_16491,N_16707);
and U19492 (N_19492,N_16477,N_16642);
nor U19493 (N_19493,N_16298,N_15312);
xnor U19494 (N_19494,N_16011,N_15449);
nand U19495 (N_19495,N_15492,N_15079);
or U19496 (N_19496,N_15262,N_16148);
nand U19497 (N_19497,N_15837,N_17190);
xnor U19498 (N_19498,N_16881,N_15372);
nand U19499 (N_19499,N_17157,N_16054);
and U19500 (N_19500,N_15444,N_16986);
or U19501 (N_19501,N_16371,N_17063);
xnor U19502 (N_19502,N_15663,N_15473);
nor U19503 (N_19503,N_16597,N_15916);
nand U19504 (N_19504,N_16327,N_15203);
nand U19505 (N_19505,N_16355,N_15047);
xor U19506 (N_19506,N_17156,N_15273);
nand U19507 (N_19507,N_16743,N_16752);
nor U19508 (N_19508,N_15628,N_17101);
nor U19509 (N_19509,N_15718,N_16136);
nor U19510 (N_19510,N_16199,N_17415);
or U19511 (N_19511,N_15309,N_16302);
or U19512 (N_19512,N_16961,N_17257);
xor U19513 (N_19513,N_15524,N_16091);
nor U19514 (N_19514,N_15502,N_16535);
xor U19515 (N_19515,N_17259,N_16636);
and U19516 (N_19516,N_15142,N_17226);
nor U19517 (N_19517,N_17029,N_17401);
xnor U19518 (N_19518,N_16224,N_15480);
or U19519 (N_19519,N_15060,N_16179);
xor U19520 (N_19520,N_16584,N_15665);
or U19521 (N_19521,N_16403,N_17475);
or U19522 (N_19522,N_17034,N_17326);
nand U19523 (N_19523,N_17140,N_15329);
and U19524 (N_19524,N_15118,N_17130);
and U19525 (N_19525,N_16974,N_16371);
nor U19526 (N_19526,N_15780,N_15541);
nor U19527 (N_19527,N_15147,N_15674);
nand U19528 (N_19528,N_15192,N_15646);
or U19529 (N_19529,N_15026,N_16083);
nor U19530 (N_19530,N_16760,N_16375);
nor U19531 (N_19531,N_16574,N_17498);
xor U19532 (N_19532,N_15691,N_15909);
or U19533 (N_19533,N_17177,N_16345);
nand U19534 (N_19534,N_17153,N_15265);
and U19535 (N_19535,N_15105,N_15537);
nand U19536 (N_19536,N_16781,N_16668);
nor U19537 (N_19537,N_16370,N_15668);
nand U19538 (N_19538,N_17007,N_16025);
nand U19539 (N_19539,N_15030,N_17477);
or U19540 (N_19540,N_17117,N_15340);
and U19541 (N_19541,N_17307,N_17016);
nor U19542 (N_19542,N_16922,N_16474);
xor U19543 (N_19543,N_17149,N_15626);
or U19544 (N_19544,N_16727,N_15414);
xnor U19545 (N_19545,N_17293,N_17352);
or U19546 (N_19546,N_16689,N_15043);
and U19547 (N_19547,N_17428,N_15469);
and U19548 (N_19548,N_15675,N_15279);
nand U19549 (N_19549,N_17075,N_15198);
and U19550 (N_19550,N_16057,N_16436);
or U19551 (N_19551,N_16349,N_17468);
xnor U19552 (N_19552,N_17129,N_15270);
nand U19553 (N_19553,N_15050,N_16409);
nand U19554 (N_19554,N_15785,N_16439);
nor U19555 (N_19555,N_17467,N_16805);
and U19556 (N_19556,N_16500,N_16076);
nor U19557 (N_19557,N_17105,N_16091);
or U19558 (N_19558,N_16397,N_17336);
and U19559 (N_19559,N_17374,N_17017);
or U19560 (N_19560,N_16835,N_17132);
xnor U19561 (N_19561,N_15140,N_17281);
nor U19562 (N_19562,N_16276,N_16287);
and U19563 (N_19563,N_15203,N_15039);
nor U19564 (N_19564,N_17377,N_17462);
nor U19565 (N_19565,N_17498,N_16234);
or U19566 (N_19566,N_16431,N_16508);
nor U19567 (N_19567,N_17164,N_15608);
or U19568 (N_19568,N_15600,N_15284);
xnor U19569 (N_19569,N_17483,N_16991);
nor U19570 (N_19570,N_16953,N_15140);
or U19571 (N_19571,N_15433,N_17118);
or U19572 (N_19572,N_16979,N_15026);
or U19573 (N_19573,N_17230,N_16419);
or U19574 (N_19574,N_17153,N_16127);
xor U19575 (N_19575,N_15260,N_17054);
xnor U19576 (N_19576,N_15824,N_15748);
nor U19577 (N_19577,N_15918,N_15828);
and U19578 (N_19578,N_15159,N_15083);
nand U19579 (N_19579,N_17315,N_17394);
and U19580 (N_19580,N_16329,N_16583);
or U19581 (N_19581,N_17408,N_15236);
or U19582 (N_19582,N_15837,N_16581);
nand U19583 (N_19583,N_16126,N_16550);
or U19584 (N_19584,N_16235,N_15001);
and U19585 (N_19585,N_16695,N_15921);
nand U19586 (N_19586,N_17282,N_16131);
or U19587 (N_19587,N_15286,N_16945);
and U19588 (N_19588,N_16778,N_17457);
xor U19589 (N_19589,N_16451,N_15026);
nor U19590 (N_19590,N_16801,N_15779);
nor U19591 (N_19591,N_16331,N_15815);
or U19592 (N_19592,N_17027,N_15066);
xor U19593 (N_19593,N_16576,N_16637);
or U19594 (N_19594,N_16456,N_17113);
xnor U19595 (N_19595,N_15262,N_15721);
or U19596 (N_19596,N_15901,N_16585);
and U19597 (N_19597,N_16343,N_16255);
nor U19598 (N_19598,N_16411,N_16131);
or U19599 (N_19599,N_15090,N_15570);
nand U19600 (N_19600,N_15618,N_15422);
and U19601 (N_19601,N_16591,N_17295);
xnor U19602 (N_19602,N_16023,N_16979);
and U19603 (N_19603,N_16313,N_15134);
or U19604 (N_19604,N_15208,N_16290);
nand U19605 (N_19605,N_15485,N_15945);
and U19606 (N_19606,N_16103,N_17378);
and U19607 (N_19607,N_15104,N_17394);
xnor U19608 (N_19608,N_17107,N_17185);
nor U19609 (N_19609,N_16851,N_15180);
nor U19610 (N_19610,N_15565,N_15372);
nand U19611 (N_19611,N_17401,N_15318);
nor U19612 (N_19612,N_15207,N_17101);
and U19613 (N_19613,N_15530,N_15375);
xnor U19614 (N_19614,N_16933,N_15735);
nor U19615 (N_19615,N_16604,N_16536);
and U19616 (N_19616,N_16309,N_15774);
or U19617 (N_19617,N_17071,N_16635);
or U19618 (N_19618,N_15550,N_15935);
nor U19619 (N_19619,N_15251,N_16331);
nor U19620 (N_19620,N_16863,N_17430);
nor U19621 (N_19621,N_17042,N_15460);
or U19622 (N_19622,N_15755,N_17452);
and U19623 (N_19623,N_15050,N_16314);
and U19624 (N_19624,N_17151,N_17348);
or U19625 (N_19625,N_16208,N_15904);
and U19626 (N_19626,N_15085,N_16038);
nand U19627 (N_19627,N_15333,N_17084);
and U19628 (N_19628,N_16091,N_15748);
or U19629 (N_19629,N_17234,N_15831);
nor U19630 (N_19630,N_16548,N_16235);
nand U19631 (N_19631,N_16091,N_15971);
xnor U19632 (N_19632,N_16512,N_17152);
nor U19633 (N_19633,N_15947,N_16859);
xor U19634 (N_19634,N_16524,N_16256);
nor U19635 (N_19635,N_16562,N_15522);
xnor U19636 (N_19636,N_16223,N_17175);
nand U19637 (N_19637,N_15211,N_15321);
nand U19638 (N_19638,N_16087,N_15607);
and U19639 (N_19639,N_15100,N_16889);
or U19640 (N_19640,N_15269,N_17038);
nor U19641 (N_19641,N_15888,N_16148);
and U19642 (N_19642,N_17005,N_16121);
xor U19643 (N_19643,N_15331,N_15652);
xor U19644 (N_19644,N_16118,N_17360);
xnor U19645 (N_19645,N_15296,N_15673);
xnor U19646 (N_19646,N_17031,N_16975);
nand U19647 (N_19647,N_16383,N_15310);
and U19648 (N_19648,N_16729,N_16059);
nor U19649 (N_19649,N_15364,N_16009);
or U19650 (N_19650,N_15064,N_16471);
nor U19651 (N_19651,N_16435,N_17220);
nor U19652 (N_19652,N_15172,N_15323);
and U19653 (N_19653,N_16227,N_16223);
nand U19654 (N_19654,N_17241,N_15515);
or U19655 (N_19655,N_17000,N_16903);
xnor U19656 (N_19656,N_15808,N_15825);
nor U19657 (N_19657,N_16339,N_17352);
xor U19658 (N_19658,N_17438,N_17482);
nand U19659 (N_19659,N_17088,N_16955);
nor U19660 (N_19660,N_17451,N_15625);
and U19661 (N_19661,N_15474,N_16613);
and U19662 (N_19662,N_16151,N_17371);
nor U19663 (N_19663,N_16494,N_17084);
nor U19664 (N_19664,N_15974,N_15537);
xor U19665 (N_19665,N_16366,N_16111);
and U19666 (N_19666,N_17175,N_16483);
or U19667 (N_19667,N_16270,N_17219);
xor U19668 (N_19668,N_17274,N_16401);
nor U19669 (N_19669,N_17020,N_15047);
xnor U19670 (N_19670,N_16712,N_15125);
nor U19671 (N_19671,N_15494,N_16506);
nand U19672 (N_19672,N_16190,N_16872);
or U19673 (N_19673,N_15986,N_15029);
xnor U19674 (N_19674,N_15198,N_15811);
nand U19675 (N_19675,N_16333,N_15682);
and U19676 (N_19676,N_15184,N_16677);
xor U19677 (N_19677,N_16142,N_16771);
nor U19678 (N_19678,N_15323,N_17423);
or U19679 (N_19679,N_16806,N_15826);
and U19680 (N_19680,N_17003,N_16871);
and U19681 (N_19681,N_15138,N_15800);
xnor U19682 (N_19682,N_16902,N_17029);
xor U19683 (N_19683,N_15316,N_15100);
nand U19684 (N_19684,N_15397,N_16539);
and U19685 (N_19685,N_16544,N_16891);
nand U19686 (N_19686,N_15250,N_16496);
nand U19687 (N_19687,N_16191,N_15893);
and U19688 (N_19688,N_17327,N_17213);
and U19689 (N_19689,N_15651,N_17400);
nand U19690 (N_19690,N_16631,N_15093);
and U19691 (N_19691,N_15719,N_16611);
or U19692 (N_19692,N_15407,N_15683);
nand U19693 (N_19693,N_17116,N_15875);
or U19694 (N_19694,N_16928,N_16816);
or U19695 (N_19695,N_15624,N_15254);
nor U19696 (N_19696,N_16455,N_16536);
or U19697 (N_19697,N_15395,N_15462);
or U19698 (N_19698,N_16683,N_16229);
or U19699 (N_19699,N_15592,N_15843);
or U19700 (N_19700,N_15049,N_16565);
and U19701 (N_19701,N_16794,N_16502);
or U19702 (N_19702,N_15475,N_17492);
xor U19703 (N_19703,N_17019,N_16666);
nand U19704 (N_19704,N_16334,N_16624);
or U19705 (N_19705,N_17484,N_16385);
and U19706 (N_19706,N_15549,N_15393);
xnor U19707 (N_19707,N_16229,N_17393);
nor U19708 (N_19708,N_15880,N_16402);
and U19709 (N_19709,N_15403,N_15920);
or U19710 (N_19710,N_16196,N_15978);
xnor U19711 (N_19711,N_16078,N_15412);
or U19712 (N_19712,N_15675,N_15125);
and U19713 (N_19713,N_16439,N_15907);
and U19714 (N_19714,N_17306,N_15167);
nor U19715 (N_19715,N_15967,N_17210);
nand U19716 (N_19716,N_15301,N_15838);
nand U19717 (N_19717,N_16380,N_15146);
and U19718 (N_19718,N_17189,N_15860);
xor U19719 (N_19719,N_17262,N_16240);
and U19720 (N_19720,N_16289,N_15209);
or U19721 (N_19721,N_16851,N_17230);
nand U19722 (N_19722,N_16111,N_16666);
and U19723 (N_19723,N_16455,N_16584);
and U19724 (N_19724,N_15099,N_16425);
or U19725 (N_19725,N_17324,N_16893);
xnor U19726 (N_19726,N_17154,N_16221);
nand U19727 (N_19727,N_16899,N_15446);
nor U19728 (N_19728,N_16559,N_17099);
nor U19729 (N_19729,N_16309,N_16556);
nor U19730 (N_19730,N_15732,N_17045);
and U19731 (N_19731,N_15764,N_16056);
nor U19732 (N_19732,N_16741,N_17296);
nor U19733 (N_19733,N_15821,N_16679);
nor U19734 (N_19734,N_16657,N_16779);
xnor U19735 (N_19735,N_17359,N_15895);
nor U19736 (N_19736,N_17407,N_17104);
nor U19737 (N_19737,N_17345,N_16337);
or U19738 (N_19738,N_17040,N_17029);
or U19739 (N_19739,N_15088,N_16718);
and U19740 (N_19740,N_17356,N_17436);
and U19741 (N_19741,N_15434,N_15696);
nor U19742 (N_19742,N_15690,N_15677);
nor U19743 (N_19743,N_16586,N_17055);
nand U19744 (N_19744,N_16753,N_15217);
or U19745 (N_19745,N_17154,N_15325);
nand U19746 (N_19746,N_15770,N_15382);
or U19747 (N_19747,N_15694,N_15057);
nor U19748 (N_19748,N_16556,N_16610);
or U19749 (N_19749,N_17305,N_15051);
xor U19750 (N_19750,N_17384,N_15657);
nor U19751 (N_19751,N_17018,N_16773);
and U19752 (N_19752,N_15938,N_16622);
xor U19753 (N_19753,N_15552,N_17232);
and U19754 (N_19754,N_15605,N_16413);
nor U19755 (N_19755,N_16111,N_15885);
nor U19756 (N_19756,N_16366,N_15597);
nor U19757 (N_19757,N_16003,N_15241);
and U19758 (N_19758,N_17236,N_16031);
nand U19759 (N_19759,N_16424,N_15063);
xor U19760 (N_19760,N_17227,N_15581);
xor U19761 (N_19761,N_16186,N_16257);
nor U19762 (N_19762,N_15680,N_15443);
and U19763 (N_19763,N_16742,N_16758);
or U19764 (N_19764,N_15691,N_15104);
nand U19765 (N_19765,N_16530,N_15717);
and U19766 (N_19766,N_15040,N_16523);
nand U19767 (N_19767,N_16928,N_16375);
and U19768 (N_19768,N_15248,N_16761);
and U19769 (N_19769,N_16934,N_15777);
nor U19770 (N_19770,N_15700,N_15829);
nor U19771 (N_19771,N_17150,N_17115);
nor U19772 (N_19772,N_16920,N_15755);
xor U19773 (N_19773,N_15377,N_15732);
nand U19774 (N_19774,N_16517,N_16184);
nand U19775 (N_19775,N_15146,N_17186);
xor U19776 (N_19776,N_15472,N_16093);
or U19777 (N_19777,N_17443,N_17115);
nor U19778 (N_19778,N_16721,N_16618);
or U19779 (N_19779,N_15068,N_15120);
xnor U19780 (N_19780,N_16108,N_17258);
and U19781 (N_19781,N_15745,N_15300);
nor U19782 (N_19782,N_15509,N_16091);
nand U19783 (N_19783,N_16120,N_15053);
or U19784 (N_19784,N_15685,N_15821);
nor U19785 (N_19785,N_16857,N_15822);
or U19786 (N_19786,N_17127,N_16508);
and U19787 (N_19787,N_15050,N_15750);
or U19788 (N_19788,N_16505,N_15349);
xnor U19789 (N_19789,N_15916,N_16270);
xor U19790 (N_19790,N_15071,N_17015);
or U19791 (N_19791,N_15142,N_16735);
nand U19792 (N_19792,N_15847,N_17237);
nand U19793 (N_19793,N_15298,N_15392);
and U19794 (N_19794,N_16550,N_16033);
nor U19795 (N_19795,N_16524,N_16745);
and U19796 (N_19796,N_16066,N_16974);
and U19797 (N_19797,N_15850,N_16503);
xnor U19798 (N_19798,N_15625,N_15466);
xor U19799 (N_19799,N_16281,N_17307);
nand U19800 (N_19800,N_16415,N_17250);
xor U19801 (N_19801,N_16576,N_17400);
or U19802 (N_19802,N_15813,N_16924);
and U19803 (N_19803,N_15022,N_17041);
nand U19804 (N_19804,N_17467,N_15638);
and U19805 (N_19805,N_17496,N_15416);
xor U19806 (N_19806,N_16401,N_16840);
nor U19807 (N_19807,N_16197,N_15385);
or U19808 (N_19808,N_15894,N_15386);
xnor U19809 (N_19809,N_15238,N_15770);
xnor U19810 (N_19810,N_16876,N_15412);
nand U19811 (N_19811,N_16711,N_17492);
xor U19812 (N_19812,N_17022,N_17113);
and U19813 (N_19813,N_15528,N_17288);
nor U19814 (N_19814,N_17415,N_17256);
and U19815 (N_19815,N_17275,N_16870);
and U19816 (N_19816,N_15615,N_15225);
nand U19817 (N_19817,N_16352,N_16044);
or U19818 (N_19818,N_16504,N_15753);
xnor U19819 (N_19819,N_16862,N_16306);
or U19820 (N_19820,N_16978,N_16107);
and U19821 (N_19821,N_16440,N_17263);
or U19822 (N_19822,N_15635,N_16807);
and U19823 (N_19823,N_15606,N_15892);
xor U19824 (N_19824,N_15309,N_16740);
and U19825 (N_19825,N_16705,N_15103);
nand U19826 (N_19826,N_16234,N_15193);
and U19827 (N_19827,N_15072,N_16787);
and U19828 (N_19828,N_17076,N_15924);
nor U19829 (N_19829,N_15551,N_15193);
and U19830 (N_19830,N_16090,N_17495);
or U19831 (N_19831,N_16204,N_16730);
and U19832 (N_19832,N_15645,N_16196);
or U19833 (N_19833,N_16113,N_15993);
nand U19834 (N_19834,N_17232,N_16651);
nor U19835 (N_19835,N_16814,N_17374);
xnor U19836 (N_19836,N_15066,N_15264);
xor U19837 (N_19837,N_15029,N_15889);
nand U19838 (N_19838,N_15298,N_16356);
xor U19839 (N_19839,N_16787,N_15645);
and U19840 (N_19840,N_16999,N_15300);
or U19841 (N_19841,N_15147,N_16595);
nand U19842 (N_19842,N_15967,N_16781);
and U19843 (N_19843,N_15169,N_15699);
xnor U19844 (N_19844,N_17060,N_16239);
nand U19845 (N_19845,N_15873,N_17175);
nor U19846 (N_19846,N_16513,N_15820);
nor U19847 (N_19847,N_15767,N_15309);
nand U19848 (N_19848,N_16446,N_16990);
and U19849 (N_19849,N_17304,N_17476);
and U19850 (N_19850,N_16055,N_15095);
xnor U19851 (N_19851,N_17437,N_15809);
or U19852 (N_19852,N_16403,N_16594);
nand U19853 (N_19853,N_15886,N_15265);
or U19854 (N_19854,N_15689,N_16870);
or U19855 (N_19855,N_17175,N_16433);
nor U19856 (N_19856,N_15970,N_17061);
or U19857 (N_19857,N_17165,N_17377);
or U19858 (N_19858,N_15117,N_15884);
or U19859 (N_19859,N_15272,N_15323);
or U19860 (N_19860,N_15692,N_15156);
xnor U19861 (N_19861,N_16281,N_15973);
nand U19862 (N_19862,N_15247,N_15325);
nor U19863 (N_19863,N_16664,N_15953);
nor U19864 (N_19864,N_15381,N_17172);
or U19865 (N_19865,N_16767,N_17108);
xor U19866 (N_19866,N_15730,N_15059);
and U19867 (N_19867,N_16667,N_16353);
or U19868 (N_19868,N_15766,N_15068);
xnor U19869 (N_19869,N_15055,N_16619);
xor U19870 (N_19870,N_15697,N_15789);
xnor U19871 (N_19871,N_17297,N_16408);
and U19872 (N_19872,N_17311,N_15850);
nand U19873 (N_19873,N_16141,N_16421);
and U19874 (N_19874,N_15789,N_16600);
and U19875 (N_19875,N_16314,N_16732);
nor U19876 (N_19876,N_16775,N_16779);
or U19877 (N_19877,N_17368,N_15236);
or U19878 (N_19878,N_17203,N_15735);
nor U19879 (N_19879,N_16360,N_16980);
and U19880 (N_19880,N_16421,N_17039);
and U19881 (N_19881,N_16944,N_15268);
xor U19882 (N_19882,N_16405,N_17126);
or U19883 (N_19883,N_15727,N_16662);
and U19884 (N_19884,N_15645,N_17079);
and U19885 (N_19885,N_17424,N_15703);
and U19886 (N_19886,N_16141,N_16168);
or U19887 (N_19887,N_17318,N_16172);
xor U19888 (N_19888,N_15783,N_17020);
xnor U19889 (N_19889,N_16033,N_16404);
or U19890 (N_19890,N_16818,N_15556);
nand U19891 (N_19891,N_16500,N_16762);
or U19892 (N_19892,N_16266,N_17225);
xor U19893 (N_19893,N_15303,N_16300);
xnor U19894 (N_19894,N_15110,N_16382);
nor U19895 (N_19895,N_16404,N_16468);
xnor U19896 (N_19896,N_15580,N_17057);
or U19897 (N_19897,N_16376,N_16079);
xnor U19898 (N_19898,N_17276,N_16929);
nand U19899 (N_19899,N_16105,N_15096);
and U19900 (N_19900,N_15780,N_16429);
nand U19901 (N_19901,N_15682,N_17480);
and U19902 (N_19902,N_15012,N_17302);
nor U19903 (N_19903,N_17332,N_17304);
nor U19904 (N_19904,N_15049,N_16132);
xnor U19905 (N_19905,N_15161,N_15177);
nor U19906 (N_19906,N_17242,N_16904);
or U19907 (N_19907,N_16202,N_15721);
and U19908 (N_19908,N_16090,N_15271);
nor U19909 (N_19909,N_15233,N_16232);
xor U19910 (N_19910,N_15481,N_15689);
or U19911 (N_19911,N_15265,N_16079);
and U19912 (N_19912,N_16438,N_16209);
nand U19913 (N_19913,N_15142,N_16571);
nand U19914 (N_19914,N_15320,N_16900);
or U19915 (N_19915,N_16670,N_15377);
and U19916 (N_19916,N_15151,N_15544);
xnor U19917 (N_19917,N_16110,N_16517);
and U19918 (N_19918,N_16614,N_17085);
or U19919 (N_19919,N_17140,N_16774);
or U19920 (N_19920,N_16758,N_16209);
or U19921 (N_19921,N_16880,N_17367);
nor U19922 (N_19922,N_15618,N_15295);
and U19923 (N_19923,N_15048,N_15445);
or U19924 (N_19924,N_16528,N_16142);
or U19925 (N_19925,N_17456,N_15639);
or U19926 (N_19926,N_16235,N_17042);
and U19927 (N_19927,N_16565,N_16755);
nor U19928 (N_19928,N_15746,N_17234);
xnor U19929 (N_19929,N_15742,N_16050);
and U19930 (N_19930,N_15552,N_17095);
xor U19931 (N_19931,N_15868,N_16857);
nand U19932 (N_19932,N_15184,N_15790);
and U19933 (N_19933,N_17065,N_15783);
nand U19934 (N_19934,N_15319,N_15160);
xnor U19935 (N_19935,N_15735,N_17031);
and U19936 (N_19936,N_16213,N_16205);
xor U19937 (N_19937,N_16300,N_15049);
nand U19938 (N_19938,N_16771,N_15298);
xor U19939 (N_19939,N_16014,N_16542);
and U19940 (N_19940,N_16217,N_16472);
and U19941 (N_19941,N_15383,N_16101);
and U19942 (N_19942,N_16384,N_16687);
and U19943 (N_19943,N_15603,N_17370);
and U19944 (N_19944,N_16527,N_15811);
xor U19945 (N_19945,N_15534,N_17077);
or U19946 (N_19946,N_15709,N_15177);
and U19947 (N_19947,N_17154,N_16576);
nor U19948 (N_19948,N_15614,N_15125);
and U19949 (N_19949,N_15494,N_16015);
nor U19950 (N_19950,N_16892,N_15587);
or U19951 (N_19951,N_15422,N_16604);
and U19952 (N_19952,N_17345,N_15380);
nor U19953 (N_19953,N_17398,N_15006);
nor U19954 (N_19954,N_15674,N_15208);
nand U19955 (N_19955,N_16345,N_16027);
xnor U19956 (N_19956,N_17100,N_16862);
or U19957 (N_19957,N_15276,N_16253);
nor U19958 (N_19958,N_15289,N_17110);
or U19959 (N_19959,N_16121,N_15949);
nand U19960 (N_19960,N_16600,N_15827);
nand U19961 (N_19961,N_15108,N_15805);
xor U19962 (N_19962,N_16895,N_16274);
nand U19963 (N_19963,N_17353,N_15238);
xnor U19964 (N_19964,N_16380,N_16171);
and U19965 (N_19965,N_15577,N_17455);
nor U19966 (N_19966,N_16470,N_16157);
and U19967 (N_19967,N_16784,N_16986);
or U19968 (N_19968,N_17183,N_17450);
and U19969 (N_19969,N_15056,N_16311);
and U19970 (N_19970,N_17060,N_15768);
and U19971 (N_19971,N_15831,N_15448);
and U19972 (N_19972,N_16734,N_17490);
and U19973 (N_19973,N_15591,N_15031);
nand U19974 (N_19974,N_17162,N_16044);
and U19975 (N_19975,N_17174,N_16261);
or U19976 (N_19976,N_15279,N_15833);
xor U19977 (N_19977,N_17258,N_15799);
nand U19978 (N_19978,N_17402,N_16171);
xor U19979 (N_19979,N_16305,N_17100);
nand U19980 (N_19980,N_16880,N_15439);
nand U19981 (N_19981,N_16338,N_15281);
and U19982 (N_19982,N_15879,N_16201);
nand U19983 (N_19983,N_16357,N_17072);
nor U19984 (N_19984,N_16945,N_15103);
or U19985 (N_19985,N_15611,N_15720);
xnor U19986 (N_19986,N_15659,N_17155);
nand U19987 (N_19987,N_15433,N_16474);
xor U19988 (N_19988,N_16335,N_16074);
nand U19989 (N_19989,N_15230,N_15589);
and U19990 (N_19990,N_15501,N_16785);
nand U19991 (N_19991,N_17154,N_17292);
nor U19992 (N_19992,N_16055,N_15861);
nor U19993 (N_19993,N_15640,N_17199);
nor U19994 (N_19994,N_15911,N_17373);
or U19995 (N_19995,N_17253,N_15921);
xor U19996 (N_19996,N_15496,N_17183);
nand U19997 (N_19997,N_16904,N_16076);
nor U19998 (N_19998,N_16953,N_17316);
or U19999 (N_19999,N_16920,N_16095);
or U20000 (N_20000,N_19139,N_18138);
nand U20001 (N_20001,N_18851,N_18969);
xor U20002 (N_20002,N_19166,N_19907);
xnor U20003 (N_20003,N_19651,N_18697);
or U20004 (N_20004,N_18781,N_18113);
xor U20005 (N_20005,N_18007,N_19060);
nand U20006 (N_20006,N_19583,N_19495);
nand U20007 (N_20007,N_17993,N_19592);
nor U20008 (N_20008,N_18247,N_18924);
nand U20009 (N_20009,N_17701,N_17914);
and U20010 (N_20010,N_18988,N_18661);
nor U20011 (N_20011,N_17806,N_18585);
or U20012 (N_20012,N_19349,N_19393);
and U20013 (N_20013,N_17540,N_17997);
and U20014 (N_20014,N_18572,N_18491);
nand U20015 (N_20015,N_18684,N_18885);
nor U20016 (N_20016,N_19532,N_18335);
and U20017 (N_20017,N_19229,N_18358);
nand U20018 (N_20018,N_17791,N_19730);
or U20019 (N_20019,N_18478,N_19710);
nand U20020 (N_20020,N_18529,N_19672);
nand U20021 (N_20021,N_18463,N_19786);
nand U20022 (N_20022,N_19205,N_18584);
xor U20023 (N_20023,N_17891,N_17962);
nor U20024 (N_20024,N_19752,N_18670);
or U20025 (N_20025,N_19751,N_19951);
and U20026 (N_20026,N_18418,N_19719);
xor U20027 (N_20027,N_19785,N_18811);
nor U20028 (N_20028,N_18215,N_19674);
or U20029 (N_20029,N_19222,N_19180);
nand U20030 (N_20030,N_18411,N_18373);
and U20031 (N_20031,N_19648,N_19124);
xnor U20032 (N_20032,N_17775,N_18688);
nand U20033 (N_20033,N_18231,N_17665);
nor U20034 (N_20034,N_18472,N_19377);
or U20035 (N_20035,N_19069,N_17821);
nor U20036 (N_20036,N_19714,N_19977);
and U20037 (N_20037,N_18429,N_19811);
or U20038 (N_20038,N_17835,N_19311);
or U20039 (N_20039,N_19632,N_17880);
nor U20040 (N_20040,N_18184,N_19586);
xor U20041 (N_20041,N_19999,N_17867);
xnor U20042 (N_20042,N_17520,N_18250);
nor U20043 (N_20043,N_18100,N_18590);
or U20044 (N_20044,N_17838,N_18334);
nor U20045 (N_20045,N_19019,N_19138);
nor U20046 (N_20046,N_19870,N_18467);
and U20047 (N_20047,N_18237,N_19112);
or U20048 (N_20048,N_19410,N_18962);
nor U20049 (N_20049,N_17839,N_19104);
xnor U20050 (N_20050,N_18818,N_19319);
nand U20051 (N_20051,N_18202,N_18852);
and U20052 (N_20052,N_18944,N_18689);
nand U20053 (N_20053,N_19929,N_19770);
or U20054 (N_20054,N_19483,N_19667);
nor U20055 (N_20055,N_18239,N_18181);
xor U20056 (N_20056,N_18014,N_19800);
nor U20057 (N_20057,N_18238,N_17904);
or U20058 (N_20058,N_18897,N_17535);
nand U20059 (N_20059,N_17521,N_17717);
or U20060 (N_20060,N_19150,N_19740);
xnor U20061 (N_20061,N_18667,N_19265);
nand U20062 (N_20062,N_19956,N_18768);
nand U20063 (N_20063,N_19169,N_17895);
or U20064 (N_20064,N_18639,N_18451);
nand U20065 (N_20065,N_17833,N_18991);
or U20066 (N_20066,N_18772,N_18106);
nor U20067 (N_20067,N_19781,N_17897);
xnor U20068 (N_20068,N_18120,N_18724);
nor U20069 (N_20069,N_18265,N_18864);
xnor U20070 (N_20070,N_18406,N_19245);
xor U20071 (N_20071,N_17952,N_19590);
or U20072 (N_20072,N_19942,N_19325);
and U20073 (N_20073,N_19878,N_18384);
xnor U20074 (N_20074,N_18034,N_18921);
and U20075 (N_20075,N_19728,N_19454);
or U20076 (N_20076,N_18176,N_19181);
xnor U20077 (N_20077,N_18179,N_17947);
and U20078 (N_20078,N_19986,N_18353);
and U20079 (N_20079,N_18337,N_19537);
nand U20080 (N_20080,N_17832,N_18425);
xnor U20081 (N_20081,N_18409,N_19820);
nand U20082 (N_20082,N_17888,N_18031);
or U20083 (N_20083,N_17913,N_19402);
or U20084 (N_20084,N_19877,N_18715);
nand U20085 (N_20085,N_19187,N_19436);
and U20086 (N_20086,N_17544,N_19677);
and U20087 (N_20087,N_19041,N_19481);
nand U20088 (N_20088,N_18047,N_19463);
nor U20089 (N_20089,N_17564,N_19991);
or U20090 (N_20090,N_19294,N_19054);
nor U20091 (N_20091,N_17935,N_19633);
or U20092 (N_20092,N_19178,N_17575);
nor U20093 (N_20093,N_19865,N_18342);
and U20094 (N_20094,N_19589,N_19601);
nor U20095 (N_20095,N_18344,N_18687);
xor U20096 (N_20096,N_19350,N_19538);
nand U20097 (N_20097,N_19716,N_18412);
xnor U20098 (N_20098,N_19237,N_19957);
nand U20099 (N_20099,N_18111,N_18044);
nor U20100 (N_20100,N_18055,N_17527);
or U20101 (N_20101,N_17639,N_18320);
nand U20102 (N_20102,N_18492,N_19638);
and U20103 (N_20103,N_19221,N_18038);
and U20104 (N_20104,N_19493,N_18448);
or U20105 (N_20105,N_19812,N_19827);
and U20106 (N_20106,N_19389,N_18295);
or U20107 (N_20107,N_17941,N_18980);
and U20108 (N_20108,N_18009,N_17679);
or U20109 (N_20109,N_17518,N_19539);
nor U20110 (N_20110,N_17594,N_19012);
nor U20111 (N_20111,N_19329,N_18096);
nand U20112 (N_20112,N_18499,N_19969);
and U20113 (N_20113,N_18614,N_18836);
nand U20114 (N_20114,N_19806,N_17657);
or U20115 (N_20115,N_18892,N_17814);
nand U20116 (N_20116,N_17534,N_18881);
nand U20117 (N_20117,N_19650,N_18501);
xnor U20118 (N_20118,N_19510,N_19459);
or U20119 (N_20119,N_19364,N_19433);
and U20120 (N_20120,N_17852,N_18821);
xor U20121 (N_20121,N_19765,N_19700);
and U20122 (N_20122,N_18175,N_19090);
nand U20123 (N_20123,N_17735,N_17647);
or U20124 (N_20124,N_18075,N_17558);
nand U20125 (N_20125,N_18895,N_19074);
nand U20126 (N_20126,N_19879,N_19305);
nor U20127 (N_20127,N_18975,N_19157);
and U20128 (N_20128,N_19995,N_19231);
or U20129 (N_20129,N_17848,N_19524);
or U20130 (N_20130,N_19557,N_17863);
and U20131 (N_20131,N_17680,N_17632);
xor U20132 (N_20132,N_17996,N_18999);
nand U20133 (N_20133,N_19262,N_19982);
or U20134 (N_20134,N_18720,N_19769);
nor U20135 (N_20135,N_18555,N_18681);
xnor U20136 (N_20136,N_18502,N_18475);
or U20137 (N_20137,N_18466,N_19772);
or U20138 (N_20138,N_19375,N_19232);
or U20139 (N_20139,N_17696,N_19331);
or U20140 (N_20140,N_19994,N_18006);
or U20141 (N_20141,N_18336,N_17596);
xnor U20142 (N_20142,N_18759,N_19379);
nor U20143 (N_20143,N_17536,N_17732);
and U20144 (N_20144,N_19779,N_18745);
or U20145 (N_20145,N_18274,N_17511);
nor U20146 (N_20146,N_19776,N_17514);
or U20147 (N_20147,N_18669,N_19608);
and U20148 (N_20148,N_18364,N_17936);
or U20149 (N_20149,N_19937,N_19545);
nand U20150 (N_20150,N_17506,N_18654);
and U20151 (N_20151,N_19013,N_19212);
and U20152 (N_20152,N_19475,N_17651);
nand U20153 (N_20153,N_17633,N_18310);
xnor U20154 (N_20154,N_18838,N_17650);
and U20155 (N_20155,N_19131,N_18297);
nand U20156 (N_20156,N_18622,N_19746);
xnor U20157 (N_20157,N_18432,N_18693);
and U20158 (N_20158,N_18293,N_17807);
and U20159 (N_20159,N_17840,N_18495);
or U20160 (N_20160,N_18443,N_18690);
nand U20161 (N_20161,N_19499,N_18696);
and U20162 (N_20162,N_19582,N_19300);
nand U20163 (N_20163,N_18087,N_17551);
xnor U20164 (N_20164,N_17804,N_18990);
xnor U20165 (N_20165,N_18767,N_18685);
nand U20166 (N_20166,N_18379,N_19693);
nor U20167 (N_20167,N_19189,N_18996);
xnor U20168 (N_20168,N_18504,N_18934);
xnor U20169 (N_20169,N_17720,N_18797);
nand U20170 (N_20170,N_19471,N_17513);
or U20171 (N_20171,N_19891,N_18556);
xnor U20172 (N_20172,N_19277,N_18810);
or U20173 (N_20173,N_18731,N_18882);
or U20174 (N_20174,N_18166,N_17582);
and U20175 (N_20175,N_18388,N_18997);
nor U20176 (N_20176,N_18779,N_19952);
nor U20177 (N_20177,N_19107,N_18813);
xnor U20178 (N_20178,N_19501,N_18082);
nand U20179 (N_20179,N_19466,N_19126);
nor U20180 (N_20180,N_18056,N_19861);
or U20181 (N_20181,N_17771,N_19120);
nand U20182 (N_20182,N_18800,N_19954);
xnor U20183 (N_20183,N_17860,N_18732);
and U20184 (N_20184,N_17861,N_19831);
and U20185 (N_20185,N_19488,N_19975);
or U20186 (N_20186,N_18394,N_19981);
or U20187 (N_20187,N_18780,N_17764);
nor U20188 (N_20188,N_19965,N_17757);
and U20189 (N_20189,N_18704,N_19932);
nand U20190 (N_20190,N_18444,N_17811);
nand U20191 (N_20191,N_19596,N_17773);
nand U20192 (N_20192,N_19431,N_18508);
or U20193 (N_20193,N_19449,N_17500);
nor U20194 (N_20194,N_19190,N_17682);
and U20195 (N_20195,N_19992,N_19960);
and U20196 (N_20196,N_18190,N_17963);
and U20197 (N_20197,N_18987,N_18116);
xor U20198 (N_20198,N_19563,N_19272);
nand U20199 (N_20199,N_19111,N_19269);
xnor U20200 (N_20200,N_18782,N_19233);
and U20201 (N_20201,N_19970,N_17882);
nor U20202 (N_20202,N_18099,N_17510);
and U20203 (N_20203,N_17747,N_19415);
nor U20204 (N_20204,N_17966,N_18307);
or U20205 (N_20205,N_17868,N_18363);
or U20206 (N_20206,N_19898,N_19308);
nor U20207 (N_20207,N_18544,N_18794);
or U20208 (N_20208,N_18579,N_19635);
xor U20209 (N_20209,N_18899,N_17956);
nor U20210 (N_20210,N_18597,N_17528);
and U20211 (N_20211,N_19346,N_19749);
and U20212 (N_20212,N_18553,N_18378);
nor U20213 (N_20213,N_19408,N_17587);
nand U20214 (N_20214,N_19451,N_19915);
nor U20215 (N_20215,N_18867,N_19182);
xor U20216 (N_20216,N_18018,N_19084);
nand U20217 (N_20217,N_19260,N_19892);
nand U20218 (N_20218,N_18000,N_18294);
xnor U20219 (N_20219,N_18900,N_18634);
nor U20220 (N_20220,N_18257,N_18568);
xor U20221 (N_20221,N_17601,N_18619);
and U20222 (N_20222,N_17624,N_18357);
or U20223 (N_20223,N_19526,N_19903);
or U20224 (N_20224,N_17504,N_19747);
or U20225 (N_20225,N_19142,N_19599);
nor U20226 (N_20226,N_17827,N_18527);
and U20227 (N_20227,N_17671,N_19533);
nor U20228 (N_20228,N_18906,N_18612);
nand U20229 (N_20229,N_19480,N_18855);
nor U20230 (N_20230,N_19708,N_17899);
nor U20231 (N_20231,N_17569,N_18941);
or U20232 (N_20232,N_19964,N_19924);
xor U20233 (N_20233,N_19341,N_18517);
or U20234 (N_20234,N_19902,N_19843);
or U20235 (N_20235,N_17611,N_18538);
xnor U20236 (N_20236,N_19134,N_19647);
or U20237 (N_20237,N_19679,N_18136);
nand U20238 (N_20238,N_17695,N_18386);
or U20239 (N_20239,N_18420,N_19604);
xnor U20240 (N_20240,N_19511,N_19249);
xnor U20241 (N_20241,N_18322,N_18982);
nor U20242 (N_20242,N_17925,N_18172);
nor U20243 (N_20243,N_17669,N_18230);
and U20244 (N_20244,N_19624,N_19218);
or U20245 (N_20245,N_19477,N_17825);
and U20246 (N_20246,N_19219,N_19543);
and U20247 (N_20247,N_19816,N_19479);
nor U20248 (N_20248,N_18737,N_19641);
nand U20249 (N_20249,N_18620,N_18046);
nor U20250 (N_20250,N_19010,N_19284);
nor U20251 (N_20251,N_17523,N_18316);
nor U20252 (N_20252,N_18227,N_19400);
xnor U20253 (N_20253,N_19795,N_19239);
nand U20254 (N_20254,N_18277,N_18659);
nand U20255 (N_20255,N_17922,N_17842);
or U20256 (N_20256,N_19884,N_17859);
and U20257 (N_20257,N_18383,N_17749);
xor U20258 (N_20258,N_18927,N_19860);
and U20259 (N_20259,N_19684,N_17876);
or U20260 (N_20260,N_19023,N_17593);
and U20261 (N_20261,N_18188,N_18993);
xnor U20262 (N_20262,N_19057,N_18734);
nor U20263 (N_20263,N_19984,N_18194);
or U20264 (N_20264,N_19602,N_19029);
nand U20265 (N_20265,N_19257,N_17724);
nor U20266 (N_20266,N_18677,N_19723);
and U20267 (N_20267,N_19489,N_18998);
nor U20268 (N_20268,N_18850,N_18786);
or U20269 (N_20269,N_19732,N_17627);
and U20270 (N_20270,N_18127,N_18793);
or U20271 (N_20271,N_19939,N_18091);
or U20272 (N_20272,N_19299,N_19027);
nand U20273 (N_20273,N_19047,N_19348);
xor U20274 (N_20274,N_19611,N_18380);
xnor U20275 (N_20275,N_19612,N_17585);
or U20276 (N_20276,N_19594,N_18647);
nand U20277 (N_20277,N_19922,N_18260);
xor U20278 (N_20278,N_19711,N_18566);
nor U20279 (N_20279,N_18776,N_18173);
and U20280 (N_20280,N_18936,N_19704);
nand U20281 (N_20281,N_19871,N_19911);
or U20282 (N_20282,N_19807,N_17630);
nand U20283 (N_20283,N_18147,N_18914);
or U20284 (N_20284,N_18083,N_17998);
or U20285 (N_20285,N_17945,N_17755);
or U20286 (N_20286,N_18185,N_19653);
nor U20287 (N_20287,N_18447,N_19670);
or U20288 (N_20288,N_18493,N_17649);
or U20289 (N_20289,N_18598,N_19979);
or U20290 (N_20290,N_18079,N_18796);
nor U20291 (N_20291,N_18626,N_18266);
or U20292 (N_20292,N_19976,N_18326);
nand U20293 (N_20293,N_18050,N_19031);
and U20294 (N_20294,N_19564,N_17946);
nand U20295 (N_20295,N_19804,N_19035);
nor U20296 (N_20296,N_17870,N_17855);
xor U20297 (N_20297,N_19467,N_18445);
nor U20298 (N_20298,N_18259,N_19634);
or U20299 (N_20299,N_19442,N_18558);
nor U20300 (N_20300,N_19598,N_17526);
nor U20301 (N_20301,N_19462,N_19355);
and U20302 (N_20302,N_19452,N_19154);
nand U20303 (N_20303,N_17730,N_19021);
and U20304 (N_20304,N_17708,N_19793);
and U20305 (N_20305,N_19396,N_19872);
and U20306 (N_20306,N_18905,N_19387);
nand U20307 (N_20307,N_19017,N_19369);
nand U20308 (N_20308,N_17603,N_19550);
nand U20309 (N_20309,N_17532,N_19067);
nor U20310 (N_20310,N_19314,N_18604);
nor U20311 (N_20311,N_19439,N_17815);
and U20312 (N_20312,N_19327,N_18072);
xor U20313 (N_20313,N_17616,N_18902);
xor U20314 (N_20314,N_17698,N_17589);
nor U20315 (N_20315,N_18049,N_19864);
and U20316 (N_20316,N_19874,N_19148);
and U20317 (N_20317,N_18783,N_18407);
nand U20318 (N_20318,N_18929,N_19642);
xor U20319 (N_20319,N_17769,N_19223);
and U20320 (N_20320,N_19996,N_19398);
xor U20321 (N_20321,N_18655,N_17813);
nand U20322 (N_20322,N_17509,N_19914);
and U20323 (N_20323,N_18925,N_18738);
xnor U20324 (N_20324,N_19853,N_19644);
and U20325 (N_20325,N_18153,N_19848);
nor U20326 (N_20326,N_18862,N_19159);
xor U20327 (N_20327,N_19832,N_18931);
or U20328 (N_20328,N_18649,N_18933);
and U20329 (N_20329,N_18740,N_17705);
nand U20330 (N_20330,N_19668,N_17798);
xor U20331 (N_20331,N_17722,N_17772);
nor U20332 (N_20332,N_17921,N_19630);
or U20333 (N_20333,N_19803,N_19815);
and U20334 (N_20334,N_18709,N_18304);
or U20335 (N_20335,N_18305,N_18891);
nor U20336 (N_20336,N_19141,N_17726);
and U20337 (N_20337,N_18024,N_18291);
nor U20338 (N_20338,N_18419,N_19842);
nand U20339 (N_20339,N_17553,N_18947);
nand U20340 (N_20340,N_19916,N_19328);
nor U20341 (N_20341,N_18986,N_19572);
nand U20342 (N_20342,N_19427,N_19617);
nand U20343 (N_20343,N_19102,N_19930);
or U20344 (N_20344,N_17697,N_18245);
and U20345 (N_20345,N_17971,N_19064);
xnor U20346 (N_20346,N_19568,N_18742);
nor U20347 (N_20347,N_19496,N_19628);
or U20348 (N_20348,N_19026,N_18920);
or U20349 (N_20349,N_17915,N_19565);
xor U20350 (N_20350,N_19151,N_19339);
or U20351 (N_20351,N_19130,N_17841);
and U20352 (N_20352,N_17706,N_19390);
and U20353 (N_20353,N_17955,N_19822);
or U20354 (N_20354,N_17723,N_18037);
and U20355 (N_20355,N_18702,N_17677);
and U20356 (N_20356,N_18972,N_18516);
and U20357 (N_20357,N_18828,N_18530);
nor U20358 (N_20358,N_18645,N_18002);
and U20359 (N_20359,N_17763,N_18076);
nand U20360 (N_20360,N_17887,N_19555);
nand U20361 (N_20361,N_18756,N_17664);
and U20362 (N_20362,N_19541,N_19940);
or U20363 (N_20363,N_19153,N_17940);
or U20364 (N_20364,N_17683,N_19446);
xnor U20365 (N_20365,N_17741,N_19256);
nand U20366 (N_20366,N_18424,N_18799);
or U20367 (N_20367,N_18979,N_18343);
or U20368 (N_20368,N_18030,N_17944);
nor U20369 (N_20369,N_18139,N_19040);
and U20370 (N_20370,N_19571,N_18019);
xnor U20371 (N_20371,N_18576,N_19629);
nor U20372 (N_20372,N_18701,N_17727);
nor U20373 (N_20373,N_18833,N_18118);
and U20374 (N_20374,N_18964,N_19472);
nand U20375 (N_20375,N_18122,N_18303);
nand U20376 (N_20376,N_18656,N_17533);
nor U20377 (N_20377,N_18532,N_19172);
nand U20378 (N_20378,N_19458,N_19455);
xnor U20379 (N_20379,N_18916,N_17783);
and U20380 (N_20380,N_18984,N_18052);
xnor U20381 (N_20381,N_19756,N_18888);
xnor U20382 (N_20382,N_18368,N_18637);
or U20383 (N_20383,N_18437,N_18073);
nand U20384 (N_20384,N_18801,N_18121);
and U20385 (N_20385,N_18267,N_19391);
or U20386 (N_20386,N_18423,N_19145);
and U20387 (N_20387,N_18610,N_18698);
or U20388 (N_20388,N_18108,N_17994);
nor U20389 (N_20389,N_19137,N_18819);
nor U20390 (N_20390,N_18101,N_18562);
xnor U20391 (N_20391,N_19133,N_19998);
and U20392 (N_20392,N_19213,N_17742);
nand U20393 (N_20393,N_19217,N_17767);
or U20394 (N_20394,N_18981,N_19420);
and U20395 (N_20395,N_18646,N_18137);
and U20396 (N_20396,N_19424,N_18735);
nand U20397 (N_20397,N_17902,N_18422);
and U20398 (N_20398,N_18695,N_18020);
nand U20399 (N_20399,N_19168,N_18683);
nor U20400 (N_20400,N_19609,N_19814);
nand U20401 (N_20401,N_19712,N_19661);
nand U20402 (N_20402,N_19535,N_18525);
and U20403 (N_20403,N_18351,N_19081);
nor U20404 (N_20404,N_18456,N_19173);
and U20405 (N_20405,N_19573,N_18027);
nand U20406 (N_20406,N_18365,N_19241);
nor U20407 (N_20407,N_19666,N_18376);
nor U20408 (N_20408,N_18829,N_18324);
and U20409 (N_20409,N_17907,N_17995);
nand U20410 (N_20410,N_19839,N_18890);
and U20411 (N_20411,N_19456,N_19099);
and U20412 (N_20412,N_18489,N_19063);
xor U20413 (N_20413,N_19618,N_19438);
xnor U20414 (N_20414,N_19216,N_17615);
or U20415 (N_20415,N_17610,N_19404);
xor U20416 (N_20416,N_19657,N_18170);
and U20417 (N_20417,N_18860,N_18658);
nand U20418 (N_20418,N_17824,N_18408);
and U20419 (N_20419,N_17886,N_19514);
xor U20420 (N_20420,N_18486,N_19373);
nand U20421 (N_20421,N_17605,N_19579);
nor U20422 (N_20422,N_19973,N_18029);
nor U20423 (N_20423,N_18983,N_19847);
or U20424 (N_20424,N_19506,N_17595);
nand U20425 (N_20425,N_18391,N_17794);
and U20426 (N_20426,N_19255,N_19201);
nand U20427 (N_20427,N_18884,N_18716);
nand U20428 (N_20428,N_19008,N_18948);
nor U20429 (N_20429,N_19748,N_19692);
xor U20430 (N_20430,N_18707,N_18141);
nand U20431 (N_20431,N_18651,N_17588);
nand U20432 (N_20432,N_17505,N_17927);
nor U20433 (N_20433,N_19515,N_17800);
and U20434 (N_20434,N_18323,N_18211);
xnor U20435 (N_20435,N_18097,N_19702);
or U20436 (N_20436,N_18494,N_17684);
xor U20437 (N_20437,N_19696,N_18333);
xnor U20438 (N_20438,N_17617,N_18839);
and U20439 (N_20439,N_18465,N_17954);
and U20440 (N_20440,N_17854,N_18203);
nand U20441 (N_20441,N_19904,N_18945);
nand U20442 (N_20442,N_18678,N_19253);
or U20443 (N_20443,N_19819,N_17782);
nand U20444 (N_20444,N_19323,N_18774);
nor U20445 (N_20445,N_17643,N_18816);
xnor U20446 (N_20446,N_19947,N_17933);
nor U20447 (N_20447,N_18404,N_19562);
nor U20448 (N_20448,N_19509,N_19654);
xor U20449 (N_20449,N_19695,N_19966);
nor U20450 (N_20450,N_18258,N_18569);
xor U20451 (N_20451,N_19206,N_18160);
xnor U20452 (N_20452,N_17711,N_19238);
and U20453 (N_20453,N_17721,N_17831);
nand U20454 (N_20454,N_18356,N_18275);
or U20455 (N_20455,N_19636,N_19724);
or U20456 (N_20456,N_17686,N_18795);
or U20457 (N_20457,N_17576,N_19673);
or U20458 (N_20458,N_17803,N_19614);
nand U20459 (N_20459,N_19215,N_19890);
nor U20460 (N_20460,N_18458,N_19588);
or U20461 (N_20461,N_18280,N_18727);
nor U20462 (N_20462,N_19324,N_19517);
nand U20463 (N_20463,N_19283,N_19755);
nor U20464 (N_20464,N_18961,N_18497);
or U20465 (N_20465,N_19616,N_17818);
nand U20466 (N_20466,N_17908,N_17795);
nor U20467 (N_20467,N_18802,N_19859);
xor U20468 (N_20468,N_19419,N_19108);
nor U20469 (N_20469,N_17538,N_19896);
xnor U20470 (N_20470,N_19523,N_17893);
xnor U20471 (N_20471,N_18045,N_19658);
or U20472 (N_20472,N_18086,N_17758);
xor U20473 (N_20473,N_17619,N_19336);
and U20474 (N_20474,N_19251,N_18403);
or U20475 (N_20475,N_18169,N_18146);
and U20476 (N_20476,N_17618,N_19610);
and U20477 (N_20477,N_17837,N_18736);
nor U20478 (N_20478,N_19337,N_18606);
nor U20479 (N_20479,N_17916,N_18582);
and U20480 (N_20480,N_19286,N_18325);
xnor U20481 (N_20481,N_18967,N_18417);
nor U20482 (N_20482,N_19980,N_19204);
nor U20483 (N_20483,N_19775,N_18071);
nor U20484 (N_20484,N_19113,N_18600);
or U20485 (N_20485,N_18178,N_19764);
and U20486 (N_20486,N_18381,N_18236);
nand U20487 (N_20487,N_17752,N_19018);
nand U20488 (N_20488,N_18207,N_19725);
xor U20489 (N_20489,N_18157,N_18542);
and U20490 (N_20490,N_19095,N_17728);
xnor U20491 (N_20491,N_19170,N_19797);
nor U20492 (N_20492,N_18503,N_19681);
nand U20493 (N_20493,N_19720,N_18453);
nand U20494 (N_20494,N_19773,N_19753);
xor U20495 (N_20495,N_19362,N_18570);
and U20496 (N_20496,N_18928,N_19005);
and U20497 (N_20497,N_19913,N_17612);
xnor U20498 (N_20498,N_17709,N_19050);
nand U20499 (N_20499,N_18148,N_19056);
or U20500 (N_20500,N_19068,N_19174);
and U20501 (N_20501,N_17968,N_17719);
nand U20502 (N_20502,N_18825,N_18717);
nand U20503 (N_20503,N_18095,N_17739);
nor U20504 (N_20504,N_19485,N_19745);
or U20505 (N_20505,N_17864,N_17858);
nor U20506 (N_20506,N_17550,N_18640);
or U20507 (N_20507,N_19352,N_18309);
nand U20508 (N_20508,N_17799,N_18135);
nand U20509 (N_20509,N_19025,N_18387);
xnor U20510 (N_20510,N_19392,N_19162);
xor U20511 (N_20511,N_17943,N_17761);
nand U20512 (N_20512,N_18197,N_18213);
nor U20513 (N_20513,N_18482,N_17898);
nor U20514 (N_20514,N_17953,N_19258);
nor U20515 (N_20515,N_19179,N_17743);
nor U20516 (N_20516,N_18298,N_19766);
nor U20517 (N_20517,N_19395,N_17602);
nor U20518 (N_20518,N_18588,N_17637);
or U20519 (N_20519,N_19844,N_17573);
nand U20520 (N_20520,N_17844,N_18512);
nor U20521 (N_20521,N_18565,N_18930);
or U20522 (N_20522,N_19697,N_19409);
or U20523 (N_20523,N_18995,N_19707);
or U20524 (N_20524,N_18806,N_18217);
and U20525 (N_20525,N_18515,N_18586);
nand U20526 (N_20526,N_19276,N_18041);
nor U20527 (N_20527,N_18976,N_19689);
nand U20528 (N_20528,N_19263,N_18061);
xor U20529 (N_20529,N_18468,N_19909);
nand U20530 (N_20530,N_18765,N_18533);
xor U20531 (N_20531,N_19278,N_18421);
nor U20532 (N_20532,N_18416,N_18270);
or U20533 (N_20533,N_19058,N_19288);
and U20534 (N_20534,N_18222,N_19492);
xor U20535 (N_20535,N_18665,N_18522);
and U20536 (N_20536,N_19910,N_18674);
nand U20537 (N_20537,N_18873,N_19821);
or U20538 (N_20538,N_18865,N_18908);
or U20539 (N_20539,N_18105,N_19705);
nand U20540 (N_20540,N_18399,N_18926);
nor U20541 (N_20541,N_18165,N_17760);
or U20542 (N_20542,N_18395,N_18957);
and U20543 (N_20543,N_19437,N_17568);
xnor U20544 (N_20544,N_18474,N_19825);
and U20545 (N_20545,N_18744,N_19291);
or U20546 (N_20546,N_17592,N_17985);
nand U20547 (N_20547,N_19421,N_17851);
nand U20548 (N_20548,N_19273,N_19354);
and U20549 (N_20549,N_18263,N_19576);
nor U20550 (N_20550,N_19198,N_18537);
nor U20551 (N_20551,N_17972,N_18278);
and U20552 (N_20552,N_18487,N_18591);
and U20553 (N_20553,N_17759,N_19518);
and U20554 (N_20554,N_18439,N_19962);
xnor U20555 (N_20555,N_19771,N_18452);
nor U20556 (N_20556,N_19663,N_18712);
nand U20557 (N_20557,N_19385,N_18753);
xnor U20558 (N_20558,N_17516,N_18354);
nor U20559 (N_20559,N_18971,N_18163);
or U20560 (N_20560,N_17675,N_18535);
or U20561 (N_20561,N_19188,N_18382);
nor U20562 (N_20562,N_18286,N_17857);
xor U20563 (N_20563,N_18159,N_18460);
and U20564 (N_20564,N_19655,N_18193);
or U20565 (N_20565,N_17912,N_18663);
nand U20566 (N_20566,N_17889,N_18161);
nor U20567 (N_20567,N_18235,N_19580);
nor U20568 (N_20568,N_19155,N_17625);
nor U20569 (N_20569,N_18151,N_17905);
or U20570 (N_20570,N_17552,N_19270);
nor U20571 (N_20571,N_18594,N_19944);
xor U20572 (N_20572,N_18123,N_18104);
and U20573 (N_20573,N_18226,N_18077);
or U20574 (N_20574,N_17812,N_19567);
nand U20575 (N_20575,N_18048,N_18638);
nand U20576 (N_20576,N_19334,N_18396);
xnor U20577 (N_20577,N_18923,N_18229);
or U20578 (N_20578,N_17901,N_19465);
xnor U20579 (N_20579,N_19297,N_17676);
or U20580 (N_20580,N_17978,N_17571);
nor U20581 (N_20581,N_17746,N_17903);
xnor U20582 (N_20582,N_19993,N_17961);
or U20583 (N_20583,N_19729,N_18004);
nand U20584 (N_20584,N_19744,N_18345);
or U20585 (N_20585,N_19326,N_18608);
or U20586 (N_20586,N_18630,N_17980);
xnor U20587 (N_20587,N_17938,N_19742);
or U20588 (N_20588,N_19378,N_17733);
and U20589 (N_20589,N_17744,N_17776);
or U20590 (N_20590,N_18671,N_19316);
or U20591 (N_20591,N_19837,N_17975);
and U20592 (N_20592,N_17930,N_19279);
and U20593 (N_20593,N_19382,N_19988);
xor U20594 (N_20594,N_19484,N_19443);
nand U20595 (N_20595,N_19768,N_18033);
nand U20596 (N_20596,N_17729,N_19955);
xor U20597 (N_20597,N_18743,N_18904);
or U20598 (N_20598,N_19282,N_19220);
nor U20599 (N_20599,N_18283,N_19250);
nor U20600 (N_20600,N_19246,N_17873);
nand U20601 (N_20601,N_19071,N_19912);
nor U20602 (N_20602,N_19280,N_18546);
nor U20603 (N_20603,N_18605,N_18893);
or U20604 (N_20604,N_18150,N_18787);
and U20605 (N_20605,N_18506,N_19889);
nand U20606 (N_20606,N_19358,N_17700);
xor U20607 (N_20607,N_17622,N_18015);
xnor U20608 (N_20608,N_18549,N_18167);
nand U20609 (N_20609,N_18431,N_17574);
or U20610 (N_20610,N_17879,N_17856);
nor U20611 (N_20611,N_18329,N_18602);
or U20612 (N_20612,N_19195,N_17638);
nor U20613 (N_20613,N_19440,N_17648);
or U20614 (N_20614,N_19214,N_17929);
nor U20615 (N_20615,N_19504,N_19403);
xor U20616 (N_20616,N_18672,N_18832);
or U20617 (N_20617,N_19548,N_19838);
or U20618 (N_20618,N_18869,N_18158);
or U20619 (N_20619,N_19461,N_18090);
xor U20620 (N_20620,N_17658,N_19422);
and U20621 (N_20621,N_18628,N_17502);
and U20622 (N_20622,N_19900,N_19801);
and U20623 (N_20623,N_18223,N_17939);
or U20624 (N_20624,N_17614,N_18994);
xor U20625 (N_20625,N_19123,N_17718);
or U20626 (N_20626,N_19149,N_18911);
or U20627 (N_20627,N_18093,N_18221);
or U20628 (N_20628,N_18450,N_17539);
nor U20629 (N_20629,N_18039,N_19886);
or U20630 (N_20630,N_18843,N_17693);
nor U20631 (N_20631,N_17987,N_17805);
or U20632 (N_20632,N_18524,N_19925);
nor U20633 (N_20633,N_19474,N_18632);
xnor U20634 (N_20634,N_19669,N_17928);
and U20635 (N_20635,N_18571,N_18523);
xor U20636 (N_20636,N_17584,N_19826);
and U20637 (N_20637,N_17607,N_19317);
or U20638 (N_20638,N_18583,N_19863);
or U20639 (N_20639,N_18498,N_19209);
nor U20640 (N_20640,N_19428,N_19109);
xnor U20641 (N_20641,N_19866,N_18228);
xnor U20642 (N_20642,N_17716,N_19678);
nor U20643 (N_20643,N_18279,N_19927);
xnor U20644 (N_20644,N_18011,N_18328);
or U20645 (N_20645,N_19507,N_19303);
xnor U20646 (N_20646,N_18708,N_18866);
or U20647 (N_20647,N_19384,N_17923);
nand U20648 (N_20648,N_17517,N_19619);
and U20649 (N_20649,N_18617,N_19649);
or U20650 (N_20650,N_19132,N_19353);
xor U20651 (N_20651,N_19478,N_19167);
nor U20652 (N_20652,N_18918,N_18301);
nand U20653 (N_20653,N_18346,N_19743);
nand U20654 (N_20654,N_19321,N_19491);
nand U20655 (N_20655,N_19805,N_18218);
xor U20656 (N_20656,N_18730,N_18664);
nand U20657 (N_20657,N_17885,N_17846);
and U20658 (N_20658,N_17692,N_18392);
xor U20659 (N_20659,N_19600,N_19052);
xor U20660 (N_20660,N_19085,N_19397);
xnor U20661 (N_20661,N_19252,N_19121);
or U20662 (N_20662,N_19858,N_18454);
nand U20663 (N_20663,N_18629,N_19709);
nand U20664 (N_20664,N_18385,N_19399);
nor U20665 (N_20665,N_19470,N_19577);
nand U20666 (N_20666,N_17754,N_18191);
or U20667 (N_20667,N_18718,N_19553);
nand U20668 (N_20668,N_18773,N_19062);
and U20669 (N_20669,N_19505,N_18350);
and U20670 (N_20670,N_18713,N_18854);
or U20671 (N_20671,N_18642,N_19591);
or U20672 (N_20672,N_18935,N_18909);
nor U20673 (N_20673,N_19365,N_18204);
xnor U20674 (N_20674,N_19103,N_19236);
nand U20675 (N_20675,N_17642,N_17640);
and U20676 (N_20676,N_19468,N_18288);
xor U20677 (N_20677,N_18434,N_19376);
and U20678 (N_20678,N_18240,N_19224);
nor U20679 (N_20679,N_18254,N_17653);
or U20680 (N_20680,N_18074,N_18970);
nand U20681 (N_20681,N_18341,N_17817);
and U20682 (N_20682,N_18607,N_19156);
or U20683 (N_20683,N_19098,N_19441);
nor U20684 (N_20684,N_17756,N_19038);
nand U20685 (N_20685,N_17557,N_18886);
or U20686 (N_20686,N_19028,N_17519);
or U20687 (N_20687,N_18192,N_19762);
xnor U20688 (N_20688,N_19597,N_18081);
nand U20689 (N_20689,N_18815,N_18130);
or U20690 (N_20690,N_19953,N_19417);
or U20691 (N_20691,N_19578,N_18282);
nand U20692 (N_20692,N_19401,N_19758);
or U20693 (N_20693,N_18728,N_17969);
nor U20694 (N_20694,N_19868,N_18917);
xor U20695 (N_20695,N_18248,N_19799);
nor U20696 (N_20696,N_18511,N_18155);
or U20697 (N_20697,N_18117,N_18949);
and U20698 (N_20698,N_19144,N_19645);
nor U20699 (N_20699,N_18901,N_19033);
nor U20700 (N_20700,N_18053,N_17865);
xnor U20701 (N_20701,N_17786,N_17964);
and U20702 (N_20702,N_19841,N_17577);
nand U20703 (N_20703,N_17820,N_19185);
or U20704 (N_20704,N_19014,N_18859);
nor U20705 (N_20705,N_19091,N_19881);
or U20706 (N_20706,N_17570,N_18317);
or U20707 (N_20707,N_17667,N_17790);
nand U20708 (N_20708,N_19360,N_18748);
xnor U20709 (N_20709,N_19032,N_18820);
nor U20710 (N_20710,N_17977,N_18940);
nand U20711 (N_20711,N_19734,N_19593);
or U20712 (N_20712,N_19007,N_19100);
or U20713 (N_20713,N_19367,N_18128);
xnor U20714 (N_20714,N_17656,N_18413);
nand U20715 (N_20715,N_18846,N_19070);
nand U20716 (N_20716,N_18861,N_18131);
xnor U20717 (N_20717,N_18256,N_18433);
xor U20718 (N_20718,N_18789,N_18518);
nand U20719 (N_20719,N_18114,N_19818);
nand U20720 (N_20720,N_17565,N_18311);
or U20721 (N_20721,N_17566,N_18863);
nor U20722 (N_20722,N_17715,N_18164);
nand U20723 (N_20723,N_19552,N_17714);
nand U20724 (N_20724,N_19426,N_19834);
nor U20725 (N_20725,N_19363,N_19694);
and U20726 (N_20726,N_18574,N_18415);
nor U20727 (N_20727,N_18932,N_17801);
xnor U20728 (N_20728,N_18599,N_17973);
or U20729 (N_20729,N_19351,N_18960);
xor U20730 (N_20730,N_19603,N_18809);
or U20731 (N_20731,N_19830,N_17770);
nor U20732 (N_20732,N_19897,N_19244);
and U20733 (N_20733,N_18631,N_18913);
xnor U20734 (N_20734,N_19024,N_19383);
xor U20735 (N_20735,N_17542,N_18872);
xor U20736 (N_20736,N_19450,N_18390);
and U20737 (N_20737,N_19464,N_17670);
xnor U20738 (N_20738,N_17515,N_18374);
nor U20739 (N_20739,N_17869,N_17606);
xnor U20740 (N_20740,N_19796,N_19503);
or U20741 (N_20741,N_19356,N_18946);
nand U20742 (N_20742,N_18561,N_18243);
nand U20743 (N_20743,N_17674,N_19094);
xnor U20744 (N_20744,N_18253,N_19931);
or U20745 (N_20745,N_19357,N_18306);
nor U20746 (N_20746,N_17849,N_18220);
xor U20747 (N_20747,N_18627,N_19368);
and U20748 (N_20748,N_17554,N_19682);
nor U20749 (N_20749,N_18719,N_18234);
xor U20750 (N_20750,N_17545,N_18847);
or U20751 (N_20751,N_18224,N_19715);
nor U20752 (N_20752,N_19546,N_19048);
xor U20753 (N_20753,N_19075,N_18679);
xnor U20754 (N_20754,N_17668,N_18261);
and U20755 (N_20755,N_19307,N_18623);
or U20756 (N_20756,N_19974,N_18741);
nand U20757 (N_20757,N_19445,N_17850);
xor U20758 (N_20758,N_17979,N_19880);
xor U20759 (N_20759,N_19225,N_17703);
xor U20760 (N_20760,N_18042,N_19022);
xor U20761 (N_20761,N_18302,N_18367);
nand U20762 (N_20762,N_19767,N_19152);
xor U20763 (N_20763,N_18308,N_17789);
nand U20764 (N_20764,N_18577,N_18963);
nand U20765 (N_20765,N_19338,N_19574);
and U20766 (N_20766,N_17866,N_18563);
xor U20767 (N_20767,N_18296,N_18775);
and U20768 (N_20768,N_17762,N_17646);
and U20769 (N_20769,N_17591,N_18401);
or U20770 (N_20770,N_17753,N_19342);
xor U20771 (N_20771,N_17750,N_19936);
nor U20772 (N_20772,N_19203,N_19448);
nor U20773 (N_20773,N_19717,N_18182);
nand U20774 (N_20774,N_17712,N_19122);
or U20775 (N_20775,N_19318,N_19926);
nor U20776 (N_20776,N_17529,N_18281);
and U20777 (N_20777,N_18823,N_18109);
nor U20778 (N_20778,N_19731,N_17877);
or U20779 (N_20779,N_19310,N_19665);
nand U20780 (N_20780,N_18485,N_19606);
nor U20781 (N_20781,N_17704,N_19158);
xor U20782 (N_20782,N_17626,N_17641);
and U20783 (N_20783,N_18156,N_18769);
nor U20784 (N_20784,N_18880,N_18771);
or U20785 (N_20785,N_19065,N_17699);
xor U20786 (N_20786,N_18022,N_17652);
and U20787 (N_20787,N_17634,N_19498);
xor U20788 (N_20788,N_19943,N_19116);
and U20789 (N_20789,N_19497,N_19978);
and U20790 (N_20790,N_17862,N_19226);
xor U20791 (N_20791,N_19983,N_18547);
nor U20792 (N_20792,N_17934,N_19595);
and U20793 (N_20793,N_17911,N_19016);
nor U20794 (N_20794,N_17631,N_17900);
xor U20795 (N_20795,N_19824,N_17681);
or U20796 (N_20796,N_19512,N_17531);
and U20797 (N_20797,N_18922,N_17942);
xor U20798 (N_20798,N_18440,N_19500);
xnor U20799 (N_20799,N_18154,N_19621);
nand U20800 (N_20800,N_18766,N_18919);
and U20801 (N_20801,N_19118,N_18269);
nand U20802 (N_20802,N_17777,N_19322);
and U20803 (N_20803,N_19676,N_17822);
nand U20804 (N_20804,N_19846,N_18125);
nor U20805 (N_20805,N_18084,N_18603);
and U20806 (N_20806,N_18339,N_17884);
or U20807 (N_20807,N_17689,N_19631);
and U20808 (N_20808,N_17983,N_19004);
xor U20809 (N_20809,N_19001,N_19845);
xor U20810 (N_20810,N_19165,N_18955);
xor U20811 (N_20811,N_19873,N_19790);
nand U20812 (N_20812,N_19200,N_18564);
or U20813 (N_20813,N_19997,N_19301);
or U20814 (N_20814,N_18694,N_17563);
and U20815 (N_20815,N_18198,N_19083);
xnor U20816 (N_20816,N_18012,N_17678);
nor U20817 (N_20817,N_18611,N_18876);
nand U20818 (N_20818,N_18966,N_19950);
xor U20819 (N_20819,N_18196,N_18040);
xor U20820 (N_20820,N_19275,N_18287);
or U20821 (N_20821,N_19888,N_19652);
or U20822 (N_20822,N_18273,N_17853);
nand U20823 (N_20823,N_18624,N_19059);
or U20824 (N_20824,N_19434,N_19809);
and U20825 (N_20825,N_19271,N_19211);
nor U20826 (N_20826,N_19061,N_18264);
nand U20827 (N_20827,N_19534,N_17937);
nand U20828 (N_20828,N_18080,N_19585);
or U20829 (N_20829,N_17808,N_18580);
xor U20830 (N_20830,N_18244,N_18703);
xor U20831 (N_20831,N_18062,N_19101);
and U20832 (N_20832,N_19044,N_18208);
xnor U20833 (N_20833,N_18812,N_18369);
or U20834 (N_20834,N_18938,N_19416);
xnor U20835 (N_20835,N_19267,N_19429);
or U20836 (N_20836,N_19306,N_18807);
or U20837 (N_20837,N_19519,N_18249);
and U20838 (N_20838,N_18573,N_17875);
nor U20839 (N_20839,N_17883,N_18449);
xnor U20840 (N_20840,N_18973,N_18199);
nand U20841 (N_20841,N_18746,N_19857);
or U20842 (N_20842,N_19959,N_17736);
and U20843 (N_20843,N_18377,N_18026);
nor U20844 (N_20844,N_19372,N_19508);
nand U20845 (N_20845,N_19627,N_19302);
xnor U20846 (N_20846,N_18536,N_17826);
or U20847 (N_20847,N_17560,N_18625);
nor U20848 (N_20848,N_19640,N_17819);
and U20849 (N_20849,N_18729,N_18592);
or U20850 (N_20850,N_18496,N_19030);
nor U20851 (N_20851,N_19569,N_17702);
xor U20852 (N_20852,N_18609,N_19808);
or U20853 (N_20853,N_18559,N_18070);
and U20854 (N_20854,N_18480,N_19760);
and U20855 (N_20855,N_18232,N_19852);
or U20856 (N_20856,N_18143,N_19082);
nor U20857 (N_20857,N_19197,N_19092);
or U20858 (N_20858,N_19242,N_19851);
or U20859 (N_20859,N_18803,N_19043);
xnor U20860 (N_20860,N_17999,N_18635);
and U20861 (N_20861,N_17713,N_19413);
nor U20862 (N_20862,N_18710,N_19359);
or U20863 (N_20863,N_18540,N_18519);
and U20864 (N_20864,N_19894,N_18777);
and U20865 (N_20865,N_19683,N_17590);
or U20866 (N_20866,N_18513,N_19829);
and U20867 (N_20867,N_18410,N_19675);
nor U20868 (N_20868,N_17992,N_19869);
xnor U20869 (N_20869,N_17572,N_19558);
and U20870 (N_20870,N_18330,N_18484);
and U20871 (N_20871,N_17673,N_18589);
xor U20872 (N_20872,N_18285,N_19287);
and U20873 (N_20873,N_19656,N_18219);
xnor U20874 (N_20874,N_17644,N_18770);
nor U20875 (N_20875,N_18575,N_19893);
or U20876 (N_20876,N_17636,N_19087);
or U20877 (N_20877,N_19584,N_18457);
nand U20878 (N_20878,N_19989,N_19193);
and U20879 (N_20879,N_19295,N_18871);
or U20880 (N_20880,N_19266,N_17694);
and U20881 (N_20881,N_18845,N_19208);
or U20882 (N_20882,N_19549,N_18723);
nor U20883 (N_20883,N_18066,N_18430);
or U20884 (N_20884,N_18092,N_17546);
or U20885 (N_20885,N_18098,N_19370);
nand U20886 (N_20886,N_18814,N_18435);
nand U20887 (N_20887,N_18332,N_19259);
and U20888 (N_20888,N_17710,N_18554);
xor U20889 (N_20889,N_18500,N_19750);
nand U20890 (N_20890,N_18035,N_18013);
nor U20891 (N_20891,N_17748,N_19895);
nand U20892 (N_20892,N_18894,N_17924);
or U20893 (N_20893,N_18760,N_18187);
nand U20894 (N_20894,N_18842,N_18673);
and U20895 (N_20895,N_17892,N_19011);
nand U20896 (N_20896,N_19987,N_19304);
and U20897 (N_20897,N_18241,N_19088);
or U20898 (N_20898,N_19777,N_19575);
and U20899 (N_20899,N_18214,N_18552);
or U20900 (N_20900,N_18848,N_18758);
and U20901 (N_20901,N_17816,N_17779);
nor U20902 (N_20902,N_17556,N_19625);
nand U20903 (N_20903,N_18739,N_18389);
xor U20904 (N_20904,N_18290,N_18666);
nand U20905 (N_20905,N_17988,N_18686);
nor U20906 (N_20906,N_18059,N_18692);
or U20907 (N_20907,N_19347,N_19918);
or U20908 (N_20908,N_19671,N_18132);
and U20909 (N_20909,N_17785,N_17662);
nor U20910 (N_20910,N_19147,N_19340);
or U20911 (N_20911,N_17950,N_19254);
and U20912 (N_20912,N_17932,N_19615);
or U20913 (N_20913,N_18005,N_17734);
xnor U20914 (N_20914,N_17666,N_18856);
nand U20915 (N_20915,N_17530,N_19963);
nor U20916 (N_20916,N_18764,N_18889);
and U20917 (N_20917,N_19854,N_19361);
xor U20918 (N_20918,N_18476,N_17909);
xnor U20919 (N_20919,N_17525,N_19281);
and U20920 (N_20920,N_18464,N_17918);
nor U20921 (N_20921,N_18805,N_18505);
nor U20922 (N_20922,N_18459,N_18315);
nor U20923 (N_20923,N_19836,N_19080);
or U20924 (N_20924,N_18835,N_18102);
or U20925 (N_20925,N_19366,N_19536);
nor U20926 (N_20926,N_19235,N_18140);
xnor U20927 (N_20927,N_18216,N_17561);
xnor U20928 (N_20928,N_17685,N_18785);
xor U20929 (N_20929,N_19146,N_19097);
xnor U20930 (N_20930,N_17906,N_19540);
or U20931 (N_20931,N_18089,N_19690);
nor U20932 (N_20932,N_17982,N_19002);
nor U20933 (N_20933,N_18462,N_19105);
or U20934 (N_20934,N_18110,N_18514);
or U20935 (N_20935,N_18790,N_18907);
nand U20936 (N_20936,N_18587,N_18481);
or U20937 (N_20937,N_17843,N_18706);
xor U20938 (N_20938,N_19513,N_18348);
nand U20939 (N_20939,N_17690,N_18206);
nand U20940 (N_20940,N_19660,N_19581);
nand U20941 (N_20941,N_17548,N_18397);
nor U20942 (N_20942,N_19551,N_18749);
or U20943 (N_20943,N_19186,N_19386);
nand U20944 (N_20944,N_18548,N_18284);
or U20945 (N_20945,N_18471,N_19135);
or U20946 (N_20946,N_18757,N_19176);
xor U20947 (N_20947,N_18010,N_18750);
and U20948 (N_20948,N_17896,N_18088);
or U20949 (N_20949,N_18129,N_17597);
or U20950 (N_20950,N_19529,N_19177);
nor U20951 (N_20951,N_19971,N_18455);
and U20952 (N_20952,N_17949,N_19928);
xnor U20953 (N_20953,N_17562,N_18233);
and U20954 (N_20954,N_19883,N_18107);
or U20955 (N_20955,N_17967,N_19110);
nor U20956 (N_20956,N_19407,N_17654);
nand U20957 (N_20957,N_18276,N_17828);
and U20958 (N_20958,N_18292,N_19309);
nor U20959 (N_20959,N_17830,N_19486);
nor U20960 (N_20960,N_17635,N_18183);
xnor U20961 (N_20961,N_18319,N_19106);
xor U20962 (N_20962,N_18898,N_17580);
or U20963 (N_20963,N_18711,N_19783);
nand U20964 (N_20964,N_19313,N_17507);
nor U20965 (N_20965,N_19791,N_18726);
nor U20966 (N_20966,N_19637,N_19086);
nor U20967 (N_20967,N_19453,N_18212);
nor U20968 (N_20968,N_17599,N_18479);
and U20969 (N_20969,N_19330,N_17960);
nand U20970 (N_20970,N_18360,N_18370);
nand U20971 (N_20971,N_18017,N_17629);
nand U20972 (N_20972,N_19522,N_18953);
and U20973 (N_20973,N_18119,N_17663);
or U20974 (N_20974,N_18355,N_17512);
or U20975 (N_20975,N_18251,N_17501);
or U20976 (N_20976,N_18668,N_19516);
nand U20977 (N_20977,N_18539,N_18762);
nor U20978 (N_20978,N_18595,N_18442);
or U20979 (N_20979,N_19066,N_17547);
xor U20980 (N_20980,N_19227,N_19686);
nor U20981 (N_20981,N_19072,N_19199);
and U20982 (N_20982,N_18142,N_18331);
and U20983 (N_20983,N_17613,N_19802);
xor U20984 (N_20984,N_17583,N_19945);
xnor U20985 (N_20985,N_19089,N_19620);
or U20986 (N_20986,N_17810,N_17768);
nand U20987 (N_20987,N_19905,N_18942);
or U20988 (N_20988,N_18978,N_17829);
xnor U20989 (N_20989,N_17847,N_18593);
or U20990 (N_20990,N_19680,N_18063);
or U20991 (N_20991,N_19292,N_17579);
xor U20992 (N_20992,N_18103,N_19093);
and U20993 (N_20993,N_19160,N_19990);
or U20994 (N_20994,N_18755,N_19228);
and U20995 (N_20995,N_17659,N_18078);
nor U20996 (N_20996,N_18543,N_19444);
nor U20997 (N_20997,N_19345,N_18189);
nor U20998 (N_20998,N_19230,N_18550);
or U20999 (N_20999,N_19412,N_18974);
nor U21000 (N_21000,N_18939,N_18054);
nand U21001 (N_21001,N_17965,N_19754);
or U21002 (N_21002,N_19034,N_19763);
and U21003 (N_21003,N_19482,N_17508);
and U21004 (N_21004,N_18126,N_19374);
xnor U21005 (N_21005,N_19261,N_18567);
nor U21006 (N_21006,N_18912,N_19855);
and U21007 (N_21007,N_18043,N_17792);
or U21008 (N_21008,N_19788,N_17555);
xnor U21009 (N_21009,N_19333,N_19274);
and U21010 (N_21010,N_19958,N_17959);
xor U21011 (N_21011,N_19520,N_17503);
and U21012 (N_21012,N_18992,N_17751);
and U21013 (N_21013,N_17766,N_19727);
xnor U21014 (N_21014,N_17874,N_19411);
xnor U21015 (N_21015,N_18791,N_17991);
xnor U21016 (N_21016,N_18822,N_17687);
and U21017 (N_21017,N_19985,N_18528);
or U21018 (N_21018,N_18300,N_18844);
nor U21019 (N_21019,N_18675,N_17926);
or U21020 (N_21020,N_18321,N_19119);
xor U21021 (N_21021,N_19935,N_18761);
and U21022 (N_21022,N_18312,N_19920);
nor U21023 (N_21023,N_18134,N_19908);
or U21024 (N_21024,N_19175,N_19849);
nor U21025 (N_21025,N_18581,N_18618);
and U21026 (N_21026,N_19418,N_17740);
xor U21027 (N_21027,N_18903,N_19078);
or U21028 (N_21028,N_18003,N_18680);
xor U21029 (N_21029,N_18937,N_17981);
or U21030 (N_21030,N_19554,N_17951);
nor U21031 (N_21031,N_18950,N_17745);
nand U21032 (N_21032,N_17802,N_18951);
nand U21033 (N_21033,N_19432,N_19343);
and U21034 (N_21034,N_17797,N_18124);
xor U21035 (N_21035,N_18792,N_18145);
or U21036 (N_21036,N_19921,N_19948);
nor U21037 (N_21037,N_19045,N_17549);
nor U21038 (N_21038,N_17598,N_18177);
xor U21039 (N_21039,N_19128,N_19794);
nor U21040 (N_21040,N_18834,N_19813);
nor U21041 (N_21041,N_19240,N_18650);
or U21042 (N_21042,N_18910,N_19127);
xor U21043 (N_21043,N_19703,N_19046);
and U21044 (N_21044,N_19823,N_18883);
xnor U21045 (N_21045,N_19882,N_19020);
xnor U21046 (N_21046,N_19782,N_19285);
and U21047 (N_21047,N_18868,N_18877);
nor U21048 (N_21048,N_19530,N_19566);
nor U21049 (N_21049,N_19243,N_19210);
or U21050 (N_21050,N_18643,N_19191);
and U21051 (N_21051,N_19039,N_18171);
nand U21052 (N_21052,N_19171,N_19196);
nor U21053 (N_21053,N_19296,N_19833);
nor U21054 (N_21054,N_18021,N_18488);
nand U21055 (N_21055,N_18023,N_18531);
or U21056 (N_21056,N_18831,N_18956);
nand U21057 (N_21057,N_19544,N_18699);
xor U21058 (N_21058,N_17957,N_19556);
and U21059 (N_21059,N_18808,N_19706);
nand U21060 (N_21060,N_17765,N_18721);
xor U21061 (N_21061,N_19761,N_19115);
and U21062 (N_21062,N_18441,N_17731);
nor U21063 (N_21063,N_18133,N_18327);
nand U21064 (N_21064,N_17920,N_18313);
nand U21065 (N_21065,N_18747,N_19460);
xnor U21066 (N_21066,N_17543,N_19933);
nand U21067 (N_21067,N_19423,N_17586);
nand U21068 (N_21068,N_17781,N_18837);
and U21069 (N_21069,N_18225,N_18691);
or U21070 (N_21070,N_19810,N_19490);
and U21071 (N_21071,N_19828,N_18959);
nand U21072 (N_21072,N_19371,N_18613);
nor U21073 (N_21073,N_19856,N_18008);
nand U21074 (N_21074,N_17707,N_18700);
nor U21075 (N_21075,N_18427,N_18112);
xnor U21076 (N_21076,N_19817,N_19605);
and U21077 (N_21077,N_18470,N_17836);
or U21078 (N_21078,N_19435,N_19850);
and U21079 (N_21079,N_18060,N_18144);
and U21080 (N_21080,N_19476,N_19718);
and U21081 (N_21081,N_18200,N_17623);
or U21082 (N_21082,N_19289,N_19867);
nor U21083 (N_21083,N_18338,N_18057);
nand U21084 (N_21084,N_19739,N_17919);
nor U21085 (N_21085,N_19320,N_18168);
nand U21086 (N_21086,N_18186,N_18028);
and U21087 (N_21087,N_18058,N_19447);
nor U21088 (N_21088,N_19006,N_18754);
or U21089 (N_21089,N_18733,N_19687);
xor U21090 (N_21090,N_17990,N_19234);
nand U21091 (N_21091,N_17958,N_19143);
xor U21092 (N_21092,N_18826,N_17604);
xnor U21093 (N_21093,N_18051,N_19570);
and U21094 (N_21094,N_17655,N_18085);
nor U21095 (N_21095,N_18958,N_18347);
or U21096 (N_21096,N_19736,N_18473);
and U21097 (N_21097,N_19161,N_17784);
nor U21098 (N_21098,N_19009,N_18115);
or U21099 (N_21099,N_19691,N_18751);
and U21100 (N_21100,N_19136,N_18262);
and U21101 (N_21101,N_18393,N_18340);
and U21102 (N_21102,N_18682,N_17609);
and U21103 (N_21103,N_18246,N_18375);
and U21104 (N_21104,N_18824,N_18676);
and U21105 (N_21105,N_19840,N_18428);
xor U21106 (N_21106,N_19876,N_19502);
and U21107 (N_21107,N_18557,N_18657);
nor U21108 (N_21108,N_19315,N_19003);
or U21109 (N_21109,N_18857,N_17541);
xnor U21110 (N_21110,N_18414,N_18601);
or U21111 (N_21111,N_18660,N_18242);
nand U21112 (N_21112,N_18483,N_17989);
nand U21113 (N_21113,N_18025,N_18318);
nand U21114 (N_21114,N_18965,N_18840);
nor U21115 (N_21115,N_17872,N_17834);
nor U21116 (N_21116,N_18149,N_17974);
or U21117 (N_21117,N_17871,N_19053);
or U21118 (N_21118,N_19531,N_18551);
xnor U21119 (N_21119,N_19587,N_17725);
nor U21120 (N_21120,N_17559,N_19643);
and U21121 (N_21121,N_19698,N_19425);
and U21122 (N_21122,N_19380,N_18520);
nor U21123 (N_21123,N_19184,N_19000);
or U21124 (N_21124,N_19015,N_19051);
nor U21125 (N_21125,N_19487,N_19125);
xor U21126 (N_21126,N_19607,N_18887);
xnor U21127 (N_21127,N_19381,N_19901);
nand U21128 (N_21128,N_18778,N_19887);
or U21129 (N_21129,N_17986,N_19664);
nor U21130 (N_21130,N_19780,N_18205);
nor U21131 (N_21131,N_18361,N_18094);
xor U21132 (N_21132,N_18152,N_19798);
nor U21133 (N_21133,N_18633,N_19076);
and U21134 (N_21134,N_18545,N_17894);
and U21135 (N_21135,N_19757,N_18438);
xnor U21136 (N_21136,N_17845,N_17737);
and U21137 (N_21137,N_19613,N_18648);
xor U21138 (N_21138,N_18752,N_19737);
nor U21139 (N_21139,N_18268,N_19639);
xor U21140 (N_21140,N_19713,N_17620);
nand U21141 (N_21141,N_18725,N_19096);
or U21142 (N_21142,N_18989,N_18490);
nand U21143 (N_21143,N_17796,N_19778);
nor U21144 (N_21144,N_19701,N_18461);
nor U21145 (N_21145,N_17660,N_18372);
nor U21146 (N_21146,N_18841,N_19037);
xor U21147 (N_21147,N_18830,N_17809);
or U21148 (N_21148,N_18209,N_19164);
nand U21149 (N_21149,N_19248,N_19114);
xnor U21150 (N_21150,N_18636,N_19077);
or U21151 (N_21151,N_19906,N_17621);
nand U21152 (N_21152,N_19247,N_18436);
and U21153 (N_21153,N_19626,N_18314);
xor U21154 (N_21154,N_17878,N_19388);
and U21155 (N_21155,N_19961,N_18943);
and U21156 (N_21156,N_19117,N_19688);
nor U21157 (N_21157,N_19547,N_19735);
nor U21158 (N_21158,N_18798,N_18064);
xor U21159 (N_21159,N_18534,N_17970);
xnor U21160 (N_21160,N_18289,N_17787);
nand U21161 (N_21161,N_18477,N_19457);
xor U21162 (N_21162,N_19941,N_18400);
or U21163 (N_21163,N_19036,N_19049);
and U21164 (N_21164,N_19335,N_19741);
or U21165 (N_21165,N_18858,N_17788);
xnor U21166 (N_21166,N_17881,N_18968);
xnor U21167 (N_21167,N_17778,N_19899);
nand U21168 (N_21168,N_19699,N_19787);
and U21169 (N_21169,N_18371,N_17780);
or U21170 (N_21170,N_18398,N_18510);
nand U21171 (N_21171,N_19738,N_19430);
nor U21172 (N_21172,N_19662,N_19726);
nand U21173 (N_21173,N_17537,N_19525);
nor U21174 (N_21174,N_19685,N_19312);
xnor U21175 (N_21175,N_18653,N_18615);
nor U21176 (N_21176,N_18446,N_19792);
and U21177 (N_21177,N_18662,N_17672);
nand U21178 (N_21178,N_19332,N_19862);
nand U21179 (N_21179,N_19293,N_18870);
and U21180 (N_21180,N_19721,N_19494);
xnor U21181 (N_21181,N_18952,N_18405);
or U21182 (N_21182,N_19835,N_18271);
xnor U21183 (N_21183,N_18299,N_19789);
nand U21184 (N_21184,N_18714,N_17645);
nor U21185 (N_21185,N_19344,N_18879);
xor U21186 (N_21186,N_18853,N_18016);
or U21187 (N_21187,N_18067,N_18827);
nand U21188 (N_21188,N_18366,N_19659);
nand U21189 (N_21189,N_17931,N_19406);
and U21190 (N_21190,N_18652,N_17823);
xnor U21191 (N_21191,N_19559,N_18032);
nor U21192 (N_21192,N_18426,N_17774);
or U21193 (N_21193,N_19521,N_17688);
or U21194 (N_21194,N_19192,N_19527);
or U21195 (N_21195,N_18616,N_18849);
xor U21196 (N_21196,N_18174,N_19774);
nand U21197 (N_21197,N_19919,N_18722);
or U21198 (N_21198,N_17976,N_19268);
nand U21199 (N_21199,N_17628,N_17917);
or U21200 (N_21200,N_18521,N_19968);
nor U21201 (N_21201,N_17793,N_17890);
or U21202 (N_21202,N_19207,N_19298);
nor U21203 (N_21203,N_19528,N_18352);
xor U21204 (N_21204,N_19949,N_19561);
xor U21205 (N_21205,N_19917,N_19055);
nor U21206 (N_21206,N_19923,N_17984);
and U21207 (N_21207,N_18272,N_19202);
and U21208 (N_21208,N_18362,N_19967);
and U21209 (N_21209,N_19938,N_17738);
xnor U21210 (N_21210,N_17948,N_17910);
nand U21211 (N_21211,N_18349,N_17522);
and U21212 (N_21212,N_19469,N_19972);
nor U21213 (N_21213,N_19560,N_17524);
nand U21214 (N_21214,N_18644,N_18896);
nand U21215 (N_21215,N_19129,N_18763);
or U21216 (N_21216,N_18180,N_18069);
nand U21217 (N_21217,N_19946,N_18252);
nor U21218 (N_21218,N_18641,N_18874);
nor U21219 (N_21219,N_18784,N_18954);
or U21220 (N_21220,N_17691,N_19759);
xnor U21221 (N_21221,N_18915,N_18977);
xor U21222 (N_21222,N_17608,N_19623);
and U21223 (N_21223,N_19414,N_17567);
or U21224 (N_21224,N_18804,N_18788);
or U21225 (N_21225,N_18985,N_19163);
or U21226 (N_21226,N_19722,N_18402);
xnor U21227 (N_21227,N_19875,N_18560);
xnor U21228 (N_21228,N_17581,N_19934);
nand U21229 (N_21229,N_19733,N_18469);
nand U21230 (N_21230,N_18526,N_18068);
xnor U21231 (N_21231,N_18578,N_18195);
nand U21232 (N_21232,N_18210,N_18036);
and U21233 (N_21233,N_18509,N_18255);
xor U21234 (N_21234,N_18817,N_18596);
nand U21235 (N_21235,N_19473,N_17661);
or U21236 (N_21236,N_18875,N_18541);
nand U21237 (N_21237,N_18201,N_18001);
nor U21238 (N_21238,N_18359,N_19542);
or U21239 (N_21239,N_19264,N_19079);
or U21240 (N_21240,N_19622,N_18507);
and U21241 (N_21241,N_19140,N_19646);
nor U21242 (N_21242,N_19194,N_17578);
or U21243 (N_21243,N_19183,N_19394);
and U21244 (N_21244,N_19073,N_18065);
nand U21245 (N_21245,N_17600,N_19885);
xor U21246 (N_21246,N_19405,N_18162);
or U21247 (N_21247,N_19042,N_18705);
nor U21248 (N_21248,N_19290,N_18621);
and U21249 (N_21249,N_19784,N_18878);
or U21250 (N_21250,N_19062,N_17954);
or U21251 (N_21251,N_18498,N_19243);
nor U21252 (N_21252,N_17678,N_17941);
xnor U21253 (N_21253,N_19497,N_18405);
or U21254 (N_21254,N_19573,N_19356);
or U21255 (N_21255,N_18049,N_17891);
nand U21256 (N_21256,N_18140,N_19536);
and U21257 (N_21257,N_17603,N_19838);
xnor U21258 (N_21258,N_17543,N_19253);
xor U21259 (N_21259,N_18498,N_17699);
nand U21260 (N_21260,N_19714,N_19452);
nor U21261 (N_21261,N_17573,N_17791);
xnor U21262 (N_21262,N_19615,N_19885);
nand U21263 (N_21263,N_19111,N_19558);
nand U21264 (N_21264,N_19136,N_19185);
xnor U21265 (N_21265,N_19095,N_18536);
nor U21266 (N_21266,N_18009,N_19021);
nor U21267 (N_21267,N_19682,N_19186);
nor U21268 (N_21268,N_19274,N_19925);
or U21269 (N_21269,N_19670,N_18668);
nor U21270 (N_21270,N_18511,N_18825);
or U21271 (N_21271,N_18194,N_18075);
nor U21272 (N_21272,N_19604,N_18892);
or U21273 (N_21273,N_19781,N_18296);
nand U21274 (N_21274,N_18246,N_17658);
nor U21275 (N_21275,N_18444,N_18523);
or U21276 (N_21276,N_19890,N_18715);
xor U21277 (N_21277,N_18938,N_17751);
xnor U21278 (N_21278,N_17932,N_19849);
nor U21279 (N_21279,N_18219,N_18592);
nor U21280 (N_21280,N_18969,N_18546);
and U21281 (N_21281,N_18394,N_19477);
or U21282 (N_21282,N_19893,N_19127);
or U21283 (N_21283,N_18897,N_19088);
nand U21284 (N_21284,N_18582,N_19571);
nand U21285 (N_21285,N_18903,N_19747);
nand U21286 (N_21286,N_17800,N_18716);
or U21287 (N_21287,N_18860,N_17723);
nor U21288 (N_21288,N_18339,N_18326);
nor U21289 (N_21289,N_18820,N_18809);
xor U21290 (N_21290,N_18645,N_19849);
or U21291 (N_21291,N_17805,N_17735);
nor U21292 (N_21292,N_17653,N_17718);
nor U21293 (N_21293,N_18763,N_17886);
and U21294 (N_21294,N_18107,N_19168);
xnor U21295 (N_21295,N_19266,N_18977);
nand U21296 (N_21296,N_17979,N_18735);
xnor U21297 (N_21297,N_18146,N_18936);
and U21298 (N_21298,N_18896,N_17745);
xnor U21299 (N_21299,N_18971,N_17597);
xor U21300 (N_21300,N_19816,N_18093);
nand U21301 (N_21301,N_17712,N_19408);
nand U21302 (N_21302,N_19824,N_18019);
nor U21303 (N_21303,N_19696,N_17722);
or U21304 (N_21304,N_17732,N_17613);
xor U21305 (N_21305,N_19459,N_19314);
nand U21306 (N_21306,N_18311,N_17988);
or U21307 (N_21307,N_17723,N_17503);
nand U21308 (N_21308,N_18066,N_18855);
xor U21309 (N_21309,N_17693,N_18795);
xnor U21310 (N_21310,N_19619,N_18779);
and U21311 (N_21311,N_19353,N_18139);
and U21312 (N_21312,N_19018,N_18493);
or U21313 (N_21313,N_18933,N_19453);
nor U21314 (N_21314,N_19301,N_18067);
xor U21315 (N_21315,N_18919,N_18831);
or U21316 (N_21316,N_19411,N_19335);
xnor U21317 (N_21317,N_19770,N_19116);
and U21318 (N_21318,N_17742,N_17874);
or U21319 (N_21319,N_18100,N_18103);
nand U21320 (N_21320,N_18163,N_18105);
nand U21321 (N_21321,N_18133,N_18436);
nand U21322 (N_21322,N_18825,N_19433);
nand U21323 (N_21323,N_19230,N_19927);
and U21324 (N_21324,N_19242,N_18819);
and U21325 (N_21325,N_18713,N_18018);
and U21326 (N_21326,N_17898,N_19599);
xor U21327 (N_21327,N_18819,N_18001);
xnor U21328 (N_21328,N_18207,N_19595);
xor U21329 (N_21329,N_17674,N_19671);
nand U21330 (N_21330,N_19994,N_18245);
nor U21331 (N_21331,N_17934,N_18301);
and U21332 (N_21332,N_17840,N_18753);
and U21333 (N_21333,N_17747,N_19342);
xor U21334 (N_21334,N_18833,N_19365);
or U21335 (N_21335,N_19657,N_19354);
nor U21336 (N_21336,N_19381,N_19560);
xor U21337 (N_21337,N_17776,N_19413);
xor U21338 (N_21338,N_18480,N_19058);
nor U21339 (N_21339,N_19958,N_19499);
nand U21340 (N_21340,N_19952,N_19271);
or U21341 (N_21341,N_19519,N_18954);
and U21342 (N_21342,N_19063,N_19779);
nand U21343 (N_21343,N_19517,N_18046);
nor U21344 (N_21344,N_18724,N_18005);
nor U21345 (N_21345,N_18874,N_19350);
xnor U21346 (N_21346,N_19231,N_19977);
and U21347 (N_21347,N_17507,N_18529);
and U21348 (N_21348,N_19377,N_19043);
xnor U21349 (N_21349,N_18393,N_19780);
or U21350 (N_21350,N_18680,N_17553);
xnor U21351 (N_21351,N_19973,N_18611);
or U21352 (N_21352,N_17612,N_18134);
nor U21353 (N_21353,N_19035,N_19571);
xnor U21354 (N_21354,N_19671,N_17653);
xnor U21355 (N_21355,N_17591,N_18309);
or U21356 (N_21356,N_19417,N_18655);
xnor U21357 (N_21357,N_18883,N_18362);
and U21358 (N_21358,N_18805,N_18795);
or U21359 (N_21359,N_18204,N_19500);
nor U21360 (N_21360,N_19363,N_19393);
nand U21361 (N_21361,N_18917,N_19191);
xnor U21362 (N_21362,N_19641,N_18708);
nand U21363 (N_21363,N_18373,N_19913);
and U21364 (N_21364,N_18141,N_18736);
nand U21365 (N_21365,N_19203,N_17802);
nand U21366 (N_21366,N_18657,N_18540);
or U21367 (N_21367,N_17945,N_17849);
nand U21368 (N_21368,N_19732,N_19396);
xor U21369 (N_21369,N_18655,N_18740);
nand U21370 (N_21370,N_18640,N_18052);
and U21371 (N_21371,N_17585,N_19871);
and U21372 (N_21372,N_18863,N_17584);
nand U21373 (N_21373,N_18799,N_19122);
xnor U21374 (N_21374,N_18804,N_17666);
and U21375 (N_21375,N_18857,N_19980);
nor U21376 (N_21376,N_17922,N_18117);
xnor U21377 (N_21377,N_19023,N_17680);
and U21378 (N_21378,N_17674,N_17505);
xor U21379 (N_21379,N_19223,N_18829);
nand U21380 (N_21380,N_18994,N_19989);
or U21381 (N_21381,N_18115,N_18687);
nand U21382 (N_21382,N_18554,N_19194);
and U21383 (N_21383,N_18383,N_18789);
nor U21384 (N_21384,N_18261,N_18534);
nand U21385 (N_21385,N_19211,N_19871);
nor U21386 (N_21386,N_18763,N_19516);
nand U21387 (N_21387,N_19725,N_18233);
or U21388 (N_21388,N_18016,N_18134);
or U21389 (N_21389,N_18570,N_18362);
or U21390 (N_21390,N_19129,N_18735);
and U21391 (N_21391,N_19101,N_17525);
nor U21392 (N_21392,N_19553,N_17729);
nand U21393 (N_21393,N_19839,N_17706);
xnor U21394 (N_21394,N_19611,N_19103);
and U21395 (N_21395,N_18636,N_19435);
xor U21396 (N_21396,N_19856,N_18494);
and U21397 (N_21397,N_19255,N_17506);
or U21398 (N_21398,N_19646,N_17608);
xor U21399 (N_21399,N_17688,N_19982);
xor U21400 (N_21400,N_17871,N_18904);
nor U21401 (N_21401,N_19109,N_17575);
and U21402 (N_21402,N_17810,N_19656);
nor U21403 (N_21403,N_17768,N_17987);
or U21404 (N_21404,N_19773,N_17543);
or U21405 (N_21405,N_17888,N_19769);
and U21406 (N_21406,N_17623,N_17659);
or U21407 (N_21407,N_18149,N_18337);
nand U21408 (N_21408,N_18101,N_17873);
nor U21409 (N_21409,N_18395,N_19062);
nand U21410 (N_21410,N_17912,N_18022);
or U21411 (N_21411,N_18011,N_19141);
and U21412 (N_21412,N_17666,N_19528);
and U21413 (N_21413,N_19193,N_18564);
nor U21414 (N_21414,N_18395,N_18532);
and U21415 (N_21415,N_18922,N_18706);
nand U21416 (N_21416,N_18242,N_17767);
xnor U21417 (N_21417,N_18137,N_17656);
nand U21418 (N_21418,N_19021,N_17559);
nand U21419 (N_21419,N_19408,N_18223);
xnor U21420 (N_21420,N_18375,N_19169);
nand U21421 (N_21421,N_17689,N_19215);
xnor U21422 (N_21422,N_19943,N_18397);
or U21423 (N_21423,N_17935,N_18893);
nand U21424 (N_21424,N_19635,N_18631);
nand U21425 (N_21425,N_17655,N_19534);
nand U21426 (N_21426,N_18023,N_18487);
nor U21427 (N_21427,N_18997,N_18792);
nand U21428 (N_21428,N_18656,N_19762);
xnor U21429 (N_21429,N_18906,N_19696);
or U21430 (N_21430,N_18863,N_17725);
nor U21431 (N_21431,N_18343,N_19064);
or U21432 (N_21432,N_18320,N_19063);
or U21433 (N_21433,N_17940,N_18880);
nor U21434 (N_21434,N_17625,N_17562);
xnor U21435 (N_21435,N_17577,N_17948);
and U21436 (N_21436,N_17837,N_18573);
and U21437 (N_21437,N_19925,N_18737);
xor U21438 (N_21438,N_17581,N_19804);
and U21439 (N_21439,N_17725,N_18260);
and U21440 (N_21440,N_18733,N_18384);
nand U21441 (N_21441,N_19937,N_18477);
nor U21442 (N_21442,N_19446,N_17850);
nand U21443 (N_21443,N_18315,N_19511);
or U21444 (N_21444,N_19949,N_18240);
xor U21445 (N_21445,N_19909,N_19171);
or U21446 (N_21446,N_18034,N_19319);
or U21447 (N_21447,N_19522,N_18690);
and U21448 (N_21448,N_18423,N_18130);
xor U21449 (N_21449,N_19451,N_18896);
nor U21450 (N_21450,N_18364,N_18472);
nor U21451 (N_21451,N_18753,N_18364);
nor U21452 (N_21452,N_19916,N_19240);
xnor U21453 (N_21453,N_18384,N_17848);
xnor U21454 (N_21454,N_19320,N_19174);
xnor U21455 (N_21455,N_19533,N_19339);
xnor U21456 (N_21456,N_18668,N_17545);
or U21457 (N_21457,N_17570,N_18574);
xnor U21458 (N_21458,N_19436,N_19955);
nand U21459 (N_21459,N_19867,N_19590);
nand U21460 (N_21460,N_17576,N_19999);
and U21461 (N_21461,N_19822,N_18526);
or U21462 (N_21462,N_19928,N_19589);
or U21463 (N_21463,N_19562,N_18860);
and U21464 (N_21464,N_18797,N_18343);
xor U21465 (N_21465,N_17773,N_19464);
xnor U21466 (N_21466,N_17505,N_18524);
or U21467 (N_21467,N_17908,N_19817);
xor U21468 (N_21468,N_19302,N_18783);
or U21469 (N_21469,N_19254,N_18308);
xnor U21470 (N_21470,N_18781,N_18892);
nor U21471 (N_21471,N_19964,N_19650);
xnor U21472 (N_21472,N_19382,N_19046);
or U21473 (N_21473,N_18224,N_18023);
nand U21474 (N_21474,N_19616,N_19516);
xor U21475 (N_21475,N_19160,N_17730);
xnor U21476 (N_21476,N_18638,N_19876);
nand U21477 (N_21477,N_18793,N_18172);
nand U21478 (N_21478,N_17527,N_18966);
xor U21479 (N_21479,N_19493,N_18661);
nand U21480 (N_21480,N_18314,N_19432);
and U21481 (N_21481,N_19212,N_18719);
nand U21482 (N_21482,N_18324,N_19826);
or U21483 (N_21483,N_18526,N_18210);
nor U21484 (N_21484,N_18695,N_18688);
nand U21485 (N_21485,N_19768,N_19708);
and U21486 (N_21486,N_17912,N_19612);
nand U21487 (N_21487,N_18181,N_18342);
xor U21488 (N_21488,N_18830,N_18764);
xnor U21489 (N_21489,N_19891,N_19710);
and U21490 (N_21490,N_17673,N_18027);
or U21491 (N_21491,N_18175,N_18404);
nand U21492 (N_21492,N_19976,N_18275);
and U21493 (N_21493,N_17633,N_18018);
or U21494 (N_21494,N_19629,N_18761);
and U21495 (N_21495,N_19910,N_19054);
nor U21496 (N_21496,N_18111,N_18237);
nand U21497 (N_21497,N_18372,N_17641);
and U21498 (N_21498,N_19855,N_18725);
xnor U21499 (N_21499,N_18202,N_18599);
nand U21500 (N_21500,N_18672,N_19933);
nor U21501 (N_21501,N_19939,N_18924);
nor U21502 (N_21502,N_17808,N_19722);
xor U21503 (N_21503,N_19451,N_19403);
xor U21504 (N_21504,N_18056,N_18071);
or U21505 (N_21505,N_18535,N_17719);
xor U21506 (N_21506,N_18092,N_19952);
and U21507 (N_21507,N_18522,N_18836);
nor U21508 (N_21508,N_18673,N_19893);
and U21509 (N_21509,N_18283,N_19660);
xnor U21510 (N_21510,N_19046,N_17726);
xor U21511 (N_21511,N_18611,N_18340);
or U21512 (N_21512,N_18716,N_19569);
nand U21513 (N_21513,N_19129,N_19779);
or U21514 (N_21514,N_19051,N_18258);
nor U21515 (N_21515,N_19691,N_17995);
nor U21516 (N_21516,N_19139,N_18539);
and U21517 (N_21517,N_18655,N_19267);
nor U21518 (N_21518,N_18525,N_17543);
xnor U21519 (N_21519,N_17567,N_18729);
xnor U21520 (N_21520,N_18623,N_19252);
xor U21521 (N_21521,N_18322,N_17714);
or U21522 (N_21522,N_19890,N_19351);
nand U21523 (N_21523,N_19791,N_19776);
nor U21524 (N_21524,N_19669,N_19384);
nor U21525 (N_21525,N_18486,N_18923);
and U21526 (N_21526,N_19149,N_19695);
or U21527 (N_21527,N_18061,N_18183);
or U21528 (N_21528,N_18644,N_19232);
and U21529 (N_21529,N_19980,N_18564);
nand U21530 (N_21530,N_17660,N_18546);
nor U21531 (N_21531,N_19067,N_19361);
xnor U21532 (N_21532,N_18379,N_19564);
nand U21533 (N_21533,N_19453,N_18144);
nor U21534 (N_21534,N_19601,N_19086);
or U21535 (N_21535,N_18726,N_18161);
nand U21536 (N_21536,N_18685,N_19571);
or U21537 (N_21537,N_18158,N_18175);
nor U21538 (N_21538,N_18428,N_19566);
nor U21539 (N_21539,N_19753,N_18025);
nand U21540 (N_21540,N_18955,N_18048);
nand U21541 (N_21541,N_19637,N_18576);
and U21542 (N_21542,N_19867,N_19323);
and U21543 (N_21543,N_18153,N_18626);
nand U21544 (N_21544,N_17889,N_19065);
and U21545 (N_21545,N_19748,N_18574);
nor U21546 (N_21546,N_19534,N_19139);
xnor U21547 (N_21547,N_19569,N_18580);
and U21548 (N_21548,N_19270,N_18103);
nand U21549 (N_21549,N_19092,N_19659);
nor U21550 (N_21550,N_19290,N_17532);
and U21551 (N_21551,N_19218,N_19316);
and U21552 (N_21552,N_19646,N_19021);
and U21553 (N_21553,N_17725,N_17735);
nor U21554 (N_21554,N_17591,N_18047);
xnor U21555 (N_21555,N_17651,N_19145);
nand U21556 (N_21556,N_19906,N_17630);
nand U21557 (N_21557,N_17856,N_19912);
nand U21558 (N_21558,N_19381,N_17967);
xor U21559 (N_21559,N_18470,N_17819);
nand U21560 (N_21560,N_19438,N_19368);
nand U21561 (N_21561,N_17811,N_19441);
xnor U21562 (N_21562,N_18433,N_18323);
xor U21563 (N_21563,N_18412,N_19899);
xor U21564 (N_21564,N_17835,N_17682);
nand U21565 (N_21565,N_19892,N_18410);
xnor U21566 (N_21566,N_19598,N_18288);
xor U21567 (N_21567,N_17932,N_18927);
and U21568 (N_21568,N_18095,N_19638);
or U21569 (N_21569,N_17771,N_18291);
xor U21570 (N_21570,N_19375,N_17847);
nand U21571 (N_21571,N_17915,N_18208);
and U21572 (N_21572,N_18975,N_19590);
nor U21573 (N_21573,N_19494,N_17551);
xnor U21574 (N_21574,N_18638,N_18994);
nand U21575 (N_21575,N_19987,N_17625);
nor U21576 (N_21576,N_18679,N_19756);
nand U21577 (N_21577,N_19314,N_18087);
and U21578 (N_21578,N_18079,N_18964);
xor U21579 (N_21579,N_18619,N_17565);
xor U21580 (N_21580,N_18312,N_18795);
xor U21581 (N_21581,N_17949,N_18022);
xor U21582 (N_21582,N_19670,N_18564);
nor U21583 (N_21583,N_17934,N_17720);
nor U21584 (N_21584,N_18186,N_19441);
or U21585 (N_21585,N_17958,N_19841);
nor U21586 (N_21586,N_19323,N_19667);
or U21587 (N_21587,N_19214,N_18365);
or U21588 (N_21588,N_18719,N_17690);
nor U21589 (N_21589,N_17960,N_19835);
or U21590 (N_21590,N_19482,N_18508);
nor U21591 (N_21591,N_18091,N_19551);
nand U21592 (N_21592,N_17674,N_19314);
nor U21593 (N_21593,N_18751,N_18326);
and U21594 (N_21594,N_18320,N_18097);
or U21595 (N_21595,N_19026,N_18061);
nor U21596 (N_21596,N_18316,N_18503);
or U21597 (N_21597,N_19538,N_19982);
xor U21598 (N_21598,N_18885,N_18484);
xor U21599 (N_21599,N_19081,N_19554);
xor U21600 (N_21600,N_18366,N_18358);
and U21601 (N_21601,N_18723,N_17759);
and U21602 (N_21602,N_18164,N_19586);
or U21603 (N_21603,N_18774,N_19196);
or U21604 (N_21604,N_18164,N_19276);
nor U21605 (N_21605,N_19257,N_19630);
nand U21606 (N_21606,N_19998,N_19923);
nand U21607 (N_21607,N_19081,N_18256);
xnor U21608 (N_21608,N_19586,N_18961);
or U21609 (N_21609,N_19102,N_18134);
xor U21610 (N_21610,N_18821,N_19502);
and U21611 (N_21611,N_18432,N_19222);
nor U21612 (N_21612,N_17754,N_17888);
xor U21613 (N_21613,N_18322,N_19631);
nand U21614 (N_21614,N_18261,N_18242);
xor U21615 (N_21615,N_19905,N_18256);
or U21616 (N_21616,N_19933,N_18350);
nand U21617 (N_21617,N_18594,N_17747);
nor U21618 (N_21618,N_18556,N_17886);
xor U21619 (N_21619,N_19209,N_18791);
nor U21620 (N_21620,N_19188,N_18986);
xor U21621 (N_21621,N_19555,N_18461);
nand U21622 (N_21622,N_17769,N_18349);
xnor U21623 (N_21623,N_18299,N_17650);
and U21624 (N_21624,N_19107,N_19701);
xnor U21625 (N_21625,N_19042,N_18492);
xnor U21626 (N_21626,N_18055,N_19316);
and U21627 (N_21627,N_18627,N_19456);
nor U21628 (N_21628,N_19164,N_18311);
nor U21629 (N_21629,N_18146,N_18031);
nor U21630 (N_21630,N_17925,N_19196);
and U21631 (N_21631,N_19409,N_19568);
xor U21632 (N_21632,N_17575,N_18431);
or U21633 (N_21633,N_19972,N_17891);
xor U21634 (N_21634,N_18268,N_19889);
xor U21635 (N_21635,N_19992,N_19147);
xnor U21636 (N_21636,N_18758,N_19738);
xor U21637 (N_21637,N_18448,N_18469);
xnor U21638 (N_21638,N_19731,N_18126);
and U21639 (N_21639,N_18216,N_17860);
nor U21640 (N_21640,N_17781,N_18665);
xnor U21641 (N_21641,N_18930,N_19426);
nand U21642 (N_21642,N_19959,N_18512);
and U21643 (N_21643,N_19265,N_17660);
nand U21644 (N_21644,N_19383,N_19215);
or U21645 (N_21645,N_18666,N_18354);
nand U21646 (N_21646,N_17976,N_19139);
nand U21647 (N_21647,N_19501,N_19823);
xor U21648 (N_21648,N_18946,N_17730);
or U21649 (N_21649,N_19451,N_18305);
or U21650 (N_21650,N_18585,N_19786);
and U21651 (N_21651,N_19929,N_17592);
xor U21652 (N_21652,N_18831,N_18514);
and U21653 (N_21653,N_18366,N_17551);
nor U21654 (N_21654,N_19006,N_19305);
and U21655 (N_21655,N_18093,N_18886);
nand U21656 (N_21656,N_18397,N_19616);
xor U21657 (N_21657,N_17793,N_17923);
nand U21658 (N_21658,N_18463,N_18494);
xnor U21659 (N_21659,N_18136,N_19984);
xnor U21660 (N_21660,N_19478,N_19847);
xor U21661 (N_21661,N_19385,N_18793);
xnor U21662 (N_21662,N_19603,N_18591);
xnor U21663 (N_21663,N_19514,N_19321);
nor U21664 (N_21664,N_19890,N_18809);
nor U21665 (N_21665,N_18343,N_17597);
or U21666 (N_21666,N_18119,N_18477);
xor U21667 (N_21667,N_19405,N_17647);
xor U21668 (N_21668,N_19136,N_19048);
nor U21669 (N_21669,N_19812,N_17784);
xnor U21670 (N_21670,N_18201,N_19607);
nand U21671 (N_21671,N_17529,N_18398);
or U21672 (N_21672,N_19973,N_19556);
nand U21673 (N_21673,N_19294,N_18662);
nand U21674 (N_21674,N_19169,N_19715);
or U21675 (N_21675,N_19859,N_19669);
and U21676 (N_21676,N_19039,N_18802);
nand U21677 (N_21677,N_19296,N_17907);
xor U21678 (N_21678,N_18170,N_18082);
xnor U21679 (N_21679,N_19983,N_18415);
and U21680 (N_21680,N_18878,N_19386);
or U21681 (N_21681,N_17524,N_18821);
nor U21682 (N_21682,N_18414,N_19355);
and U21683 (N_21683,N_18631,N_19836);
xnor U21684 (N_21684,N_19954,N_17503);
xor U21685 (N_21685,N_19459,N_19039);
nor U21686 (N_21686,N_19876,N_17652);
xnor U21687 (N_21687,N_18494,N_19970);
nor U21688 (N_21688,N_18428,N_17716);
and U21689 (N_21689,N_19136,N_19429);
nand U21690 (N_21690,N_17733,N_18262);
nand U21691 (N_21691,N_19796,N_17601);
nand U21692 (N_21692,N_18202,N_18098);
xor U21693 (N_21693,N_17534,N_18529);
and U21694 (N_21694,N_18194,N_19891);
nor U21695 (N_21695,N_18708,N_19238);
nand U21696 (N_21696,N_18747,N_19407);
and U21697 (N_21697,N_17800,N_17705);
or U21698 (N_21698,N_19725,N_19928);
or U21699 (N_21699,N_19286,N_19293);
or U21700 (N_21700,N_19272,N_19818);
or U21701 (N_21701,N_17580,N_18819);
nand U21702 (N_21702,N_19931,N_18326);
and U21703 (N_21703,N_19792,N_18816);
and U21704 (N_21704,N_17797,N_19065);
and U21705 (N_21705,N_19512,N_18252);
nand U21706 (N_21706,N_18088,N_17503);
nand U21707 (N_21707,N_19326,N_19495);
or U21708 (N_21708,N_17950,N_18450);
xor U21709 (N_21709,N_18421,N_18513);
and U21710 (N_21710,N_18598,N_19954);
xor U21711 (N_21711,N_17854,N_19070);
xnor U21712 (N_21712,N_17771,N_18979);
or U21713 (N_21713,N_18583,N_17979);
and U21714 (N_21714,N_18444,N_17526);
or U21715 (N_21715,N_17559,N_18404);
nand U21716 (N_21716,N_18554,N_19269);
nor U21717 (N_21717,N_18042,N_19186);
or U21718 (N_21718,N_18858,N_17611);
nand U21719 (N_21719,N_18006,N_18503);
xor U21720 (N_21720,N_18167,N_18823);
or U21721 (N_21721,N_19139,N_19080);
or U21722 (N_21722,N_19937,N_17827);
or U21723 (N_21723,N_19317,N_18019);
nor U21724 (N_21724,N_18507,N_18037);
nor U21725 (N_21725,N_19543,N_18884);
nor U21726 (N_21726,N_18358,N_19884);
nor U21727 (N_21727,N_19550,N_17848);
nor U21728 (N_21728,N_19003,N_19916);
nor U21729 (N_21729,N_18473,N_19328);
nand U21730 (N_21730,N_18313,N_18439);
or U21731 (N_21731,N_19911,N_17987);
xnor U21732 (N_21732,N_19717,N_18050);
and U21733 (N_21733,N_17671,N_18227);
and U21734 (N_21734,N_17944,N_17783);
and U21735 (N_21735,N_19430,N_19695);
or U21736 (N_21736,N_19231,N_18755);
and U21737 (N_21737,N_18482,N_19109);
nand U21738 (N_21738,N_18968,N_18247);
or U21739 (N_21739,N_19320,N_18551);
nor U21740 (N_21740,N_19101,N_17589);
xor U21741 (N_21741,N_18545,N_19536);
xnor U21742 (N_21742,N_19997,N_19399);
and U21743 (N_21743,N_19380,N_19885);
nor U21744 (N_21744,N_17782,N_18082);
and U21745 (N_21745,N_17700,N_19532);
and U21746 (N_21746,N_17765,N_17783);
and U21747 (N_21747,N_17606,N_17602);
and U21748 (N_21748,N_18301,N_19156);
nand U21749 (N_21749,N_19191,N_17909);
or U21750 (N_21750,N_18495,N_18489);
xnor U21751 (N_21751,N_18220,N_17527);
xnor U21752 (N_21752,N_18732,N_18199);
nand U21753 (N_21753,N_18340,N_18753);
and U21754 (N_21754,N_19798,N_19696);
nand U21755 (N_21755,N_19002,N_17614);
xor U21756 (N_21756,N_18394,N_18767);
and U21757 (N_21757,N_19292,N_17639);
or U21758 (N_21758,N_18951,N_18350);
nand U21759 (N_21759,N_17623,N_19954);
nand U21760 (N_21760,N_18995,N_19748);
nor U21761 (N_21761,N_18010,N_19963);
nor U21762 (N_21762,N_19995,N_18118);
and U21763 (N_21763,N_18957,N_19216);
or U21764 (N_21764,N_19647,N_17967);
xor U21765 (N_21765,N_18769,N_18517);
or U21766 (N_21766,N_19708,N_18988);
xnor U21767 (N_21767,N_18512,N_19753);
nand U21768 (N_21768,N_19759,N_18685);
and U21769 (N_21769,N_19237,N_18653);
or U21770 (N_21770,N_18511,N_17689);
and U21771 (N_21771,N_19014,N_18360);
xnor U21772 (N_21772,N_18048,N_19871);
nand U21773 (N_21773,N_18260,N_17504);
xor U21774 (N_21774,N_19602,N_17679);
and U21775 (N_21775,N_18868,N_19741);
or U21776 (N_21776,N_18760,N_17762);
xor U21777 (N_21777,N_19041,N_17886);
or U21778 (N_21778,N_18298,N_19196);
nand U21779 (N_21779,N_19327,N_17891);
or U21780 (N_21780,N_17518,N_18531);
or U21781 (N_21781,N_18276,N_17514);
xor U21782 (N_21782,N_18365,N_18364);
and U21783 (N_21783,N_18616,N_17946);
xnor U21784 (N_21784,N_17681,N_18901);
or U21785 (N_21785,N_18770,N_18904);
and U21786 (N_21786,N_18866,N_17736);
nand U21787 (N_21787,N_18728,N_18716);
nand U21788 (N_21788,N_18328,N_18690);
nand U21789 (N_21789,N_19424,N_18837);
nand U21790 (N_21790,N_18047,N_19592);
or U21791 (N_21791,N_18904,N_17953);
nand U21792 (N_21792,N_19776,N_18355);
xor U21793 (N_21793,N_18776,N_18681);
or U21794 (N_21794,N_19074,N_17721);
nand U21795 (N_21795,N_19400,N_19083);
nor U21796 (N_21796,N_17671,N_17975);
nor U21797 (N_21797,N_17755,N_18929);
or U21798 (N_21798,N_18796,N_19031);
xnor U21799 (N_21799,N_19090,N_18621);
and U21800 (N_21800,N_18059,N_17521);
or U21801 (N_21801,N_17518,N_19404);
or U21802 (N_21802,N_18248,N_18353);
and U21803 (N_21803,N_17576,N_18766);
nor U21804 (N_21804,N_18643,N_19882);
xnor U21805 (N_21805,N_17883,N_18212);
nand U21806 (N_21806,N_19877,N_18046);
nand U21807 (N_21807,N_18837,N_17662);
and U21808 (N_21808,N_19501,N_19554);
nor U21809 (N_21809,N_19889,N_18688);
or U21810 (N_21810,N_19495,N_18103);
nor U21811 (N_21811,N_19162,N_17878);
nor U21812 (N_21812,N_19737,N_18330);
nand U21813 (N_21813,N_19222,N_17825);
and U21814 (N_21814,N_19015,N_19928);
or U21815 (N_21815,N_19544,N_19885);
nand U21816 (N_21816,N_19411,N_18383);
or U21817 (N_21817,N_18570,N_18621);
nand U21818 (N_21818,N_19152,N_18875);
xnor U21819 (N_21819,N_18982,N_18710);
or U21820 (N_21820,N_19534,N_18902);
xor U21821 (N_21821,N_19766,N_19310);
and U21822 (N_21822,N_19144,N_19682);
or U21823 (N_21823,N_19002,N_19304);
nor U21824 (N_21824,N_17502,N_19990);
and U21825 (N_21825,N_19287,N_19709);
nand U21826 (N_21826,N_19280,N_18730);
nand U21827 (N_21827,N_19753,N_19876);
nand U21828 (N_21828,N_18231,N_19933);
nand U21829 (N_21829,N_18400,N_19525);
nor U21830 (N_21830,N_17890,N_18436);
nor U21831 (N_21831,N_19387,N_18997);
nor U21832 (N_21832,N_19670,N_18658);
nand U21833 (N_21833,N_17779,N_18473);
or U21834 (N_21834,N_18667,N_19692);
nand U21835 (N_21835,N_18413,N_17584);
nand U21836 (N_21836,N_19822,N_17741);
xor U21837 (N_21837,N_18588,N_18351);
and U21838 (N_21838,N_18178,N_18002);
nor U21839 (N_21839,N_19819,N_19423);
and U21840 (N_21840,N_19143,N_17920);
xor U21841 (N_21841,N_19035,N_18549);
or U21842 (N_21842,N_19273,N_18023);
xnor U21843 (N_21843,N_19160,N_19972);
nand U21844 (N_21844,N_17843,N_19378);
and U21845 (N_21845,N_18022,N_18386);
nand U21846 (N_21846,N_18304,N_17900);
or U21847 (N_21847,N_19896,N_18875);
or U21848 (N_21848,N_18284,N_19701);
nor U21849 (N_21849,N_19344,N_19182);
nor U21850 (N_21850,N_18864,N_19009);
xnor U21851 (N_21851,N_18232,N_18807);
and U21852 (N_21852,N_17943,N_19031);
or U21853 (N_21853,N_19595,N_18319);
xnor U21854 (N_21854,N_18435,N_17799);
nor U21855 (N_21855,N_18650,N_19924);
and U21856 (N_21856,N_18070,N_19817);
nor U21857 (N_21857,N_19257,N_18712);
nor U21858 (N_21858,N_18926,N_18389);
or U21859 (N_21859,N_17693,N_18642);
or U21860 (N_21860,N_18002,N_18318);
or U21861 (N_21861,N_19742,N_19787);
or U21862 (N_21862,N_19972,N_19267);
nor U21863 (N_21863,N_18281,N_17629);
and U21864 (N_21864,N_18631,N_18536);
and U21865 (N_21865,N_18837,N_19924);
nand U21866 (N_21866,N_19404,N_18470);
nand U21867 (N_21867,N_18298,N_18014);
xnor U21868 (N_21868,N_17827,N_18352);
nor U21869 (N_21869,N_19869,N_19849);
or U21870 (N_21870,N_17706,N_17710);
xnor U21871 (N_21871,N_18265,N_17812);
xnor U21872 (N_21872,N_18080,N_19318);
nor U21873 (N_21873,N_17614,N_19351);
and U21874 (N_21874,N_19318,N_19702);
nand U21875 (N_21875,N_19645,N_19688);
and U21876 (N_21876,N_17590,N_19503);
nand U21877 (N_21877,N_17722,N_18399);
nand U21878 (N_21878,N_19327,N_19120);
nor U21879 (N_21879,N_18433,N_19166);
and U21880 (N_21880,N_17779,N_17520);
nor U21881 (N_21881,N_17864,N_19251);
nor U21882 (N_21882,N_17713,N_19295);
or U21883 (N_21883,N_18337,N_18324);
or U21884 (N_21884,N_17889,N_17673);
nand U21885 (N_21885,N_18693,N_19003);
xnor U21886 (N_21886,N_18048,N_18994);
xnor U21887 (N_21887,N_17587,N_18458);
xnor U21888 (N_21888,N_18418,N_18310);
nor U21889 (N_21889,N_18567,N_18311);
and U21890 (N_21890,N_18508,N_18188);
and U21891 (N_21891,N_18378,N_17669);
nor U21892 (N_21892,N_19210,N_18364);
xnor U21893 (N_21893,N_19019,N_19637);
nor U21894 (N_21894,N_18204,N_18323);
nand U21895 (N_21895,N_19444,N_17849);
nor U21896 (N_21896,N_19359,N_18616);
nor U21897 (N_21897,N_17592,N_19537);
nand U21898 (N_21898,N_19773,N_19694);
nor U21899 (N_21899,N_17584,N_19962);
or U21900 (N_21900,N_19067,N_17719);
and U21901 (N_21901,N_18926,N_19676);
nand U21902 (N_21902,N_19081,N_18568);
xor U21903 (N_21903,N_19709,N_18687);
nand U21904 (N_21904,N_17501,N_18724);
and U21905 (N_21905,N_19283,N_17846);
xnor U21906 (N_21906,N_18422,N_18386);
and U21907 (N_21907,N_18306,N_19875);
or U21908 (N_21908,N_17851,N_17906);
and U21909 (N_21909,N_19455,N_17658);
nor U21910 (N_21910,N_19103,N_18996);
nand U21911 (N_21911,N_18529,N_18924);
and U21912 (N_21912,N_19709,N_18190);
nand U21913 (N_21913,N_17532,N_18949);
nor U21914 (N_21914,N_19583,N_18505);
nor U21915 (N_21915,N_18762,N_18430);
and U21916 (N_21916,N_18705,N_18613);
xnor U21917 (N_21917,N_17522,N_17592);
nand U21918 (N_21918,N_19802,N_19921);
or U21919 (N_21919,N_17903,N_19643);
or U21920 (N_21920,N_18958,N_19500);
nand U21921 (N_21921,N_17778,N_19453);
or U21922 (N_21922,N_18604,N_17503);
xnor U21923 (N_21923,N_18209,N_19650);
or U21924 (N_21924,N_18122,N_19066);
nand U21925 (N_21925,N_18960,N_18683);
or U21926 (N_21926,N_17914,N_17521);
nand U21927 (N_21927,N_17548,N_18281);
xor U21928 (N_21928,N_19857,N_19213);
and U21929 (N_21929,N_17641,N_17774);
nor U21930 (N_21930,N_18066,N_19993);
xnor U21931 (N_21931,N_18292,N_19518);
and U21932 (N_21932,N_18834,N_18398);
xnor U21933 (N_21933,N_19226,N_19174);
xor U21934 (N_21934,N_17931,N_17959);
and U21935 (N_21935,N_18431,N_17901);
xor U21936 (N_21936,N_18843,N_17762);
xnor U21937 (N_21937,N_19169,N_18219);
nor U21938 (N_21938,N_18418,N_19470);
nand U21939 (N_21939,N_18214,N_18114);
and U21940 (N_21940,N_19742,N_19795);
xnor U21941 (N_21941,N_19343,N_17779);
and U21942 (N_21942,N_19258,N_17636);
xnor U21943 (N_21943,N_19755,N_18820);
or U21944 (N_21944,N_17732,N_19646);
nand U21945 (N_21945,N_19553,N_19350);
or U21946 (N_21946,N_17854,N_18029);
nor U21947 (N_21947,N_19490,N_19890);
xnor U21948 (N_21948,N_18583,N_17613);
xnor U21949 (N_21949,N_18550,N_18497);
xor U21950 (N_21950,N_19955,N_18645);
nand U21951 (N_21951,N_18696,N_17783);
nand U21952 (N_21952,N_18068,N_19159);
or U21953 (N_21953,N_18146,N_19354);
and U21954 (N_21954,N_17721,N_18347);
xnor U21955 (N_21955,N_19129,N_18651);
xnor U21956 (N_21956,N_19817,N_17543);
and U21957 (N_21957,N_18872,N_18241);
or U21958 (N_21958,N_18041,N_19716);
or U21959 (N_21959,N_19154,N_17647);
xnor U21960 (N_21960,N_18093,N_18690);
or U21961 (N_21961,N_19721,N_18241);
and U21962 (N_21962,N_19530,N_18214);
or U21963 (N_21963,N_19287,N_19090);
xnor U21964 (N_21964,N_18331,N_18303);
xnor U21965 (N_21965,N_19120,N_19603);
and U21966 (N_21966,N_17664,N_19148);
and U21967 (N_21967,N_18499,N_17605);
and U21968 (N_21968,N_19454,N_18135);
and U21969 (N_21969,N_19659,N_18351);
or U21970 (N_21970,N_18361,N_19940);
or U21971 (N_21971,N_19745,N_19212);
nand U21972 (N_21972,N_19128,N_19013);
xnor U21973 (N_21973,N_19965,N_19277);
nand U21974 (N_21974,N_19814,N_17995);
nand U21975 (N_21975,N_19779,N_19826);
and U21976 (N_21976,N_19219,N_17880);
nor U21977 (N_21977,N_17643,N_19726);
nor U21978 (N_21978,N_19023,N_17542);
or U21979 (N_21979,N_18766,N_18849);
and U21980 (N_21980,N_17893,N_18470);
xor U21981 (N_21981,N_19052,N_18534);
and U21982 (N_21982,N_18271,N_18189);
or U21983 (N_21983,N_19519,N_18384);
and U21984 (N_21984,N_19894,N_19263);
xor U21985 (N_21985,N_17692,N_17642);
and U21986 (N_21986,N_19691,N_17737);
or U21987 (N_21987,N_17760,N_18946);
and U21988 (N_21988,N_19918,N_19021);
nor U21989 (N_21989,N_18054,N_19854);
and U21990 (N_21990,N_19680,N_18561);
xor U21991 (N_21991,N_18206,N_19172);
or U21992 (N_21992,N_18044,N_19463);
or U21993 (N_21993,N_19332,N_17505);
xnor U21994 (N_21994,N_19646,N_17910);
or U21995 (N_21995,N_17741,N_18783);
or U21996 (N_21996,N_18148,N_18262);
nand U21997 (N_21997,N_18413,N_17928);
nand U21998 (N_21998,N_17596,N_18098);
and U21999 (N_21999,N_18595,N_19467);
or U22000 (N_22000,N_18548,N_19907);
and U22001 (N_22001,N_18475,N_19263);
or U22002 (N_22002,N_19788,N_19703);
nor U22003 (N_22003,N_19284,N_18685);
nand U22004 (N_22004,N_19185,N_18248);
nor U22005 (N_22005,N_19874,N_17908);
or U22006 (N_22006,N_19918,N_18381);
nand U22007 (N_22007,N_18720,N_19896);
and U22008 (N_22008,N_19279,N_19440);
xnor U22009 (N_22009,N_19457,N_19099);
nor U22010 (N_22010,N_19378,N_19593);
and U22011 (N_22011,N_18908,N_19374);
nand U22012 (N_22012,N_19010,N_19152);
nor U22013 (N_22013,N_19580,N_17509);
and U22014 (N_22014,N_18663,N_17994);
or U22015 (N_22015,N_19719,N_19897);
or U22016 (N_22016,N_18512,N_17969);
or U22017 (N_22017,N_19113,N_18509);
and U22018 (N_22018,N_18065,N_19882);
nor U22019 (N_22019,N_18643,N_18124);
xnor U22020 (N_22020,N_18879,N_19081);
and U22021 (N_22021,N_19573,N_19194);
xor U22022 (N_22022,N_19280,N_18822);
or U22023 (N_22023,N_18493,N_19612);
nor U22024 (N_22024,N_19812,N_19781);
nor U22025 (N_22025,N_18053,N_19461);
xor U22026 (N_22026,N_19297,N_19035);
nand U22027 (N_22027,N_19403,N_19514);
nor U22028 (N_22028,N_19059,N_19208);
xor U22029 (N_22029,N_19527,N_18931);
or U22030 (N_22030,N_18344,N_18276);
nand U22031 (N_22031,N_19569,N_18502);
nor U22032 (N_22032,N_18423,N_18539);
or U22033 (N_22033,N_19518,N_18060);
nand U22034 (N_22034,N_17886,N_19810);
and U22035 (N_22035,N_17706,N_17611);
xnor U22036 (N_22036,N_17804,N_19674);
nor U22037 (N_22037,N_19348,N_17671);
or U22038 (N_22038,N_19797,N_17790);
or U22039 (N_22039,N_18471,N_19840);
xor U22040 (N_22040,N_18955,N_18493);
nor U22041 (N_22041,N_17992,N_19103);
xor U22042 (N_22042,N_19056,N_18085);
and U22043 (N_22043,N_19307,N_18593);
xor U22044 (N_22044,N_18312,N_19368);
or U22045 (N_22045,N_17540,N_18098);
or U22046 (N_22046,N_18043,N_17921);
nand U22047 (N_22047,N_19058,N_17644);
or U22048 (N_22048,N_19692,N_19462);
or U22049 (N_22049,N_18263,N_17956);
and U22050 (N_22050,N_17662,N_18591);
nand U22051 (N_22051,N_18561,N_19076);
nor U22052 (N_22052,N_19424,N_17839);
or U22053 (N_22053,N_17799,N_19761);
nor U22054 (N_22054,N_17960,N_18582);
or U22055 (N_22055,N_18120,N_17939);
nand U22056 (N_22056,N_18352,N_19244);
or U22057 (N_22057,N_19924,N_17790);
nand U22058 (N_22058,N_18744,N_19339);
and U22059 (N_22059,N_17640,N_19604);
nand U22060 (N_22060,N_19191,N_19400);
or U22061 (N_22061,N_17625,N_17890);
and U22062 (N_22062,N_17775,N_19959);
nor U22063 (N_22063,N_18278,N_18695);
nand U22064 (N_22064,N_19823,N_18871);
or U22065 (N_22065,N_17904,N_19407);
xor U22066 (N_22066,N_18290,N_18357);
or U22067 (N_22067,N_19856,N_17609);
nor U22068 (N_22068,N_17739,N_19508);
xnor U22069 (N_22069,N_19503,N_18638);
and U22070 (N_22070,N_17686,N_18585);
or U22071 (N_22071,N_19272,N_19737);
nor U22072 (N_22072,N_19360,N_18178);
nor U22073 (N_22073,N_19126,N_18327);
nand U22074 (N_22074,N_17770,N_19367);
or U22075 (N_22075,N_17720,N_18910);
and U22076 (N_22076,N_19045,N_19006);
nor U22077 (N_22077,N_18528,N_18281);
nand U22078 (N_22078,N_19865,N_19517);
nand U22079 (N_22079,N_19761,N_18427);
nand U22080 (N_22080,N_18960,N_17761);
nor U22081 (N_22081,N_17891,N_19011);
and U22082 (N_22082,N_19135,N_18835);
nor U22083 (N_22083,N_17770,N_19055);
nor U22084 (N_22084,N_18486,N_19448);
xnor U22085 (N_22085,N_17882,N_19562);
and U22086 (N_22086,N_17701,N_18067);
nor U22087 (N_22087,N_17587,N_18184);
nand U22088 (N_22088,N_18757,N_19396);
nand U22089 (N_22089,N_19378,N_19221);
or U22090 (N_22090,N_17846,N_18699);
nand U22091 (N_22091,N_19039,N_18868);
xor U22092 (N_22092,N_17537,N_19602);
nand U22093 (N_22093,N_18521,N_18850);
and U22094 (N_22094,N_18624,N_19561);
nand U22095 (N_22095,N_18603,N_18079);
or U22096 (N_22096,N_18816,N_19893);
or U22097 (N_22097,N_18283,N_17613);
or U22098 (N_22098,N_19219,N_18736);
or U22099 (N_22099,N_19260,N_19736);
xnor U22100 (N_22100,N_19016,N_18284);
or U22101 (N_22101,N_17961,N_19171);
or U22102 (N_22102,N_19991,N_19920);
xnor U22103 (N_22103,N_19805,N_18805);
nor U22104 (N_22104,N_18916,N_17654);
and U22105 (N_22105,N_17789,N_19528);
xor U22106 (N_22106,N_19617,N_18459);
and U22107 (N_22107,N_17842,N_18597);
and U22108 (N_22108,N_18253,N_19044);
nand U22109 (N_22109,N_19701,N_17795);
nor U22110 (N_22110,N_18847,N_19816);
nor U22111 (N_22111,N_19069,N_18575);
or U22112 (N_22112,N_18297,N_18686);
nand U22113 (N_22113,N_18984,N_19741);
and U22114 (N_22114,N_18935,N_18029);
and U22115 (N_22115,N_18332,N_17736);
or U22116 (N_22116,N_18710,N_18953);
nor U22117 (N_22117,N_17808,N_19693);
or U22118 (N_22118,N_17943,N_18706);
or U22119 (N_22119,N_19294,N_19719);
or U22120 (N_22120,N_19006,N_17804);
and U22121 (N_22121,N_19408,N_18608);
nor U22122 (N_22122,N_18904,N_18072);
nor U22123 (N_22123,N_19203,N_18858);
and U22124 (N_22124,N_19294,N_18060);
or U22125 (N_22125,N_18188,N_19536);
xnor U22126 (N_22126,N_19308,N_19948);
xnor U22127 (N_22127,N_19492,N_18548);
nand U22128 (N_22128,N_18162,N_17865);
and U22129 (N_22129,N_18948,N_17863);
xnor U22130 (N_22130,N_18795,N_19967);
nand U22131 (N_22131,N_19377,N_18754);
xnor U22132 (N_22132,N_19656,N_18220);
nand U22133 (N_22133,N_17572,N_18618);
xor U22134 (N_22134,N_18760,N_18032);
and U22135 (N_22135,N_18048,N_18847);
and U22136 (N_22136,N_17790,N_18541);
and U22137 (N_22137,N_18722,N_18501);
nand U22138 (N_22138,N_18818,N_19544);
xor U22139 (N_22139,N_19928,N_18225);
nor U22140 (N_22140,N_18902,N_17641);
nor U22141 (N_22141,N_19587,N_19639);
xor U22142 (N_22142,N_18401,N_18347);
nor U22143 (N_22143,N_19913,N_18559);
nor U22144 (N_22144,N_19006,N_19984);
or U22145 (N_22145,N_18901,N_17723);
nand U22146 (N_22146,N_18275,N_19693);
and U22147 (N_22147,N_19001,N_19811);
nand U22148 (N_22148,N_18603,N_19111);
nand U22149 (N_22149,N_19807,N_19276);
xnor U22150 (N_22150,N_17782,N_18386);
or U22151 (N_22151,N_19676,N_19735);
or U22152 (N_22152,N_18342,N_17898);
and U22153 (N_22153,N_18471,N_18290);
xnor U22154 (N_22154,N_19502,N_19559);
and U22155 (N_22155,N_19920,N_19306);
xnor U22156 (N_22156,N_19600,N_18859);
xor U22157 (N_22157,N_19220,N_19202);
and U22158 (N_22158,N_17725,N_19829);
or U22159 (N_22159,N_18756,N_19127);
and U22160 (N_22160,N_18024,N_18719);
or U22161 (N_22161,N_18329,N_19290);
nand U22162 (N_22162,N_19240,N_18161);
nor U22163 (N_22163,N_17729,N_18340);
or U22164 (N_22164,N_19698,N_19087);
nor U22165 (N_22165,N_19233,N_18299);
and U22166 (N_22166,N_18113,N_19092);
xor U22167 (N_22167,N_19282,N_18323);
nor U22168 (N_22168,N_19055,N_19435);
or U22169 (N_22169,N_19402,N_17619);
nand U22170 (N_22170,N_18232,N_18251);
nand U22171 (N_22171,N_18427,N_17538);
nor U22172 (N_22172,N_18518,N_19944);
xor U22173 (N_22173,N_18211,N_19196);
or U22174 (N_22174,N_17743,N_19029);
and U22175 (N_22175,N_18169,N_17584);
or U22176 (N_22176,N_19358,N_19708);
or U22177 (N_22177,N_18910,N_18680);
xor U22178 (N_22178,N_19736,N_18822);
and U22179 (N_22179,N_17996,N_18202);
xor U22180 (N_22180,N_17578,N_19525);
or U22181 (N_22181,N_19795,N_17822);
nand U22182 (N_22182,N_19748,N_17971);
or U22183 (N_22183,N_18038,N_18911);
xor U22184 (N_22184,N_19429,N_17784);
xnor U22185 (N_22185,N_18055,N_18867);
and U22186 (N_22186,N_18253,N_19174);
or U22187 (N_22187,N_19804,N_19961);
and U22188 (N_22188,N_17531,N_18768);
nand U22189 (N_22189,N_19515,N_19244);
xor U22190 (N_22190,N_19880,N_18998);
nand U22191 (N_22191,N_18923,N_17954);
and U22192 (N_22192,N_18763,N_18849);
xnor U22193 (N_22193,N_19487,N_19267);
xor U22194 (N_22194,N_18555,N_18151);
nor U22195 (N_22195,N_19345,N_17681);
nand U22196 (N_22196,N_18915,N_19542);
and U22197 (N_22197,N_19482,N_19727);
nand U22198 (N_22198,N_19087,N_19208);
nor U22199 (N_22199,N_17566,N_19313);
and U22200 (N_22200,N_17669,N_18546);
nor U22201 (N_22201,N_18192,N_17935);
nand U22202 (N_22202,N_19576,N_18466);
and U22203 (N_22203,N_19783,N_18029);
nand U22204 (N_22204,N_18035,N_18777);
or U22205 (N_22205,N_18388,N_19204);
or U22206 (N_22206,N_17701,N_19979);
and U22207 (N_22207,N_19509,N_18597);
and U22208 (N_22208,N_19016,N_18411);
nand U22209 (N_22209,N_19805,N_18077);
nor U22210 (N_22210,N_18475,N_18657);
nand U22211 (N_22211,N_18141,N_17909);
nand U22212 (N_22212,N_18050,N_19119);
and U22213 (N_22213,N_19467,N_19409);
nor U22214 (N_22214,N_18886,N_17857);
nand U22215 (N_22215,N_18464,N_19837);
xnor U22216 (N_22216,N_17809,N_19737);
nand U22217 (N_22217,N_17728,N_18231);
or U22218 (N_22218,N_18104,N_19231);
nor U22219 (N_22219,N_19688,N_18667);
nand U22220 (N_22220,N_18880,N_17911);
nor U22221 (N_22221,N_18175,N_19212);
nor U22222 (N_22222,N_19007,N_19997);
and U22223 (N_22223,N_19106,N_18965);
xor U22224 (N_22224,N_19748,N_19118);
and U22225 (N_22225,N_18769,N_18635);
nand U22226 (N_22226,N_17775,N_17762);
and U22227 (N_22227,N_19920,N_19091);
nand U22228 (N_22228,N_19702,N_18693);
nand U22229 (N_22229,N_18124,N_19371);
nand U22230 (N_22230,N_19067,N_18804);
nand U22231 (N_22231,N_19752,N_17727);
and U22232 (N_22232,N_17541,N_17919);
xnor U22233 (N_22233,N_18712,N_18203);
nor U22234 (N_22234,N_18427,N_17559);
xor U22235 (N_22235,N_17976,N_19187);
nand U22236 (N_22236,N_18279,N_17988);
nor U22237 (N_22237,N_19023,N_17597);
nor U22238 (N_22238,N_18013,N_19214);
nand U22239 (N_22239,N_17925,N_19304);
nor U22240 (N_22240,N_19150,N_19854);
and U22241 (N_22241,N_18818,N_17607);
or U22242 (N_22242,N_19655,N_19032);
xor U22243 (N_22243,N_19454,N_19175);
nor U22244 (N_22244,N_18539,N_17752);
or U22245 (N_22245,N_19707,N_19948);
xor U22246 (N_22246,N_18190,N_18437);
nor U22247 (N_22247,N_19826,N_18844);
and U22248 (N_22248,N_19584,N_19354);
nor U22249 (N_22249,N_19155,N_18700);
nand U22250 (N_22250,N_19088,N_19213);
nand U22251 (N_22251,N_19587,N_19164);
nor U22252 (N_22252,N_19041,N_18393);
nand U22253 (N_22253,N_19145,N_18976);
nor U22254 (N_22254,N_19155,N_18290);
or U22255 (N_22255,N_19851,N_19801);
and U22256 (N_22256,N_19985,N_17740);
xnor U22257 (N_22257,N_18603,N_17792);
xnor U22258 (N_22258,N_17502,N_19902);
xnor U22259 (N_22259,N_18025,N_19388);
and U22260 (N_22260,N_19097,N_17871);
nor U22261 (N_22261,N_19691,N_17525);
and U22262 (N_22262,N_19657,N_17523);
and U22263 (N_22263,N_19001,N_17957);
nor U22264 (N_22264,N_19032,N_19625);
nor U22265 (N_22265,N_17598,N_18489);
and U22266 (N_22266,N_18370,N_19123);
and U22267 (N_22267,N_19013,N_18184);
and U22268 (N_22268,N_19355,N_18213);
nor U22269 (N_22269,N_18186,N_18758);
or U22270 (N_22270,N_19957,N_19035);
or U22271 (N_22271,N_18659,N_17708);
nand U22272 (N_22272,N_18193,N_19162);
and U22273 (N_22273,N_17876,N_19661);
xor U22274 (N_22274,N_17570,N_19973);
nand U22275 (N_22275,N_19159,N_18204);
nand U22276 (N_22276,N_17868,N_18844);
xnor U22277 (N_22277,N_19290,N_18456);
xnor U22278 (N_22278,N_19655,N_19318);
or U22279 (N_22279,N_19848,N_18946);
nor U22280 (N_22280,N_18354,N_18840);
nand U22281 (N_22281,N_18497,N_18799);
or U22282 (N_22282,N_17671,N_17838);
or U22283 (N_22283,N_18928,N_18052);
nor U22284 (N_22284,N_18697,N_18459);
xnor U22285 (N_22285,N_18017,N_19823);
nor U22286 (N_22286,N_18356,N_17985);
nand U22287 (N_22287,N_18096,N_18857);
xor U22288 (N_22288,N_19509,N_18259);
nand U22289 (N_22289,N_19980,N_17872);
and U22290 (N_22290,N_19044,N_18466);
xnor U22291 (N_22291,N_19894,N_19415);
and U22292 (N_22292,N_19293,N_17923);
or U22293 (N_22293,N_17561,N_19801);
or U22294 (N_22294,N_19803,N_19731);
xor U22295 (N_22295,N_18291,N_18143);
and U22296 (N_22296,N_18539,N_17550);
and U22297 (N_22297,N_18396,N_19745);
and U22298 (N_22298,N_19671,N_18720);
nor U22299 (N_22299,N_18489,N_19371);
xor U22300 (N_22300,N_17629,N_18372);
xnor U22301 (N_22301,N_17771,N_18523);
or U22302 (N_22302,N_17628,N_19255);
or U22303 (N_22303,N_18444,N_18627);
xnor U22304 (N_22304,N_18932,N_17822);
nand U22305 (N_22305,N_18495,N_19939);
or U22306 (N_22306,N_19431,N_19904);
and U22307 (N_22307,N_18725,N_18540);
and U22308 (N_22308,N_17610,N_17944);
xor U22309 (N_22309,N_18488,N_19449);
and U22310 (N_22310,N_19352,N_19940);
nand U22311 (N_22311,N_19259,N_18884);
xor U22312 (N_22312,N_17546,N_18559);
xor U22313 (N_22313,N_18036,N_19819);
nand U22314 (N_22314,N_18670,N_17919);
nand U22315 (N_22315,N_17709,N_19535);
nor U22316 (N_22316,N_18651,N_17916);
and U22317 (N_22317,N_18873,N_19478);
nor U22318 (N_22318,N_18200,N_18671);
nand U22319 (N_22319,N_17749,N_19192);
and U22320 (N_22320,N_19194,N_18517);
xnor U22321 (N_22321,N_18800,N_18796);
or U22322 (N_22322,N_18764,N_19634);
or U22323 (N_22323,N_18213,N_19054);
and U22324 (N_22324,N_18860,N_19626);
and U22325 (N_22325,N_19017,N_18391);
and U22326 (N_22326,N_17927,N_19807);
nor U22327 (N_22327,N_17682,N_19400);
nand U22328 (N_22328,N_19261,N_19041);
nor U22329 (N_22329,N_17938,N_18030);
nor U22330 (N_22330,N_18803,N_18972);
and U22331 (N_22331,N_19753,N_18161);
nand U22332 (N_22332,N_18910,N_18702);
and U22333 (N_22333,N_19943,N_18851);
xnor U22334 (N_22334,N_18309,N_18596);
nor U22335 (N_22335,N_18434,N_17738);
and U22336 (N_22336,N_17570,N_19285);
xnor U22337 (N_22337,N_18391,N_19922);
nand U22338 (N_22338,N_18491,N_18197);
nand U22339 (N_22339,N_19320,N_19004);
or U22340 (N_22340,N_18195,N_19495);
nand U22341 (N_22341,N_19905,N_19103);
nor U22342 (N_22342,N_19873,N_19265);
or U22343 (N_22343,N_17892,N_19091);
xor U22344 (N_22344,N_18365,N_17583);
and U22345 (N_22345,N_17886,N_19766);
and U22346 (N_22346,N_18409,N_17964);
xor U22347 (N_22347,N_19825,N_18710);
nor U22348 (N_22348,N_19297,N_18929);
xor U22349 (N_22349,N_18253,N_17628);
nor U22350 (N_22350,N_19838,N_19006);
or U22351 (N_22351,N_19434,N_18161);
nor U22352 (N_22352,N_19174,N_19814);
nand U22353 (N_22353,N_18403,N_17736);
xor U22354 (N_22354,N_18719,N_19280);
xor U22355 (N_22355,N_18947,N_17687);
xnor U22356 (N_22356,N_17830,N_17508);
nand U22357 (N_22357,N_18972,N_18870);
nor U22358 (N_22358,N_19714,N_18072);
nand U22359 (N_22359,N_18368,N_18263);
nor U22360 (N_22360,N_19787,N_18052);
and U22361 (N_22361,N_17657,N_18040);
nand U22362 (N_22362,N_18559,N_17882);
xor U22363 (N_22363,N_18408,N_19302);
nor U22364 (N_22364,N_18353,N_18225);
nor U22365 (N_22365,N_17885,N_18549);
xnor U22366 (N_22366,N_17975,N_19507);
or U22367 (N_22367,N_18012,N_18320);
nor U22368 (N_22368,N_18395,N_18103);
and U22369 (N_22369,N_19678,N_18191);
nand U22370 (N_22370,N_19819,N_18687);
nor U22371 (N_22371,N_18448,N_18136);
nand U22372 (N_22372,N_19967,N_19236);
nand U22373 (N_22373,N_17984,N_17696);
and U22374 (N_22374,N_18991,N_19499);
nor U22375 (N_22375,N_19859,N_19580);
nor U22376 (N_22376,N_19886,N_18100);
or U22377 (N_22377,N_18030,N_18949);
and U22378 (N_22378,N_19107,N_18719);
xor U22379 (N_22379,N_18142,N_18358);
or U22380 (N_22380,N_17916,N_19917);
nor U22381 (N_22381,N_18000,N_19584);
or U22382 (N_22382,N_19565,N_19463);
and U22383 (N_22383,N_19773,N_19738);
xor U22384 (N_22384,N_18677,N_19893);
or U22385 (N_22385,N_17576,N_17540);
and U22386 (N_22386,N_19203,N_18476);
or U22387 (N_22387,N_18423,N_19277);
xnor U22388 (N_22388,N_18096,N_18030);
xnor U22389 (N_22389,N_18126,N_17715);
nand U22390 (N_22390,N_17853,N_19935);
or U22391 (N_22391,N_19418,N_19986);
nand U22392 (N_22392,N_19527,N_18560);
xor U22393 (N_22393,N_18897,N_18438);
or U22394 (N_22394,N_17710,N_19031);
nand U22395 (N_22395,N_17858,N_19089);
nor U22396 (N_22396,N_19555,N_19964);
or U22397 (N_22397,N_19042,N_18610);
xnor U22398 (N_22398,N_17546,N_17788);
nor U22399 (N_22399,N_19530,N_19694);
nand U22400 (N_22400,N_17932,N_19230);
and U22401 (N_22401,N_19230,N_18218);
nor U22402 (N_22402,N_19509,N_19126);
nor U22403 (N_22403,N_19079,N_18595);
nor U22404 (N_22404,N_19498,N_17678);
or U22405 (N_22405,N_18134,N_17567);
nand U22406 (N_22406,N_19203,N_18540);
and U22407 (N_22407,N_18625,N_19922);
or U22408 (N_22408,N_19065,N_19446);
nor U22409 (N_22409,N_19824,N_19237);
and U22410 (N_22410,N_19433,N_19669);
nor U22411 (N_22411,N_19003,N_19016);
xor U22412 (N_22412,N_18066,N_19737);
xor U22413 (N_22413,N_19686,N_18659);
nor U22414 (N_22414,N_18741,N_18108);
nand U22415 (N_22415,N_17851,N_19693);
xor U22416 (N_22416,N_19013,N_18356);
xnor U22417 (N_22417,N_19983,N_17829);
and U22418 (N_22418,N_19198,N_19830);
or U22419 (N_22419,N_19512,N_19166);
and U22420 (N_22420,N_19588,N_18482);
or U22421 (N_22421,N_19390,N_17994);
or U22422 (N_22422,N_19771,N_17809);
xor U22423 (N_22423,N_17727,N_19868);
and U22424 (N_22424,N_19883,N_18038);
nand U22425 (N_22425,N_19547,N_18453);
or U22426 (N_22426,N_17732,N_17824);
and U22427 (N_22427,N_17505,N_19006);
or U22428 (N_22428,N_18328,N_18239);
nor U22429 (N_22429,N_18449,N_19486);
nor U22430 (N_22430,N_19815,N_18390);
and U22431 (N_22431,N_19154,N_19756);
or U22432 (N_22432,N_18515,N_18867);
nand U22433 (N_22433,N_18103,N_17929);
nand U22434 (N_22434,N_17692,N_18574);
nor U22435 (N_22435,N_18675,N_18029);
xnor U22436 (N_22436,N_17768,N_19389);
nor U22437 (N_22437,N_18848,N_17928);
xor U22438 (N_22438,N_19731,N_18127);
and U22439 (N_22439,N_18407,N_18512);
or U22440 (N_22440,N_17557,N_19092);
nor U22441 (N_22441,N_19901,N_19725);
or U22442 (N_22442,N_19065,N_19418);
nor U22443 (N_22443,N_17513,N_19166);
nand U22444 (N_22444,N_18980,N_19151);
or U22445 (N_22445,N_19138,N_18372);
nand U22446 (N_22446,N_17532,N_18614);
or U22447 (N_22447,N_19763,N_18839);
xnor U22448 (N_22448,N_17629,N_18931);
nand U22449 (N_22449,N_19682,N_19358);
nand U22450 (N_22450,N_18989,N_18596);
nand U22451 (N_22451,N_18039,N_18927);
and U22452 (N_22452,N_19524,N_19051);
nand U22453 (N_22453,N_17560,N_18468);
nor U22454 (N_22454,N_18986,N_17787);
nand U22455 (N_22455,N_19592,N_18176);
nor U22456 (N_22456,N_17869,N_19780);
nor U22457 (N_22457,N_18068,N_18770);
or U22458 (N_22458,N_19006,N_18841);
nor U22459 (N_22459,N_17735,N_17991);
or U22460 (N_22460,N_17702,N_18624);
nand U22461 (N_22461,N_19973,N_19078);
or U22462 (N_22462,N_18923,N_17732);
and U22463 (N_22463,N_19466,N_19326);
or U22464 (N_22464,N_18811,N_19161);
or U22465 (N_22465,N_18851,N_18753);
nor U22466 (N_22466,N_17810,N_19569);
nor U22467 (N_22467,N_18015,N_19119);
nor U22468 (N_22468,N_18597,N_18467);
nor U22469 (N_22469,N_19361,N_18920);
nor U22470 (N_22470,N_19773,N_19948);
nand U22471 (N_22471,N_19657,N_19910);
nand U22472 (N_22472,N_17649,N_19055);
nand U22473 (N_22473,N_19648,N_18661);
or U22474 (N_22474,N_17853,N_17952);
xor U22475 (N_22475,N_17691,N_18375);
and U22476 (N_22476,N_19526,N_18114);
nand U22477 (N_22477,N_18384,N_17899);
nor U22478 (N_22478,N_17544,N_17736);
nand U22479 (N_22479,N_18875,N_19357);
xnor U22480 (N_22480,N_18232,N_17849);
xnor U22481 (N_22481,N_17967,N_18073);
xnor U22482 (N_22482,N_19195,N_19897);
and U22483 (N_22483,N_19239,N_19369);
and U22484 (N_22484,N_18600,N_19987);
nor U22485 (N_22485,N_18013,N_19596);
xor U22486 (N_22486,N_19214,N_19027);
nand U22487 (N_22487,N_17828,N_18221);
or U22488 (N_22488,N_17587,N_17527);
nor U22489 (N_22489,N_17628,N_17796);
and U22490 (N_22490,N_18510,N_19224);
nor U22491 (N_22491,N_19148,N_19708);
or U22492 (N_22492,N_19244,N_19363);
or U22493 (N_22493,N_19649,N_17866);
xor U22494 (N_22494,N_19788,N_18742);
or U22495 (N_22495,N_19757,N_17599);
xor U22496 (N_22496,N_18839,N_17511);
or U22497 (N_22497,N_17718,N_18888);
xnor U22498 (N_22498,N_18599,N_19263);
nand U22499 (N_22499,N_18101,N_19899);
and U22500 (N_22500,N_20577,N_20129);
xor U22501 (N_22501,N_21380,N_21736);
and U22502 (N_22502,N_20218,N_20581);
xnor U22503 (N_22503,N_20001,N_21682);
nand U22504 (N_22504,N_21909,N_21841);
or U22505 (N_22505,N_20009,N_20529);
nand U22506 (N_22506,N_21735,N_20892);
xnor U22507 (N_22507,N_22297,N_21318);
nand U22508 (N_22508,N_20840,N_21052);
nor U22509 (N_22509,N_20962,N_20929);
and U22510 (N_22510,N_21045,N_22138);
nand U22511 (N_22511,N_21913,N_21410);
nand U22512 (N_22512,N_21604,N_20977);
and U22513 (N_22513,N_22038,N_22027);
xnor U22514 (N_22514,N_20028,N_21474);
or U22515 (N_22515,N_20361,N_21647);
nand U22516 (N_22516,N_22026,N_20660);
nand U22517 (N_22517,N_20592,N_22196);
nor U22518 (N_22518,N_20334,N_20704);
or U22519 (N_22519,N_20553,N_21070);
or U22520 (N_22520,N_20425,N_20494);
or U22521 (N_22521,N_20765,N_21681);
nor U22522 (N_22522,N_20923,N_21138);
nor U22523 (N_22523,N_21182,N_21870);
nor U22524 (N_22524,N_22085,N_22193);
xnor U22525 (N_22525,N_20434,N_20318);
xor U22526 (N_22526,N_20648,N_20042);
nand U22527 (N_22527,N_21499,N_22135);
and U22528 (N_22528,N_22343,N_22492);
or U22529 (N_22529,N_21373,N_20467);
and U22530 (N_22530,N_21446,N_20645);
nand U22531 (N_22531,N_22228,N_21547);
and U22532 (N_22532,N_20754,N_20774);
nand U22533 (N_22533,N_21825,N_22314);
and U22534 (N_22534,N_22336,N_22438);
and U22535 (N_22535,N_21588,N_20813);
nand U22536 (N_22536,N_21031,N_22452);
and U22537 (N_22537,N_21353,N_20498);
nand U22538 (N_22538,N_21814,N_21622);
nor U22539 (N_22539,N_21077,N_20811);
and U22540 (N_22540,N_21886,N_20300);
or U22541 (N_22541,N_22088,N_21765);
or U22542 (N_22542,N_21206,N_21450);
xnor U22543 (N_22543,N_22060,N_21256);
or U22544 (N_22544,N_21329,N_20513);
nand U22545 (N_22545,N_20210,N_22280);
nand U22546 (N_22546,N_20304,N_21720);
nand U22547 (N_22547,N_20053,N_20531);
xor U22548 (N_22548,N_22068,N_21012);
nor U22549 (N_22549,N_21295,N_20777);
xnor U22550 (N_22550,N_21107,N_21283);
and U22551 (N_22551,N_20082,N_20104);
and U22552 (N_22552,N_20688,N_22232);
xor U22553 (N_22553,N_21649,N_20446);
nand U22554 (N_22554,N_21459,N_20881);
and U22555 (N_22555,N_22041,N_22016);
nand U22556 (N_22556,N_22165,N_20794);
nand U22557 (N_22557,N_22414,N_20672);
or U22558 (N_22558,N_21974,N_20909);
or U22559 (N_22559,N_20181,N_20044);
xnor U22560 (N_22560,N_21756,N_21580);
nor U22561 (N_22561,N_21451,N_20297);
nor U22562 (N_22562,N_21927,N_20547);
or U22563 (N_22563,N_22058,N_21425);
nand U22564 (N_22564,N_20430,N_22428);
or U22565 (N_22565,N_20667,N_21670);
xnor U22566 (N_22566,N_21141,N_22052);
xor U22567 (N_22567,N_22001,N_21963);
nor U22568 (N_22568,N_20600,N_22406);
nand U22569 (N_22569,N_20429,N_20955);
xnor U22570 (N_22570,N_20359,N_20842);
xnor U22571 (N_22571,N_21265,N_21101);
and U22572 (N_22572,N_22344,N_20603);
and U22573 (N_22573,N_22277,N_21055);
nor U22574 (N_22574,N_21009,N_22104);
xnor U22575 (N_22575,N_20591,N_22474);
and U22576 (N_22576,N_20900,N_21395);
nor U22577 (N_22577,N_21934,N_20673);
and U22578 (N_22578,N_21457,N_20327);
and U22579 (N_22579,N_20311,N_20906);
nor U22580 (N_22580,N_21638,N_21312);
and U22581 (N_22581,N_21118,N_21019);
nor U22582 (N_22582,N_20993,N_21300);
nand U22583 (N_22583,N_21179,N_20098);
xnor U22584 (N_22584,N_20611,N_21452);
and U22585 (N_22585,N_22031,N_22323);
or U22586 (N_22586,N_21015,N_20081);
xor U22587 (N_22587,N_20431,N_20762);
nor U22588 (N_22588,N_21316,N_21067);
nor U22589 (N_22589,N_22212,N_21091);
xor U22590 (N_22590,N_20108,N_20134);
nor U22591 (N_22591,N_22442,N_22434);
or U22592 (N_22592,N_20230,N_20883);
and U22593 (N_22593,N_21247,N_21060);
xor U22594 (N_22594,N_20473,N_21117);
or U22595 (N_22595,N_22288,N_20199);
nand U22596 (N_22596,N_21990,N_21073);
nor U22597 (N_22597,N_21342,N_22171);
nand U22598 (N_22598,N_20781,N_20320);
or U22599 (N_22599,N_21630,N_21878);
nor U22600 (N_22600,N_20812,N_21786);
xnor U22601 (N_22601,N_20907,N_20661);
xor U22602 (N_22602,N_21520,N_21777);
or U22603 (N_22603,N_21359,N_20045);
nor U22604 (N_22604,N_20856,N_20882);
nand U22605 (N_22605,N_22412,N_21332);
or U22606 (N_22606,N_20666,N_21176);
and U22607 (N_22607,N_22271,N_21608);
nor U22608 (N_22608,N_20254,N_21656);
nand U22609 (N_22609,N_20072,N_22258);
xor U22610 (N_22610,N_21793,N_22380);
xor U22611 (N_22611,N_20367,N_21851);
nor U22612 (N_22612,N_20274,N_21954);
nand U22613 (N_22613,N_22285,N_22101);
nor U22614 (N_22614,N_21912,N_20036);
or U22615 (N_22615,N_22305,N_20744);
xnor U22616 (N_22616,N_21533,N_21360);
or U22617 (N_22617,N_21370,N_20202);
xnor U22618 (N_22618,N_22453,N_20634);
nor U22619 (N_22619,N_22313,N_20564);
or U22620 (N_22620,N_20100,N_20285);
xor U22621 (N_22621,N_22022,N_20890);
nor U22622 (N_22622,N_20951,N_22109);
nor U22623 (N_22623,N_21619,N_21253);
or U22624 (N_22624,N_20879,N_21394);
nor U22625 (N_22625,N_21086,N_22354);
nand U22626 (N_22626,N_20459,N_21613);
and U22627 (N_22627,N_21739,N_20133);
nand U22628 (N_22628,N_21609,N_22231);
and U22629 (N_22629,N_20049,N_20699);
and U22630 (N_22630,N_21578,N_21694);
xor U22631 (N_22631,N_22291,N_20269);
or U22632 (N_22632,N_21791,N_20166);
or U22633 (N_22633,N_20745,N_21099);
nand U22634 (N_22634,N_20983,N_21328);
and U22635 (N_22635,N_20286,N_21291);
or U22636 (N_22636,N_20959,N_22136);
xnor U22637 (N_22637,N_20864,N_20270);
xnor U22638 (N_22638,N_21530,N_21235);
or U22639 (N_22639,N_20272,N_20313);
xnor U22640 (N_22640,N_20821,N_20557);
or U22641 (N_22641,N_22451,N_20556);
and U22642 (N_22642,N_20610,N_21354);
nor U22643 (N_22643,N_22437,N_20022);
and U22644 (N_22644,N_22098,N_20719);
nor U22645 (N_22645,N_20299,N_21333);
xnor U22646 (N_22646,N_21460,N_20417);
and U22647 (N_22647,N_20364,N_20120);
nand U22648 (N_22648,N_21476,N_22011);
or U22649 (N_22649,N_20213,N_20469);
or U22650 (N_22650,N_20766,N_22373);
xnor U22651 (N_22651,N_21174,N_20362);
xnor U22652 (N_22652,N_20623,N_21819);
nor U22653 (N_22653,N_20308,N_22301);
and U22654 (N_22654,N_21445,N_21541);
or U22655 (N_22655,N_22478,N_21136);
and U22656 (N_22656,N_21214,N_20388);
and U22657 (N_22657,N_21033,N_20889);
xor U22658 (N_22658,N_21614,N_20348);
nor U22659 (N_22659,N_22468,N_21740);
and U22660 (N_22660,N_21782,N_20246);
xnor U22661 (N_22661,N_22126,N_22421);
xor U22662 (N_22662,N_20898,N_21896);
xnor U22663 (N_22663,N_21434,N_21687);
and U22664 (N_22664,N_22218,N_21148);
and U22665 (N_22665,N_20323,N_22097);
and U22666 (N_22666,N_20208,N_20708);
nand U22667 (N_22667,N_21339,N_20152);
nor U22668 (N_22668,N_21241,N_22309);
or U22669 (N_22669,N_20078,N_20131);
or U22670 (N_22670,N_21779,N_20891);
nor U22671 (N_22671,N_21254,N_21942);
xor U22672 (N_22672,N_20160,N_21728);
nand U22673 (N_22673,N_21723,N_21673);
nand U22674 (N_22674,N_22195,N_22310);
and U22675 (N_22675,N_21566,N_20852);
nand U22676 (N_22676,N_20482,N_22164);
or U22677 (N_22677,N_21659,N_22008);
and U22678 (N_22678,N_22348,N_21442);
nand U22679 (N_22679,N_21243,N_22071);
and U22680 (N_22680,N_21481,N_22418);
nor U22681 (N_22681,N_22176,N_21496);
xor U22682 (N_22682,N_22106,N_20717);
and U22683 (N_22683,N_21518,N_22062);
nor U22684 (N_22684,N_20893,N_20665);
or U22685 (N_22685,N_22485,N_20390);
nor U22686 (N_22686,N_21879,N_20669);
nand U22687 (N_22687,N_21775,N_21586);
or U22688 (N_22688,N_21192,N_20468);
nor U22689 (N_22689,N_20488,N_21207);
or U22690 (N_22690,N_21422,N_20822);
or U22691 (N_22691,N_20394,N_20176);
xor U22692 (N_22692,N_20055,N_20989);
nor U22693 (N_22693,N_21095,N_20032);
xor U22694 (N_22694,N_22172,N_20377);
xor U22695 (N_22695,N_20229,N_22283);
nor U22696 (N_22696,N_21358,N_20143);
nand U22697 (N_22697,N_22167,N_20451);
xor U22698 (N_22698,N_21710,N_20373);
nand U22699 (N_22699,N_21552,N_20271);
xnor U22700 (N_22700,N_20601,N_20521);
nand U22701 (N_22701,N_20150,N_21123);
and U22702 (N_22702,N_22214,N_21028);
nor U22703 (N_22703,N_20408,N_20355);
or U22704 (N_22704,N_21323,N_20105);
xor U22705 (N_22705,N_20743,N_22411);
nand U22706 (N_22706,N_22099,N_21575);
and U22707 (N_22707,N_20858,N_20870);
nand U22708 (N_22708,N_22180,N_20985);
xor U22709 (N_22709,N_20259,N_22252);
xor U22710 (N_22710,N_21036,N_20153);
xor U22711 (N_22711,N_21041,N_22043);
xor U22712 (N_22712,N_21596,N_21688);
xor U22713 (N_22713,N_22364,N_21536);
or U22714 (N_22714,N_22251,N_20282);
nor U22715 (N_22715,N_21577,N_21257);
or U22716 (N_22716,N_20051,N_20728);
and U22717 (N_22717,N_20800,N_20792);
nor U22718 (N_22718,N_20747,N_21967);
xnor U22719 (N_22719,N_22381,N_21737);
xor U22720 (N_22720,N_22037,N_21936);
nor U22721 (N_22721,N_20445,N_20470);
or U22722 (N_22722,N_21309,N_21859);
or U22723 (N_22723,N_20426,N_20647);
xnor U22724 (N_22724,N_21832,N_21803);
and U22725 (N_22725,N_21306,N_20530);
and U22726 (N_22726,N_21854,N_21845);
nand U22727 (N_22727,N_22239,N_21054);
and U22728 (N_22728,N_21898,N_21755);
nor U22729 (N_22729,N_21984,N_20604);
nand U22730 (N_22730,N_21806,N_21471);
or U22731 (N_22731,N_20074,N_22307);
and U22732 (N_22732,N_20077,N_21116);
nand U22733 (N_22733,N_21004,N_20808);
or U22734 (N_22734,N_20216,N_22467);
and U22735 (N_22735,N_22465,N_20768);
or U22736 (N_22736,N_22202,N_20056);
and U22737 (N_22737,N_20412,N_22420);
and U22738 (N_22738,N_21121,N_20099);
nand U22739 (N_22739,N_20795,N_21925);
xor U22740 (N_22740,N_21502,N_21559);
nand U22741 (N_22741,N_20837,N_20371);
or U22742 (N_22742,N_22475,N_20796);
xor U22743 (N_22743,N_20292,N_21260);
nor U22744 (N_22744,N_21715,N_21140);
nor U22745 (N_22745,N_20294,N_20903);
or U22746 (N_22746,N_20515,N_21556);
nor U22747 (N_22747,N_21891,N_21464);
nand U22748 (N_22748,N_20861,N_20155);
nand U22749 (N_22749,N_20884,N_20386);
nand U22750 (N_22750,N_22227,N_21341);
nor U22751 (N_22751,N_21821,N_20170);
and U22752 (N_22752,N_21708,N_22042);
xor U22753 (N_22753,N_21709,N_21027);
nand U22754 (N_22754,N_21824,N_21108);
xnor U22755 (N_22755,N_22394,N_21144);
or U22756 (N_22756,N_21155,N_21805);
and U22757 (N_22757,N_20917,N_21510);
and U22758 (N_22758,N_21551,N_21043);
and U22759 (N_22759,N_20875,N_21945);
nor U22760 (N_22760,N_21846,N_20999);
or U22761 (N_22761,N_20162,N_21753);
nand U22762 (N_22762,N_21109,N_20751);
and U22763 (N_22763,N_21096,N_20366);
nor U22764 (N_22764,N_21853,N_22372);
xnor U22765 (N_22765,N_20406,N_21635);
xnor U22766 (N_22766,N_21920,N_22400);
xnor U22767 (N_22767,N_20310,N_22413);
nor U22768 (N_22768,N_20514,N_22132);
or U22769 (N_22769,N_22386,N_21959);
nor U22770 (N_22770,N_20849,N_20065);
or U22771 (N_22771,N_20102,N_20476);
xnor U22772 (N_22772,N_21906,N_22090);
and U22773 (N_22773,N_20084,N_20646);
nor U22774 (N_22774,N_21218,N_20025);
and U22775 (N_22775,N_20433,N_21553);
xor U22776 (N_22776,N_22112,N_20125);
xor U22777 (N_22777,N_21584,N_20877);
xnor U22778 (N_22778,N_21587,N_22130);
or U22779 (N_22779,N_20350,N_20635);
and U22780 (N_22780,N_20097,N_21669);
nor U22781 (N_22781,N_20141,N_21336);
and U22782 (N_22782,N_20670,N_20071);
or U22783 (N_22783,N_22255,N_21432);
nor U22784 (N_22784,N_21868,N_21075);
or U22785 (N_22785,N_21980,N_20041);
nand U22786 (N_22786,N_21381,N_22382);
and U22787 (N_22787,N_20659,N_22084);
and U22788 (N_22788,N_22279,N_20260);
and U22789 (N_22789,N_21162,N_20438);
and U22790 (N_22790,N_20011,N_21124);
and U22791 (N_22791,N_22377,N_22319);
nor U22792 (N_22792,N_20954,N_22312);
and U22793 (N_22793,N_21883,N_20561);
or U22794 (N_22794,N_20804,N_21711);
nor U22795 (N_22795,N_20620,N_21978);
and U22796 (N_22796,N_20154,N_21529);
nor U22797 (N_22797,N_20772,N_22150);
nor U22798 (N_22798,N_20679,N_20926);
xor U22799 (N_22799,N_21494,N_21897);
or U22800 (N_22800,N_21595,N_21001);
nor U22801 (N_22801,N_21764,N_21674);
or U22802 (N_22802,N_21910,N_21335);
nand U22803 (N_22803,N_20157,N_21382);
xnor U22804 (N_22804,N_20324,N_20033);
nor U22805 (N_22805,N_21693,N_21372);
nand U22806 (N_22806,N_21125,N_20958);
or U22807 (N_22807,N_21215,N_20135);
nor U22808 (N_22808,N_20465,N_21221);
xnor U22809 (N_22809,N_20136,N_22148);
or U22810 (N_22810,N_21119,N_21479);
xnor U22811 (N_22811,N_20060,N_20655);
xnor U22812 (N_22812,N_20554,N_21849);
or U22813 (N_22813,N_20683,N_21894);
and U22814 (N_22814,N_20625,N_21960);
and U22815 (N_22815,N_22267,N_20585);
nor U22816 (N_22816,N_20549,N_20110);
and U22817 (N_22817,N_22069,N_22229);
or U22818 (N_22818,N_20880,N_20351);
xor U22819 (N_22819,N_20826,N_20988);
or U22820 (N_22820,N_21789,N_20798);
nand U22821 (N_22821,N_21792,N_21597);
nand U22822 (N_22822,N_20574,N_22222);
xor U22823 (N_22823,N_21524,N_21620);
and U22824 (N_22824,N_21734,N_20247);
and U22825 (N_22825,N_20705,N_20191);
nand U22826 (N_22826,N_22054,N_20690);
nor U22827 (N_22827,N_21396,N_20061);
nand U22828 (N_22828,N_20702,N_22146);
or U22829 (N_22829,N_20998,N_21000);
nand U22830 (N_22830,N_21126,N_21132);
or U22831 (N_22831,N_20922,N_22487);
nor U22832 (N_22832,N_20005,N_20908);
nor U22833 (N_22833,N_22094,N_21863);
nor U22834 (N_22834,N_20018,N_20040);
or U22835 (N_22835,N_21969,N_20149);
and U22836 (N_22836,N_20587,N_22157);
or U22837 (N_22837,N_21486,N_20689);
nor U22838 (N_22838,N_21563,N_20048);
nor U22839 (N_22839,N_20178,N_22213);
xor U22840 (N_22840,N_21292,N_21252);
and U22841 (N_22841,N_20478,N_20818);
and U22842 (N_22842,N_21852,N_20663);
and U22843 (N_22843,N_21817,N_21271);
and U22844 (N_22844,N_20642,N_20085);
nor U22845 (N_22845,N_21818,N_21829);
nand U22846 (N_22846,N_20037,N_22378);
nor U22847 (N_22847,N_22431,N_20267);
nand U22848 (N_22848,N_21873,N_21637);
or U22849 (N_22849,N_20961,N_22224);
or U22850 (N_22850,N_21187,N_22324);
and U22851 (N_22851,N_20714,N_22159);
nor U22852 (N_22852,N_20671,N_22115);
or U22853 (N_22853,N_20725,N_20523);
and U22854 (N_22854,N_21287,N_22466);
xor U22855 (N_22855,N_20944,N_20677);
or U22856 (N_22856,N_22100,N_20896);
or U22857 (N_22857,N_22489,N_21196);
or U22858 (N_22858,N_22091,N_21475);
xnor U22859 (N_22859,N_21895,N_21188);
nand U22860 (N_22860,N_20746,N_21134);
nor U22861 (N_22861,N_21634,N_20385);
and U22862 (N_22862,N_22429,N_20769);
and U22863 (N_22863,N_21881,N_20692);
nand U22864 (N_22864,N_21268,N_20797);
or U22865 (N_22865,N_20629,N_21893);
and U22866 (N_22866,N_21083,N_22419);
and U22867 (N_22867,N_20615,N_21244);
xor U22868 (N_22868,N_21010,N_22326);
or U22869 (N_22869,N_20967,N_21800);
and U22870 (N_22870,N_22342,N_21992);
and U22871 (N_22871,N_21228,N_22347);
nor U22872 (N_22872,N_20636,N_21810);
or U22873 (N_22873,N_20779,N_21049);
and U22874 (N_22874,N_20475,N_22220);
xnor U22875 (N_22875,N_20164,N_21546);
and U22876 (N_22876,N_20584,N_21506);
or U22877 (N_22877,N_20707,N_20314);
or U22878 (N_22878,N_21568,N_20833);
nor U22879 (N_22879,N_20114,N_21515);
xor U22880 (N_22880,N_20730,N_20376);
xnor U22881 (N_22881,N_21864,N_20978);
nor U22882 (N_22882,N_21828,N_20123);
nor U22883 (N_22883,N_21362,N_20532);
nand U22884 (N_22884,N_21098,N_21477);
xnor U22885 (N_22885,N_21466,N_22033);
xnor U22886 (N_22886,N_21406,N_21264);
or U22887 (N_22887,N_21717,N_21219);
xor U22888 (N_22888,N_20863,N_20328);
and U22889 (N_22889,N_21538,N_20681);
or U22890 (N_22890,N_20484,N_22483);
or U22891 (N_22891,N_22120,N_21962);
xnor U22892 (N_22892,N_21512,N_20325);
nor U22893 (N_22893,N_21478,N_20767);
nor U22894 (N_22894,N_20653,N_22029);
or U22895 (N_22895,N_21463,N_20510);
nor U22896 (N_22896,N_20541,N_20843);
nor U22897 (N_22897,N_22404,N_22108);
and U22898 (N_22898,N_20450,N_21650);
nor U22899 (N_22899,N_20474,N_22484);
or U22900 (N_22900,N_22238,N_21748);
xnor U22901 (N_22901,N_21589,N_21885);
nor U22902 (N_22902,N_20773,N_21663);
xor U22903 (N_22903,N_20215,N_20219);
xor U22904 (N_22904,N_20546,N_22306);
or U22905 (N_22905,N_22278,N_20419);
or U22906 (N_22906,N_21198,N_21289);
and U22907 (N_22907,N_20619,N_21042);
nand U22908 (N_22908,N_21495,N_22082);
and U22909 (N_22909,N_22092,N_20609);
and U22910 (N_22910,N_20887,N_21263);
xnor U22911 (N_22911,N_22446,N_20369);
xor U22912 (N_22912,N_20997,N_21002);
nand U22913 (N_22913,N_20248,N_22236);
and U22914 (N_22914,N_20301,N_21473);
xnor U22915 (N_22915,N_20543,N_20685);
xor U22916 (N_22916,N_21497,N_21628);
xor U22917 (N_22917,N_22166,N_21351);
and U22918 (N_22918,N_20046,N_22175);
or U22919 (N_22919,N_22287,N_20396);
nand U22920 (N_22920,N_21298,N_20206);
and U22921 (N_22921,N_21046,N_21716);
xnor U22922 (N_22922,N_22013,N_20456);
xnor U22923 (N_22923,N_20780,N_22367);
xor U22924 (N_22924,N_21581,N_21923);
and U22925 (N_22925,N_21714,N_20158);
xnor U22926 (N_22926,N_21816,N_21697);
and U22927 (N_22927,N_22203,N_22253);
nor U22928 (N_22928,N_20872,N_22034);
or U22929 (N_22929,N_21472,N_21456);
or U22930 (N_22930,N_20168,N_20365);
xnor U22931 (N_22931,N_22294,N_22044);
nor U22932 (N_22932,N_21030,N_21783);
nand U22933 (N_22933,N_22331,N_21607);
and U22934 (N_22934,N_20461,N_20742);
nor U22935 (N_22935,N_22012,N_20816);
xnor U22936 (N_22936,N_22030,N_20857);
nand U22937 (N_22937,N_21937,N_21641);
nand U22938 (N_22938,N_21742,N_20502);
and U22939 (N_22939,N_21233,N_20241);
nand U22940 (N_22940,N_21461,N_21744);
and U22941 (N_22941,N_20920,N_21114);
xnor U22942 (N_22942,N_22245,N_21409);
or U22943 (N_22943,N_21350,N_20536);
and U22944 (N_22944,N_22260,N_21498);
nor U22945 (N_22945,N_21149,N_22035);
nor U22946 (N_22946,N_20643,N_20976);
xnor U22947 (N_22947,N_21880,N_20913);
nor U22948 (N_22948,N_21593,N_21013);
or U22949 (N_22949,N_21245,N_22444);
and U22950 (N_22950,N_20522,N_22237);
nor U22951 (N_22951,N_20678,N_20177);
xnor U22952 (N_22952,N_20566,N_22028);
nor U22953 (N_22953,N_20187,N_22308);
and U22954 (N_22954,N_21848,N_20752);
xnor U22955 (N_22955,N_21801,N_21542);
nand U22956 (N_22956,N_22241,N_21008);
and U22957 (N_22957,N_20198,N_20126);
and U22958 (N_22958,N_20664,N_22210);
nor U22959 (N_22959,N_21211,N_21195);
nand U22960 (N_22960,N_21385,N_20483);
nor U22961 (N_22961,N_22185,N_20088);
nor U22962 (N_22962,N_20627,N_21110);
and U22963 (N_22963,N_21066,N_20223);
xor U22964 (N_22964,N_21904,N_20256);
and U22965 (N_22965,N_20021,N_21751);
nor U22966 (N_22966,N_21860,N_21725);
xor U22967 (N_22967,N_21743,N_22254);
nor U22968 (N_22968,N_21976,N_21501);
nand U22969 (N_22969,N_20638,N_21051);
nor U22970 (N_22970,N_22074,N_20945);
nand U22971 (N_22971,N_21201,N_21706);
xnor U22972 (N_22972,N_22114,N_20594);
and U22973 (N_22973,N_20321,N_20287);
nand U22974 (N_22974,N_21150,N_22334);
or U22975 (N_22975,N_20694,N_20031);
nand U22976 (N_22976,N_21651,N_20791);
nand U22977 (N_22977,N_21965,N_22477);
nor U22978 (N_22978,N_20240,N_20375);
or U22979 (N_22979,N_20137,N_20266);
and U22980 (N_22980,N_20545,N_20731);
and U22981 (N_22981,N_21319,N_21284);
nand U22982 (N_22982,N_22234,N_22168);
nor U22983 (N_22983,N_20517,N_21642);
nor U22984 (N_22984,N_22072,N_22118);
or U22985 (N_22985,N_22204,N_20016);
and U22986 (N_22986,N_20721,N_21662);
or U22987 (N_22987,N_20356,N_20535);
nor U22988 (N_22988,N_20576,N_20111);
xor U22989 (N_22989,N_20302,N_20966);
nor U22990 (N_22990,N_22405,N_20613);
nor U22991 (N_22991,N_21003,N_22458);
xnor U22992 (N_22992,N_21203,N_20934);
or U22993 (N_22993,N_20251,N_22360);
nand U22994 (N_22994,N_20866,N_21946);
xor U22995 (N_22995,N_20075,N_20802);
nand U22996 (N_22996,N_20212,N_22263);
nor U22997 (N_22997,N_21212,N_20886);
nand U22998 (N_22998,N_22350,N_21624);
and U22999 (N_22999,N_20119,N_22407);
xnor U23000 (N_23000,N_22415,N_20221);
or U23001 (N_23001,N_21334,N_21441);
xnor U23002 (N_23002,N_20736,N_22087);
nor U23003 (N_23003,N_21059,N_20495);
and U23004 (N_23004,N_22445,N_21420);
nor U23005 (N_23005,N_21240,N_20398);
nor U23006 (N_23006,N_21857,N_20607);
and U23007 (N_23007,N_20440,N_22051);
nand U23008 (N_23008,N_20165,N_22143);
nand U23009 (N_23009,N_21557,N_21683);
and U23010 (N_23010,N_20552,N_20740);
xnor U23011 (N_23011,N_20783,N_22395);
nor U23012 (N_23012,N_20622,N_21151);
xnor U23013 (N_23013,N_21161,N_22303);
xor U23014 (N_23014,N_20015,N_20651);
nor U23015 (N_23015,N_22351,N_20253);
nand U23016 (N_23016,N_21229,N_20404);
or U23017 (N_23017,N_20234,N_21190);
or U23018 (N_23018,N_22206,N_22048);
xor U23019 (N_23019,N_21238,N_20173);
xnor U23020 (N_23020,N_20828,N_20293);
xor U23021 (N_23021,N_20466,N_20534);
or U23022 (N_23022,N_20511,N_22470);
xor U23023 (N_23023,N_20374,N_21331);
nor U23024 (N_23024,N_21811,N_21636);
xor U23025 (N_23025,N_20941,N_21443);
and U23026 (N_23026,N_22289,N_20414);
nand U23027 (N_23027,N_21482,N_21266);
and U23028 (N_23028,N_20012,N_21167);
and U23029 (N_23029,N_20087,N_20194);
nor U23030 (N_23030,N_21407,N_21752);
nand U23031 (N_23031,N_22261,N_20986);
xor U23032 (N_23032,N_20668,N_21402);
or U23033 (N_23033,N_20393,N_21591);
nand U23034 (N_23034,N_21809,N_20010);
nor U23035 (N_23035,N_21692,N_22399);
nor U23036 (N_23036,N_20039,N_21367);
nor U23037 (N_23037,N_20481,N_21202);
or U23038 (N_23038,N_22004,N_20217);
nor U23039 (N_23039,N_21889,N_21232);
and U23040 (N_23040,N_20338,N_22329);
or U23041 (N_23041,N_22003,N_21509);
nand U23042 (N_23042,N_20641,N_22436);
nand U23043 (N_23043,N_20539,N_20733);
xor U23044 (N_23044,N_21166,N_20298);
nor U23045 (N_23045,N_20453,N_20151);
and U23046 (N_23046,N_21991,N_22223);
or U23047 (N_23047,N_20598,N_21135);
nor U23048 (N_23048,N_21986,N_20499);
xnor U23049 (N_23049,N_21955,N_21901);
xor U23050 (N_23050,N_21772,N_20370);
nor U23051 (N_23051,N_21325,N_21177);
xor U23052 (N_23052,N_21778,N_22425);
xor U23053 (N_23053,N_21184,N_22113);
xnor U23054 (N_23054,N_20487,N_20841);
xor U23055 (N_23055,N_21774,N_21153);
nand U23056 (N_23056,N_22457,N_20096);
nand U23057 (N_23057,N_22243,N_21677);
and U23058 (N_23058,N_21388,N_21217);
xnor U23059 (N_23059,N_21199,N_21914);
or U23060 (N_23060,N_21251,N_21672);
and U23061 (N_23061,N_20953,N_20947);
nand U23062 (N_23062,N_21280,N_20086);
xor U23063 (N_23063,N_21754,N_21200);
or U23064 (N_23064,N_21983,N_21102);
nand U23065 (N_23065,N_21771,N_21550);
xor U23066 (N_23066,N_21820,N_22219);
or U23067 (N_23067,N_22361,N_20871);
nor U23068 (N_23068,N_20252,N_21269);
or U23069 (N_23069,N_20427,N_21944);
xor U23070 (N_23070,N_22182,N_21892);
nand U23071 (N_23071,N_22345,N_21865);
and U23072 (N_23072,N_21761,N_21639);
xor U23073 (N_23073,N_22341,N_20332);
nor U23074 (N_23074,N_20512,N_21837);
nand U23075 (N_23075,N_21666,N_21576);
nand U23076 (N_23076,N_21194,N_21802);
and U23077 (N_23077,N_21917,N_20054);
xnor U23078 (N_23078,N_20211,N_21320);
and U23079 (N_23079,N_21977,N_21696);
and U23080 (N_23080,N_22005,N_22123);
nor U23081 (N_23081,N_20333,N_22387);
nand U23082 (N_23082,N_21979,N_20058);
nor U23083 (N_23083,N_21209,N_20537);
nand U23084 (N_23084,N_21741,N_20491);
and U23085 (N_23085,N_20995,N_20258);
xnor U23086 (N_23086,N_20336,N_20876);
nand U23087 (N_23087,N_21259,N_20027);
xor U23088 (N_23088,N_21667,N_21302);
nor U23089 (N_23089,N_20277,N_20528);
nand U23090 (N_23090,N_21590,N_22482);
xnor U23091 (N_23091,N_21064,N_21713);
nand U23092 (N_23092,N_20930,N_22246);
nand U23093 (N_23093,N_21862,N_22353);
and U23094 (N_23094,N_20633,N_20847);
and U23095 (N_23095,N_20914,N_20326);
or U23096 (N_23096,N_20146,N_20910);
nand U23097 (N_23097,N_20583,N_22276);
and U23098 (N_23098,N_22472,N_21392);
and U23099 (N_23099,N_20068,N_21794);
and U23100 (N_23100,N_21226,N_22298);
and U23101 (N_23101,N_20250,N_20987);
nor U23102 (N_23102,N_20919,N_21299);
and U23103 (N_23103,N_22036,N_20720);
xnor U23104 (N_23104,N_21627,N_21258);
or U23105 (N_23105,N_22019,N_20693);
or U23106 (N_23106,N_20614,N_20589);
and U23107 (N_23107,N_21830,N_20948);
nand U23108 (N_23108,N_21902,N_22275);
xnor U23109 (N_23109,N_20503,N_21534);
and U23110 (N_23110,N_22186,N_20464);
nand U23111 (N_23111,N_22107,N_21267);
nor U23112 (N_23112,N_21807,N_21159);
nor U23113 (N_23113,N_21480,N_21447);
xnor U23114 (N_23114,N_20138,N_21931);
nand U23115 (N_23115,N_22391,N_21007);
xor U23116 (N_23116,N_22017,N_22075);
and U23117 (N_23117,N_21038,N_21032);
nor U23118 (N_23118,N_21170,N_21554);
and U23119 (N_23119,N_21998,N_22128);
nand U23120 (N_23120,N_20019,N_21703);
or U23121 (N_23121,N_20381,N_20089);
or U23122 (N_23122,N_20582,N_21301);
or U23123 (N_23123,N_20706,N_22163);
or U23124 (N_23124,N_20263,N_21952);
xor U23125 (N_23125,N_22142,N_21103);
or U23126 (N_23126,N_20268,N_21605);
nor U23127 (N_23127,N_20479,N_21888);
nand U23128 (N_23128,N_21623,N_20389);
and U23129 (N_23129,N_21058,N_21872);
nand U23130 (N_23130,N_21664,N_22462);
nor U23131 (N_23131,N_22281,N_20764);
xnor U23132 (N_23132,N_22032,N_21652);
or U23133 (N_23133,N_21842,N_20824);
nand U23134 (N_23134,N_20749,N_20755);
and U23135 (N_23135,N_21561,N_21433);
nor U23136 (N_23136,N_20288,N_22295);
nor U23137 (N_23137,N_21645,N_22173);
nor U23138 (N_23138,N_21866,N_21618);
xnor U23139 (N_23139,N_20563,N_21970);
nor U23140 (N_23140,N_20691,N_20597);
nor U23141 (N_23141,N_21758,N_21448);
nor U23142 (N_23142,N_20276,N_21834);
nand U23143 (N_23143,N_21053,N_20063);
and U23144 (N_23144,N_21485,N_20630);
xnor U23145 (N_23145,N_21376,N_22476);
xnor U23146 (N_23146,N_21957,N_21242);
and U23147 (N_23147,N_22131,N_22355);
nand U23148 (N_23148,N_20992,N_21361);
and U23149 (N_23149,N_20257,N_20172);
and U23150 (N_23150,N_20095,N_21890);
xor U23151 (N_23151,N_21427,N_20423);
xnor U23152 (N_23152,N_20675,N_21080);
nor U23153 (N_23153,N_20454,N_20565);
and U23154 (N_23154,N_21186,N_20608);
xnor U23155 (N_23155,N_20312,N_21185);
or U23156 (N_23156,N_20652,N_22264);
nand U23157 (N_23157,N_20008,N_21569);
or U23158 (N_23158,N_22486,N_20912);
nand U23159 (N_23159,N_21327,N_21784);
nor U23160 (N_23160,N_21523,N_21078);
or U23161 (N_23161,N_21062,N_20569);
xnor U23162 (N_23162,N_21056,N_22014);
nor U23163 (N_23163,N_21469,N_21173);
nand U23164 (N_23164,N_21018,N_21436);
nand U23165 (N_23165,N_21788,N_21317);
or U23166 (N_23166,N_20189,N_20859);
and U23167 (N_23167,N_21843,N_20595);
nor U23168 (N_23168,N_22181,N_21171);
nand U23169 (N_23169,N_21956,N_21532);
xnor U23170 (N_23170,N_20209,N_20497);
and U23171 (N_23171,N_21668,N_21705);
xor U23172 (N_23172,N_20562,N_22063);
nand U23173 (N_23173,N_21330,N_21612);
nor U23174 (N_23174,N_21130,N_20785);
nand U23175 (N_23175,N_22250,N_20701);
or U23176 (N_23176,N_20145,N_20835);
xnor U23177 (N_23177,N_21163,N_21374);
nor U23178 (N_23178,N_20723,N_22449);
or U23179 (N_23179,N_21437,N_21763);
nand U23180 (N_23180,N_20070,N_21371);
and U23181 (N_23181,N_21521,N_20410);
xor U23182 (N_23182,N_22338,N_21296);
xor U23183 (N_23183,N_21648,N_21505);
and U23184 (N_23184,N_21850,N_21449);
nand U23185 (N_23185,N_20303,N_21246);
nand U23186 (N_23186,N_20091,N_21543);
and U23187 (N_23187,N_20939,N_21522);
nand U23188 (N_23188,N_22145,N_20411);
or U23189 (N_23189,N_21384,N_21766);
xor U23190 (N_23190,N_21704,N_21164);
and U23191 (N_23191,N_21231,N_21024);
nor U23192 (N_23192,N_21653,N_20486);
nand U23193 (N_23193,N_22282,N_20850);
and U23194 (N_23194,N_20232,N_20624);
nand U23195 (N_23195,N_20965,N_22257);
nor U23196 (N_23196,N_22495,N_20413);
nand U23197 (N_23197,N_20378,N_20382);
and U23198 (N_23198,N_21017,N_21113);
or U23199 (N_23199,N_21285,N_21719);
nor U23200 (N_23200,N_21785,N_21104);
or U23201 (N_23201,N_20422,N_22357);
or U23202 (N_23202,N_22249,N_20757);
xnor U23203 (N_23203,N_22156,N_20349);
xnor U23204 (N_23204,N_22293,N_21465);
nor U23205 (N_23205,N_22169,N_20567);
or U23206 (N_23206,N_20860,N_21290);
nand U23207 (N_23207,N_21592,N_20076);
or U23208 (N_23208,N_20750,N_22117);
and U23209 (N_23209,N_20231,N_21029);
or U23210 (N_23210,N_20810,N_20420);
or U23211 (N_23211,N_21903,N_20339);
nand U23212 (N_23212,N_20975,N_22317);
and U23213 (N_23213,N_20463,N_20727);
xnor U23214 (N_23214,N_21129,N_20825);
nand U23215 (N_23215,N_21462,N_21583);
xnor U23216 (N_23216,N_20969,N_21982);
or U23217 (N_23217,N_20829,N_20342);
or U23218 (N_23218,N_20806,N_21087);
or U23219 (N_23219,N_21308,N_21397);
or U23220 (N_23220,N_21326,N_21143);
nor U23221 (N_23221,N_22435,N_22299);
nor U23222 (N_23222,N_21508,N_20973);
and U23223 (N_23223,N_21695,N_21665);
or U23224 (N_23224,N_21943,N_22006);
nand U23225 (N_23225,N_20379,N_22337);
nor U23226 (N_23226,N_22359,N_22315);
nor U23227 (N_23227,N_22497,N_20776);
and U23228 (N_23228,N_22392,N_20343);
nor U23229 (N_23229,N_20280,N_21759);
nor U23230 (N_23230,N_21796,N_21127);
xnor U23231 (N_23231,N_22356,N_21421);
and U23232 (N_23232,N_20399,N_20204);
and U23233 (N_23233,N_22388,N_20265);
xnor U23234 (N_23234,N_20026,N_20904);
and U23235 (N_23235,N_21631,N_21646);
nor U23236 (N_23236,N_21154,N_21152);
or U23237 (N_23237,N_20237,N_21403);
or U23238 (N_23238,N_21429,N_22021);
nand U23239 (N_23239,N_20586,N_22247);
or U23240 (N_23240,N_21389,N_20606);
or U23241 (N_23241,N_20275,N_20803);
nor U23242 (N_23242,N_21369,N_22040);
nand U23243 (N_23243,N_21678,N_22339);
or U23244 (N_23244,N_21453,N_22368);
or U23245 (N_23245,N_20296,N_21994);
nand U23246 (N_23246,N_21718,N_21511);
xor U23247 (N_23247,N_21020,N_21676);
and U23248 (N_23248,N_21549,N_21224);
nand U23249 (N_23249,N_21707,N_22205);
or U23250 (N_23250,N_22333,N_21364);
or U23251 (N_23251,N_21050,N_20402);
xnor U23252 (N_23252,N_20200,N_22144);
nor U23253 (N_23253,N_21571,N_22369);
or U23254 (N_23254,N_20580,N_21900);
nor U23255 (N_23255,N_21958,N_20942);
or U23256 (N_23256,N_21489,N_21230);
nor U23257 (N_23257,N_21025,N_20435);
nor U23258 (N_23258,N_22493,N_21349);
xnor U23259 (N_23259,N_21517,N_21137);
and U23260 (N_23260,N_22189,N_21540);
nor U23261 (N_23261,N_21216,N_22061);
and U23262 (N_23262,N_21527,N_21798);
or U23263 (N_23263,N_22056,N_21833);
or U23264 (N_23264,N_22015,N_21249);
nand U23265 (N_23265,N_22322,N_20222);
or U23266 (N_23266,N_20330,N_20935);
and U23267 (N_23267,N_21005,N_21691);
nand U23268 (N_23268,N_21236,N_20617);
or U23269 (N_23269,N_21823,N_20703);
or U23270 (N_23270,N_20169,N_21699);
or U23271 (N_23271,N_21321,N_20496);
nand U23272 (N_23272,N_21131,N_21181);
nor U23273 (N_23273,N_21921,N_21822);
and U23274 (N_23274,N_22443,N_21911);
or U23275 (N_23275,N_21191,N_20621);
or U23276 (N_23276,N_20401,N_21011);
nand U23277 (N_23277,N_22093,N_20193);
xor U23278 (N_23278,N_20855,N_21128);
xnor U23279 (N_23279,N_20972,N_21686);
and U23280 (N_23280,N_22340,N_21640);
or U23281 (N_23281,N_21492,N_20090);
or U23282 (N_23282,N_22498,N_21156);
nor U23283 (N_23283,N_21602,N_21386);
or U23284 (N_23284,N_20830,N_20639);
nor U23285 (N_23285,N_22174,N_22240);
nand U23286 (N_23286,N_21572,N_22045);
and U23287 (N_23287,N_20943,N_21072);
or U23288 (N_23288,N_20674,N_21262);
nor U23289 (N_23289,N_20124,N_20322);
or U23290 (N_23290,N_21223,N_20013);
nor U23291 (N_23291,N_21724,N_20452);
or U23292 (N_23292,N_22200,N_20784);
nor U23293 (N_23293,N_21120,N_20729);
nand U23294 (N_23294,N_21074,N_20748);
nor U23295 (N_23295,N_20605,N_20017);
nand U23296 (N_23296,N_21769,N_22430);
xnor U23297 (N_23297,N_22208,N_21874);
nor U23298 (N_23298,N_20109,N_21276);
nand U23299 (N_23299,N_20233,N_21303);
xor U23300 (N_23300,N_21685,N_21180);
or U23301 (N_23301,N_22393,N_20925);
and U23302 (N_23302,N_20968,N_22262);
nor U23303 (N_23303,N_21006,N_20067);
nor U23304 (N_23304,N_20186,N_21278);
and U23305 (N_23305,N_20462,N_21617);
nor U23306 (N_23306,N_21165,N_21454);
nor U23307 (N_23307,N_20000,N_22149);
or U23308 (N_23308,N_20680,N_20441);
or U23309 (N_23309,N_20034,N_22096);
or U23310 (N_23310,N_22268,N_21189);
nor U23311 (N_23311,N_21414,N_22147);
xor U23312 (N_23312,N_20874,N_20264);
xnor U23313 (N_23313,N_22211,N_20519);
xnor U23314 (N_23314,N_22197,N_21525);
or U23315 (N_23315,N_21147,N_22055);
nand U23316 (N_23316,N_22479,N_21057);
or U23317 (N_23317,N_21146,N_20024);
or U23318 (N_23318,N_21924,N_21621);
nor U23319 (N_23319,N_21411,N_20424);
xor U23320 (N_23320,N_22119,N_21981);
nand U23321 (N_23321,N_21438,N_22460);
and U23322 (N_23322,N_21658,N_21804);
nand U23323 (N_23323,N_21044,N_21953);
or U23324 (N_23324,N_20658,N_20383);
xor U23325 (N_23325,N_20862,N_20654);
nand U23326 (N_23326,N_21985,N_22179);
nor U23327 (N_23327,N_20885,N_21951);
or U23328 (N_23328,N_20540,N_20738);
nand U23329 (N_23329,N_20092,N_21100);
nand U23330 (N_23330,N_22178,N_22207);
xnor U23331 (N_23331,N_21169,N_21915);
nor U23332 (N_23332,N_21877,N_20093);
xnor U23333 (N_23333,N_20437,N_21929);
xnor U23334 (N_23334,N_20834,N_20139);
and U23335 (N_23335,N_21797,N_21770);
or U23336 (N_23336,N_21111,N_20559);
or U23337 (N_23337,N_21698,N_20380);
nand U23338 (N_23338,N_20132,N_21455);
or U23339 (N_23339,N_20573,N_20354);
or U23340 (N_23340,N_21484,N_20981);
or U23341 (N_23341,N_22335,N_21996);
nand U23342 (N_23342,N_20905,N_22362);
nand U23343 (N_23343,N_20501,N_21366);
or U23344 (N_23344,N_20428,N_20195);
nor U23345 (N_23345,N_22296,N_21094);
and U23346 (N_23346,N_21905,N_22491);
nor U23347 (N_23347,N_20316,N_21887);
nor U23348 (N_23348,N_20963,N_22316);
nor U23349 (N_23349,N_21413,N_20006);
and U23350 (N_23350,N_22402,N_21884);
and U23351 (N_23351,N_22050,N_21871);
or U23352 (N_23352,N_20932,N_22162);
and U23353 (N_23353,N_22439,N_22158);
nor U23354 (N_23354,N_21600,N_20924);
nor U23355 (N_23355,N_20121,N_20698);
nand U23356 (N_23356,N_21272,N_21444);
nor U23357 (N_23357,N_22376,N_22139);
nand U23358 (N_23358,N_20447,N_22127);
or U23359 (N_23359,N_20347,N_20578);
nand U23360 (N_23360,N_20760,N_21157);
or U23361 (N_23361,N_21916,N_21799);
nand U23362 (N_23362,N_20449,N_22433);
nand U23363 (N_23363,N_22424,N_20043);
and U23364 (N_23364,N_22134,N_21560);
xor U23365 (N_23365,N_21611,N_21293);
or U23366 (N_23366,N_21275,N_22217);
nand U23367 (N_23367,N_22024,N_22464);
xnor U23368 (N_23368,N_20946,N_20415);
and U23369 (N_23369,N_22079,N_20392);
nor U23370 (N_23370,N_21615,N_20057);
and U23371 (N_23371,N_22463,N_20713);
nand U23372 (N_23372,N_21016,N_22201);
xor U23373 (N_23373,N_21324,N_22073);
nor U23374 (N_23374,N_22116,N_20631);
nand U23375 (N_23375,N_22192,N_21644);
nand U23376 (N_23376,N_21585,N_20846);
nand U23377 (N_23377,N_20147,N_22473);
nand U23378 (N_23378,N_21762,N_20261);
nor U23379 (N_23379,N_22383,N_21610);
xnor U23380 (N_23380,N_20492,N_21213);
xnor U23381 (N_23381,N_22046,N_20448);
and U23382 (N_23382,N_20555,N_22125);
and U23383 (N_23383,N_21625,N_20485);
xnor U23384 (N_23384,N_22111,N_22009);
nor U23385 (N_23385,N_20741,N_20201);
nand U23386 (N_23386,N_20832,N_21919);
or U23387 (N_23387,N_21768,N_20640);
nor U23388 (N_23388,N_20558,N_21106);
nand U23389 (N_23389,N_20337,N_22396);
nand U23390 (N_23390,N_20004,N_20697);
and U23391 (N_23391,N_22408,N_22161);
xnor U23392 (N_23392,N_20761,N_21399);
and U23393 (N_23393,N_20759,N_22025);
or U23394 (N_23394,N_20506,N_21470);
nor U23395 (N_23395,N_21702,N_22459);
xor U23396 (N_23396,N_22235,N_22230);
xor U23397 (N_23397,N_20938,N_20183);
xnor U23398 (N_23398,N_22066,N_20279);
nor U23399 (N_23399,N_20524,N_22057);
xnor U23400 (N_23400,N_21222,N_20551);
and U23401 (N_23401,N_20344,N_20710);
nand U23402 (N_23402,N_22187,N_21305);
and U23403 (N_23403,N_22321,N_21579);
nor U23404 (N_23404,N_20895,N_22242);
and U23405 (N_23405,N_20358,N_21654);
nor U23406 (N_23406,N_21926,N_21700);
nor U23407 (N_23407,N_20083,N_20518);
or U23408 (N_23408,N_20853,N_21738);
or U23409 (N_23409,N_21105,N_20409);
and U23410 (N_23410,N_21726,N_21928);
nor U23411 (N_23411,N_20979,N_21021);
nand U23412 (N_23412,N_22121,N_20928);
nand U23413 (N_23413,N_20700,N_21279);
nor U23414 (N_23414,N_22154,N_21068);
or U23415 (N_23415,N_21047,N_22286);
and U23416 (N_23416,N_21037,N_20443);
and U23417 (N_23417,N_22270,N_20838);
nand U23418 (N_23418,N_22363,N_20684);
nor U23419 (N_23419,N_20516,N_21767);
xor U23420 (N_23420,N_21337,N_21721);
nor U23421 (N_23421,N_22365,N_21344);
and U23422 (N_23422,N_22274,N_20888);
nand U23423 (N_23423,N_21680,N_21733);
xnor U23424 (N_23424,N_21760,N_22103);
nand U23425 (N_23425,N_20644,N_21689);
nand U23426 (N_23426,N_20950,N_21918);
or U23427 (N_23427,N_20805,N_20756);
nand U23428 (N_23428,N_21145,N_21168);
nand U23429 (N_23429,N_22494,N_21993);
or U23430 (N_23430,N_21089,N_20763);
nor U23431 (N_23431,N_22349,N_22023);
xor U23432 (N_23432,N_22304,N_22160);
and U23433 (N_23433,N_21225,N_20179);
nand U23434 (N_23434,N_21061,N_20616);
and U23435 (N_23435,N_21379,N_20128);
or U23436 (N_23436,N_22078,N_22488);
or U23437 (N_23437,N_21175,N_21526);
nand U23438 (N_23438,N_22330,N_20363);
or U23439 (N_23439,N_21197,N_20695);
nor U23440 (N_23440,N_21307,N_21836);
nand U23441 (N_23441,N_22151,N_20771);
nor U23442 (N_23442,N_20820,N_20982);
nand U23443 (N_23443,N_21039,N_21428);
or U23444 (N_23444,N_21408,N_21861);
or U23445 (N_23445,N_21286,N_20782);
nor U23446 (N_23446,N_22371,N_20127);
and U23447 (N_23447,N_21255,N_20873);
xnor U23448 (N_23448,N_20844,N_21398);
nor U23449 (N_23449,N_21014,N_21417);
nand U23450 (N_23450,N_20550,N_20662);
xor U23451 (N_23451,N_20228,N_22384);
and U23452 (N_23452,N_21838,N_20185);
nor U23453 (N_23453,N_20712,N_21281);
and U23454 (N_23454,N_20686,N_21390);
or U23455 (N_23455,N_21606,N_22480);
nor U23456 (N_23456,N_20118,N_22358);
xor U23457 (N_23457,N_21729,N_21935);
or U23458 (N_23458,N_20650,N_20817);
xor U23459 (N_23459,N_21419,N_21537);
and U23460 (N_23460,N_21297,N_22065);
or U23461 (N_23461,N_21947,N_20509);
xnor U23462 (N_23462,N_22272,N_20188);
and U23463 (N_23463,N_21950,N_20094);
xnor U23464 (N_23464,N_20593,N_20637);
nand U23465 (N_23465,N_21023,N_21193);
nand U23466 (N_23466,N_22049,N_21528);
nor U23467 (N_23467,N_21626,N_20175);
nor U23468 (N_23468,N_21400,N_22332);
and U23469 (N_23469,N_20144,N_22496);
nand U23470 (N_23470,N_20421,N_22124);
nand U23471 (N_23471,N_20167,N_21727);
and U23472 (N_23472,N_21085,N_20718);
nor U23473 (N_23473,N_20921,N_22102);
nand U23474 (N_23474,N_21972,N_20050);
nand U23475 (N_23475,N_21535,N_21907);
or U23476 (N_23476,N_21431,N_22077);
and U23477 (N_23477,N_21679,N_21988);
xor U23478 (N_23478,N_20542,N_22273);
nor U23479 (N_23479,N_22020,N_21412);
or U23480 (N_23480,N_22427,N_20726);
or U23481 (N_23481,N_21876,N_20073);
nand U23482 (N_23482,N_22190,N_21088);
nand U23483 (N_23483,N_20735,N_21415);
nor U23484 (N_23484,N_21172,N_20869);
nor U23485 (N_23485,N_22409,N_21749);
nor U23486 (N_23486,N_22226,N_21544);
nor U23487 (N_23487,N_20570,N_20931);
or U23488 (N_23488,N_21112,N_20649);
nor U23489 (N_23489,N_21932,N_21092);
nand U23490 (N_23490,N_20819,N_21570);
xor U23491 (N_23491,N_21435,N_22199);
and U23492 (N_23492,N_20196,N_21122);
nand U23493 (N_23493,N_20273,N_21430);
nor U23494 (N_23494,N_20319,N_22221);
nor U23495 (N_23495,N_22416,N_21840);
and U23496 (N_23496,N_21730,N_22385);
nand U23497 (N_23497,N_21599,N_20952);
nand U23498 (N_23498,N_21933,N_20295);
xnor U23499 (N_23499,N_21355,N_20807);
xor U23500 (N_23500,N_20458,N_21282);
and U23501 (N_23501,N_21304,N_20477);
nor U23502 (N_23502,N_20971,N_20418);
and U23503 (N_23503,N_20190,N_20020);
or U23504 (N_23504,N_21084,N_20457);
and U23505 (N_23505,N_20315,N_21383);
xor U23506 (N_23506,N_20148,N_22155);
xor U23507 (N_23507,N_20472,N_21340);
nor U23508 (N_23508,N_20839,N_22248);
nor U23509 (N_23509,N_22007,N_20628);
and U23510 (N_23510,N_21391,N_20901);
and U23511 (N_23511,N_20360,N_21973);
or U23512 (N_23512,N_20214,N_21093);
nand U23513 (N_23513,N_20236,N_22346);
and U23514 (N_23514,N_20854,N_21961);
or U23515 (N_23515,N_21069,N_20226);
and U23516 (N_23516,N_20865,N_21418);
or U23517 (N_23517,N_20305,N_21081);
nor U23518 (N_23518,N_21220,N_20436);
nor U23519 (N_23519,N_22039,N_20526);
xor U23520 (N_23520,N_20715,N_20030);
and U23521 (N_23521,N_20352,N_21227);
nor U23522 (N_23522,N_21657,N_21065);
or U23523 (N_23523,N_21827,N_21975);
or U23524 (N_23524,N_20960,N_21210);
xor U23525 (N_23525,N_20079,N_20956);
nor U23526 (N_23526,N_20823,N_21487);
nor U23527 (N_23527,N_21787,N_20739);
and U23528 (N_23528,N_21750,N_20814);
nor U23529 (N_23529,N_21855,N_22302);
and U23530 (N_23530,N_20245,N_22067);
and U23531 (N_23531,N_20416,N_21277);
nand U23532 (N_23532,N_20788,N_21813);
nand U23533 (N_23533,N_21513,N_21063);
xnor U23534 (N_23534,N_20003,N_21310);
nor U23535 (N_23535,N_21311,N_20568);
and U23536 (N_23536,N_22225,N_20403);
xnor U23537 (N_23537,N_21208,N_20758);
xor U23538 (N_23538,N_21773,N_22423);
nand U23539 (N_23539,N_22216,N_20724);
or U23540 (N_23540,N_20990,N_20579);
and U23541 (N_23541,N_20106,N_22198);
nor U23542 (N_23542,N_20192,N_20964);
and U23543 (N_23543,N_20911,N_21555);
or U23544 (N_23544,N_22284,N_20937);
nor U23545 (N_23545,N_20460,N_22448);
and U23546 (N_23546,N_20799,N_20927);
or U23547 (N_23547,N_21747,N_21467);
xor U23548 (N_23548,N_20340,N_20612);
nand U23549 (N_23549,N_20656,N_20341);
or U23550 (N_23550,N_21997,N_21338);
nand U23551 (N_23551,N_21616,N_21882);
or U23552 (N_23552,N_20171,N_20117);
and U23553 (N_23553,N_21856,N_20239);
or U23554 (N_23554,N_20140,N_21776);
or U23555 (N_23555,N_20682,N_22370);
xor U23556 (N_23556,N_21071,N_21826);
or U23557 (N_23557,N_20384,N_21930);
and U23558 (N_23558,N_22432,N_20789);
nor U23559 (N_23559,N_21288,N_20289);
nor U23560 (N_23560,N_22215,N_21567);
and U23561 (N_23561,N_20845,N_21315);
and U23562 (N_23562,N_21675,N_21661);
nor U23563 (N_23563,N_20307,N_20243);
or U23564 (N_23564,N_21204,N_21352);
nand U23565 (N_23565,N_22086,N_22183);
and U23566 (N_23566,N_21035,N_21504);
nor U23567 (N_23567,N_22256,N_22447);
nor U23568 (N_23568,N_20116,N_20397);
nor U23569 (N_23569,N_20933,N_22318);
nor U23570 (N_23570,N_22070,N_20062);
xor U23571 (N_23571,N_20080,N_20602);
xnor U23572 (N_23572,N_20836,N_22440);
xnor U23573 (N_23573,N_20281,N_21598);
and U23574 (N_23574,N_20493,N_22366);
or U23575 (N_23575,N_21971,N_20560);
and U23576 (N_23576,N_22426,N_21239);
and U23577 (N_23577,N_21133,N_21048);
nor U23578 (N_23578,N_21401,N_22417);
nand U23579 (N_23579,N_21835,N_21234);
or U23580 (N_23580,N_20867,N_20357);
nand U23581 (N_23581,N_21548,N_20851);
and U23582 (N_23582,N_21780,N_20023);
and U23583 (N_23583,N_21558,N_20227);
and U23584 (N_23584,N_21343,N_20599);
or U23585 (N_23585,N_20918,N_20687);
nand U23586 (N_23586,N_22194,N_22471);
nor U23587 (N_23587,N_22233,N_20786);
or U23588 (N_23588,N_22327,N_21483);
nand U23589 (N_23589,N_20207,N_21079);
xnor U23590 (N_23590,N_20527,N_20572);
or U23591 (N_23591,N_21815,N_21115);
nand U23592 (N_23592,N_20490,N_20957);
and U23593 (N_23593,N_20827,N_20112);
and U23594 (N_23594,N_22375,N_20897);
or U23595 (N_23595,N_22140,N_21458);
xor U23596 (N_23596,N_22018,N_21899);
xnor U23597 (N_23597,N_21562,N_20122);
and U23598 (N_23598,N_22209,N_20249);
nand U23599 (N_23599,N_22191,N_20991);
xor U23600 (N_23600,N_22481,N_22325);
nand U23601 (N_23601,N_21539,N_22010);
or U23602 (N_23602,N_20197,N_21938);
and U23603 (N_23603,N_20734,N_20996);
or U23604 (N_23604,N_22177,N_22129);
nor U23605 (N_23605,N_22081,N_20626);
or U23606 (N_23606,N_20916,N_21643);
nand U23607 (N_23607,N_20224,N_21378);
nor U23608 (N_23608,N_21722,N_20894);
and U23609 (N_23609,N_20161,N_20244);
nand U23610 (N_23610,N_20657,N_20115);
xor U23611 (N_23611,N_21468,N_21440);
or U23612 (N_23612,N_20775,N_22410);
and U23613 (N_23613,N_20059,N_20444);
xnor U23614 (N_23614,N_22064,N_20290);
or U23615 (N_23615,N_22083,N_20283);
nor U23616 (N_23616,N_20815,N_20317);
nor U23617 (N_23617,N_21274,N_22469);
or U23618 (N_23618,N_22300,N_21660);
nand U23619 (N_23619,N_20711,N_21922);
and U23620 (N_23620,N_22397,N_21987);
nor U23621 (N_23621,N_20235,N_21313);
xor U23622 (N_23622,N_21516,N_21519);
xor U23623 (N_23623,N_21795,N_21139);
and U23624 (N_23624,N_21142,N_21158);
nor U23625 (N_23625,N_22352,N_21949);
and U23626 (N_23626,N_20480,N_20066);
and U23627 (N_23627,N_21491,N_21205);
xor U23628 (N_23628,N_22047,N_20291);
xor U23629 (N_23629,N_22499,N_20052);
or U23630 (N_23630,N_21745,N_20538);
and U23631 (N_23631,N_20395,N_21831);
and U23632 (N_23632,N_21594,N_21387);
and U23633 (N_23633,N_20709,N_21500);
nand U23634 (N_23634,N_20368,N_22269);
nand U23635 (N_23635,N_22456,N_20508);
nand U23636 (N_23636,N_21393,N_21812);
or U23637 (N_23637,N_22133,N_20590);
and U23638 (N_23638,N_20387,N_22328);
xor U23639 (N_23639,N_21250,N_21503);
nand U23640 (N_23640,N_21424,N_22152);
nor U23641 (N_23641,N_21514,N_20801);
and U23642 (N_23642,N_21989,N_22110);
nor U23643 (N_23643,N_20353,N_22095);
xnor U23644 (N_23644,N_22379,N_20533);
or U23645 (N_23645,N_22259,N_20069);
nor U23646 (N_23646,N_20868,N_22080);
nor U23647 (N_23647,N_21690,N_21839);
or U23648 (N_23648,N_21939,N_21404);
and U23649 (N_23649,N_20507,N_20471);
nand U23650 (N_23650,N_21966,N_20575);
xor U23651 (N_23651,N_22059,N_21603);
or U23652 (N_23652,N_20329,N_20064);
nor U23653 (N_23653,N_20035,N_21034);
nor U23654 (N_23654,N_20676,N_20588);
nor U23655 (N_23655,N_20544,N_21847);
nand U23656 (N_23656,N_20238,N_21941);
nand U23657 (N_23657,N_21493,N_20346);
xnor U23658 (N_23658,N_20505,N_22053);
or U23659 (N_23659,N_20878,N_20007);
xor U23660 (N_23660,N_20262,N_20182);
nor U23661 (N_23661,N_21808,N_22320);
nor U23662 (N_23662,N_22170,N_21582);
xor U23663 (N_23663,N_21082,N_20915);
xor U23664 (N_23664,N_21712,N_20984);
xnor U23665 (N_23665,N_20793,N_21731);
or U23666 (N_23666,N_22455,N_20632);
or U23667 (N_23667,N_22089,N_20489);
xor U23668 (N_23668,N_21531,N_22002);
nor U23669 (N_23669,N_21377,N_20571);
or U23670 (N_23670,N_22454,N_20439);
xnor U23671 (N_23671,N_20790,N_21701);
xor U23672 (N_23672,N_21365,N_21574);
and U23673 (N_23673,N_21790,N_20107);
or U23674 (N_23674,N_22266,N_20504);
nand U23675 (N_23675,N_20455,N_20716);
xor U23676 (N_23676,N_21968,N_21405);
nand U23677 (N_23677,N_21248,N_21964);
and U23678 (N_23678,N_20405,N_22137);
nand U23679 (N_23679,N_21183,N_20400);
and U23680 (N_23680,N_20156,N_20520);
and U23681 (N_23681,N_20113,N_20974);
nor U23682 (N_23682,N_22000,N_20242);
or U23683 (N_23683,N_21426,N_20970);
nor U23684 (N_23684,N_21026,N_21348);
nand U23685 (N_23685,N_21040,N_21684);
nor U23686 (N_23686,N_21270,N_20994);
or U23687 (N_23687,N_20142,N_20163);
nand U23688 (N_23688,N_21237,N_20831);
or U23689 (N_23689,N_20809,N_21178);
xnor U23690 (N_23690,N_21363,N_20278);
and U23691 (N_23691,N_20159,N_22265);
xnor U23692 (N_23692,N_21545,N_21999);
or U23693 (N_23693,N_22450,N_21314);
xnor U23694 (N_23694,N_21601,N_20101);
nor U23695 (N_23695,N_20180,N_21273);
xnor U23696 (N_23696,N_21346,N_21507);
and U23697 (N_23697,N_22374,N_21022);
and U23698 (N_23698,N_21347,N_22122);
xnor U23699 (N_23699,N_20103,N_20778);
xor U23700 (N_23700,N_21633,N_20029);
or U23701 (N_23701,N_21844,N_21357);
xor U23702 (N_23702,N_20225,N_21345);
xor U23703 (N_23703,N_20899,N_20203);
nand U23704 (N_23704,N_20902,N_20407);
and U23705 (N_23705,N_20596,N_20205);
or U23706 (N_23706,N_22441,N_21375);
and U23707 (N_23707,N_20345,N_22290);
or U23708 (N_23708,N_21294,N_21948);
nor U23709 (N_23709,N_22076,N_20184);
or U23710 (N_23710,N_20770,N_22188);
xnor U23711 (N_23711,N_21781,N_20940);
or U23712 (N_23712,N_22244,N_20848);
or U23713 (N_23713,N_20432,N_21746);
nand U23714 (N_23714,N_21629,N_21573);
nor U23715 (N_23715,N_20335,N_21995);
and U23716 (N_23716,N_21858,N_22184);
and U23717 (N_23717,N_21423,N_20372);
and U23718 (N_23718,N_20391,N_20130);
or U23719 (N_23719,N_22292,N_20936);
or U23720 (N_23720,N_20047,N_20618);
nor U23721 (N_23721,N_20220,N_21869);
xor U23722 (N_23722,N_22153,N_21160);
nor U23723 (N_23723,N_22389,N_21655);
or U23724 (N_23724,N_20980,N_21416);
and U23725 (N_23725,N_20284,N_21908);
nor U23726 (N_23726,N_21632,N_21565);
xor U23727 (N_23727,N_21732,N_22461);
or U23728 (N_23728,N_20174,N_20753);
xor U23729 (N_23729,N_21097,N_20525);
and U23730 (N_23730,N_20331,N_21671);
xor U23731 (N_23731,N_21488,N_21940);
and U23732 (N_23732,N_21368,N_22141);
xnor U23733 (N_23733,N_21439,N_20548);
xor U23734 (N_23734,N_21564,N_21757);
xnor U23735 (N_23735,N_22390,N_20696);
nand U23736 (N_23736,N_21356,N_20014);
and U23737 (N_23737,N_22403,N_20002);
or U23738 (N_23738,N_20038,N_22422);
xor U23739 (N_23739,N_21490,N_20500);
or U23740 (N_23740,N_20306,N_20442);
xnor U23741 (N_23741,N_20722,N_20732);
nor U23742 (N_23742,N_20737,N_21322);
nand U23743 (N_23743,N_22311,N_21076);
nand U23744 (N_23744,N_21867,N_21261);
nor U23745 (N_23745,N_22105,N_22398);
xnor U23746 (N_23746,N_21090,N_22401);
or U23747 (N_23747,N_20949,N_22490);
xnor U23748 (N_23748,N_20309,N_20255);
nor U23749 (N_23749,N_20787,N_21875);
xnor U23750 (N_23750,N_21561,N_21443);
or U23751 (N_23751,N_20223,N_20747);
xnor U23752 (N_23752,N_21653,N_20855);
nand U23753 (N_23753,N_21755,N_21074);
nand U23754 (N_23754,N_21178,N_21466);
nand U23755 (N_23755,N_22109,N_20424);
xnor U23756 (N_23756,N_20300,N_21504);
or U23757 (N_23757,N_20388,N_20243);
nor U23758 (N_23758,N_20016,N_20234);
or U23759 (N_23759,N_22289,N_21351);
nor U23760 (N_23760,N_20024,N_20638);
nor U23761 (N_23761,N_20094,N_20200);
and U23762 (N_23762,N_21439,N_20892);
nand U23763 (N_23763,N_21186,N_20218);
and U23764 (N_23764,N_20178,N_21973);
nor U23765 (N_23765,N_21643,N_21421);
or U23766 (N_23766,N_20153,N_20816);
and U23767 (N_23767,N_22169,N_22148);
xor U23768 (N_23768,N_22279,N_20523);
nand U23769 (N_23769,N_20848,N_20668);
nand U23770 (N_23770,N_22151,N_21532);
nand U23771 (N_23771,N_21259,N_20352);
nor U23772 (N_23772,N_21569,N_20148);
xor U23773 (N_23773,N_21592,N_22300);
nor U23774 (N_23774,N_22269,N_21810);
nor U23775 (N_23775,N_21506,N_20802);
and U23776 (N_23776,N_21769,N_20533);
xnor U23777 (N_23777,N_21672,N_21293);
or U23778 (N_23778,N_22315,N_20262);
nor U23779 (N_23779,N_22141,N_20595);
xnor U23780 (N_23780,N_22134,N_21109);
xnor U23781 (N_23781,N_22354,N_20403);
and U23782 (N_23782,N_20952,N_20971);
nor U23783 (N_23783,N_22459,N_20766);
xor U23784 (N_23784,N_21154,N_20900);
or U23785 (N_23785,N_20460,N_21004);
nand U23786 (N_23786,N_21091,N_20339);
nand U23787 (N_23787,N_22398,N_21674);
nor U23788 (N_23788,N_22218,N_21992);
or U23789 (N_23789,N_20009,N_20523);
nand U23790 (N_23790,N_22175,N_20135);
xor U23791 (N_23791,N_21989,N_20321);
nand U23792 (N_23792,N_21412,N_20885);
or U23793 (N_23793,N_22339,N_20650);
or U23794 (N_23794,N_22160,N_21834);
xnor U23795 (N_23795,N_21563,N_21851);
nor U23796 (N_23796,N_21085,N_21422);
or U23797 (N_23797,N_20653,N_21602);
or U23798 (N_23798,N_20521,N_20580);
or U23799 (N_23799,N_21343,N_21106);
nor U23800 (N_23800,N_21095,N_20496);
xnor U23801 (N_23801,N_20168,N_20071);
xor U23802 (N_23802,N_21601,N_21772);
xor U23803 (N_23803,N_21676,N_20322);
or U23804 (N_23804,N_20175,N_21721);
and U23805 (N_23805,N_20354,N_20781);
and U23806 (N_23806,N_22233,N_21538);
nand U23807 (N_23807,N_22455,N_21711);
xor U23808 (N_23808,N_20799,N_20752);
nor U23809 (N_23809,N_21146,N_21601);
nor U23810 (N_23810,N_20612,N_20996);
xor U23811 (N_23811,N_20507,N_21185);
xnor U23812 (N_23812,N_22473,N_21127);
nand U23813 (N_23813,N_21868,N_20846);
nor U23814 (N_23814,N_21974,N_22319);
xor U23815 (N_23815,N_21866,N_20443);
nor U23816 (N_23816,N_21854,N_22380);
xnor U23817 (N_23817,N_20667,N_20689);
or U23818 (N_23818,N_22120,N_21913);
or U23819 (N_23819,N_22462,N_20608);
or U23820 (N_23820,N_21565,N_21590);
and U23821 (N_23821,N_21307,N_20798);
or U23822 (N_23822,N_21319,N_21529);
nor U23823 (N_23823,N_22320,N_20035);
nor U23824 (N_23824,N_20228,N_21314);
nand U23825 (N_23825,N_20650,N_21040);
xnor U23826 (N_23826,N_21669,N_21912);
nor U23827 (N_23827,N_20828,N_21390);
nor U23828 (N_23828,N_20555,N_22171);
or U23829 (N_23829,N_20038,N_20763);
nor U23830 (N_23830,N_21976,N_21623);
xor U23831 (N_23831,N_21797,N_21130);
and U23832 (N_23832,N_20085,N_22141);
xor U23833 (N_23833,N_20969,N_22163);
nand U23834 (N_23834,N_22348,N_20992);
nand U23835 (N_23835,N_21378,N_20796);
nor U23836 (N_23836,N_21211,N_20090);
nand U23837 (N_23837,N_21360,N_20537);
xor U23838 (N_23838,N_21510,N_22352);
or U23839 (N_23839,N_20902,N_22317);
nand U23840 (N_23840,N_21015,N_20571);
xnor U23841 (N_23841,N_21241,N_20540);
nand U23842 (N_23842,N_20933,N_20797);
xor U23843 (N_23843,N_20945,N_22210);
nand U23844 (N_23844,N_20637,N_20460);
nor U23845 (N_23845,N_20322,N_22243);
nand U23846 (N_23846,N_20591,N_20336);
xor U23847 (N_23847,N_20590,N_22249);
and U23848 (N_23848,N_22361,N_21255);
xnor U23849 (N_23849,N_20813,N_20230);
xnor U23850 (N_23850,N_21150,N_20902);
xnor U23851 (N_23851,N_22188,N_21039);
and U23852 (N_23852,N_21698,N_20773);
and U23853 (N_23853,N_21083,N_21896);
nand U23854 (N_23854,N_21665,N_21844);
or U23855 (N_23855,N_20069,N_21853);
nor U23856 (N_23856,N_22476,N_21038);
nor U23857 (N_23857,N_21908,N_20308);
nand U23858 (N_23858,N_20352,N_20841);
nand U23859 (N_23859,N_20499,N_21209);
and U23860 (N_23860,N_21270,N_22080);
or U23861 (N_23861,N_21890,N_22182);
and U23862 (N_23862,N_21520,N_21795);
xor U23863 (N_23863,N_22475,N_21515);
and U23864 (N_23864,N_21481,N_20728);
or U23865 (N_23865,N_21734,N_22230);
nand U23866 (N_23866,N_21376,N_21102);
nand U23867 (N_23867,N_21814,N_21297);
and U23868 (N_23868,N_22416,N_20947);
xnor U23869 (N_23869,N_20511,N_21580);
xor U23870 (N_23870,N_21312,N_21372);
or U23871 (N_23871,N_21615,N_21215);
nand U23872 (N_23872,N_22008,N_22346);
and U23873 (N_23873,N_20655,N_22492);
and U23874 (N_23874,N_21532,N_20434);
nand U23875 (N_23875,N_22337,N_20096);
nor U23876 (N_23876,N_21089,N_21972);
nor U23877 (N_23877,N_22164,N_20922);
nand U23878 (N_23878,N_21911,N_20513);
or U23879 (N_23879,N_20248,N_21535);
xnor U23880 (N_23880,N_21300,N_21478);
or U23881 (N_23881,N_20570,N_20925);
xnor U23882 (N_23882,N_21713,N_22235);
or U23883 (N_23883,N_22390,N_22159);
xnor U23884 (N_23884,N_22179,N_20964);
xnor U23885 (N_23885,N_20433,N_21802);
and U23886 (N_23886,N_20082,N_22051);
xnor U23887 (N_23887,N_20020,N_20432);
and U23888 (N_23888,N_21213,N_20126);
or U23889 (N_23889,N_20380,N_20541);
and U23890 (N_23890,N_20827,N_22143);
xnor U23891 (N_23891,N_20410,N_20917);
or U23892 (N_23892,N_21330,N_21637);
and U23893 (N_23893,N_20397,N_21709);
nand U23894 (N_23894,N_21129,N_21528);
and U23895 (N_23895,N_21256,N_22174);
and U23896 (N_23896,N_21030,N_21020);
xnor U23897 (N_23897,N_21720,N_21358);
nand U23898 (N_23898,N_21152,N_20614);
nand U23899 (N_23899,N_21740,N_20612);
nor U23900 (N_23900,N_20805,N_22052);
nor U23901 (N_23901,N_20689,N_20883);
or U23902 (N_23902,N_22381,N_21638);
nand U23903 (N_23903,N_20454,N_21358);
and U23904 (N_23904,N_21353,N_21452);
and U23905 (N_23905,N_20937,N_20681);
and U23906 (N_23906,N_21654,N_20517);
xnor U23907 (N_23907,N_20127,N_20921);
or U23908 (N_23908,N_20525,N_21393);
nand U23909 (N_23909,N_21879,N_20084);
and U23910 (N_23910,N_20617,N_21844);
nor U23911 (N_23911,N_20973,N_21803);
xor U23912 (N_23912,N_20933,N_20136);
nor U23913 (N_23913,N_20765,N_22163);
nand U23914 (N_23914,N_20154,N_20492);
nor U23915 (N_23915,N_20226,N_21647);
or U23916 (N_23916,N_22170,N_20867);
nand U23917 (N_23917,N_20636,N_21647);
nand U23918 (N_23918,N_22339,N_20152);
xnor U23919 (N_23919,N_20298,N_20481);
and U23920 (N_23920,N_21365,N_22347);
xor U23921 (N_23921,N_21683,N_21256);
xnor U23922 (N_23922,N_20655,N_22128);
or U23923 (N_23923,N_20261,N_21029);
nand U23924 (N_23924,N_22169,N_20571);
xnor U23925 (N_23925,N_22260,N_22294);
or U23926 (N_23926,N_21714,N_21716);
nand U23927 (N_23927,N_20034,N_20226);
or U23928 (N_23928,N_22095,N_20500);
nor U23929 (N_23929,N_21694,N_21788);
nor U23930 (N_23930,N_22110,N_21329);
or U23931 (N_23931,N_21331,N_20055);
nand U23932 (N_23932,N_21142,N_20600);
nor U23933 (N_23933,N_21371,N_22080);
xor U23934 (N_23934,N_20700,N_20583);
xor U23935 (N_23935,N_21999,N_20241);
and U23936 (N_23936,N_21625,N_21621);
nor U23937 (N_23937,N_21188,N_20135);
or U23938 (N_23938,N_22061,N_21604);
nor U23939 (N_23939,N_21592,N_21121);
and U23940 (N_23940,N_20099,N_21292);
nand U23941 (N_23941,N_20166,N_20649);
nor U23942 (N_23942,N_22158,N_20916);
nand U23943 (N_23943,N_22011,N_20623);
nand U23944 (N_23944,N_20411,N_22414);
xnor U23945 (N_23945,N_21906,N_20133);
nand U23946 (N_23946,N_20680,N_21938);
nand U23947 (N_23947,N_21277,N_20021);
nor U23948 (N_23948,N_22059,N_20921);
nand U23949 (N_23949,N_20760,N_22143);
or U23950 (N_23950,N_20640,N_20194);
xor U23951 (N_23951,N_20993,N_22040);
or U23952 (N_23952,N_22195,N_20823);
nor U23953 (N_23953,N_21532,N_20135);
xor U23954 (N_23954,N_21977,N_20727);
and U23955 (N_23955,N_21126,N_20215);
or U23956 (N_23956,N_21641,N_20421);
or U23957 (N_23957,N_21676,N_21094);
and U23958 (N_23958,N_20871,N_21354);
and U23959 (N_23959,N_21922,N_21005);
nor U23960 (N_23960,N_20359,N_22479);
or U23961 (N_23961,N_20083,N_20763);
xnor U23962 (N_23962,N_21448,N_21297);
nor U23963 (N_23963,N_21496,N_22371);
xnor U23964 (N_23964,N_20915,N_22048);
nor U23965 (N_23965,N_22198,N_20962);
nand U23966 (N_23966,N_22323,N_21595);
or U23967 (N_23967,N_20027,N_22456);
or U23968 (N_23968,N_21796,N_20534);
nand U23969 (N_23969,N_20537,N_20614);
or U23970 (N_23970,N_21724,N_21026);
nor U23971 (N_23971,N_21538,N_21370);
xnor U23972 (N_23972,N_20326,N_22250);
nand U23973 (N_23973,N_21589,N_21050);
nor U23974 (N_23974,N_21330,N_21970);
nor U23975 (N_23975,N_22398,N_22354);
and U23976 (N_23976,N_20849,N_20551);
or U23977 (N_23977,N_20470,N_21781);
and U23978 (N_23978,N_21809,N_21561);
or U23979 (N_23979,N_22498,N_20336);
nor U23980 (N_23980,N_21115,N_22422);
nand U23981 (N_23981,N_22401,N_21376);
xor U23982 (N_23982,N_21735,N_20937);
nand U23983 (N_23983,N_20036,N_20392);
or U23984 (N_23984,N_20086,N_21478);
xnor U23985 (N_23985,N_22338,N_20715);
nand U23986 (N_23986,N_21772,N_21807);
nor U23987 (N_23987,N_20301,N_20577);
xor U23988 (N_23988,N_20096,N_21787);
nand U23989 (N_23989,N_21457,N_21743);
nor U23990 (N_23990,N_22168,N_21986);
and U23991 (N_23991,N_22309,N_21995);
nand U23992 (N_23992,N_21578,N_21679);
nor U23993 (N_23993,N_21637,N_20302);
and U23994 (N_23994,N_21771,N_20466);
xor U23995 (N_23995,N_21033,N_20440);
and U23996 (N_23996,N_21316,N_20852);
nand U23997 (N_23997,N_21853,N_20085);
or U23998 (N_23998,N_20478,N_21151);
and U23999 (N_23999,N_22434,N_21154);
nor U24000 (N_24000,N_20599,N_20047);
or U24001 (N_24001,N_20621,N_22107);
or U24002 (N_24002,N_20722,N_21800);
xnor U24003 (N_24003,N_21669,N_21767);
nor U24004 (N_24004,N_21405,N_22295);
xnor U24005 (N_24005,N_20032,N_21329);
and U24006 (N_24006,N_21718,N_20490);
nand U24007 (N_24007,N_20805,N_21983);
nand U24008 (N_24008,N_20740,N_21385);
or U24009 (N_24009,N_21128,N_21084);
xor U24010 (N_24010,N_21737,N_22369);
xnor U24011 (N_24011,N_22279,N_21420);
and U24012 (N_24012,N_20976,N_20450);
nand U24013 (N_24013,N_20874,N_20455);
xnor U24014 (N_24014,N_21049,N_20756);
nand U24015 (N_24015,N_21621,N_20915);
and U24016 (N_24016,N_20976,N_21732);
or U24017 (N_24017,N_20360,N_21774);
or U24018 (N_24018,N_21829,N_22191);
or U24019 (N_24019,N_20504,N_21699);
xnor U24020 (N_24020,N_21983,N_20798);
or U24021 (N_24021,N_21181,N_21389);
and U24022 (N_24022,N_21855,N_21460);
nand U24023 (N_24023,N_20978,N_20641);
nor U24024 (N_24024,N_22306,N_21652);
or U24025 (N_24025,N_20629,N_20614);
nand U24026 (N_24026,N_22036,N_20228);
xor U24027 (N_24027,N_21217,N_22368);
xnor U24028 (N_24028,N_22496,N_22186);
xnor U24029 (N_24029,N_21892,N_21758);
and U24030 (N_24030,N_22424,N_21334);
and U24031 (N_24031,N_22387,N_20779);
nand U24032 (N_24032,N_20424,N_22135);
xor U24033 (N_24033,N_21737,N_20444);
nor U24034 (N_24034,N_20765,N_21828);
or U24035 (N_24035,N_20987,N_21838);
xor U24036 (N_24036,N_21655,N_20211);
nor U24037 (N_24037,N_20338,N_21775);
nor U24038 (N_24038,N_20608,N_20887);
nor U24039 (N_24039,N_22346,N_20499);
nor U24040 (N_24040,N_21052,N_20519);
nor U24041 (N_24041,N_20997,N_22354);
xor U24042 (N_24042,N_22279,N_22152);
nand U24043 (N_24043,N_21349,N_20676);
and U24044 (N_24044,N_21908,N_22011);
xnor U24045 (N_24045,N_22247,N_22255);
and U24046 (N_24046,N_22369,N_20994);
and U24047 (N_24047,N_21691,N_21131);
xnor U24048 (N_24048,N_22169,N_21915);
nor U24049 (N_24049,N_20124,N_22230);
or U24050 (N_24050,N_20185,N_20092);
nor U24051 (N_24051,N_20172,N_20407);
xor U24052 (N_24052,N_22215,N_21595);
nor U24053 (N_24053,N_20201,N_21262);
nand U24054 (N_24054,N_21104,N_21704);
and U24055 (N_24055,N_22489,N_20715);
and U24056 (N_24056,N_21868,N_21675);
xnor U24057 (N_24057,N_21425,N_20299);
nor U24058 (N_24058,N_21542,N_20372);
or U24059 (N_24059,N_21595,N_22260);
xnor U24060 (N_24060,N_20116,N_20784);
or U24061 (N_24061,N_22482,N_22214);
or U24062 (N_24062,N_20703,N_22402);
and U24063 (N_24063,N_22027,N_21094);
nand U24064 (N_24064,N_20369,N_22111);
and U24065 (N_24065,N_21112,N_21838);
nand U24066 (N_24066,N_21778,N_21373);
xor U24067 (N_24067,N_22435,N_20608);
and U24068 (N_24068,N_21896,N_20463);
xnor U24069 (N_24069,N_21074,N_21583);
nor U24070 (N_24070,N_20900,N_21233);
nor U24071 (N_24071,N_21935,N_22139);
nor U24072 (N_24072,N_20195,N_21802);
nand U24073 (N_24073,N_20588,N_21811);
nor U24074 (N_24074,N_21447,N_20815);
nand U24075 (N_24075,N_21712,N_21440);
nand U24076 (N_24076,N_21274,N_22175);
nor U24077 (N_24077,N_20777,N_20440);
nor U24078 (N_24078,N_20454,N_20445);
nand U24079 (N_24079,N_22094,N_22025);
nor U24080 (N_24080,N_21108,N_21883);
and U24081 (N_24081,N_21914,N_21936);
xor U24082 (N_24082,N_21294,N_21148);
xor U24083 (N_24083,N_22030,N_21614);
nand U24084 (N_24084,N_21633,N_20289);
nand U24085 (N_24085,N_21119,N_22435);
xnor U24086 (N_24086,N_22485,N_22301);
nor U24087 (N_24087,N_22420,N_20564);
xor U24088 (N_24088,N_22322,N_21625);
nand U24089 (N_24089,N_20032,N_21810);
and U24090 (N_24090,N_21179,N_20240);
or U24091 (N_24091,N_20288,N_21709);
or U24092 (N_24092,N_21901,N_22236);
or U24093 (N_24093,N_22316,N_21483);
or U24094 (N_24094,N_20225,N_21206);
or U24095 (N_24095,N_22348,N_20173);
nand U24096 (N_24096,N_21829,N_20337);
nor U24097 (N_24097,N_21740,N_20459);
xor U24098 (N_24098,N_22025,N_21633);
or U24099 (N_24099,N_21344,N_22241);
xor U24100 (N_24100,N_22440,N_20687);
or U24101 (N_24101,N_20033,N_21404);
nand U24102 (N_24102,N_20360,N_21685);
nor U24103 (N_24103,N_21799,N_20485);
nor U24104 (N_24104,N_20386,N_21467);
and U24105 (N_24105,N_21283,N_20236);
nand U24106 (N_24106,N_20039,N_20187);
and U24107 (N_24107,N_22354,N_22379);
nand U24108 (N_24108,N_21841,N_20742);
nor U24109 (N_24109,N_22270,N_22494);
nor U24110 (N_24110,N_21490,N_21609);
nor U24111 (N_24111,N_21473,N_21672);
and U24112 (N_24112,N_22008,N_21052);
xor U24113 (N_24113,N_22039,N_21581);
nand U24114 (N_24114,N_20343,N_21915);
nor U24115 (N_24115,N_21386,N_20273);
nor U24116 (N_24116,N_20471,N_21292);
or U24117 (N_24117,N_21004,N_20878);
xnor U24118 (N_24118,N_20468,N_21134);
nor U24119 (N_24119,N_21230,N_22233);
or U24120 (N_24120,N_20601,N_21316);
xor U24121 (N_24121,N_20134,N_20852);
xor U24122 (N_24122,N_20441,N_21334);
nor U24123 (N_24123,N_20030,N_21932);
nand U24124 (N_24124,N_21883,N_20356);
and U24125 (N_24125,N_20194,N_20339);
xnor U24126 (N_24126,N_20639,N_21683);
nand U24127 (N_24127,N_21242,N_20228);
xnor U24128 (N_24128,N_20026,N_21915);
and U24129 (N_24129,N_21091,N_21292);
nor U24130 (N_24130,N_21320,N_20934);
nand U24131 (N_24131,N_22276,N_21133);
nand U24132 (N_24132,N_21209,N_21688);
xnor U24133 (N_24133,N_21794,N_22225);
or U24134 (N_24134,N_21137,N_21668);
nand U24135 (N_24135,N_21561,N_20828);
nor U24136 (N_24136,N_21591,N_22102);
and U24137 (N_24137,N_20563,N_22417);
xnor U24138 (N_24138,N_22182,N_20666);
nand U24139 (N_24139,N_20523,N_20251);
or U24140 (N_24140,N_20959,N_22372);
or U24141 (N_24141,N_21304,N_22433);
nand U24142 (N_24142,N_20771,N_22458);
nor U24143 (N_24143,N_22321,N_21092);
or U24144 (N_24144,N_22223,N_21581);
or U24145 (N_24145,N_21843,N_22433);
or U24146 (N_24146,N_22222,N_20593);
or U24147 (N_24147,N_20040,N_22276);
nand U24148 (N_24148,N_21407,N_20408);
nand U24149 (N_24149,N_20209,N_20746);
nand U24150 (N_24150,N_22273,N_21240);
or U24151 (N_24151,N_22033,N_20984);
xnor U24152 (N_24152,N_22167,N_20112);
and U24153 (N_24153,N_21575,N_21784);
xor U24154 (N_24154,N_21388,N_21024);
nand U24155 (N_24155,N_21543,N_20559);
nor U24156 (N_24156,N_22417,N_21376);
and U24157 (N_24157,N_21814,N_21553);
nor U24158 (N_24158,N_20056,N_20235);
or U24159 (N_24159,N_20292,N_20688);
or U24160 (N_24160,N_21312,N_22418);
xor U24161 (N_24161,N_21244,N_20165);
xnor U24162 (N_24162,N_20373,N_22168);
or U24163 (N_24163,N_22391,N_20522);
nand U24164 (N_24164,N_21834,N_21756);
xor U24165 (N_24165,N_20199,N_21902);
or U24166 (N_24166,N_21474,N_20237);
and U24167 (N_24167,N_20173,N_21387);
nor U24168 (N_24168,N_20689,N_21965);
or U24169 (N_24169,N_21958,N_21915);
nor U24170 (N_24170,N_20508,N_20421);
or U24171 (N_24171,N_20245,N_20937);
nor U24172 (N_24172,N_21502,N_21297);
xor U24173 (N_24173,N_21365,N_21457);
and U24174 (N_24174,N_20949,N_22354);
nand U24175 (N_24175,N_22246,N_21328);
xor U24176 (N_24176,N_21088,N_22172);
nor U24177 (N_24177,N_21395,N_22402);
or U24178 (N_24178,N_22087,N_21265);
and U24179 (N_24179,N_21773,N_20851);
or U24180 (N_24180,N_20361,N_20888);
nand U24181 (N_24181,N_21069,N_22497);
nor U24182 (N_24182,N_20109,N_21526);
xor U24183 (N_24183,N_22225,N_20379);
nand U24184 (N_24184,N_21867,N_21524);
and U24185 (N_24185,N_21360,N_21850);
nand U24186 (N_24186,N_20797,N_21555);
nor U24187 (N_24187,N_21973,N_20897);
or U24188 (N_24188,N_21046,N_20481);
and U24189 (N_24189,N_21929,N_20421);
xnor U24190 (N_24190,N_22479,N_20765);
or U24191 (N_24191,N_22166,N_20387);
xnor U24192 (N_24192,N_22483,N_21896);
xor U24193 (N_24193,N_21464,N_21693);
or U24194 (N_24194,N_22179,N_20399);
xor U24195 (N_24195,N_21131,N_21040);
or U24196 (N_24196,N_20384,N_21720);
xor U24197 (N_24197,N_20775,N_20154);
nand U24198 (N_24198,N_21119,N_22178);
and U24199 (N_24199,N_22144,N_21107);
or U24200 (N_24200,N_22207,N_21215);
nand U24201 (N_24201,N_20985,N_21401);
xor U24202 (N_24202,N_22187,N_21872);
nor U24203 (N_24203,N_22160,N_20759);
nand U24204 (N_24204,N_20391,N_20641);
nand U24205 (N_24205,N_21529,N_20477);
and U24206 (N_24206,N_21297,N_21474);
nand U24207 (N_24207,N_20982,N_22300);
nand U24208 (N_24208,N_21070,N_20966);
and U24209 (N_24209,N_20633,N_21372);
nor U24210 (N_24210,N_21156,N_21718);
nor U24211 (N_24211,N_21140,N_22414);
and U24212 (N_24212,N_22325,N_21207);
or U24213 (N_24213,N_21391,N_21390);
or U24214 (N_24214,N_21386,N_22086);
nand U24215 (N_24215,N_20769,N_20753);
and U24216 (N_24216,N_21920,N_21878);
nand U24217 (N_24217,N_20303,N_20547);
or U24218 (N_24218,N_21000,N_21388);
xor U24219 (N_24219,N_22179,N_22334);
or U24220 (N_24220,N_21849,N_21138);
xor U24221 (N_24221,N_21245,N_20128);
and U24222 (N_24222,N_21667,N_21967);
nor U24223 (N_24223,N_21354,N_20824);
nand U24224 (N_24224,N_22106,N_21770);
and U24225 (N_24225,N_20422,N_20048);
nand U24226 (N_24226,N_20444,N_22462);
or U24227 (N_24227,N_21246,N_20003);
nor U24228 (N_24228,N_21198,N_21112);
nor U24229 (N_24229,N_21385,N_20664);
nand U24230 (N_24230,N_21501,N_20086);
nor U24231 (N_24231,N_20969,N_20391);
xor U24232 (N_24232,N_21328,N_20844);
or U24233 (N_24233,N_20052,N_20280);
or U24234 (N_24234,N_21454,N_22395);
and U24235 (N_24235,N_20825,N_22402);
and U24236 (N_24236,N_20785,N_20357);
and U24237 (N_24237,N_20334,N_20694);
nor U24238 (N_24238,N_21174,N_21853);
and U24239 (N_24239,N_22236,N_21767);
xor U24240 (N_24240,N_21029,N_21844);
nor U24241 (N_24241,N_20444,N_21603);
or U24242 (N_24242,N_21250,N_21622);
and U24243 (N_24243,N_21603,N_20720);
xnor U24244 (N_24244,N_20111,N_20874);
nor U24245 (N_24245,N_20003,N_20495);
and U24246 (N_24246,N_20627,N_20966);
and U24247 (N_24247,N_20909,N_22089);
nor U24248 (N_24248,N_21620,N_21090);
nor U24249 (N_24249,N_21661,N_20042);
nor U24250 (N_24250,N_20341,N_20248);
or U24251 (N_24251,N_22239,N_22444);
and U24252 (N_24252,N_21493,N_20727);
or U24253 (N_24253,N_22135,N_20189);
or U24254 (N_24254,N_21347,N_21902);
nand U24255 (N_24255,N_22298,N_20266);
nand U24256 (N_24256,N_21999,N_21680);
nor U24257 (N_24257,N_20510,N_20556);
and U24258 (N_24258,N_21920,N_21717);
xor U24259 (N_24259,N_20575,N_21997);
nand U24260 (N_24260,N_21890,N_22331);
or U24261 (N_24261,N_22048,N_21823);
nand U24262 (N_24262,N_22080,N_20187);
and U24263 (N_24263,N_21408,N_22241);
nor U24264 (N_24264,N_22412,N_22276);
nand U24265 (N_24265,N_21668,N_22270);
nand U24266 (N_24266,N_20120,N_20379);
and U24267 (N_24267,N_21634,N_20866);
or U24268 (N_24268,N_21751,N_20734);
and U24269 (N_24269,N_20500,N_22454);
and U24270 (N_24270,N_20297,N_20169);
or U24271 (N_24271,N_21167,N_20906);
and U24272 (N_24272,N_21044,N_21792);
and U24273 (N_24273,N_21088,N_22365);
xnor U24274 (N_24274,N_22400,N_21187);
xnor U24275 (N_24275,N_22312,N_20708);
nand U24276 (N_24276,N_20621,N_21308);
nor U24277 (N_24277,N_21812,N_20867);
or U24278 (N_24278,N_22179,N_20109);
xor U24279 (N_24279,N_22368,N_20379);
nor U24280 (N_24280,N_20263,N_21909);
and U24281 (N_24281,N_20600,N_21890);
xnor U24282 (N_24282,N_21503,N_22152);
nand U24283 (N_24283,N_22003,N_20615);
nand U24284 (N_24284,N_20649,N_21719);
nand U24285 (N_24285,N_21024,N_21597);
nand U24286 (N_24286,N_20662,N_22297);
nand U24287 (N_24287,N_22092,N_20250);
or U24288 (N_24288,N_21061,N_21147);
and U24289 (N_24289,N_21861,N_22042);
nor U24290 (N_24290,N_21973,N_21326);
nand U24291 (N_24291,N_20617,N_20363);
or U24292 (N_24292,N_21585,N_21651);
nor U24293 (N_24293,N_22136,N_20431);
xor U24294 (N_24294,N_20538,N_20906);
nor U24295 (N_24295,N_20341,N_20692);
xor U24296 (N_24296,N_20032,N_20795);
or U24297 (N_24297,N_20296,N_20273);
or U24298 (N_24298,N_21283,N_21089);
nor U24299 (N_24299,N_21765,N_21856);
and U24300 (N_24300,N_21852,N_20264);
nor U24301 (N_24301,N_21842,N_22080);
xor U24302 (N_24302,N_21902,N_21571);
and U24303 (N_24303,N_21735,N_22113);
nor U24304 (N_24304,N_20635,N_21405);
and U24305 (N_24305,N_20737,N_21570);
nand U24306 (N_24306,N_21305,N_21540);
nor U24307 (N_24307,N_21411,N_21878);
or U24308 (N_24308,N_21301,N_21970);
xnor U24309 (N_24309,N_22113,N_20435);
or U24310 (N_24310,N_20539,N_21508);
xnor U24311 (N_24311,N_20642,N_21311);
nor U24312 (N_24312,N_21895,N_20783);
xnor U24313 (N_24313,N_21768,N_22042);
nor U24314 (N_24314,N_22109,N_22207);
or U24315 (N_24315,N_21048,N_22122);
nor U24316 (N_24316,N_20148,N_21783);
xor U24317 (N_24317,N_20389,N_21964);
and U24318 (N_24318,N_22201,N_20086);
xor U24319 (N_24319,N_20357,N_20783);
or U24320 (N_24320,N_20944,N_20574);
xnor U24321 (N_24321,N_20265,N_20361);
or U24322 (N_24322,N_21838,N_21534);
xnor U24323 (N_24323,N_20201,N_21098);
nor U24324 (N_24324,N_21270,N_21808);
or U24325 (N_24325,N_20553,N_22218);
nand U24326 (N_24326,N_21641,N_20209);
xor U24327 (N_24327,N_20338,N_20649);
or U24328 (N_24328,N_20220,N_20232);
or U24329 (N_24329,N_21896,N_22146);
nor U24330 (N_24330,N_20713,N_21228);
or U24331 (N_24331,N_20058,N_20445);
nor U24332 (N_24332,N_21378,N_20913);
and U24333 (N_24333,N_21361,N_22311);
nand U24334 (N_24334,N_22308,N_20293);
and U24335 (N_24335,N_22378,N_20220);
nand U24336 (N_24336,N_22040,N_21381);
nand U24337 (N_24337,N_20653,N_21495);
and U24338 (N_24338,N_21897,N_20971);
and U24339 (N_24339,N_21939,N_21854);
or U24340 (N_24340,N_21789,N_20992);
or U24341 (N_24341,N_20316,N_21868);
nand U24342 (N_24342,N_20270,N_20803);
or U24343 (N_24343,N_20566,N_21835);
and U24344 (N_24344,N_20640,N_20146);
and U24345 (N_24345,N_20837,N_21181);
or U24346 (N_24346,N_21689,N_22380);
nor U24347 (N_24347,N_20002,N_21998);
nor U24348 (N_24348,N_20067,N_20718);
xor U24349 (N_24349,N_20042,N_22283);
nand U24350 (N_24350,N_22259,N_22451);
nor U24351 (N_24351,N_22163,N_22232);
and U24352 (N_24352,N_20487,N_20124);
nor U24353 (N_24353,N_20484,N_20003);
nor U24354 (N_24354,N_20432,N_20069);
and U24355 (N_24355,N_22297,N_20545);
and U24356 (N_24356,N_21710,N_22014);
nand U24357 (N_24357,N_20816,N_21747);
and U24358 (N_24358,N_20217,N_22136);
or U24359 (N_24359,N_20347,N_20509);
or U24360 (N_24360,N_21313,N_22467);
or U24361 (N_24361,N_21722,N_21121);
or U24362 (N_24362,N_20133,N_21116);
and U24363 (N_24363,N_20355,N_21780);
nand U24364 (N_24364,N_22145,N_21049);
or U24365 (N_24365,N_22485,N_22446);
and U24366 (N_24366,N_21987,N_21570);
xnor U24367 (N_24367,N_22396,N_20442);
or U24368 (N_24368,N_22013,N_22377);
nor U24369 (N_24369,N_22254,N_22083);
nand U24370 (N_24370,N_21082,N_20025);
nand U24371 (N_24371,N_21810,N_21864);
xor U24372 (N_24372,N_21563,N_20132);
nand U24373 (N_24373,N_22275,N_22495);
and U24374 (N_24374,N_20831,N_20701);
xnor U24375 (N_24375,N_21159,N_20659);
nor U24376 (N_24376,N_21041,N_20446);
and U24377 (N_24377,N_20827,N_20549);
or U24378 (N_24378,N_21594,N_21940);
xnor U24379 (N_24379,N_21494,N_21211);
or U24380 (N_24380,N_21798,N_21826);
xor U24381 (N_24381,N_20077,N_20381);
xnor U24382 (N_24382,N_20398,N_20548);
xor U24383 (N_24383,N_20200,N_21105);
or U24384 (N_24384,N_20699,N_20927);
nor U24385 (N_24385,N_21459,N_21650);
xnor U24386 (N_24386,N_21498,N_22101);
nor U24387 (N_24387,N_20530,N_20477);
and U24388 (N_24388,N_20823,N_22057);
nand U24389 (N_24389,N_21035,N_22036);
and U24390 (N_24390,N_21170,N_20115);
nand U24391 (N_24391,N_22066,N_21970);
xor U24392 (N_24392,N_20980,N_20932);
nor U24393 (N_24393,N_21216,N_21814);
and U24394 (N_24394,N_20992,N_20418);
nand U24395 (N_24395,N_21880,N_21295);
nor U24396 (N_24396,N_20603,N_22124);
xnor U24397 (N_24397,N_21216,N_20782);
xnor U24398 (N_24398,N_20092,N_20233);
nor U24399 (N_24399,N_20522,N_20338);
xnor U24400 (N_24400,N_21671,N_21299);
xnor U24401 (N_24401,N_20458,N_20212);
nand U24402 (N_24402,N_21125,N_20887);
and U24403 (N_24403,N_22434,N_21743);
or U24404 (N_24404,N_21134,N_21153);
nor U24405 (N_24405,N_22006,N_20642);
nand U24406 (N_24406,N_20640,N_21047);
xnor U24407 (N_24407,N_22380,N_22394);
nor U24408 (N_24408,N_22226,N_21943);
and U24409 (N_24409,N_20020,N_22024);
or U24410 (N_24410,N_20642,N_22149);
nor U24411 (N_24411,N_21233,N_20507);
or U24412 (N_24412,N_22048,N_22438);
nor U24413 (N_24413,N_21582,N_21399);
xor U24414 (N_24414,N_21485,N_22204);
nand U24415 (N_24415,N_22164,N_22315);
nor U24416 (N_24416,N_21876,N_20102);
and U24417 (N_24417,N_21568,N_20843);
xnor U24418 (N_24418,N_20743,N_22184);
nand U24419 (N_24419,N_22410,N_21394);
nor U24420 (N_24420,N_20547,N_21411);
xor U24421 (N_24421,N_20634,N_20741);
nand U24422 (N_24422,N_20531,N_21171);
and U24423 (N_24423,N_21772,N_21884);
nand U24424 (N_24424,N_22049,N_22075);
xnor U24425 (N_24425,N_20876,N_22288);
xnor U24426 (N_24426,N_21056,N_21755);
nor U24427 (N_24427,N_20679,N_21160);
xnor U24428 (N_24428,N_20842,N_21889);
nor U24429 (N_24429,N_20082,N_22337);
xnor U24430 (N_24430,N_21530,N_21156);
or U24431 (N_24431,N_20689,N_20260);
xor U24432 (N_24432,N_21001,N_21786);
xor U24433 (N_24433,N_20339,N_22099);
xnor U24434 (N_24434,N_20225,N_22200);
or U24435 (N_24435,N_20304,N_21585);
nor U24436 (N_24436,N_20468,N_20008);
xor U24437 (N_24437,N_21531,N_20575);
and U24438 (N_24438,N_22436,N_21231);
xnor U24439 (N_24439,N_20045,N_21714);
xnor U24440 (N_24440,N_20897,N_21015);
and U24441 (N_24441,N_21101,N_20520);
and U24442 (N_24442,N_21753,N_21124);
and U24443 (N_24443,N_20149,N_21629);
or U24444 (N_24444,N_21477,N_22267);
or U24445 (N_24445,N_21368,N_21959);
or U24446 (N_24446,N_21552,N_20878);
xor U24447 (N_24447,N_21741,N_20101);
or U24448 (N_24448,N_21087,N_22476);
or U24449 (N_24449,N_20826,N_20730);
nand U24450 (N_24450,N_21575,N_22000);
and U24451 (N_24451,N_21855,N_20127);
xnor U24452 (N_24452,N_20056,N_22403);
nand U24453 (N_24453,N_22429,N_20628);
xnor U24454 (N_24454,N_20664,N_21860);
xnor U24455 (N_24455,N_22359,N_22081);
nand U24456 (N_24456,N_20055,N_22103);
nand U24457 (N_24457,N_20337,N_20587);
and U24458 (N_24458,N_20702,N_21721);
or U24459 (N_24459,N_22031,N_21174);
and U24460 (N_24460,N_20166,N_20140);
and U24461 (N_24461,N_21199,N_21810);
xor U24462 (N_24462,N_20242,N_20489);
or U24463 (N_24463,N_22210,N_20992);
and U24464 (N_24464,N_22118,N_20005);
nand U24465 (N_24465,N_21825,N_21253);
nand U24466 (N_24466,N_20994,N_22189);
nor U24467 (N_24467,N_20966,N_21901);
xnor U24468 (N_24468,N_20801,N_21624);
or U24469 (N_24469,N_22384,N_20819);
and U24470 (N_24470,N_20260,N_20308);
nand U24471 (N_24471,N_20315,N_21034);
nor U24472 (N_24472,N_21911,N_21532);
or U24473 (N_24473,N_22494,N_20511);
nand U24474 (N_24474,N_21112,N_22418);
xnor U24475 (N_24475,N_20022,N_20827);
and U24476 (N_24476,N_21384,N_21683);
nor U24477 (N_24477,N_20540,N_20850);
and U24478 (N_24478,N_20413,N_21724);
nand U24479 (N_24479,N_22293,N_22110);
or U24480 (N_24480,N_20693,N_20095);
xnor U24481 (N_24481,N_20329,N_20092);
and U24482 (N_24482,N_22424,N_21465);
nor U24483 (N_24483,N_22303,N_20772);
xnor U24484 (N_24484,N_21783,N_20845);
and U24485 (N_24485,N_22224,N_21045);
and U24486 (N_24486,N_20708,N_21478);
xor U24487 (N_24487,N_21952,N_20740);
or U24488 (N_24488,N_21332,N_20560);
nor U24489 (N_24489,N_20962,N_20669);
xor U24490 (N_24490,N_22137,N_22265);
and U24491 (N_24491,N_20321,N_20129);
xnor U24492 (N_24492,N_20393,N_20835);
nand U24493 (N_24493,N_20160,N_21710);
nor U24494 (N_24494,N_20989,N_20438);
nand U24495 (N_24495,N_20211,N_20185);
nand U24496 (N_24496,N_20682,N_20063);
or U24497 (N_24497,N_20736,N_22174);
nand U24498 (N_24498,N_21042,N_20267);
nand U24499 (N_24499,N_20566,N_22206);
and U24500 (N_24500,N_21015,N_21774);
xnor U24501 (N_24501,N_22002,N_20489);
and U24502 (N_24502,N_22490,N_20236);
nor U24503 (N_24503,N_22366,N_22306);
or U24504 (N_24504,N_22398,N_21508);
nand U24505 (N_24505,N_22471,N_21767);
nor U24506 (N_24506,N_21964,N_20435);
and U24507 (N_24507,N_21335,N_20538);
nor U24508 (N_24508,N_22314,N_22036);
xor U24509 (N_24509,N_20426,N_21303);
nand U24510 (N_24510,N_21052,N_21318);
nand U24511 (N_24511,N_22175,N_20928);
nand U24512 (N_24512,N_21379,N_21377);
nor U24513 (N_24513,N_22043,N_22360);
nand U24514 (N_24514,N_21834,N_21038);
or U24515 (N_24515,N_22094,N_20859);
xor U24516 (N_24516,N_20448,N_20832);
nor U24517 (N_24517,N_21009,N_20609);
and U24518 (N_24518,N_21128,N_20361);
and U24519 (N_24519,N_21222,N_22170);
or U24520 (N_24520,N_22246,N_21848);
nand U24521 (N_24521,N_21048,N_21405);
xnor U24522 (N_24522,N_20251,N_21972);
nor U24523 (N_24523,N_21156,N_20802);
xor U24524 (N_24524,N_22490,N_21210);
nor U24525 (N_24525,N_21122,N_20595);
xnor U24526 (N_24526,N_20459,N_21691);
xor U24527 (N_24527,N_21835,N_21871);
nor U24528 (N_24528,N_22306,N_20912);
or U24529 (N_24529,N_21756,N_22254);
or U24530 (N_24530,N_20545,N_21305);
xnor U24531 (N_24531,N_20827,N_22313);
and U24532 (N_24532,N_22103,N_20928);
or U24533 (N_24533,N_21815,N_20724);
and U24534 (N_24534,N_21741,N_20009);
nor U24535 (N_24535,N_21412,N_20057);
xnor U24536 (N_24536,N_20661,N_20178);
and U24537 (N_24537,N_21820,N_20252);
or U24538 (N_24538,N_20346,N_20580);
xor U24539 (N_24539,N_20578,N_21739);
and U24540 (N_24540,N_21279,N_20746);
nor U24541 (N_24541,N_21612,N_20681);
nor U24542 (N_24542,N_20906,N_21380);
nand U24543 (N_24543,N_20958,N_20108);
nor U24544 (N_24544,N_20531,N_20702);
nor U24545 (N_24545,N_20828,N_21885);
xnor U24546 (N_24546,N_22165,N_21770);
and U24547 (N_24547,N_21912,N_20217);
xor U24548 (N_24548,N_20972,N_20710);
or U24549 (N_24549,N_21295,N_20720);
xor U24550 (N_24550,N_20111,N_21934);
or U24551 (N_24551,N_20471,N_20370);
and U24552 (N_24552,N_20463,N_20217);
xor U24553 (N_24553,N_21249,N_21414);
xnor U24554 (N_24554,N_21579,N_20471);
and U24555 (N_24555,N_21488,N_20297);
nor U24556 (N_24556,N_21329,N_21593);
nand U24557 (N_24557,N_20968,N_20635);
or U24558 (N_24558,N_21106,N_22221);
or U24559 (N_24559,N_20709,N_20890);
or U24560 (N_24560,N_20869,N_22263);
xnor U24561 (N_24561,N_21175,N_22115);
and U24562 (N_24562,N_20808,N_22193);
nor U24563 (N_24563,N_22140,N_22130);
or U24564 (N_24564,N_20595,N_20541);
or U24565 (N_24565,N_21184,N_20389);
nor U24566 (N_24566,N_20522,N_21650);
xnor U24567 (N_24567,N_20146,N_22053);
nand U24568 (N_24568,N_21134,N_21923);
xnor U24569 (N_24569,N_21534,N_20570);
and U24570 (N_24570,N_20843,N_21018);
and U24571 (N_24571,N_20113,N_22240);
nor U24572 (N_24572,N_21421,N_20745);
nor U24573 (N_24573,N_20076,N_21668);
xor U24574 (N_24574,N_20939,N_21752);
nor U24575 (N_24575,N_20545,N_22262);
nor U24576 (N_24576,N_22243,N_20791);
and U24577 (N_24577,N_22064,N_20697);
and U24578 (N_24578,N_21865,N_21538);
xnor U24579 (N_24579,N_20041,N_21558);
nand U24580 (N_24580,N_22332,N_21199);
nor U24581 (N_24581,N_21240,N_21028);
and U24582 (N_24582,N_20169,N_22427);
or U24583 (N_24583,N_21524,N_21374);
nor U24584 (N_24584,N_21032,N_22001);
nor U24585 (N_24585,N_21263,N_20773);
xnor U24586 (N_24586,N_20459,N_21538);
xnor U24587 (N_24587,N_20874,N_20549);
xnor U24588 (N_24588,N_21792,N_20288);
or U24589 (N_24589,N_22336,N_21280);
nand U24590 (N_24590,N_22468,N_21118);
xnor U24591 (N_24591,N_20249,N_21816);
xnor U24592 (N_24592,N_20401,N_21395);
and U24593 (N_24593,N_21159,N_21928);
and U24594 (N_24594,N_21117,N_20782);
nor U24595 (N_24595,N_20386,N_20841);
nor U24596 (N_24596,N_22431,N_20687);
nor U24597 (N_24597,N_20235,N_20513);
or U24598 (N_24598,N_22167,N_21067);
or U24599 (N_24599,N_22039,N_20754);
and U24600 (N_24600,N_22205,N_21209);
nor U24601 (N_24601,N_21934,N_21065);
nand U24602 (N_24602,N_20842,N_21597);
nor U24603 (N_24603,N_22168,N_20781);
nor U24604 (N_24604,N_22140,N_20256);
and U24605 (N_24605,N_21243,N_21080);
and U24606 (N_24606,N_21967,N_22008);
or U24607 (N_24607,N_20691,N_21053);
and U24608 (N_24608,N_21271,N_20826);
and U24609 (N_24609,N_21947,N_21032);
or U24610 (N_24610,N_21050,N_20586);
and U24611 (N_24611,N_21060,N_21828);
nand U24612 (N_24612,N_22015,N_20398);
or U24613 (N_24613,N_20936,N_20918);
or U24614 (N_24614,N_20438,N_21907);
nor U24615 (N_24615,N_20095,N_20247);
xor U24616 (N_24616,N_20295,N_21550);
and U24617 (N_24617,N_21444,N_22330);
and U24618 (N_24618,N_21122,N_20047);
and U24619 (N_24619,N_21839,N_22375);
xnor U24620 (N_24620,N_21898,N_20724);
nand U24621 (N_24621,N_20122,N_21025);
nor U24622 (N_24622,N_20091,N_22354);
or U24623 (N_24623,N_20193,N_22078);
nor U24624 (N_24624,N_22102,N_20020);
nor U24625 (N_24625,N_21568,N_21723);
or U24626 (N_24626,N_21589,N_20371);
nand U24627 (N_24627,N_21953,N_21201);
xor U24628 (N_24628,N_21613,N_22018);
or U24629 (N_24629,N_21658,N_20318);
and U24630 (N_24630,N_21729,N_21486);
nor U24631 (N_24631,N_21239,N_22424);
or U24632 (N_24632,N_21099,N_20464);
or U24633 (N_24633,N_20280,N_20324);
xor U24634 (N_24634,N_21401,N_20812);
nor U24635 (N_24635,N_20374,N_20331);
xnor U24636 (N_24636,N_20123,N_20331);
and U24637 (N_24637,N_20937,N_22241);
xor U24638 (N_24638,N_20435,N_22361);
nor U24639 (N_24639,N_21097,N_21004);
nor U24640 (N_24640,N_20785,N_20268);
xor U24641 (N_24641,N_22451,N_20108);
and U24642 (N_24642,N_22307,N_20571);
and U24643 (N_24643,N_20334,N_22342);
xnor U24644 (N_24644,N_20915,N_20664);
xnor U24645 (N_24645,N_22409,N_22152);
or U24646 (N_24646,N_21128,N_20987);
nand U24647 (N_24647,N_22021,N_20832);
nand U24648 (N_24648,N_22169,N_22134);
xnor U24649 (N_24649,N_22293,N_20278);
or U24650 (N_24650,N_22344,N_20866);
nor U24651 (N_24651,N_20279,N_21708);
nor U24652 (N_24652,N_21048,N_22379);
nand U24653 (N_24653,N_22013,N_21248);
and U24654 (N_24654,N_20247,N_21941);
and U24655 (N_24655,N_22470,N_21053);
xor U24656 (N_24656,N_20670,N_20505);
or U24657 (N_24657,N_22228,N_20696);
nor U24658 (N_24658,N_22194,N_20127);
or U24659 (N_24659,N_21803,N_21278);
and U24660 (N_24660,N_20564,N_21140);
and U24661 (N_24661,N_21110,N_20597);
nand U24662 (N_24662,N_21403,N_21695);
or U24663 (N_24663,N_20643,N_21717);
nand U24664 (N_24664,N_22010,N_21431);
nor U24665 (N_24665,N_21416,N_21233);
nor U24666 (N_24666,N_22356,N_22325);
and U24667 (N_24667,N_20327,N_20163);
and U24668 (N_24668,N_20610,N_21343);
nand U24669 (N_24669,N_21762,N_21727);
and U24670 (N_24670,N_20729,N_21816);
nor U24671 (N_24671,N_20961,N_20656);
nand U24672 (N_24672,N_22012,N_20474);
nor U24673 (N_24673,N_20969,N_20967);
nand U24674 (N_24674,N_22005,N_20435);
and U24675 (N_24675,N_22368,N_21100);
xnor U24676 (N_24676,N_21774,N_22181);
xnor U24677 (N_24677,N_22026,N_21721);
nor U24678 (N_24678,N_20094,N_22009);
nor U24679 (N_24679,N_22175,N_20644);
nand U24680 (N_24680,N_20150,N_21913);
or U24681 (N_24681,N_22229,N_20531);
nor U24682 (N_24682,N_22271,N_21786);
nand U24683 (N_24683,N_20618,N_21389);
xor U24684 (N_24684,N_21344,N_22054);
and U24685 (N_24685,N_22213,N_21374);
xnor U24686 (N_24686,N_21284,N_20245);
and U24687 (N_24687,N_20911,N_21634);
nor U24688 (N_24688,N_20673,N_22026);
or U24689 (N_24689,N_22224,N_21604);
and U24690 (N_24690,N_21673,N_21984);
and U24691 (N_24691,N_20941,N_20303);
xnor U24692 (N_24692,N_20537,N_21317);
nand U24693 (N_24693,N_21352,N_22424);
nand U24694 (N_24694,N_20576,N_20120);
and U24695 (N_24695,N_21180,N_21811);
nand U24696 (N_24696,N_21618,N_20565);
nand U24697 (N_24697,N_21182,N_21547);
nand U24698 (N_24698,N_21474,N_20941);
xor U24699 (N_24699,N_21324,N_21056);
nor U24700 (N_24700,N_22123,N_20628);
xnor U24701 (N_24701,N_21874,N_20873);
or U24702 (N_24702,N_22408,N_20429);
nand U24703 (N_24703,N_20612,N_21896);
and U24704 (N_24704,N_21718,N_21077);
or U24705 (N_24705,N_22427,N_20682);
nand U24706 (N_24706,N_20148,N_20770);
nor U24707 (N_24707,N_21112,N_21534);
xor U24708 (N_24708,N_21128,N_22446);
and U24709 (N_24709,N_20945,N_20935);
or U24710 (N_24710,N_20690,N_20939);
nand U24711 (N_24711,N_21316,N_22034);
and U24712 (N_24712,N_20510,N_22171);
nor U24713 (N_24713,N_21771,N_20903);
xor U24714 (N_24714,N_21611,N_21887);
or U24715 (N_24715,N_21335,N_21802);
or U24716 (N_24716,N_20192,N_20235);
and U24717 (N_24717,N_21123,N_21099);
or U24718 (N_24718,N_21652,N_20134);
or U24719 (N_24719,N_21714,N_20962);
or U24720 (N_24720,N_20221,N_21051);
xor U24721 (N_24721,N_20506,N_20451);
nor U24722 (N_24722,N_20464,N_21432);
and U24723 (N_24723,N_22056,N_20356);
or U24724 (N_24724,N_20824,N_22238);
and U24725 (N_24725,N_22483,N_20127);
xnor U24726 (N_24726,N_21754,N_20093);
and U24727 (N_24727,N_22102,N_20344);
nor U24728 (N_24728,N_20642,N_20712);
nand U24729 (N_24729,N_20516,N_20383);
xor U24730 (N_24730,N_22247,N_21286);
nor U24731 (N_24731,N_21314,N_20171);
xor U24732 (N_24732,N_21232,N_20103);
nand U24733 (N_24733,N_22039,N_20349);
nand U24734 (N_24734,N_21612,N_22064);
nand U24735 (N_24735,N_22249,N_21150);
and U24736 (N_24736,N_21731,N_20671);
nand U24737 (N_24737,N_20694,N_20877);
and U24738 (N_24738,N_22051,N_21532);
xor U24739 (N_24739,N_20502,N_21280);
or U24740 (N_24740,N_21052,N_21251);
and U24741 (N_24741,N_21344,N_20285);
nand U24742 (N_24742,N_21648,N_21695);
and U24743 (N_24743,N_21481,N_22325);
nand U24744 (N_24744,N_20476,N_20074);
xor U24745 (N_24745,N_22345,N_20651);
nand U24746 (N_24746,N_20136,N_22439);
or U24747 (N_24747,N_20384,N_22486);
xnor U24748 (N_24748,N_20371,N_21641);
and U24749 (N_24749,N_20504,N_20666);
nand U24750 (N_24750,N_20047,N_21349);
nand U24751 (N_24751,N_21487,N_22065);
xor U24752 (N_24752,N_20547,N_21300);
nor U24753 (N_24753,N_21361,N_20307);
xor U24754 (N_24754,N_21603,N_21643);
xnor U24755 (N_24755,N_21177,N_22280);
xor U24756 (N_24756,N_20395,N_20987);
xor U24757 (N_24757,N_22430,N_20958);
nor U24758 (N_24758,N_20663,N_21325);
or U24759 (N_24759,N_20203,N_21911);
xor U24760 (N_24760,N_22042,N_22281);
xor U24761 (N_24761,N_21218,N_20154);
xnor U24762 (N_24762,N_22083,N_21186);
nand U24763 (N_24763,N_21222,N_20093);
nor U24764 (N_24764,N_20527,N_22311);
nor U24765 (N_24765,N_21494,N_21931);
xnor U24766 (N_24766,N_20189,N_21300);
xor U24767 (N_24767,N_20282,N_22495);
nand U24768 (N_24768,N_20004,N_20357);
nor U24769 (N_24769,N_20724,N_20098);
nand U24770 (N_24770,N_21722,N_22287);
nor U24771 (N_24771,N_21282,N_20962);
and U24772 (N_24772,N_20646,N_20235);
nor U24773 (N_24773,N_21476,N_21602);
xor U24774 (N_24774,N_22073,N_20568);
or U24775 (N_24775,N_20679,N_20557);
nor U24776 (N_24776,N_21854,N_22486);
and U24777 (N_24777,N_21573,N_21378);
nor U24778 (N_24778,N_21394,N_20346);
xnor U24779 (N_24779,N_21705,N_20540);
xor U24780 (N_24780,N_20820,N_21146);
and U24781 (N_24781,N_21103,N_20559);
and U24782 (N_24782,N_21566,N_21385);
or U24783 (N_24783,N_21018,N_22371);
or U24784 (N_24784,N_21648,N_22177);
or U24785 (N_24785,N_21053,N_21645);
nor U24786 (N_24786,N_21501,N_20286);
xnor U24787 (N_24787,N_21195,N_22229);
or U24788 (N_24788,N_21178,N_20678);
nand U24789 (N_24789,N_21468,N_20565);
nand U24790 (N_24790,N_20351,N_20284);
xnor U24791 (N_24791,N_20653,N_21024);
nor U24792 (N_24792,N_22038,N_22387);
or U24793 (N_24793,N_21815,N_20538);
xnor U24794 (N_24794,N_21012,N_20938);
or U24795 (N_24795,N_21857,N_22227);
xnor U24796 (N_24796,N_22016,N_22080);
and U24797 (N_24797,N_21569,N_20248);
and U24798 (N_24798,N_22157,N_21410);
nor U24799 (N_24799,N_21821,N_20557);
xnor U24800 (N_24800,N_20058,N_20541);
xnor U24801 (N_24801,N_22123,N_22064);
nor U24802 (N_24802,N_20075,N_20410);
and U24803 (N_24803,N_21674,N_21022);
xor U24804 (N_24804,N_21755,N_21026);
xor U24805 (N_24805,N_21837,N_20847);
or U24806 (N_24806,N_22453,N_21665);
nand U24807 (N_24807,N_22218,N_21587);
nand U24808 (N_24808,N_20684,N_20379);
and U24809 (N_24809,N_21141,N_21023);
xor U24810 (N_24810,N_22180,N_20109);
and U24811 (N_24811,N_21272,N_20890);
nand U24812 (N_24812,N_21646,N_20525);
xnor U24813 (N_24813,N_21388,N_20755);
or U24814 (N_24814,N_21735,N_22482);
and U24815 (N_24815,N_20238,N_20675);
or U24816 (N_24816,N_21102,N_20699);
and U24817 (N_24817,N_20824,N_21496);
nor U24818 (N_24818,N_21744,N_21223);
and U24819 (N_24819,N_20873,N_21384);
nor U24820 (N_24820,N_21023,N_22006);
nand U24821 (N_24821,N_20557,N_21763);
nand U24822 (N_24822,N_21720,N_21263);
nand U24823 (N_24823,N_20865,N_21927);
or U24824 (N_24824,N_20955,N_20295);
nand U24825 (N_24825,N_20781,N_22355);
nor U24826 (N_24826,N_21660,N_20382);
nor U24827 (N_24827,N_21001,N_21244);
and U24828 (N_24828,N_20138,N_21810);
xor U24829 (N_24829,N_20117,N_20459);
xor U24830 (N_24830,N_21744,N_20354);
and U24831 (N_24831,N_20348,N_21747);
nand U24832 (N_24832,N_20282,N_22164);
and U24833 (N_24833,N_20696,N_22411);
or U24834 (N_24834,N_20173,N_20239);
and U24835 (N_24835,N_21437,N_21121);
xor U24836 (N_24836,N_22048,N_21330);
nor U24837 (N_24837,N_21008,N_21129);
nor U24838 (N_24838,N_20076,N_21630);
nand U24839 (N_24839,N_21690,N_21851);
and U24840 (N_24840,N_20016,N_21873);
and U24841 (N_24841,N_20757,N_22301);
or U24842 (N_24842,N_21100,N_21676);
nand U24843 (N_24843,N_22080,N_20240);
or U24844 (N_24844,N_22386,N_20928);
xnor U24845 (N_24845,N_22378,N_21604);
nor U24846 (N_24846,N_21510,N_21977);
or U24847 (N_24847,N_22044,N_20588);
and U24848 (N_24848,N_20176,N_21057);
and U24849 (N_24849,N_21361,N_21424);
and U24850 (N_24850,N_20307,N_22435);
nand U24851 (N_24851,N_22263,N_22371);
xnor U24852 (N_24852,N_20524,N_22310);
nand U24853 (N_24853,N_22493,N_22164);
nand U24854 (N_24854,N_20437,N_21507);
nand U24855 (N_24855,N_21305,N_22232);
nand U24856 (N_24856,N_21162,N_22028);
xor U24857 (N_24857,N_21007,N_21141);
or U24858 (N_24858,N_21421,N_21874);
nand U24859 (N_24859,N_20180,N_21244);
or U24860 (N_24860,N_22351,N_20329);
nand U24861 (N_24861,N_20858,N_21125);
and U24862 (N_24862,N_20461,N_20952);
xnor U24863 (N_24863,N_20289,N_20510);
and U24864 (N_24864,N_21556,N_20652);
or U24865 (N_24865,N_21851,N_20636);
and U24866 (N_24866,N_20574,N_21241);
or U24867 (N_24867,N_22445,N_21579);
and U24868 (N_24868,N_21727,N_21038);
nand U24869 (N_24869,N_20364,N_21542);
nand U24870 (N_24870,N_20354,N_20920);
or U24871 (N_24871,N_22304,N_22498);
xnor U24872 (N_24872,N_21755,N_21479);
xor U24873 (N_24873,N_21249,N_20284);
and U24874 (N_24874,N_20845,N_21273);
nor U24875 (N_24875,N_20046,N_22232);
nor U24876 (N_24876,N_22181,N_22300);
nor U24877 (N_24877,N_20954,N_22176);
nand U24878 (N_24878,N_20654,N_22012);
or U24879 (N_24879,N_21694,N_22366);
xnor U24880 (N_24880,N_21575,N_20410);
and U24881 (N_24881,N_21110,N_20030);
or U24882 (N_24882,N_20852,N_20053);
or U24883 (N_24883,N_20814,N_20165);
xnor U24884 (N_24884,N_21802,N_22118);
and U24885 (N_24885,N_21366,N_21216);
xor U24886 (N_24886,N_21406,N_20997);
and U24887 (N_24887,N_21474,N_22470);
nand U24888 (N_24888,N_22081,N_21937);
or U24889 (N_24889,N_21639,N_21357);
and U24890 (N_24890,N_22098,N_22462);
nand U24891 (N_24891,N_21728,N_20551);
and U24892 (N_24892,N_20695,N_22248);
xor U24893 (N_24893,N_22227,N_20963);
or U24894 (N_24894,N_20345,N_20295);
and U24895 (N_24895,N_20348,N_21348);
or U24896 (N_24896,N_21493,N_21864);
or U24897 (N_24897,N_21716,N_22099);
nand U24898 (N_24898,N_21197,N_20552);
and U24899 (N_24899,N_20786,N_21073);
and U24900 (N_24900,N_20711,N_20501);
and U24901 (N_24901,N_20455,N_21946);
xnor U24902 (N_24902,N_20719,N_20950);
xnor U24903 (N_24903,N_22447,N_21156);
and U24904 (N_24904,N_20881,N_22423);
nor U24905 (N_24905,N_21796,N_22466);
or U24906 (N_24906,N_21598,N_20918);
or U24907 (N_24907,N_22422,N_20990);
and U24908 (N_24908,N_22435,N_20336);
xor U24909 (N_24909,N_21638,N_21420);
and U24910 (N_24910,N_22029,N_21280);
nand U24911 (N_24911,N_20022,N_21526);
nor U24912 (N_24912,N_21685,N_20730);
and U24913 (N_24913,N_22454,N_20207);
or U24914 (N_24914,N_21046,N_22316);
nand U24915 (N_24915,N_22390,N_21798);
xor U24916 (N_24916,N_22207,N_21607);
nand U24917 (N_24917,N_20983,N_20099);
xor U24918 (N_24918,N_21577,N_21497);
nor U24919 (N_24919,N_21132,N_21300);
xor U24920 (N_24920,N_22474,N_20375);
nor U24921 (N_24921,N_20323,N_20997);
and U24922 (N_24922,N_20756,N_21487);
nor U24923 (N_24923,N_20103,N_20721);
nand U24924 (N_24924,N_21905,N_21587);
xnor U24925 (N_24925,N_20367,N_20518);
and U24926 (N_24926,N_21776,N_20718);
and U24927 (N_24927,N_21059,N_20866);
xor U24928 (N_24928,N_20978,N_22161);
or U24929 (N_24929,N_21186,N_21703);
nand U24930 (N_24930,N_20270,N_21792);
or U24931 (N_24931,N_20747,N_20858);
nor U24932 (N_24932,N_20681,N_21418);
and U24933 (N_24933,N_21402,N_22155);
nand U24934 (N_24934,N_21394,N_20483);
and U24935 (N_24935,N_20577,N_20222);
nand U24936 (N_24936,N_21290,N_22294);
and U24937 (N_24937,N_21492,N_22157);
or U24938 (N_24938,N_20566,N_20485);
nand U24939 (N_24939,N_21877,N_22453);
xnor U24940 (N_24940,N_20431,N_20764);
nor U24941 (N_24941,N_21281,N_21768);
or U24942 (N_24942,N_20830,N_21299);
xor U24943 (N_24943,N_22139,N_20161);
and U24944 (N_24944,N_21784,N_22279);
nand U24945 (N_24945,N_20681,N_20699);
nor U24946 (N_24946,N_22294,N_21475);
xnor U24947 (N_24947,N_22129,N_20478);
xor U24948 (N_24948,N_21330,N_21304);
xnor U24949 (N_24949,N_21847,N_22418);
nor U24950 (N_24950,N_20670,N_22317);
and U24951 (N_24951,N_21639,N_20843);
xnor U24952 (N_24952,N_22184,N_20153);
nor U24953 (N_24953,N_21442,N_20652);
or U24954 (N_24954,N_20011,N_20260);
and U24955 (N_24955,N_20962,N_21646);
and U24956 (N_24956,N_20400,N_21025);
or U24957 (N_24957,N_22070,N_20989);
and U24958 (N_24958,N_22208,N_21265);
and U24959 (N_24959,N_22071,N_20718);
nand U24960 (N_24960,N_20360,N_20442);
nand U24961 (N_24961,N_21621,N_20204);
xnor U24962 (N_24962,N_22002,N_20937);
and U24963 (N_24963,N_22225,N_20193);
nand U24964 (N_24964,N_21872,N_20117);
and U24965 (N_24965,N_22296,N_20965);
nor U24966 (N_24966,N_20953,N_21672);
xnor U24967 (N_24967,N_20791,N_20952);
xnor U24968 (N_24968,N_21709,N_21584);
and U24969 (N_24969,N_22258,N_22222);
and U24970 (N_24970,N_21759,N_20063);
xnor U24971 (N_24971,N_20783,N_20088);
and U24972 (N_24972,N_21969,N_21926);
nand U24973 (N_24973,N_20110,N_20341);
nand U24974 (N_24974,N_21996,N_21224);
nor U24975 (N_24975,N_22259,N_20079);
xnor U24976 (N_24976,N_21825,N_20781);
or U24977 (N_24977,N_21262,N_21331);
nor U24978 (N_24978,N_21757,N_21511);
xnor U24979 (N_24979,N_20299,N_21118);
nor U24980 (N_24980,N_21088,N_20319);
xnor U24981 (N_24981,N_20500,N_22248);
or U24982 (N_24982,N_20734,N_22127);
or U24983 (N_24983,N_22359,N_20573);
nand U24984 (N_24984,N_20853,N_22444);
nand U24985 (N_24985,N_21534,N_20448);
nand U24986 (N_24986,N_22099,N_22283);
or U24987 (N_24987,N_22498,N_20358);
nand U24988 (N_24988,N_20898,N_20518);
and U24989 (N_24989,N_21660,N_21316);
xor U24990 (N_24990,N_22001,N_22485);
or U24991 (N_24991,N_21723,N_20390);
xnor U24992 (N_24992,N_21419,N_21995);
and U24993 (N_24993,N_21903,N_20816);
nor U24994 (N_24994,N_21638,N_22364);
xor U24995 (N_24995,N_21541,N_20049);
nand U24996 (N_24996,N_22247,N_20344);
nand U24997 (N_24997,N_21365,N_21030);
nand U24998 (N_24998,N_21538,N_20679);
xor U24999 (N_24999,N_20103,N_21512);
nand U25000 (N_25000,N_24859,N_24827);
and U25001 (N_25001,N_23794,N_24573);
or U25002 (N_25002,N_23524,N_24338);
nor U25003 (N_25003,N_24000,N_24942);
nor U25004 (N_25004,N_23217,N_24111);
nor U25005 (N_25005,N_24253,N_22608);
and U25006 (N_25006,N_22819,N_24516);
nand U25007 (N_25007,N_24985,N_22615);
nor U25008 (N_25008,N_23955,N_23812);
or U25009 (N_25009,N_23868,N_23537);
or U25010 (N_25010,N_24416,N_23791);
xor U25011 (N_25011,N_23765,N_22523);
and U25012 (N_25012,N_24280,N_22578);
xnor U25013 (N_25013,N_23725,N_23432);
xnor U25014 (N_25014,N_22740,N_24397);
and U25015 (N_25015,N_24854,N_23134);
or U25016 (N_25016,N_24479,N_23672);
nor U25017 (N_25017,N_24410,N_24939);
nor U25018 (N_25018,N_24222,N_23427);
nand U25019 (N_25019,N_23161,N_23856);
or U25020 (N_25020,N_24219,N_24216);
nor U25021 (N_25021,N_23169,N_23355);
nor U25022 (N_25022,N_23899,N_24078);
or U25023 (N_25023,N_24190,N_23224);
or U25024 (N_25024,N_22911,N_23942);
nor U25025 (N_25025,N_24169,N_23944);
xnor U25026 (N_25026,N_24591,N_23552);
nand U25027 (N_25027,N_24242,N_22513);
or U25028 (N_25028,N_22734,N_24756);
and U25029 (N_25029,N_22776,N_23421);
and U25030 (N_25030,N_23632,N_23097);
nor U25031 (N_25031,N_23437,N_23888);
xor U25032 (N_25032,N_24973,N_24692);
and U25033 (N_25033,N_22864,N_24911);
or U25034 (N_25034,N_23368,N_24173);
nand U25035 (N_25035,N_22573,N_23068);
nor U25036 (N_25036,N_23860,N_23153);
xnor U25037 (N_25037,N_23016,N_23685);
or U25038 (N_25038,N_22759,N_24440);
nor U25039 (N_25039,N_23830,N_24131);
nand U25040 (N_25040,N_22801,N_23814);
xnor U25041 (N_25041,N_23608,N_24370);
nand U25042 (N_25042,N_23138,N_22550);
nand U25043 (N_25043,N_23444,N_24639);
nor U25044 (N_25044,N_22521,N_22793);
or U25045 (N_25045,N_23197,N_24200);
or U25046 (N_25046,N_23542,N_24385);
or U25047 (N_25047,N_24977,N_24503);
nor U25048 (N_25048,N_23329,N_24753);
xor U25049 (N_25049,N_23648,N_23879);
xor U25050 (N_25050,N_24777,N_24271);
nand U25051 (N_25051,N_22913,N_22874);
xnor U25052 (N_25052,N_22947,N_23350);
nor U25053 (N_25053,N_24109,N_23757);
nor U25054 (N_25054,N_23460,N_23715);
nand U25055 (N_25055,N_22824,N_24912);
xnor U25056 (N_25056,N_24733,N_22748);
and U25057 (N_25057,N_24134,N_23305);
or U25058 (N_25058,N_23494,N_22778);
nor U25059 (N_25059,N_23146,N_24436);
and U25060 (N_25060,N_23484,N_24211);
xor U25061 (N_25061,N_24629,N_23095);
or U25062 (N_25062,N_24090,N_23967);
and U25063 (N_25063,N_23292,N_24940);
nor U25064 (N_25064,N_24158,N_24205);
or U25065 (N_25065,N_23275,N_22587);
or U25066 (N_25066,N_24027,N_23324);
or U25067 (N_25067,N_23042,N_24605);
nor U25068 (N_25068,N_23160,N_24291);
and U25069 (N_25069,N_24540,N_24059);
nand U25070 (N_25070,N_23144,N_24630);
nor U25071 (N_25071,N_22526,N_24313);
xnor U25072 (N_25072,N_22943,N_22939);
and U25073 (N_25073,N_24672,N_24582);
and U25074 (N_25074,N_22690,N_23020);
nor U25075 (N_25075,N_23583,N_24910);
nor U25076 (N_25076,N_24054,N_22953);
xnor U25077 (N_25077,N_24818,N_24719);
nor U25078 (N_25078,N_24862,N_23943);
nor U25079 (N_25079,N_23154,N_24956);
xor U25080 (N_25080,N_23807,N_23049);
or U25081 (N_25081,N_24126,N_24736);
nand U25082 (N_25082,N_23553,N_24043);
and U25083 (N_25083,N_23591,N_24673);
or U25084 (N_25084,N_23993,N_23257);
nand U25085 (N_25085,N_22955,N_24287);
nand U25086 (N_25086,N_22525,N_22832);
nand U25087 (N_25087,N_22685,N_23143);
xor U25088 (N_25088,N_23239,N_24607);
and U25089 (N_25089,N_23587,N_24814);
and U25090 (N_25090,N_22678,N_23266);
nand U25091 (N_25091,N_23433,N_24441);
xnor U25092 (N_25092,N_24514,N_24895);
xor U25093 (N_25093,N_23914,N_22940);
and U25094 (N_25094,N_24524,N_23036);
nor U25095 (N_25095,N_23751,N_22712);
xnor U25096 (N_25096,N_24567,N_24921);
and U25097 (N_25097,N_23237,N_24218);
or U25098 (N_25098,N_23832,N_23697);
xnor U25099 (N_25099,N_24909,N_24010);
nor U25100 (N_25100,N_24477,N_24473);
xor U25101 (N_25101,N_22956,N_22806);
nand U25102 (N_25102,N_23392,N_23195);
or U25103 (N_25103,N_24778,N_24716);
or U25104 (N_25104,N_24206,N_22975);
or U25105 (N_25105,N_23530,N_23130);
or U25106 (N_25106,N_24933,N_24641);
xor U25107 (N_25107,N_24492,N_23098);
nor U25108 (N_25108,N_23376,N_22727);
xnor U25109 (N_25109,N_24847,N_23935);
and U25110 (N_25110,N_23182,N_23582);
nand U25111 (N_25111,N_24358,N_23528);
and U25112 (N_25112,N_23414,N_23459);
and U25113 (N_25113,N_24668,N_23829);
nor U25114 (N_25114,N_24915,N_22950);
and U25115 (N_25115,N_22596,N_24811);
xor U25116 (N_25116,N_23615,N_24214);
xor U25117 (N_25117,N_24678,N_23395);
or U25118 (N_25118,N_24596,N_23145);
and U25119 (N_25119,N_23311,N_24870);
and U25120 (N_25120,N_23901,N_23453);
nor U25121 (N_25121,N_24504,N_22559);
and U25122 (N_25122,N_24741,N_24030);
and U25123 (N_25123,N_24293,N_24715);
or U25124 (N_25124,N_23805,N_23096);
xor U25125 (N_25125,N_22898,N_24860);
nand U25126 (N_25126,N_23880,N_24331);
and U25127 (N_25127,N_24693,N_22630);
or U25128 (N_25128,N_22610,N_23842);
nor U25129 (N_25129,N_24375,N_22612);
or U25130 (N_25130,N_22676,N_23649);
nor U25131 (N_25131,N_23398,N_24355);
nor U25132 (N_25132,N_23164,N_22501);
or U25133 (N_25133,N_24459,N_22570);
xnor U25134 (N_25134,N_24257,N_23597);
or U25135 (N_25135,N_22538,N_24978);
and U25136 (N_25136,N_23917,N_23304);
xnor U25137 (N_25137,N_23462,N_24664);
or U25138 (N_25138,N_23560,N_23293);
xor U25139 (N_25139,N_24703,N_22990);
nand U25140 (N_25140,N_23319,N_24137);
nor U25141 (N_25141,N_22873,N_22901);
or U25142 (N_25142,N_24241,N_23354);
or U25143 (N_25143,N_23902,N_24974);
and U25144 (N_25144,N_24221,N_23698);
or U25145 (N_25145,N_23924,N_23541);
xor U25146 (N_25146,N_23823,N_22849);
or U25147 (N_25147,N_23442,N_23385);
nor U25148 (N_25148,N_23473,N_22771);
nand U25149 (N_25149,N_24725,N_23105);
and U25150 (N_25150,N_23334,N_22962);
xnor U25151 (N_25151,N_24101,N_23115);
nor U25152 (N_25152,N_22772,N_24277);
nor U25153 (N_25153,N_22731,N_23107);
xnor U25154 (N_25154,N_24770,N_22633);
and U25155 (N_25155,N_22826,N_24553);
nand U25156 (N_25156,N_24143,N_23526);
nor U25157 (N_25157,N_24651,N_24275);
and U25158 (N_25158,N_23635,N_23236);
nor U25159 (N_25159,N_24944,N_23147);
nor U25160 (N_25160,N_24543,N_22683);
nor U25161 (N_25161,N_23116,N_22909);
and U25162 (N_25162,N_24259,N_23041);
and U25163 (N_25163,N_23710,N_24129);
nor U25164 (N_25164,N_22507,N_22841);
xnor U25165 (N_25165,N_24835,N_23844);
nor U25166 (N_25166,N_24794,N_22858);
nor U25167 (N_25167,N_22511,N_23780);
xor U25168 (N_25168,N_24759,N_23282);
and U25169 (N_25169,N_23203,N_24527);
and U25170 (N_25170,N_23678,N_24658);
or U25171 (N_25171,N_22620,N_23731);
nand U25172 (N_25172,N_23847,N_23643);
nor U25173 (N_25173,N_22992,N_24743);
or U25174 (N_25174,N_23746,N_24157);
and U25175 (N_25175,N_23288,N_24614);
or U25176 (N_25176,N_24979,N_24633);
xnor U25177 (N_25177,N_23216,N_24491);
nor U25178 (N_25178,N_22613,N_23506);
nand U25179 (N_25179,N_24718,N_24768);
and U25180 (N_25180,N_22800,N_23483);
or U25181 (N_25181,N_23656,N_24426);
nand U25182 (N_25182,N_24676,N_24339);
xnor U25183 (N_25183,N_22694,N_23843);
nand U25184 (N_25184,N_24976,N_22605);
and U25185 (N_25185,N_23492,N_22998);
and U25186 (N_25186,N_24579,N_22933);
and U25187 (N_25187,N_24738,N_23748);
or U25188 (N_25188,N_23362,N_24040);
and U25189 (N_25189,N_23638,N_24354);
and U25190 (N_25190,N_24082,N_22805);
nor U25191 (N_25191,N_24904,N_24493);
and U25192 (N_25192,N_23119,N_22838);
nor U25193 (N_25193,N_24168,N_24024);
and U25194 (N_25194,N_22624,N_23665);
or U25195 (N_25195,N_24992,N_24038);
xor U25196 (N_25196,N_23776,N_24728);
nor U25197 (N_25197,N_24954,N_24993);
xnor U25198 (N_25198,N_24807,N_23796);
nor U25199 (N_25199,N_22946,N_24379);
nor U25200 (N_25200,N_23332,N_24212);
nand U25201 (N_25201,N_24531,N_24826);
nand U25202 (N_25202,N_23808,N_23787);
and U25203 (N_25203,N_22653,N_23007);
xnor U25204 (N_25204,N_23799,N_22686);
nor U25205 (N_25205,N_24470,N_22815);
and U25206 (N_25206,N_24505,N_24347);
nor U25207 (N_25207,N_23185,N_24453);
nand U25208 (N_25208,N_24843,N_24310);
or U25209 (N_25209,N_23610,N_23853);
nand U25210 (N_25210,N_23015,N_24273);
nor U25211 (N_25211,N_24717,N_23439);
nor U25212 (N_25212,N_23269,N_22662);
nand U25213 (N_25213,N_24618,N_22867);
or U25214 (N_25214,N_22958,N_24930);
and U25215 (N_25215,N_24866,N_22660);
and U25216 (N_25216,N_22986,N_23858);
and U25217 (N_25217,N_22546,N_23106);
xor U25218 (N_25218,N_23629,N_24266);
nand U25219 (N_25219,N_23574,N_22517);
xnor U25220 (N_25220,N_23060,N_22606);
xor U25221 (N_25221,N_23152,N_22993);
nand U25222 (N_25222,N_24946,N_24822);
nand U25223 (N_25223,N_24653,N_23864);
and U25224 (N_25224,N_24346,N_24029);
xor U25225 (N_25225,N_24194,N_23463);
or U25226 (N_25226,N_23579,N_23733);
or U25227 (N_25227,N_23131,N_23456);
xnor U25228 (N_25228,N_23214,N_24398);
or U25229 (N_25229,N_23085,N_23268);
xor U25230 (N_25230,N_22965,N_23838);
or U25231 (N_25231,N_24447,N_23002);
and U25232 (N_25232,N_24467,N_23947);
nand U25233 (N_25233,N_23906,N_24230);
nand U25234 (N_25234,N_23309,N_24550);
nor U25235 (N_25235,N_24886,N_23938);
and U25236 (N_25236,N_24409,N_23952);
nor U25237 (N_25237,N_22903,N_24274);
nand U25238 (N_25238,N_24456,N_23622);
nor U25239 (N_25239,N_24463,N_24051);
and U25240 (N_25240,N_24305,N_24971);
nor U25241 (N_25241,N_24279,N_22941);
nor U25242 (N_25242,N_23065,N_24713);
or U25243 (N_25243,N_24431,N_24041);
and U25244 (N_25244,N_22961,N_22899);
and U25245 (N_25245,N_24314,N_24751);
and U25246 (N_25246,N_23310,N_23979);
nor U25247 (N_25247,N_24989,N_23990);
xnor U25248 (N_25248,N_22549,N_23531);
and U25249 (N_25249,N_24581,N_23170);
xnor U25250 (N_25250,N_23986,N_23230);
or U25251 (N_25251,N_23254,N_23692);
xnor U25252 (N_25252,N_24711,N_22652);
xor U25253 (N_25253,N_24649,N_23274);
or U25254 (N_25254,N_23148,N_22808);
xor U25255 (N_25255,N_22807,N_22700);
nor U25256 (N_25256,N_24325,N_24892);
nand U25257 (N_25257,N_24709,N_24003);
and U25258 (N_25258,N_24695,N_22739);
nor U25259 (N_25259,N_23504,N_23301);
xor U25260 (N_25260,N_22580,N_24351);
nand U25261 (N_25261,N_24154,N_23669);
or U25262 (N_25262,N_23207,N_24964);
nor U25263 (N_25263,N_23894,N_24813);
nand U25264 (N_25264,N_24675,N_23364);
and U25265 (N_25265,N_23684,N_24320);
or U25266 (N_25266,N_22868,N_24302);
nor U25267 (N_25267,N_24850,N_22904);
and U25268 (N_25268,N_24619,N_24642);
nand U25269 (N_25269,N_22637,N_24622);
and U25270 (N_25270,N_22619,N_23509);
nor U25271 (N_25271,N_22649,N_23871);
nor U25272 (N_25272,N_22905,N_23194);
and U25273 (N_25273,N_24660,N_23937);
nand U25274 (N_25274,N_23486,N_22856);
xor U25275 (N_25275,N_23175,N_24311);
or U25276 (N_25276,N_23136,N_23229);
xor U25277 (N_25277,N_24704,N_24654);
xor U25278 (N_25278,N_24262,N_23886);
nor U25279 (N_25279,N_22894,N_24153);
or U25280 (N_25280,N_23777,N_22750);
or U25281 (N_25281,N_23718,N_23074);
and U25282 (N_25282,N_22522,N_24833);
and U25283 (N_25283,N_24900,N_23455);
and U25284 (N_25284,N_23353,N_24335);
or U25285 (N_25285,N_24585,N_24487);
nand U25286 (N_25286,N_22846,N_24421);
and U25287 (N_25287,N_23225,N_23916);
xnor U25288 (N_25288,N_23601,N_23032);
and U25289 (N_25289,N_22921,N_23186);
nor U25290 (N_25290,N_24472,N_24737);
and U25291 (N_25291,N_24445,N_23763);
xnor U25292 (N_25292,N_23682,N_24094);
nand U25293 (N_25293,N_24250,N_24840);
nor U25294 (N_25294,N_23448,N_23501);
nor U25295 (N_25295,N_24799,N_22591);
nor U25296 (N_25296,N_23910,N_23854);
xor U25297 (N_25297,N_23277,N_24106);
or U25298 (N_25298,N_22770,N_24975);
xnor U25299 (N_25299,N_24369,N_23641);
nand U25300 (N_25300,N_24970,N_24880);
or U25301 (N_25301,N_24851,N_24967);
xnor U25302 (N_25302,N_22803,N_24981);
xor U25303 (N_25303,N_24261,N_24511);
xnor U25304 (N_25304,N_23975,N_24239);
xnor U25305 (N_25305,N_24730,N_23800);
nand U25306 (N_25306,N_24044,N_24202);
or U25307 (N_25307,N_23768,N_24837);
and U25308 (N_25308,N_23845,N_23245);
and U25309 (N_25309,N_23837,N_23810);
xor U25310 (N_25310,N_23778,N_24571);
or U25311 (N_25311,N_23365,N_22987);
and U25312 (N_25312,N_23171,N_22812);
xnor U25313 (N_25313,N_24532,N_23966);
or U25314 (N_25314,N_24958,N_23781);
and U25315 (N_25315,N_24136,N_23846);
and U25316 (N_25316,N_23464,N_23892);
or U25317 (N_25317,N_22635,N_23034);
and U25318 (N_25318,N_24902,N_23936);
nor U25319 (N_25319,N_24080,N_23720);
xor U25320 (N_25320,N_24742,N_23836);
and U25321 (N_25321,N_23030,N_24008);
nand U25322 (N_25322,N_23811,N_22818);
nand U25323 (N_25323,N_24545,N_24175);
xnor U25324 (N_25324,N_24914,N_23828);
and U25325 (N_25325,N_22566,N_23806);
or U25326 (N_25326,N_23256,N_24663);
nor U25327 (N_25327,N_23430,N_22680);
or U25328 (N_25328,N_23103,N_23358);
or U25329 (N_25329,N_22688,N_23278);
xnor U25330 (N_25330,N_23037,N_23928);
xor U25331 (N_25331,N_23485,N_23387);
nor U25332 (N_25332,N_22758,N_23525);
xor U25333 (N_25333,N_23381,N_22532);
and U25334 (N_25334,N_24036,N_22543);
nor U25335 (N_25335,N_24359,N_24986);
xnor U25336 (N_25336,N_24923,N_23918);
and U25337 (N_25337,N_24110,N_24365);
nor U25338 (N_25338,N_23699,N_23613);
and U25339 (N_25339,N_24712,N_22707);
xor U25340 (N_25340,N_23227,N_23571);
or U25341 (N_25341,N_23407,N_24072);
nand U25342 (N_25342,N_24443,N_23080);
xor U25343 (N_25343,N_24330,N_23294);
or U25344 (N_25344,N_23188,N_24011);
or U25345 (N_25345,N_23921,N_24118);
nor U25346 (N_25346,N_23729,N_22879);
nor U25347 (N_25347,N_22565,N_23951);
and U25348 (N_25348,N_22720,N_24417);
or U25349 (N_25349,N_24179,N_24052);
or U25350 (N_25350,N_24662,N_23945);
nor U25351 (N_25351,N_22969,N_22972);
nand U25352 (N_25352,N_23544,N_24322);
or U25353 (N_25353,N_23258,N_23403);
nand U25354 (N_25354,N_24983,N_23389);
nor U25355 (N_25355,N_24522,N_22840);
nor U25356 (N_25356,N_24210,N_23576);
and U25357 (N_25357,N_23200,N_23084);
xor U25358 (N_25358,N_23673,N_23140);
or U25359 (N_25359,N_24195,N_23420);
or U25360 (N_25360,N_24708,N_24382);
or U25361 (N_25361,N_24005,N_22974);
and U25362 (N_25362,N_23912,N_24523);
nand U25363 (N_25363,N_23377,N_22675);
and U25364 (N_25364,N_23046,N_24317);
or U25365 (N_25365,N_24217,N_24296);
nor U25366 (N_25366,N_24035,N_23862);
nor U25367 (N_25367,N_24160,N_23409);
nand U25368 (N_25368,N_23510,N_24601);
or U25369 (N_25369,N_22670,N_22790);
xnor U25370 (N_25370,N_23356,N_23003);
xnor U25371 (N_25371,N_22533,N_22666);
xor U25372 (N_25372,N_22945,N_22509);
xnor U25373 (N_25373,N_23336,N_22908);
nor U25374 (N_25374,N_23434,N_23428);
and U25375 (N_25375,N_24181,N_24161);
and U25376 (N_25376,N_23331,N_23066);
nor U25377 (N_25377,N_24513,N_24509);
and U25378 (N_25378,N_23663,N_22744);
xnor U25379 (N_25379,N_24433,N_24095);
nand U25380 (N_25380,N_23999,N_22892);
nor U25381 (N_25381,N_24114,N_22985);
and U25382 (N_25382,N_23991,N_24411);
nor U25383 (N_25383,N_23840,N_24931);
nand U25384 (N_25384,N_24105,N_22855);
nand U25385 (N_25385,N_23841,N_23686);
nor U25386 (N_25386,N_23543,N_24739);
and U25387 (N_25387,N_24427,N_24278);
or U25388 (N_25388,N_22561,N_23750);
nor U25389 (N_25389,N_24502,N_24224);
and U25390 (N_25390,N_23548,N_23861);
nand U25391 (N_25391,N_23797,N_24243);
or U25392 (N_25392,N_24235,N_23690);
nor U25393 (N_25393,N_24481,N_24474);
nor U25394 (N_25394,N_23404,N_22502);
xnor U25395 (N_25395,N_24371,N_22520);
and U25396 (N_25396,N_24785,N_24557);
nand U25397 (N_25397,N_23004,N_23734);
nor U25398 (N_25398,N_24220,N_22515);
nor U25399 (N_25399,N_24796,N_24932);
nand U25400 (N_25400,N_24583,N_24594);
nor U25401 (N_25401,N_23295,N_22703);
or U25402 (N_25402,N_24058,N_24284);
nand U25403 (N_25403,N_22569,N_23063);
nor U25404 (N_25404,N_23057,N_22788);
xor U25405 (N_25405,N_23232,N_23931);
or U25406 (N_25406,N_23196,N_24661);
and U25407 (N_25407,N_24680,N_24155);
and U25408 (N_25408,N_22641,N_24165);
xnor U25409 (N_25409,N_23067,N_24201);
xnor U25410 (N_25410,N_24039,N_23934);
nand U25411 (N_25411,N_24758,N_24632);
or U25412 (N_25412,N_23675,N_24774);
nand U25413 (N_25413,N_23818,N_23174);
or U25414 (N_25414,N_23318,N_23578);
or U25415 (N_25415,N_24290,N_23025);
xnor U25416 (N_25416,N_23372,N_24117);
nand U25417 (N_25417,N_23337,N_23658);
nand U25418 (N_25418,N_22746,N_23634);
or U25419 (N_25419,N_22631,N_22982);
xor U25420 (N_25420,N_23618,N_23189);
or U25421 (N_25421,N_23960,N_24199);
nor U25422 (N_25422,N_23754,N_23803);
nand U25423 (N_25423,N_24797,N_24750);
xnor U25424 (N_25424,N_24576,N_24123);
or U25425 (N_25425,N_23090,N_24282);
and U25426 (N_25426,N_24084,N_24593);
and U25427 (N_25427,N_22816,N_24616);
xnor U25428 (N_25428,N_24352,N_22668);
nand U25429 (N_25429,N_24067,N_23240);
nand U25430 (N_25430,N_23361,N_22752);
and U25431 (N_25431,N_23774,N_24390);
or U25432 (N_25432,N_23941,N_23770);
xor U25433 (N_25433,N_24326,N_24223);
nor U25434 (N_25434,N_22843,N_23101);
nor U25435 (N_25435,N_23617,N_22888);
nand U25436 (N_25436,N_22718,N_22713);
nand U25437 (N_25437,N_23469,N_23416);
nand U25438 (N_25438,N_24723,N_24125);
nor U25439 (N_25439,N_24204,N_23338);
nand U25440 (N_25440,N_24871,N_24432);
or U25441 (N_25441,N_22671,N_22640);
nand U25442 (N_25442,N_23633,N_24802);
and U25443 (N_25443,N_24446,N_23447);
and U25444 (N_25444,N_24260,N_23426);
xor U25445 (N_25445,N_23939,N_23547);
nand U25446 (N_25446,N_23047,N_22827);
nand U25447 (N_25447,N_23133,N_24381);
xnor U25448 (N_25448,N_24578,N_22743);
or U25449 (N_25449,N_23482,N_23904);
or U25450 (N_25450,N_22760,N_22556);
and U25451 (N_25451,N_24400,N_24720);
and U25452 (N_25452,N_24244,N_24306);
nand U25453 (N_25453,N_23619,N_23243);
nor U25454 (N_25454,N_24636,N_23141);
nand U25455 (N_25455,N_23645,N_23497);
nor U25456 (N_25456,N_23711,N_23166);
nand U25457 (N_25457,N_23566,N_23406);
and U25458 (N_25458,N_24450,N_22954);
xnor U25459 (N_25459,N_24113,N_22667);
and U25460 (N_25460,N_23824,N_23739);
nand U25461 (N_25461,N_24392,N_24233);
or U25462 (N_25462,N_24748,N_24948);
nand U25463 (N_25463,N_22747,N_22621);
or U25464 (N_25464,N_23260,N_23514);
nor U25465 (N_25465,N_23073,N_22777);
nor U25466 (N_25466,N_24620,N_24542);
xnor U25467 (N_25467,N_22585,N_23527);
xnor U25468 (N_25468,N_24142,N_24990);
or U25469 (N_25469,N_24635,N_23985);
xor U25470 (N_25470,N_22651,N_23759);
and U25471 (N_25471,N_23822,N_22603);
or U25472 (N_25472,N_24791,N_24089);
xnor U25473 (N_25473,N_24138,N_22541);
nor U25474 (N_25474,N_23369,N_22897);
nand U25475 (N_25475,N_22853,N_23054);
or U25476 (N_25476,N_24648,N_24878);
or U25477 (N_25477,N_24286,N_23695);
nand U25478 (N_25478,N_24897,N_24903);
and U25479 (N_25479,N_24740,N_24256);
nand U25480 (N_25480,N_24413,N_23965);
nand U25481 (N_25481,N_23883,N_22614);
or U25482 (N_25482,N_24565,N_24874);
or U25483 (N_25483,N_23767,N_23412);
and U25484 (N_25484,N_24691,N_24096);
nand U25485 (N_25485,N_23359,N_23250);
or U25486 (N_25486,N_23363,N_22529);
xnor U25487 (N_25487,N_24085,N_24070);
nand U25488 (N_25488,N_24529,N_22823);
and U25489 (N_25489,N_24829,N_23586);
nor U25490 (N_25490,N_23184,N_24927);
or U25491 (N_25491,N_23594,N_23241);
nand U25492 (N_25492,N_24422,N_24879);
xor U25493 (N_25493,N_22684,N_24198);
xnor U25494 (N_25494,N_23383,N_23333);
xnor U25495 (N_25495,N_22835,N_23556);
or U25496 (N_25496,N_23159,N_23761);
nand U25497 (N_25497,N_22852,N_24499);
or U25498 (N_25498,N_23373,N_23078);
and U25499 (N_25499,N_23263,N_23192);
and U25500 (N_25500,N_23172,N_24536);
nor U25501 (N_25501,N_23538,N_24133);
nand U25502 (N_25502,N_23687,N_23328);
nor U25503 (N_25503,N_24535,N_23435);
xnor U25504 (N_25504,N_24185,N_24624);
nor U25505 (N_25505,N_24570,N_23018);
and U25506 (N_25506,N_24657,N_22751);
or U25507 (N_25507,N_22851,N_24073);
and U25508 (N_25508,N_22755,N_23450);
or U25509 (N_25509,N_23874,N_24882);
and U25510 (N_25510,N_23231,N_24528);
or U25511 (N_25511,N_24587,N_22978);
nand U25512 (N_25512,N_23242,N_24762);
or U25513 (N_25513,N_24053,N_22527);
xnor U25514 (N_25514,N_23335,N_24176);
nand U25515 (N_25515,N_23555,N_22791);
nor U25516 (N_25516,N_23178,N_24434);
and U25517 (N_25517,N_22725,N_22545);
xor U25518 (N_25518,N_22655,N_24615);
or U25519 (N_25519,N_24883,N_24561);
xor U25520 (N_25520,N_23091,N_24569);
nor U25521 (N_25521,N_23664,N_23563);
and U25522 (N_25522,N_23551,N_23826);
or U25523 (N_25523,N_23343,N_23458);
xnor U25524 (N_25524,N_23992,N_22721);
nand U25525 (N_25525,N_23998,N_22787);
and U25526 (N_25526,N_24395,N_23076);
or U25527 (N_25527,N_24809,N_22799);
nor U25528 (N_25528,N_23121,N_24380);
or U25529 (N_25529,N_23728,N_22822);
xnor U25530 (N_25530,N_23151,N_23532);
or U25531 (N_25531,N_23930,N_22850);
or U25532 (N_25532,N_23714,N_24497);
and U25533 (N_25533,N_24066,N_24469);
xor U25534 (N_25534,N_22576,N_22773);
or U25535 (N_25535,N_22883,N_24077);
or U25536 (N_25536,N_23323,N_24821);
nand U25537 (N_25537,N_22768,N_22643);
or U25538 (N_25538,N_22553,N_24462);
nor U25539 (N_25539,N_23261,N_22918);
and U25540 (N_25540,N_23518,N_24189);
xnor U25541 (N_25541,N_23651,N_24247);
xnor U25542 (N_25542,N_23491,N_22936);
xnor U25543 (N_25543,N_23536,N_24994);
or U25544 (N_25544,N_24270,N_22957);
and U25545 (N_25545,N_24079,N_23911);
xor U25546 (N_25546,N_22592,N_24793);
nand U25547 (N_25547,N_24498,N_22726);
or U25548 (N_25548,N_24858,N_23820);
and U25549 (N_25549,N_22648,N_23218);
and U25550 (N_25550,N_23740,N_23308);
and U25551 (N_25551,N_24182,N_23953);
and U25552 (N_25552,N_23440,N_22586);
or U25553 (N_25553,N_24876,N_24959);
xnor U25554 (N_25554,N_23962,N_24922);
or U25555 (N_25555,N_24018,N_22730);
and U25556 (N_25556,N_23755,N_23521);
and U25557 (N_25557,N_24172,N_22988);
nand U25558 (N_25558,N_23344,N_23388);
nand U25559 (N_25559,N_23747,N_24823);
nor U25560 (N_25560,N_23700,N_23300);
or U25561 (N_25561,N_24393,N_23284);
xor U25562 (N_25562,N_24183,N_22861);
nand U25563 (N_25563,N_24437,N_22948);
and U25564 (N_25564,N_24323,N_22654);
xnor U25565 (N_25565,N_23006,N_22862);
nor U25566 (N_25566,N_24890,N_23212);
nor U25567 (N_25567,N_23315,N_24515);
or U25568 (N_25568,N_24603,N_24329);
and U25569 (N_25569,N_24512,N_22949);
xnor U25570 (N_25570,N_23813,N_24068);
nand U25571 (N_25571,N_22583,N_23783);
nor U25572 (N_25572,N_23997,N_23994);
nor U25573 (N_25573,N_24403,N_23964);
or U25574 (N_25574,N_23082,N_24324);
xnor U25575 (N_25575,N_24404,N_23452);
nor U25576 (N_25576,N_24406,N_24001);
xnor U25577 (N_25577,N_23375,N_22500);
or U25578 (N_25578,N_24401,N_23801);
xor U25579 (N_25579,N_23443,N_23671);
nand U25580 (N_25580,N_22983,N_22875);
xor U25581 (N_25581,N_23623,N_23535);
and U25582 (N_25582,N_23611,N_24891);
and U25583 (N_25583,N_23961,N_23925);
and U25584 (N_25584,N_22728,N_22537);
or U25585 (N_25585,N_24608,N_23048);
nand U25586 (N_25586,N_24905,N_24009);
nor U25587 (N_25587,N_23550,N_22692);
or U25588 (N_25588,N_23357,N_24215);
xnor U25589 (N_25589,N_22540,N_24151);
nor U25590 (N_25590,N_23575,N_23627);
xnor U25591 (N_25591,N_24853,N_23855);
nand U25592 (N_25592,N_23259,N_24804);
xnor U25593 (N_25593,N_23508,N_24081);
nand U25594 (N_25594,N_24048,N_23540);
nand U25595 (N_25595,N_24962,N_24026);
nor U25596 (N_25596,N_24965,N_22589);
or U25597 (N_25597,N_24782,N_22842);
xor U25598 (N_25598,N_23884,N_23339);
nand U25599 (N_25599,N_24953,N_22704);
or U25600 (N_25600,N_23745,N_23727);
nor U25601 (N_25601,N_22745,N_22632);
or U25602 (N_25602,N_23124,N_22995);
nand U25603 (N_25603,N_23620,N_24251);
and U25604 (N_25604,N_24655,N_24466);
nand U25605 (N_25605,N_24391,N_24063);
xnor U25606 (N_25606,N_24815,N_22564);
nand U25607 (N_25607,N_24006,N_22705);
or U25608 (N_25608,N_24609,N_23721);
xnor U25609 (N_25609,N_23081,N_23976);
nand U25610 (N_25610,N_23396,N_24637);
or U25611 (N_25611,N_22782,N_23341);
nand U25612 (N_25612,N_24069,N_22627);
xor U25613 (N_25613,N_23983,N_22588);
and U25614 (N_25614,N_23996,N_24501);
nand U25615 (N_25615,N_23903,N_22754);
xor U25616 (N_25616,N_22865,N_23271);
xor U25617 (N_25617,N_24414,N_22968);
nand U25618 (N_25618,N_23870,N_24568);
or U25619 (N_25619,N_23599,N_24560);
or U25620 (N_25620,N_23219,N_23604);
or U25621 (N_25621,N_24276,N_23816);
or U25622 (N_25622,N_24424,N_24808);
nand U25623 (N_25623,N_23696,N_24760);
nor U25624 (N_25624,N_24087,N_22659);
xnor U25625 (N_25625,N_23595,N_22536);
or U25626 (N_25626,N_24104,N_23973);
and U25627 (N_25627,N_22572,N_24945);
nor U25628 (N_25628,N_24538,N_23589);
nand U25629 (N_25629,N_23609,N_24208);
nor U25630 (N_25630,N_22567,N_24298);
nand U25631 (N_25631,N_24745,N_22929);
nand U25632 (N_25632,N_23417,N_22924);
nor U25633 (N_25633,N_24289,N_23122);
and U25634 (N_25634,N_24803,N_24460);
nand U25635 (N_25635,N_22780,N_24789);
xor U25636 (N_25636,N_22575,N_22639);
xnor U25637 (N_25637,N_23522,N_24541);
and U25638 (N_25638,N_22584,N_23157);
or U25639 (N_25639,N_23024,N_23423);
and U25640 (N_25640,N_23351,N_23878);
and U25641 (N_25641,N_22866,N_23393);
and U25642 (N_25642,N_24255,N_23863);
or U25643 (N_25643,N_23790,N_24881);
and U25644 (N_25644,N_22798,N_24597);
and U25645 (N_25645,N_24766,N_23554);
nor U25646 (N_25646,N_23716,N_23908);
nand U25647 (N_25647,N_23299,N_23349);
nor U25648 (N_25648,N_24696,N_23652);
and U25649 (N_25649,N_23726,N_22989);
xor U25650 (N_25650,N_23126,N_24203);
or U25651 (N_25651,N_23529,N_22966);
xor U25652 (N_25652,N_23471,N_23083);
and U25653 (N_25653,N_22679,N_23558);
or U25654 (N_25654,N_23399,N_24226);
or U25655 (N_25655,N_24488,N_22604);
nand U25656 (N_25656,N_23001,N_24519);
xor U25657 (N_25657,N_23100,N_23108);
nor U25658 (N_25658,N_24689,N_24457);
nand U25659 (N_25659,N_24046,N_24107);
nand U25660 (N_25660,N_22682,N_24520);
and U25661 (N_25661,N_24225,N_24402);
nor U25662 (N_25662,N_23736,N_24783);
nand U25663 (N_25663,N_23565,N_24484);
or U25664 (N_25664,N_24301,N_24345);
and U25665 (N_25665,N_23457,N_23325);
xnor U25666 (N_25666,N_23749,N_23590);
and U25667 (N_25667,N_24014,N_24562);
or U25668 (N_25668,N_23272,N_24634);
nand U25669 (N_25669,N_24754,N_23033);
nor U25670 (N_25670,N_23958,N_24316);
and U25671 (N_25671,N_24139,N_24559);
and U25672 (N_25672,N_24478,N_24998);
nand U25673 (N_25673,N_23744,N_23499);
xor U25674 (N_25674,N_23223,N_22890);
or U25675 (N_25675,N_24145,N_24149);
and U25676 (N_25676,N_24480,N_22979);
xnor U25677 (N_25677,N_22786,N_22926);
and U25678 (N_25678,N_23640,N_24489);
or U25679 (N_25679,N_24412,N_24638);
or U25680 (N_25680,N_24336,N_23825);
nor U25681 (N_25681,N_24817,N_24606);
nand U25682 (N_25682,N_23559,N_23630);
or U25683 (N_25683,N_23445,N_23612);
nor U25684 (N_25684,N_24150,N_24088);
nor U25685 (N_25685,N_23470,N_23382);
xnor U25686 (N_25686,N_24588,N_24589);
and U25687 (N_25687,N_23592,N_23760);
nor U25688 (N_25688,N_24957,N_22741);
and U25689 (N_25689,N_24340,N_22810);
and U25690 (N_25690,N_24996,N_23907);
or U25691 (N_25691,N_22552,N_23167);
xnor U25692 (N_25692,N_23756,N_23636);
nor U25693 (N_25693,N_23253,N_24801);
or U25694 (N_25694,N_24299,N_24574);
or U25695 (N_25695,N_24686,N_23210);
or U25696 (N_25696,N_23281,N_24969);
nand U25697 (N_25697,N_23400,N_24677);
or U25698 (N_25698,N_24045,N_22702);
nand U25699 (N_25699,N_23580,N_24611);
nor U25700 (N_25700,N_22938,N_23342);
or U25701 (N_25701,N_22887,N_23588);
nand U25702 (N_25702,N_24972,N_23753);
xor U25703 (N_25703,N_22919,N_23173);
nand U25704 (N_25704,N_22503,N_23429);
nand U25705 (N_25705,N_22560,N_22834);
nand U25706 (N_25706,N_24924,N_24949);
xor U25707 (N_25707,N_23511,N_23379);
and U25708 (N_25708,N_24420,N_23005);
or U25709 (N_25709,N_23202,N_24374);
nor U25710 (N_25710,N_23132,N_24701);
and U25711 (N_25711,N_24360,N_24075);
and U25712 (N_25712,N_23653,N_23413);
nand U25713 (N_25713,N_22784,N_22764);
and U25714 (N_25714,N_23370,N_23276);
and U25715 (N_25715,N_23752,N_24644);
and U25716 (N_25716,N_23940,N_22696);
and U25717 (N_25717,N_23732,N_23926);
nand U25718 (N_25718,N_24951,N_22997);
nand U25719 (N_25719,N_22761,N_24093);
nand U25720 (N_25720,N_24631,N_24968);
nand U25721 (N_25721,N_23517,N_23674);
nor U25722 (N_25722,N_23495,N_24297);
xor U25723 (N_25723,N_22881,N_22937);
and U25724 (N_25724,N_22625,N_24368);
and U25725 (N_25725,N_23391,N_23163);
nor U25726 (N_25726,N_23798,N_22594);
nor U25727 (N_25727,N_23900,N_24156);
nand U25728 (N_25728,N_23340,N_24580);
xnor U25729 (N_25729,N_24396,N_24544);
xnor U25730 (N_25730,N_24454,N_24572);
or U25731 (N_25731,N_24849,N_23549);
xnor U25732 (N_25732,N_23298,N_24076);
or U25733 (N_25733,N_22973,N_23089);
and U25734 (N_25734,N_23616,N_23366);
and U25735 (N_25735,N_23454,N_22644);
nor U25736 (N_25736,N_23849,N_23422);
nand U25737 (N_25737,N_22763,N_23625);
nor U25738 (N_25738,N_22794,N_23978);
nor U25739 (N_25739,N_24925,N_22870);
nand U25740 (N_25740,N_23719,N_24510);
nor U25741 (N_25741,N_22698,N_24438);
xnor U25742 (N_25742,N_24258,N_22999);
nor U25743 (N_25743,N_23923,N_23221);
or U25744 (N_25744,N_24452,N_24373);
and U25745 (N_25745,N_24281,N_24312);
or U25746 (N_25746,N_24050,N_23201);
and U25747 (N_25747,N_24057,N_24697);
nor U25748 (N_25748,N_24999,N_23804);
nor U25749 (N_25749,N_22600,N_24841);
nand U25750 (N_25750,N_23762,N_22736);
or U25751 (N_25751,N_24896,N_24863);
or U25752 (N_25752,N_24698,N_24091);
and U25753 (N_25753,N_23642,N_22717);
and U25754 (N_25754,N_24518,N_23927);
nor U25755 (N_25755,N_22844,N_24685);
nor U25756 (N_25756,N_24442,N_23679);
or U25757 (N_25757,N_23929,N_24034);
and U25758 (N_25758,N_23614,N_23970);
and U25759 (N_25759,N_24800,N_22889);
or U25760 (N_25760,N_23345,N_22872);
nor U25761 (N_25761,N_22942,N_23915);
or U25762 (N_25762,N_23873,N_23821);
nand U25763 (N_25763,N_23893,N_24755);
or U25764 (N_25764,N_22893,N_24461);
or U25765 (N_25765,N_23621,N_23053);
nand U25766 (N_25766,N_24229,N_24928);
xnor U25767 (N_25767,N_23730,N_24625);
and U25768 (N_25768,N_23424,N_22765);
or U25769 (N_25769,N_24399,N_23307);
and U25770 (N_25770,N_23498,N_24681);
and U25771 (N_25771,N_24772,N_23905);
or U25772 (N_25772,N_22506,N_23322);
nor U25773 (N_25773,N_23561,N_23070);
and U25774 (N_25774,N_23220,N_22753);
xnor U25775 (N_25775,N_23624,N_23657);
and U25776 (N_25776,N_23386,N_22699);
nand U25777 (N_25777,N_24507,N_23038);
xor U25778 (N_25778,N_24875,N_23028);
or U25779 (N_25779,N_23316,N_22689);
nand U25780 (N_25780,N_23988,N_22638);
nor U25781 (N_25781,N_23572,N_24548);
or U25782 (N_25782,N_24020,N_23909);
nand U25783 (N_25783,N_23897,N_24135);
and U25784 (N_25784,N_22902,N_23488);
nand U25785 (N_25785,N_23769,N_23436);
nor U25786 (N_25786,N_23287,N_23513);
nand U25787 (N_25787,N_23865,N_23071);
nand U25788 (N_25788,N_23431,N_24721);
nand U25789 (N_25789,N_23771,N_23102);
xnor U25790 (N_25790,N_22833,N_23378);
nand U25791 (N_25791,N_23035,N_24032);
and U25792 (N_25792,N_23735,N_23285);
nand U25793 (N_25793,N_24471,N_24458);
nor U25794 (N_25794,N_24269,N_24747);
or U25795 (N_25795,N_24929,N_23467);
nor U25796 (N_25796,N_23507,N_23766);
nor U25797 (N_25797,N_24671,N_24584);
or U25798 (N_25798,N_24861,N_22863);
nor U25799 (N_25799,N_22504,N_23792);
nor U25800 (N_25800,N_23198,N_23410);
nor U25801 (N_25801,N_22544,N_23374);
nor U25802 (N_25802,N_22896,N_23127);
or U25803 (N_25803,N_23044,N_22512);
and U25804 (N_25804,N_22963,N_24174);
and U25805 (N_25805,N_24309,N_24288);
or U25806 (N_25806,N_23043,N_23051);
and U25807 (N_25807,N_23693,N_22535);
xor U25808 (N_25808,N_22677,N_24383);
or U25809 (N_25809,N_23981,N_23248);
nor U25810 (N_25810,N_22907,N_22674);
or U25811 (N_25811,N_23061,N_22642);
xnor U25812 (N_25812,N_23859,N_24771);
and U25813 (N_25813,N_23093,N_23390);
and U25814 (N_25814,N_23779,N_24292);
and U25815 (N_25815,N_23360,N_24746);
xnor U25816 (N_25816,N_24765,N_22952);
and U25817 (N_25817,N_24735,N_22735);
nand U25818 (N_25818,N_23773,N_24901);
nor U25819 (N_25819,N_24966,N_24852);
nand U25820 (N_25820,N_23534,N_23706);
nor U25821 (N_25821,N_23584,N_22809);
and U25822 (N_25822,N_24363,N_24019);
and U25823 (N_25823,N_22960,N_23019);
and U25824 (N_25824,N_22781,N_23602);
xor U25825 (N_25825,N_23441,N_24016);
xnor U25826 (N_25826,N_24418,N_24367);
xor U25827 (N_25827,N_24405,N_24083);
nor U25828 (N_25828,N_22792,N_22716);
xnor U25829 (N_25829,N_23139,N_23503);
or U25830 (N_25830,N_24537,N_23977);
and U25831 (N_25831,N_23087,N_22837);
nor U25832 (N_25832,N_24683,N_24788);
nor U25833 (N_25833,N_24232,N_24546);
and U25834 (N_25834,N_24604,N_24982);
or U25835 (N_25835,N_23135,N_24757);
nand U25836 (N_25836,N_24435,N_23303);
or U25837 (N_25837,N_23099,N_24684);
xnor U25838 (N_25838,N_22885,N_24690);
nor U25839 (N_25839,N_23948,N_23113);
and U25840 (N_25840,N_23831,N_23827);
xnor U25841 (N_25841,N_24688,N_23782);
nor U25842 (N_25842,N_24795,N_23605);
nor U25843 (N_25843,N_24237,N_24556);
and U25844 (N_25844,N_23570,N_24207);
or U25845 (N_25845,N_22534,N_24595);
nor U25846 (N_25846,N_23887,N_24665);
nand U25847 (N_25847,N_22971,N_24761);
or U25848 (N_25848,N_22796,N_22859);
nand U25849 (N_25849,N_24779,N_24495);
xnor U25850 (N_25850,N_24476,N_22917);
or U25851 (N_25851,N_23596,N_23567);
nor U25852 (N_25852,N_24372,N_24127);
nor U25853 (N_25853,N_23291,N_22912);
or U25854 (N_25854,N_24408,N_24773);
nand U25855 (N_25855,N_22593,N_24295);
nor U25856 (N_25856,N_24963,N_23233);
and U25857 (N_25857,N_24384,N_22839);
nand U25858 (N_25858,N_23306,N_23724);
and U25859 (N_25859,N_24577,N_23933);
nor U25860 (N_25860,N_23764,N_23069);
and U25861 (N_25861,N_24042,N_23834);
xor U25862 (N_25862,N_23738,N_23795);
nand U25863 (N_25863,N_23502,N_23743);
xor U25864 (N_25864,N_23817,N_23017);
xnor U25865 (N_25865,N_23950,N_24015);
or U25866 (N_25866,N_22860,N_23670);
and U25867 (N_25867,N_23701,N_22518);
or U25868 (N_25868,N_22656,N_23898);
xnor U25869 (N_25869,N_24997,N_24191);
and U25870 (N_25870,N_24700,N_23954);
or U25871 (N_25871,N_22845,N_24913);
xor U25872 (N_25872,N_23302,N_22616);
or U25873 (N_25873,N_22884,N_23222);
nor U25874 (N_25874,N_24564,N_23000);
xor U25875 (N_25875,N_23519,N_23009);
nand U25876 (N_25876,N_24353,N_23603);
nor U25877 (N_25877,N_23691,N_24667);
and U25878 (N_25878,N_23209,N_23788);
or U25879 (N_25879,N_24337,N_24049);
nor U25880 (N_25880,N_24028,N_23707);
xnor U25881 (N_25881,N_24061,N_23920);
nand U25882 (N_25882,N_23118,N_23449);
nand U25883 (N_25883,N_22991,N_24500);
and U25884 (N_25884,N_24549,N_23265);
and U25885 (N_25885,N_23411,N_24832);
and U25886 (N_25886,N_23191,N_24097);
or U25887 (N_25887,N_22687,N_24193);
nand U25888 (N_25888,N_23205,N_23639);
xnor U25889 (N_25889,N_24388,N_22708);
nand U25890 (N_25890,N_22617,N_23251);
or U25891 (N_25891,N_24121,N_24991);
and U25892 (N_25892,N_24845,N_24980);
xnor U25893 (N_25893,N_24707,N_22516);
or U25894 (N_25894,N_23668,N_24386);
nor U25895 (N_25895,N_24805,N_22925);
and U25896 (N_25896,N_23881,N_23270);
xor U25897 (N_25897,N_23833,N_22508);
and U25898 (N_25898,N_23348,N_23255);
and U25899 (N_25899,N_22769,N_23314);
nor U25900 (N_25900,N_24820,N_22599);
nand U25901 (N_25901,N_24245,N_22665);
nor U25902 (N_25902,N_24071,N_22555);
xnor U25903 (N_25903,N_23949,N_22737);
xnor U25904 (N_25904,N_23246,N_23857);
nand U25905 (N_25905,N_24037,N_24152);
nor U25906 (N_25906,N_22869,N_23703);
and U25907 (N_25907,N_22914,N_24465);
xnor U25908 (N_25908,N_24767,N_22548);
nand U25909 (N_25909,N_24496,N_24887);
nand U25910 (N_25910,N_24332,N_22562);
xnor U25911 (N_25911,N_22854,N_23014);
nand U25912 (N_25912,N_23021,N_22906);
or U25913 (N_25913,N_24341,N_24490);
and U25914 (N_25914,N_22577,N_22967);
and U25915 (N_25915,N_23226,N_23283);
nand U25916 (N_25916,N_22542,N_24327);
or U25917 (N_25917,N_24423,N_22706);
or U25918 (N_25918,N_24647,N_22880);
or U25919 (N_25919,N_23026,N_24486);
xor U25920 (N_25920,N_23165,N_23980);
and U25921 (N_25921,N_22814,N_23475);
and U25922 (N_25922,N_22915,N_24065);
or U25923 (N_25923,N_22927,N_24448);
nand U25924 (N_25924,N_23713,N_24873);
nand U25925 (N_25925,N_24623,N_22732);
or U25926 (N_25926,N_22505,N_24025);
nand U25927 (N_25927,N_24825,N_23027);
nor U25928 (N_25928,N_23142,N_23479);
xor U25929 (N_25929,N_23598,N_23313);
xnor U25930 (N_25930,N_23474,N_23650);
or U25931 (N_25931,N_23867,N_24836);
nand U25932 (N_25932,N_22813,N_22622);
nand U25933 (N_25933,N_22994,N_22710);
xor U25934 (N_25934,N_23694,N_22775);
nand U25935 (N_25935,N_23451,N_23408);
nand U25936 (N_25936,N_23199,N_22691);
and U25937 (N_25937,N_24936,N_24627);
xnor U25938 (N_25938,N_23418,N_23689);
nand U25939 (N_25939,N_24164,N_24598);
nor U25940 (N_25940,N_24056,N_23712);
nand U25941 (N_25941,N_24961,N_22733);
xnor U25942 (N_25942,N_24439,N_24227);
nor U25943 (N_25943,N_24387,N_23600);
xnor U25944 (N_25944,N_24180,N_22646);
nor U25945 (N_25945,N_23472,N_24307);
nor U25946 (N_25946,N_24007,N_24699);
or U25947 (N_25947,N_23500,N_22657);
or U25948 (N_25948,N_24839,N_23562);
and U25949 (N_25949,N_24669,N_22590);
nand U25950 (N_25950,N_22597,N_24159);
and U25951 (N_25951,N_24494,N_23557);
nand U25952 (N_25952,N_24357,N_23876);
and U25953 (N_25953,N_23480,N_22871);
or U25954 (N_25954,N_23112,N_23465);
or U25955 (N_25955,N_24906,N_23023);
and U25956 (N_25956,N_22959,N_22877);
nor U25957 (N_25957,N_24884,N_22601);
xnor U25958 (N_25958,N_24263,N_23647);
or U25959 (N_25959,N_24907,N_24834);
or U25960 (N_25960,N_23659,N_24926);
nor U25961 (N_25961,N_22722,N_24342);
nor U25962 (N_25962,N_22664,N_22817);
or U25963 (N_25963,N_22563,N_24300);
xor U25964 (N_25964,N_24062,N_23737);
nor U25965 (N_25965,N_22762,N_24621);
or U25966 (N_25966,N_23913,N_24248);
and U25967 (N_25967,N_24455,N_24344);
xor U25968 (N_25968,N_24670,N_23176);
nor U25969 (N_25969,N_22996,N_22658);
or U25970 (N_25970,N_23438,N_24786);
or U25971 (N_25971,N_24167,N_23280);
and U25972 (N_25972,N_23181,N_23128);
or U25973 (N_25973,N_23676,N_23262);
nor U25974 (N_25974,N_23963,N_24430);
nor U25975 (N_25975,N_22719,N_23520);
or U25976 (N_25976,N_24682,N_23539);
nor U25977 (N_25977,N_22920,N_22626);
nor U25978 (N_25978,N_23180,N_23394);
and U25979 (N_25979,N_23974,N_24526);
and U25980 (N_25980,N_24319,N_24240);
or U25981 (N_25981,N_24356,N_22900);
xnor U25982 (N_25982,N_22766,N_22661);
nor U25983 (N_25983,N_24140,N_23789);
or U25984 (N_25984,N_24377,N_24415);
xor U25985 (N_25985,N_22519,N_24952);
nand U25986 (N_25986,N_23839,N_23056);
nor U25987 (N_25987,N_24586,N_22767);
nor U25988 (N_25988,N_23114,N_23666);
and U25989 (N_25989,N_24885,N_23187);
xor U25990 (N_25990,N_24419,N_23505);
nand U25991 (N_25991,N_23179,N_23347);
or U25992 (N_25992,N_24916,N_24192);
nor U25993 (N_25993,N_23793,N_24525);
nor U25994 (N_25994,N_24177,N_24378);
or U25995 (N_25995,N_22882,N_23628);
xnor U25996 (N_25996,N_24566,N_24141);
nand U25997 (N_25997,N_24394,N_24362);
and U25998 (N_25998,N_24249,N_24893);
nor U25999 (N_25999,N_24099,N_22628);
nor U26000 (N_26000,N_24643,N_23489);
and U26001 (N_26001,N_23723,N_24694);
nand U26002 (N_26002,N_23722,N_23031);
nand U26003 (N_26003,N_24120,N_23680);
and U26004 (N_26004,N_24197,N_22964);
and U26005 (N_26005,N_23785,N_24012);
nand U26006 (N_26006,N_24710,N_24033);
nand U26007 (N_26007,N_23249,N_23802);
nor U26008 (N_26008,N_23968,N_23235);
xor U26009 (N_26009,N_23059,N_22558);
nand U26010 (N_26010,N_24366,N_23312);
and U26011 (N_26011,N_23346,N_24047);
nand U26012 (N_26012,N_24343,N_23819);
or U26013 (N_26013,N_24819,N_24334);
nand U26014 (N_26014,N_23667,N_24687);
nand U26015 (N_26015,N_24539,N_24124);
or U26016 (N_26016,N_24268,N_22729);
nor U26017 (N_26017,N_24533,N_23742);
or U26018 (N_26018,N_24517,N_23593);
and U26019 (N_26019,N_24563,N_22886);
nand U26020 (N_26020,N_22828,N_23238);
nand U26021 (N_26021,N_23569,N_23286);
nand U26022 (N_26022,N_24872,N_23490);
or U26023 (N_26023,N_24726,N_24147);
and U26024 (N_26024,N_22785,N_22931);
xor U26025 (N_26025,N_24132,N_23247);
xor U26026 (N_26026,N_22857,N_24449);
nand U26027 (N_26027,N_24888,N_23895);
nand U26028 (N_26028,N_23972,N_22723);
xnor U26029 (N_26029,N_24272,N_24444);
nor U26030 (N_26030,N_23190,N_22779);
or U26031 (N_26031,N_22820,N_24919);
xor U26032 (N_26032,N_23110,N_22524);
xnor U26033 (N_26033,N_22738,N_24763);
and U26034 (N_26034,N_24792,N_23320);
nand U26035 (N_26035,N_23872,N_23008);
xnor U26036 (N_26036,N_24119,N_24869);
and U26037 (N_26037,N_24787,N_22821);
nand U26038 (N_26038,N_24846,N_24727);
xor U26039 (N_26039,N_23208,N_22669);
or U26040 (N_26040,N_22528,N_24652);
and U26041 (N_26041,N_22981,N_23573);
or U26042 (N_26042,N_23088,N_24196);
nor U26043 (N_26043,N_23850,N_24602);
or U26044 (N_26044,N_23969,N_23213);
nor U26045 (N_26045,N_23677,N_23264);
nor U26046 (N_26046,N_24017,N_23045);
xnor U26047 (N_26047,N_23626,N_23158);
or U26048 (N_26048,N_23606,N_23384);
xor U26049 (N_26049,N_23050,N_24729);
nand U26050 (N_26050,N_24315,N_24995);
or U26051 (N_26051,N_24238,N_23984);
or U26052 (N_26052,N_23380,N_22701);
nand U26053 (N_26053,N_22836,N_23206);
and U26054 (N_26054,N_24831,N_23156);
nand U26055 (N_26055,N_24102,N_23137);
xnor U26056 (N_26056,N_24868,N_22554);
and U26057 (N_26057,N_23646,N_22673);
or U26058 (N_26058,N_24798,N_24613);
and U26059 (N_26059,N_24806,N_24950);
and U26060 (N_26060,N_22647,N_24551);
or U26061 (N_26061,N_23546,N_24482);
xnor U26062 (N_26062,N_22848,N_24830);
nor U26063 (N_26063,N_24485,N_23446);
and U26064 (N_26064,N_23919,N_23183);
nor U26065 (N_26065,N_24186,N_22980);
nor U26066 (N_26066,N_24002,N_24844);
and U26067 (N_26067,N_24144,N_24769);
xnor U26068 (N_26068,N_23772,N_24162);
nor U26069 (N_26069,N_23215,N_23077);
and U26070 (N_26070,N_24937,N_23104);
or U26071 (N_26071,N_24988,N_23890);
xnor U26072 (N_26072,N_22742,N_23419);
nand U26073 (N_26073,N_22618,N_24810);
xnor U26074 (N_26074,N_23564,N_22568);
nand U26075 (N_26075,N_22634,N_24575);
nand U26076 (N_26076,N_24130,N_23995);
xor U26077 (N_26077,N_23289,N_24389);
or U26078 (N_26078,N_22847,N_24333);
xnor U26079 (N_26079,N_23989,N_24984);
nand U26080 (N_26080,N_24108,N_23129);
or U26081 (N_26081,N_24348,N_23848);
xor U26082 (N_26082,N_24267,N_22830);
or U26083 (N_26083,N_24731,N_24812);
nand U26084 (N_26084,N_23094,N_24590);
nand U26085 (N_26085,N_22672,N_23661);
nor U26086 (N_26086,N_23064,N_22514);
xor U26087 (N_26087,N_24064,N_23244);
and U26088 (N_26088,N_24022,N_23852);
xnor U26089 (N_26089,N_23013,N_22693);
and U26090 (N_26090,N_22811,N_24781);
or U26091 (N_26091,N_23869,N_23125);
nand U26092 (N_26092,N_23758,N_23011);
nor U26093 (N_26093,N_23896,N_24187);
nor U26094 (N_26094,N_22650,N_23402);
and U26095 (N_26095,N_22783,N_23637);
and U26096 (N_26096,N_22697,N_22934);
nor U26097 (N_26097,N_24506,N_24361);
nand U26098 (N_26098,N_23367,N_22645);
nand U26099 (N_26099,N_23040,N_23875);
nand U26100 (N_26100,N_24554,N_22714);
and U26101 (N_26101,N_23851,N_24364);
and U26102 (N_26102,N_24283,N_23055);
nand U26103 (N_26103,N_24744,N_23815);
and U26104 (N_26104,N_24838,N_23415);
xor U26105 (N_26105,N_24857,N_22795);
and U26106 (N_26106,N_22595,N_24599);
and U26107 (N_26107,N_24451,N_24234);
xor U26108 (N_26108,N_24285,N_22531);
and U26109 (N_26109,N_24617,N_24894);
xor U26110 (N_26110,N_22695,N_23644);
and U26111 (N_26111,N_22935,N_24021);
nand U26112 (N_26112,N_24254,N_24060);
or U26113 (N_26113,N_24530,N_23461);
nor U26114 (N_26114,N_24103,N_23956);
and U26115 (N_26115,N_23052,N_22829);
xor U26116 (N_26116,N_24112,N_24166);
and U26117 (N_26117,N_23123,N_24610);
nor U26118 (N_26118,N_22757,N_24889);
nor U26119 (N_26119,N_22602,N_23092);
and U26120 (N_26120,N_24645,N_23523);
or U26121 (N_26121,N_23496,N_23468);
nand U26122 (N_26122,N_23704,N_23039);
or U26123 (N_26123,N_22629,N_23545);
and U26124 (N_26124,N_24626,N_24246);
nand U26125 (N_26125,N_22891,N_23971);
nand U26126 (N_26126,N_22831,N_22802);
or U26127 (N_26127,N_24098,N_23866);
nand U26128 (N_26128,N_23321,N_24534);
nor U26129 (N_26129,N_24856,N_23681);
nor U26130 (N_26130,N_23478,N_23117);
and U26131 (N_26131,N_22579,N_24350);
xor U26132 (N_26132,N_24816,N_24659);
or U26133 (N_26133,N_24547,N_24349);
xor U26134 (N_26134,N_24867,N_23662);
and U26135 (N_26135,N_24475,N_22977);
and U26136 (N_26136,N_22928,N_23922);
nand U26137 (N_26137,N_24425,N_24592);
or U26138 (N_26138,N_24265,N_24184);
xnor U26139 (N_26139,N_22930,N_23273);
nand U26140 (N_26140,N_24650,N_24612);
nand U26141 (N_26141,N_24706,N_24236);
xnor U26142 (N_26142,N_23075,N_24115);
nor U26143 (N_26143,N_23786,N_23889);
nor U26144 (N_26144,N_24666,N_24264);
or U26145 (N_26145,N_24521,N_24674);
and U26146 (N_26146,N_23317,N_22581);
nor U26147 (N_26147,N_22984,N_22715);
or U26148 (N_26148,N_23109,N_24209);
and U26149 (N_26149,N_23477,N_23708);
xnor U26150 (N_26150,N_24734,N_23330);
nand U26151 (N_26151,N_24148,N_22547);
nand U26152 (N_26152,N_22923,N_22598);
nor U26153 (N_26153,N_23149,N_24031);
xnor U26154 (N_26154,N_22623,N_24934);
and U26155 (N_26155,N_23012,N_23326);
and U26156 (N_26156,N_24171,N_23957);
or U26157 (N_26157,N_24508,N_22789);
nand U26158 (N_26158,N_23660,N_22825);
nand U26159 (N_26159,N_22895,N_24918);
or U26160 (N_26160,N_24640,N_23267);
nor U26161 (N_26161,N_24775,N_23476);
or U26162 (N_26162,N_23297,N_24679);
nor U26163 (N_26163,N_23705,N_24304);
or U26164 (N_26164,N_24086,N_23010);
and U26165 (N_26165,N_24092,N_23835);
xnor U26166 (N_26166,N_23775,N_23581);
or U26167 (N_26167,N_22749,N_24714);
and U26168 (N_26168,N_23515,N_24938);
and U26169 (N_26169,N_23397,N_22922);
or U26170 (N_26170,N_23891,N_23882);
nand U26171 (N_26171,N_24600,N_22609);
nand U26172 (N_26172,N_24464,N_24074);
nor U26173 (N_26173,N_24702,N_24228);
nor U26174 (N_26174,N_22571,N_24188);
or U26175 (N_26175,N_24328,N_23512);
nor U26176 (N_26176,N_24941,N_23029);
or U26177 (N_26177,N_24023,N_22951);
nor U26178 (N_26178,N_23631,N_24935);
xnor U26179 (N_26179,N_22932,N_23296);
and U26180 (N_26180,N_23234,N_23959);
and U26181 (N_26181,N_22582,N_23425);
nand U26182 (N_26182,N_24252,N_24163);
nor U26183 (N_26183,N_24213,N_22711);
xor U26184 (N_26184,N_24646,N_24848);
and U26185 (N_26185,N_23062,N_23058);
and U26186 (N_26186,N_23568,N_23204);
xnor U26187 (N_26187,N_23466,N_24100);
nand U26188 (N_26188,N_24294,N_24908);
nor U26189 (N_26189,N_23120,N_22916);
or U26190 (N_26190,N_22551,N_22944);
nor U26191 (N_26191,N_23290,N_24824);
xor U26192 (N_26192,N_24170,N_24628);
and U26193 (N_26193,N_23279,N_24558);
xor U26194 (N_26194,N_24128,N_24004);
nor U26195 (N_26195,N_24877,N_23405);
xor U26196 (N_26196,N_24428,N_23162);
or U26197 (N_26197,N_23072,N_23177);
xnor U26198 (N_26198,N_23168,N_24231);
and U26199 (N_26199,N_24828,N_22910);
nor U26200 (N_26200,N_24943,N_24376);
nand U26201 (N_26201,N_24898,N_23193);
or U26202 (N_26202,N_23885,N_24483);
xor U26203 (N_26203,N_23607,N_23946);
xnor U26204 (N_26204,N_23987,N_23741);
nand U26205 (N_26205,N_23655,N_23709);
nand U26206 (N_26206,N_23252,N_24178);
and U26207 (N_26207,N_24855,N_24308);
nand U26208 (N_26208,N_24842,N_24013);
nor U26209 (N_26209,N_22574,N_23577);
and U26210 (N_26210,N_24555,N_24318);
nor U26211 (N_26211,N_23352,N_24899);
nand U26212 (N_26212,N_24780,N_23702);
xnor U26213 (N_26213,N_24764,N_22724);
or U26214 (N_26214,N_22663,N_23533);
nor U26215 (N_26215,N_23079,N_23481);
xnor U26216 (N_26216,N_24784,N_22970);
nor U26217 (N_26217,N_23932,N_23022);
or U26218 (N_26218,N_24722,N_23493);
nor U26219 (N_26219,N_23150,N_22681);
nand U26220 (N_26220,N_24705,N_24790);
xor U26221 (N_26221,N_22804,N_24303);
nand U26222 (N_26222,N_22878,N_24732);
xnor U26223 (N_26223,N_24960,N_24920);
xor U26224 (N_26224,N_23877,N_24146);
and U26225 (N_26225,N_24865,N_22876);
xor U26226 (N_26226,N_23784,N_24321);
nor U26227 (N_26227,N_24468,N_22557);
xnor U26228 (N_26228,N_23111,N_24724);
nand U26229 (N_26229,N_24947,N_22774);
nand U26230 (N_26230,N_24776,N_24955);
xnor U26231 (N_26231,N_24752,N_24917);
and U26232 (N_26232,N_22709,N_22611);
and U26233 (N_26233,N_23688,N_22510);
xor U26234 (N_26234,N_24749,N_23487);
xor U26235 (N_26235,N_23228,N_23809);
and U26236 (N_26236,N_23155,N_23982);
nor U26237 (N_26237,N_23516,N_24407);
nand U26238 (N_26238,N_23086,N_24055);
nand U26239 (N_26239,N_23371,N_24116);
or U26240 (N_26240,N_22976,N_22607);
nand U26241 (N_26241,N_22756,N_23211);
xor U26242 (N_26242,N_23654,N_23327);
or U26243 (N_26243,N_24429,N_22530);
nor U26244 (N_26244,N_24987,N_23401);
and U26245 (N_26245,N_23585,N_24122);
nand U26246 (N_26246,N_24864,N_22539);
xor U26247 (N_26247,N_23683,N_22797);
or U26248 (N_26248,N_24656,N_22636);
xor U26249 (N_26249,N_24552,N_23717);
nand U26250 (N_26250,N_24665,N_23200);
nand U26251 (N_26251,N_22642,N_24553);
nand U26252 (N_26252,N_23388,N_22987);
xor U26253 (N_26253,N_24764,N_22943);
nand U26254 (N_26254,N_23642,N_24079);
or U26255 (N_26255,N_23890,N_23365);
or U26256 (N_26256,N_22544,N_24145);
xnor U26257 (N_26257,N_22975,N_22811);
or U26258 (N_26258,N_22553,N_22536);
nor U26259 (N_26259,N_22761,N_24314);
or U26260 (N_26260,N_24099,N_22727);
nor U26261 (N_26261,N_23267,N_23364);
and U26262 (N_26262,N_24173,N_24692);
xor U26263 (N_26263,N_24314,N_23225);
xor U26264 (N_26264,N_22595,N_24247);
xor U26265 (N_26265,N_22688,N_23995);
or U26266 (N_26266,N_24367,N_23216);
and U26267 (N_26267,N_23606,N_24619);
nand U26268 (N_26268,N_23660,N_23599);
nor U26269 (N_26269,N_24932,N_23651);
nor U26270 (N_26270,N_23754,N_24567);
nand U26271 (N_26271,N_22516,N_24244);
nand U26272 (N_26272,N_22803,N_23942);
or U26273 (N_26273,N_23709,N_24165);
or U26274 (N_26274,N_23572,N_24963);
nor U26275 (N_26275,N_24620,N_24038);
and U26276 (N_26276,N_22813,N_23991);
nor U26277 (N_26277,N_24824,N_23045);
or U26278 (N_26278,N_23066,N_23696);
and U26279 (N_26279,N_22528,N_23691);
and U26280 (N_26280,N_23961,N_24469);
nand U26281 (N_26281,N_23183,N_24409);
nand U26282 (N_26282,N_24323,N_24031);
nand U26283 (N_26283,N_24372,N_24821);
nand U26284 (N_26284,N_22976,N_23805);
or U26285 (N_26285,N_23575,N_24794);
nand U26286 (N_26286,N_24882,N_23893);
and U26287 (N_26287,N_23862,N_22991);
or U26288 (N_26288,N_23686,N_23217);
nor U26289 (N_26289,N_22641,N_23086);
xor U26290 (N_26290,N_23589,N_22720);
nand U26291 (N_26291,N_23331,N_24409);
or U26292 (N_26292,N_24200,N_24597);
nand U26293 (N_26293,N_22901,N_23168);
nand U26294 (N_26294,N_24636,N_22874);
nand U26295 (N_26295,N_23939,N_22780);
and U26296 (N_26296,N_23886,N_24564);
xnor U26297 (N_26297,N_24192,N_23326);
or U26298 (N_26298,N_24287,N_23196);
nand U26299 (N_26299,N_24985,N_22832);
and U26300 (N_26300,N_23424,N_24087);
nor U26301 (N_26301,N_24160,N_23499);
xor U26302 (N_26302,N_23737,N_23189);
or U26303 (N_26303,N_23839,N_24325);
or U26304 (N_26304,N_24631,N_22762);
nor U26305 (N_26305,N_24975,N_24757);
and U26306 (N_26306,N_24565,N_24237);
xor U26307 (N_26307,N_22824,N_23065);
nor U26308 (N_26308,N_22578,N_22635);
and U26309 (N_26309,N_24085,N_24982);
and U26310 (N_26310,N_23157,N_22742);
xnor U26311 (N_26311,N_24503,N_22943);
nand U26312 (N_26312,N_24374,N_23689);
and U26313 (N_26313,N_23754,N_23031);
nor U26314 (N_26314,N_23974,N_23676);
xnor U26315 (N_26315,N_23980,N_24183);
nor U26316 (N_26316,N_22864,N_24469);
xnor U26317 (N_26317,N_24451,N_23405);
or U26318 (N_26318,N_24669,N_22702);
xnor U26319 (N_26319,N_24266,N_24864);
or U26320 (N_26320,N_24683,N_24636);
nand U26321 (N_26321,N_22936,N_22941);
xnor U26322 (N_26322,N_22551,N_22928);
and U26323 (N_26323,N_22821,N_24212);
nor U26324 (N_26324,N_22579,N_22727);
and U26325 (N_26325,N_24864,N_22765);
nand U26326 (N_26326,N_24532,N_22909);
nor U26327 (N_26327,N_23218,N_24487);
xor U26328 (N_26328,N_23810,N_23622);
xor U26329 (N_26329,N_24111,N_23774);
nor U26330 (N_26330,N_24831,N_24255);
and U26331 (N_26331,N_24402,N_23305);
or U26332 (N_26332,N_22520,N_23388);
and U26333 (N_26333,N_24016,N_24082);
nor U26334 (N_26334,N_24164,N_23578);
xor U26335 (N_26335,N_23502,N_24530);
nand U26336 (N_26336,N_24759,N_22635);
nand U26337 (N_26337,N_23260,N_22732);
and U26338 (N_26338,N_23729,N_23194);
nor U26339 (N_26339,N_22983,N_23521);
or U26340 (N_26340,N_22899,N_22886);
and U26341 (N_26341,N_22506,N_24388);
xnor U26342 (N_26342,N_23399,N_24242);
or U26343 (N_26343,N_24823,N_24306);
and U26344 (N_26344,N_23083,N_24409);
xor U26345 (N_26345,N_23569,N_24097);
or U26346 (N_26346,N_24483,N_24664);
xor U26347 (N_26347,N_23944,N_22624);
nand U26348 (N_26348,N_23084,N_24382);
and U26349 (N_26349,N_23363,N_24158);
or U26350 (N_26350,N_24787,N_23048);
xnor U26351 (N_26351,N_22736,N_22881);
nand U26352 (N_26352,N_23929,N_23075);
nor U26353 (N_26353,N_24145,N_23958);
nand U26354 (N_26354,N_24667,N_24941);
xnor U26355 (N_26355,N_22556,N_22656);
nor U26356 (N_26356,N_24589,N_22978);
or U26357 (N_26357,N_23573,N_24998);
xor U26358 (N_26358,N_24640,N_22651);
and U26359 (N_26359,N_22842,N_24281);
or U26360 (N_26360,N_23977,N_22805);
xnor U26361 (N_26361,N_23896,N_22853);
nand U26362 (N_26362,N_24336,N_23823);
and U26363 (N_26363,N_24271,N_23440);
nor U26364 (N_26364,N_23905,N_24077);
nand U26365 (N_26365,N_23532,N_22905);
or U26366 (N_26366,N_24282,N_23450);
nand U26367 (N_26367,N_22790,N_24661);
xor U26368 (N_26368,N_23304,N_24392);
xnor U26369 (N_26369,N_23722,N_22889);
xor U26370 (N_26370,N_23075,N_22980);
and U26371 (N_26371,N_24073,N_23992);
nor U26372 (N_26372,N_23380,N_24127);
nor U26373 (N_26373,N_24381,N_23075);
xor U26374 (N_26374,N_23972,N_23832);
xor U26375 (N_26375,N_22951,N_22654);
or U26376 (N_26376,N_23037,N_22569);
nor U26377 (N_26377,N_22906,N_23490);
and U26378 (N_26378,N_23074,N_23814);
or U26379 (N_26379,N_22814,N_23232);
and U26380 (N_26380,N_23704,N_24317);
or U26381 (N_26381,N_23597,N_22939);
or U26382 (N_26382,N_23705,N_22542);
or U26383 (N_26383,N_22909,N_23034);
and U26384 (N_26384,N_24300,N_22949);
and U26385 (N_26385,N_24197,N_23908);
xnor U26386 (N_26386,N_24371,N_24799);
nand U26387 (N_26387,N_22771,N_24002);
nand U26388 (N_26388,N_23172,N_24288);
or U26389 (N_26389,N_24573,N_24089);
xor U26390 (N_26390,N_24409,N_23462);
nor U26391 (N_26391,N_23733,N_24272);
nor U26392 (N_26392,N_24667,N_23503);
xnor U26393 (N_26393,N_23249,N_24107);
xor U26394 (N_26394,N_23228,N_24976);
nand U26395 (N_26395,N_23025,N_22676);
and U26396 (N_26396,N_23881,N_23570);
nor U26397 (N_26397,N_24863,N_22991);
and U26398 (N_26398,N_24622,N_23262);
and U26399 (N_26399,N_24583,N_22570);
nand U26400 (N_26400,N_24569,N_22997);
xnor U26401 (N_26401,N_22686,N_24114);
and U26402 (N_26402,N_23244,N_23440);
and U26403 (N_26403,N_22763,N_22900);
or U26404 (N_26404,N_23546,N_24961);
xor U26405 (N_26405,N_24385,N_23236);
nand U26406 (N_26406,N_22996,N_23440);
nor U26407 (N_26407,N_24467,N_22919);
and U26408 (N_26408,N_23562,N_22672);
nor U26409 (N_26409,N_24606,N_24942);
nand U26410 (N_26410,N_23333,N_22905);
and U26411 (N_26411,N_22749,N_24627);
nand U26412 (N_26412,N_24061,N_23873);
and U26413 (N_26413,N_23726,N_22797);
and U26414 (N_26414,N_23436,N_24901);
nor U26415 (N_26415,N_23044,N_22706);
xnor U26416 (N_26416,N_23472,N_23803);
nand U26417 (N_26417,N_24495,N_23702);
nor U26418 (N_26418,N_23967,N_24646);
and U26419 (N_26419,N_22961,N_23323);
nand U26420 (N_26420,N_23767,N_22773);
nand U26421 (N_26421,N_23984,N_24696);
or U26422 (N_26422,N_23960,N_24993);
xnor U26423 (N_26423,N_22710,N_23521);
nand U26424 (N_26424,N_22543,N_22559);
or U26425 (N_26425,N_23513,N_22967);
nand U26426 (N_26426,N_22639,N_24486);
nor U26427 (N_26427,N_23936,N_22834);
nor U26428 (N_26428,N_23423,N_22948);
or U26429 (N_26429,N_24730,N_22969);
nand U26430 (N_26430,N_23087,N_22513);
xor U26431 (N_26431,N_23565,N_23839);
or U26432 (N_26432,N_23981,N_23608);
and U26433 (N_26433,N_23792,N_23069);
xnor U26434 (N_26434,N_23686,N_22503);
nand U26435 (N_26435,N_22612,N_24765);
nand U26436 (N_26436,N_23255,N_24747);
and U26437 (N_26437,N_24317,N_22959);
or U26438 (N_26438,N_24305,N_23623);
nor U26439 (N_26439,N_22681,N_24441);
xnor U26440 (N_26440,N_22642,N_23360);
xor U26441 (N_26441,N_23172,N_24598);
or U26442 (N_26442,N_22729,N_23721);
or U26443 (N_26443,N_22881,N_22508);
nor U26444 (N_26444,N_23493,N_24869);
xor U26445 (N_26445,N_23171,N_23871);
nand U26446 (N_26446,N_22960,N_24081);
or U26447 (N_26447,N_24972,N_24651);
nand U26448 (N_26448,N_23368,N_23077);
nor U26449 (N_26449,N_22602,N_24364);
nor U26450 (N_26450,N_23531,N_22611);
xnor U26451 (N_26451,N_22949,N_23587);
nand U26452 (N_26452,N_24601,N_23339);
and U26453 (N_26453,N_23565,N_24686);
or U26454 (N_26454,N_22890,N_24563);
xor U26455 (N_26455,N_24136,N_23405);
and U26456 (N_26456,N_23821,N_23524);
xnor U26457 (N_26457,N_22521,N_23684);
and U26458 (N_26458,N_22658,N_23203);
and U26459 (N_26459,N_23402,N_23632);
and U26460 (N_26460,N_24742,N_23172);
nand U26461 (N_26461,N_23773,N_22670);
xnor U26462 (N_26462,N_23608,N_23027);
nand U26463 (N_26463,N_24313,N_23924);
nand U26464 (N_26464,N_24770,N_24452);
or U26465 (N_26465,N_23702,N_24050);
nor U26466 (N_26466,N_24361,N_22782);
nor U26467 (N_26467,N_24684,N_22696);
and U26468 (N_26468,N_23211,N_24004);
nor U26469 (N_26469,N_23425,N_23480);
xnor U26470 (N_26470,N_23139,N_23755);
xor U26471 (N_26471,N_23659,N_22579);
xnor U26472 (N_26472,N_24283,N_23449);
nand U26473 (N_26473,N_22585,N_22500);
nand U26474 (N_26474,N_22623,N_23897);
nor U26475 (N_26475,N_23747,N_24427);
or U26476 (N_26476,N_23550,N_24359);
nor U26477 (N_26477,N_23775,N_23966);
nand U26478 (N_26478,N_23158,N_23028);
nor U26479 (N_26479,N_22848,N_23713);
nor U26480 (N_26480,N_22760,N_23266);
nand U26481 (N_26481,N_22758,N_24528);
nand U26482 (N_26482,N_23398,N_23712);
nand U26483 (N_26483,N_23410,N_24118);
and U26484 (N_26484,N_24733,N_24638);
and U26485 (N_26485,N_24396,N_22940);
and U26486 (N_26486,N_22937,N_23964);
and U26487 (N_26487,N_22715,N_23918);
and U26488 (N_26488,N_23171,N_24761);
nand U26489 (N_26489,N_24893,N_23395);
nand U26490 (N_26490,N_22852,N_23501);
nand U26491 (N_26491,N_23975,N_24378);
or U26492 (N_26492,N_23276,N_24382);
and U26493 (N_26493,N_23493,N_23563);
and U26494 (N_26494,N_22872,N_23677);
xor U26495 (N_26495,N_24792,N_22754);
or U26496 (N_26496,N_24329,N_24834);
nand U26497 (N_26497,N_23352,N_24603);
nor U26498 (N_26498,N_23778,N_24436);
nor U26499 (N_26499,N_22822,N_24273);
or U26500 (N_26500,N_24362,N_23330);
and U26501 (N_26501,N_24016,N_24470);
nor U26502 (N_26502,N_23763,N_24307);
or U26503 (N_26503,N_22810,N_23240);
or U26504 (N_26504,N_23474,N_23583);
xor U26505 (N_26505,N_24635,N_24696);
nand U26506 (N_26506,N_24385,N_24144);
nand U26507 (N_26507,N_22805,N_22559);
nor U26508 (N_26508,N_24715,N_24705);
and U26509 (N_26509,N_23234,N_22679);
or U26510 (N_26510,N_24707,N_23585);
and U26511 (N_26511,N_23950,N_23898);
nand U26512 (N_26512,N_23519,N_23879);
nand U26513 (N_26513,N_23005,N_24227);
xnor U26514 (N_26514,N_24191,N_22642);
nor U26515 (N_26515,N_22560,N_24913);
nor U26516 (N_26516,N_22656,N_22863);
xnor U26517 (N_26517,N_22759,N_24088);
nor U26518 (N_26518,N_22628,N_23296);
xnor U26519 (N_26519,N_24738,N_24252);
xor U26520 (N_26520,N_24769,N_24154);
or U26521 (N_26521,N_24930,N_24508);
or U26522 (N_26522,N_22811,N_23539);
and U26523 (N_26523,N_24525,N_23288);
nand U26524 (N_26524,N_24910,N_24270);
or U26525 (N_26525,N_22519,N_24019);
and U26526 (N_26526,N_23525,N_22575);
or U26527 (N_26527,N_22504,N_22999);
or U26528 (N_26528,N_23698,N_24575);
nor U26529 (N_26529,N_23482,N_23046);
or U26530 (N_26530,N_23980,N_23257);
nand U26531 (N_26531,N_24972,N_24039);
nand U26532 (N_26532,N_23910,N_23322);
nor U26533 (N_26533,N_23021,N_24317);
nand U26534 (N_26534,N_24404,N_24191);
nor U26535 (N_26535,N_23558,N_24210);
xor U26536 (N_26536,N_24378,N_22824);
nand U26537 (N_26537,N_23142,N_24007);
xor U26538 (N_26538,N_23683,N_22760);
and U26539 (N_26539,N_24267,N_23150);
and U26540 (N_26540,N_22873,N_24704);
nor U26541 (N_26541,N_23005,N_24382);
nor U26542 (N_26542,N_24280,N_23667);
and U26543 (N_26543,N_23123,N_24100);
or U26544 (N_26544,N_24932,N_22724);
nor U26545 (N_26545,N_23286,N_23000);
nor U26546 (N_26546,N_23511,N_24618);
or U26547 (N_26547,N_24288,N_22609);
nor U26548 (N_26548,N_23804,N_23829);
or U26549 (N_26549,N_22681,N_22892);
nand U26550 (N_26550,N_24135,N_23238);
nor U26551 (N_26551,N_24065,N_22884);
nor U26552 (N_26552,N_23767,N_22899);
or U26553 (N_26553,N_23563,N_22777);
and U26554 (N_26554,N_23009,N_22903);
and U26555 (N_26555,N_22929,N_23407);
and U26556 (N_26556,N_23010,N_24351);
nor U26557 (N_26557,N_23983,N_23563);
and U26558 (N_26558,N_23940,N_24652);
nor U26559 (N_26559,N_24639,N_24706);
and U26560 (N_26560,N_22503,N_24344);
nand U26561 (N_26561,N_23356,N_22577);
xor U26562 (N_26562,N_22899,N_23084);
nor U26563 (N_26563,N_22689,N_22951);
nand U26564 (N_26564,N_23897,N_23337);
and U26565 (N_26565,N_22533,N_24307);
or U26566 (N_26566,N_23419,N_24916);
or U26567 (N_26567,N_23360,N_22884);
xor U26568 (N_26568,N_22927,N_23102);
nor U26569 (N_26569,N_23917,N_22764);
xnor U26570 (N_26570,N_22514,N_24048);
xnor U26571 (N_26571,N_22930,N_22621);
nor U26572 (N_26572,N_24745,N_24286);
nor U26573 (N_26573,N_23056,N_23764);
nand U26574 (N_26574,N_22645,N_22622);
nor U26575 (N_26575,N_24669,N_22969);
or U26576 (N_26576,N_24206,N_22686);
nor U26577 (N_26577,N_22815,N_22648);
or U26578 (N_26578,N_23720,N_23853);
nor U26579 (N_26579,N_23296,N_23678);
and U26580 (N_26580,N_22678,N_23058);
nand U26581 (N_26581,N_24687,N_23293);
or U26582 (N_26582,N_23999,N_24289);
nand U26583 (N_26583,N_24294,N_24438);
xnor U26584 (N_26584,N_22943,N_23051);
and U26585 (N_26585,N_23362,N_22704);
nor U26586 (N_26586,N_23603,N_23073);
or U26587 (N_26587,N_23988,N_22683);
xor U26588 (N_26588,N_23161,N_22650);
or U26589 (N_26589,N_24021,N_23291);
nand U26590 (N_26590,N_24748,N_23307);
and U26591 (N_26591,N_22506,N_23525);
and U26592 (N_26592,N_22944,N_22624);
or U26593 (N_26593,N_24449,N_23758);
nor U26594 (N_26594,N_24480,N_24870);
nor U26595 (N_26595,N_24403,N_23978);
nand U26596 (N_26596,N_23456,N_24819);
xor U26597 (N_26597,N_22583,N_23034);
nor U26598 (N_26598,N_23462,N_23730);
nor U26599 (N_26599,N_22933,N_24161);
xor U26600 (N_26600,N_24370,N_24702);
nand U26601 (N_26601,N_22738,N_24840);
or U26602 (N_26602,N_23035,N_23805);
nor U26603 (N_26603,N_24629,N_23914);
nand U26604 (N_26604,N_22642,N_23439);
nand U26605 (N_26605,N_24820,N_22771);
xnor U26606 (N_26606,N_23625,N_24624);
nand U26607 (N_26607,N_24357,N_23559);
xor U26608 (N_26608,N_23254,N_23044);
nor U26609 (N_26609,N_24937,N_23361);
nor U26610 (N_26610,N_24260,N_23534);
or U26611 (N_26611,N_24551,N_24535);
nand U26612 (N_26612,N_23482,N_23630);
xnor U26613 (N_26613,N_23154,N_22726);
and U26614 (N_26614,N_24899,N_24747);
and U26615 (N_26615,N_24205,N_22557);
nor U26616 (N_26616,N_23515,N_23631);
xor U26617 (N_26617,N_22944,N_24311);
xor U26618 (N_26618,N_23106,N_24495);
and U26619 (N_26619,N_24936,N_24984);
nor U26620 (N_26620,N_23806,N_23584);
nor U26621 (N_26621,N_24149,N_24285);
xnor U26622 (N_26622,N_24392,N_22610);
nor U26623 (N_26623,N_23710,N_22812);
nand U26624 (N_26624,N_24007,N_23809);
xor U26625 (N_26625,N_22577,N_23393);
nand U26626 (N_26626,N_23823,N_23335);
nand U26627 (N_26627,N_23961,N_24449);
or U26628 (N_26628,N_23494,N_22534);
nor U26629 (N_26629,N_23784,N_23319);
nor U26630 (N_26630,N_22769,N_24900);
nand U26631 (N_26631,N_24193,N_24805);
nor U26632 (N_26632,N_24927,N_23486);
or U26633 (N_26633,N_23862,N_23128);
and U26634 (N_26634,N_24921,N_22731);
nand U26635 (N_26635,N_24588,N_22795);
nand U26636 (N_26636,N_24593,N_23242);
or U26637 (N_26637,N_22611,N_23943);
or U26638 (N_26638,N_23552,N_23714);
and U26639 (N_26639,N_23298,N_24847);
nand U26640 (N_26640,N_22894,N_22750);
nor U26641 (N_26641,N_23531,N_24287);
nand U26642 (N_26642,N_24325,N_23251);
xor U26643 (N_26643,N_23113,N_23425);
xor U26644 (N_26644,N_24542,N_22803);
xor U26645 (N_26645,N_24296,N_22512);
nor U26646 (N_26646,N_24572,N_23502);
nand U26647 (N_26647,N_23551,N_24129);
nor U26648 (N_26648,N_24028,N_23534);
nor U26649 (N_26649,N_24775,N_23742);
xnor U26650 (N_26650,N_23597,N_24732);
nand U26651 (N_26651,N_24849,N_24487);
xnor U26652 (N_26652,N_22641,N_23008);
or U26653 (N_26653,N_24795,N_24191);
nand U26654 (N_26654,N_24338,N_23645);
nor U26655 (N_26655,N_23525,N_23528);
or U26656 (N_26656,N_22793,N_23466);
and U26657 (N_26657,N_24903,N_22504);
xor U26658 (N_26658,N_22586,N_22535);
xnor U26659 (N_26659,N_23850,N_22593);
xnor U26660 (N_26660,N_23991,N_23154);
nand U26661 (N_26661,N_24758,N_23538);
nand U26662 (N_26662,N_24679,N_24782);
or U26663 (N_26663,N_24742,N_23002);
or U26664 (N_26664,N_23654,N_23857);
and U26665 (N_26665,N_23000,N_22993);
and U26666 (N_26666,N_24049,N_24855);
and U26667 (N_26667,N_24633,N_24421);
nor U26668 (N_26668,N_22654,N_24734);
nand U26669 (N_26669,N_23540,N_23185);
and U26670 (N_26670,N_24413,N_24867);
xnor U26671 (N_26671,N_23867,N_22540);
nand U26672 (N_26672,N_23389,N_24136);
nor U26673 (N_26673,N_22662,N_24744);
nor U26674 (N_26674,N_23912,N_22905);
nor U26675 (N_26675,N_22734,N_23202);
nand U26676 (N_26676,N_23623,N_24822);
or U26677 (N_26677,N_23572,N_24342);
nand U26678 (N_26678,N_23286,N_23768);
xnor U26679 (N_26679,N_23127,N_22544);
xnor U26680 (N_26680,N_24890,N_23141);
xnor U26681 (N_26681,N_23623,N_24175);
and U26682 (N_26682,N_22546,N_23984);
nor U26683 (N_26683,N_23518,N_24029);
or U26684 (N_26684,N_24966,N_22815);
nor U26685 (N_26685,N_24164,N_24722);
nand U26686 (N_26686,N_24133,N_24390);
xnor U26687 (N_26687,N_23286,N_23816);
nand U26688 (N_26688,N_23313,N_24367);
and U26689 (N_26689,N_24485,N_24685);
and U26690 (N_26690,N_23828,N_23256);
nand U26691 (N_26691,N_23540,N_23455);
nor U26692 (N_26692,N_23987,N_23077);
nor U26693 (N_26693,N_24400,N_24001);
and U26694 (N_26694,N_23906,N_24567);
and U26695 (N_26695,N_23120,N_24605);
or U26696 (N_26696,N_23241,N_23990);
xnor U26697 (N_26697,N_23827,N_24996);
or U26698 (N_26698,N_24523,N_22875);
or U26699 (N_26699,N_24264,N_24339);
or U26700 (N_26700,N_23257,N_24177);
and U26701 (N_26701,N_24180,N_23077);
xor U26702 (N_26702,N_24648,N_24183);
xor U26703 (N_26703,N_22631,N_23566);
nand U26704 (N_26704,N_23671,N_22612);
nand U26705 (N_26705,N_23412,N_23951);
or U26706 (N_26706,N_24203,N_24630);
and U26707 (N_26707,N_24854,N_24935);
nand U26708 (N_26708,N_24871,N_24499);
nor U26709 (N_26709,N_24571,N_23155);
and U26710 (N_26710,N_23289,N_23610);
and U26711 (N_26711,N_24153,N_24740);
and U26712 (N_26712,N_23387,N_23364);
and U26713 (N_26713,N_23315,N_24951);
and U26714 (N_26714,N_24613,N_23718);
and U26715 (N_26715,N_22531,N_23917);
xor U26716 (N_26716,N_24458,N_24351);
and U26717 (N_26717,N_24596,N_24061);
nor U26718 (N_26718,N_23967,N_23191);
nor U26719 (N_26719,N_22845,N_23387);
and U26720 (N_26720,N_23031,N_23764);
nor U26721 (N_26721,N_23753,N_24998);
nand U26722 (N_26722,N_24410,N_23124);
nor U26723 (N_26723,N_22990,N_24770);
and U26724 (N_26724,N_24897,N_24893);
nor U26725 (N_26725,N_23277,N_24204);
or U26726 (N_26726,N_23417,N_24161);
nand U26727 (N_26727,N_24166,N_22810);
nand U26728 (N_26728,N_23312,N_24029);
and U26729 (N_26729,N_23770,N_23018);
and U26730 (N_26730,N_23638,N_24336);
nor U26731 (N_26731,N_23966,N_24074);
and U26732 (N_26732,N_22972,N_23605);
and U26733 (N_26733,N_22661,N_24843);
xor U26734 (N_26734,N_22508,N_24371);
xnor U26735 (N_26735,N_22698,N_24347);
nor U26736 (N_26736,N_24795,N_22558);
xor U26737 (N_26737,N_23003,N_23286);
xnor U26738 (N_26738,N_23260,N_23009);
and U26739 (N_26739,N_24442,N_24265);
nand U26740 (N_26740,N_22826,N_24298);
nor U26741 (N_26741,N_23221,N_24780);
and U26742 (N_26742,N_23029,N_24149);
or U26743 (N_26743,N_23450,N_24727);
or U26744 (N_26744,N_23075,N_24025);
nor U26745 (N_26745,N_23107,N_22935);
or U26746 (N_26746,N_22549,N_22876);
and U26747 (N_26747,N_23997,N_22803);
and U26748 (N_26748,N_23747,N_22835);
xnor U26749 (N_26749,N_24808,N_23916);
and U26750 (N_26750,N_24549,N_23033);
nand U26751 (N_26751,N_23176,N_23876);
and U26752 (N_26752,N_22725,N_24391);
xnor U26753 (N_26753,N_23874,N_23756);
nand U26754 (N_26754,N_22695,N_24242);
or U26755 (N_26755,N_24834,N_24082);
and U26756 (N_26756,N_24871,N_24385);
xnor U26757 (N_26757,N_24146,N_24859);
xor U26758 (N_26758,N_22630,N_24198);
and U26759 (N_26759,N_24024,N_23028);
and U26760 (N_26760,N_24674,N_23928);
nand U26761 (N_26761,N_23632,N_23852);
nor U26762 (N_26762,N_23603,N_24400);
xnor U26763 (N_26763,N_23561,N_24421);
and U26764 (N_26764,N_24001,N_24953);
nand U26765 (N_26765,N_23829,N_22698);
nor U26766 (N_26766,N_23621,N_22605);
nor U26767 (N_26767,N_24454,N_23825);
xor U26768 (N_26768,N_23958,N_24305);
nor U26769 (N_26769,N_22820,N_24918);
and U26770 (N_26770,N_22829,N_24360);
xor U26771 (N_26771,N_24819,N_24295);
nor U26772 (N_26772,N_23542,N_24921);
or U26773 (N_26773,N_23434,N_23100);
nand U26774 (N_26774,N_23406,N_23123);
nor U26775 (N_26775,N_23225,N_23031);
or U26776 (N_26776,N_23688,N_23454);
or U26777 (N_26777,N_24278,N_23807);
or U26778 (N_26778,N_23478,N_23961);
and U26779 (N_26779,N_23396,N_24615);
or U26780 (N_26780,N_23152,N_23889);
xnor U26781 (N_26781,N_22918,N_24392);
nor U26782 (N_26782,N_23736,N_24253);
nand U26783 (N_26783,N_23840,N_22524);
nand U26784 (N_26784,N_24844,N_23330);
xnor U26785 (N_26785,N_24962,N_23717);
nor U26786 (N_26786,N_23903,N_24776);
or U26787 (N_26787,N_23897,N_23025);
nand U26788 (N_26788,N_23916,N_24257);
nor U26789 (N_26789,N_22512,N_24781);
nor U26790 (N_26790,N_24890,N_24320);
or U26791 (N_26791,N_23649,N_24472);
xnor U26792 (N_26792,N_24354,N_24041);
nand U26793 (N_26793,N_23860,N_24576);
or U26794 (N_26794,N_23633,N_24762);
or U26795 (N_26795,N_23485,N_24913);
xnor U26796 (N_26796,N_23000,N_23441);
or U26797 (N_26797,N_22825,N_22592);
or U26798 (N_26798,N_24744,N_22807);
or U26799 (N_26799,N_23986,N_24324);
and U26800 (N_26800,N_24210,N_23772);
nor U26801 (N_26801,N_22764,N_23221);
xor U26802 (N_26802,N_24281,N_22537);
or U26803 (N_26803,N_23429,N_24687);
xor U26804 (N_26804,N_22514,N_23538);
nand U26805 (N_26805,N_24633,N_23936);
and U26806 (N_26806,N_23145,N_22955);
nor U26807 (N_26807,N_22606,N_22590);
xnor U26808 (N_26808,N_22962,N_24254);
nand U26809 (N_26809,N_22817,N_22958);
or U26810 (N_26810,N_24010,N_24437);
nand U26811 (N_26811,N_23046,N_24261);
nand U26812 (N_26812,N_24241,N_24177);
xnor U26813 (N_26813,N_24212,N_24521);
nor U26814 (N_26814,N_23132,N_23648);
nor U26815 (N_26815,N_24188,N_22800);
nand U26816 (N_26816,N_23693,N_23352);
and U26817 (N_26817,N_24182,N_22936);
and U26818 (N_26818,N_22959,N_23137);
nand U26819 (N_26819,N_24763,N_24052);
or U26820 (N_26820,N_23321,N_23951);
nor U26821 (N_26821,N_22972,N_23373);
and U26822 (N_26822,N_24003,N_24660);
nor U26823 (N_26823,N_24073,N_23380);
nor U26824 (N_26824,N_22858,N_23742);
nand U26825 (N_26825,N_24047,N_24433);
or U26826 (N_26826,N_23175,N_23369);
nor U26827 (N_26827,N_23018,N_22951);
nor U26828 (N_26828,N_23722,N_23249);
xor U26829 (N_26829,N_24718,N_24977);
nor U26830 (N_26830,N_23529,N_24014);
or U26831 (N_26831,N_22642,N_23928);
and U26832 (N_26832,N_24153,N_23320);
xor U26833 (N_26833,N_23772,N_23059);
and U26834 (N_26834,N_23870,N_24790);
or U26835 (N_26835,N_24405,N_22849);
nand U26836 (N_26836,N_23354,N_24934);
and U26837 (N_26837,N_22885,N_22611);
nand U26838 (N_26838,N_23019,N_22676);
nand U26839 (N_26839,N_23145,N_24798);
or U26840 (N_26840,N_23858,N_22888);
xnor U26841 (N_26841,N_24100,N_23352);
nand U26842 (N_26842,N_23210,N_22782);
or U26843 (N_26843,N_23949,N_24295);
or U26844 (N_26844,N_24776,N_24450);
nor U26845 (N_26845,N_24654,N_22537);
or U26846 (N_26846,N_24932,N_24850);
and U26847 (N_26847,N_22718,N_23264);
nand U26848 (N_26848,N_23374,N_24099);
xor U26849 (N_26849,N_22734,N_23702);
nand U26850 (N_26850,N_24572,N_24711);
nand U26851 (N_26851,N_24722,N_22934);
or U26852 (N_26852,N_22509,N_23322);
nand U26853 (N_26853,N_22573,N_23829);
nor U26854 (N_26854,N_23913,N_22835);
and U26855 (N_26855,N_22640,N_24950);
and U26856 (N_26856,N_24209,N_23537);
nand U26857 (N_26857,N_24564,N_23236);
or U26858 (N_26858,N_24110,N_24362);
or U26859 (N_26859,N_23281,N_23452);
nor U26860 (N_26860,N_23457,N_23759);
and U26861 (N_26861,N_23910,N_23307);
or U26862 (N_26862,N_24297,N_24468);
xnor U26863 (N_26863,N_22781,N_22772);
nor U26864 (N_26864,N_22667,N_24834);
nand U26865 (N_26865,N_23964,N_24253);
nor U26866 (N_26866,N_24701,N_23066);
or U26867 (N_26867,N_24709,N_24794);
nor U26868 (N_26868,N_24572,N_23554);
nor U26869 (N_26869,N_23976,N_24821);
or U26870 (N_26870,N_23565,N_24765);
or U26871 (N_26871,N_23483,N_24950);
nor U26872 (N_26872,N_24625,N_24812);
xnor U26873 (N_26873,N_22600,N_23310);
nor U26874 (N_26874,N_23395,N_24137);
nand U26875 (N_26875,N_23527,N_23658);
nor U26876 (N_26876,N_23135,N_23995);
or U26877 (N_26877,N_23574,N_23244);
nor U26878 (N_26878,N_24828,N_22999);
nand U26879 (N_26879,N_22963,N_24530);
nor U26880 (N_26880,N_22942,N_23334);
and U26881 (N_26881,N_24149,N_22677);
and U26882 (N_26882,N_22892,N_23884);
nor U26883 (N_26883,N_23396,N_24680);
xor U26884 (N_26884,N_23102,N_24750);
nor U26885 (N_26885,N_24837,N_24613);
xor U26886 (N_26886,N_23801,N_23931);
or U26887 (N_26887,N_22958,N_23700);
or U26888 (N_26888,N_23098,N_22807);
and U26889 (N_26889,N_23192,N_23574);
nor U26890 (N_26890,N_23575,N_22907);
xnor U26891 (N_26891,N_24871,N_23471);
nand U26892 (N_26892,N_22908,N_23034);
and U26893 (N_26893,N_23109,N_24325);
nand U26894 (N_26894,N_23373,N_23911);
nand U26895 (N_26895,N_24343,N_24754);
xnor U26896 (N_26896,N_24690,N_24553);
nand U26897 (N_26897,N_22560,N_23496);
nor U26898 (N_26898,N_24521,N_22788);
xor U26899 (N_26899,N_24681,N_23404);
and U26900 (N_26900,N_23007,N_23873);
nor U26901 (N_26901,N_24167,N_24913);
xor U26902 (N_26902,N_22773,N_24056);
and U26903 (N_26903,N_24357,N_23394);
nand U26904 (N_26904,N_23393,N_22766);
and U26905 (N_26905,N_22594,N_23930);
xnor U26906 (N_26906,N_24110,N_24008);
nand U26907 (N_26907,N_23006,N_22982);
nor U26908 (N_26908,N_24327,N_24106);
or U26909 (N_26909,N_22729,N_24032);
or U26910 (N_26910,N_24518,N_24196);
nor U26911 (N_26911,N_23746,N_24745);
xor U26912 (N_26912,N_23522,N_23914);
nand U26913 (N_26913,N_23695,N_24327);
nor U26914 (N_26914,N_24636,N_24595);
or U26915 (N_26915,N_24737,N_23238);
nand U26916 (N_26916,N_22730,N_22822);
nand U26917 (N_26917,N_23857,N_22763);
nand U26918 (N_26918,N_24724,N_23682);
xnor U26919 (N_26919,N_23992,N_24617);
xnor U26920 (N_26920,N_24936,N_22695);
nor U26921 (N_26921,N_23640,N_24731);
nor U26922 (N_26922,N_24110,N_22629);
nor U26923 (N_26923,N_24877,N_23407);
nor U26924 (N_26924,N_23152,N_24882);
xor U26925 (N_26925,N_22652,N_23992);
xnor U26926 (N_26926,N_22902,N_23812);
nand U26927 (N_26927,N_24196,N_24434);
and U26928 (N_26928,N_24274,N_23369);
and U26929 (N_26929,N_23355,N_24819);
and U26930 (N_26930,N_24505,N_24511);
nand U26931 (N_26931,N_24625,N_23787);
or U26932 (N_26932,N_22973,N_22872);
nor U26933 (N_26933,N_24150,N_24594);
and U26934 (N_26934,N_24934,N_23966);
xnor U26935 (N_26935,N_22999,N_22937);
nor U26936 (N_26936,N_23702,N_23875);
and U26937 (N_26937,N_23881,N_23592);
xor U26938 (N_26938,N_24225,N_23057);
and U26939 (N_26939,N_24394,N_23324);
nor U26940 (N_26940,N_24248,N_22813);
nor U26941 (N_26941,N_23468,N_22812);
xnor U26942 (N_26942,N_23514,N_24197);
and U26943 (N_26943,N_23385,N_24344);
nor U26944 (N_26944,N_23602,N_24218);
nand U26945 (N_26945,N_23838,N_23687);
or U26946 (N_26946,N_23849,N_23829);
nand U26947 (N_26947,N_22731,N_22745);
xor U26948 (N_26948,N_22943,N_24190);
nand U26949 (N_26949,N_22814,N_23799);
and U26950 (N_26950,N_22852,N_23198);
nor U26951 (N_26951,N_24453,N_22673);
or U26952 (N_26952,N_24336,N_23082);
nand U26953 (N_26953,N_23976,N_22730);
nor U26954 (N_26954,N_23691,N_22575);
nand U26955 (N_26955,N_24097,N_24609);
or U26956 (N_26956,N_23128,N_24270);
nor U26957 (N_26957,N_23443,N_23562);
xnor U26958 (N_26958,N_24544,N_23415);
or U26959 (N_26959,N_24170,N_24127);
or U26960 (N_26960,N_23765,N_24190);
xnor U26961 (N_26961,N_22677,N_22802);
nor U26962 (N_26962,N_23937,N_24849);
xnor U26963 (N_26963,N_22855,N_22876);
xor U26964 (N_26964,N_22982,N_24524);
or U26965 (N_26965,N_24509,N_22532);
nand U26966 (N_26966,N_24176,N_23635);
and U26967 (N_26967,N_23435,N_24094);
nor U26968 (N_26968,N_22516,N_23767);
nand U26969 (N_26969,N_24002,N_23114);
or U26970 (N_26970,N_22635,N_24758);
xor U26971 (N_26971,N_24439,N_23761);
xnor U26972 (N_26972,N_23405,N_23476);
nor U26973 (N_26973,N_22537,N_24937);
nor U26974 (N_26974,N_24208,N_23853);
nor U26975 (N_26975,N_24475,N_22855);
or U26976 (N_26976,N_23743,N_24574);
nand U26977 (N_26977,N_23624,N_23865);
xnor U26978 (N_26978,N_22991,N_22778);
and U26979 (N_26979,N_23372,N_23980);
xnor U26980 (N_26980,N_24767,N_23169);
nand U26981 (N_26981,N_24189,N_24114);
or U26982 (N_26982,N_24432,N_22740);
or U26983 (N_26983,N_23779,N_24662);
nand U26984 (N_26984,N_22988,N_22878);
nand U26985 (N_26985,N_24315,N_22826);
xnor U26986 (N_26986,N_24151,N_24097);
nand U26987 (N_26987,N_22751,N_23324);
nor U26988 (N_26988,N_24878,N_24406);
and U26989 (N_26989,N_22814,N_24056);
nor U26990 (N_26990,N_24781,N_22900);
xnor U26991 (N_26991,N_24348,N_23804);
and U26992 (N_26992,N_24912,N_24562);
nand U26993 (N_26993,N_23349,N_22516);
nor U26994 (N_26994,N_24327,N_23624);
nor U26995 (N_26995,N_22939,N_24123);
or U26996 (N_26996,N_24786,N_23988);
nor U26997 (N_26997,N_23911,N_23220);
or U26998 (N_26998,N_23888,N_22983);
and U26999 (N_26999,N_23522,N_24899);
xnor U27000 (N_27000,N_24925,N_23708);
or U27001 (N_27001,N_23511,N_23090);
nand U27002 (N_27002,N_24223,N_24375);
xor U27003 (N_27003,N_24801,N_23275);
nand U27004 (N_27004,N_23161,N_24355);
or U27005 (N_27005,N_22612,N_22983);
or U27006 (N_27006,N_24229,N_24168);
or U27007 (N_27007,N_23598,N_23851);
and U27008 (N_27008,N_24026,N_23135);
nand U27009 (N_27009,N_24836,N_23193);
and U27010 (N_27010,N_22773,N_22600);
nand U27011 (N_27011,N_23783,N_22894);
nor U27012 (N_27012,N_24587,N_22805);
nand U27013 (N_27013,N_23774,N_23632);
or U27014 (N_27014,N_24741,N_22869);
nand U27015 (N_27015,N_23278,N_23267);
nor U27016 (N_27016,N_22734,N_24320);
xor U27017 (N_27017,N_22511,N_24414);
xor U27018 (N_27018,N_24339,N_24474);
xor U27019 (N_27019,N_22823,N_23580);
nor U27020 (N_27020,N_23818,N_24601);
or U27021 (N_27021,N_24412,N_24860);
xor U27022 (N_27022,N_24929,N_23040);
and U27023 (N_27023,N_23708,N_22811);
nor U27024 (N_27024,N_23151,N_23790);
xnor U27025 (N_27025,N_23450,N_24520);
nor U27026 (N_27026,N_24481,N_24821);
or U27027 (N_27027,N_22653,N_22879);
nand U27028 (N_27028,N_22595,N_23819);
nand U27029 (N_27029,N_23331,N_24614);
or U27030 (N_27030,N_24323,N_23110);
and U27031 (N_27031,N_23742,N_23736);
and U27032 (N_27032,N_23677,N_24868);
nand U27033 (N_27033,N_24696,N_22753);
and U27034 (N_27034,N_24958,N_24270);
or U27035 (N_27035,N_22573,N_23130);
xor U27036 (N_27036,N_23658,N_23514);
nand U27037 (N_27037,N_23993,N_23219);
and U27038 (N_27038,N_23102,N_24740);
xnor U27039 (N_27039,N_24720,N_22612);
xor U27040 (N_27040,N_23627,N_24272);
nor U27041 (N_27041,N_24708,N_24164);
nand U27042 (N_27042,N_23433,N_23100);
and U27043 (N_27043,N_23655,N_23563);
xor U27044 (N_27044,N_24616,N_23223);
and U27045 (N_27045,N_22985,N_23597);
xnor U27046 (N_27046,N_24905,N_22995);
xor U27047 (N_27047,N_24290,N_23163);
or U27048 (N_27048,N_24045,N_23041);
or U27049 (N_27049,N_22856,N_23974);
nor U27050 (N_27050,N_24270,N_23460);
nand U27051 (N_27051,N_24151,N_23013);
xnor U27052 (N_27052,N_22910,N_22904);
nor U27053 (N_27053,N_23776,N_24767);
nand U27054 (N_27054,N_23700,N_22814);
nand U27055 (N_27055,N_23864,N_22504);
and U27056 (N_27056,N_24482,N_23016);
or U27057 (N_27057,N_24070,N_23822);
xnor U27058 (N_27058,N_23329,N_24673);
nor U27059 (N_27059,N_23943,N_23144);
nor U27060 (N_27060,N_23177,N_24039);
nor U27061 (N_27061,N_23337,N_23480);
nand U27062 (N_27062,N_22946,N_24365);
xnor U27063 (N_27063,N_23180,N_23486);
and U27064 (N_27064,N_23147,N_24786);
xnor U27065 (N_27065,N_24628,N_23998);
nor U27066 (N_27066,N_24944,N_24108);
nand U27067 (N_27067,N_24433,N_22826);
nor U27068 (N_27068,N_24766,N_24381);
xor U27069 (N_27069,N_22655,N_24051);
nor U27070 (N_27070,N_23584,N_23920);
or U27071 (N_27071,N_24831,N_23539);
and U27072 (N_27072,N_24671,N_23675);
nand U27073 (N_27073,N_24346,N_23032);
nand U27074 (N_27074,N_24925,N_24309);
xor U27075 (N_27075,N_23794,N_24575);
or U27076 (N_27076,N_22752,N_23908);
nor U27077 (N_27077,N_23055,N_22549);
xnor U27078 (N_27078,N_24466,N_24994);
and U27079 (N_27079,N_24248,N_23007);
nor U27080 (N_27080,N_24782,N_23766);
and U27081 (N_27081,N_24224,N_23125);
nor U27082 (N_27082,N_23940,N_24399);
nor U27083 (N_27083,N_24136,N_24828);
xor U27084 (N_27084,N_22957,N_23868);
or U27085 (N_27085,N_23968,N_23233);
xnor U27086 (N_27086,N_23250,N_23915);
nor U27087 (N_27087,N_24749,N_22962);
nor U27088 (N_27088,N_23513,N_22628);
xnor U27089 (N_27089,N_24031,N_22868);
nand U27090 (N_27090,N_23591,N_24195);
xnor U27091 (N_27091,N_22920,N_22963);
nand U27092 (N_27092,N_24568,N_24343);
and U27093 (N_27093,N_24289,N_24158);
nand U27094 (N_27094,N_24855,N_22846);
xor U27095 (N_27095,N_24765,N_23159);
nor U27096 (N_27096,N_23828,N_22840);
xor U27097 (N_27097,N_24054,N_22533);
nand U27098 (N_27098,N_24194,N_22539);
or U27099 (N_27099,N_23141,N_24998);
nand U27100 (N_27100,N_22750,N_23655);
xor U27101 (N_27101,N_23668,N_22888);
nand U27102 (N_27102,N_24223,N_23922);
xor U27103 (N_27103,N_24253,N_24846);
and U27104 (N_27104,N_22604,N_22707);
or U27105 (N_27105,N_23424,N_22631);
nor U27106 (N_27106,N_23549,N_24969);
xnor U27107 (N_27107,N_22500,N_22767);
nor U27108 (N_27108,N_24932,N_23224);
and U27109 (N_27109,N_22537,N_23129);
and U27110 (N_27110,N_23429,N_22951);
or U27111 (N_27111,N_24631,N_22987);
nor U27112 (N_27112,N_24624,N_23401);
xnor U27113 (N_27113,N_24810,N_22735);
xor U27114 (N_27114,N_24147,N_23901);
nand U27115 (N_27115,N_23278,N_23100);
and U27116 (N_27116,N_24889,N_23647);
xnor U27117 (N_27117,N_22587,N_24054);
or U27118 (N_27118,N_24703,N_22708);
xor U27119 (N_27119,N_23315,N_22854);
nand U27120 (N_27120,N_22992,N_22864);
or U27121 (N_27121,N_23981,N_24727);
or U27122 (N_27122,N_24484,N_23201);
and U27123 (N_27123,N_22895,N_24855);
or U27124 (N_27124,N_23004,N_23658);
nor U27125 (N_27125,N_24874,N_24108);
xor U27126 (N_27126,N_24933,N_24413);
and U27127 (N_27127,N_24202,N_24243);
or U27128 (N_27128,N_23465,N_23835);
or U27129 (N_27129,N_22597,N_23759);
nor U27130 (N_27130,N_23425,N_23631);
nor U27131 (N_27131,N_24098,N_24882);
nand U27132 (N_27132,N_23735,N_24655);
xor U27133 (N_27133,N_24667,N_24241);
nand U27134 (N_27134,N_24409,N_24178);
and U27135 (N_27135,N_24922,N_22869);
or U27136 (N_27136,N_24258,N_22504);
nor U27137 (N_27137,N_24773,N_24992);
xnor U27138 (N_27138,N_23423,N_23127);
xor U27139 (N_27139,N_24469,N_23413);
or U27140 (N_27140,N_24220,N_24703);
nand U27141 (N_27141,N_24974,N_23908);
nand U27142 (N_27142,N_22781,N_22807);
nand U27143 (N_27143,N_23880,N_23454);
nand U27144 (N_27144,N_24628,N_24598);
xnor U27145 (N_27145,N_23574,N_22737);
nor U27146 (N_27146,N_23439,N_24537);
xnor U27147 (N_27147,N_23814,N_24563);
or U27148 (N_27148,N_22501,N_24454);
and U27149 (N_27149,N_23873,N_22613);
xnor U27150 (N_27150,N_24301,N_24794);
nand U27151 (N_27151,N_24077,N_24265);
or U27152 (N_27152,N_22849,N_23648);
and U27153 (N_27153,N_24082,N_24991);
nor U27154 (N_27154,N_22754,N_23371);
nand U27155 (N_27155,N_23308,N_23922);
nor U27156 (N_27156,N_23008,N_24687);
nor U27157 (N_27157,N_24812,N_23725);
xor U27158 (N_27158,N_23914,N_24834);
or U27159 (N_27159,N_23249,N_24311);
xnor U27160 (N_27160,N_23691,N_22863);
xnor U27161 (N_27161,N_23026,N_22872);
xor U27162 (N_27162,N_22899,N_23410);
nand U27163 (N_27163,N_22821,N_24608);
nor U27164 (N_27164,N_24465,N_23558);
or U27165 (N_27165,N_24110,N_24256);
nor U27166 (N_27166,N_23426,N_23361);
or U27167 (N_27167,N_24544,N_23690);
or U27168 (N_27168,N_23596,N_23200);
nand U27169 (N_27169,N_23297,N_23181);
or U27170 (N_27170,N_23779,N_24540);
or U27171 (N_27171,N_23902,N_24890);
nand U27172 (N_27172,N_22992,N_23369);
xor U27173 (N_27173,N_24398,N_23161);
xor U27174 (N_27174,N_23517,N_23013);
nor U27175 (N_27175,N_22666,N_24790);
nor U27176 (N_27176,N_24108,N_23011);
nand U27177 (N_27177,N_24993,N_23847);
and U27178 (N_27178,N_22972,N_23394);
xnor U27179 (N_27179,N_24979,N_23810);
nand U27180 (N_27180,N_24217,N_23256);
or U27181 (N_27181,N_23782,N_24753);
and U27182 (N_27182,N_23861,N_22658);
xnor U27183 (N_27183,N_22907,N_22931);
xnor U27184 (N_27184,N_23236,N_23515);
and U27185 (N_27185,N_24403,N_23021);
or U27186 (N_27186,N_24376,N_24552);
and U27187 (N_27187,N_24240,N_23272);
and U27188 (N_27188,N_23678,N_23832);
nor U27189 (N_27189,N_23154,N_22904);
nor U27190 (N_27190,N_23303,N_22572);
and U27191 (N_27191,N_23282,N_23161);
xnor U27192 (N_27192,N_24466,N_22757);
nor U27193 (N_27193,N_23124,N_22582);
or U27194 (N_27194,N_23105,N_23024);
nor U27195 (N_27195,N_24520,N_22537);
xor U27196 (N_27196,N_22748,N_24904);
or U27197 (N_27197,N_23022,N_24352);
nor U27198 (N_27198,N_24134,N_23676);
xor U27199 (N_27199,N_22568,N_24297);
nor U27200 (N_27200,N_23328,N_23071);
and U27201 (N_27201,N_24230,N_23704);
or U27202 (N_27202,N_23959,N_23657);
or U27203 (N_27203,N_23640,N_23726);
and U27204 (N_27204,N_24604,N_23635);
xor U27205 (N_27205,N_23802,N_22987);
or U27206 (N_27206,N_23719,N_23735);
or U27207 (N_27207,N_22720,N_22852);
and U27208 (N_27208,N_22956,N_23486);
nor U27209 (N_27209,N_24738,N_24976);
nand U27210 (N_27210,N_22566,N_24523);
nand U27211 (N_27211,N_23715,N_23647);
or U27212 (N_27212,N_24555,N_23173);
nor U27213 (N_27213,N_23422,N_23888);
nor U27214 (N_27214,N_23407,N_22960);
nand U27215 (N_27215,N_24127,N_22731);
nand U27216 (N_27216,N_23318,N_24839);
and U27217 (N_27217,N_23586,N_23029);
and U27218 (N_27218,N_23395,N_22971);
nand U27219 (N_27219,N_24290,N_23033);
nor U27220 (N_27220,N_23136,N_23508);
nand U27221 (N_27221,N_24648,N_22650);
xnor U27222 (N_27222,N_24321,N_22960);
and U27223 (N_27223,N_22944,N_23513);
and U27224 (N_27224,N_24862,N_22663);
nand U27225 (N_27225,N_23561,N_23944);
and U27226 (N_27226,N_22922,N_22618);
nor U27227 (N_27227,N_24408,N_23406);
and U27228 (N_27228,N_24174,N_22834);
nand U27229 (N_27229,N_24640,N_24777);
and U27230 (N_27230,N_23977,N_23314);
xor U27231 (N_27231,N_24974,N_22829);
xnor U27232 (N_27232,N_24662,N_23258);
xnor U27233 (N_27233,N_24244,N_24101);
or U27234 (N_27234,N_23095,N_22741);
xor U27235 (N_27235,N_24885,N_24341);
nor U27236 (N_27236,N_23803,N_22562);
xor U27237 (N_27237,N_24781,N_24059);
xor U27238 (N_27238,N_23006,N_24399);
nand U27239 (N_27239,N_22657,N_24431);
xnor U27240 (N_27240,N_23756,N_22815);
nor U27241 (N_27241,N_24246,N_22640);
xor U27242 (N_27242,N_22735,N_23334);
and U27243 (N_27243,N_22865,N_23920);
nor U27244 (N_27244,N_23227,N_24204);
or U27245 (N_27245,N_24668,N_23397);
nand U27246 (N_27246,N_22579,N_22563);
nor U27247 (N_27247,N_24821,N_22878);
nand U27248 (N_27248,N_22965,N_22660);
and U27249 (N_27249,N_24335,N_23109);
nand U27250 (N_27250,N_23488,N_24655);
nand U27251 (N_27251,N_23960,N_23902);
and U27252 (N_27252,N_24169,N_24493);
and U27253 (N_27253,N_23656,N_24407);
and U27254 (N_27254,N_24564,N_23405);
and U27255 (N_27255,N_23473,N_24955);
or U27256 (N_27256,N_23046,N_23188);
and U27257 (N_27257,N_24454,N_22713);
nor U27258 (N_27258,N_24420,N_22606);
nand U27259 (N_27259,N_23115,N_22615);
nor U27260 (N_27260,N_24607,N_24198);
nor U27261 (N_27261,N_23267,N_24423);
xor U27262 (N_27262,N_23640,N_24746);
nor U27263 (N_27263,N_24730,N_24575);
nor U27264 (N_27264,N_24938,N_22684);
and U27265 (N_27265,N_23201,N_24686);
or U27266 (N_27266,N_24965,N_24654);
or U27267 (N_27267,N_22558,N_24890);
or U27268 (N_27268,N_24699,N_24055);
or U27269 (N_27269,N_23710,N_23284);
or U27270 (N_27270,N_24095,N_24661);
or U27271 (N_27271,N_23586,N_23669);
nor U27272 (N_27272,N_24357,N_23676);
nor U27273 (N_27273,N_23525,N_24219);
xor U27274 (N_27274,N_22539,N_24987);
or U27275 (N_27275,N_23044,N_24152);
nor U27276 (N_27276,N_24929,N_24776);
nand U27277 (N_27277,N_23457,N_24226);
nand U27278 (N_27278,N_23930,N_24382);
xor U27279 (N_27279,N_22980,N_24780);
or U27280 (N_27280,N_22904,N_23583);
nand U27281 (N_27281,N_23645,N_23303);
nor U27282 (N_27282,N_24817,N_22552);
or U27283 (N_27283,N_23126,N_23787);
or U27284 (N_27284,N_24914,N_23473);
nand U27285 (N_27285,N_23910,N_24149);
and U27286 (N_27286,N_22842,N_24997);
nor U27287 (N_27287,N_22706,N_23151);
nand U27288 (N_27288,N_24422,N_22597);
or U27289 (N_27289,N_24488,N_24749);
xor U27290 (N_27290,N_22697,N_22708);
nand U27291 (N_27291,N_22952,N_24803);
nor U27292 (N_27292,N_23340,N_24353);
nor U27293 (N_27293,N_23328,N_22857);
nor U27294 (N_27294,N_24495,N_22816);
and U27295 (N_27295,N_24996,N_23339);
and U27296 (N_27296,N_22713,N_23700);
or U27297 (N_27297,N_23676,N_23178);
and U27298 (N_27298,N_23784,N_24850);
or U27299 (N_27299,N_23332,N_23881);
nor U27300 (N_27300,N_24671,N_23456);
xor U27301 (N_27301,N_24909,N_23534);
or U27302 (N_27302,N_24918,N_24934);
or U27303 (N_27303,N_22951,N_24826);
or U27304 (N_27304,N_23219,N_23899);
nand U27305 (N_27305,N_24724,N_23451);
and U27306 (N_27306,N_23704,N_23612);
nand U27307 (N_27307,N_23271,N_23460);
xnor U27308 (N_27308,N_22570,N_24453);
and U27309 (N_27309,N_24589,N_23334);
or U27310 (N_27310,N_24410,N_24995);
nor U27311 (N_27311,N_24098,N_23767);
and U27312 (N_27312,N_22949,N_23216);
nor U27313 (N_27313,N_24045,N_24991);
nand U27314 (N_27314,N_24942,N_24614);
nand U27315 (N_27315,N_23096,N_24469);
nand U27316 (N_27316,N_23529,N_24670);
or U27317 (N_27317,N_23521,N_23144);
nand U27318 (N_27318,N_23263,N_23423);
nand U27319 (N_27319,N_22579,N_24017);
xor U27320 (N_27320,N_24621,N_24288);
or U27321 (N_27321,N_22864,N_23750);
nand U27322 (N_27322,N_23084,N_24467);
or U27323 (N_27323,N_24568,N_23899);
nand U27324 (N_27324,N_23230,N_23575);
nand U27325 (N_27325,N_24049,N_23141);
xnor U27326 (N_27326,N_23815,N_23746);
and U27327 (N_27327,N_24344,N_23669);
and U27328 (N_27328,N_24051,N_22840);
or U27329 (N_27329,N_23559,N_22525);
nand U27330 (N_27330,N_24097,N_23391);
xnor U27331 (N_27331,N_23452,N_23959);
nor U27332 (N_27332,N_23605,N_24448);
nor U27333 (N_27333,N_24614,N_24501);
and U27334 (N_27334,N_24825,N_22949);
and U27335 (N_27335,N_24403,N_24636);
nor U27336 (N_27336,N_23340,N_23349);
or U27337 (N_27337,N_23901,N_22696);
nand U27338 (N_27338,N_23254,N_23776);
nor U27339 (N_27339,N_24678,N_23659);
nor U27340 (N_27340,N_22795,N_22882);
and U27341 (N_27341,N_23171,N_23195);
xnor U27342 (N_27342,N_24422,N_22652);
nor U27343 (N_27343,N_22593,N_24072);
xor U27344 (N_27344,N_23219,N_23083);
xnor U27345 (N_27345,N_24204,N_22755);
xor U27346 (N_27346,N_24430,N_23018);
nand U27347 (N_27347,N_24683,N_23151);
nor U27348 (N_27348,N_24634,N_24100);
nor U27349 (N_27349,N_22676,N_24628);
xor U27350 (N_27350,N_23320,N_22909);
and U27351 (N_27351,N_24930,N_24444);
nand U27352 (N_27352,N_24747,N_24180);
xnor U27353 (N_27353,N_24154,N_24926);
nor U27354 (N_27354,N_22995,N_24738);
nand U27355 (N_27355,N_24033,N_23401);
xor U27356 (N_27356,N_23653,N_23255);
and U27357 (N_27357,N_23448,N_23803);
and U27358 (N_27358,N_23579,N_24563);
or U27359 (N_27359,N_22730,N_24559);
nand U27360 (N_27360,N_23297,N_23228);
or U27361 (N_27361,N_23402,N_23127);
or U27362 (N_27362,N_24675,N_23353);
and U27363 (N_27363,N_24371,N_24582);
nand U27364 (N_27364,N_24595,N_22974);
nor U27365 (N_27365,N_23882,N_23900);
nor U27366 (N_27366,N_24112,N_24600);
xnor U27367 (N_27367,N_24196,N_24491);
or U27368 (N_27368,N_23862,N_24173);
or U27369 (N_27369,N_24526,N_24103);
nand U27370 (N_27370,N_23695,N_24125);
and U27371 (N_27371,N_23707,N_23809);
nand U27372 (N_27372,N_23787,N_24950);
or U27373 (N_27373,N_24094,N_22967);
nor U27374 (N_27374,N_23335,N_23026);
nor U27375 (N_27375,N_22809,N_23743);
or U27376 (N_27376,N_23318,N_23228);
nor U27377 (N_27377,N_23712,N_23643);
nand U27378 (N_27378,N_24429,N_22578);
and U27379 (N_27379,N_24146,N_24935);
nor U27380 (N_27380,N_24444,N_22737);
xnor U27381 (N_27381,N_23729,N_22936);
xor U27382 (N_27382,N_23591,N_23175);
or U27383 (N_27383,N_24622,N_24235);
or U27384 (N_27384,N_23990,N_23082);
xor U27385 (N_27385,N_22755,N_23395);
and U27386 (N_27386,N_22599,N_23587);
nand U27387 (N_27387,N_23443,N_24612);
xnor U27388 (N_27388,N_22817,N_23001);
xnor U27389 (N_27389,N_24874,N_23562);
or U27390 (N_27390,N_22915,N_24742);
or U27391 (N_27391,N_24638,N_23869);
and U27392 (N_27392,N_23735,N_23248);
xnor U27393 (N_27393,N_24037,N_24601);
or U27394 (N_27394,N_24003,N_24166);
nand U27395 (N_27395,N_23810,N_22597);
nand U27396 (N_27396,N_23588,N_23438);
or U27397 (N_27397,N_23414,N_22963);
xnor U27398 (N_27398,N_22663,N_23150);
nand U27399 (N_27399,N_23404,N_24788);
and U27400 (N_27400,N_24417,N_24576);
or U27401 (N_27401,N_24864,N_23042);
nand U27402 (N_27402,N_23920,N_24954);
nand U27403 (N_27403,N_24159,N_24418);
and U27404 (N_27404,N_24683,N_23594);
nand U27405 (N_27405,N_22727,N_22818);
xnor U27406 (N_27406,N_24383,N_22619);
nor U27407 (N_27407,N_23831,N_23750);
nand U27408 (N_27408,N_23654,N_23955);
nor U27409 (N_27409,N_24780,N_22668);
nand U27410 (N_27410,N_24675,N_23285);
and U27411 (N_27411,N_24113,N_24758);
and U27412 (N_27412,N_23607,N_23068);
xnor U27413 (N_27413,N_22753,N_22515);
xor U27414 (N_27414,N_22888,N_24038);
nand U27415 (N_27415,N_22747,N_23673);
xnor U27416 (N_27416,N_24961,N_24650);
nor U27417 (N_27417,N_22824,N_24552);
or U27418 (N_27418,N_23210,N_22961);
and U27419 (N_27419,N_24680,N_24377);
nand U27420 (N_27420,N_24835,N_22631);
nor U27421 (N_27421,N_24481,N_23045);
nor U27422 (N_27422,N_22587,N_23941);
and U27423 (N_27423,N_24235,N_22508);
xnor U27424 (N_27424,N_23350,N_24744);
or U27425 (N_27425,N_23116,N_23921);
xor U27426 (N_27426,N_24718,N_24170);
nor U27427 (N_27427,N_22958,N_24586);
and U27428 (N_27428,N_24028,N_23909);
xnor U27429 (N_27429,N_24115,N_24654);
or U27430 (N_27430,N_22855,N_24702);
xor U27431 (N_27431,N_24957,N_24017);
nor U27432 (N_27432,N_24453,N_23137);
nor U27433 (N_27433,N_23825,N_24852);
and U27434 (N_27434,N_24942,N_24781);
and U27435 (N_27435,N_23671,N_23647);
and U27436 (N_27436,N_22964,N_23192);
or U27437 (N_27437,N_23046,N_22718);
nor U27438 (N_27438,N_23366,N_23037);
xnor U27439 (N_27439,N_22662,N_23418);
xor U27440 (N_27440,N_23946,N_24607);
xor U27441 (N_27441,N_23143,N_24063);
or U27442 (N_27442,N_24997,N_23583);
xnor U27443 (N_27443,N_23549,N_24766);
xnor U27444 (N_27444,N_23513,N_22878);
and U27445 (N_27445,N_23097,N_23799);
nand U27446 (N_27446,N_23974,N_23622);
or U27447 (N_27447,N_24947,N_23200);
or U27448 (N_27448,N_23963,N_24004);
nor U27449 (N_27449,N_22684,N_23197);
xor U27450 (N_27450,N_24959,N_23398);
or U27451 (N_27451,N_23234,N_22932);
nor U27452 (N_27452,N_22688,N_24732);
and U27453 (N_27453,N_23759,N_23324);
and U27454 (N_27454,N_23746,N_23139);
nor U27455 (N_27455,N_24151,N_23592);
nand U27456 (N_27456,N_22582,N_23809);
or U27457 (N_27457,N_24272,N_24584);
nor U27458 (N_27458,N_23203,N_23833);
nand U27459 (N_27459,N_23210,N_22769);
xor U27460 (N_27460,N_23019,N_24062);
and U27461 (N_27461,N_22711,N_23604);
or U27462 (N_27462,N_24794,N_23379);
and U27463 (N_27463,N_23678,N_23681);
nor U27464 (N_27464,N_24807,N_23774);
xor U27465 (N_27465,N_23145,N_23160);
and U27466 (N_27466,N_22526,N_23631);
xor U27467 (N_27467,N_23390,N_22970);
nor U27468 (N_27468,N_23664,N_22623);
or U27469 (N_27469,N_24178,N_23419);
xnor U27470 (N_27470,N_23879,N_24021);
or U27471 (N_27471,N_22601,N_22652);
xnor U27472 (N_27472,N_24869,N_22783);
xor U27473 (N_27473,N_23453,N_24918);
and U27474 (N_27474,N_24057,N_23582);
or U27475 (N_27475,N_23526,N_23064);
and U27476 (N_27476,N_23602,N_23031);
and U27477 (N_27477,N_22895,N_24750);
xnor U27478 (N_27478,N_23201,N_23383);
nand U27479 (N_27479,N_22666,N_23962);
xor U27480 (N_27480,N_24053,N_23363);
or U27481 (N_27481,N_22671,N_23205);
nand U27482 (N_27482,N_22937,N_23821);
xor U27483 (N_27483,N_23088,N_23757);
xnor U27484 (N_27484,N_22769,N_23559);
nand U27485 (N_27485,N_23242,N_24650);
and U27486 (N_27486,N_24535,N_23168);
nand U27487 (N_27487,N_22666,N_23714);
nor U27488 (N_27488,N_23754,N_24443);
nand U27489 (N_27489,N_22933,N_24888);
nand U27490 (N_27490,N_22863,N_22520);
xnor U27491 (N_27491,N_24838,N_23445);
and U27492 (N_27492,N_24902,N_23817);
and U27493 (N_27493,N_24123,N_23062);
or U27494 (N_27494,N_24925,N_24901);
xor U27495 (N_27495,N_24875,N_23895);
xor U27496 (N_27496,N_23397,N_24401);
xor U27497 (N_27497,N_23534,N_24129);
nand U27498 (N_27498,N_23020,N_24516);
xnor U27499 (N_27499,N_22570,N_23499);
nand U27500 (N_27500,N_25852,N_25856);
nand U27501 (N_27501,N_26412,N_25502);
and U27502 (N_27502,N_26908,N_27286);
nor U27503 (N_27503,N_27427,N_26974);
nand U27504 (N_27504,N_26151,N_26738);
and U27505 (N_27505,N_26785,N_26773);
nor U27506 (N_27506,N_27225,N_26178);
nor U27507 (N_27507,N_26382,N_26887);
nor U27508 (N_27508,N_25529,N_25698);
xor U27509 (N_27509,N_25935,N_27245);
and U27510 (N_27510,N_26111,N_27033);
and U27511 (N_27511,N_25289,N_26112);
and U27512 (N_27512,N_25052,N_26638);
or U27513 (N_27513,N_27470,N_25549);
xnor U27514 (N_27514,N_27422,N_26371);
nand U27515 (N_27515,N_25039,N_26649);
nand U27516 (N_27516,N_26374,N_25714);
or U27517 (N_27517,N_27122,N_25636);
or U27518 (N_27518,N_26637,N_26142);
and U27519 (N_27519,N_27175,N_26916);
xnor U27520 (N_27520,N_25304,N_25813);
or U27521 (N_27521,N_26500,N_26018);
nor U27522 (N_27522,N_26823,N_25885);
xor U27523 (N_27523,N_26107,N_25035);
nand U27524 (N_27524,N_27359,N_26568);
and U27525 (N_27525,N_25803,N_25620);
nand U27526 (N_27526,N_26671,N_25559);
nand U27527 (N_27527,N_25306,N_26566);
or U27528 (N_27528,N_25275,N_25458);
or U27529 (N_27529,N_25783,N_26700);
xnor U27530 (N_27530,N_25579,N_26059);
nor U27531 (N_27531,N_27307,N_27370);
nor U27532 (N_27532,N_26460,N_26850);
and U27533 (N_27533,N_25341,N_25878);
xnor U27534 (N_27534,N_25122,N_27116);
and U27535 (N_27535,N_25450,N_27143);
or U27536 (N_27536,N_27151,N_27378);
nand U27537 (N_27537,N_25524,N_26524);
and U27538 (N_27538,N_25354,N_25821);
nor U27539 (N_27539,N_25745,N_26867);
and U27540 (N_27540,N_27062,N_25733);
nand U27541 (N_27541,N_26354,N_26222);
nor U27542 (N_27542,N_25608,N_25105);
nor U27543 (N_27543,N_26701,N_25888);
or U27544 (N_27544,N_27227,N_25463);
and U27545 (N_27545,N_26716,N_27110);
or U27546 (N_27546,N_25682,N_26387);
xnor U27547 (N_27547,N_26602,N_25180);
and U27548 (N_27548,N_26323,N_26426);
xnor U27549 (N_27549,N_26596,N_26648);
nor U27550 (N_27550,N_25164,N_26183);
nand U27551 (N_27551,N_27156,N_26318);
or U27552 (N_27552,N_25941,N_26960);
or U27553 (N_27553,N_27094,N_25490);
or U27554 (N_27554,N_25124,N_27445);
xor U27555 (N_27555,N_27018,N_25240);
xor U27556 (N_27556,N_27403,N_26032);
nor U27557 (N_27557,N_25276,N_27322);
nor U27558 (N_27558,N_26001,N_26084);
nand U27559 (N_27559,N_27252,N_26975);
or U27560 (N_27560,N_25368,N_26071);
or U27561 (N_27561,N_25247,N_25446);
nor U27562 (N_27562,N_26155,N_27390);
and U27563 (N_27563,N_26834,N_26761);
nor U27564 (N_27564,N_27148,N_26582);
xnor U27565 (N_27565,N_25238,N_27329);
or U27566 (N_27566,N_26856,N_26606);
or U27567 (N_27567,N_25233,N_26280);
or U27568 (N_27568,N_26527,N_26288);
nor U27569 (N_27569,N_25989,N_27406);
xor U27570 (N_27570,N_27089,N_27379);
or U27571 (N_27571,N_26368,N_26999);
xnor U27572 (N_27572,N_26099,N_26423);
nor U27573 (N_27573,N_26874,N_26547);
nand U27574 (N_27574,N_26829,N_25471);
xnor U27575 (N_27575,N_25789,N_27028);
and U27576 (N_27576,N_27185,N_25319);
or U27577 (N_27577,N_26956,N_27004);
or U27578 (N_27578,N_25717,N_25676);
or U27579 (N_27579,N_25861,N_25774);
xnor U27580 (N_27580,N_25205,N_26242);
and U27581 (N_27581,N_27292,N_27120);
nand U27582 (N_27582,N_27298,N_25936);
nor U27583 (N_27583,N_25815,N_26519);
and U27584 (N_27584,N_25970,N_27451);
xnor U27585 (N_27585,N_25896,N_25484);
xnor U27586 (N_27586,N_25506,N_25401);
and U27587 (N_27587,N_25903,N_26505);
nor U27588 (N_27588,N_27366,N_25080);
and U27589 (N_27589,N_26977,N_26234);
nor U27590 (N_27590,N_27396,N_26133);
and U27591 (N_27591,N_26381,N_26724);
and U27592 (N_27592,N_25499,N_25396);
and U27593 (N_27593,N_27358,N_26255);
and U27594 (N_27594,N_27325,N_25414);
nor U27595 (N_27595,N_27141,N_25239);
nor U27596 (N_27596,N_25925,N_25601);
nand U27597 (N_27597,N_25104,N_26243);
or U27598 (N_27598,N_26838,N_26082);
nor U27599 (N_27599,N_25175,N_25792);
nor U27600 (N_27600,N_26055,N_26418);
nand U27601 (N_27601,N_25027,N_26160);
xnor U27602 (N_27602,N_26231,N_27069);
xor U27603 (N_27603,N_25103,N_27481);
xnor U27604 (N_27604,N_25556,N_26942);
nor U27605 (N_27605,N_26275,N_26149);
nor U27606 (N_27606,N_27401,N_26410);
xor U27607 (N_27607,N_25706,N_26427);
nor U27608 (N_27608,N_27263,N_25918);
and U27609 (N_27609,N_27165,N_26129);
and U27610 (N_27610,N_25822,N_25966);
nor U27611 (N_27611,N_27454,N_27385);
and U27612 (N_27612,N_27248,N_25436);
nand U27613 (N_27613,N_27027,N_25974);
or U27614 (N_27614,N_26370,N_25649);
nand U27615 (N_27615,N_25864,N_26390);
and U27616 (N_27616,N_25668,N_25791);
and U27617 (N_27617,N_26168,N_25592);
and U27618 (N_27618,N_25426,N_27301);
or U27619 (N_27619,N_26109,N_25554);
xor U27620 (N_27620,N_26170,N_25063);
and U27621 (N_27621,N_26403,N_25320);
and U27622 (N_27622,N_26310,N_26186);
xnor U27623 (N_27623,N_26538,N_25500);
nor U27624 (N_27624,N_27186,N_25111);
or U27625 (N_27625,N_26817,N_26904);
nand U27626 (N_27626,N_25527,N_25470);
and U27627 (N_27627,N_26517,N_25981);
nand U27628 (N_27628,N_25193,N_26120);
xor U27629 (N_27629,N_26575,N_26025);
nor U27630 (N_27630,N_26080,N_26273);
and U27631 (N_27631,N_27324,N_26430);
xor U27632 (N_27632,N_25190,N_27228);
nand U27633 (N_27633,N_27063,N_25539);
xor U27634 (N_27634,N_26585,N_26683);
nand U27635 (N_27635,N_25841,N_26348);
and U27636 (N_27636,N_27434,N_26413);
and U27637 (N_27637,N_25351,N_27169);
and U27638 (N_27638,N_26507,N_26910);
and U27639 (N_27639,N_26384,N_25750);
or U27640 (N_27640,N_26281,N_27467);
and U27641 (N_27641,N_27450,N_26973);
and U27642 (N_27642,N_25708,N_26366);
or U27643 (N_27643,N_27455,N_26475);
or U27644 (N_27644,N_25317,N_26534);
nor U27645 (N_27645,N_26420,N_27220);
nor U27646 (N_27646,N_27285,N_26639);
or U27647 (N_27647,N_27345,N_27281);
and U27648 (N_27648,N_26301,N_27187);
nand U27649 (N_27649,N_25646,N_25525);
nor U27650 (N_27650,N_25173,N_25727);
nand U27651 (N_27651,N_26576,N_26786);
xor U27652 (N_27652,N_26965,N_25011);
or U27653 (N_27653,N_26959,N_25267);
or U27654 (N_27654,N_26051,N_26136);
nand U27655 (N_27655,N_25514,N_26503);
nor U27656 (N_27656,N_27022,N_25732);
or U27657 (N_27657,N_25736,N_26611);
xor U27658 (N_27658,N_25263,N_26666);
and U27659 (N_27659,N_25623,N_26378);
xnor U27660 (N_27660,N_26035,N_25756);
nor U27661 (N_27661,N_25975,N_25906);
nor U27662 (N_27662,N_25101,N_27279);
nand U27663 (N_27663,N_25467,N_27420);
xnor U27664 (N_27664,N_26556,N_25921);
nor U27665 (N_27665,N_25369,N_26217);
nor U27666 (N_27666,N_27289,N_25560);
xor U27667 (N_27667,N_26802,N_25587);
or U27668 (N_27668,N_26809,N_26141);
or U27669 (N_27669,N_26140,N_27191);
and U27670 (N_27670,N_25285,N_27466);
nor U27671 (N_27671,N_26501,N_26165);
or U27672 (N_27672,N_27226,N_26912);
nor U27673 (N_27673,N_26945,N_25438);
and U27674 (N_27674,N_25187,N_26295);
or U27675 (N_27675,N_26755,N_25230);
nand U27676 (N_27676,N_27108,N_25007);
nor U27677 (N_27677,N_25749,N_27178);
or U27678 (N_27678,N_26157,N_25626);
nor U27679 (N_27679,N_25863,N_26261);
nor U27680 (N_27680,N_25225,N_26669);
nor U27681 (N_27681,N_25672,N_27476);
nand U27682 (N_27682,N_25911,N_25729);
nor U27683 (N_27683,N_25871,N_25115);
nand U27684 (N_27684,N_25360,N_26346);
xor U27685 (N_27685,N_27332,N_25330);
and U27686 (N_27686,N_25352,N_27121);
nor U27687 (N_27687,N_25015,N_26437);
and U27688 (N_27688,N_25421,N_25678);
nor U27689 (N_27689,N_25880,N_25066);
and U27690 (N_27690,N_25325,N_26890);
nand U27691 (N_27691,N_26735,N_25283);
nor U27692 (N_27692,N_25082,N_26008);
xnor U27693 (N_27693,N_25804,N_27180);
or U27694 (N_27694,N_26487,N_26610);
and U27695 (N_27695,N_26810,N_25472);
and U27696 (N_27696,N_25479,N_25023);
or U27697 (N_27697,N_25894,N_26961);
or U27698 (N_27698,N_25252,N_26282);
nand U27699 (N_27699,N_27200,N_27086);
xor U27700 (N_27700,N_26176,N_26642);
and U27701 (N_27701,N_26303,N_26340);
nor U27702 (N_27702,N_27229,N_26407);
xnor U27703 (N_27703,N_27419,N_26495);
nand U27704 (N_27704,N_25003,N_25146);
xnor U27705 (N_27705,N_25399,N_25533);
nand U27706 (N_27706,N_26546,N_26909);
nand U27707 (N_27707,N_26167,N_26074);
or U27708 (N_27708,N_27382,N_27354);
xnor U27709 (N_27709,N_25816,N_27374);
xor U27710 (N_27710,N_25215,N_26360);
or U27711 (N_27711,N_27269,N_26329);
xor U27712 (N_27712,N_25231,N_25221);
nor U27713 (N_27713,N_27368,N_27192);
xnor U27714 (N_27714,N_26774,N_27430);
nor U27715 (N_27715,N_25395,N_25223);
nor U27716 (N_27716,N_25168,N_26341);
nor U27717 (N_27717,N_25162,N_25688);
nor U27718 (N_27718,N_27312,N_27413);
xor U27719 (N_27719,N_27237,N_27243);
and U27720 (N_27720,N_27458,N_26251);
and U27721 (N_27721,N_25144,N_26296);
or U27722 (N_27722,N_25327,N_25140);
xor U27723 (N_27723,N_26298,N_26190);
or U27724 (N_27724,N_27314,N_26383);
and U27725 (N_27725,N_25488,N_25602);
or U27726 (N_27726,N_27397,N_26322);
or U27727 (N_27727,N_27235,N_26088);
nand U27728 (N_27728,N_25632,N_27495);
or U27729 (N_27729,N_27162,N_25843);
nand U27730 (N_27730,N_25228,N_25345);
nand U27731 (N_27731,N_25652,N_26240);
xor U27732 (N_27732,N_25990,N_27473);
and U27733 (N_27733,N_27484,N_26249);
nand U27734 (N_27734,N_25161,N_25687);
and U27735 (N_27735,N_26828,N_25110);
nand U27736 (N_27736,N_25107,N_26202);
nand U27737 (N_27737,N_26164,N_25847);
and U27738 (N_27738,N_25637,N_26122);
nor U27739 (N_27739,N_26808,N_25674);
nor U27740 (N_27740,N_25301,N_26499);
xnor U27741 (N_27741,N_25788,N_26731);
or U27742 (N_27742,N_25967,N_27124);
and U27743 (N_27743,N_26653,N_26210);
nor U27744 (N_27744,N_27318,N_25814);
or U27745 (N_27745,N_27246,N_25895);
xnor U27746 (N_27746,N_25834,N_27215);
nor U27747 (N_27747,N_25157,N_27111);
xor U27748 (N_27748,N_25435,N_26715);
xnor U27749 (N_27749,N_27347,N_26045);
nor U27750 (N_27750,N_26416,N_27060);
xor U27751 (N_27751,N_26599,N_25286);
nor U27752 (N_27752,N_26570,N_26897);
xnor U27753 (N_27753,N_25313,N_27303);
nand U27754 (N_27754,N_25246,N_25884);
nor U27755 (N_27755,N_25070,N_25242);
nor U27756 (N_27756,N_25516,N_27153);
and U27757 (N_27757,N_27115,N_26078);
or U27758 (N_27758,N_25937,N_26705);
or U27759 (N_27759,N_25483,N_27188);
and U27760 (N_27760,N_27030,N_26652);
or U27761 (N_27761,N_25326,N_25389);
nor U27762 (N_27762,N_27166,N_25163);
nand U27763 (N_27763,N_26733,N_26698);
xnor U27764 (N_27764,N_25938,N_27440);
or U27765 (N_27765,N_26866,N_25358);
and U27766 (N_27766,N_26748,N_26336);
xnor U27767 (N_27767,N_26727,N_26893);
nor U27768 (N_27768,N_25184,N_27049);
nor U27769 (N_27769,N_27230,N_25808);
nor U27770 (N_27770,N_26692,N_25314);
nor U27771 (N_27771,N_25734,N_25604);
nor U27772 (N_27772,N_26284,N_26935);
xnor U27773 (N_27773,N_25139,N_27136);
nand U27774 (N_27774,N_25372,N_25202);
or U27775 (N_27775,N_25462,N_27411);
nor U27776 (N_27776,N_27483,N_25532);
nor U27777 (N_27777,N_26860,N_25060);
xor U27778 (N_27778,N_26830,N_27276);
and U27779 (N_27779,N_26597,N_26216);
nor U27780 (N_27780,N_26446,N_25630);
nand U27781 (N_27781,N_26473,N_26472);
and U27782 (N_27782,N_26937,N_25445);
or U27783 (N_27783,N_25848,N_26220);
xnor U27784 (N_27784,N_25405,N_26214);
nand U27785 (N_27785,N_27485,N_26797);
nand U27786 (N_27786,N_26532,N_27195);
and U27787 (N_27787,N_25192,N_26985);
nand U27788 (N_27788,N_25645,N_26299);
and U27789 (N_27789,N_25511,N_25819);
nand U27790 (N_27790,N_25618,N_26722);
nand U27791 (N_27791,N_26837,N_26425);
nand U27792 (N_27792,N_26957,N_25662);
and U27793 (N_27793,N_25159,N_26745);
xnor U27794 (N_27794,N_26219,N_25826);
xnor U27795 (N_27795,N_25947,N_27438);
nand U27796 (N_27796,N_26414,N_26392);
or U27797 (N_27797,N_27134,N_26225);
and U27798 (N_27798,N_26728,N_25014);
nand U27799 (N_27799,N_26496,N_26911);
xor U27800 (N_27800,N_26144,N_25866);
nor U27801 (N_27801,N_25628,N_26889);
xnor U27802 (N_27802,N_25901,N_26247);
nor U27803 (N_27803,N_25174,N_25831);
or U27804 (N_27804,N_25795,N_26087);
nor U27805 (N_27805,N_25984,N_26946);
nor U27806 (N_27806,N_25065,N_25868);
nor U27807 (N_27807,N_26337,N_25128);
or U27808 (N_27808,N_27418,N_25555);
xnor U27809 (N_27809,N_25547,N_25218);
nor U27810 (N_27810,N_25050,N_25125);
xor U27811 (N_27811,N_27017,N_25069);
and U27812 (N_27812,N_26976,N_26094);
xor U27813 (N_27813,N_25042,N_25134);
nor U27814 (N_27814,N_26030,N_26763);
or U27815 (N_27815,N_27071,N_26949);
xor U27816 (N_27816,N_25116,N_26840);
nand U27817 (N_27817,N_25933,N_26885);
or U27818 (N_27818,N_26269,N_25631);
or U27819 (N_27819,N_26987,N_26300);
nand U27820 (N_27820,N_25338,N_25810);
or U27821 (N_27821,N_26806,N_26708);
or U27822 (N_27822,N_26609,N_25659);
or U27823 (N_27823,N_26581,N_26017);
nand U27824 (N_27824,N_27216,N_26940);
and U27825 (N_27825,N_26293,N_26042);
nand U27826 (N_27826,N_27005,N_26654);
nor U27827 (N_27827,N_26743,N_26053);
nand U27828 (N_27828,N_25558,N_25725);
nor U27829 (N_27829,N_26833,N_27428);
xor U27830 (N_27830,N_25030,N_26022);
xnor U27831 (N_27831,N_26510,N_26864);
nand U27832 (N_27832,N_26695,N_26297);
xnor U27833 (N_27833,N_27497,N_25366);
nor U27834 (N_27834,N_27061,N_25748);
nand U27835 (N_27835,N_26097,N_26043);
xor U27836 (N_27836,N_27321,N_25318);
xor U27837 (N_27837,N_26702,N_25546);
xnor U27838 (N_27838,N_26574,N_25764);
and U27839 (N_27839,N_27241,N_26616);
nand U27840 (N_27840,N_27369,N_26402);
and U27841 (N_27841,N_26233,N_26213);
nor U27842 (N_27842,N_27362,N_27257);
nor U27843 (N_27843,N_25158,N_25609);
xnor U27844 (N_27844,N_26464,N_25759);
xor U27845 (N_27845,N_25208,N_25026);
nor U27846 (N_27846,N_25206,N_25518);
nand U27847 (N_27847,N_25009,N_27492);
nor U27848 (N_27848,N_25695,N_26302);
nand U27849 (N_27849,N_25403,N_27078);
nor U27850 (N_27850,N_25566,N_25054);
nor U27851 (N_27851,N_27389,N_26955);
nor U27852 (N_27852,N_27337,N_25927);
nand U27853 (N_27853,N_26205,N_25942);
nand U27854 (N_27854,N_27057,N_27488);
and U27855 (N_27855,N_25417,N_25295);
nor U27856 (N_27856,N_27471,N_27144);
xor U27857 (N_27857,N_25016,N_26057);
and U27858 (N_27858,N_25680,N_25777);
xnor U27859 (N_27859,N_27393,N_25033);
or U27860 (N_27860,N_25944,N_27376);
or U27861 (N_27861,N_26812,N_25606);
nor U27862 (N_27862,N_27453,N_25145);
or U27863 (N_27863,N_25076,N_27327);
nand U27864 (N_27864,N_27331,N_26285);
nor U27865 (N_27865,N_25770,N_25635);
nor U27866 (N_27866,N_25957,N_26752);
nor U27867 (N_27867,N_27223,N_26522);
or U27868 (N_27868,N_27163,N_25504);
xnor U27869 (N_27869,N_26765,N_27334);
or U27870 (N_27870,N_26684,N_25420);
nand U27871 (N_27871,N_25771,N_27035);
xnor U27872 (N_27872,N_27361,N_25355);
or U27873 (N_27873,N_27048,N_25365);
nand U27874 (N_27874,N_25167,N_25322);
and U27875 (N_27875,N_25605,N_27105);
xor U27876 (N_27876,N_26673,N_26680);
nand U27877 (N_27877,N_25336,N_27260);
or U27878 (N_27878,N_26608,N_26778);
nand U27879 (N_27879,N_26863,N_27489);
xnor U27880 (N_27880,N_26641,N_25270);
xor U27881 (N_27881,N_27308,N_25386);
xnor U27882 (N_27882,N_25411,N_26750);
nor U27883 (N_27883,N_25377,N_25044);
and U27884 (N_27884,N_25744,N_26450);
nand U27885 (N_27885,N_26441,N_25155);
and U27886 (N_27886,N_27140,N_27297);
or U27887 (N_27887,N_27363,N_26550);
xor U27888 (N_27888,N_25526,N_26782);
or U27889 (N_27889,N_27042,N_26855);
nand U27890 (N_27890,N_27386,N_25394);
and U27891 (N_27891,N_25669,N_26714);
or U27892 (N_27892,N_25715,N_26805);
nor U27893 (N_27893,N_27414,N_27015);
xnor U27894 (N_27894,N_25917,N_27256);
nand U27895 (N_27895,N_25100,N_25207);
nand U27896 (N_27896,N_25404,N_26011);
nand U27897 (N_27897,N_25999,N_25711);
xor U27898 (N_27898,N_26125,N_26995);
nand U27899 (N_27899,N_27351,N_26455);
and U27900 (N_27900,N_26888,N_26344);
nor U27901 (N_27901,N_26332,N_25964);
and U27902 (N_27902,N_25055,N_26646);
xor U27903 (N_27903,N_25874,N_25459);
xnor U27904 (N_27904,N_26206,N_26900);
nand U27905 (N_27905,N_26447,N_26918);
and U27906 (N_27906,N_26342,N_25873);
xor U27907 (N_27907,N_27290,N_26431);
nor U27908 (N_27908,N_26274,N_25805);
nor U27909 (N_27909,N_25651,N_25169);
nand U27910 (N_27910,N_27395,N_25031);
or U27911 (N_27911,N_26138,N_26056);
or U27912 (N_27912,N_25222,N_25992);
nor U27913 (N_27913,N_25235,N_26256);
nor U27914 (N_27914,N_26166,N_27213);
xor U27915 (N_27915,N_25603,N_26419);
xor U27916 (N_27916,N_25910,N_25965);
xor U27917 (N_27917,N_26770,N_26380);
nor U27918 (N_27918,N_25277,N_25817);
or U27919 (N_27919,N_26796,N_26253);
xor U27920 (N_27920,N_25025,N_26983);
and U27921 (N_27921,N_25485,N_27055);
and U27922 (N_27922,N_27019,N_25705);
xnor U27923 (N_27923,N_26497,N_25127);
and U27924 (N_27924,N_26925,N_25448);
xor U27925 (N_27925,N_26981,N_26291);
nand U27926 (N_27926,N_26947,N_25746);
nor U27927 (N_27927,N_25923,N_26046);
nand U27928 (N_27928,N_26559,N_26506);
and U27929 (N_27929,N_26819,N_25929);
and U27930 (N_27930,N_25022,N_26906);
xor U27931 (N_27931,N_27209,N_26619);
or U27932 (N_27932,N_27335,N_25634);
nor U27933 (N_27933,N_26580,N_26706);
and U27934 (N_27934,N_26182,N_25294);
xnor U27935 (N_27935,N_26072,N_25362);
or U27936 (N_27936,N_25198,N_27082);
or U27937 (N_27937,N_26886,N_25045);
and U27938 (N_27938,N_26461,N_26553);
or U27939 (N_27939,N_27387,N_26191);
nor U27940 (N_27940,N_26411,N_26579);
nor U27941 (N_27941,N_25909,N_27020);
nor U27942 (N_27942,N_25523,N_27013);
and U27943 (N_27943,N_25621,N_25130);
or U27944 (N_27944,N_25742,N_25995);
nand U27945 (N_27945,N_26662,N_26645);
xnor U27946 (N_27946,N_26783,N_26816);
nor U27947 (N_27947,N_25945,N_26744);
nand U27948 (N_27948,N_26734,N_25926);
nand U27949 (N_27949,N_26758,N_26365);
nor U27950 (N_27950,N_25281,N_26345);
xor U27951 (N_27951,N_25638,N_27486);
nand U27952 (N_27952,N_25633,N_27432);
or U27953 (N_27953,N_25391,N_25660);
nor U27954 (N_27954,N_26560,N_26913);
and U27955 (N_27955,N_26607,N_26180);
and U27956 (N_27956,N_25266,N_27469);
and U27957 (N_27957,N_26793,N_25721);
or U27958 (N_27958,N_25612,N_26789);
and U27959 (N_27959,N_26749,N_26349);
nor U27960 (N_27960,N_26620,N_25179);
nor U27961 (N_27961,N_26333,N_27462);
nor U27962 (N_27962,N_26244,N_26063);
and U27963 (N_27963,N_25794,N_26868);
and U27964 (N_27964,N_25288,N_25265);
nor U27965 (N_27965,N_26398,N_26875);
or U27966 (N_27966,N_25954,N_25433);
or U27967 (N_27967,N_26721,N_25466);
nor U27968 (N_27968,N_26037,N_26978);
xor U27969 (N_27969,N_26312,N_25961);
nor U27970 (N_27970,N_26651,N_25024);
xnor U27971 (N_27971,N_25800,N_27066);
xnor U27972 (N_27972,N_25064,N_26338);
nand U27973 (N_27973,N_26896,N_26415);
or U27974 (N_27974,N_26264,N_26801);
or U27975 (N_27975,N_27371,N_25160);
or U27976 (N_27976,N_25005,N_25456);
and U27977 (N_27977,N_25084,N_26803);
or U27978 (N_27978,N_27433,N_26542);
nor U27979 (N_27979,N_26870,N_25441);
xor U27980 (N_27980,N_26040,N_26814);
xnor U27981 (N_27981,N_26543,N_26308);
nor U27982 (N_27982,N_25509,N_26998);
and U27983 (N_27983,N_26936,N_25565);
and U27984 (N_27984,N_25912,N_26377);
xor U27985 (N_27985,N_27400,N_25296);
xnor U27986 (N_27986,N_26229,N_26276);
and U27987 (N_27987,N_25889,N_25661);
nor U27988 (N_27988,N_26760,N_25418);
xnor U27989 (N_27989,N_25280,N_26577);
nor U27990 (N_27990,N_26267,N_25536);
nand U27991 (N_27991,N_27081,N_25806);
or U27992 (N_27992,N_26372,N_25272);
nor U27993 (N_27993,N_27160,N_25416);
nor U27994 (N_27994,N_25166,N_27349);
nor U27995 (N_27995,N_26169,N_26179);
nor U27996 (N_27996,N_26873,N_26313);
xnor U27997 (N_27997,N_25350,N_25148);
and U27998 (N_27998,N_26391,N_27341);
nand U27999 (N_27999,N_25178,N_25213);
nand U28000 (N_28000,N_25686,N_26531);
and U28001 (N_28001,N_25182,N_26979);
nand U28002 (N_28002,N_26211,N_26127);
nor U28003 (N_28003,N_27088,N_25802);
xnor U28004 (N_28004,N_27282,N_25407);
xnor U28005 (N_28005,N_25305,N_25581);
nand U28006 (N_28006,N_25969,N_27067);
or U28007 (N_28007,N_25097,N_26096);
and U28008 (N_28008,N_27380,N_25844);
nor U28009 (N_28009,N_27093,N_26730);
nand U28010 (N_28010,N_27340,N_25960);
nor U28011 (N_28011,N_26661,N_26010);
or U28012 (N_28012,N_26736,N_25402);
nor U28013 (N_28013,N_25872,N_26675);
nand U28014 (N_28014,N_26159,N_25758);
or U28015 (N_28015,N_25654,N_25542);
xor U28016 (N_28016,N_26379,N_27074);
or U28017 (N_28017,N_26404,N_27219);
and U28018 (N_28018,N_26024,N_26287);
nor U28019 (N_28019,N_26328,N_25996);
nand U28020 (N_28020,N_26396,N_27034);
or U28021 (N_28021,N_26048,N_25507);
nor U28022 (N_28022,N_26436,N_27271);
or U28023 (N_28023,N_25057,N_27099);
nand U28024 (N_28024,N_26658,N_26331);
and U28025 (N_28025,N_26515,N_26509);
nand U28026 (N_28026,N_25924,N_27346);
nor U28027 (N_28027,N_25172,N_26564);
or U28028 (N_28028,N_25679,N_25364);
xnor U28029 (N_28029,N_26239,N_25557);
nor U28030 (N_28030,N_25486,N_25702);
nand U28031 (N_28031,N_27348,N_25567);
or U28032 (N_28032,N_26676,N_26625);
xor U28033 (N_28033,N_26327,N_25836);
xor U28034 (N_28034,N_26739,N_25922);
xnor U28035 (N_28035,N_27442,N_26089);
nor U28036 (N_28036,N_26173,N_26145);
nor U28037 (N_28037,N_27439,N_25227);
xnor U28038 (N_28038,N_26586,N_26077);
and U28039 (N_28039,N_26064,N_26093);
xnor U28040 (N_28040,N_26201,N_25855);
or U28041 (N_28041,N_25328,N_25979);
nor U28042 (N_28042,N_25857,N_25034);
and U28043 (N_28043,N_26720,N_27065);
xnor U28044 (N_28044,N_27443,N_26952);
nand U28045 (N_28045,N_26631,N_26938);
or U28046 (N_28046,N_26776,N_25971);
nor U28047 (N_28047,N_25123,N_26226);
and U28048 (N_28048,N_26316,N_25582);
or U28049 (N_28049,N_25473,N_25062);
nor U28050 (N_28050,N_27272,N_26083);
nor U28051 (N_28051,N_25259,N_25839);
nand U28052 (N_28052,N_26036,N_25290);
xnor U28053 (N_28053,N_26386,N_26292);
xnor U28054 (N_28054,N_25689,N_26871);
or U28055 (N_28055,N_26304,N_25982);
and U28056 (N_28056,N_25616,N_25308);
nand U28057 (N_28057,N_25273,N_27189);
or U28058 (N_28058,N_26408,N_27254);
xor U28059 (N_28059,N_26667,N_26044);
or U28060 (N_28060,N_26948,N_26511);
nor U28061 (N_28061,N_25939,N_26822);
or U28062 (N_28062,N_27026,N_25703);
xor U28063 (N_28063,N_27375,N_26593);
or U28064 (N_28064,N_27465,N_27392);
and U28065 (N_28065,N_25211,N_25958);
and U28066 (N_28066,N_25457,N_27487);
and U28067 (N_28067,N_27043,N_26121);
and U28068 (N_28068,N_26512,N_25870);
nand U28069 (N_28069,N_25752,N_26126);
nor U28070 (N_28070,N_26931,N_26449);
nor U28071 (N_28071,N_26682,N_26452);
nand U28072 (N_28072,N_26848,N_26583);
nor U28073 (N_28073,N_26993,N_27326);
nor U28074 (N_28074,N_26650,N_26192);
and U28075 (N_28075,N_25226,N_25931);
nand U28076 (N_28076,N_26525,N_26482);
and U28077 (N_28077,N_25194,N_25598);
and U28078 (N_28078,N_25666,N_25150);
nor U28079 (N_28079,N_25956,N_25801);
xnor U28080 (N_28080,N_26713,N_25188);
nor U28081 (N_28081,N_25754,N_25032);
or U28082 (N_28082,N_25037,N_25131);
and U28083 (N_28083,N_25012,N_25419);
and U28084 (N_28084,N_25200,N_25846);
xor U28085 (N_28085,N_25837,N_25349);
xnor U28086 (N_28086,N_25643,N_26401);
and U28087 (N_28087,N_25112,N_25465);
xnor U28088 (N_28088,N_26200,N_26395);
nor U28089 (N_28089,N_26681,N_25284);
xnor U28090 (N_28090,N_25832,N_26221);
or U28091 (N_28091,N_27158,N_26618);
and U28092 (N_28092,N_26154,N_26921);
or U28093 (N_28093,N_26521,N_26962);
xor U28094 (N_28094,N_25040,N_25701);
nand U28095 (N_28095,N_27221,N_27448);
and U28096 (N_28096,N_25553,N_27232);
and U28097 (N_28097,N_25699,N_25665);
nand U28098 (N_28098,N_27184,N_25807);
or U28099 (N_28099,N_26563,N_25424);
nand U28100 (N_28100,N_26246,N_26571);
and U28101 (N_28101,N_25998,N_25449);
or U28102 (N_28102,N_26230,N_26516);
and U28103 (N_28103,N_25622,N_27155);
and U28104 (N_28104,N_25118,N_26248);
nand U28105 (N_28105,N_26257,N_25455);
nand U28106 (N_28106,N_25953,N_25482);
and U28107 (N_28107,N_25186,N_26847);
and U28108 (N_28108,N_26076,N_25256);
and U28109 (N_28109,N_27304,N_26081);
nand U28110 (N_28110,N_26068,N_26788);
xnor U28111 (N_28111,N_25738,N_25339);
xor U28112 (N_28112,N_26134,N_25596);
nand U28113 (N_28113,N_25410,N_26520);
or U28114 (N_28114,N_26798,N_25430);
or U28115 (N_28115,N_25156,N_26989);
nor U28116 (N_28116,N_25385,N_26901);
or U28117 (N_28117,N_26314,N_25614);
nand U28118 (N_28118,N_27264,N_27193);
and U28119 (N_28119,N_25914,N_25983);
or U28120 (N_28120,N_25893,N_26005);
xnor U28121 (N_28121,N_25343,N_25469);
xor U28122 (N_28122,N_25095,N_25657);
nor U28123 (N_28123,N_27404,N_25584);
and U28124 (N_28124,N_26095,N_25574);
or U28125 (N_28125,N_26457,N_26604);
or U28126 (N_28126,N_25153,N_25219);
xor U28127 (N_28127,N_25291,N_25988);
or U28128 (N_28128,N_25769,N_25902);
and U28129 (N_28129,N_25346,N_27224);
nand U28130 (N_28130,N_26643,N_25881);
or U28131 (N_28131,N_26771,N_27295);
and U28132 (N_28132,N_26878,N_27283);
nor U28133 (N_28133,N_27003,N_25720);
nor U28134 (N_28134,N_26709,N_25568);
or U28135 (N_28135,N_25775,N_25919);
and U28136 (N_28136,N_26373,N_25061);
nor U28137 (N_28137,N_25117,N_27016);
or U28138 (N_28138,N_27182,N_25443);
nand U28139 (N_28139,N_27316,N_26478);
and U28140 (N_28140,N_25378,N_27266);
nand U28141 (N_28141,N_25773,N_26474);
or U28142 (N_28142,N_26266,N_26883);
nor U28143 (N_28143,N_26861,N_25591);
xor U28144 (N_28144,N_25897,N_27142);
or U28145 (N_28145,N_27125,N_26784);
nand U28146 (N_28146,N_25898,N_26898);
nand U28147 (N_28147,N_26013,N_26442);
or U28148 (N_28148,N_27152,N_25658);
and U28149 (N_28149,N_26751,N_27457);
xnor U28150 (N_28150,N_26635,N_26723);
and U28151 (N_28151,N_27288,N_25697);
or U28152 (N_28152,N_26350,N_25610);
and U28153 (N_28153,N_26086,N_25722);
nand U28154 (N_28154,N_26687,N_26845);
nor U28155 (N_28155,N_26467,N_27472);
or U28156 (N_28156,N_27429,N_25743);
and U28157 (N_28157,N_27236,N_26023);
or U28158 (N_28158,N_25757,N_25972);
nor U28159 (N_28159,N_27435,N_25333);
or U28160 (N_28160,N_25323,N_25489);
xnor U28161 (N_28161,N_26634,N_25384);
nor U28162 (N_28162,N_26656,N_27460);
nand U28163 (N_28163,N_25712,N_26678);
xnor U28164 (N_28164,N_26766,N_27173);
xnor U28165 (N_28165,N_26456,N_27176);
and U28166 (N_28166,N_26006,N_27249);
nor U28167 (N_28167,N_26459,N_26335);
nand U28168 (N_28168,N_25959,N_26352);
or U28169 (N_28169,N_25973,N_26363);
and U28170 (N_28170,N_27421,N_26311);
or U28171 (N_28171,N_26184,N_25250);
nand U28172 (N_28172,N_25877,N_26502);
and U28173 (N_28173,N_27291,N_25640);
xor U28174 (N_28174,N_26518,N_26188);
or U28175 (N_28175,N_26513,N_27006);
nor U28176 (N_28176,N_26212,N_25108);
nor U28177 (N_28177,N_27000,N_26630);
and U28178 (N_28178,N_25503,N_26800);
or U28179 (N_28179,N_26674,N_25120);
or U28180 (N_28180,N_25269,N_26417);
nor U28181 (N_28181,N_25010,N_26768);
and U28182 (N_28182,N_27367,N_27355);
and U28183 (N_28183,N_25020,N_25860);
xnor U28184 (N_28184,N_26660,N_26928);
nand U28185 (N_28185,N_26278,N_25617);
xor U28186 (N_28186,N_25051,N_25370);
nor U28187 (N_28187,N_26835,N_25595);
or U28188 (N_28188,N_27463,N_25570);
nand U28189 (N_28189,N_26326,N_26102);
nor U28190 (N_28190,N_25262,N_26903);
nor U28191 (N_28191,N_26021,N_27270);
xnor U28192 (N_28192,N_26194,N_26307);
xnor U28193 (N_28193,N_26424,N_25422);
or U28194 (N_28194,N_25563,N_26986);
or U28195 (N_28195,N_25440,N_25761);
xnor U28196 (N_28196,N_25347,N_27333);
xor U28197 (N_28197,N_26679,N_27207);
xnor U28198 (N_28198,N_26185,N_25887);
nand U28199 (N_28199,N_26548,N_27131);
and U28200 (N_28200,N_26769,N_27102);
or U28201 (N_28201,N_25423,N_25952);
nor U28202 (N_28202,N_25028,N_26153);
nor U28203 (N_28203,N_26272,N_26567);
nand U28204 (N_28204,N_25079,N_25495);
nor U28205 (N_28205,N_26990,N_26792);
nor U28206 (N_28206,N_26554,N_25677);
nor U28207 (N_28207,N_26544,N_26196);
or U28208 (N_28208,N_25940,N_26358);
nor U28209 (N_28209,N_27356,N_25827);
nor U28210 (N_28210,N_25976,N_26058);
nand U28211 (N_28211,N_27336,N_26849);
xnor U28212 (N_28212,N_27064,N_26926);
and U28213 (N_28213,N_27080,N_25993);
or U28214 (N_28214,N_25838,N_27296);
nor U28215 (N_28215,N_25387,N_27408);
or U28216 (N_28216,N_25098,N_25491);
xor U28217 (N_28217,N_26807,N_27101);
nor U28218 (N_28218,N_25367,N_27343);
nor U28219 (N_28219,N_26174,N_26429);
nor U28220 (N_28220,N_25879,N_25041);
xor U28221 (N_28221,N_27197,N_26541);
and U28222 (N_28222,N_26237,N_26624);
xnor U28223 (N_28223,N_27100,N_25056);
nor U28224 (N_28224,N_26846,N_25681);
nor U28225 (N_28225,N_26440,N_25381);
and U28226 (N_28226,N_26529,N_25828);
xor U28227 (N_28227,N_25876,N_25962);
and U28228 (N_28228,N_27205,N_27014);
and U28229 (N_28229,N_25737,N_25390);
nor U28230 (N_28230,N_25348,N_26139);
nor U28231 (N_28231,N_27407,N_27130);
nand U28232 (N_28232,N_27106,N_26491);
xnor U28233 (N_28233,N_26357,N_26879);
nor U28234 (N_28234,N_26877,N_26636);
or U28235 (N_28235,N_25292,N_25480);
nand U28236 (N_28236,N_26841,N_27417);
or U28237 (N_28237,N_27330,N_25641);
xor U28238 (N_28238,N_25908,N_27372);
nor U28239 (N_28239,N_27447,N_26199);
and U28240 (N_28240,N_25077,N_27183);
or U28241 (N_28241,N_25408,N_25282);
and U28242 (N_28242,N_26070,N_26108);
nand U28243 (N_28243,N_25515,N_26762);
or U28244 (N_28244,N_27317,N_25268);
xor U28245 (N_28245,N_27315,N_27275);
xnor U28246 (N_28246,N_26696,N_27135);
and U28247 (N_28247,N_27052,N_25611);
xnor U28248 (N_28248,N_25704,N_26694);
or U28249 (N_28249,N_25017,N_26137);
and U28250 (N_28250,N_27468,N_25891);
or U28251 (N_28251,N_25531,N_26476);
nand U28252 (N_28252,N_26836,N_27262);
and U28253 (N_28253,N_25724,N_26062);
or U28254 (N_28254,N_25540,N_25224);
and U28255 (N_28255,N_25655,N_27036);
or U28256 (N_28256,N_25376,N_27113);
or U28257 (N_28257,N_26958,N_26919);
nand U28258 (N_28258,N_27046,N_25751);
or U28259 (N_28259,N_26876,N_25916);
nor U28260 (N_28260,N_26309,N_26626);
nand U28261 (N_28261,N_26772,N_27278);
and U28262 (N_28262,N_26647,N_26523);
nand U28263 (N_28263,N_25453,N_27352);
or U28264 (N_28264,N_25522,N_25642);
and U28265 (N_28265,N_25329,N_25243);
nand U28266 (N_28266,N_25950,N_26818);
and U28267 (N_28267,N_27274,N_26982);
and U28268 (N_28268,N_25088,N_26477);
or U28269 (N_28269,N_25835,N_25615);
xor U28270 (N_28270,N_25388,N_26558);
nor U28271 (N_28271,N_27037,N_26128);
and U28272 (N_28272,N_25586,N_25997);
xnor U28273 (N_28273,N_26880,N_25883);
or U28274 (N_28274,N_26533,N_25550);
and U28275 (N_28275,N_27360,N_26815);
and U28276 (N_28276,N_26351,N_26612);
and U28277 (N_28277,N_25287,N_26343);
nand U28278 (N_28278,N_25899,N_25517);
nor U28279 (N_28279,N_26627,N_27280);
nor U28280 (N_28280,N_27002,N_26915);
nor U28281 (N_28281,N_26657,N_25728);
or U28282 (N_28282,N_25825,N_25723);
and U28283 (N_28283,N_26465,N_26555);
and U28284 (N_28284,N_26813,N_26254);
nor U28285 (N_28285,N_25371,N_25002);
nor U28286 (N_28286,N_27456,N_27070);
or U28287 (N_28287,N_27044,N_26428);
or U28288 (N_28288,N_25129,N_27032);
or U28289 (N_28289,N_26294,N_25497);
nand U28290 (N_28290,N_27206,N_26632);
and U28291 (N_28291,N_26688,N_25693);
nor U28292 (N_28292,N_26163,N_26584);
nand U28293 (N_28293,N_26881,N_26146);
nor U28294 (N_28294,N_25718,N_26105);
nor U28295 (N_28295,N_26376,N_27464);
and U28296 (N_28296,N_25432,N_25383);
nand U28297 (N_28297,N_27273,N_25840);
and U28298 (N_28298,N_26677,N_26060);
nand U28299 (N_28299,N_25913,N_26486);
nor U28300 (N_28300,N_26717,N_25968);
and U28301 (N_28301,N_26601,N_26594);
nor U28302 (N_28302,N_27268,N_25075);
xnor U28303 (N_28303,N_25374,N_25152);
xor U28304 (N_28304,N_25099,N_27194);
and U28305 (N_28305,N_26038,N_27010);
xor U28306 (N_28306,N_26075,N_25508);
or U28307 (N_28307,N_25113,N_27234);
nor U28308 (N_28308,N_27402,N_25406);
or U28309 (N_28309,N_26711,N_25232);
nand U28310 (N_28310,N_25114,N_26549);
nor U28311 (N_28311,N_27068,N_26277);
or U28312 (N_28312,N_25400,N_25151);
and U28313 (N_28313,N_25589,N_26049);
nor U28314 (N_28314,N_27491,N_27058);
nand U28315 (N_28315,N_26397,N_27050);
xnor U28316 (N_28316,N_27478,N_27040);
nand U28317 (N_28317,N_25862,N_25561);
or U28318 (N_28318,N_25946,N_26469);
nand U28319 (N_28319,N_26994,N_26858);
or U28320 (N_28320,N_25253,N_26764);
or U28321 (N_28321,N_26347,N_26924);
xnor U28322 (N_28322,N_26862,N_25074);
nand U28323 (N_28323,N_26162,N_25444);
xnor U28324 (N_28324,N_26895,N_25671);
or U28325 (N_28325,N_25018,N_27073);
nand U28326 (N_28326,N_26433,N_27405);
nor U28327 (N_28327,N_25216,N_26334);
xor U28328 (N_28328,N_25425,N_26172);
and U28329 (N_28329,N_25236,N_25244);
and U28330 (N_28330,N_26355,N_25613);
or U28331 (N_28331,N_25335,N_25102);
nand U28332 (N_28332,N_25823,N_27425);
or U28333 (N_28333,N_25431,N_26353);
and U28334 (N_28334,N_26927,N_27498);
or U28335 (N_28335,N_26562,N_27127);
nand U28336 (N_28336,N_26364,N_26844);
nor U28337 (N_28337,N_26732,N_25767);
xnor U28338 (N_28338,N_27190,N_26115);
nand U28339 (N_28339,N_26468,N_26699);
nand U28340 (N_28340,N_26621,N_25036);
nand U28341 (N_28341,N_25171,N_25991);
nand U28342 (N_28342,N_25780,N_27147);
xnor U28343 (N_28343,N_26359,N_27202);
nor U28344 (N_28344,N_25487,N_26123);
and U28345 (N_28345,N_25859,N_26020);
xor U28346 (N_28346,N_25004,N_25251);
and U28347 (N_28347,N_26444,N_25019);
and U28348 (N_28348,N_26628,N_27210);
nand U28349 (N_28349,N_26710,N_27137);
or U28350 (N_28350,N_27287,N_25475);
or U28351 (N_28351,N_26934,N_25278);
xor U28352 (N_28352,N_27446,N_26481);
nor U28353 (N_28353,N_27119,N_26485);
and U28354 (N_28354,N_25569,N_25829);
nor U28355 (N_28355,N_27299,N_26622);
xnor U28356 (N_28356,N_26385,N_25867);
xor U28357 (N_28357,N_26152,N_25726);
nor U28358 (N_28358,N_26795,N_26238);
or U28359 (N_28359,N_25985,N_25987);
xor U28360 (N_28360,N_25534,N_27171);
or U28361 (N_28361,N_26147,N_26445);
and U28362 (N_28362,N_27277,N_27079);
nor U28363 (N_28363,N_26223,N_26530);
xor U28364 (N_28364,N_26175,N_27394);
xor U28365 (N_28365,N_27409,N_26132);
and U28366 (N_28366,N_25716,N_27305);
nand U28367 (N_28367,N_27424,N_26375);
or U28368 (N_28368,N_27384,N_27161);
nor U28369 (N_28369,N_26970,N_26389);
nand U28370 (N_28370,N_26104,N_26203);
nor U28371 (N_28371,N_25356,N_26016);
or U28372 (N_28372,N_25261,N_27423);
or U28373 (N_28373,N_27107,N_25977);
nor U28374 (N_28374,N_27267,N_26279);
and U28375 (N_28375,N_27416,N_27415);
and U28376 (N_28376,N_26725,N_25842);
nor U28377 (N_28377,N_26767,N_25778);
and U28378 (N_28378,N_26719,N_26831);
xor U28379 (N_28379,N_27126,N_27109);
nand U28380 (N_28380,N_27001,N_25673);
or U28381 (N_28381,N_25766,N_25691);
nor U28382 (N_28382,N_26780,N_25454);
xnor U28383 (N_28383,N_26827,N_25217);
nor U28384 (N_28384,N_26589,N_26592);
nand U28385 (N_28385,N_25214,N_25310);
and U28386 (N_28386,N_26034,N_26991);
xor U28387 (N_28387,N_25185,N_25183);
and U28388 (N_28388,N_25255,N_26966);
and U28389 (N_28389,N_25544,N_26790);
and U28390 (N_28390,N_25851,N_26690);
and U28391 (N_28391,N_25779,N_26545);
and U28392 (N_28392,N_25078,N_25176);
nor U28393 (N_28393,N_25357,N_26753);
nor U28394 (N_28394,N_25229,N_27259);
nor U28395 (N_28395,N_26090,N_25713);
nand U28396 (N_28396,N_25434,N_25833);
and U28397 (N_28397,N_25468,N_26930);
or U28398 (N_28398,N_25955,N_25963);
nand U28399 (N_28399,N_25809,N_25038);
or U28400 (N_28400,N_26843,N_26623);
nand U28401 (N_28401,N_26852,N_26434);
or U28402 (N_28402,N_25683,N_25249);
nor U28403 (N_28403,N_25776,N_25886);
nor U28404 (N_28404,N_26742,N_25510);
or U28405 (N_28405,N_25029,N_26740);
and U28406 (N_28406,N_27494,N_26484);
nand U28407 (N_28407,N_26065,N_25302);
xor U28408 (N_28408,N_25375,N_26092);
nor U28409 (N_28409,N_25978,N_26061);
nor U28410 (N_28410,N_26882,N_27181);
and U28411 (N_28411,N_25543,N_27167);
xnor U28412 (N_28412,N_27199,N_27087);
and U28413 (N_28413,N_26757,N_26236);
xor U28414 (N_28414,N_26598,N_27072);
xor U28415 (N_28415,N_25000,N_26463);
or U28416 (N_28416,N_25663,N_27426);
nand U28417 (N_28417,N_26595,N_27208);
and U28418 (N_28418,N_27059,N_27009);
nand U28419 (N_28419,N_26605,N_26047);
xor U28420 (N_28420,N_26393,N_26208);
or U28421 (N_28421,N_26189,N_25165);
or U28422 (N_28422,N_26019,N_26435);
nand U28423 (N_28423,N_26655,N_25460);
and U28424 (N_28424,N_25793,N_25477);
or U28425 (N_28425,N_26907,N_25994);
nand U28426 (N_28426,N_25141,N_25690);
and U28427 (N_28427,N_25513,N_26665);
nor U28428 (N_28428,N_26317,N_25189);
or U28429 (N_28429,N_25639,N_26321);
and U28430 (N_28430,N_27399,N_25787);
or U28431 (N_28431,N_26235,N_25461);
nand U28432 (N_28432,N_26114,N_26283);
nand U28433 (N_28433,N_26917,N_25585);
and U28434 (N_28434,N_26421,N_26839);
xor U28435 (N_28435,N_27383,N_26052);
nor U28436 (N_28436,N_27231,N_26968);
or U28437 (N_28437,N_27118,N_27477);
nor U28438 (N_28438,N_27320,N_27496);
nand U28439 (N_28439,N_25299,N_25237);
xor U28440 (N_28440,N_25739,N_25311);
xnor U28441 (N_28441,N_26488,N_25552);
nor U28442 (N_28442,N_25071,N_25048);
and U28443 (N_28443,N_27365,N_26270);
and U28444 (N_28444,N_27239,N_26069);
and U28445 (N_28445,N_25293,N_27146);
and U28446 (N_28446,N_26483,N_26324);
or U28447 (N_28447,N_26600,N_26103);
nor U28448 (N_28448,N_25109,N_25572);
and U28449 (N_28449,N_25904,N_27490);
or U28450 (N_28450,N_26027,N_25786);
xnor U28451 (N_28451,N_25537,N_26033);
or U28452 (N_28452,N_25824,N_26118);
nor U28453 (N_28453,N_25915,N_27076);
nor U28454 (N_28454,N_26480,N_26997);
or U28455 (N_28455,N_25501,N_26029);
nand U28456 (N_28456,N_26902,N_25656);
xor U28457 (N_28457,N_25948,N_26207);
or U28458 (N_28458,N_26339,N_27212);
nor U28459 (N_28459,N_26209,N_27373);
or U28460 (N_28460,N_26922,N_25332);
nand U28461 (N_28461,N_26629,N_27344);
nand U28462 (N_28462,N_27431,N_26869);
nand U28463 (N_28463,N_25442,N_26933);
nor U28464 (N_28464,N_27007,N_26002);
and U28465 (N_28465,N_27310,N_27258);
and U28466 (N_28466,N_25498,N_25429);
or U28467 (N_28467,N_26422,N_25625);
and U28468 (N_28468,N_25321,N_25760);
and U28469 (N_28469,N_26539,N_26250);
and U28470 (N_28470,N_27479,N_25220);
and U28471 (N_28471,N_26156,N_26490);
and U28472 (N_28472,N_26113,N_26181);
nand U28473 (N_28473,N_26668,N_27128);
or U28474 (N_28474,N_25049,N_25307);
nand U28475 (N_28475,N_25191,N_26899);
nand U28476 (N_28476,N_26551,N_25135);
xnor U28477 (N_28477,N_25578,N_26670);
nor U28478 (N_28478,N_27154,N_25784);
nand U28479 (N_28479,N_25315,N_27164);
or U28480 (N_28480,N_26148,N_25685);
xnor U28481 (N_28481,N_26718,N_25428);
and U28482 (N_28482,N_26262,N_27265);
nor U28483 (N_28483,N_26920,N_26085);
or U28484 (N_28484,N_26315,N_25951);
and U28485 (N_28485,N_27045,N_26158);
or U28486 (N_28486,N_26409,N_25607);
nor U28487 (N_28487,N_27092,N_26259);
and U28488 (N_28488,N_26799,N_27168);
and U28489 (N_28489,N_26039,N_25363);
xnor U28490 (N_28490,N_27437,N_26644);
and U28491 (N_28491,N_25058,N_26195);
xnor U28492 (N_28492,N_26101,N_26003);
nand U28493 (N_28493,N_25869,N_25907);
nor U28494 (N_28494,N_26073,N_26150);
xor U28495 (N_28495,N_25298,N_25694);
nor U28496 (N_28496,N_26857,N_26590);
nand U28497 (N_28497,N_26439,N_25521);
and U28498 (N_28498,N_25260,N_26663);
xnor U28499 (N_28499,N_27157,N_25875);
xor U28500 (N_28500,N_26842,N_26536);
nor U28501 (N_28501,N_27056,N_27023);
or U28502 (N_28502,N_26493,N_27253);
nor U28503 (N_28503,N_26290,N_26640);
or U28504 (N_28504,N_25980,N_25264);
and U28505 (N_28505,N_26972,N_26106);
or U28506 (N_28506,N_25573,N_27284);
or U28507 (N_28507,N_25106,N_27313);
or U28508 (N_28508,N_26131,N_27075);
nand U28509 (N_28509,N_26865,N_25594);
nor U28510 (N_28510,N_25415,N_26470);
or U28511 (N_28511,N_26950,N_27244);
xnor U28512 (N_28512,N_26241,N_25548);
xor U28513 (N_28513,N_27114,N_26686);
and U28514 (N_28514,N_25629,N_27051);
or U28515 (N_28515,N_26825,N_25476);
xnor U28516 (N_28516,N_27388,N_25094);
xnor U28517 (N_28517,N_26832,N_25845);
nand U28518 (N_28518,N_26227,N_26726);
nor U28519 (N_28519,N_26462,N_25700);
and U28520 (N_28520,N_26471,N_27139);
nor U28521 (N_28521,N_25735,N_26617);
and U28522 (N_28522,N_25133,N_25001);
or U28523 (N_28523,N_27047,N_25492);
nor U28524 (N_28524,N_25818,N_26967);
or U28525 (N_28525,N_26672,N_25297);
and U28526 (N_28526,N_25528,N_25138);
xor U28527 (N_28527,N_27170,N_27091);
nand U28528 (N_28528,N_27095,N_25212);
xnor U28529 (N_28529,N_25089,N_26859);
nor U28530 (N_28530,N_25409,N_27214);
nor U28531 (N_28531,N_27112,N_25684);
and U28532 (N_28532,N_27218,N_25006);
xnor U28533 (N_28533,N_26578,N_26091);
xor U28534 (N_28534,N_26388,N_26325);
nand U28535 (N_28535,N_26232,N_25830);
xnor U28536 (N_28536,N_25379,N_25373);
nand U28537 (N_28537,N_27240,N_27008);
or U28538 (N_28538,N_26054,N_26704);
nand U28539 (N_28539,N_27025,N_25707);
xnor U28540 (N_28540,N_26824,N_26754);
nor U28541 (N_28541,N_25147,N_26050);
and U28542 (N_28542,N_27096,N_25849);
nand U28543 (N_28543,N_25530,N_26306);
and U28544 (N_28544,N_25279,N_27293);
or U28545 (N_28545,N_26851,N_26004);
and U28546 (N_28546,N_26432,N_25344);
nand U28547 (N_28547,N_27011,N_25412);
nor U28548 (N_28548,N_27499,N_27377);
and U28549 (N_28549,N_26996,N_25731);
and U28550 (N_28550,N_26453,N_25930);
or U28551 (N_28551,N_26953,N_27104);
and U28552 (N_28552,N_25181,N_27097);
or U28553 (N_28553,N_27222,N_27449);
or U28554 (N_28554,N_26565,N_25121);
nand U28555 (N_28555,N_26320,N_27123);
nor U28556 (N_28556,N_25392,N_25303);
nor U28557 (N_28557,N_27129,N_27159);
and U28558 (N_28558,N_25593,N_26964);
xor U28559 (N_28559,N_26014,N_25170);
nor U28560 (N_28560,N_25334,N_25730);
nor U28561 (N_28561,N_26361,N_26697);
nor U28562 (N_28562,N_26260,N_26498);
nor U28563 (N_28563,N_25900,N_25890);
xor U28564 (N_28564,N_27090,N_27024);
nand U28565 (N_28565,N_26526,N_25464);
nand U28566 (N_28566,N_27342,N_27177);
and U28567 (N_28567,N_25324,N_27444);
xor U28568 (N_28568,N_26204,N_26535);
xnor U28569 (N_28569,N_25072,N_25670);
or U28570 (N_28570,N_26399,N_25493);
or U28571 (N_28571,N_26664,N_26362);
nand U28572 (N_28572,N_26941,N_26826);
xor U28573 (N_28573,N_26712,N_27242);
xnor U28574 (N_28574,N_27474,N_25086);
and U28575 (N_28575,N_26537,N_25853);
xnor U28576 (N_28576,N_26591,N_25505);
nand U28577 (N_28577,N_27255,N_26197);
nor U28578 (N_28578,N_26066,N_25920);
xor U28579 (N_28579,N_27410,N_26009);
xnor U28580 (N_28580,N_25763,N_27441);
and U28581 (N_28581,N_26271,N_25675);
xnor U28582 (N_28582,N_25949,N_25047);
nor U28583 (N_28583,N_26587,N_26130);
or U28584 (N_28584,N_26561,N_27233);
and U28585 (N_28585,N_26557,N_25085);
and U28586 (N_28586,N_25741,N_25359);
nor U28587 (N_28587,N_25013,N_27098);
nor U28588 (N_28588,N_25245,N_26573);
and U28589 (N_28589,N_25382,N_27338);
or U28590 (N_28590,N_25337,N_25398);
nand U28591 (N_28591,N_25647,N_27039);
nor U28592 (N_28592,N_26741,N_25627);
xor U28593 (N_28593,N_26161,N_25580);
xor U28594 (N_28594,N_26685,N_26528);
or U28595 (N_28595,N_25538,N_26804);
nand U28596 (N_28596,N_26615,N_27261);
xor U28597 (N_28597,N_25340,N_25090);
xnor U28598 (N_28598,N_25478,N_26394);
or U28599 (N_28599,N_25648,N_26193);
nand U28600 (N_28600,N_25755,N_26963);
xnor U28601 (N_28601,N_25241,N_25439);
xor U28602 (N_28602,N_26369,N_27196);
nand U28603 (N_28603,N_25781,N_26905);
nor U28604 (N_28604,N_27294,N_27436);
or U28605 (N_28605,N_25154,N_26872);
nor U28606 (N_28606,N_25820,N_26703);
nor U28607 (N_28607,N_25091,N_25353);
or U28608 (N_28608,N_25447,N_25892);
nor U28609 (N_28609,N_26775,N_26263);
and U28610 (N_28610,N_26951,N_25119);
nor U28611 (N_28611,N_25785,N_26746);
xor U28612 (N_28612,N_25667,N_26438);
nand U28613 (N_28613,N_27306,N_27038);
nand U28614 (N_28614,N_26451,N_26821);
and U28615 (N_28615,N_27461,N_26228);
nor U28616 (N_28616,N_27381,N_25209);
nor U28617 (N_28617,N_26892,N_26689);
nor U28618 (N_28618,N_26100,N_26569);
and U28619 (N_28619,N_26939,N_26367);
nor U28620 (N_28620,N_25692,N_26954);
or U28621 (N_28621,N_25854,N_27323);
and U28622 (N_28622,N_26135,N_26215);
and U28623 (N_28623,N_25149,N_27459);
and U28624 (N_28624,N_26289,N_25571);
nand U28625 (N_28625,N_25397,N_25201);
or U28626 (N_28626,N_26448,N_25653);
or U28627 (N_28627,N_26984,N_26265);
xnor U28628 (N_28628,N_25494,N_25143);
or U28629 (N_28629,N_25588,N_25452);
xor U28630 (N_28630,N_27150,N_26489);
nand U28631 (N_28631,N_25812,N_26603);
nor U28632 (N_28632,N_25765,N_26504);
nand U28633 (N_28633,N_25747,N_27145);
xor U28634 (N_28634,N_26177,N_26171);
nor U28635 (N_28635,N_25619,N_25905);
or U28636 (N_28636,N_25551,N_25142);
xnor U28637 (N_28637,N_25380,N_26479);
nor U28638 (N_28638,N_25248,N_25083);
xor U28639 (N_28639,N_26759,N_26781);
or U28640 (N_28640,N_25053,N_26633);
nand U28641 (N_28641,N_25342,N_27201);
nor U28642 (N_28642,N_27198,N_27250);
and U28643 (N_28643,N_25316,N_25577);
or U28644 (N_28644,N_27339,N_27138);
nor U28645 (N_28645,N_25197,N_25932);
xor U28646 (N_28646,N_25093,N_27041);
xor U28647 (N_28647,N_25562,N_27482);
and U28648 (N_28648,N_27054,N_25575);
or U28649 (N_28649,N_25541,N_26026);
nor U28650 (N_28650,N_25772,N_27391);
nand U28651 (N_28651,N_26224,N_26330);
and U28652 (N_28652,N_27021,N_25858);
nand U28653 (N_28653,N_26268,N_26820);
and U28654 (N_28654,N_27238,N_25545);
nor U28655 (N_28655,N_27319,N_25710);
nand U28656 (N_28656,N_26454,N_27053);
and U28657 (N_28657,N_26187,N_27302);
nor U28658 (N_28658,N_25798,N_26218);
nand U28659 (N_28659,N_25865,N_25762);
or U28660 (N_28660,N_26458,N_25583);
and U28661 (N_28661,N_26405,N_26988);
and U28662 (N_28662,N_25081,N_25073);
or U28663 (N_28663,N_25046,N_27132);
nor U28664 (N_28664,N_27083,N_25021);
xor U28665 (N_28665,N_26969,N_26811);
xnor U28666 (N_28666,N_25943,N_26779);
nand U28667 (N_28667,N_27217,N_26110);
xor U28668 (N_28668,N_25624,N_25199);
or U28669 (N_28669,N_26944,N_26117);
and U28670 (N_28670,N_26914,N_27357);
and U28671 (N_28671,N_26614,N_27029);
nor U28672 (N_28672,N_27174,N_25696);
nor U28673 (N_28673,N_26693,N_27172);
xor U28674 (N_28674,N_25768,N_25309);
nor U28675 (N_28675,N_25600,N_25719);
nand U28676 (N_28676,N_26492,N_27031);
nand U28677 (N_28677,N_25928,N_26540);
or U28678 (N_28678,N_27364,N_26258);
nor U28679 (N_28679,N_27179,N_26737);
and U28680 (N_28680,N_26286,N_27300);
and U28681 (N_28681,N_25254,N_26007);
or U28682 (N_28682,N_26000,N_26508);
nor U28683 (N_28683,N_26943,N_27493);
nand U28684 (N_28684,N_26031,N_25597);
nor U28685 (N_28685,N_26787,N_26891);
nor U28686 (N_28686,N_25882,N_25986);
nor U28687 (N_28687,N_26932,N_25564);
or U28688 (N_28688,N_27398,N_26791);
xnor U28689 (N_28689,N_27133,N_25753);
and U28690 (N_28690,N_26067,N_26012);
or U28691 (N_28691,N_25067,N_25799);
nand U28692 (N_28692,N_26992,N_26659);
xnor U28693 (N_28693,N_25092,N_25043);
nand U28694 (N_28694,N_26406,N_25257);
or U28695 (N_28695,N_27353,N_27412);
nor U28696 (N_28696,N_25300,N_25137);
nor U28697 (N_28697,N_25195,N_26552);
nor U28698 (N_28698,N_25177,N_26124);
and U28699 (N_28699,N_25590,N_26747);
or U28700 (N_28700,N_26466,N_25393);
xnor U28701 (N_28701,N_26707,N_25331);
nor U28702 (N_28702,N_25782,N_25437);
nor U28703 (N_28703,N_26143,N_25519);
nor U28704 (N_28704,N_27204,N_26494);
nand U28705 (N_28705,N_26514,N_26929);
and U28706 (N_28706,N_27247,N_25204);
xor U28707 (N_28707,N_27149,N_25644);
nor U28708 (N_28708,N_25413,N_25096);
nand U28709 (N_28709,N_26041,N_27475);
nor U28710 (N_28710,N_25068,N_27103);
xnor U28711 (N_28711,N_26400,N_25087);
nand U28712 (N_28712,N_25811,N_25132);
and U28713 (N_28713,N_26116,N_26119);
nand U28714 (N_28714,N_27350,N_26015);
or U28715 (N_28715,N_27328,N_26923);
nand U28716 (N_28716,N_27084,N_27012);
nand U28717 (N_28717,N_25136,N_26853);
nand U28718 (N_28718,N_27085,N_26588);
and U28719 (N_28719,N_26028,N_27452);
xor U28720 (N_28720,N_27117,N_27311);
and U28721 (N_28721,N_27309,N_26356);
and U28722 (N_28722,N_26794,N_25234);
nand U28723 (N_28723,N_26305,N_25496);
xnor U28724 (N_28724,N_26854,N_25258);
xor U28725 (N_28725,N_26572,N_25210);
nand U28726 (N_28726,N_25481,N_27211);
or U28727 (N_28727,N_25650,N_25664);
and U28728 (N_28728,N_26691,N_26980);
nand U28729 (N_28729,N_27077,N_25576);
nor U28730 (N_28730,N_26777,N_26756);
nand U28731 (N_28731,N_25535,N_25451);
or U28732 (N_28732,N_25740,N_25126);
nor U28733 (N_28733,N_25520,N_25474);
nand U28734 (N_28734,N_25196,N_26884);
and U28735 (N_28735,N_26319,N_26971);
and U28736 (N_28736,N_25709,N_25797);
xnor U28737 (N_28737,N_25796,N_25203);
nand U28738 (N_28738,N_27251,N_27203);
xnor U28739 (N_28739,N_26252,N_25790);
xor U28740 (N_28740,N_26894,N_25850);
nor U28741 (N_28741,N_26098,N_26079);
nor U28742 (N_28742,N_26198,N_25008);
and U28743 (N_28743,N_25427,N_25934);
nor U28744 (N_28744,N_26245,N_25512);
nor U28745 (N_28745,N_26443,N_27480);
and U28746 (N_28746,N_25599,N_25312);
nand U28747 (N_28747,N_25271,N_25361);
or U28748 (N_28748,N_25059,N_26613);
or U28749 (N_28749,N_26729,N_25274);
and U28750 (N_28750,N_26382,N_25738);
nor U28751 (N_28751,N_26763,N_25510);
and U28752 (N_28752,N_25290,N_25475);
and U28753 (N_28753,N_26914,N_26074);
nand U28754 (N_28754,N_25576,N_27068);
nor U28755 (N_28755,N_25829,N_26044);
nand U28756 (N_28756,N_26536,N_25186);
and U28757 (N_28757,N_25594,N_26712);
xor U28758 (N_28758,N_25188,N_25716);
nor U28759 (N_28759,N_27414,N_26283);
and U28760 (N_28760,N_27143,N_26610);
nand U28761 (N_28761,N_26967,N_25162);
nor U28762 (N_28762,N_27302,N_26800);
nand U28763 (N_28763,N_26322,N_25432);
or U28764 (N_28764,N_26920,N_25679);
and U28765 (N_28765,N_26061,N_26783);
nor U28766 (N_28766,N_25970,N_25758);
xnor U28767 (N_28767,N_26195,N_25578);
nand U28768 (N_28768,N_25662,N_26024);
nand U28769 (N_28769,N_27173,N_25952);
or U28770 (N_28770,N_26478,N_26418);
nand U28771 (N_28771,N_26478,N_25197);
nor U28772 (N_28772,N_26940,N_26401);
and U28773 (N_28773,N_27058,N_25282);
nor U28774 (N_28774,N_27216,N_26458);
xnor U28775 (N_28775,N_26402,N_27201);
or U28776 (N_28776,N_25645,N_25910);
nand U28777 (N_28777,N_26257,N_25430);
and U28778 (N_28778,N_25796,N_27490);
nor U28779 (N_28779,N_26496,N_25192);
xor U28780 (N_28780,N_26344,N_25831);
nand U28781 (N_28781,N_25946,N_27055);
nor U28782 (N_28782,N_25530,N_26312);
and U28783 (N_28783,N_27176,N_26281);
nand U28784 (N_28784,N_25943,N_26307);
xor U28785 (N_28785,N_25694,N_26340);
nand U28786 (N_28786,N_26100,N_25594);
or U28787 (N_28787,N_27307,N_26518);
and U28788 (N_28788,N_26318,N_26920);
xor U28789 (N_28789,N_26063,N_25093);
xnor U28790 (N_28790,N_25731,N_26316);
or U28791 (N_28791,N_26642,N_27376);
xnor U28792 (N_28792,N_26111,N_26118);
nor U28793 (N_28793,N_25406,N_26873);
nand U28794 (N_28794,N_27152,N_25707);
or U28795 (N_28795,N_27337,N_27034);
nor U28796 (N_28796,N_25623,N_25819);
nand U28797 (N_28797,N_26181,N_25368);
nor U28798 (N_28798,N_26851,N_26766);
xor U28799 (N_28799,N_27206,N_27020);
and U28800 (N_28800,N_25104,N_27238);
or U28801 (N_28801,N_25460,N_27438);
nand U28802 (N_28802,N_25350,N_27365);
nor U28803 (N_28803,N_26491,N_26264);
nand U28804 (N_28804,N_26389,N_26913);
xor U28805 (N_28805,N_25497,N_25986);
xnor U28806 (N_28806,N_27269,N_25648);
nand U28807 (N_28807,N_26833,N_25608);
nor U28808 (N_28808,N_27360,N_26241);
xnor U28809 (N_28809,N_25222,N_26901);
nor U28810 (N_28810,N_26278,N_26370);
nand U28811 (N_28811,N_27019,N_26923);
nand U28812 (N_28812,N_25947,N_25301);
or U28813 (N_28813,N_27399,N_26235);
and U28814 (N_28814,N_26044,N_25369);
xnor U28815 (N_28815,N_27218,N_25454);
nor U28816 (N_28816,N_25979,N_26852);
xnor U28817 (N_28817,N_26604,N_25824);
and U28818 (N_28818,N_26400,N_27051);
and U28819 (N_28819,N_25271,N_25184);
nor U28820 (N_28820,N_27400,N_26839);
or U28821 (N_28821,N_25129,N_25772);
and U28822 (N_28822,N_27220,N_26023);
or U28823 (N_28823,N_27117,N_25389);
xor U28824 (N_28824,N_26508,N_25402);
and U28825 (N_28825,N_26009,N_26316);
nor U28826 (N_28826,N_25650,N_25412);
xor U28827 (N_28827,N_25612,N_25195);
or U28828 (N_28828,N_25994,N_26449);
xor U28829 (N_28829,N_26424,N_26258);
nor U28830 (N_28830,N_25263,N_26923);
and U28831 (N_28831,N_27024,N_27061);
nor U28832 (N_28832,N_27379,N_27265);
and U28833 (N_28833,N_27052,N_25599);
and U28834 (N_28834,N_27386,N_26259);
and U28835 (N_28835,N_26791,N_26663);
nor U28836 (N_28836,N_25457,N_27126);
nor U28837 (N_28837,N_26236,N_26630);
nor U28838 (N_28838,N_27301,N_26465);
or U28839 (N_28839,N_26095,N_27407);
xnor U28840 (N_28840,N_26978,N_25113);
nand U28841 (N_28841,N_25908,N_27174);
or U28842 (N_28842,N_26795,N_26848);
and U28843 (N_28843,N_25872,N_26527);
or U28844 (N_28844,N_26757,N_26776);
nor U28845 (N_28845,N_26784,N_26518);
nor U28846 (N_28846,N_25686,N_25941);
xor U28847 (N_28847,N_25613,N_26064);
and U28848 (N_28848,N_25375,N_25871);
nor U28849 (N_28849,N_25031,N_26382);
or U28850 (N_28850,N_26149,N_26521);
and U28851 (N_28851,N_26815,N_26452);
and U28852 (N_28852,N_27058,N_25443);
nor U28853 (N_28853,N_26090,N_25169);
or U28854 (N_28854,N_26882,N_25181);
and U28855 (N_28855,N_27439,N_26604);
nand U28856 (N_28856,N_26019,N_27409);
and U28857 (N_28857,N_25488,N_26177);
and U28858 (N_28858,N_26212,N_26983);
nor U28859 (N_28859,N_26282,N_27338);
xnor U28860 (N_28860,N_25562,N_26458);
nand U28861 (N_28861,N_27142,N_25611);
nand U28862 (N_28862,N_25720,N_26660);
nand U28863 (N_28863,N_26607,N_25341);
xor U28864 (N_28864,N_26113,N_26024);
or U28865 (N_28865,N_26297,N_26566);
xor U28866 (N_28866,N_27035,N_25070);
and U28867 (N_28867,N_26961,N_26296);
xor U28868 (N_28868,N_26216,N_26226);
nand U28869 (N_28869,N_25850,N_26613);
nand U28870 (N_28870,N_25179,N_26204);
nor U28871 (N_28871,N_27096,N_27213);
nand U28872 (N_28872,N_25617,N_25894);
nand U28873 (N_28873,N_26118,N_26781);
and U28874 (N_28874,N_26480,N_26932);
nand U28875 (N_28875,N_27236,N_25576);
or U28876 (N_28876,N_27280,N_26807);
nor U28877 (N_28877,N_25083,N_26793);
nor U28878 (N_28878,N_26765,N_25781);
xnor U28879 (N_28879,N_26888,N_25602);
xor U28880 (N_28880,N_25520,N_27480);
or U28881 (N_28881,N_25568,N_25395);
and U28882 (N_28882,N_27484,N_25873);
xnor U28883 (N_28883,N_26219,N_26406);
nand U28884 (N_28884,N_26430,N_25893);
or U28885 (N_28885,N_26389,N_25838);
or U28886 (N_28886,N_27099,N_26661);
and U28887 (N_28887,N_27220,N_25780);
xnor U28888 (N_28888,N_26607,N_26469);
nand U28889 (N_28889,N_26166,N_26248);
xor U28890 (N_28890,N_26764,N_25146);
nand U28891 (N_28891,N_26181,N_25686);
nand U28892 (N_28892,N_26210,N_25942);
nand U28893 (N_28893,N_26981,N_27086);
and U28894 (N_28894,N_25952,N_26464);
and U28895 (N_28895,N_26891,N_25312);
and U28896 (N_28896,N_25151,N_25879);
or U28897 (N_28897,N_25377,N_26309);
nor U28898 (N_28898,N_25347,N_25769);
and U28899 (N_28899,N_26973,N_26865);
xor U28900 (N_28900,N_25252,N_25683);
or U28901 (N_28901,N_26990,N_25164);
xnor U28902 (N_28902,N_26625,N_25863);
and U28903 (N_28903,N_26338,N_25831);
xor U28904 (N_28904,N_27211,N_25111);
or U28905 (N_28905,N_26889,N_26236);
xor U28906 (N_28906,N_26274,N_25858);
nor U28907 (N_28907,N_25002,N_27251);
nor U28908 (N_28908,N_26792,N_26823);
or U28909 (N_28909,N_25696,N_26348);
xnor U28910 (N_28910,N_27495,N_25725);
nand U28911 (N_28911,N_25402,N_25504);
xnor U28912 (N_28912,N_27175,N_27043);
xnor U28913 (N_28913,N_26702,N_26555);
and U28914 (N_28914,N_25437,N_26638);
and U28915 (N_28915,N_26038,N_25867);
nand U28916 (N_28916,N_26671,N_27144);
xnor U28917 (N_28917,N_26551,N_25571);
or U28918 (N_28918,N_27399,N_25575);
nand U28919 (N_28919,N_26487,N_25042);
nor U28920 (N_28920,N_26034,N_25684);
and U28921 (N_28921,N_26651,N_27081);
nand U28922 (N_28922,N_27152,N_27417);
xnor U28923 (N_28923,N_27236,N_26302);
nand U28924 (N_28924,N_27295,N_25074);
or U28925 (N_28925,N_26644,N_26050);
nand U28926 (N_28926,N_25311,N_27058);
or U28927 (N_28927,N_27354,N_25161);
nor U28928 (N_28928,N_26074,N_26359);
nor U28929 (N_28929,N_26789,N_25910);
nor U28930 (N_28930,N_25824,N_25204);
nor U28931 (N_28931,N_25753,N_27374);
nand U28932 (N_28932,N_26301,N_26284);
or U28933 (N_28933,N_26308,N_26670);
and U28934 (N_28934,N_26416,N_25465);
nand U28935 (N_28935,N_25131,N_26661);
nand U28936 (N_28936,N_26487,N_27257);
and U28937 (N_28937,N_26017,N_26487);
or U28938 (N_28938,N_27175,N_26427);
xnor U28939 (N_28939,N_27185,N_25761);
and U28940 (N_28940,N_27468,N_25342);
xnor U28941 (N_28941,N_25944,N_25873);
and U28942 (N_28942,N_27348,N_26391);
nand U28943 (N_28943,N_26473,N_26154);
xor U28944 (N_28944,N_27247,N_25893);
or U28945 (N_28945,N_27117,N_27163);
nand U28946 (N_28946,N_26268,N_26290);
nor U28947 (N_28947,N_25411,N_25679);
nand U28948 (N_28948,N_25914,N_25994);
xor U28949 (N_28949,N_25084,N_26912);
nand U28950 (N_28950,N_25762,N_26197);
nor U28951 (N_28951,N_27290,N_26674);
nor U28952 (N_28952,N_25673,N_25329);
nor U28953 (N_28953,N_26564,N_26507);
and U28954 (N_28954,N_26317,N_27079);
nor U28955 (N_28955,N_25120,N_26955);
nand U28956 (N_28956,N_25754,N_27288);
nand U28957 (N_28957,N_25971,N_26651);
xnor U28958 (N_28958,N_27057,N_27013);
nor U28959 (N_28959,N_25299,N_25482);
or U28960 (N_28960,N_27187,N_25950);
xnor U28961 (N_28961,N_25785,N_25833);
nor U28962 (N_28962,N_27190,N_27412);
nor U28963 (N_28963,N_27077,N_26475);
and U28964 (N_28964,N_25221,N_25766);
nor U28965 (N_28965,N_27035,N_26809);
xor U28966 (N_28966,N_27339,N_26141);
and U28967 (N_28967,N_27082,N_25657);
nor U28968 (N_28968,N_25965,N_26030);
or U28969 (N_28969,N_26703,N_25136);
nand U28970 (N_28970,N_27213,N_25123);
nand U28971 (N_28971,N_26523,N_25795);
nand U28972 (N_28972,N_26475,N_26859);
xnor U28973 (N_28973,N_27172,N_26722);
and U28974 (N_28974,N_26323,N_27478);
nand U28975 (N_28975,N_25648,N_25104);
nand U28976 (N_28976,N_26954,N_26380);
nor U28977 (N_28977,N_26177,N_25439);
or U28978 (N_28978,N_26148,N_26327);
nand U28979 (N_28979,N_25040,N_26230);
or U28980 (N_28980,N_27180,N_25451);
and U28981 (N_28981,N_25776,N_26282);
or U28982 (N_28982,N_26140,N_26422);
nor U28983 (N_28983,N_26216,N_26368);
and U28984 (N_28984,N_25670,N_25869);
nand U28985 (N_28985,N_25247,N_25896);
nand U28986 (N_28986,N_26044,N_25576);
nor U28987 (N_28987,N_26793,N_26097);
nor U28988 (N_28988,N_25812,N_26040);
and U28989 (N_28989,N_25547,N_27367);
xor U28990 (N_28990,N_25280,N_25663);
xor U28991 (N_28991,N_25760,N_26698);
nand U28992 (N_28992,N_25628,N_25721);
xor U28993 (N_28993,N_26994,N_27062);
nor U28994 (N_28994,N_27022,N_25489);
nand U28995 (N_28995,N_25696,N_26374);
nor U28996 (N_28996,N_25022,N_25451);
and U28997 (N_28997,N_25840,N_26413);
and U28998 (N_28998,N_25135,N_26010);
and U28999 (N_28999,N_26560,N_27231);
nand U29000 (N_29000,N_27477,N_27444);
and U29001 (N_29001,N_26737,N_25072);
xnor U29002 (N_29002,N_27162,N_26986);
nand U29003 (N_29003,N_25296,N_26942);
nand U29004 (N_29004,N_26465,N_26143);
and U29005 (N_29005,N_27047,N_26904);
nor U29006 (N_29006,N_25861,N_25811);
xor U29007 (N_29007,N_25589,N_26401);
and U29008 (N_29008,N_27041,N_25954);
nand U29009 (N_29009,N_25022,N_25389);
nand U29010 (N_29010,N_25016,N_25662);
nand U29011 (N_29011,N_26383,N_27065);
nand U29012 (N_29012,N_27181,N_26529);
nand U29013 (N_29013,N_26645,N_25408);
and U29014 (N_29014,N_27068,N_27492);
nor U29015 (N_29015,N_25070,N_25160);
and U29016 (N_29016,N_26206,N_26916);
or U29017 (N_29017,N_25861,N_25233);
and U29018 (N_29018,N_25577,N_25526);
and U29019 (N_29019,N_25485,N_26270);
nor U29020 (N_29020,N_27347,N_26141);
xor U29021 (N_29021,N_25016,N_25594);
and U29022 (N_29022,N_25400,N_26496);
nand U29023 (N_29023,N_27381,N_25002);
nor U29024 (N_29024,N_26925,N_26013);
xor U29025 (N_29025,N_25874,N_25398);
xor U29026 (N_29026,N_25775,N_26521);
nor U29027 (N_29027,N_25337,N_26301);
and U29028 (N_29028,N_25046,N_27185);
nor U29029 (N_29029,N_26121,N_25299);
xnor U29030 (N_29030,N_26637,N_25347);
nor U29031 (N_29031,N_27427,N_27193);
xor U29032 (N_29032,N_25742,N_26118);
nand U29033 (N_29033,N_25637,N_26484);
nand U29034 (N_29034,N_27180,N_25052);
or U29035 (N_29035,N_25018,N_27335);
nand U29036 (N_29036,N_26327,N_25555);
or U29037 (N_29037,N_25195,N_25148);
and U29038 (N_29038,N_25790,N_25003);
or U29039 (N_29039,N_25529,N_26592);
and U29040 (N_29040,N_25434,N_27403);
and U29041 (N_29041,N_25598,N_27258);
nor U29042 (N_29042,N_27156,N_26299);
nor U29043 (N_29043,N_26860,N_25028);
or U29044 (N_29044,N_27385,N_25700);
xnor U29045 (N_29045,N_25706,N_26448);
or U29046 (N_29046,N_25143,N_27456);
nor U29047 (N_29047,N_27497,N_26377);
or U29048 (N_29048,N_27300,N_27125);
xor U29049 (N_29049,N_25851,N_26928);
and U29050 (N_29050,N_26859,N_26771);
and U29051 (N_29051,N_25579,N_27220);
or U29052 (N_29052,N_26403,N_25315);
or U29053 (N_29053,N_25700,N_26051);
nand U29054 (N_29054,N_27105,N_26563);
nor U29055 (N_29055,N_27274,N_26376);
or U29056 (N_29056,N_25910,N_25849);
nor U29057 (N_29057,N_25379,N_26302);
or U29058 (N_29058,N_26014,N_25629);
xnor U29059 (N_29059,N_26067,N_25256);
or U29060 (N_29060,N_25801,N_25095);
nand U29061 (N_29061,N_25222,N_27251);
and U29062 (N_29062,N_27182,N_27491);
nor U29063 (N_29063,N_25756,N_25787);
nor U29064 (N_29064,N_26214,N_26370);
or U29065 (N_29065,N_27231,N_25851);
xor U29066 (N_29066,N_26730,N_26812);
nand U29067 (N_29067,N_25281,N_25614);
and U29068 (N_29068,N_25555,N_26434);
nor U29069 (N_29069,N_25785,N_26859);
xor U29070 (N_29070,N_25411,N_27090);
nand U29071 (N_29071,N_27095,N_25383);
or U29072 (N_29072,N_25815,N_25803);
nor U29073 (N_29073,N_27311,N_25842);
xor U29074 (N_29074,N_26345,N_27080);
or U29075 (N_29075,N_26648,N_27158);
or U29076 (N_29076,N_25564,N_25257);
nor U29077 (N_29077,N_26591,N_25679);
and U29078 (N_29078,N_25642,N_26225);
nand U29079 (N_29079,N_27002,N_25872);
or U29080 (N_29080,N_25284,N_25069);
xnor U29081 (N_29081,N_25459,N_25118);
xor U29082 (N_29082,N_26126,N_25443);
or U29083 (N_29083,N_26246,N_25276);
nor U29084 (N_29084,N_26439,N_26219);
xor U29085 (N_29085,N_25870,N_27062);
xnor U29086 (N_29086,N_26532,N_27071);
nand U29087 (N_29087,N_27437,N_26200);
nand U29088 (N_29088,N_25818,N_26801);
nor U29089 (N_29089,N_25356,N_25628);
or U29090 (N_29090,N_27258,N_25821);
nor U29091 (N_29091,N_25651,N_26163);
or U29092 (N_29092,N_26769,N_25386);
and U29093 (N_29093,N_26429,N_27238);
nand U29094 (N_29094,N_27239,N_25890);
xnor U29095 (N_29095,N_25089,N_25399);
and U29096 (N_29096,N_25502,N_26800);
or U29097 (N_29097,N_25754,N_25134);
nand U29098 (N_29098,N_26554,N_26902);
xor U29099 (N_29099,N_25905,N_26010);
nor U29100 (N_29100,N_27169,N_27095);
and U29101 (N_29101,N_26759,N_25945);
and U29102 (N_29102,N_25210,N_26605);
xor U29103 (N_29103,N_27321,N_26532);
nor U29104 (N_29104,N_26330,N_26051);
or U29105 (N_29105,N_25563,N_25438);
nor U29106 (N_29106,N_26434,N_26190);
and U29107 (N_29107,N_25827,N_25759);
nand U29108 (N_29108,N_26557,N_25586);
nand U29109 (N_29109,N_25237,N_25338);
xor U29110 (N_29110,N_25837,N_25523);
or U29111 (N_29111,N_27421,N_25279);
nor U29112 (N_29112,N_25280,N_27296);
xor U29113 (N_29113,N_27257,N_26068);
and U29114 (N_29114,N_25918,N_25485);
nor U29115 (N_29115,N_26797,N_26071);
nor U29116 (N_29116,N_27277,N_26104);
nor U29117 (N_29117,N_27282,N_27462);
and U29118 (N_29118,N_26025,N_26116);
nand U29119 (N_29119,N_25607,N_25554);
xor U29120 (N_29120,N_25398,N_27142);
or U29121 (N_29121,N_26059,N_26261);
xor U29122 (N_29122,N_25254,N_26837);
nand U29123 (N_29123,N_25485,N_26189);
or U29124 (N_29124,N_27308,N_26206);
nor U29125 (N_29125,N_27370,N_26491);
or U29126 (N_29126,N_25672,N_27020);
nor U29127 (N_29127,N_25490,N_26441);
nand U29128 (N_29128,N_25172,N_26831);
xnor U29129 (N_29129,N_26490,N_26518);
xnor U29130 (N_29130,N_26914,N_26406);
and U29131 (N_29131,N_26035,N_26786);
xor U29132 (N_29132,N_26561,N_25836);
and U29133 (N_29133,N_26732,N_27293);
nand U29134 (N_29134,N_25934,N_26830);
and U29135 (N_29135,N_25219,N_27443);
and U29136 (N_29136,N_27109,N_25751);
xnor U29137 (N_29137,N_25600,N_26886);
xnor U29138 (N_29138,N_25226,N_26831);
xnor U29139 (N_29139,N_25758,N_26413);
nand U29140 (N_29140,N_25734,N_25793);
nand U29141 (N_29141,N_25773,N_27467);
nand U29142 (N_29142,N_26870,N_26199);
nand U29143 (N_29143,N_25560,N_25739);
nor U29144 (N_29144,N_25258,N_27283);
xor U29145 (N_29145,N_25549,N_27478);
nand U29146 (N_29146,N_26358,N_27389);
xnor U29147 (N_29147,N_27018,N_25088);
xor U29148 (N_29148,N_25654,N_25491);
xor U29149 (N_29149,N_25062,N_25677);
or U29150 (N_29150,N_27384,N_25894);
nand U29151 (N_29151,N_25398,N_26431);
and U29152 (N_29152,N_26799,N_27139);
nor U29153 (N_29153,N_26122,N_26642);
and U29154 (N_29154,N_26726,N_25762);
nor U29155 (N_29155,N_25499,N_26237);
or U29156 (N_29156,N_26717,N_25485);
xor U29157 (N_29157,N_25498,N_27238);
nor U29158 (N_29158,N_25845,N_26142);
or U29159 (N_29159,N_27293,N_25124);
and U29160 (N_29160,N_25230,N_26736);
xor U29161 (N_29161,N_25487,N_27309);
or U29162 (N_29162,N_25749,N_25398);
nand U29163 (N_29163,N_26050,N_27234);
xor U29164 (N_29164,N_26354,N_27171);
nand U29165 (N_29165,N_25683,N_25559);
nand U29166 (N_29166,N_27394,N_25431);
nand U29167 (N_29167,N_25161,N_25800);
xnor U29168 (N_29168,N_27021,N_25899);
nor U29169 (N_29169,N_25919,N_27265);
or U29170 (N_29170,N_26557,N_27271);
and U29171 (N_29171,N_25761,N_26974);
and U29172 (N_29172,N_25431,N_26310);
and U29173 (N_29173,N_26464,N_25378);
nand U29174 (N_29174,N_26931,N_26647);
and U29175 (N_29175,N_26292,N_26090);
nor U29176 (N_29176,N_25351,N_26789);
and U29177 (N_29177,N_27013,N_25535);
xor U29178 (N_29178,N_27125,N_26722);
xor U29179 (N_29179,N_27434,N_25505);
xor U29180 (N_29180,N_25367,N_26123);
nor U29181 (N_29181,N_26289,N_25835);
and U29182 (N_29182,N_26119,N_25003);
nand U29183 (N_29183,N_25558,N_25636);
nor U29184 (N_29184,N_25672,N_26197);
nor U29185 (N_29185,N_25687,N_25117);
xnor U29186 (N_29186,N_25955,N_25437);
nand U29187 (N_29187,N_26614,N_26717);
nand U29188 (N_29188,N_26108,N_25777);
nor U29189 (N_29189,N_26559,N_27044);
or U29190 (N_29190,N_27413,N_26115);
or U29191 (N_29191,N_25280,N_26238);
xnor U29192 (N_29192,N_26300,N_26530);
nor U29193 (N_29193,N_27444,N_25094);
nand U29194 (N_29194,N_25437,N_26670);
nor U29195 (N_29195,N_25529,N_26596);
nand U29196 (N_29196,N_26653,N_26381);
and U29197 (N_29197,N_25046,N_26966);
nor U29198 (N_29198,N_26640,N_25911);
nor U29199 (N_29199,N_25635,N_26932);
and U29200 (N_29200,N_25976,N_25190);
xor U29201 (N_29201,N_25433,N_26454);
nand U29202 (N_29202,N_25300,N_26664);
nor U29203 (N_29203,N_26578,N_25591);
nor U29204 (N_29204,N_26106,N_26997);
nand U29205 (N_29205,N_25240,N_25878);
nor U29206 (N_29206,N_26802,N_26941);
or U29207 (N_29207,N_26048,N_27118);
xnor U29208 (N_29208,N_25202,N_26322);
and U29209 (N_29209,N_25458,N_26692);
nor U29210 (N_29210,N_26225,N_27079);
and U29211 (N_29211,N_25627,N_27368);
and U29212 (N_29212,N_26744,N_26581);
xor U29213 (N_29213,N_27129,N_25697);
nor U29214 (N_29214,N_27389,N_25225);
and U29215 (N_29215,N_25529,N_25568);
or U29216 (N_29216,N_27248,N_25377);
nand U29217 (N_29217,N_26217,N_25421);
nor U29218 (N_29218,N_26264,N_26354);
xor U29219 (N_29219,N_26429,N_26129);
xor U29220 (N_29220,N_27187,N_26073);
xor U29221 (N_29221,N_26247,N_25080);
nor U29222 (N_29222,N_25378,N_27166);
or U29223 (N_29223,N_26794,N_27464);
nor U29224 (N_29224,N_26166,N_26192);
or U29225 (N_29225,N_25971,N_27118);
and U29226 (N_29226,N_25650,N_26267);
nand U29227 (N_29227,N_25962,N_26302);
and U29228 (N_29228,N_26848,N_27273);
and U29229 (N_29229,N_26692,N_25501);
xor U29230 (N_29230,N_25340,N_25581);
nor U29231 (N_29231,N_26567,N_27454);
nor U29232 (N_29232,N_27380,N_25242);
and U29233 (N_29233,N_25245,N_25659);
xor U29234 (N_29234,N_25400,N_26397);
nand U29235 (N_29235,N_25592,N_26627);
nor U29236 (N_29236,N_27398,N_27146);
or U29237 (N_29237,N_25259,N_26841);
nand U29238 (N_29238,N_27077,N_25371);
or U29239 (N_29239,N_25282,N_25905);
nand U29240 (N_29240,N_26329,N_25075);
nor U29241 (N_29241,N_25312,N_25774);
and U29242 (N_29242,N_26985,N_26930);
or U29243 (N_29243,N_25028,N_25217);
or U29244 (N_29244,N_27023,N_27177);
xor U29245 (N_29245,N_25660,N_26033);
and U29246 (N_29246,N_27215,N_26703);
nand U29247 (N_29247,N_27019,N_26986);
nor U29248 (N_29248,N_26075,N_27306);
nor U29249 (N_29249,N_26294,N_25375);
or U29250 (N_29250,N_25469,N_25313);
nor U29251 (N_29251,N_27197,N_25404);
nor U29252 (N_29252,N_25133,N_25891);
nor U29253 (N_29253,N_25555,N_26078);
and U29254 (N_29254,N_26529,N_26349);
nor U29255 (N_29255,N_26321,N_26257);
nor U29256 (N_29256,N_26791,N_25489);
or U29257 (N_29257,N_25973,N_26820);
or U29258 (N_29258,N_27371,N_25895);
and U29259 (N_29259,N_26100,N_25425);
nor U29260 (N_29260,N_25665,N_26960);
or U29261 (N_29261,N_26628,N_26904);
xnor U29262 (N_29262,N_27194,N_26557);
nand U29263 (N_29263,N_27279,N_25316);
xnor U29264 (N_29264,N_26520,N_26003);
and U29265 (N_29265,N_25172,N_26953);
nand U29266 (N_29266,N_26961,N_26716);
nand U29267 (N_29267,N_26309,N_26017);
nor U29268 (N_29268,N_27081,N_25951);
nor U29269 (N_29269,N_25937,N_27246);
and U29270 (N_29270,N_26300,N_26203);
xor U29271 (N_29271,N_25053,N_27439);
nor U29272 (N_29272,N_25164,N_27343);
or U29273 (N_29273,N_26367,N_26625);
nand U29274 (N_29274,N_25921,N_26433);
xnor U29275 (N_29275,N_27359,N_25111);
and U29276 (N_29276,N_27116,N_27445);
xnor U29277 (N_29277,N_26737,N_26611);
nor U29278 (N_29278,N_25607,N_27431);
or U29279 (N_29279,N_27348,N_25865);
xnor U29280 (N_29280,N_26877,N_25800);
nor U29281 (N_29281,N_25453,N_25428);
and U29282 (N_29282,N_26092,N_27375);
nand U29283 (N_29283,N_25420,N_26495);
and U29284 (N_29284,N_27296,N_26108);
xor U29285 (N_29285,N_25571,N_25857);
and U29286 (N_29286,N_27124,N_26317);
xor U29287 (N_29287,N_26456,N_25442);
xor U29288 (N_29288,N_25238,N_26025);
xnor U29289 (N_29289,N_25384,N_25985);
or U29290 (N_29290,N_26478,N_25768);
nor U29291 (N_29291,N_25798,N_27371);
or U29292 (N_29292,N_26874,N_25717);
and U29293 (N_29293,N_26221,N_27412);
xnor U29294 (N_29294,N_26753,N_26195);
and U29295 (N_29295,N_27168,N_25240);
and U29296 (N_29296,N_26113,N_25994);
and U29297 (N_29297,N_25713,N_26898);
xor U29298 (N_29298,N_26570,N_25178);
nand U29299 (N_29299,N_27488,N_25538);
or U29300 (N_29300,N_27261,N_27428);
nor U29301 (N_29301,N_27197,N_26923);
or U29302 (N_29302,N_26516,N_25033);
nor U29303 (N_29303,N_25757,N_26816);
nor U29304 (N_29304,N_26212,N_26845);
nand U29305 (N_29305,N_26336,N_25264);
and U29306 (N_29306,N_26288,N_25697);
nand U29307 (N_29307,N_26839,N_27305);
or U29308 (N_29308,N_25788,N_25049);
or U29309 (N_29309,N_26674,N_27167);
nand U29310 (N_29310,N_26918,N_26739);
nand U29311 (N_29311,N_26523,N_26894);
nor U29312 (N_29312,N_26945,N_26356);
and U29313 (N_29313,N_25657,N_25897);
or U29314 (N_29314,N_25163,N_27354);
or U29315 (N_29315,N_25335,N_26174);
and U29316 (N_29316,N_25752,N_25229);
xnor U29317 (N_29317,N_26000,N_25563);
nor U29318 (N_29318,N_27094,N_25170);
and U29319 (N_29319,N_25174,N_27058);
xor U29320 (N_29320,N_25232,N_25122);
nand U29321 (N_29321,N_27253,N_27116);
nor U29322 (N_29322,N_26018,N_27319);
nor U29323 (N_29323,N_26462,N_26791);
nor U29324 (N_29324,N_26411,N_26723);
nor U29325 (N_29325,N_25821,N_26990);
and U29326 (N_29326,N_26363,N_25101);
and U29327 (N_29327,N_25666,N_26987);
and U29328 (N_29328,N_25794,N_26525);
or U29329 (N_29329,N_25331,N_26298);
nor U29330 (N_29330,N_26571,N_25837);
xnor U29331 (N_29331,N_26536,N_25800);
nand U29332 (N_29332,N_25044,N_27442);
nand U29333 (N_29333,N_27384,N_27491);
nand U29334 (N_29334,N_25800,N_27288);
nor U29335 (N_29335,N_25191,N_25517);
and U29336 (N_29336,N_27392,N_27346);
nand U29337 (N_29337,N_26197,N_25354);
and U29338 (N_29338,N_25598,N_26295);
or U29339 (N_29339,N_26756,N_25019);
nand U29340 (N_29340,N_25052,N_27124);
nor U29341 (N_29341,N_25228,N_27259);
nand U29342 (N_29342,N_26452,N_26496);
nor U29343 (N_29343,N_25127,N_25895);
or U29344 (N_29344,N_25196,N_27161);
and U29345 (N_29345,N_25836,N_25849);
or U29346 (N_29346,N_25287,N_26624);
or U29347 (N_29347,N_26097,N_25949);
nor U29348 (N_29348,N_27449,N_27097);
or U29349 (N_29349,N_25041,N_26222);
xor U29350 (N_29350,N_25510,N_25466);
nor U29351 (N_29351,N_27143,N_26248);
xor U29352 (N_29352,N_26271,N_27417);
xor U29353 (N_29353,N_26056,N_26968);
and U29354 (N_29354,N_26938,N_26263);
and U29355 (N_29355,N_26599,N_27193);
xnor U29356 (N_29356,N_25283,N_27421);
or U29357 (N_29357,N_25549,N_26903);
nand U29358 (N_29358,N_26896,N_25290);
or U29359 (N_29359,N_26804,N_26248);
nand U29360 (N_29360,N_27451,N_26560);
xnor U29361 (N_29361,N_26600,N_25308);
nor U29362 (N_29362,N_25024,N_26928);
or U29363 (N_29363,N_26723,N_26580);
and U29364 (N_29364,N_26327,N_25275);
nor U29365 (N_29365,N_27354,N_25221);
or U29366 (N_29366,N_26877,N_27184);
or U29367 (N_29367,N_25622,N_25612);
and U29368 (N_29368,N_27159,N_26049);
nand U29369 (N_29369,N_25869,N_26132);
or U29370 (N_29370,N_27348,N_25804);
xnor U29371 (N_29371,N_26958,N_25185);
and U29372 (N_29372,N_25438,N_25576);
nor U29373 (N_29373,N_25390,N_25784);
nor U29374 (N_29374,N_25289,N_26396);
xor U29375 (N_29375,N_26219,N_26771);
nand U29376 (N_29376,N_27251,N_26127);
and U29377 (N_29377,N_26420,N_25471);
and U29378 (N_29378,N_25105,N_25540);
and U29379 (N_29379,N_25986,N_27175);
xnor U29380 (N_29380,N_27041,N_25583);
nand U29381 (N_29381,N_25124,N_25634);
or U29382 (N_29382,N_25605,N_26733);
and U29383 (N_29383,N_25005,N_25028);
or U29384 (N_29384,N_27301,N_26068);
nand U29385 (N_29385,N_25232,N_26567);
nand U29386 (N_29386,N_26648,N_25477);
nor U29387 (N_29387,N_26082,N_25865);
nor U29388 (N_29388,N_26653,N_25896);
nor U29389 (N_29389,N_26293,N_26701);
xnor U29390 (N_29390,N_26660,N_25467);
nor U29391 (N_29391,N_26311,N_26070);
and U29392 (N_29392,N_27493,N_25878);
xnor U29393 (N_29393,N_26988,N_25506);
and U29394 (N_29394,N_25014,N_25271);
and U29395 (N_29395,N_25233,N_27258);
xor U29396 (N_29396,N_27165,N_26690);
nand U29397 (N_29397,N_25075,N_26415);
nand U29398 (N_29398,N_25798,N_25537);
and U29399 (N_29399,N_25630,N_27416);
nand U29400 (N_29400,N_27176,N_26891);
nor U29401 (N_29401,N_26669,N_26109);
and U29402 (N_29402,N_26608,N_25093);
nor U29403 (N_29403,N_26013,N_27161);
nand U29404 (N_29404,N_26230,N_25501);
xor U29405 (N_29405,N_25672,N_27250);
nor U29406 (N_29406,N_25411,N_25756);
or U29407 (N_29407,N_25276,N_25686);
nand U29408 (N_29408,N_27218,N_26573);
nand U29409 (N_29409,N_26999,N_26331);
nor U29410 (N_29410,N_26531,N_25077);
and U29411 (N_29411,N_25385,N_26720);
or U29412 (N_29412,N_25520,N_26603);
and U29413 (N_29413,N_26361,N_25485);
nand U29414 (N_29414,N_25684,N_25918);
xnor U29415 (N_29415,N_26926,N_26810);
nor U29416 (N_29416,N_25491,N_26865);
nor U29417 (N_29417,N_26430,N_25666);
xor U29418 (N_29418,N_25894,N_26126);
xor U29419 (N_29419,N_26812,N_26111);
nand U29420 (N_29420,N_27235,N_26004);
nor U29421 (N_29421,N_25003,N_27161);
and U29422 (N_29422,N_27267,N_27308);
or U29423 (N_29423,N_26451,N_27255);
and U29424 (N_29424,N_27453,N_25899);
nand U29425 (N_29425,N_26041,N_26030);
or U29426 (N_29426,N_26158,N_26041);
or U29427 (N_29427,N_26345,N_25914);
or U29428 (N_29428,N_26185,N_25975);
xnor U29429 (N_29429,N_25314,N_25410);
or U29430 (N_29430,N_25390,N_25719);
nor U29431 (N_29431,N_25857,N_26957);
xnor U29432 (N_29432,N_26240,N_27125);
nor U29433 (N_29433,N_26941,N_27364);
and U29434 (N_29434,N_25589,N_25421);
nor U29435 (N_29435,N_26678,N_26782);
nand U29436 (N_29436,N_26562,N_27040);
xnor U29437 (N_29437,N_27066,N_26380);
or U29438 (N_29438,N_26156,N_25835);
xor U29439 (N_29439,N_26149,N_26794);
or U29440 (N_29440,N_26196,N_26987);
nor U29441 (N_29441,N_27323,N_26495);
and U29442 (N_29442,N_26491,N_25967);
and U29443 (N_29443,N_25921,N_25099);
and U29444 (N_29444,N_26607,N_26928);
nor U29445 (N_29445,N_26061,N_25153);
or U29446 (N_29446,N_26116,N_26730);
or U29447 (N_29447,N_25718,N_27232);
or U29448 (N_29448,N_27449,N_26915);
or U29449 (N_29449,N_25059,N_25210);
and U29450 (N_29450,N_27004,N_27082);
nor U29451 (N_29451,N_26728,N_26675);
nor U29452 (N_29452,N_27305,N_25681);
nand U29453 (N_29453,N_25956,N_27206);
xor U29454 (N_29454,N_26902,N_25679);
nand U29455 (N_29455,N_26713,N_25424);
xnor U29456 (N_29456,N_26522,N_25175);
or U29457 (N_29457,N_27442,N_26405);
nand U29458 (N_29458,N_26946,N_26595);
nor U29459 (N_29459,N_25737,N_27336);
and U29460 (N_29460,N_26244,N_26891);
nand U29461 (N_29461,N_27415,N_27450);
xor U29462 (N_29462,N_27264,N_26855);
nand U29463 (N_29463,N_26256,N_26725);
nand U29464 (N_29464,N_26789,N_26668);
nand U29465 (N_29465,N_27359,N_26667);
xor U29466 (N_29466,N_25378,N_27049);
xor U29467 (N_29467,N_26479,N_25393);
and U29468 (N_29468,N_26108,N_26633);
xnor U29469 (N_29469,N_26281,N_25057);
nand U29470 (N_29470,N_25716,N_26022);
and U29471 (N_29471,N_26452,N_25346);
and U29472 (N_29472,N_26985,N_25330);
xor U29473 (N_29473,N_25751,N_26421);
xnor U29474 (N_29474,N_26416,N_26380);
nand U29475 (N_29475,N_26007,N_26166);
or U29476 (N_29476,N_25062,N_25252);
or U29477 (N_29477,N_25536,N_25390);
xor U29478 (N_29478,N_25665,N_27119);
or U29479 (N_29479,N_27378,N_25653);
nand U29480 (N_29480,N_27376,N_25521);
and U29481 (N_29481,N_26479,N_25296);
nor U29482 (N_29482,N_26975,N_26433);
nor U29483 (N_29483,N_25884,N_26924);
or U29484 (N_29484,N_26570,N_25661);
nand U29485 (N_29485,N_25649,N_26295);
nor U29486 (N_29486,N_27271,N_26934);
nand U29487 (N_29487,N_25509,N_26169);
xor U29488 (N_29488,N_26973,N_27491);
xnor U29489 (N_29489,N_25341,N_26569);
nand U29490 (N_29490,N_27244,N_25857);
nor U29491 (N_29491,N_25345,N_27029);
nor U29492 (N_29492,N_27122,N_25799);
nand U29493 (N_29493,N_26431,N_25526);
xor U29494 (N_29494,N_26509,N_25848);
xnor U29495 (N_29495,N_26323,N_25730);
and U29496 (N_29496,N_25134,N_27426);
nor U29497 (N_29497,N_25516,N_26598);
xnor U29498 (N_29498,N_27336,N_26590);
nand U29499 (N_29499,N_25494,N_26915);
and U29500 (N_29500,N_26700,N_26063);
nor U29501 (N_29501,N_26625,N_26863);
or U29502 (N_29502,N_26135,N_27276);
nor U29503 (N_29503,N_26302,N_26753);
or U29504 (N_29504,N_25005,N_25023);
and U29505 (N_29505,N_25811,N_27028);
or U29506 (N_29506,N_26642,N_25729);
and U29507 (N_29507,N_26049,N_27147);
or U29508 (N_29508,N_25715,N_27148);
and U29509 (N_29509,N_26259,N_27146);
and U29510 (N_29510,N_26263,N_27032);
nand U29511 (N_29511,N_27349,N_26485);
or U29512 (N_29512,N_25923,N_25362);
and U29513 (N_29513,N_25922,N_27299);
or U29514 (N_29514,N_25327,N_26447);
nand U29515 (N_29515,N_26970,N_26003);
nand U29516 (N_29516,N_25111,N_27414);
nor U29517 (N_29517,N_26609,N_25952);
and U29518 (N_29518,N_27383,N_25321);
nand U29519 (N_29519,N_26642,N_25632);
or U29520 (N_29520,N_27131,N_26794);
or U29521 (N_29521,N_26370,N_27190);
nor U29522 (N_29522,N_25255,N_25028);
or U29523 (N_29523,N_25575,N_26827);
xnor U29524 (N_29524,N_25252,N_25352);
or U29525 (N_29525,N_27289,N_26148);
or U29526 (N_29526,N_25464,N_27325);
nor U29527 (N_29527,N_25743,N_27223);
or U29528 (N_29528,N_26043,N_25684);
and U29529 (N_29529,N_25398,N_26753);
or U29530 (N_29530,N_25461,N_25978);
xor U29531 (N_29531,N_25314,N_25936);
nand U29532 (N_29532,N_26989,N_25663);
nand U29533 (N_29533,N_25450,N_26083);
xor U29534 (N_29534,N_25248,N_27383);
or U29535 (N_29535,N_25537,N_26161);
nor U29536 (N_29536,N_27258,N_27207);
and U29537 (N_29537,N_27289,N_26747);
and U29538 (N_29538,N_26101,N_27182);
and U29539 (N_29539,N_26600,N_25142);
or U29540 (N_29540,N_25339,N_25973);
nand U29541 (N_29541,N_26603,N_26452);
and U29542 (N_29542,N_26293,N_27283);
xor U29543 (N_29543,N_26520,N_26379);
or U29544 (N_29544,N_25697,N_25427);
nand U29545 (N_29545,N_25450,N_27458);
or U29546 (N_29546,N_25160,N_25970);
xnor U29547 (N_29547,N_27221,N_25004);
or U29548 (N_29548,N_25833,N_25022);
nor U29549 (N_29549,N_25311,N_26675);
xor U29550 (N_29550,N_25988,N_27334);
xnor U29551 (N_29551,N_27124,N_26451);
nor U29552 (N_29552,N_25847,N_26185);
or U29553 (N_29553,N_26566,N_26207);
xnor U29554 (N_29554,N_25418,N_27209);
nor U29555 (N_29555,N_25097,N_25934);
nor U29556 (N_29556,N_26081,N_25298);
xnor U29557 (N_29557,N_25165,N_25236);
nand U29558 (N_29558,N_26970,N_26774);
nand U29559 (N_29559,N_27243,N_25514);
xnor U29560 (N_29560,N_25493,N_25742);
and U29561 (N_29561,N_25875,N_25931);
nor U29562 (N_29562,N_27242,N_26938);
or U29563 (N_29563,N_26488,N_27223);
or U29564 (N_29564,N_25078,N_25403);
xor U29565 (N_29565,N_27010,N_26228);
or U29566 (N_29566,N_27465,N_25426);
nor U29567 (N_29567,N_26894,N_27124);
xnor U29568 (N_29568,N_27119,N_25983);
nor U29569 (N_29569,N_25486,N_26061);
xor U29570 (N_29570,N_25142,N_26051);
nand U29571 (N_29571,N_25615,N_27262);
or U29572 (N_29572,N_27495,N_25682);
nor U29573 (N_29573,N_27269,N_27196);
nand U29574 (N_29574,N_27046,N_26138);
nor U29575 (N_29575,N_25563,N_26442);
and U29576 (N_29576,N_27340,N_27328);
nor U29577 (N_29577,N_26829,N_26396);
or U29578 (N_29578,N_25411,N_26818);
or U29579 (N_29579,N_27316,N_27242);
or U29580 (N_29580,N_26647,N_26009);
or U29581 (N_29581,N_25888,N_26334);
xnor U29582 (N_29582,N_26230,N_26597);
nand U29583 (N_29583,N_25895,N_26354);
and U29584 (N_29584,N_26149,N_26732);
and U29585 (N_29585,N_25529,N_26640);
nand U29586 (N_29586,N_25712,N_25233);
xnor U29587 (N_29587,N_27176,N_25038);
nor U29588 (N_29588,N_26932,N_25332);
and U29589 (N_29589,N_25540,N_26090);
xor U29590 (N_29590,N_27394,N_25631);
nor U29591 (N_29591,N_25576,N_26034);
xor U29592 (N_29592,N_25223,N_26474);
nand U29593 (N_29593,N_25541,N_26556);
xor U29594 (N_29594,N_26100,N_25755);
nand U29595 (N_29595,N_26374,N_26818);
or U29596 (N_29596,N_26473,N_27388);
or U29597 (N_29597,N_26127,N_25974);
nand U29598 (N_29598,N_25890,N_26854);
or U29599 (N_29599,N_25107,N_25620);
or U29600 (N_29600,N_26643,N_26424);
nand U29601 (N_29601,N_26333,N_26294);
nor U29602 (N_29602,N_26702,N_26669);
xnor U29603 (N_29603,N_27356,N_26370);
nor U29604 (N_29604,N_25456,N_26119);
and U29605 (N_29605,N_25295,N_27367);
or U29606 (N_29606,N_25940,N_26166);
xor U29607 (N_29607,N_26505,N_26915);
and U29608 (N_29608,N_27289,N_26107);
nand U29609 (N_29609,N_25719,N_26063);
xnor U29610 (N_29610,N_26605,N_27129);
or U29611 (N_29611,N_26015,N_26901);
nor U29612 (N_29612,N_25313,N_26374);
xnor U29613 (N_29613,N_25692,N_25904);
xnor U29614 (N_29614,N_25560,N_26354);
or U29615 (N_29615,N_25409,N_25560);
and U29616 (N_29616,N_26503,N_27330);
and U29617 (N_29617,N_25549,N_25008);
nand U29618 (N_29618,N_26133,N_26093);
or U29619 (N_29619,N_25797,N_26158);
xnor U29620 (N_29620,N_26635,N_25578);
nor U29621 (N_29621,N_26252,N_26150);
xnor U29622 (N_29622,N_26052,N_25613);
and U29623 (N_29623,N_25302,N_26840);
and U29624 (N_29624,N_25030,N_27082);
xor U29625 (N_29625,N_27043,N_26033);
xor U29626 (N_29626,N_25992,N_25045);
and U29627 (N_29627,N_27352,N_26784);
xnor U29628 (N_29628,N_25760,N_27316);
nor U29629 (N_29629,N_25158,N_25587);
xor U29630 (N_29630,N_26318,N_26493);
xnor U29631 (N_29631,N_25960,N_25588);
nand U29632 (N_29632,N_26903,N_26384);
and U29633 (N_29633,N_26069,N_25120);
or U29634 (N_29634,N_26245,N_26037);
or U29635 (N_29635,N_25264,N_26835);
and U29636 (N_29636,N_25909,N_25699);
xor U29637 (N_29637,N_27410,N_26901);
nor U29638 (N_29638,N_26670,N_27423);
nand U29639 (N_29639,N_26310,N_25678);
xor U29640 (N_29640,N_26321,N_25660);
or U29641 (N_29641,N_27344,N_25474);
xnor U29642 (N_29642,N_25630,N_26815);
and U29643 (N_29643,N_26313,N_26136);
xor U29644 (N_29644,N_25387,N_25642);
nor U29645 (N_29645,N_25049,N_26192);
xnor U29646 (N_29646,N_26110,N_25003);
nor U29647 (N_29647,N_25093,N_27466);
nand U29648 (N_29648,N_25157,N_26970);
nor U29649 (N_29649,N_26193,N_26331);
nand U29650 (N_29650,N_25951,N_25588);
nand U29651 (N_29651,N_25437,N_27002);
nand U29652 (N_29652,N_25366,N_26466);
xnor U29653 (N_29653,N_25346,N_27070);
or U29654 (N_29654,N_25284,N_25348);
nor U29655 (N_29655,N_25874,N_26356);
nand U29656 (N_29656,N_25862,N_27303);
nand U29657 (N_29657,N_26742,N_26898);
and U29658 (N_29658,N_26225,N_25412);
nand U29659 (N_29659,N_27481,N_26739);
and U29660 (N_29660,N_25793,N_25910);
nor U29661 (N_29661,N_27108,N_25675);
nand U29662 (N_29662,N_27213,N_25942);
nand U29663 (N_29663,N_25878,N_25163);
or U29664 (N_29664,N_26456,N_25642);
and U29665 (N_29665,N_26811,N_26788);
nor U29666 (N_29666,N_26848,N_26948);
and U29667 (N_29667,N_26115,N_26916);
xnor U29668 (N_29668,N_26054,N_26822);
or U29669 (N_29669,N_27496,N_26771);
nor U29670 (N_29670,N_26278,N_26531);
nor U29671 (N_29671,N_27234,N_26874);
nand U29672 (N_29672,N_26466,N_26497);
nand U29673 (N_29673,N_26193,N_27128);
nand U29674 (N_29674,N_26306,N_27329);
or U29675 (N_29675,N_27495,N_25525);
xnor U29676 (N_29676,N_25190,N_27044);
xnor U29677 (N_29677,N_25616,N_25301);
and U29678 (N_29678,N_27491,N_25842);
nand U29679 (N_29679,N_26415,N_26037);
nor U29680 (N_29680,N_26002,N_25503);
nor U29681 (N_29681,N_25766,N_26605);
or U29682 (N_29682,N_26523,N_25591);
and U29683 (N_29683,N_25720,N_26152);
nor U29684 (N_29684,N_25740,N_27422);
and U29685 (N_29685,N_25813,N_26940);
xor U29686 (N_29686,N_27310,N_27422);
xnor U29687 (N_29687,N_25522,N_26499);
xor U29688 (N_29688,N_26574,N_25864);
xor U29689 (N_29689,N_26713,N_27168);
or U29690 (N_29690,N_26981,N_26208);
or U29691 (N_29691,N_25282,N_26466);
xnor U29692 (N_29692,N_25543,N_27159);
or U29693 (N_29693,N_25634,N_25968);
xnor U29694 (N_29694,N_25019,N_26699);
and U29695 (N_29695,N_25726,N_25169);
and U29696 (N_29696,N_26065,N_27499);
xnor U29697 (N_29697,N_26017,N_25430);
nand U29698 (N_29698,N_26614,N_25776);
nand U29699 (N_29699,N_25135,N_25483);
and U29700 (N_29700,N_26481,N_25700);
and U29701 (N_29701,N_26865,N_25330);
or U29702 (N_29702,N_25985,N_26518);
and U29703 (N_29703,N_26840,N_26823);
nor U29704 (N_29704,N_25564,N_25943);
and U29705 (N_29705,N_27341,N_26626);
nor U29706 (N_29706,N_26540,N_26996);
or U29707 (N_29707,N_26287,N_27051);
or U29708 (N_29708,N_26862,N_26167);
or U29709 (N_29709,N_25274,N_26782);
nor U29710 (N_29710,N_26427,N_26267);
nand U29711 (N_29711,N_26575,N_25637);
and U29712 (N_29712,N_27398,N_27150);
nor U29713 (N_29713,N_25879,N_25009);
or U29714 (N_29714,N_25261,N_27011);
nand U29715 (N_29715,N_25604,N_27327);
nor U29716 (N_29716,N_26985,N_26316);
and U29717 (N_29717,N_26790,N_25293);
xnor U29718 (N_29718,N_26289,N_26852);
or U29719 (N_29719,N_26352,N_26132);
or U29720 (N_29720,N_26007,N_25240);
and U29721 (N_29721,N_26152,N_26092);
xor U29722 (N_29722,N_27169,N_25498);
and U29723 (N_29723,N_26866,N_25059);
or U29724 (N_29724,N_25467,N_25056);
nor U29725 (N_29725,N_25056,N_27328);
xnor U29726 (N_29726,N_25212,N_26934);
nor U29727 (N_29727,N_26522,N_26002);
nor U29728 (N_29728,N_25350,N_26308);
nor U29729 (N_29729,N_26665,N_27205);
xor U29730 (N_29730,N_26375,N_27270);
xnor U29731 (N_29731,N_27207,N_25693);
nor U29732 (N_29732,N_27000,N_27216);
or U29733 (N_29733,N_25699,N_27341);
nand U29734 (N_29734,N_27449,N_26206);
xor U29735 (N_29735,N_27377,N_26064);
or U29736 (N_29736,N_27132,N_26368);
nand U29737 (N_29737,N_26076,N_26389);
xnor U29738 (N_29738,N_25661,N_26742);
nor U29739 (N_29739,N_25498,N_25642);
xor U29740 (N_29740,N_25181,N_25714);
and U29741 (N_29741,N_27075,N_25464);
nand U29742 (N_29742,N_27340,N_26369);
and U29743 (N_29743,N_25054,N_25988);
nor U29744 (N_29744,N_27342,N_26446);
nand U29745 (N_29745,N_27198,N_27428);
or U29746 (N_29746,N_27350,N_26167);
and U29747 (N_29747,N_25001,N_27246);
or U29748 (N_29748,N_25353,N_25728);
xor U29749 (N_29749,N_25979,N_25142);
xnor U29750 (N_29750,N_25424,N_27129);
and U29751 (N_29751,N_26382,N_26141);
xor U29752 (N_29752,N_25360,N_25834);
nand U29753 (N_29753,N_25503,N_27229);
and U29754 (N_29754,N_25281,N_25907);
and U29755 (N_29755,N_27258,N_25649);
or U29756 (N_29756,N_25709,N_25828);
nand U29757 (N_29757,N_25878,N_26125);
xnor U29758 (N_29758,N_25194,N_27461);
and U29759 (N_29759,N_26511,N_26090);
nor U29760 (N_29760,N_25693,N_26670);
or U29761 (N_29761,N_26187,N_25580);
and U29762 (N_29762,N_26105,N_26701);
or U29763 (N_29763,N_26582,N_27234);
nor U29764 (N_29764,N_26419,N_27464);
nor U29765 (N_29765,N_26122,N_25229);
nor U29766 (N_29766,N_25710,N_25733);
xor U29767 (N_29767,N_27038,N_25278);
or U29768 (N_29768,N_25581,N_26433);
nor U29769 (N_29769,N_25250,N_26388);
xnor U29770 (N_29770,N_25239,N_26532);
nand U29771 (N_29771,N_25231,N_25869);
or U29772 (N_29772,N_27024,N_26599);
xor U29773 (N_29773,N_26234,N_26720);
and U29774 (N_29774,N_25633,N_25406);
nor U29775 (N_29775,N_27114,N_25209);
nor U29776 (N_29776,N_25008,N_26318);
xnor U29777 (N_29777,N_25885,N_27354);
and U29778 (N_29778,N_25053,N_25188);
and U29779 (N_29779,N_26942,N_27225);
nand U29780 (N_29780,N_25498,N_27377);
nand U29781 (N_29781,N_25552,N_25498);
nand U29782 (N_29782,N_27408,N_25210);
nand U29783 (N_29783,N_25428,N_26418);
xnor U29784 (N_29784,N_26325,N_26513);
xor U29785 (N_29785,N_26326,N_26832);
xnor U29786 (N_29786,N_26629,N_26568);
and U29787 (N_29787,N_27361,N_27328);
nor U29788 (N_29788,N_26310,N_25409);
nor U29789 (N_29789,N_26247,N_25103);
nand U29790 (N_29790,N_26202,N_26790);
or U29791 (N_29791,N_25943,N_25738);
and U29792 (N_29792,N_25305,N_26523);
nor U29793 (N_29793,N_26914,N_26754);
and U29794 (N_29794,N_25266,N_25743);
xnor U29795 (N_29795,N_25626,N_27461);
and U29796 (N_29796,N_26047,N_26171);
nand U29797 (N_29797,N_25615,N_25359);
or U29798 (N_29798,N_25230,N_26958);
or U29799 (N_29799,N_25925,N_25937);
xor U29800 (N_29800,N_25524,N_26755);
or U29801 (N_29801,N_26017,N_27294);
nor U29802 (N_29802,N_27187,N_25437);
nand U29803 (N_29803,N_26446,N_25381);
nor U29804 (N_29804,N_26093,N_26470);
or U29805 (N_29805,N_25071,N_25782);
nand U29806 (N_29806,N_26940,N_26214);
nand U29807 (N_29807,N_26727,N_26850);
or U29808 (N_29808,N_25618,N_26803);
nand U29809 (N_29809,N_26068,N_25707);
xnor U29810 (N_29810,N_27320,N_27223);
nand U29811 (N_29811,N_26423,N_26022);
nor U29812 (N_29812,N_26592,N_25391);
xnor U29813 (N_29813,N_25526,N_25269);
xnor U29814 (N_29814,N_25294,N_27096);
nand U29815 (N_29815,N_27307,N_27086);
nor U29816 (N_29816,N_25308,N_25800);
nor U29817 (N_29817,N_25205,N_25573);
xor U29818 (N_29818,N_27399,N_25450);
xor U29819 (N_29819,N_26310,N_27326);
nor U29820 (N_29820,N_26042,N_27016);
and U29821 (N_29821,N_26736,N_25156);
nor U29822 (N_29822,N_26359,N_26431);
nor U29823 (N_29823,N_25749,N_25392);
xnor U29824 (N_29824,N_25037,N_26072);
xnor U29825 (N_29825,N_26493,N_26342);
or U29826 (N_29826,N_25390,N_25262);
xnor U29827 (N_29827,N_25635,N_26428);
and U29828 (N_29828,N_25775,N_26037);
and U29829 (N_29829,N_27289,N_26902);
or U29830 (N_29830,N_26117,N_25220);
nor U29831 (N_29831,N_26150,N_26931);
nor U29832 (N_29832,N_25321,N_25762);
nand U29833 (N_29833,N_25948,N_26925);
xnor U29834 (N_29834,N_25572,N_25199);
or U29835 (N_29835,N_26802,N_27021);
nand U29836 (N_29836,N_25639,N_27059);
nor U29837 (N_29837,N_27454,N_26194);
or U29838 (N_29838,N_26016,N_25375);
nand U29839 (N_29839,N_26566,N_25483);
nor U29840 (N_29840,N_26273,N_25053);
nand U29841 (N_29841,N_25679,N_26793);
and U29842 (N_29842,N_27281,N_26620);
nor U29843 (N_29843,N_25253,N_25727);
xor U29844 (N_29844,N_25917,N_25565);
xnor U29845 (N_29845,N_25355,N_25795);
nor U29846 (N_29846,N_27110,N_25612);
and U29847 (N_29847,N_26296,N_26496);
and U29848 (N_29848,N_26785,N_25568);
and U29849 (N_29849,N_27186,N_26738);
nand U29850 (N_29850,N_26834,N_27497);
xor U29851 (N_29851,N_25522,N_27051);
and U29852 (N_29852,N_26728,N_27292);
xnor U29853 (N_29853,N_26396,N_25139);
nand U29854 (N_29854,N_26513,N_27193);
and U29855 (N_29855,N_25761,N_25519);
and U29856 (N_29856,N_26985,N_25323);
or U29857 (N_29857,N_25408,N_25172);
nor U29858 (N_29858,N_27354,N_27399);
nor U29859 (N_29859,N_27435,N_27431);
and U29860 (N_29860,N_25587,N_26594);
xor U29861 (N_29861,N_25836,N_26868);
or U29862 (N_29862,N_26912,N_25776);
xor U29863 (N_29863,N_26075,N_25276);
and U29864 (N_29864,N_26108,N_27383);
nor U29865 (N_29865,N_26767,N_26726);
nor U29866 (N_29866,N_26760,N_25446);
nor U29867 (N_29867,N_26385,N_25658);
and U29868 (N_29868,N_26624,N_25418);
nand U29869 (N_29869,N_25788,N_27301);
or U29870 (N_29870,N_25449,N_26593);
and U29871 (N_29871,N_26774,N_26159);
and U29872 (N_29872,N_27132,N_25830);
xor U29873 (N_29873,N_26725,N_26371);
nor U29874 (N_29874,N_25697,N_25966);
or U29875 (N_29875,N_26063,N_25629);
xor U29876 (N_29876,N_25507,N_26685);
and U29877 (N_29877,N_26801,N_26922);
nor U29878 (N_29878,N_27104,N_25475);
nand U29879 (N_29879,N_26560,N_26930);
and U29880 (N_29880,N_25119,N_26939);
or U29881 (N_29881,N_26846,N_27126);
xor U29882 (N_29882,N_27474,N_25469);
nand U29883 (N_29883,N_26815,N_26723);
nand U29884 (N_29884,N_25227,N_25651);
or U29885 (N_29885,N_26749,N_27025);
or U29886 (N_29886,N_27096,N_25485);
nand U29887 (N_29887,N_26377,N_26475);
nand U29888 (N_29888,N_27214,N_26818);
xnor U29889 (N_29889,N_26416,N_26785);
and U29890 (N_29890,N_25888,N_26851);
and U29891 (N_29891,N_27451,N_26820);
xnor U29892 (N_29892,N_25619,N_27247);
xor U29893 (N_29893,N_26004,N_26256);
and U29894 (N_29894,N_27345,N_25102);
or U29895 (N_29895,N_26102,N_25727);
nor U29896 (N_29896,N_27076,N_26270);
nand U29897 (N_29897,N_27154,N_27306);
nor U29898 (N_29898,N_25069,N_25612);
nand U29899 (N_29899,N_26977,N_25696);
or U29900 (N_29900,N_25164,N_25768);
and U29901 (N_29901,N_26397,N_26408);
nand U29902 (N_29902,N_26791,N_25462);
or U29903 (N_29903,N_26789,N_25930);
and U29904 (N_29904,N_26010,N_26224);
nor U29905 (N_29905,N_25822,N_25686);
nand U29906 (N_29906,N_26415,N_27032);
or U29907 (N_29907,N_25746,N_25385);
xor U29908 (N_29908,N_25531,N_25542);
nand U29909 (N_29909,N_26640,N_26737);
nand U29910 (N_29910,N_27384,N_25129);
nand U29911 (N_29911,N_27462,N_26789);
xnor U29912 (N_29912,N_26033,N_25489);
nor U29913 (N_29913,N_26277,N_25301);
nor U29914 (N_29914,N_25988,N_26626);
nor U29915 (N_29915,N_26055,N_26713);
nor U29916 (N_29916,N_26157,N_25885);
and U29917 (N_29917,N_25468,N_26905);
and U29918 (N_29918,N_25072,N_25891);
nor U29919 (N_29919,N_26122,N_27122);
nor U29920 (N_29920,N_26830,N_25236);
nand U29921 (N_29921,N_26522,N_26077);
nand U29922 (N_29922,N_26353,N_26062);
or U29923 (N_29923,N_25077,N_25175);
and U29924 (N_29924,N_27012,N_26072);
nor U29925 (N_29925,N_27311,N_25720);
or U29926 (N_29926,N_26247,N_25993);
xnor U29927 (N_29927,N_26644,N_26232);
or U29928 (N_29928,N_27351,N_26022);
or U29929 (N_29929,N_26585,N_27386);
xor U29930 (N_29930,N_25409,N_25798);
xor U29931 (N_29931,N_26613,N_25621);
nand U29932 (N_29932,N_25983,N_26033);
nand U29933 (N_29933,N_25587,N_26901);
and U29934 (N_29934,N_25082,N_26505);
nor U29935 (N_29935,N_26525,N_25514);
and U29936 (N_29936,N_26180,N_25320);
and U29937 (N_29937,N_26195,N_26469);
and U29938 (N_29938,N_26148,N_26736);
nor U29939 (N_29939,N_27402,N_26343);
and U29940 (N_29940,N_26982,N_27051);
xor U29941 (N_29941,N_27088,N_26766);
or U29942 (N_29942,N_26157,N_26970);
or U29943 (N_29943,N_26950,N_25477);
or U29944 (N_29944,N_25719,N_25914);
or U29945 (N_29945,N_26597,N_25938);
nor U29946 (N_29946,N_27236,N_27335);
xor U29947 (N_29947,N_26924,N_25256);
xor U29948 (N_29948,N_26048,N_26562);
or U29949 (N_29949,N_26027,N_26379);
and U29950 (N_29950,N_25455,N_25908);
xor U29951 (N_29951,N_26843,N_27395);
and U29952 (N_29952,N_25718,N_25746);
nor U29953 (N_29953,N_26804,N_26226);
nor U29954 (N_29954,N_26390,N_26685);
or U29955 (N_29955,N_25281,N_25392);
nand U29956 (N_29956,N_27003,N_27223);
nor U29957 (N_29957,N_25623,N_26128);
and U29958 (N_29958,N_27034,N_25869);
xor U29959 (N_29959,N_25082,N_25035);
and U29960 (N_29960,N_25645,N_26215);
nand U29961 (N_29961,N_26327,N_25654);
xor U29962 (N_29962,N_26861,N_26121);
xnor U29963 (N_29963,N_26179,N_26251);
nand U29964 (N_29964,N_25180,N_25518);
and U29965 (N_29965,N_25012,N_25780);
or U29966 (N_29966,N_26196,N_27366);
and U29967 (N_29967,N_26163,N_25027);
or U29968 (N_29968,N_25254,N_26526);
nand U29969 (N_29969,N_26501,N_27388);
or U29970 (N_29970,N_25627,N_25155);
nor U29971 (N_29971,N_26311,N_26389);
nand U29972 (N_29972,N_26057,N_25468);
and U29973 (N_29973,N_27189,N_25461);
xnor U29974 (N_29974,N_26569,N_27152);
xnor U29975 (N_29975,N_26749,N_25574);
nand U29976 (N_29976,N_25750,N_25593);
nand U29977 (N_29977,N_25070,N_26565);
and U29978 (N_29978,N_26190,N_26611);
and U29979 (N_29979,N_25295,N_26898);
and U29980 (N_29980,N_26217,N_26508);
xnor U29981 (N_29981,N_25867,N_27093);
and U29982 (N_29982,N_27404,N_26720);
or U29983 (N_29983,N_26891,N_25316);
nand U29984 (N_29984,N_26439,N_26120);
nor U29985 (N_29985,N_25223,N_27407);
xor U29986 (N_29986,N_27072,N_25178);
or U29987 (N_29987,N_25812,N_26670);
nor U29988 (N_29988,N_26916,N_26942);
nor U29989 (N_29989,N_26727,N_25825);
nor U29990 (N_29990,N_26396,N_25804);
and U29991 (N_29991,N_25155,N_26348);
and U29992 (N_29992,N_25623,N_27123);
nor U29993 (N_29993,N_25491,N_25606);
and U29994 (N_29994,N_27203,N_27080);
xnor U29995 (N_29995,N_25972,N_26887);
xnor U29996 (N_29996,N_25369,N_27249);
nand U29997 (N_29997,N_26071,N_26914);
nor U29998 (N_29998,N_25520,N_26171);
or U29999 (N_29999,N_25292,N_25535);
xnor U30000 (N_30000,N_27641,N_27543);
nor U30001 (N_30001,N_29929,N_27876);
or U30002 (N_30002,N_28249,N_29757);
xnor U30003 (N_30003,N_27820,N_29676);
nor U30004 (N_30004,N_28765,N_28733);
nor U30005 (N_30005,N_28118,N_29762);
nor U30006 (N_30006,N_28583,N_29182);
xnor U30007 (N_30007,N_27802,N_28231);
xor U30008 (N_30008,N_27628,N_29086);
or U30009 (N_30009,N_28885,N_28225);
nand U30010 (N_30010,N_27880,N_29355);
and U30011 (N_30011,N_29284,N_28565);
or U30012 (N_30012,N_28900,N_27702);
nand U30013 (N_30013,N_29026,N_29982);
nand U30014 (N_30014,N_29326,N_28581);
and U30015 (N_30015,N_29393,N_29138);
xor U30016 (N_30016,N_29611,N_29339);
and U30017 (N_30017,N_29560,N_29065);
nor U30018 (N_30018,N_29937,N_29570);
nand U30019 (N_30019,N_29195,N_29750);
nor U30020 (N_30020,N_29583,N_28999);
xnor U30021 (N_30021,N_29928,N_27668);
xor U30022 (N_30022,N_29966,N_28797);
and U30023 (N_30023,N_29502,N_27715);
xnor U30024 (N_30024,N_28020,N_29740);
xnor U30025 (N_30025,N_28587,N_28075);
nor U30026 (N_30026,N_28402,N_28428);
xnor U30027 (N_30027,N_28189,N_29069);
nor U30028 (N_30028,N_28171,N_28140);
nand U30029 (N_30029,N_27741,N_27546);
and U30030 (N_30030,N_28853,N_29429);
xor U30031 (N_30031,N_28701,N_29745);
or U30032 (N_30032,N_28337,N_28837);
or U30033 (N_30033,N_27530,N_29246);
nor U30034 (N_30034,N_27701,N_28568);
or U30035 (N_30035,N_29374,N_28083);
and U30036 (N_30036,N_27653,N_27629);
xnor U30037 (N_30037,N_28324,N_29903);
and U30038 (N_30038,N_29948,N_29634);
xor U30039 (N_30039,N_28247,N_28041);
and U30040 (N_30040,N_27966,N_28584);
xnor U30041 (N_30041,N_29964,N_28120);
or U30042 (N_30042,N_29522,N_27679);
nand U30043 (N_30043,N_29555,N_27719);
nand U30044 (N_30044,N_28112,N_28699);
nand U30045 (N_30045,N_29513,N_29818);
nor U30046 (N_30046,N_28170,N_27821);
xor U30047 (N_30047,N_29987,N_29702);
nor U30048 (N_30048,N_29409,N_28614);
nor U30049 (N_30049,N_29465,N_28436);
and U30050 (N_30050,N_28062,N_28310);
and U30051 (N_30051,N_29358,N_28743);
nand U30052 (N_30052,N_28259,N_28946);
xnor U30053 (N_30053,N_27758,N_28117);
nor U30054 (N_30054,N_28246,N_28983);
nand U30055 (N_30055,N_27924,N_29161);
xnor U30056 (N_30056,N_29667,N_29243);
nand U30057 (N_30057,N_28443,N_29410);
nand U30058 (N_30058,N_28716,N_29835);
xnor U30059 (N_30059,N_29067,N_29994);
nor U30060 (N_30060,N_28215,N_28113);
xor U30061 (N_30061,N_27774,N_28490);
and U30062 (N_30062,N_28632,N_29211);
nand U30063 (N_30063,N_28509,N_29654);
and U30064 (N_30064,N_28579,N_27982);
or U30065 (N_30065,N_29594,N_28292);
xor U30066 (N_30066,N_28839,N_28732);
and U30067 (N_30067,N_28939,N_28407);
or U30068 (N_30068,N_28116,N_29830);
nand U30069 (N_30069,N_29181,N_28236);
or U30070 (N_30070,N_28227,N_28448);
nor U30071 (N_30071,N_28143,N_27515);
nor U30072 (N_30072,N_28412,N_28220);
nand U30073 (N_30073,N_28858,N_29581);
nand U30074 (N_30074,N_29106,N_27650);
or U30075 (N_30075,N_28274,N_28195);
and U30076 (N_30076,N_29552,N_28491);
and U30077 (N_30077,N_28234,N_28954);
nand U30078 (N_30078,N_28929,N_29005);
or U30079 (N_30079,N_29970,N_29126);
nand U30080 (N_30080,N_27816,N_29864);
and U30081 (N_30081,N_29021,N_29691);
or U30082 (N_30082,N_28869,N_28350);
or U30083 (N_30083,N_28627,N_28023);
nand U30084 (N_30084,N_29045,N_28639);
nand U30085 (N_30085,N_29041,N_28437);
nor U30086 (N_30086,N_29427,N_29879);
nand U30087 (N_30087,N_29669,N_29638);
xor U30088 (N_30088,N_29647,N_28389);
nand U30089 (N_30089,N_28940,N_28164);
nand U30090 (N_30090,N_29871,N_29598);
xnor U30091 (N_30091,N_27926,N_28744);
or U30092 (N_30092,N_27936,N_28703);
xor U30093 (N_30093,N_28003,N_27992);
nor U30094 (N_30094,N_29798,N_29807);
nand U30095 (N_30095,N_29518,N_29420);
nor U30096 (N_30096,N_29257,N_28862);
nand U30097 (N_30097,N_28567,N_27755);
nor U30098 (N_30098,N_28530,N_28365);
and U30099 (N_30099,N_29276,N_29331);
nand U30100 (N_30100,N_28128,N_27670);
nand U30101 (N_30101,N_28185,N_28950);
and U30102 (N_30102,N_27549,N_28492);
or U30103 (N_30103,N_28630,N_28846);
nor U30104 (N_30104,N_29505,N_28408);
nor U30105 (N_30105,N_29817,N_29956);
nor U30106 (N_30106,N_29279,N_29372);
or U30107 (N_30107,N_29946,N_28756);
or U30108 (N_30108,N_28049,N_28764);
or U30109 (N_30109,N_29703,N_28966);
xnor U30110 (N_30110,N_27999,N_29576);
or U30111 (N_30111,N_27511,N_29862);
or U30112 (N_30112,N_27827,N_29605);
nand U30113 (N_30113,N_27858,N_28758);
and U30114 (N_30114,N_28620,N_28551);
nand U30115 (N_30115,N_28386,N_28729);
nor U30116 (N_30116,N_29778,N_29042);
xnor U30117 (N_30117,N_27792,N_29655);
xnor U30118 (N_30118,N_27911,N_28461);
xor U30119 (N_30119,N_27797,N_28129);
nand U30120 (N_30120,N_28349,N_28072);
xor U30121 (N_30121,N_29878,N_28156);
or U30122 (N_30122,N_27839,N_28155);
or U30123 (N_30123,N_29474,N_29436);
nor U30124 (N_30124,N_29311,N_28086);
and U30125 (N_30125,N_29530,N_28816);
nand U30126 (N_30126,N_29547,N_29422);
nor U30127 (N_30127,N_29678,N_28714);
nor U30128 (N_30128,N_29336,N_28652);
nor U30129 (N_30129,N_29932,N_28243);
xor U30130 (N_30130,N_28099,N_28887);
or U30131 (N_30131,N_29764,N_28256);
nand U30132 (N_30132,N_29240,N_28146);
nor U30133 (N_30133,N_28500,N_28042);
xnor U30134 (N_30134,N_27994,N_29219);
nor U30135 (N_30135,N_28269,N_29218);
nor U30136 (N_30136,N_28242,N_27788);
and U30137 (N_30137,N_29991,N_29664);
nand U30138 (N_30138,N_27939,N_28859);
xnor U30139 (N_30139,N_29743,N_27824);
nand U30140 (N_30140,N_27739,N_28449);
and U30141 (N_30141,N_28844,N_27913);
and U30142 (N_30142,N_28495,N_29484);
xnor U30143 (N_30143,N_28683,N_28138);
nor U30144 (N_30144,N_29854,N_27748);
xor U30145 (N_30145,N_27882,N_29093);
and U30146 (N_30146,N_28606,N_28822);
xnor U30147 (N_30147,N_27932,N_29824);
xor U30148 (N_30148,N_29385,N_29738);
xor U30149 (N_30149,N_27749,N_28961);
and U30150 (N_30150,N_28089,N_27840);
or U30151 (N_30151,N_28895,N_28253);
nor U30152 (N_30152,N_28665,N_29147);
or U30153 (N_30153,N_29012,N_28297);
nand U30154 (N_30154,N_28860,N_29969);
nand U30155 (N_30155,N_29345,N_28254);
nor U30156 (N_30156,N_29488,N_29592);
and U30157 (N_30157,N_28807,N_27675);
nand U30158 (N_30158,N_28369,N_27895);
and U30159 (N_30159,N_28209,N_29054);
xnor U30160 (N_30160,N_29601,N_29875);
and U30161 (N_30161,N_28188,N_29618);
nand U30162 (N_30162,N_29085,N_28158);
nor U30163 (N_30163,N_28087,N_28941);
and U30164 (N_30164,N_28442,N_29228);
and U30165 (N_30165,N_29914,N_29828);
xor U30166 (N_30166,N_27615,N_27518);
nand U30167 (N_30167,N_29399,N_28842);
nand U30168 (N_30168,N_29172,N_29370);
and U30169 (N_30169,N_28051,N_29863);
or U30170 (N_30170,N_29538,N_29074);
or U30171 (N_30171,N_29723,N_29827);
nor U30172 (N_30172,N_29023,N_29585);
nor U30173 (N_30173,N_29857,N_28498);
nand U30174 (N_30174,N_28291,N_29789);
and U30175 (N_30175,N_27981,N_29758);
or U30176 (N_30176,N_28791,N_28897);
nor U30177 (N_30177,N_28507,N_27985);
nand U30178 (N_30178,N_29213,N_27754);
or U30179 (N_30179,N_29842,N_28589);
xnor U30180 (N_30180,N_28539,N_27892);
xor U30181 (N_30181,N_27815,N_28841);
or U30182 (N_30182,N_29548,N_29471);
nor U30183 (N_30183,N_29114,N_27909);
and U30184 (N_30184,N_27517,N_28675);
and U30185 (N_30185,N_27953,N_29721);
xnor U30186 (N_30186,N_28226,N_28692);
and U30187 (N_30187,N_28060,N_29531);
nand U30188 (N_30188,N_27676,N_28239);
and U30189 (N_30189,N_27712,N_29203);
and U30190 (N_30190,N_28727,N_29155);
nand U30191 (N_30191,N_29623,N_28988);
nor U30192 (N_30192,N_29404,N_28906);
or U30193 (N_30193,N_29603,N_28237);
nor U30194 (N_30194,N_28278,N_28682);
or U30195 (N_30195,N_28981,N_28302);
or U30196 (N_30196,N_29917,N_29645);
nand U30197 (N_30197,N_28817,N_27962);
nor U30198 (N_30198,N_27584,N_28531);
nand U30199 (N_30199,N_29796,N_29148);
nor U30200 (N_30200,N_27760,N_28308);
or U30201 (N_30201,N_29786,N_29774);
xor U30202 (N_30202,N_29048,N_27655);
xor U30203 (N_30203,N_29032,N_28355);
or U30204 (N_30204,N_27567,N_28248);
and U30205 (N_30205,N_28423,N_28706);
nand U30206 (N_30206,N_27979,N_27886);
or U30207 (N_30207,N_29325,N_29597);
nor U30208 (N_30208,N_29280,N_28715);
nor U30209 (N_30209,N_29259,N_29584);
nor U30210 (N_30210,N_29532,N_29935);
nor U30211 (N_30211,N_27734,N_28640);
or U30212 (N_30212,N_27885,N_27875);
and U30213 (N_30213,N_27989,N_29865);
or U30214 (N_30214,N_29099,N_29558);
nand U30215 (N_30215,N_28329,N_27878);
and U30216 (N_30216,N_28053,N_28997);
xnor U30217 (N_30217,N_29298,N_29950);
and U30218 (N_30218,N_29707,N_29299);
and U30219 (N_30219,N_28690,N_28725);
and U30220 (N_30220,N_28331,N_29156);
and U30221 (N_30221,N_29630,N_29710);
or U30222 (N_30222,N_29641,N_29307);
xnor U30223 (N_30223,N_28938,N_27845);
nand U30224 (N_30224,N_29260,N_27678);
nor U30225 (N_30225,N_28205,N_29814);
xor U30226 (N_30226,N_27529,N_27569);
nand U30227 (N_30227,N_29556,N_27532);
nand U30228 (N_30228,N_29995,N_29251);
nand U30229 (N_30229,N_28984,N_28528);
nor U30230 (N_30230,N_28043,N_29081);
and U30231 (N_30231,N_27935,N_27938);
or U30232 (N_30232,N_28502,N_28212);
xor U30233 (N_30233,N_28504,N_27578);
and U30234 (N_30234,N_29639,N_27697);
nor U30235 (N_30235,N_27680,N_28616);
and U30236 (N_30236,N_28258,N_28126);
xor U30237 (N_30237,N_28081,N_28252);
nor U30238 (N_30238,N_28121,N_28417);
nand U30239 (N_30239,N_29868,N_29826);
nor U30240 (N_30240,N_28338,N_29608);
and U30241 (N_30241,N_27705,N_29491);
and U30242 (N_30242,N_28625,N_28019);
and U30243 (N_30243,N_28775,N_28615);
and U30244 (N_30244,N_29015,N_27575);
nor U30245 (N_30245,N_27786,N_28933);
or U30246 (N_30246,N_27978,N_29196);
nand U30247 (N_30247,N_29766,N_29342);
xor U30248 (N_30248,N_28012,N_29869);
or U30249 (N_30249,N_28857,N_28580);
or U30250 (N_30250,N_29121,N_27681);
nor U30251 (N_30251,N_29697,N_29199);
and U30252 (N_30252,N_28216,N_28367);
or U30253 (N_30253,N_28918,N_29263);
nand U30254 (N_30254,N_29470,N_29289);
xor U30255 (N_30255,N_28371,N_27894);
or U30256 (N_30256,N_28034,N_29706);
xnor U30257 (N_30257,N_29273,N_28325);
or U30258 (N_30258,N_29557,N_28293);
and U30259 (N_30259,N_28629,N_28908);
and U30260 (N_30260,N_28124,N_27706);
nor U30261 (N_30261,N_29449,N_29340);
or U30262 (N_30262,N_28336,N_27506);
nand U30263 (N_30263,N_28809,N_28920);
xnor U30264 (N_30264,N_28578,N_27730);
nor U30265 (N_30265,N_27535,N_29978);
xor U30266 (N_30266,N_29636,N_29812);
nand U30267 (N_30267,N_28183,N_29511);
or U30268 (N_30268,N_28965,N_28169);
nand U30269 (N_30269,N_29642,N_29785);
xnor U30270 (N_30270,N_29759,N_27718);
nand U30271 (N_30271,N_29400,N_29687);
xnor U30272 (N_30272,N_29271,N_29799);
or U30273 (N_30273,N_27544,N_28586);
nor U30274 (N_30274,N_29406,N_29163);
nor U30275 (N_30275,N_27862,N_28280);
or U30276 (N_30276,N_28240,N_28610);
nand U30277 (N_30277,N_28400,N_27829);
nand U30278 (N_30278,N_29795,N_27647);
or U30279 (N_30279,N_27625,N_27975);
nand U30280 (N_30280,N_29787,N_29305);
or U30281 (N_30281,N_29487,N_29709);
and U30282 (N_30282,N_28322,N_28264);
or U30283 (N_30283,N_27804,N_27574);
or U30284 (N_30284,N_28284,N_27656);
nor U30285 (N_30285,N_28218,N_29619);
xor U30286 (N_30286,N_29128,N_27539);
and U30287 (N_30287,N_29770,N_29159);
and U30288 (N_30288,N_29316,N_28262);
nand U30289 (N_30289,N_29900,N_29523);
nand U30290 (N_30290,N_29103,N_28330);
nor U30291 (N_30291,N_28326,N_27841);
nand U30292 (N_30292,N_28393,N_27686);
or U30293 (N_30293,N_28229,N_29413);
xor U30294 (N_30294,N_28320,N_28711);
or U30295 (N_30295,N_29816,N_27607);
and U30296 (N_30296,N_28193,N_29380);
xor U30297 (N_30297,N_29674,N_28410);
and U30298 (N_30298,N_27639,N_29292);
nor U30299 (N_30299,N_27777,N_29977);
nor U30300 (N_30300,N_29483,N_29751);
xor U30301 (N_30301,N_29076,N_29028);
xnor U30302 (N_30302,N_27799,N_29823);
nand U30303 (N_30303,N_28401,N_28295);
nor U30304 (N_30304,N_27587,N_27551);
nor U30305 (N_30305,N_29407,N_27609);
nand U30306 (N_30306,N_29694,N_27907);
xnor U30307 (N_30307,N_28406,N_29108);
xor U30308 (N_30308,N_29784,N_28840);
nor U30309 (N_30309,N_29190,N_29847);
nand U30310 (N_30310,N_27643,N_28752);
and U30311 (N_30311,N_28207,N_29446);
nand U30312 (N_30312,N_29539,N_28646);
nor U30313 (N_30313,N_29025,N_28912);
xor U30314 (N_30314,N_28135,N_29973);
nand U30315 (N_30315,N_29221,N_28079);
nand U30316 (N_30316,N_29442,N_28647);
nand U30317 (N_30317,N_29120,N_27996);
xnor U30318 (N_30318,N_28190,N_28778);
and U30319 (N_30319,N_28546,N_27770);
or U30320 (N_30320,N_29614,N_27874);
and U30321 (N_30321,N_27708,N_27500);
nand U30322 (N_30322,N_27794,N_28137);
and U30323 (N_30323,N_28708,N_29281);
xor U30324 (N_30324,N_29888,N_29653);
or U30325 (N_30325,N_29070,N_29658);
nor U30326 (N_30326,N_27509,N_27649);
or U30327 (N_30327,N_27921,N_29278);
and U30328 (N_30328,N_27901,N_28497);
or U30329 (N_30329,N_29509,N_28222);
or U30330 (N_30330,N_28718,N_28092);
nand U30331 (N_30331,N_29017,N_28516);
nand U30332 (N_30332,N_27793,N_27555);
nor U30333 (N_30333,N_29902,N_28694);
or U30334 (N_30334,N_28179,N_28317);
nor U30335 (N_30335,N_29606,N_29495);
nand U30336 (N_30336,N_29177,N_29665);
nor U30337 (N_30337,N_28010,N_29733);
and U30338 (N_30338,N_29423,N_28709);
or U30339 (N_30339,N_28696,N_27965);
xor U30340 (N_30340,N_28390,N_27943);
xor U30341 (N_30341,N_27957,N_28747);
nand U30342 (N_30342,N_29717,N_27764);
or U30343 (N_30343,N_28000,N_29082);
and U30344 (N_30344,N_29980,N_29383);
xor U30345 (N_30345,N_27685,N_29401);
and U30346 (N_30346,N_29515,N_28953);
xnor U30347 (N_30347,N_27906,N_28031);
xnor U30348 (N_30348,N_29482,N_28499);
and U30349 (N_30349,N_28199,N_29782);
nand U30350 (N_30350,N_29927,N_29735);
and U30351 (N_30351,N_29250,N_29417);
xnor U30352 (N_30352,N_28339,N_27564);
nor U30353 (N_30353,N_29747,N_29002);
nand U30354 (N_30354,N_28110,N_28174);
nand U30355 (N_30355,N_28739,N_28313);
or U30356 (N_30356,N_29035,N_28348);
xor U30357 (N_30357,N_28656,N_28039);
nor U30358 (N_30358,N_27828,N_29506);
and U30359 (N_30359,N_28182,N_29957);
nand U30360 (N_30360,N_29097,N_27881);
nor U30361 (N_30361,N_27613,N_29892);
xor U30362 (N_30362,N_29525,N_28166);
and U30363 (N_30363,N_28806,N_28456);
nand U30364 (N_30364,N_28357,N_27769);
xor U30365 (N_30365,N_28352,N_29512);
nor U30366 (N_30366,N_28303,N_28761);
nor U30367 (N_30367,N_27780,N_29650);
xor U30368 (N_30368,N_27597,N_28035);
nor U30369 (N_30369,N_29640,N_29403);
and U30370 (N_30370,N_27580,N_28780);
and U30371 (N_30371,N_29529,N_27915);
nand U30372 (N_30372,N_28021,N_28460);
nor U30373 (N_30373,N_28511,N_27790);
nand U30374 (N_30374,N_28687,N_28299);
and U30375 (N_30375,N_27648,N_27731);
or U30376 (N_30376,N_29337,N_28028);
nor U30377 (N_30377,N_27813,N_27504);
and U30378 (N_30378,N_29949,N_29850);
and U30379 (N_30379,N_28872,N_29677);
nand U30380 (N_30380,N_27902,N_29036);
xor U30381 (N_30381,N_28421,N_28657);
or U30382 (N_30382,N_27767,N_28469);
or U30383 (N_30383,N_28852,N_29992);
and U30384 (N_30384,N_28880,N_27916);
or U30385 (N_30385,N_28341,N_29965);
nor U30386 (N_30386,N_29118,N_28047);
xnor U30387 (N_30387,N_29202,N_28686);
nor U30388 (N_30388,N_29149,N_27644);
nor U30389 (N_30389,N_28728,N_27634);
and U30390 (N_30390,N_27756,N_28309);
and U30391 (N_30391,N_27520,N_28554);
nand U30392 (N_30392,N_29631,N_27617);
nor U30393 (N_30393,N_27958,N_29498);
and U30394 (N_30394,N_29941,N_28446);
nor U30395 (N_30395,N_28152,N_28544);
or U30396 (N_30396,N_29428,N_29976);
and U30397 (N_30397,N_27960,N_29477);
nand U30398 (N_30398,N_29908,N_27903);
nor U30399 (N_30399,N_28843,N_27736);
nand U30400 (N_30400,N_29347,N_28992);
and U30401 (N_30401,N_28574,N_28015);
nand U30402 (N_30402,N_27733,N_27823);
and U30403 (N_30403,N_27727,N_28004);
nor U30404 (N_30404,N_29373,N_27796);
or U30405 (N_30405,N_29312,N_28975);
or U30406 (N_30406,N_27667,N_27877);
nor U30407 (N_30407,N_28288,N_27853);
xor U30408 (N_30408,N_28069,N_27514);
nor U30409 (N_30409,N_29226,N_29510);
xor U30410 (N_30410,N_28628,N_27872);
or U30411 (N_30411,N_29646,N_29845);
nand U30412 (N_30412,N_28821,N_28132);
xnor U30413 (N_30413,N_28702,N_29115);
xnor U30414 (N_30414,N_28560,N_29390);
or U30415 (N_30415,N_28864,N_29885);
and U30416 (N_30416,N_28789,N_28524);
nand U30417 (N_30417,N_28766,N_27620);
nor U30418 (N_30418,N_29180,N_28296);
and U30419 (N_30419,N_29194,N_29480);
nor U30420 (N_30420,N_29999,N_29604);
or U30421 (N_30421,N_28381,N_27889);
or U30422 (N_30422,N_27807,N_29744);
nand U30423 (N_30423,N_29541,N_28076);
nor U30424 (N_30424,N_28202,N_27990);
nand U30425 (N_30425,N_28693,N_28312);
and U30426 (N_30426,N_27969,N_28065);
xor U30427 (N_30427,N_29535,N_27707);
or U30428 (N_30428,N_28748,N_29910);
xor U30429 (N_30429,N_28001,N_28707);
and U30430 (N_30430,N_28377,N_28548);
xnor U30431 (N_30431,N_28082,N_27808);
nor U30432 (N_30432,N_29124,N_28925);
xnor U30433 (N_30433,N_29426,N_29320);
nand U30434 (N_30434,N_28726,N_28213);
and U30435 (N_30435,N_29627,N_29820);
or U30436 (N_30436,N_28995,N_27724);
nor U30437 (N_30437,N_29107,N_27523);
and U30438 (N_30438,N_28103,N_29979);
xnor U30439 (N_30439,N_29524,N_28814);
and U30440 (N_30440,N_29375,N_28123);
nand U30441 (N_30441,N_29494,N_29644);
or U30442 (N_30442,N_28452,N_28052);
nor U30443 (N_30443,N_28197,N_27687);
or U30444 (N_30444,N_28275,N_29262);
xor U30445 (N_30445,N_29092,N_28416);
or U30446 (N_30446,N_29971,N_29274);
or U30447 (N_30447,N_28763,N_29170);
nor U30448 (N_30448,N_29688,N_29139);
xor U30449 (N_30449,N_29327,N_29398);
and U30450 (N_30450,N_29365,N_29109);
and U30451 (N_30451,N_29323,N_27851);
or U30452 (N_30452,N_28411,N_28985);
xor U30453 (N_30453,N_27883,N_28148);
xor U30454 (N_30454,N_28136,N_28691);
and U30455 (N_30455,N_29224,N_29113);
or U30456 (N_30456,N_29329,N_28645);
nor U30457 (N_30457,N_29780,N_28904);
nand U30458 (N_30458,N_29475,N_28597);
and U30459 (N_30459,N_29414,N_28631);
nor U30460 (N_30460,N_29127,N_27891);
nor U30461 (N_30461,N_29467,N_29071);
nor U30462 (N_30462,N_27785,N_28886);
nand U30463 (N_30463,N_28316,N_28059);
and U30464 (N_30464,N_29010,N_29652);
nand U30465 (N_30465,N_29689,N_28802);
xor U30466 (N_30466,N_28378,N_27801);
and U30467 (N_30467,N_28613,N_29217);
xnor U30468 (N_30468,N_27690,N_28865);
and U30469 (N_30469,N_28098,N_28623);
or U30470 (N_30470,N_29135,N_29684);
nand U30471 (N_30471,N_29479,N_28327);
and U30472 (N_30472,N_29073,N_27611);
nor U30473 (N_30473,N_27608,N_28032);
and U30474 (N_30474,N_29258,N_29241);
nand U30475 (N_30475,N_29571,N_27726);
xor U30476 (N_30476,N_29366,N_28750);
nand U30477 (N_30477,N_29526,N_29503);
nand U30478 (N_30478,N_28467,N_28368);
xnor U30479 (N_30479,N_28422,N_29111);
nand U30480 (N_30480,N_29551,N_29169);
xor U30481 (N_30481,N_27592,N_27689);
xor U30482 (N_30482,N_29154,N_27873);
or U30483 (N_30483,N_29926,N_27513);
nand U30484 (N_30484,N_28783,N_27923);
xnor U30485 (N_30485,N_28977,N_29204);
and U30486 (N_30486,N_28463,N_28306);
and U30487 (N_30487,N_28907,N_29379);
or U30488 (N_30488,N_28978,N_29974);
nor U30489 (N_30489,N_29668,N_28605);
and U30490 (N_30490,N_28387,N_29376);
or U30491 (N_30491,N_27540,N_28871);
nor U30492 (N_30492,N_28160,N_28251);
nor U30493 (N_30493,N_29497,N_29421);
nand U30494 (N_30494,N_29047,N_28277);
nor U30495 (N_30495,N_29846,N_28923);
or U30496 (N_30496,N_28618,N_27833);
and U30497 (N_30497,N_27809,N_29063);
and U30498 (N_30498,N_27927,N_29849);
nor U30499 (N_30499,N_27860,N_29635);
xor U30500 (N_30500,N_28782,N_29430);
or U30501 (N_30501,N_29517,N_27723);
and U30502 (N_30502,N_28757,N_28730);
or U30503 (N_30503,N_27627,N_28561);
or U30504 (N_30504,N_29876,N_27750);
nor U30505 (N_30505,N_28829,N_27624);
xor U30506 (N_30506,N_28959,N_29767);
and U30507 (N_30507,N_29916,N_28315);
nor U30508 (N_30508,N_27983,N_28483);
nand U30509 (N_30509,N_27897,N_29612);
and U30510 (N_30510,N_29095,N_29453);
and U30511 (N_30511,N_29637,N_29141);
nand U30512 (N_30512,N_27605,N_28547);
nor U30513 (N_30513,N_29853,N_28228);
nand U30514 (N_30514,N_29056,N_27541);
and U30515 (N_30515,N_29350,N_29593);
and U30516 (N_30516,N_29920,N_28255);
xnor U30517 (N_30517,N_28710,N_28068);
xor U30518 (N_30518,N_29729,N_29024);
xnor U30519 (N_30519,N_27646,N_27973);
nand U30520 (N_30520,N_29416,N_28529);
and U30521 (N_30521,N_29282,N_27738);
or U30522 (N_30522,N_27728,N_27595);
or U30523 (N_30523,N_28913,N_29133);
or U30524 (N_30524,N_28311,N_28787);
nand U30525 (N_30525,N_28464,N_29116);
nor U30526 (N_30526,N_28964,N_29772);
nor U30527 (N_30527,N_29049,N_27711);
nand U30528 (N_30528,N_28196,N_27729);
and U30529 (N_30529,N_29563,N_28753);
and U30530 (N_30530,N_29072,N_27910);
nand U30531 (N_30531,N_27568,N_29055);
xnor U30532 (N_30532,N_29448,N_28563);
xnor U30533 (N_30533,N_28366,N_29607);
and U30534 (N_30534,N_27566,N_28643);
xor U30535 (N_30535,N_29947,N_28803);
nand U30536 (N_30536,N_29715,N_29394);
nor U30537 (N_30537,N_29245,N_29867);
nor U30538 (N_30538,N_27614,N_27834);
or U30539 (N_30539,N_28382,N_29157);
xnor U30540 (N_30540,N_28608,N_29424);
or U30541 (N_30541,N_28917,N_28485);
xor U30542 (N_30542,N_27908,N_29819);
nor U30543 (N_30543,N_28607,N_29096);
nand U30544 (N_30544,N_27735,N_29136);
nand U30545 (N_30545,N_29938,N_28811);
nand U30546 (N_30546,N_29419,N_29469);
or U30547 (N_30547,N_27814,N_27914);
nand U30548 (N_30548,N_28119,N_27576);
xor U30549 (N_30549,N_29629,N_27635);
nand U30550 (N_30550,N_29922,N_28636);
nor U30551 (N_30551,N_28232,N_27616);
nor U30552 (N_30552,N_29628,N_29815);
nor U30553 (N_30553,N_28905,N_28279);
xnor U30554 (N_30554,N_29175,N_27665);
nor U30555 (N_30555,N_29564,N_29520);
and U30556 (N_30556,N_29285,N_28724);
or U30557 (N_30557,N_28376,N_29661);
nand U30558 (N_30558,N_29174,N_28663);
nand U30559 (N_30559,N_29624,N_29295);
or U30560 (N_30560,N_29314,N_28805);
xnor U30561 (N_30561,N_28142,N_29371);
nor U30562 (N_30562,N_27512,N_28235);
xnor U30563 (N_30563,N_28354,N_29942);
nand U30564 (N_30564,N_28967,N_29184);
nor U30565 (N_30565,N_28045,N_29580);
or U30566 (N_30566,N_29763,N_29913);
and U30567 (N_30567,N_27812,N_29131);
xor U30568 (N_30568,N_28935,N_28562);
nor U30569 (N_30569,N_28233,N_29860);
or U30570 (N_30570,N_29330,N_28545);
nor U30571 (N_30571,N_28972,N_29132);
or U30572 (N_30572,N_28176,N_28037);
nor U30573 (N_30573,N_27717,N_27652);
or U30574 (N_30574,N_28719,N_28698);
nor U30575 (N_30575,N_28391,N_29804);
or U30576 (N_30576,N_28187,N_28109);
and U30577 (N_30577,N_28432,N_27550);
nor U30578 (N_30578,N_27664,N_28475);
and U30579 (N_30579,N_29098,N_27842);
nor U30580 (N_30580,N_28881,N_28633);
nand U30581 (N_30581,N_27838,N_29951);
xor U30582 (N_30582,N_29649,N_28833);
nand U30583 (N_30583,N_29573,N_27571);
and U30584 (N_30584,N_28818,N_27700);
xor U30585 (N_30585,N_28238,N_29732);
xor U30586 (N_30586,N_28874,N_28191);
nand U30587 (N_30587,N_27961,N_28267);
nand U30588 (N_30588,N_27538,N_28866);
xor U30589 (N_30589,N_28321,N_29384);
nor U30590 (N_30590,N_28741,N_27673);
nor U30591 (N_30591,N_28828,N_27947);
or U30592 (N_30592,N_29445,N_29310);
and U30593 (N_30593,N_29088,N_28362);
nor U30594 (N_30594,N_28655,N_28388);
nor U30595 (N_30595,N_27928,N_27888);
xnor U30596 (N_30596,N_29792,N_28962);
or U30597 (N_30597,N_28532,N_28470);
xnor U30598 (N_30598,N_28734,N_29447);
and U30599 (N_30599,N_28575,N_28549);
nor U30600 (N_30600,N_29364,N_28477);
and U30601 (N_30601,N_29061,N_28749);
or U30602 (N_30602,N_29328,N_29287);
or U30603 (N_30603,N_28175,N_29589);
and U30604 (N_30604,N_29050,N_29921);
or U30605 (N_30605,N_28909,N_28928);
nor U30606 (N_30606,N_29466,N_28944);
xor U30607 (N_30607,N_29158,N_29968);
nor U30608 (N_30608,N_29338,N_28515);
and U30609 (N_30609,N_28241,N_29229);
or U30610 (N_30610,N_28040,N_27871);
or U30611 (N_30611,N_27671,N_27941);
nor U30612 (N_30612,N_27784,N_27582);
and U30613 (N_30613,N_28230,N_29206);
xor U30614 (N_30614,N_28479,N_27835);
or U30615 (N_30615,N_28772,N_28482);
nor U30616 (N_30616,N_27995,N_27606);
xor U30617 (N_30617,N_29000,N_27946);
xor U30618 (N_30618,N_29444,N_28108);
xnor U30619 (N_30619,N_28945,N_28705);
and U30620 (N_30620,N_29761,N_29134);
and U30621 (N_30621,N_27588,N_29771);
xor U30622 (N_30622,N_28779,N_28998);
nor U30623 (N_30623,N_29011,N_27870);
nor U30624 (N_30624,N_28294,N_29493);
and U30625 (N_30625,N_29288,N_27556);
nor U30626 (N_30626,N_28914,N_28493);
nor U30627 (N_30627,N_28541,N_27638);
nor U30628 (N_30628,N_29696,N_27630);
or U30629 (N_30629,N_28650,N_28314);
and U30630 (N_30630,N_29858,N_27692);
nand U30631 (N_30631,N_27722,N_27688);
or U30632 (N_30632,N_28523,N_27803);
nor U30633 (N_30633,N_27956,N_29212);
or U30634 (N_30634,N_27855,N_28157);
and U30635 (N_30635,N_27594,N_29615);
xnor U30636 (N_30636,N_28024,N_29432);
and U30637 (N_30637,N_29844,N_29391);
xor U30638 (N_30638,N_28740,N_29290);
xor U30639 (N_30639,N_29486,N_29253);
and U30640 (N_30640,N_29754,N_28396);
nand U30641 (N_30641,N_28014,N_29006);
nor U30642 (N_30642,N_28679,N_28768);
and U30643 (N_30643,N_27940,N_28002);
nand U30644 (N_30644,N_29700,N_29725);
nand U30645 (N_30645,N_28224,N_27968);
nor U30646 (N_30646,N_29007,N_29341);
or U30647 (N_30647,N_27537,N_28883);
xor U30648 (N_30648,N_27768,N_29753);
nand U30649 (N_30649,N_29013,N_27972);
or U30650 (N_30650,N_29368,N_28825);
nand U30651 (N_30651,N_29294,N_27589);
and U30652 (N_30652,N_29363,N_27524);
or U30653 (N_30653,N_29222,N_28901);
nor U30654 (N_30654,N_27997,N_28776);
nand U30655 (N_30655,N_28085,N_28556);
and U30656 (N_30656,N_29760,N_29680);
or U30657 (N_30657,N_28165,N_27984);
or U30658 (N_30658,N_28557,N_27552);
nand U30659 (N_30659,N_29296,N_28990);
or U30660 (N_30660,N_27744,N_29322);
and U30661 (N_30661,N_29476,N_28659);
and U30662 (N_30662,N_28210,N_28214);
and U30663 (N_30663,N_27830,N_28622);
xnor U30664 (N_30664,N_27577,N_28521);
and U30665 (N_30665,N_28029,N_29599);
xnor U30666 (N_30666,N_28697,N_28484);
xor U30667 (N_30667,N_28804,N_29572);
nor U30668 (N_30668,N_29381,N_29388);
or U30669 (N_30669,N_29062,N_27825);
xnor U30670 (N_30670,N_29711,N_28777);
nor U30671 (N_30671,N_28384,N_28717);
or U30672 (N_30672,N_28153,N_27547);
or U30673 (N_30673,N_28667,N_29472);
nor U30674 (N_30674,N_28680,N_29119);
or U30675 (N_30675,N_29958,N_29411);
nor U30676 (N_30676,N_28459,N_27849);
nor U30677 (N_30677,N_29825,N_27721);
and U30678 (N_30678,N_28638,N_29713);
and U30679 (N_30679,N_28512,N_29838);
xor U30680 (N_30680,N_27852,N_27586);
nand U30681 (N_30681,N_27752,N_28055);
xnor U30682 (N_30682,N_28334,N_27740);
and U30683 (N_30683,N_28932,N_29832);
nand U30684 (N_30684,N_29016,N_29064);
nor U30685 (N_30685,N_29722,N_29905);
xnor U30686 (N_30686,N_28927,N_29939);
nor U30687 (N_30687,N_29235,N_29779);
xor U30688 (N_30688,N_29038,N_27848);
nor U30689 (N_30689,N_28644,N_29952);
or U30690 (N_30690,N_29931,N_28017);
xnor U30691 (N_30691,N_29490,N_29270);
nand U30692 (N_30692,N_28877,N_29736);
nand U30693 (N_30693,N_27945,N_28444);
nor U30694 (N_30694,N_29836,N_28875);
and U30695 (N_30695,N_29435,N_28520);
xnor U30696 (N_30696,N_28301,N_28257);
and U30697 (N_30697,N_27636,N_29909);
xnor U30698 (N_30698,N_27971,N_28451);
or U30699 (N_30699,N_27952,N_28180);
nand U30700 (N_30700,N_29343,N_29675);
and U30701 (N_30701,N_28415,N_28091);
nor U30702 (N_30702,N_28672,N_29233);
nand U30703 (N_30703,N_29151,N_29283);
or U30704 (N_30704,N_29499,N_29911);
xor U30705 (N_30705,N_28018,N_28364);
or U30706 (N_30706,N_28572,N_28754);
and U30707 (N_30707,N_29460,N_28184);
nand U30708 (N_30708,N_28480,N_29621);
nand U30709 (N_30709,N_28527,N_28799);
nor U30710 (N_30710,N_29481,N_28038);
xor U30711 (N_30711,N_27602,N_27837);
xnor U30712 (N_30712,N_27791,N_27612);
or U30713 (N_30713,N_29955,N_27659);
nand U30714 (N_30714,N_29353,N_28061);
xnor U30715 (N_30715,N_29369,N_27757);
and U30716 (N_30716,N_27970,N_29352);
and U30717 (N_30717,N_27980,N_27562);
nor U30718 (N_30718,N_28582,N_28139);
nand U30719 (N_30719,N_28131,N_27501);
and U30720 (N_30720,N_29620,N_27779);
nand U30721 (N_30721,N_27963,N_29516);
nor U30722 (N_30722,N_28162,N_28133);
xnor U30723 (N_30723,N_28538,N_29501);
xor U30724 (N_30724,N_27536,N_27766);
or U30725 (N_30725,N_28973,N_27773);
and U30726 (N_30726,N_27782,N_29458);
xor U30727 (N_30727,N_29996,N_28008);
nand U30728 (N_30728,N_28380,N_28426);
or U30729 (N_30729,N_27682,N_29898);
or U30730 (N_30730,N_28960,N_29919);
or U30731 (N_30731,N_28591,N_27818);
or U30732 (N_30732,N_29657,N_28849);
xnor U30733 (N_30733,N_27662,N_27977);
nor U30734 (N_30734,N_27534,N_28370);
or U30735 (N_30735,N_29418,N_29457);
and U30736 (N_30736,N_29090,N_27918);
nand U30737 (N_30737,N_28245,N_28181);
or U30738 (N_30738,N_28770,N_29893);
nand U30739 (N_30739,N_28674,N_28731);
nand U30740 (N_30740,N_28427,N_28942);
or U30741 (N_30741,N_29144,N_29841);
nand U30742 (N_30742,N_27789,N_29625);
nand U30743 (N_30743,N_28333,N_27864);
and U30744 (N_30744,N_29705,N_27548);
and U30745 (N_30745,N_28892,N_27522);
xor U30746 (N_30746,N_27573,N_28543);
xnor U30747 (N_30747,N_28742,N_29104);
nand U30748 (N_30748,N_27619,N_27545);
or U30749 (N_30749,N_28078,N_28077);
nor U30750 (N_30750,N_29443,N_29719);
and U30751 (N_30751,N_29060,N_28669);
nand U30752 (N_30752,N_28425,N_29693);
or U30753 (N_30753,N_28101,N_27674);
or U30754 (N_30754,N_29089,N_29261);
xnor U30755 (N_30755,N_29209,N_28429);
and U30756 (N_30756,N_27765,N_27747);
and U30757 (N_30757,N_28145,N_28383);
xnor U30758 (N_30758,N_28343,N_29507);
nand U30759 (N_30759,N_28013,N_28801);
nor U30760 (N_30760,N_28056,N_29769);
nand U30761 (N_30761,N_27933,N_29234);
nor U30762 (N_30762,N_28223,N_27585);
and U30763 (N_30763,N_29768,N_29960);
nand U30764 (N_30764,N_28473,N_29324);
or U30765 (N_30765,N_28106,N_29492);
or U30766 (N_30766,N_29334,N_29137);
or U30767 (N_30767,N_28458,N_29901);
xor U30768 (N_30768,N_28353,N_29236);
nor U30769 (N_30769,N_27948,N_29359);
nor U30770 (N_30770,N_29102,N_28738);
nor U30771 (N_30771,N_29277,N_28058);
and U30772 (N_30772,N_28592,N_27904);
nor U30773 (N_30773,N_28026,N_27542);
xnor U30774 (N_30774,N_27810,N_28735);
or U30775 (N_30775,N_29873,N_27699);
nor U30776 (N_30776,N_29191,N_28571);
and U30777 (N_30777,N_27857,N_27593);
and U30778 (N_30778,N_28952,N_29200);
xnor U30779 (N_30779,N_27732,N_29861);
nor U30780 (N_30780,N_28637,N_29168);
nand U30781 (N_30781,N_27658,N_28600);
xor U30782 (N_30782,N_27900,N_28594);
and U30783 (N_30783,N_28537,N_28486);
nand U30784 (N_30784,N_27920,N_29988);
or U30785 (N_30785,N_28093,N_29833);
xor U30786 (N_30786,N_29626,N_29008);
nand U30787 (N_30787,N_29150,N_28700);
xor U30788 (N_30788,N_28064,N_28658);
or U30789 (N_30789,N_28794,N_29963);
nand U30790 (N_30790,N_29575,N_28088);
nor U30791 (N_30791,N_29004,N_28057);
or U30792 (N_30792,N_28030,N_28850);
and U30793 (N_30793,N_28769,N_29536);
or U30794 (N_30794,N_29663,N_27669);
xor U30795 (N_30795,N_29521,N_27683);
nand U30796 (N_30796,N_28134,N_28281);
or U30797 (N_30797,N_29101,N_29877);
nor U30798 (N_30798,N_28465,N_29389);
or U30799 (N_30799,N_29189,N_28634);
nand U30800 (N_30800,N_28027,N_29890);
and U30801 (N_30801,N_28434,N_28919);
nor U30802 (N_30802,N_28558,N_28173);
nand U30803 (N_30803,N_29587,N_29566);
or U30804 (N_30804,N_27976,N_28934);
nand U30805 (N_30805,N_29439,N_27618);
or U30806 (N_30806,N_28481,N_27521);
or U30807 (N_30807,N_29275,N_27703);
xor U30808 (N_30808,N_29361,N_29332);
nand U30809 (N_30809,N_29716,N_29001);
and U30810 (N_30810,N_29822,N_28819);
and U30811 (N_30811,N_29075,N_28899);
nor U30812 (N_30812,N_29112,N_29775);
or U30813 (N_30813,N_29546,N_27631);
xor U30814 (N_30814,N_29883,N_29904);
or U30815 (N_30815,N_29923,N_28271);
xnor U30816 (N_30816,N_27565,N_29933);
xor U30817 (N_30817,N_29333,N_29171);
xnor U30818 (N_30818,N_28399,N_27987);
nor U30819 (N_30819,N_28149,N_29033);
xor U30820 (N_30820,N_27942,N_27929);
and U30821 (N_30821,N_29756,N_27826);
or U30822 (N_30822,N_28868,N_27709);
and U30823 (N_30823,N_29724,N_27831);
nor U30824 (N_30824,N_29809,N_28194);
xor U30825 (N_30825,N_28094,N_28454);
or U30826 (N_30826,N_29582,N_28854);
xnor U30827 (N_30827,N_29972,N_28878);
xor U30828 (N_30828,N_29248,N_28890);
nor U30829 (N_30829,N_29348,N_27693);
xor U30830 (N_30830,N_29834,N_28851);
nand U30831 (N_30831,N_29989,N_29527);
nand U30832 (N_30832,N_28372,N_29238);
nand U30833 (N_30833,N_27596,N_29776);
nand U30834 (N_30834,N_29058,N_28662);
xnor U30835 (N_30835,N_29843,N_27884);
xor U30836 (N_30836,N_28125,N_29528);
and U30837 (N_30837,N_29304,N_29440);
nand U30838 (N_30838,N_29230,N_28095);
nor U30839 (N_30839,N_29895,N_28505);
and U30840 (N_30840,N_28873,N_29728);
or U30841 (N_30841,N_28564,N_28345);
nor U30842 (N_30842,N_29456,N_28996);
nor U30843 (N_30843,N_28746,N_27599);
and U30844 (N_30844,N_29318,N_29193);
and U30845 (N_30845,N_27917,N_27771);
xnor U30846 (N_30846,N_28323,N_27974);
or U30847 (N_30847,N_29319,N_27503);
or U30848 (N_30848,N_29925,N_28784);
nand U30849 (N_30849,N_28090,N_28888);
or U30850 (N_30850,N_28947,N_29550);
xnor U30851 (N_30851,N_29609,N_28161);
and U30852 (N_30852,N_28217,N_27832);
or U30853 (N_30853,N_27879,N_28598);
xor U30854 (N_30854,N_28266,N_29272);
and U30855 (N_30855,N_28178,N_29591);
xnor U30856 (N_30856,N_28487,N_27600);
or U30857 (N_30857,N_29651,N_28603);
or U30858 (N_30858,N_27583,N_29496);
nor U30859 (N_30859,N_27640,N_28767);
nor U30860 (N_30860,N_28599,N_28263);
nand U30861 (N_30861,N_29806,N_29872);
or U30862 (N_30862,N_27581,N_29485);
xor U30863 (N_30863,N_29313,N_28689);
xor U30864 (N_30864,N_28648,N_28666);
nand U30865 (N_30865,N_29561,N_29975);
nor U30866 (N_30866,N_28462,N_29679);
xnor U30867 (N_30867,N_27775,N_27654);
xnor U30868 (N_30868,N_29265,N_27787);
and U30869 (N_30869,N_28177,N_29269);
and U30870 (N_30870,N_29737,N_27937);
xnor U30871 (N_30871,N_28540,N_28827);
xor U30872 (N_30872,N_28830,N_28150);
and U30873 (N_30873,N_28147,N_28737);
and U30874 (N_30874,N_28861,N_29291);
and U30875 (N_30875,N_29146,N_28619);
nand U30876 (N_30876,N_29602,N_29160);
and U30877 (N_30877,N_28066,N_28453);
and U30878 (N_30878,N_28845,N_29223);
or U30879 (N_30879,N_28414,N_27955);
nand U30880 (N_30880,N_28398,N_29220);
nor U30881 (N_30881,N_29039,N_28163);
or U30882 (N_30882,N_28590,N_29455);
nor U30883 (N_30883,N_28834,N_28046);
nor U30884 (N_30884,N_28810,N_28513);
nand U30885 (N_30885,N_28798,N_29286);
and U30886 (N_30886,N_29083,N_29986);
xnor U30887 (N_30887,N_29936,N_29405);
xnor U30888 (N_30888,N_27890,N_28438);
nor U30889 (N_30889,N_27930,N_28514);
nor U30890 (N_30890,N_29953,N_28926);
nand U30891 (N_30891,N_29100,N_29438);
nand U30892 (N_30892,N_28503,N_29020);
nand U30893 (N_30893,N_27553,N_29802);
or U30894 (N_30894,N_28272,N_27572);
nand U30895 (N_30895,N_28937,N_29068);
or U30896 (N_30896,N_28870,N_28781);
and U30897 (N_30897,N_29256,N_28550);
xnor U30898 (N_30898,N_29633,N_29354);
or U30899 (N_30899,N_28604,N_29415);
xnor U30900 (N_30900,N_27637,N_28681);
xnor U30901 (N_30901,N_29586,N_29362);
xor U30902 (N_30902,N_27742,N_27762);
and U30903 (N_30903,N_27591,N_28910);
nor U30904 (N_30904,N_28836,N_29301);
and U30905 (N_30905,N_29643,N_29018);
or U30906 (N_30906,N_27867,N_28100);
and U30907 (N_30907,N_29855,N_28921);
nor U30908 (N_30908,N_27781,N_29335);
nand U30909 (N_30909,N_28884,N_29478);
xor U30910 (N_30910,N_28668,N_29306);
and U30911 (N_30911,N_28340,N_28342);
and U30912 (N_30912,N_27846,N_29533);
nor U30913 (N_30913,N_28795,N_29268);
or U30914 (N_30914,N_29632,N_28609);
nor U30915 (N_30915,N_29886,N_29382);
or U30916 (N_30916,N_28951,N_29790);
xor U30917 (N_30917,N_29357,N_28420);
and U30918 (N_30918,N_29367,N_27633);
and U30919 (N_30919,N_28375,N_27986);
nor U30920 (N_30920,N_28007,N_27795);
and U30921 (N_30921,N_28468,N_28307);
xnor U30922 (N_30922,N_29617,N_28496);
and U30923 (N_30923,N_29315,N_29590);
xnor U30924 (N_30924,N_28204,N_29569);
nor U30925 (N_30925,N_29117,N_29317);
or U30926 (N_30926,N_29188,N_27753);
or U30927 (N_30927,N_28409,N_27531);
and U30928 (N_30928,N_28374,N_29091);
nand U30929 (N_30929,N_28855,N_29232);
and U30930 (N_30930,N_29392,N_29749);
nand U30931 (N_30931,N_29356,N_28602);
nand U30932 (N_30932,N_29164,N_29681);
xnor U30933 (N_30933,N_28304,N_27850);
nand U30934 (N_30934,N_29185,N_29870);
nand U30935 (N_30935,N_29534,N_27710);
and U30936 (N_30936,N_29377,N_28641);
or U30937 (N_30937,N_27806,N_28356);
nand U30938 (N_30938,N_28265,N_28522);
xnor U30939 (N_30939,N_28654,N_28745);
or U30940 (N_30940,N_28244,N_28506);
nand U30941 (N_30941,N_27704,N_29616);
or U30942 (N_30942,N_29808,N_28478);
and U30943 (N_30943,N_28141,N_28397);
or U30944 (N_30944,N_29046,N_27598);
and U30945 (N_30945,N_29837,N_28922);
nor U30946 (N_30946,N_28405,N_28198);
nor U30947 (N_30947,N_29848,N_27558);
xnor U30948 (N_30948,N_29293,N_28882);
or U30949 (N_30949,N_28440,N_27800);
and U30950 (N_30950,N_28832,N_27998);
xnor U30951 (N_30951,N_29659,N_29452);
xor U30952 (N_30952,N_29162,N_28517);
xnor U30953 (N_30953,N_29891,N_29600);
or U30954 (N_30954,N_27854,N_28510);
and U30955 (N_30955,N_29954,N_28612);
and U30956 (N_30956,N_29239,N_29549);
xor U30957 (N_30957,N_27869,N_29215);
nor U30958 (N_30958,N_29321,N_27868);
nor U30959 (N_30959,N_28379,N_27865);
or U30960 (N_30960,N_28071,N_29031);
xnor U30961 (N_30961,N_27622,N_29198);
xnor U30962 (N_30962,N_29690,N_27931);
xnor U30963 (N_30963,N_28424,N_28107);
xor U30964 (N_30964,N_28508,N_29682);
or U30965 (N_30965,N_29896,N_29672);
nor U30966 (N_30966,N_28273,N_28250);
xor U30967 (N_30967,N_28856,N_29130);
xor U30968 (N_30968,N_28466,N_29252);
or U30969 (N_30969,N_29029,N_28751);
nand U30970 (N_30970,N_28664,N_28488);
nor U30971 (N_30971,N_28987,N_28005);
xnor U30972 (N_30972,N_29451,N_28688);
xnor U30973 (N_30973,N_28063,N_28684);
xor U30974 (N_30974,N_27866,N_28695);
xnor U30975 (N_30975,N_28902,N_28762);
or U30976 (N_30976,N_27604,N_28318);
xnor U30977 (N_30977,N_29831,N_29894);
nand U30978 (N_30978,N_27508,N_29813);
nor U30979 (N_30979,N_28570,N_28898);
nor U30980 (N_30980,N_28104,N_28206);
nor U30981 (N_30981,N_29810,N_27507);
and U30982 (N_30982,N_28346,N_28838);
or U30983 (N_30983,N_27666,N_28305);
and U30984 (N_30984,N_29730,N_28127);
and U30985 (N_30985,N_28790,N_29906);
or U30986 (N_30986,N_29596,N_28200);
xnor U30987 (N_30987,N_28122,N_28555);
nor U30988 (N_30988,N_29123,N_28070);
and U30989 (N_30989,N_28685,N_29441);
xor U30990 (N_30990,N_28472,N_27817);
nand U30991 (N_30991,N_28976,N_28993);
nor U30992 (N_30992,N_28876,N_29537);
and U30993 (N_30993,N_28044,N_29395);
or U30994 (N_30994,N_29887,N_29186);
and U30995 (N_30995,N_27772,N_28893);
xnor U30996 (N_30996,N_27528,N_29727);
nand U30997 (N_30997,N_28601,N_28569);
nand U30998 (N_30998,N_27896,N_28813);
xnor U30999 (N_30999,N_28351,N_28800);
nor U31000 (N_31000,N_29800,N_28611);
nor U31001 (N_31001,N_27887,N_28435);
or U31002 (N_31002,N_28566,N_29489);
and U31003 (N_31003,N_28621,N_29685);
nand U31004 (N_31004,N_28670,N_28115);
or U31005 (N_31005,N_28219,N_28894);
nand U31006 (N_31006,N_29402,N_27856);
nand U31007 (N_31007,N_29985,N_29698);
xor U31008 (N_31008,N_28300,N_28788);
and U31009 (N_31009,N_28536,N_29930);
nand U31010 (N_31010,N_29197,N_28720);
or U31011 (N_31011,N_28982,N_28168);
nand U31012 (N_31012,N_28863,N_29797);
nor U31013 (N_31013,N_28036,N_28755);
or U31014 (N_31014,N_29701,N_27684);
or U31015 (N_31015,N_28671,N_29984);
nor U31016 (N_31016,N_29859,N_28450);
or U31017 (N_31017,N_27950,N_29052);
or U31018 (N_31018,N_28009,N_27626);
or U31019 (N_31019,N_28385,N_28319);
xnor U31020 (N_31020,N_28677,N_28011);
nor U31021 (N_31021,N_27661,N_27714);
xor U31022 (N_31022,N_28268,N_29748);
or U31023 (N_31023,N_29308,N_29670);
or U31024 (N_31024,N_29781,N_29145);
xnor U31025 (N_31025,N_29660,N_28721);
nor U31026 (N_31026,N_28808,N_29192);
nand U31027 (N_31027,N_28025,N_27805);
xor U31028 (N_31028,N_29346,N_28404);
nand U31029 (N_31029,N_28418,N_29143);
xnor U31030 (N_31030,N_29793,N_29829);
xor U31031 (N_31031,N_29839,N_28283);
nand U31032 (N_31032,N_27993,N_28359);
xnor U31033 (N_31033,N_28736,N_29297);
nor U31034 (N_31034,N_28635,N_29671);
and U31035 (N_31035,N_29622,N_29959);
and U31036 (N_31036,N_29794,N_28773);
or U31037 (N_31037,N_28924,N_29704);
nor U31038 (N_31038,N_29433,N_29309);
nand U31039 (N_31039,N_29648,N_28956);
nand U31040 (N_31040,N_28172,N_28963);
or U31041 (N_31041,N_29300,N_28447);
nor U31042 (N_31042,N_29079,N_29918);
nor U31043 (N_31043,N_28445,N_28519);
and U31044 (N_31044,N_27657,N_27570);
nor U31045 (N_31045,N_28347,N_28221);
or U31046 (N_31046,N_29934,N_29351);
xor U31047 (N_31047,N_27603,N_29945);
and U31048 (N_31048,N_27746,N_28430);
xor U31049 (N_31049,N_29462,N_29912);
xor U31050 (N_31050,N_27944,N_27559);
or U31051 (N_31051,N_29777,N_28431);
and U31052 (N_31052,N_29183,N_28704);
xnor U31053 (N_31053,N_28344,N_29187);
and U31054 (N_31054,N_28105,N_28111);
xnor U31055 (N_31055,N_27759,N_28760);
or U31056 (N_31056,N_28074,N_28260);
and U31057 (N_31057,N_29881,N_29255);
or U31058 (N_31058,N_27579,N_29231);
xnor U31059 (N_31059,N_29852,N_27590);
nor U31060 (N_31060,N_29851,N_27899);
and U31061 (N_31061,N_28651,N_28067);
and U31062 (N_31062,N_28048,N_27954);
and U31063 (N_31063,N_28713,N_29201);
xor U31064 (N_31064,N_28957,N_28433);
and U31065 (N_31065,N_29303,N_28016);
and U31066 (N_31066,N_27560,N_28439);
nor U31067 (N_31067,N_28203,N_29473);
nand U31068 (N_31068,N_27716,N_28889);
nor U31069 (N_31069,N_28102,N_28552);
and U31070 (N_31070,N_29961,N_28759);
nand U31071 (N_31071,N_27516,N_29943);
and U31072 (N_31072,N_29542,N_29567);
nand U31073 (N_31073,N_29176,N_28577);
nor U31074 (N_31074,N_29179,N_29866);
nor U31075 (N_31075,N_28585,N_29578);
nor U31076 (N_31076,N_28471,N_27798);
nand U31077 (N_31077,N_29783,N_27561);
and U31078 (N_31078,N_27623,N_28653);
xor U31079 (N_31079,N_29022,N_29034);
or U31080 (N_31080,N_28660,N_29408);
and U31081 (N_31081,N_28786,N_29553);
xor U31082 (N_31082,N_28276,N_29244);
or U31083 (N_31083,N_29207,N_28793);
or U31084 (N_31084,N_28812,N_29267);
nand U31085 (N_31085,N_29801,N_29811);
nor U31086 (N_31086,N_28573,N_27843);
xor U31087 (N_31087,N_29242,N_29210);
nand U31088 (N_31088,N_29746,N_29997);
and U31089 (N_31089,N_27696,N_27822);
and U31090 (N_31090,N_29205,N_29504);
xor U31091 (N_31091,N_29880,N_29755);
or U31092 (N_31092,N_29562,N_29140);
xnor U31093 (N_31093,N_27859,N_28535);
xnor U31094 (N_31094,N_29264,N_27672);
or U31095 (N_31095,N_28518,N_28211);
and U31096 (N_31096,N_29167,N_29030);
and U31097 (N_31097,N_28867,N_27776);
nor U31098 (N_31098,N_29739,N_28290);
or U31099 (N_31099,N_29500,N_29057);
xnor U31100 (N_31100,N_28474,N_28796);
nand U31101 (N_31101,N_28831,N_29662);
nand U31102 (N_31102,N_28358,N_29805);
and U31103 (N_31103,N_28792,N_28328);
xnor U31104 (N_31104,N_28154,N_29084);
xnor U31105 (N_31105,N_28525,N_28151);
or U31106 (N_31106,N_27557,N_27745);
nor U31107 (N_31107,N_28006,N_28931);
and U31108 (N_31108,N_29840,N_28771);
xnor U31109 (N_31109,N_28588,N_29907);
xor U31110 (N_31110,N_28994,N_27713);
nand U31111 (N_31111,N_29752,N_29720);
nor U31112 (N_31112,N_29666,N_28360);
xor U31113 (N_31113,N_29459,N_27763);
xor U31114 (N_31114,N_29544,N_29166);
or U31115 (N_31115,N_27811,N_27922);
and U31116 (N_31116,N_29087,N_29249);
xor U31117 (N_31117,N_28930,N_27988);
nand U31118 (N_31118,N_29434,N_29554);
nand U31119 (N_31119,N_28989,N_28991);
xor U31120 (N_31120,N_29254,N_29981);
and U31121 (N_31121,N_29454,N_28361);
nand U31122 (N_31122,N_29019,N_27898);
nand U31123 (N_31123,N_29152,N_28084);
nand U31124 (N_31124,N_29173,N_28974);
and U31125 (N_31125,N_27743,N_29683);
and U31126 (N_31126,N_28373,N_29712);
or U31127 (N_31127,N_29686,N_29009);
xnor U31128 (N_31128,N_28392,N_28970);
and U31129 (N_31129,N_27912,N_29216);
nand U31130 (N_31130,N_28593,N_28050);
nand U31131 (N_31131,N_27526,N_29237);
nor U31132 (N_31132,N_27778,N_27694);
and U31133 (N_31133,N_29129,N_29788);
nor U31134 (N_31134,N_29153,N_27991);
nor U31135 (N_31135,N_29821,N_28785);
nand U31136 (N_31136,N_29519,N_27905);
and U31137 (N_31137,N_28943,N_27925);
nor U31138 (N_31138,N_28595,N_28712);
nand U31139 (N_31139,N_29692,N_29077);
nor U31140 (N_31140,N_29899,N_28114);
nor U31141 (N_31141,N_29349,N_29803);
or U31142 (N_31142,N_28130,N_28916);
nor U31143 (N_31143,N_28948,N_27505);
nand U31144 (N_31144,N_27663,N_27525);
nand U31145 (N_31145,N_27934,N_29882);
and U31146 (N_31146,N_29066,N_28501);
or U31147 (N_31147,N_29027,N_28955);
nand U31148 (N_31148,N_29579,N_28936);
nand U31149 (N_31149,N_27610,N_29142);
and U31150 (N_31150,N_27563,N_29468);
nand U31151 (N_31151,N_29714,N_29110);
or U31152 (N_31152,N_28335,N_27554);
nor U31153 (N_31153,N_29078,N_27783);
nand U31154 (N_31154,N_29214,N_28413);
nor U31155 (N_31155,N_28455,N_27863);
nand U31156 (N_31156,N_29014,N_28282);
nor U31157 (N_31157,N_29437,N_27527);
xor U31158 (N_31158,N_28915,N_29884);
nand U31159 (N_31159,N_29178,N_28403);
xnor U31160 (N_31160,N_27949,N_29208);
nor U31161 (N_31161,N_27861,N_28642);
nor U31162 (N_31162,N_29574,N_29613);
nand U31163 (N_31163,N_29559,N_29545);
nand U31164 (N_31164,N_28080,N_27751);
xor U31165 (N_31165,N_29734,N_29386);
and U31166 (N_31166,N_27601,N_28661);
nand U31167 (N_31167,N_29741,N_27967);
and U31168 (N_31168,N_28287,N_28054);
nand U31169 (N_31169,N_29577,N_29695);
nor U31170 (N_31170,N_28911,N_28033);
nand U31171 (N_31171,N_29874,N_28576);
nand U31172 (N_31172,N_29773,N_28980);
nor U31173 (N_31173,N_29450,N_28559);
or U31174 (N_31174,N_28891,N_29967);
nand U31175 (N_31175,N_28542,N_27677);
nand U31176 (N_31176,N_27725,N_28824);
xor U31177 (N_31177,N_28270,N_27836);
xor U31178 (N_31178,N_27919,N_28879);
nor U31179 (N_31179,N_28903,N_28285);
nand U31180 (N_31180,N_29266,N_28096);
nor U31181 (N_31181,N_29425,N_28526);
or U31182 (N_31182,N_27632,N_28826);
or U31183 (N_31183,N_29412,N_28298);
or U31184 (N_31184,N_28617,N_29718);
nor U31185 (N_31185,N_28820,N_29990);
xnor U31186 (N_31186,N_27844,N_28971);
nand U31187 (N_31187,N_29856,N_29514);
nor U31188 (N_31188,N_28624,N_29998);
xnor U31189 (N_31189,N_28848,N_29588);
or U31190 (N_31190,N_27645,N_28979);
nor U31191 (N_31191,N_29105,N_29059);
nand U31192 (N_31192,N_29396,N_28774);
nand U31193 (N_31193,N_29983,N_27533);
nand U31194 (N_31194,N_28553,N_28489);
nand U31195 (N_31195,N_27695,N_29360);
and U31196 (N_31196,N_28363,N_29726);
nand U31197 (N_31197,N_28159,N_28835);
nor U31198 (N_31198,N_28596,N_28723);
and U31199 (N_31199,N_28395,N_28847);
xor U31200 (N_31200,N_28968,N_27651);
nor U31201 (N_31201,N_27510,N_29924);
nor U31202 (N_31202,N_29993,N_28186);
or U31203 (N_31203,N_29940,N_28823);
xor U31204 (N_31204,N_28534,N_29397);
nor U31205 (N_31205,N_29344,N_27819);
or U31206 (N_31206,N_27660,N_27502);
nor U31207 (N_31207,N_27847,N_28201);
nor U31208 (N_31208,N_28394,N_29125);
nor U31209 (N_31209,N_29765,N_29791);
or U31210 (N_31210,N_28626,N_29897);
or U31211 (N_31211,N_29040,N_28958);
nor U31212 (N_31212,N_29731,N_28949);
or U31213 (N_31213,N_29431,N_28208);
nand U31214 (N_31214,N_28896,N_27698);
or U31215 (N_31215,N_28494,N_28673);
and U31216 (N_31216,N_28533,N_27642);
xnor U31217 (N_31217,N_29043,N_29568);
nand U31218 (N_31218,N_29962,N_28457);
and U31219 (N_31219,N_29508,N_29053);
or U31220 (N_31220,N_28678,N_28289);
nor U31221 (N_31221,N_28441,N_29387);
and U31222 (N_31222,N_29742,N_29673);
or U31223 (N_31223,N_29094,N_28476);
xnor U31224 (N_31224,N_28073,N_29122);
xor U31225 (N_31225,N_28192,N_29463);
or U31226 (N_31226,N_28097,N_29889);
and U31227 (N_31227,N_27720,N_28419);
xor U31228 (N_31228,N_29915,N_27951);
xnor U31229 (N_31229,N_27691,N_27621);
nor U31230 (N_31230,N_29037,N_27964);
nor U31231 (N_31231,N_29051,N_28167);
nor U31232 (N_31232,N_28022,N_29944);
xor U31233 (N_31233,N_28649,N_29565);
and U31234 (N_31234,N_29225,N_29227);
or U31235 (N_31235,N_29165,N_29247);
nand U31236 (N_31236,N_27761,N_29044);
or U31237 (N_31237,N_28986,N_28261);
xor U31238 (N_31238,N_29302,N_28815);
xor U31239 (N_31239,N_28969,N_28332);
or U31240 (N_31240,N_29699,N_29543);
or U31241 (N_31241,N_29610,N_29003);
or U31242 (N_31242,N_29378,N_28144);
nor U31243 (N_31243,N_28676,N_29464);
or U31244 (N_31244,N_27959,N_27893);
and U31245 (N_31245,N_29595,N_27519);
and U31246 (N_31246,N_28722,N_29540);
nor U31247 (N_31247,N_29461,N_27737);
and U31248 (N_31248,N_29080,N_28286);
nor U31249 (N_31249,N_29656,N_29708);
and U31250 (N_31250,N_28099,N_29191);
nor U31251 (N_31251,N_28167,N_28234);
nand U31252 (N_31252,N_29937,N_29801);
nand U31253 (N_31253,N_28353,N_27877);
xor U31254 (N_31254,N_29558,N_29480);
nand U31255 (N_31255,N_28143,N_27634);
or U31256 (N_31256,N_27573,N_29606);
xor U31257 (N_31257,N_27603,N_27887);
nor U31258 (N_31258,N_29352,N_29487);
nor U31259 (N_31259,N_29426,N_28056);
or U31260 (N_31260,N_28892,N_27790);
xnor U31261 (N_31261,N_29715,N_27573);
or U31262 (N_31262,N_29988,N_28230);
or U31263 (N_31263,N_27909,N_28475);
and U31264 (N_31264,N_28605,N_29809);
nor U31265 (N_31265,N_29524,N_28233);
nor U31266 (N_31266,N_28745,N_27617);
nand U31267 (N_31267,N_27919,N_27706);
or U31268 (N_31268,N_27935,N_29068);
or U31269 (N_31269,N_29474,N_27608);
and U31270 (N_31270,N_27837,N_29407);
nand U31271 (N_31271,N_29077,N_28534);
nand U31272 (N_31272,N_29823,N_28820);
or U31273 (N_31273,N_28114,N_28266);
and U31274 (N_31274,N_28731,N_27503);
and U31275 (N_31275,N_29227,N_29032);
nor U31276 (N_31276,N_28400,N_28636);
nand U31277 (N_31277,N_29714,N_28348);
or U31278 (N_31278,N_29993,N_29716);
or U31279 (N_31279,N_29866,N_29621);
nand U31280 (N_31280,N_29511,N_28571);
nor U31281 (N_31281,N_27830,N_28907);
nor U31282 (N_31282,N_28624,N_29722);
or U31283 (N_31283,N_28313,N_29180);
xor U31284 (N_31284,N_29644,N_27581);
nand U31285 (N_31285,N_29360,N_27668);
xnor U31286 (N_31286,N_29871,N_28175);
and U31287 (N_31287,N_29210,N_28361);
xnor U31288 (N_31288,N_28168,N_28609);
and U31289 (N_31289,N_28588,N_28980);
and U31290 (N_31290,N_29537,N_28595);
xnor U31291 (N_31291,N_27712,N_29872);
or U31292 (N_31292,N_27889,N_27730);
or U31293 (N_31293,N_28499,N_29291);
xnor U31294 (N_31294,N_29878,N_27663);
xor U31295 (N_31295,N_27955,N_29500);
nor U31296 (N_31296,N_29116,N_28105);
nand U31297 (N_31297,N_29182,N_28901);
nand U31298 (N_31298,N_28799,N_28888);
xor U31299 (N_31299,N_29999,N_29075);
nor U31300 (N_31300,N_28805,N_29388);
nor U31301 (N_31301,N_28881,N_29696);
nand U31302 (N_31302,N_28561,N_28979);
xnor U31303 (N_31303,N_27830,N_28127);
nand U31304 (N_31304,N_29046,N_29132);
nor U31305 (N_31305,N_29720,N_28471);
nand U31306 (N_31306,N_27879,N_29698);
xor U31307 (N_31307,N_27668,N_29059);
and U31308 (N_31308,N_28209,N_29851);
xor U31309 (N_31309,N_29499,N_28648);
nor U31310 (N_31310,N_27740,N_28208);
or U31311 (N_31311,N_28704,N_29224);
xor U31312 (N_31312,N_29756,N_29980);
nor U31313 (N_31313,N_28481,N_28758);
xnor U31314 (N_31314,N_28150,N_28464);
or U31315 (N_31315,N_27920,N_28482);
or U31316 (N_31316,N_28758,N_28454);
and U31317 (N_31317,N_27687,N_29768);
nor U31318 (N_31318,N_29650,N_28517);
xnor U31319 (N_31319,N_28012,N_27547);
or U31320 (N_31320,N_28431,N_29256);
and U31321 (N_31321,N_27615,N_27632);
xnor U31322 (N_31322,N_29875,N_27606);
nand U31323 (N_31323,N_29691,N_27538);
nand U31324 (N_31324,N_29316,N_27549);
nor U31325 (N_31325,N_29260,N_29448);
xnor U31326 (N_31326,N_29015,N_29567);
nand U31327 (N_31327,N_28573,N_28989);
nor U31328 (N_31328,N_29561,N_29197);
xnor U31329 (N_31329,N_29768,N_28035);
or U31330 (N_31330,N_29727,N_29990);
nor U31331 (N_31331,N_28678,N_29019);
nor U31332 (N_31332,N_29463,N_29867);
xor U31333 (N_31333,N_29896,N_27895);
and U31334 (N_31334,N_28209,N_28053);
nand U31335 (N_31335,N_28253,N_28195);
or U31336 (N_31336,N_28493,N_29415);
xnor U31337 (N_31337,N_29863,N_28414);
xnor U31338 (N_31338,N_27579,N_28588);
nand U31339 (N_31339,N_28678,N_29956);
nor U31340 (N_31340,N_29806,N_29983);
and U31341 (N_31341,N_29435,N_29883);
nand U31342 (N_31342,N_28475,N_29306);
and U31343 (N_31343,N_29354,N_29626);
and U31344 (N_31344,N_29868,N_29390);
and U31345 (N_31345,N_27941,N_29558);
or U31346 (N_31346,N_28049,N_29497);
or U31347 (N_31347,N_29587,N_28956);
xor U31348 (N_31348,N_27960,N_28571);
and U31349 (N_31349,N_29593,N_28721);
nand U31350 (N_31350,N_29071,N_29224);
or U31351 (N_31351,N_27895,N_27666);
or U31352 (N_31352,N_28542,N_28603);
and U31353 (N_31353,N_29564,N_28951);
nor U31354 (N_31354,N_29618,N_29348);
nand U31355 (N_31355,N_29578,N_28280);
xor U31356 (N_31356,N_27850,N_28380);
nand U31357 (N_31357,N_28264,N_29582);
and U31358 (N_31358,N_29316,N_27522);
xor U31359 (N_31359,N_28326,N_29173);
nand U31360 (N_31360,N_28235,N_27599);
xnor U31361 (N_31361,N_28191,N_29009);
and U31362 (N_31362,N_29310,N_28431);
and U31363 (N_31363,N_29166,N_28535);
xnor U31364 (N_31364,N_28226,N_28690);
xnor U31365 (N_31365,N_29530,N_28107);
or U31366 (N_31366,N_27836,N_28444);
and U31367 (N_31367,N_29944,N_28663);
or U31368 (N_31368,N_29554,N_28397);
nand U31369 (N_31369,N_29131,N_27647);
and U31370 (N_31370,N_29419,N_29051);
nand U31371 (N_31371,N_28065,N_28855);
nor U31372 (N_31372,N_28431,N_29903);
nand U31373 (N_31373,N_29828,N_29565);
or U31374 (N_31374,N_29984,N_28878);
nor U31375 (N_31375,N_28637,N_29068);
nor U31376 (N_31376,N_29735,N_28156);
nand U31377 (N_31377,N_29012,N_28605);
xnor U31378 (N_31378,N_27808,N_29826);
and U31379 (N_31379,N_28428,N_27850);
or U31380 (N_31380,N_27801,N_28349);
or U31381 (N_31381,N_28803,N_28925);
and U31382 (N_31382,N_27954,N_28918);
and U31383 (N_31383,N_28857,N_27705);
or U31384 (N_31384,N_27576,N_28404);
xnor U31385 (N_31385,N_28189,N_29010);
xor U31386 (N_31386,N_27694,N_28452);
and U31387 (N_31387,N_28841,N_27986);
nor U31388 (N_31388,N_28703,N_27696);
nor U31389 (N_31389,N_27766,N_27885);
xor U31390 (N_31390,N_27714,N_29045);
or U31391 (N_31391,N_29503,N_28208);
or U31392 (N_31392,N_29569,N_29344);
nand U31393 (N_31393,N_28750,N_29183);
or U31394 (N_31394,N_29207,N_28751);
nor U31395 (N_31395,N_29101,N_29926);
nand U31396 (N_31396,N_27677,N_27502);
xnor U31397 (N_31397,N_29210,N_28906);
or U31398 (N_31398,N_28378,N_28384);
nand U31399 (N_31399,N_29721,N_29233);
nand U31400 (N_31400,N_28008,N_27713);
nor U31401 (N_31401,N_28636,N_29489);
or U31402 (N_31402,N_28500,N_28630);
or U31403 (N_31403,N_29597,N_28126);
nor U31404 (N_31404,N_29858,N_29981);
or U31405 (N_31405,N_29474,N_27863);
nor U31406 (N_31406,N_27754,N_29453);
and U31407 (N_31407,N_27975,N_29057);
nor U31408 (N_31408,N_27716,N_27667);
nand U31409 (N_31409,N_28565,N_29555);
xor U31410 (N_31410,N_28694,N_28001);
nand U31411 (N_31411,N_27761,N_29983);
nor U31412 (N_31412,N_29409,N_29423);
nand U31413 (N_31413,N_28087,N_29518);
and U31414 (N_31414,N_27577,N_27838);
nor U31415 (N_31415,N_27934,N_28507);
nor U31416 (N_31416,N_29394,N_28819);
nand U31417 (N_31417,N_28926,N_28887);
or U31418 (N_31418,N_28107,N_28326);
and U31419 (N_31419,N_29698,N_29395);
nand U31420 (N_31420,N_27966,N_28877);
nor U31421 (N_31421,N_27801,N_28307);
nand U31422 (N_31422,N_27726,N_29342);
and U31423 (N_31423,N_29500,N_28270);
and U31424 (N_31424,N_29960,N_28223);
nor U31425 (N_31425,N_27941,N_29422);
or U31426 (N_31426,N_27638,N_27907);
xor U31427 (N_31427,N_27921,N_29760);
nor U31428 (N_31428,N_29013,N_28574);
nor U31429 (N_31429,N_27549,N_27780);
and U31430 (N_31430,N_27561,N_29139);
and U31431 (N_31431,N_28837,N_28687);
or U31432 (N_31432,N_29033,N_27904);
xnor U31433 (N_31433,N_28854,N_28047);
nand U31434 (N_31434,N_29633,N_29689);
xor U31435 (N_31435,N_29294,N_27524);
or U31436 (N_31436,N_28794,N_27551);
and U31437 (N_31437,N_27860,N_27810);
nor U31438 (N_31438,N_29407,N_28748);
xor U31439 (N_31439,N_29362,N_27981);
nor U31440 (N_31440,N_28142,N_28596);
nand U31441 (N_31441,N_28660,N_28122);
nor U31442 (N_31442,N_28792,N_28456);
nand U31443 (N_31443,N_29239,N_29174);
and U31444 (N_31444,N_28978,N_27541);
nand U31445 (N_31445,N_29466,N_27910);
and U31446 (N_31446,N_28434,N_28022);
and U31447 (N_31447,N_28024,N_29954);
or U31448 (N_31448,N_29683,N_28648);
nor U31449 (N_31449,N_29136,N_28396);
and U31450 (N_31450,N_29994,N_28688);
nand U31451 (N_31451,N_29741,N_28611);
and U31452 (N_31452,N_28762,N_27616);
or U31453 (N_31453,N_29628,N_29466);
or U31454 (N_31454,N_29337,N_29539);
nor U31455 (N_31455,N_28415,N_29666);
nand U31456 (N_31456,N_29305,N_29916);
nand U31457 (N_31457,N_28688,N_27993);
or U31458 (N_31458,N_28342,N_28755);
or U31459 (N_31459,N_29857,N_28657);
xnor U31460 (N_31460,N_29413,N_27535);
or U31461 (N_31461,N_29065,N_28650);
nor U31462 (N_31462,N_29630,N_28382);
nand U31463 (N_31463,N_28491,N_28187);
nor U31464 (N_31464,N_28159,N_27603);
nor U31465 (N_31465,N_28316,N_29251);
or U31466 (N_31466,N_28520,N_29499);
nor U31467 (N_31467,N_28068,N_29823);
xor U31468 (N_31468,N_27565,N_29476);
nor U31469 (N_31469,N_28587,N_29819);
nand U31470 (N_31470,N_29401,N_28196);
or U31471 (N_31471,N_28133,N_27653);
nand U31472 (N_31472,N_27614,N_27664);
xor U31473 (N_31473,N_29497,N_29320);
or U31474 (N_31474,N_28077,N_28059);
or U31475 (N_31475,N_28396,N_29190);
xnor U31476 (N_31476,N_29942,N_28584);
nand U31477 (N_31477,N_28569,N_27985);
or U31478 (N_31478,N_28425,N_27931);
and U31479 (N_31479,N_28243,N_28442);
or U31480 (N_31480,N_27743,N_29155);
or U31481 (N_31481,N_28815,N_27961);
nor U31482 (N_31482,N_27727,N_27901);
nand U31483 (N_31483,N_28906,N_28387);
nand U31484 (N_31484,N_28387,N_29620);
nor U31485 (N_31485,N_28894,N_29864);
nor U31486 (N_31486,N_27575,N_27586);
nor U31487 (N_31487,N_28459,N_28645);
nand U31488 (N_31488,N_28063,N_28087);
nor U31489 (N_31489,N_27538,N_29635);
nor U31490 (N_31490,N_27700,N_28335);
nand U31491 (N_31491,N_29935,N_29160);
xor U31492 (N_31492,N_29999,N_29083);
or U31493 (N_31493,N_28500,N_28316);
and U31494 (N_31494,N_28105,N_27772);
and U31495 (N_31495,N_27888,N_29668);
nand U31496 (N_31496,N_27590,N_29616);
nand U31497 (N_31497,N_28192,N_29955);
nand U31498 (N_31498,N_29519,N_29648);
and U31499 (N_31499,N_29520,N_28342);
nand U31500 (N_31500,N_28568,N_27673);
nand U31501 (N_31501,N_28337,N_28357);
and U31502 (N_31502,N_28796,N_28748);
nand U31503 (N_31503,N_28332,N_29185);
xnor U31504 (N_31504,N_28268,N_27556);
and U31505 (N_31505,N_27673,N_28563);
xnor U31506 (N_31506,N_27806,N_28780);
xnor U31507 (N_31507,N_28199,N_27717);
or U31508 (N_31508,N_27615,N_29669);
nor U31509 (N_31509,N_28718,N_28631);
nor U31510 (N_31510,N_27794,N_27995);
and U31511 (N_31511,N_29688,N_29392);
or U31512 (N_31512,N_27607,N_28647);
nor U31513 (N_31513,N_27536,N_28177);
xor U31514 (N_31514,N_29652,N_29249);
and U31515 (N_31515,N_28523,N_28579);
nor U31516 (N_31516,N_29388,N_28868);
xnor U31517 (N_31517,N_29595,N_27915);
nor U31518 (N_31518,N_29655,N_27925);
xnor U31519 (N_31519,N_29047,N_28796);
nor U31520 (N_31520,N_27728,N_27579);
xnor U31521 (N_31521,N_27591,N_28886);
nand U31522 (N_31522,N_29117,N_28757);
nand U31523 (N_31523,N_28477,N_28696);
and U31524 (N_31524,N_27787,N_29029);
nor U31525 (N_31525,N_29573,N_27665);
and U31526 (N_31526,N_28233,N_29406);
or U31527 (N_31527,N_29607,N_29705);
and U31528 (N_31528,N_29200,N_27803);
or U31529 (N_31529,N_28210,N_28714);
and U31530 (N_31530,N_27969,N_27954);
nand U31531 (N_31531,N_29477,N_29938);
and U31532 (N_31532,N_28919,N_28739);
nand U31533 (N_31533,N_28237,N_29306);
xor U31534 (N_31534,N_28776,N_29099);
xnor U31535 (N_31535,N_28366,N_28837);
or U31536 (N_31536,N_28670,N_29175);
or U31537 (N_31537,N_29318,N_29234);
nand U31538 (N_31538,N_28855,N_29318);
and U31539 (N_31539,N_27790,N_27757);
and U31540 (N_31540,N_29713,N_29720);
nor U31541 (N_31541,N_29589,N_28279);
or U31542 (N_31542,N_27820,N_29228);
and U31543 (N_31543,N_27959,N_29405);
and U31544 (N_31544,N_28759,N_29688);
nand U31545 (N_31545,N_28854,N_27610);
and U31546 (N_31546,N_28436,N_29882);
nand U31547 (N_31547,N_29592,N_28316);
xnor U31548 (N_31548,N_28771,N_29240);
xor U31549 (N_31549,N_29837,N_28995);
xor U31550 (N_31550,N_27610,N_28635);
nand U31551 (N_31551,N_28273,N_29905);
nor U31552 (N_31552,N_27872,N_27667);
xor U31553 (N_31553,N_29333,N_27745);
nor U31554 (N_31554,N_29752,N_27601);
nand U31555 (N_31555,N_27961,N_28359);
xor U31556 (N_31556,N_29550,N_29776);
nor U31557 (N_31557,N_29562,N_28873);
and U31558 (N_31558,N_27586,N_29669);
and U31559 (N_31559,N_29525,N_29235);
xnor U31560 (N_31560,N_28308,N_27973);
nor U31561 (N_31561,N_28982,N_29393);
or U31562 (N_31562,N_27799,N_29802);
nand U31563 (N_31563,N_27965,N_27559);
nand U31564 (N_31564,N_29139,N_29722);
or U31565 (N_31565,N_28495,N_28664);
and U31566 (N_31566,N_29499,N_29097);
nor U31567 (N_31567,N_29642,N_28545);
and U31568 (N_31568,N_28334,N_29337);
xnor U31569 (N_31569,N_28304,N_27798);
nor U31570 (N_31570,N_29492,N_29903);
or U31571 (N_31571,N_28022,N_29281);
nor U31572 (N_31572,N_29911,N_29813);
or U31573 (N_31573,N_28294,N_28039);
or U31574 (N_31574,N_28536,N_29249);
nor U31575 (N_31575,N_29878,N_28711);
xor U31576 (N_31576,N_27729,N_27683);
or U31577 (N_31577,N_29821,N_28899);
or U31578 (N_31578,N_28985,N_29438);
xor U31579 (N_31579,N_28881,N_28985);
and U31580 (N_31580,N_29186,N_29945);
nand U31581 (N_31581,N_29042,N_28442);
and U31582 (N_31582,N_29974,N_28343);
nand U31583 (N_31583,N_28302,N_29106);
or U31584 (N_31584,N_28119,N_28315);
xnor U31585 (N_31585,N_27814,N_29277);
or U31586 (N_31586,N_29852,N_27746);
nand U31587 (N_31587,N_27592,N_28783);
xnor U31588 (N_31588,N_28236,N_29134);
and U31589 (N_31589,N_28278,N_28726);
and U31590 (N_31590,N_27918,N_28906);
nor U31591 (N_31591,N_28594,N_29977);
and U31592 (N_31592,N_29153,N_28050);
nor U31593 (N_31593,N_29210,N_29949);
xnor U31594 (N_31594,N_28124,N_29149);
and U31595 (N_31595,N_28302,N_28254);
nand U31596 (N_31596,N_27989,N_29806);
xor U31597 (N_31597,N_28259,N_29505);
xor U31598 (N_31598,N_29860,N_28238);
and U31599 (N_31599,N_27844,N_29901);
nor U31600 (N_31600,N_28413,N_29068);
nor U31601 (N_31601,N_28362,N_28875);
nand U31602 (N_31602,N_29733,N_29530);
nand U31603 (N_31603,N_29061,N_28357);
nor U31604 (N_31604,N_29055,N_28713);
nor U31605 (N_31605,N_29897,N_28859);
or U31606 (N_31606,N_28594,N_28943);
or U31607 (N_31607,N_27910,N_29085);
xnor U31608 (N_31608,N_28017,N_27950);
nand U31609 (N_31609,N_28776,N_28268);
nand U31610 (N_31610,N_28536,N_28874);
nand U31611 (N_31611,N_28258,N_28552);
and U31612 (N_31612,N_29266,N_29865);
or U31613 (N_31613,N_29689,N_29806);
nand U31614 (N_31614,N_28756,N_29490);
xnor U31615 (N_31615,N_28922,N_29905);
nand U31616 (N_31616,N_27628,N_29444);
and U31617 (N_31617,N_27791,N_28113);
and U31618 (N_31618,N_28839,N_29661);
and U31619 (N_31619,N_28662,N_29776);
and U31620 (N_31620,N_27755,N_29166);
nand U31621 (N_31621,N_28993,N_29955);
or U31622 (N_31622,N_28471,N_28933);
xnor U31623 (N_31623,N_29657,N_28237);
and U31624 (N_31624,N_28971,N_27726);
or U31625 (N_31625,N_29795,N_28917);
xnor U31626 (N_31626,N_29900,N_28912);
or U31627 (N_31627,N_29998,N_28057);
nor U31628 (N_31628,N_27501,N_29250);
or U31629 (N_31629,N_28639,N_28663);
or U31630 (N_31630,N_28175,N_29311);
or U31631 (N_31631,N_28618,N_29514);
xor U31632 (N_31632,N_29386,N_29489);
nor U31633 (N_31633,N_29706,N_29162);
nor U31634 (N_31634,N_28698,N_28738);
and U31635 (N_31635,N_28674,N_29179);
and U31636 (N_31636,N_27558,N_29282);
nor U31637 (N_31637,N_28681,N_28087);
and U31638 (N_31638,N_28073,N_29733);
or U31639 (N_31639,N_28558,N_29528);
nor U31640 (N_31640,N_29456,N_28475);
xnor U31641 (N_31641,N_27823,N_27760);
or U31642 (N_31642,N_28307,N_27940);
nand U31643 (N_31643,N_29342,N_29765);
or U31644 (N_31644,N_28997,N_29683);
nand U31645 (N_31645,N_28804,N_29676);
and U31646 (N_31646,N_29311,N_27540);
or U31647 (N_31647,N_28954,N_29244);
nand U31648 (N_31648,N_29903,N_29527);
and U31649 (N_31649,N_28416,N_28640);
nand U31650 (N_31650,N_27784,N_28277);
nand U31651 (N_31651,N_29098,N_29007);
nand U31652 (N_31652,N_29367,N_28355);
nor U31653 (N_31653,N_29475,N_27912);
or U31654 (N_31654,N_28576,N_29678);
xor U31655 (N_31655,N_29118,N_29924);
and U31656 (N_31656,N_27604,N_28057);
nand U31657 (N_31657,N_27966,N_28334);
xnor U31658 (N_31658,N_29858,N_28924);
xor U31659 (N_31659,N_27513,N_29705);
nor U31660 (N_31660,N_29879,N_29434);
nand U31661 (N_31661,N_29673,N_29465);
nor U31662 (N_31662,N_27835,N_28184);
nand U31663 (N_31663,N_29617,N_28566);
xor U31664 (N_31664,N_28772,N_27718);
nand U31665 (N_31665,N_27957,N_29405);
xnor U31666 (N_31666,N_28911,N_28517);
xnor U31667 (N_31667,N_29375,N_29450);
and U31668 (N_31668,N_27598,N_29166);
nand U31669 (N_31669,N_29439,N_27551);
or U31670 (N_31670,N_27825,N_29044);
nand U31671 (N_31671,N_27922,N_29708);
nor U31672 (N_31672,N_28843,N_29847);
xnor U31673 (N_31673,N_28445,N_27637);
nand U31674 (N_31674,N_29390,N_28103);
or U31675 (N_31675,N_28441,N_29644);
or U31676 (N_31676,N_29380,N_27687);
or U31677 (N_31677,N_29632,N_29826);
nand U31678 (N_31678,N_27858,N_28684);
nor U31679 (N_31679,N_28852,N_28337);
nor U31680 (N_31680,N_29624,N_29069);
and U31681 (N_31681,N_29328,N_29969);
or U31682 (N_31682,N_27857,N_28244);
nor U31683 (N_31683,N_27928,N_28523);
nand U31684 (N_31684,N_29909,N_29379);
nor U31685 (N_31685,N_29841,N_28529);
or U31686 (N_31686,N_27681,N_29819);
xor U31687 (N_31687,N_29406,N_28796);
nor U31688 (N_31688,N_28837,N_27783);
xor U31689 (N_31689,N_27841,N_29391);
and U31690 (N_31690,N_29757,N_27541);
xor U31691 (N_31691,N_27946,N_27796);
or U31692 (N_31692,N_28416,N_28996);
xor U31693 (N_31693,N_28865,N_29324);
or U31694 (N_31694,N_29758,N_29851);
xor U31695 (N_31695,N_29010,N_29007);
and U31696 (N_31696,N_27693,N_28662);
xnor U31697 (N_31697,N_27568,N_28903);
and U31698 (N_31698,N_29039,N_27984);
nor U31699 (N_31699,N_29513,N_28042);
or U31700 (N_31700,N_28762,N_29963);
or U31701 (N_31701,N_29451,N_27774);
and U31702 (N_31702,N_29919,N_27617);
or U31703 (N_31703,N_28306,N_29528);
and U31704 (N_31704,N_28339,N_28038);
nand U31705 (N_31705,N_29988,N_27610);
xnor U31706 (N_31706,N_28215,N_27826);
and U31707 (N_31707,N_29454,N_29687);
nor U31708 (N_31708,N_28902,N_29482);
nor U31709 (N_31709,N_29203,N_28867);
xor U31710 (N_31710,N_28986,N_28891);
nor U31711 (N_31711,N_29942,N_28779);
nor U31712 (N_31712,N_29247,N_28356);
nand U31713 (N_31713,N_28038,N_28077);
xor U31714 (N_31714,N_28986,N_27707);
nor U31715 (N_31715,N_29812,N_28089);
and U31716 (N_31716,N_28065,N_27543);
nor U31717 (N_31717,N_29849,N_29434);
and U31718 (N_31718,N_27610,N_29509);
and U31719 (N_31719,N_28592,N_28736);
and U31720 (N_31720,N_29972,N_27968);
or U31721 (N_31721,N_29993,N_29606);
xnor U31722 (N_31722,N_29002,N_29352);
xor U31723 (N_31723,N_28600,N_28711);
and U31724 (N_31724,N_29970,N_29141);
nand U31725 (N_31725,N_29004,N_29019);
or U31726 (N_31726,N_29324,N_28898);
nand U31727 (N_31727,N_29462,N_28169);
or U31728 (N_31728,N_28066,N_29634);
or U31729 (N_31729,N_28290,N_28717);
xnor U31730 (N_31730,N_29355,N_27554);
or U31731 (N_31731,N_27951,N_28404);
or U31732 (N_31732,N_28597,N_27972);
xnor U31733 (N_31733,N_27519,N_28125);
xnor U31734 (N_31734,N_29068,N_29840);
nor U31735 (N_31735,N_29892,N_28591);
nand U31736 (N_31736,N_27758,N_29150);
or U31737 (N_31737,N_29825,N_28805);
xor U31738 (N_31738,N_29099,N_29216);
nand U31739 (N_31739,N_28727,N_28294);
or U31740 (N_31740,N_28986,N_29684);
nand U31741 (N_31741,N_28972,N_28721);
and U31742 (N_31742,N_27905,N_29704);
xnor U31743 (N_31743,N_29508,N_28642);
xor U31744 (N_31744,N_28843,N_27789);
nand U31745 (N_31745,N_29343,N_28155);
xnor U31746 (N_31746,N_29914,N_28531);
or U31747 (N_31747,N_27827,N_29869);
nand U31748 (N_31748,N_28718,N_28886);
nand U31749 (N_31749,N_29367,N_29900);
and U31750 (N_31750,N_28054,N_28791);
and U31751 (N_31751,N_29106,N_28440);
nor U31752 (N_31752,N_28017,N_28755);
nand U31753 (N_31753,N_29789,N_28421);
nor U31754 (N_31754,N_28143,N_28333);
xnor U31755 (N_31755,N_29083,N_27854);
xor U31756 (N_31756,N_27902,N_28011);
xor U31757 (N_31757,N_29279,N_28299);
or U31758 (N_31758,N_28573,N_28769);
or U31759 (N_31759,N_29056,N_29018);
nor U31760 (N_31760,N_29491,N_27826);
nand U31761 (N_31761,N_29385,N_29040);
or U31762 (N_31762,N_29701,N_29185);
nor U31763 (N_31763,N_29144,N_29277);
nor U31764 (N_31764,N_29984,N_29588);
xor U31765 (N_31765,N_29341,N_29306);
or U31766 (N_31766,N_28247,N_29366);
and U31767 (N_31767,N_29086,N_29870);
nor U31768 (N_31768,N_28368,N_29386);
and U31769 (N_31769,N_28544,N_29999);
and U31770 (N_31770,N_29305,N_29442);
nand U31771 (N_31771,N_28508,N_27830);
or U31772 (N_31772,N_27966,N_28792);
nor U31773 (N_31773,N_28572,N_29893);
nand U31774 (N_31774,N_28765,N_29889);
nor U31775 (N_31775,N_28214,N_27971);
nor U31776 (N_31776,N_29028,N_29521);
xor U31777 (N_31777,N_28306,N_27953);
nor U31778 (N_31778,N_27809,N_28530);
and U31779 (N_31779,N_28481,N_28411);
nor U31780 (N_31780,N_28811,N_29425);
xnor U31781 (N_31781,N_28014,N_29229);
nor U31782 (N_31782,N_29481,N_27691);
nand U31783 (N_31783,N_28367,N_28437);
nand U31784 (N_31784,N_29509,N_27702);
or U31785 (N_31785,N_28880,N_28229);
xor U31786 (N_31786,N_28240,N_27928);
and U31787 (N_31787,N_28487,N_28258);
nand U31788 (N_31788,N_27976,N_29190);
or U31789 (N_31789,N_29665,N_29591);
and U31790 (N_31790,N_28840,N_29775);
xor U31791 (N_31791,N_28546,N_29484);
or U31792 (N_31792,N_28296,N_28895);
nand U31793 (N_31793,N_27752,N_28424);
or U31794 (N_31794,N_28542,N_29712);
nor U31795 (N_31795,N_29396,N_28480);
nor U31796 (N_31796,N_29575,N_27666);
xor U31797 (N_31797,N_28573,N_28823);
and U31798 (N_31798,N_27898,N_29341);
nor U31799 (N_31799,N_29756,N_29736);
nand U31800 (N_31800,N_28952,N_29449);
xor U31801 (N_31801,N_29424,N_28396);
xor U31802 (N_31802,N_29835,N_29703);
nor U31803 (N_31803,N_28437,N_29703);
nor U31804 (N_31804,N_29158,N_28750);
nor U31805 (N_31805,N_28373,N_28425);
nor U31806 (N_31806,N_28190,N_29235);
xnor U31807 (N_31807,N_28565,N_29948);
xnor U31808 (N_31808,N_29909,N_27778);
and U31809 (N_31809,N_29764,N_28024);
nor U31810 (N_31810,N_27585,N_29097);
nand U31811 (N_31811,N_29175,N_29099);
nor U31812 (N_31812,N_29432,N_29817);
nand U31813 (N_31813,N_29925,N_28826);
and U31814 (N_31814,N_28818,N_28996);
nor U31815 (N_31815,N_29794,N_29741);
and U31816 (N_31816,N_29793,N_28083);
and U31817 (N_31817,N_29502,N_28183);
and U31818 (N_31818,N_28218,N_27915);
or U31819 (N_31819,N_28716,N_28778);
or U31820 (N_31820,N_29535,N_29850);
or U31821 (N_31821,N_27891,N_28396);
and U31822 (N_31822,N_27584,N_28251);
or U31823 (N_31823,N_28742,N_29381);
nand U31824 (N_31824,N_28106,N_29667);
or U31825 (N_31825,N_29545,N_28723);
nor U31826 (N_31826,N_27618,N_29331);
nand U31827 (N_31827,N_29639,N_28010);
nand U31828 (N_31828,N_29883,N_29903);
and U31829 (N_31829,N_29330,N_28818);
xor U31830 (N_31830,N_28097,N_27989);
nand U31831 (N_31831,N_29054,N_29084);
nor U31832 (N_31832,N_28436,N_29698);
or U31833 (N_31833,N_29308,N_29648);
nand U31834 (N_31834,N_29593,N_28846);
nor U31835 (N_31835,N_28043,N_29456);
nor U31836 (N_31836,N_27547,N_27649);
xnor U31837 (N_31837,N_29515,N_27726);
xnor U31838 (N_31838,N_29036,N_29631);
nor U31839 (N_31839,N_28030,N_27612);
nor U31840 (N_31840,N_28842,N_29566);
nand U31841 (N_31841,N_28790,N_28232);
or U31842 (N_31842,N_27639,N_29464);
or U31843 (N_31843,N_29555,N_28812);
or U31844 (N_31844,N_28117,N_29267);
and U31845 (N_31845,N_28191,N_29058);
and U31846 (N_31846,N_29847,N_28793);
or U31847 (N_31847,N_28390,N_27503);
nor U31848 (N_31848,N_29441,N_29666);
xnor U31849 (N_31849,N_28348,N_29988);
xor U31850 (N_31850,N_28255,N_29070);
xnor U31851 (N_31851,N_28235,N_27986);
nor U31852 (N_31852,N_28337,N_27666);
and U31853 (N_31853,N_27555,N_29437);
or U31854 (N_31854,N_27503,N_27619);
xor U31855 (N_31855,N_29291,N_29605);
or U31856 (N_31856,N_29299,N_27593);
or U31857 (N_31857,N_28788,N_29148);
and U31858 (N_31858,N_29136,N_28611);
or U31859 (N_31859,N_28758,N_29108);
and U31860 (N_31860,N_29444,N_27655);
nor U31861 (N_31861,N_28357,N_28022);
xnor U31862 (N_31862,N_29751,N_27710);
or U31863 (N_31863,N_29594,N_28832);
nor U31864 (N_31864,N_29314,N_29493);
nand U31865 (N_31865,N_27880,N_27810);
or U31866 (N_31866,N_27909,N_29967);
or U31867 (N_31867,N_29105,N_29556);
or U31868 (N_31868,N_27613,N_29952);
nor U31869 (N_31869,N_29914,N_27931);
or U31870 (N_31870,N_28076,N_28233);
nand U31871 (N_31871,N_29350,N_29141);
xor U31872 (N_31872,N_27933,N_29805);
nand U31873 (N_31873,N_28869,N_29350);
nand U31874 (N_31874,N_28547,N_29985);
or U31875 (N_31875,N_29673,N_29031);
nor U31876 (N_31876,N_28880,N_27778);
nand U31877 (N_31877,N_28902,N_28560);
or U31878 (N_31878,N_29738,N_28745);
xor U31879 (N_31879,N_29377,N_28489);
nand U31880 (N_31880,N_29938,N_28500);
xnor U31881 (N_31881,N_27792,N_28090);
and U31882 (N_31882,N_29290,N_28050);
nor U31883 (N_31883,N_28408,N_29965);
nand U31884 (N_31884,N_28820,N_29339);
and U31885 (N_31885,N_29217,N_29275);
xor U31886 (N_31886,N_29902,N_29009);
or U31887 (N_31887,N_29277,N_28642);
and U31888 (N_31888,N_28736,N_29274);
or U31889 (N_31889,N_27678,N_28022);
xnor U31890 (N_31890,N_28071,N_29870);
and U31891 (N_31891,N_29908,N_29707);
xor U31892 (N_31892,N_28918,N_29350);
and U31893 (N_31893,N_28712,N_29281);
or U31894 (N_31894,N_27985,N_28201);
and U31895 (N_31895,N_28913,N_29031);
and U31896 (N_31896,N_29187,N_29244);
nand U31897 (N_31897,N_27512,N_29206);
nor U31898 (N_31898,N_29327,N_28565);
and U31899 (N_31899,N_29134,N_29505);
nand U31900 (N_31900,N_27563,N_28241);
nand U31901 (N_31901,N_29017,N_29659);
and U31902 (N_31902,N_27792,N_27587);
or U31903 (N_31903,N_29284,N_28907);
nor U31904 (N_31904,N_29622,N_28888);
and U31905 (N_31905,N_28598,N_28323);
nand U31906 (N_31906,N_28433,N_28257);
nand U31907 (N_31907,N_28403,N_29949);
nand U31908 (N_31908,N_29716,N_29566);
and U31909 (N_31909,N_28442,N_29711);
or U31910 (N_31910,N_29156,N_27554);
nor U31911 (N_31911,N_28069,N_28705);
xor U31912 (N_31912,N_27591,N_28897);
or U31913 (N_31913,N_28117,N_28548);
and U31914 (N_31914,N_28492,N_28369);
nand U31915 (N_31915,N_29618,N_29078);
or U31916 (N_31916,N_27807,N_28180);
and U31917 (N_31917,N_29252,N_29219);
or U31918 (N_31918,N_29892,N_28357);
or U31919 (N_31919,N_29905,N_27793);
and U31920 (N_31920,N_28437,N_29071);
nor U31921 (N_31921,N_29313,N_29644);
nor U31922 (N_31922,N_27532,N_29269);
or U31923 (N_31923,N_29488,N_28970);
or U31924 (N_31924,N_27777,N_27709);
xnor U31925 (N_31925,N_29765,N_29064);
or U31926 (N_31926,N_28218,N_28524);
and U31927 (N_31927,N_27710,N_27762);
or U31928 (N_31928,N_29887,N_29749);
nand U31929 (N_31929,N_28568,N_28581);
nor U31930 (N_31930,N_29545,N_29115);
or U31931 (N_31931,N_29604,N_29040);
or U31932 (N_31932,N_27592,N_29341);
xor U31933 (N_31933,N_27599,N_28127);
nor U31934 (N_31934,N_27501,N_28785);
and U31935 (N_31935,N_29049,N_28094);
xnor U31936 (N_31936,N_29265,N_29139);
or U31937 (N_31937,N_29817,N_27544);
xor U31938 (N_31938,N_29905,N_29785);
and U31939 (N_31939,N_27633,N_28067);
or U31940 (N_31940,N_29708,N_28935);
nor U31941 (N_31941,N_29332,N_28102);
nand U31942 (N_31942,N_29279,N_27576);
nor U31943 (N_31943,N_29833,N_27951);
nand U31944 (N_31944,N_28569,N_29069);
xnor U31945 (N_31945,N_29128,N_27970);
or U31946 (N_31946,N_29521,N_28953);
and U31947 (N_31947,N_29584,N_28582);
nand U31948 (N_31948,N_28627,N_28673);
or U31949 (N_31949,N_28638,N_29885);
nor U31950 (N_31950,N_28110,N_28836);
nand U31951 (N_31951,N_28948,N_28522);
or U31952 (N_31952,N_27778,N_28583);
xor U31953 (N_31953,N_29593,N_29885);
nor U31954 (N_31954,N_28375,N_28088);
xnor U31955 (N_31955,N_29922,N_27871);
nor U31956 (N_31956,N_28493,N_28834);
nor U31957 (N_31957,N_29678,N_28345);
xor U31958 (N_31958,N_27814,N_28980);
nand U31959 (N_31959,N_29737,N_27992);
and U31960 (N_31960,N_28564,N_29675);
nor U31961 (N_31961,N_28362,N_29438);
xnor U31962 (N_31962,N_28716,N_28791);
xor U31963 (N_31963,N_29223,N_27920);
nor U31964 (N_31964,N_27865,N_27803);
xor U31965 (N_31965,N_29654,N_29839);
or U31966 (N_31966,N_27869,N_29322);
or U31967 (N_31967,N_28634,N_29244);
xnor U31968 (N_31968,N_27567,N_28696);
and U31969 (N_31969,N_28465,N_29669);
nand U31970 (N_31970,N_28470,N_29806);
xor U31971 (N_31971,N_29670,N_28607);
nor U31972 (N_31972,N_29420,N_29259);
and U31973 (N_31973,N_29390,N_29806);
nor U31974 (N_31974,N_28280,N_27810);
xor U31975 (N_31975,N_29058,N_27549);
and U31976 (N_31976,N_27832,N_28909);
or U31977 (N_31977,N_29427,N_27753);
or U31978 (N_31978,N_29927,N_29782);
nor U31979 (N_31979,N_29229,N_29208);
nor U31980 (N_31980,N_28486,N_27912);
nand U31981 (N_31981,N_28285,N_29193);
nand U31982 (N_31982,N_28616,N_29063);
nor U31983 (N_31983,N_29165,N_29577);
xor U31984 (N_31984,N_29455,N_27901);
or U31985 (N_31985,N_29506,N_28548);
xor U31986 (N_31986,N_28254,N_28586);
nor U31987 (N_31987,N_27846,N_29818);
xnor U31988 (N_31988,N_29143,N_29470);
nand U31989 (N_31989,N_28876,N_29769);
nor U31990 (N_31990,N_28105,N_29921);
xnor U31991 (N_31991,N_28804,N_29209);
nor U31992 (N_31992,N_27550,N_27577);
nand U31993 (N_31993,N_27538,N_28372);
or U31994 (N_31994,N_29182,N_29566);
or U31995 (N_31995,N_27535,N_27531);
and U31996 (N_31996,N_28356,N_28250);
and U31997 (N_31997,N_29364,N_29143);
nor U31998 (N_31998,N_28595,N_29666);
nand U31999 (N_31999,N_29805,N_29849);
xor U32000 (N_32000,N_29082,N_29293);
nor U32001 (N_32001,N_29817,N_27599);
nor U32002 (N_32002,N_29336,N_28002);
and U32003 (N_32003,N_27600,N_27967);
nand U32004 (N_32004,N_27955,N_28657);
xnor U32005 (N_32005,N_28383,N_27803);
nand U32006 (N_32006,N_29665,N_28268);
or U32007 (N_32007,N_28637,N_28351);
or U32008 (N_32008,N_28811,N_28380);
xnor U32009 (N_32009,N_28198,N_27607);
xor U32010 (N_32010,N_27667,N_29614);
and U32011 (N_32011,N_28507,N_27660);
nand U32012 (N_32012,N_28743,N_29337);
nand U32013 (N_32013,N_29572,N_28178);
or U32014 (N_32014,N_28522,N_29902);
nand U32015 (N_32015,N_27744,N_28434);
nand U32016 (N_32016,N_28768,N_29604);
xnor U32017 (N_32017,N_27900,N_28791);
or U32018 (N_32018,N_27728,N_27993);
or U32019 (N_32019,N_29916,N_29534);
nor U32020 (N_32020,N_28027,N_28261);
or U32021 (N_32021,N_27738,N_29682);
xnor U32022 (N_32022,N_29702,N_29045);
xor U32023 (N_32023,N_29898,N_29408);
nor U32024 (N_32024,N_28465,N_28986);
and U32025 (N_32025,N_28748,N_29308);
nor U32026 (N_32026,N_29026,N_27878);
xor U32027 (N_32027,N_27793,N_28910);
nand U32028 (N_32028,N_29365,N_29395);
nor U32029 (N_32029,N_28213,N_28184);
nor U32030 (N_32030,N_29597,N_28612);
nand U32031 (N_32031,N_29411,N_28475);
or U32032 (N_32032,N_29763,N_29515);
or U32033 (N_32033,N_28262,N_27962);
nand U32034 (N_32034,N_29984,N_29215);
or U32035 (N_32035,N_29666,N_28032);
and U32036 (N_32036,N_29936,N_29250);
or U32037 (N_32037,N_28548,N_29154);
xnor U32038 (N_32038,N_27971,N_27720);
nor U32039 (N_32039,N_27845,N_29925);
and U32040 (N_32040,N_27988,N_27686);
nand U32041 (N_32041,N_27869,N_28673);
xnor U32042 (N_32042,N_27616,N_29919);
xor U32043 (N_32043,N_29845,N_28193);
xnor U32044 (N_32044,N_29933,N_28120);
xnor U32045 (N_32045,N_28212,N_27862);
or U32046 (N_32046,N_28117,N_28632);
nor U32047 (N_32047,N_29381,N_29434);
xor U32048 (N_32048,N_29497,N_28053);
and U32049 (N_32049,N_27501,N_29469);
nor U32050 (N_32050,N_29506,N_28596);
nor U32051 (N_32051,N_29977,N_28182);
nor U32052 (N_32052,N_27571,N_29860);
xnor U32053 (N_32053,N_29058,N_29037);
or U32054 (N_32054,N_29612,N_28267);
or U32055 (N_32055,N_28890,N_29955);
xnor U32056 (N_32056,N_29071,N_29411);
nor U32057 (N_32057,N_29247,N_29520);
and U32058 (N_32058,N_27870,N_29926);
nor U32059 (N_32059,N_29153,N_29658);
and U32060 (N_32060,N_29359,N_29318);
nand U32061 (N_32061,N_29002,N_28777);
or U32062 (N_32062,N_29234,N_28392);
nor U32063 (N_32063,N_28627,N_28009);
nor U32064 (N_32064,N_28332,N_29703);
nand U32065 (N_32065,N_27750,N_28799);
nor U32066 (N_32066,N_29958,N_28223);
and U32067 (N_32067,N_29305,N_29669);
nand U32068 (N_32068,N_27588,N_28995);
nand U32069 (N_32069,N_28890,N_28441);
and U32070 (N_32070,N_27660,N_29975);
xor U32071 (N_32071,N_29839,N_28919);
xor U32072 (N_32072,N_29290,N_27675);
nor U32073 (N_32073,N_29031,N_29888);
nor U32074 (N_32074,N_28711,N_29624);
xnor U32075 (N_32075,N_29975,N_29465);
xnor U32076 (N_32076,N_29068,N_28053);
nand U32077 (N_32077,N_29080,N_29434);
nand U32078 (N_32078,N_28537,N_28155);
xnor U32079 (N_32079,N_29115,N_29925);
nor U32080 (N_32080,N_27932,N_29843);
and U32081 (N_32081,N_27881,N_29550);
nor U32082 (N_32082,N_29761,N_28556);
or U32083 (N_32083,N_28968,N_29661);
nand U32084 (N_32084,N_28450,N_28584);
nor U32085 (N_32085,N_29716,N_28077);
xor U32086 (N_32086,N_29170,N_27960);
xnor U32087 (N_32087,N_28437,N_28935);
nand U32088 (N_32088,N_28943,N_29146);
xnor U32089 (N_32089,N_29868,N_28085);
or U32090 (N_32090,N_29076,N_28656);
and U32091 (N_32091,N_29012,N_29914);
nand U32092 (N_32092,N_28350,N_28432);
or U32093 (N_32093,N_28087,N_28077);
nor U32094 (N_32094,N_27744,N_28121);
xnor U32095 (N_32095,N_29179,N_28946);
nand U32096 (N_32096,N_28004,N_29712);
and U32097 (N_32097,N_28775,N_29909);
nand U32098 (N_32098,N_28918,N_27618);
nor U32099 (N_32099,N_29160,N_28263);
and U32100 (N_32100,N_29276,N_29794);
nor U32101 (N_32101,N_28349,N_29657);
nor U32102 (N_32102,N_28300,N_28006);
xor U32103 (N_32103,N_27822,N_28846);
nor U32104 (N_32104,N_27714,N_29844);
nand U32105 (N_32105,N_28864,N_29192);
xor U32106 (N_32106,N_28219,N_28279);
xnor U32107 (N_32107,N_29675,N_29742);
nor U32108 (N_32108,N_29831,N_27742);
xor U32109 (N_32109,N_28456,N_29424);
and U32110 (N_32110,N_29184,N_27550);
nand U32111 (N_32111,N_29976,N_29205);
xor U32112 (N_32112,N_28256,N_29686);
or U32113 (N_32113,N_29309,N_28029);
nor U32114 (N_32114,N_28229,N_28342);
xnor U32115 (N_32115,N_29379,N_27831);
nor U32116 (N_32116,N_28753,N_27578);
nand U32117 (N_32117,N_28284,N_28188);
and U32118 (N_32118,N_27513,N_29917);
or U32119 (N_32119,N_28364,N_28837);
nand U32120 (N_32120,N_29730,N_29724);
xor U32121 (N_32121,N_27961,N_27805);
nand U32122 (N_32122,N_28085,N_27968);
nand U32123 (N_32123,N_29591,N_29647);
nand U32124 (N_32124,N_28574,N_29646);
nor U32125 (N_32125,N_29743,N_28162);
nand U32126 (N_32126,N_27629,N_28879);
and U32127 (N_32127,N_28832,N_28984);
xnor U32128 (N_32128,N_28350,N_27747);
nand U32129 (N_32129,N_29263,N_28457);
nor U32130 (N_32130,N_29331,N_29849);
xnor U32131 (N_32131,N_29389,N_27666);
and U32132 (N_32132,N_28095,N_29935);
nand U32133 (N_32133,N_27748,N_29775);
nand U32134 (N_32134,N_29636,N_29708);
xnor U32135 (N_32135,N_29508,N_27864);
nand U32136 (N_32136,N_29558,N_28809);
nor U32137 (N_32137,N_29666,N_28071);
nand U32138 (N_32138,N_29573,N_29081);
nand U32139 (N_32139,N_29817,N_28583);
nor U32140 (N_32140,N_27562,N_27596);
nand U32141 (N_32141,N_28372,N_28589);
nand U32142 (N_32142,N_28514,N_28049);
nor U32143 (N_32143,N_28153,N_29332);
and U32144 (N_32144,N_28080,N_28889);
xnor U32145 (N_32145,N_29499,N_29703);
xnor U32146 (N_32146,N_29892,N_28300);
nor U32147 (N_32147,N_27950,N_29867);
nor U32148 (N_32148,N_28690,N_27818);
nand U32149 (N_32149,N_28170,N_28326);
xor U32150 (N_32150,N_29718,N_28089);
xor U32151 (N_32151,N_28628,N_28676);
nand U32152 (N_32152,N_28418,N_29485);
nand U32153 (N_32153,N_28131,N_29338);
or U32154 (N_32154,N_28327,N_28134);
nand U32155 (N_32155,N_29635,N_28861);
nor U32156 (N_32156,N_28504,N_28074);
nand U32157 (N_32157,N_28082,N_29153);
or U32158 (N_32158,N_27899,N_28852);
xor U32159 (N_32159,N_28873,N_28362);
or U32160 (N_32160,N_29522,N_29736);
and U32161 (N_32161,N_27901,N_29299);
and U32162 (N_32162,N_28908,N_28145);
nand U32163 (N_32163,N_29518,N_27602);
xor U32164 (N_32164,N_28368,N_27690);
nor U32165 (N_32165,N_28728,N_28447);
nor U32166 (N_32166,N_29791,N_29726);
nand U32167 (N_32167,N_27834,N_29824);
or U32168 (N_32168,N_29765,N_29486);
xor U32169 (N_32169,N_28816,N_28389);
nor U32170 (N_32170,N_28118,N_28939);
and U32171 (N_32171,N_27512,N_29394);
and U32172 (N_32172,N_29655,N_28499);
nor U32173 (N_32173,N_28371,N_28253);
or U32174 (N_32174,N_28272,N_29402);
nor U32175 (N_32175,N_27689,N_28973);
or U32176 (N_32176,N_27568,N_29402);
and U32177 (N_32177,N_27707,N_29283);
nor U32178 (N_32178,N_29575,N_27894);
or U32179 (N_32179,N_29769,N_27848);
nor U32180 (N_32180,N_29085,N_28469);
or U32181 (N_32181,N_29204,N_28437);
or U32182 (N_32182,N_29638,N_27947);
nor U32183 (N_32183,N_27536,N_29660);
nor U32184 (N_32184,N_27710,N_27989);
nand U32185 (N_32185,N_27983,N_27898);
nand U32186 (N_32186,N_27738,N_27920);
xor U32187 (N_32187,N_27639,N_29827);
xor U32188 (N_32188,N_29783,N_29736);
and U32189 (N_32189,N_27582,N_28064);
xor U32190 (N_32190,N_29934,N_29036);
and U32191 (N_32191,N_28434,N_29675);
xor U32192 (N_32192,N_29451,N_28659);
xnor U32193 (N_32193,N_27954,N_28999);
and U32194 (N_32194,N_28600,N_27580);
or U32195 (N_32195,N_29199,N_28173);
and U32196 (N_32196,N_27978,N_29890);
nor U32197 (N_32197,N_29348,N_29778);
and U32198 (N_32198,N_27730,N_28386);
or U32199 (N_32199,N_28573,N_29436);
and U32200 (N_32200,N_27927,N_29696);
nor U32201 (N_32201,N_29776,N_27653);
and U32202 (N_32202,N_28106,N_28112);
and U32203 (N_32203,N_28270,N_27953);
xor U32204 (N_32204,N_28809,N_28198);
and U32205 (N_32205,N_28026,N_29243);
nand U32206 (N_32206,N_28483,N_29453);
nand U32207 (N_32207,N_27661,N_28135);
nand U32208 (N_32208,N_28317,N_28385);
or U32209 (N_32209,N_28618,N_28122);
xnor U32210 (N_32210,N_29004,N_29712);
nor U32211 (N_32211,N_28282,N_28036);
nor U32212 (N_32212,N_28448,N_29340);
and U32213 (N_32213,N_29379,N_29589);
or U32214 (N_32214,N_29547,N_29178);
and U32215 (N_32215,N_27525,N_29818);
xnor U32216 (N_32216,N_29612,N_28437);
or U32217 (N_32217,N_29923,N_27514);
or U32218 (N_32218,N_29736,N_29578);
xnor U32219 (N_32219,N_27802,N_28271);
xnor U32220 (N_32220,N_28552,N_28301);
nor U32221 (N_32221,N_28403,N_28183);
nand U32222 (N_32222,N_27770,N_27859);
and U32223 (N_32223,N_29330,N_29172);
nor U32224 (N_32224,N_28419,N_28551);
or U32225 (N_32225,N_29812,N_27945);
nor U32226 (N_32226,N_27934,N_27877);
or U32227 (N_32227,N_29687,N_28351);
nor U32228 (N_32228,N_28931,N_28776);
nor U32229 (N_32229,N_27825,N_29509);
nand U32230 (N_32230,N_28664,N_29981);
xnor U32231 (N_32231,N_29053,N_28979);
nand U32232 (N_32232,N_28913,N_28852);
and U32233 (N_32233,N_29249,N_29437);
nand U32234 (N_32234,N_29810,N_29499);
and U32235 (N_32235,N_28700,N_27674);
xor U32236 (N_32236,N_29828,N_28628);
xnor U32237 (N_32237,N_29262,N_29738);
and U32238 (N_32238,N_28854,N_27700);
nand U32239 (N_32239,N_27742,N_28161);
or U32240 (N_32240,N_29877,N_28903);
xnor U32241 (N_32241,N_29350,N_28417);
nand U32242 (N_32242,N_28671,N_28905);
nand U32243 (N_32243,N_27718,N_28277);
nor U32244 (N_32244,N_28091,N_29847);
nor U32245 (N_32245,N_28767,N_28277);
xor U32246 (N_32246,N_29346,N_29901);
nand U32247 (N_32247,N_27532,N_27728);
nor U32248 (N_32248,N_28022,N_28785);
nor U32249 (N_32249,N_29211,N_28352);
or U32250 (N_32250,N_28351,N_27697);
xor U32251 (N_32251,N_29898,N_29828);
and U32252 (N_32252,N_27950,N_28213);
xor U32253 (N_32253,N_29252,N_28720);
nand U32254 (N_32254,N_29423,N_29566);
xor U32255 (N_32255,N_29089,N_29963);
xnor U32256 (N_32256,N_29604,N_27695);
nor U32257 (N_32257,N_29077,N_27834);
or U32258 (N_32258,N_29224,N_29956);
or U32259 (N_32259,N_29395,N_28530);
xor U32260 (N_32260,N_28041,N_29817);
and U32261 (N_32261,N_28246,N_29579);
and U32262 (N_32262,N_28564,N_28428);
and U32263 (N_32263,N_28508,N_27700);
xor U32264 (N_32264,N_28359,N_29543);
nor U32265 (N_32265,N_28281,N_28656);
or U32266 (N_32266,N_27908,N_28576);
or U32267 (N_32267,N_29672,N_27930);
xor U32268 (N_32268,N_28375,N_28223);
nor U32269 (N_32269,N_28683,N_29452);
nor U32270 (N_32270,N_27795,N_28912);
nor U32271 (N_32271,N_28902,N_29172);
nor U32272 (N_32272,N_28874,N_27899);
nor U32273 (N_32273,N_28278,N_29009);
and U32274 (N_32274,N_27698,N_28251);
nor U32275 (N_32275,N_29615,N_28120);
xor U32276 (N_32276,N_28684,N_27811);
and U32277 (N_32277,N_27743,N_29870);
and U32278 (N_32278,N_29388,N_27787);
or U32279 (N_32279,N_28018,N_28844);
xnor U32280 (N_32280,N_28105,N_29088);
and U32281 (N_32281,N_27520,N_27833);
nand U32282 (N_32282,N_29291,N_28014);
or U32283 (N_32283,N_27892,N_29902);
nand U32284 (N_32284,N_27680,N_27581);
xnor U32285 (N_32285,N_28631,N_29901);
xnor U32286 (N_32286,N_28777,N_29409);
nand U32287 (N_32287,N_29791,N_28963);
nand U32288 (N_32288,N_27652,N_28753);
and U32289 (N_32289,N_28207,N_28563);
and U32290 (N_32290,N_29420,N_28571);
or U32291 (N_32291,N_27643,N_29052);
and U32292 (N_32292,N_29520,N_27903);
nand U32293 (N_32293,N_27860,N_28698);
nor U32294 (N_32294,N_27619,N_28774);
xor U32295 (N_32295,N_28965,N_28079);
or U32296 (N_32296,N_29951,N_27997);
xnor U32297 (N_32297,N_29767,N_29090);
nor U32298 (N_32298,N_29551,N_29505);
xor U32299 (N_32299,N_28443,N_27781);
nor U32300 (N_32300,N_28785,N_28224);
xnor U32301 (N_32301,N_28374,N_27868);
nor U32302 (N_32302,N_27826,N_27715);
nand U32303 (N_32303,N_29882,N_28541);
or U32304 (N_32304,N_27983,N_29713);
xnor U32305 (N_32305,N_28371,N_27796);
xor U32306 (N_32306,N_28385,N_28015);
xor U32307 (N_32307,N_29593,N_28446);
nand U32308 (N_32308,N_28952,N_29886);
nand U32309 (N_32309,N_29818,N_29903);
nand U32310 (N_32310,N_28003,N_27725);
xnor U32311 (N_32311,N_28768,N_28119);
and U32312 (N_32312,N_29332,N_28288);
nand U32313 (N_32313,N_28786,N_28069);
or U32314 (N_32314,N_28158,N_29705);
nand U32315 (N_32315,N_28870,N_28626);
or U32316 (N_32316,N_28821,N_29107);
or U32317 (N_32317,N_29471,N_27822);
nand U32318 (N_32318,N_29295,N_28030);
or U32319 (N_32319,N_28240,N_29742);
nand U32320 (N_32320,N_28687,N_28954);
nor U32321 (N_32321,N_28748,N_28396);
nor U32322 (N_32322,N_29946,N_28840);
nor U32323 (N_32323,N_29124,N_29059);
nor U32324 (N_32324,N_28483,N_29489);
xor U32325 (N_32325,N_28600,N_29099);
nor U32326 (N_32326,N_27578,N_28769);
nand U32327 (N_32327,N_28450,N_28371);
nand U32328 (N_32328,N_27835,N_29700);
xor U32329 (N_32329,N_28064,N_27890);
and U32330 (N_32330,N_28814,N_27842);
nand U32331 (N_32331,N_28801,N_29549);
and U32332 (N_32332,N_28934,N_29624);
and U32333 (N_32333,N_28546,N_28437);
nand U32334 (N_32334,N_28416,N_28890);
nor U32335 (N_32335,N_28480,N_29097);
nand U32336 (N_32336,N_29723,N_27872);
xnor U32337 (N_32337,N_29997,N_28762);
nand U32338 (N_32338,N_29936,N_28025);
and U32339 (N_32339,N_27550,N_28263);
and U32340 (N_32340,N_29625,N_29233);
nand U32341 (N_32341,N_29142,N_28108);
nor U32342 (N_32342,N_29097,N_29889);
and U32343 (N_32343,N_27692,N_27743);
or U32344 (N_32344,N_27696,N_29894);
or U32345 (N_32345,N_29408,N_28075);
xnor U32346 (N_32346,N_28997,N_29402);
nor U32347 (N_32347,N_29580,N_29773);
nand U32348 (N_32348,N_29840,N_29993);
xor U32349 (N_32349,N_29261,N_29376);
nand U32350 (N_32350,N_27665,N_28186);
or U32351 (N_32351,N_29358,N_29107);
xor U32352 (N_32352,N_28365,N_28288);
nand U32353 (N_32353,N_29101,N_29759);
nor U32354 (N_32354,N_28247,N_27743);
or U32355 (N_32355,N_29665,N_28324);
nand U32356 (N_32356,N_27898,N_29363);
nand U32357 (N_32357,N_28383,N_28447);
nand U32358 (N_32358,N_28947,N_29573);
nand U32359 (N_32359,N_27611,N_29186);
or U32360 (N_32360,N_29475,N_27968);
xor U32361 (N_32361,N_29483,N_27764);
nor U32362 (N_32362,N_29927,N_29479);
nor U32363 (N_32363,N_29469,N_29366);
nand U32364 (N_32364,N_28413,N_27743);
and U32365 (N_32365,N_29468,N_29422);
nand U32366 (N_32366,N_29521,N_28779);
or U32367 (N_32367,N_29609,N_27512);
nand U32368 (N_32368,N_27914,N_28509);
nand U32369 (N_32369,N_28195,N_28194);
nor U32370 (N_32370,N_28310,N_27897);
nand U32371 (N_32371,N_29963,N_29844);
and U32372 (N_32372,N_29559,N_29028);
nand U32373 (N_32373,N_28510,N_28398);
nand U32374 (N_32374,N_29252,N_29145);
xor U32375 (N_32375,N_27961,N_29651);
nor U32376 (N_32376,N_29958,N_28374);
nand U32377 (N_32377,N_28062,N_28040);
or U32378 (N_32378,N_29606,N_29538);
or U32379 (N_32379,N_29606,N_28624);
xnor U32380 (N_32380,N_29970,N_28689);
xor U32381 (N_32381,N_27936,N_28686);
nand U32382 (N_32382,N_29391,N_28686);
and U32383 (N_32383,N_28571,N_27658);
and U32384 (N_32384,N_29383,N_29310);
and U32385 (N_32385,N_28734,N_27689);
nor U32386 (N_32386,N_29639,N_28383);
xnor U32387 (N_32387,N_27797,N_29086);
and U32388 (N_32388,N_29686,N_27966);
xor U32389 (N_32389,N_29634,N_28388);
nor U32390 (N_32390,N_28303,N_28815);
nor U32391 (N_32391,N_27596,N_29988);
or U32392 (N_32392,N_29447,N_28717);
or U32393 (N_32393,N_28931,N_28820);
nand U32394 (N_32394,N_29316,N_29107);
nand U32395 (N_32395,N_29647,N_29981);
nand U32396 (N_32396,N_28572,N_29355);
or U32397 (N_32397,N_29526,N_28840);
nor U32398 (N_32398,N_27682,N_28567);
nor U32399 (N_32399,N_29434,N_28320);
and U32400 (N_32400,N_29554,N_28194);
nor U32401 (N_32401,N_29612,N_29643);
xor U32402 (N_32402,N_29561,N_28049);
nor U32403 (N_32403,N_28862,N_29774);
xor U32404 (N_32404,N_29201,N_27935);
xor U32405 (N_32405,N_27667,N_27668);
nand U32406 (N_32406,N_29551,N_28026);
nand U32407 (N_32407,N_29335,N_29567);
or U32408 (N_32408,N_28731,N_27638);
or U32409 (N_32409,N_28137,N_28633);
and U32410 (N_32410,N_29182,N_27678);
nor U32411 (N_32411,N_28363,N_29983);
nor U32412 (N_32412,N_29136,N_28051);
xnor U32413 (N_32413,N_28349,N_28739);
or U32414 (N_32414,N_29650,N_29919);
xnor U32415 (N_32415,N_28656,N_28684);
nor U32416 (N_32416,N_28042,N_29383);
nand U32417 (N_32417,N_27817,N_28639);
or U32418 (N_32418,N_29818,N_28928);
xor U32419 (N_32419,N_29161,N_28110);
nand U32420 (N_32420,N_29874,N_29204);
or U32421 (N_32421,N_28566,N_28312);
and U32422 (N_32422,N_27930,N_28397);
nand U32423 (N_32423,N_27984,N_29915);
or U32424 (N_32424,N_27957,N_28567);
or U32425 (N_32425,N_27943,N_28508);
and U32426 (N_32426,N_29471,N_28582);
and U32427 (N_32427,N_27593,N_28942);
nor U32428 (N_32428,N_29904,N_29970);
xnor U32429 (N_32429,N_29116,N_29230);
nand U32430 (N_32430,N_28018,N_29332);
and U32431 (N_32431,N_27917,N_28389);
nand U32432 (N_32432,N_29293,N_29026);
and U32433 (N_32433,N_27616,N_28958);
xnor U32434 (N_32434,N_28856,N_29744);
xor U32435 (N_32435,N_29557,N_27901);
xor U32436 (N_32436,N_27659,N_28621);
or U32437 (N_32437,N_28532,N_29033);
and U32438 (N_32438,N_29420,N_29112);
nor U32439 (N_32439,N_28089,N_29628);
and U32440 (N_32440,N_27506,N_28597);
and U32441 (N_32441,N_28155,N_28855);
or U32442 (N_32442,N_28863,N_29979);
and U32443 (N_32443,N_28410,N_28890);
or U32444 (N_32444,N_27641,N_28385);
nand U32445 (N_32445,N_29142,N_28321);
nand U32446 (N_32446,N_28897,N_27618);
xnor U32447 (N_32447,N_28498,N_28269);
nor U32448 (N_32448,N_28153,N_28835);
nand U32449 (N_32449,N_29993,N_28983);
nand U32450 (N_32450,N_28083,N_28359);
xnor U32451 (N_32451,N_29135,N_27513);
xor U32452 (N_32452,N_29231,N_29997);
xor U32453 (N_32453,N_28520,N_28194);
nand U32454 (N_32454,N_28169,N_29736);
xor U32455 (N_32455,N_29533,N_28764);
or U32456 (N_32456,N_27628,N_28480);
or U32457 (N_32457,N_27638,N_29108);
nand U32458 (N_32458,N_28451,N_28749);
nand U32459 (N_32459,N_29376,N_29689);
nand U32460 (N_32460,N_27922,N_29396);
nand U32461 (N_32461,N_28975,N_29986);
and U32462 (N_32462,N_28214,N_29875);
nand U32463 (N_32463,N_27634,N_29832);
xnor U32464 (N_32464,N_29723,N_27638);
xnor U32465 (N_32465,N_27968,N_29562);
nand U32466 (N_32466,N_27689,N_27517);
nor U32467 (N_32467,N_29061,N_28418);
nand U32468 (N_32468,N_29860,N_28244);
nor U32469 (N_32469,N_29532,N_29805);
nor U32470 (N_32470,N_28161,N_27572);
nand U32471 (N_32471,N_29203,N_27601);
xor U32472 (N_32472,N_28946,N_28669);
or U32473 (N_32473,N_28456,N_28674);
xnor U32474 (N_32474,N_28823,N_29326);
nand U32475 (N_32475,N_29703,N_28706);
and U32476 (N_32476,N_28412,N_29684);
or U32477 (N_32477,N_28688,N_28164);
nor U32478 (N_32478,N_28222,N_29612);
xnor U32479 (N_32479,N_28612,N_27862);
and U32480 (N_32480,N_27795,N_29609);
nor U32481 (N_32481,N_27711,N_29859);
xor U32482 (N_32482,N_27710,N_28848);
or U32483 (N_32483,N_29334,N_29244);
and U32484 (N_32484,N_27791,N_29338);
and U32485 (N_32485,N_27514,N_28045);
or U32486 (N_32486,N_28535,N_29844);
and U32487 (N_32487,N_28012,N_29785);
nor U32488 (N_32488,N_29594,N_28079);
or U32489 (N_32489,N_28039,N_29190);
nand U32490 (N_32490,N_28545,N_29396);
and U32491 (N_32491,N_29112,N_28826);
or U32492 (N_32492,N_27554,N_27975);
nor U32493 (N_32493,N_28257,N_29174);
nor U32494 (N_32494,N_27889,N_29112);
and U32495 (N_32495,N_29065,N_28882);
and U32496 (N_32496,N_29253,N_29776);
or U32497 (N_32497,N_29955,N_27564);
or U32498 (N_32498,N_28280,N_28118);
xnor U32499 (N_32499,N_29417,N_29892);
or U32500 (N_32500,N_31363,N_32135);
and U32501 (N_32501,N_31137,N_31457);
and U32502 (N_32502,N_31000,N_31646);
xor U32503 (N_32503,N_32461,N_31287);
and U32504 (N_32504,N_30686,N_31552);
and U32505 (N_32505,N_31184,N_31855);
nor U32506 (N_32506,N_31955,N_31674);
xnor U32507 (N_32507,N_32104,N_32311);
nor U32508 (N_32508,N_32299,N_30684);
nor U32509 (N_32509,N_31577,N_31224);
nor U32510 (N_32510,N_31571,N_31528);
or U32511 (N_32511,N_31477,N_31752);
nor U32512 (N_32512,N_31433,N_32405);
and U32513 (N_32513,N_31726,N_32001);
nand U32514 (N_32514,N_31089,N_31606);
nor U32515 (N_32515,N_32181,N_30907);
nor U32516 (N_32516,N_31352,N_31374);
and U32517 (N_32517,N_32221,N_31691);
xor U32518 (N_32518,N_31605,N_32367);
xnor U32519 (N_32519,N_30170,N_31220);
or U32520 (N_32520,N_31823,N_31312);
and U32521 (N_32521,N_32368,N_31159);
and U32522 (N_32522,N_31770,N_31749);
nor U32523 (N_32523,N_30177,N_32294);
and U32524 (N_32524,N_32000,N_31621);
nand U32525 (N_32525,N_32073,N_30388);
xnor U32526 (N_32526,N_30505,N_32011);
nand U32527 (N_32527,N_30963,N_30737);
nand U32528 (N_32528,N_31190,N_31108);
nor U32529 (N_32529,N_31171,N_31035);
nor U32530 (N_32530,N_31721,N_32373);
or U32531 (N_32531,N_30249,N_30998);
xnor U32532 (N_32532,N_31705,N_30860);
or U32533 (N_32533,N_31512,N_30054);
and U32534 (N_32534,N_31780,N_31596);
nand U32535 (N_32535,N_32089,N_30329);
nand U32536 (N_32536,N_32337,N_32121);
nand U32537 (N_32537,N_30022,N_31341);
nand U32538 (N_32538,N_30234,N_32485);
xnor U32539 (N_32539,N_31075,N_32374);
nor U32540 (N_32540,N_31722,N_30052);
and U32541 (N_32541,N_30470,N_30130);
and U32542 (N_32542,N_31856,N_30131);
or U32543 (N_32543,N_32490,N_31937);
nand U32544 (N_32544,N_31858,N_30550);
xor U32545 (N_32545,N_32290,N_32193);
xnor U32546 (N_32546,N_31655,N_30809);
and U32547 (N_32547,N_31815,N_32252);
nor U32548 (N_32548,N_32454,N_30944);
and U32549 (N_32549,N_30534,N_31515);
or U32550 (N_32550,N_30261,N_30033);
or U32551 (N_32551,N_31327,N_30578);
xnor U32552 (N_32552,N_31464,N_31603);
and U32553 (N_32553,N_30367,N_32344);
xor U32554 (N_32554,N_30735,N_32075);
and U32555 (N_32555,N_31015,N_30264);
or U32556 (N_32556,N_30306,N_30113);
xor U32557 (N_32557,N_30373,N_30082);
nor U32558 (N_32558,N_31439,N_30451);
nor U32559 (N_32559,N_30986,N_31878);
nor U32560 (N_32560,N_31521,N_30493);
nor U32561 (N_32561,N_30248,N_31670);
nor U32562 (N_32562,N_31056,N_30516);
nor U32563 (N_32563,N_30283,N_31767);
xor U32564 (N_32564,N_30830,N_31591);
or U32565 (N_32565,N_30947,N_31927);
or U32566 (N_32566,N_30340,N_31185);
nand U32567 (N_32567,N_32147,N_32394);
nand U32568 (N_32568,N_30974,N_30577);
and U32569 (N_32569,N_30657,N_31066);
xnor U32570 (N_32570,N_31947,N_31310);
xnor U32571 (N_32571,N_30148,N_30927);
xnor U32572 (N_32572,N_30659,N_30140);
xnor U32573 (N_32573,N_31420,N_31095);
or U32574 (N_32574,N_30818,N_30796);
nor U32575 (N_32575,N_30730,N_30997);
nor U32576 (N_32576,N_32307,N_32232);
nand U32577 (N_32577,N_31925,N_31934);
nand U32578 (N_32578,N_31756,N_32059);
and U32579 (N_32579,N_31747,N_32464);
xnor U32580 (N_32580,N_30583,N_30894);
xor U32581 (N_32581,N_30387,N_30060);
and U32582 (N_32582,N_30910,N_30554);
nand U32583 (N_32583,N_31261,N_32164);
nand U32584 (N_32584,N_31985,N_31134);
or U32585 (N_32585,N_31008,N_30840);
nor U32586 (N_32586,N_32424,N_32284);
nor U32587 (N_32587,N_32463,N_32286);
xnor U32588 (N_32588,N_30241,N_31544);
xnor U32589 (N_32589,N_30062,N_32324);
nor U32590 (N_32590,N_31584,N_31119);
or U32591 (N_32591,N_30473,N_30202);
nand U32592 (N_32592,N_32319,N_32036);
or U32593 (N_32593,N_30069,N_31582);
nor U32594 (N_32594,N_30533,N_32034);
xnor U32595 (N_32595,N_30197,N_31434);
and U32596 (N_32596,N_30806,N_31175);
nor U32597 (N_32597,N_32240,N_30708);
or U32598 (N_32598,N_31028,N_30147);
or U32599 (N_32599,N_31006,N_32019);
xor U32600 (N_32600,N_32358,N_31792);
nor U32601 (N_32601,N_30671,N_32316);
and U32602 (N_32602,N_31317,N_30602);
nor U32603 (N_32603,N_31850,N_31902);
and U32604 (N_32604,N_31413,N_30750);
xnor U32605 (N_32605,N_32277,N_31775);
and U32606 (N_32606,N_32106,N_32486);
nand U32607 (N_32607,N_31101,N_32428);
and U32608 (N_32608,N_31063,N_32079);
and U32609 (N_32609,N_32298,N_30002);
nand U32610 (N_32610,N_31798,N_32201);
nor U32611 (N_32611,N_32229,N_30629);
nand U32612 (N_32612,N_31208,N_31094);
xnor U32613 (N_32613,N_31510,N_30865);
nor U32614 (N_32614,N_30747,N_31225);
or U32615 (N_32615,N_30742,N_32012);
or U32616 (N_32616,N_31741,N_31305);
and U32617 (N_32617,N_30316,N_31717);
nand U32618 (N_32618,N_30838,N_30711);
nor U32619 (N_32619,N_30702,N_30591);
xnor U32620 (N_32620,N_32407,N_32381);
nor U32621 (N_32621,N_30411,N_32269);
and U32622 (N_32622,N_31841,N_30851);
or U32623 (N_32623,N_31758,N_31629);
xor U32624 (N_32624,N_32355,N_31529);
nor U32625 (N_32625,N_30418,N_30395);
or U32626 (N_32626,N_32396,N_31293);
xnor U32627 (N_32627,N_32005,N_31480);
xor U32628 (N_32628,N_31479,N_31386);
xor U32629 (N_32629,N_30468,N_31398);
xor U32630 (N_32630,N_30557,N_30523);
nand U32631 (N_32631,N_30749,N_31005);
and U32632 (N_32632,N_30981,N_31860);
nand U32633 (N_32633,N_31284,N_31755);
and U32634 (N_32634,N_31820,N_31594);
nor U32635 (N_32635,N_30076,N_30128);
nor U32636 (N_32636,N_31474,N_32209);
xor U32637 (N_32637,N_31728,N_31627);
nor U32638 (N_32638,N_30712,N_31754);
nor U32639 (N_32639,N_30887,N_30462);
nor U32640 (N_32640,N_32235,N_31407);
or U32641 (N_32641,N_32223,N_30649);
nor U32642 (N_32642,N_31126,N_30275);
nand U32643 (N_32643,N_30206,N_32077);
xor U32644 (N_32644,N_30541,N_30091);
nor U32645 (N_32645,N_32226,N_30567);
nand U32646 (N_32646,N_30905,N_30169);
nor U32647 (N_32647,N_30617,N_31631);
nand U32648 (N_32648,N_30695,N_30630);
xnor U32649 (N_32649,N_32222,N_31379);
and U32650 (N_32650,N_30487,N_31421);
nor U32651 (N_32651,N_31328,N_32369);
nand U32652 (N_32652,N_31781,N_31267);
nand U32653 (N_32653,N_31482,N_30080);
nand U32654 (N_32654,N_30237,N_30495);
xnor U32655 (N_32655,N_30719,N_30697);
and U32656 (N_32656,N_31554,N_31709);
nand U32657 (N_32657,N_30520,N_32078);
or U32658 (N_32658,N_31693,N_30476);
xnor U32659 (N_32659,N_31851,N_30627);
xnor U32660 (N_32660,N_31625,N_31213);
nand U32661 (N_32661,N_30492,N_30982);
nor U32662 (N_32662,N_31389,N_30077);
and U32663 (N_32663,N_32391,N_30159);
xor U32664 (N_32664,N_30603,N_30855);
nor U32665 (N_32665,N_30104,N_31710);
nor U32666 (N_32666,N_30420,N_30506);
nand U32667 (N_32667,N_31899,N_30588);
nand U32668 (N_32668,N_30208,N_31687);
nor U32669 (N_32669,N_31809,N_30439);
and U32670 (N_32670,N_31916,N_30435);
xor U32671 (N_32671,N_31524,N_30084);
and U32672 (N_32672,N_30030,N_32283);
xnor U32673 (N_32673,N_30326,N_30394);
nand U32674 (N_32674,N_30491,N_30587);
xnor U32675 (N_32675,N_30114,N_30460);
xor U32676 (N_32676,N_31959,N_30442);
or U32677 (N_32677,N_30977,N_32158);
nand U32678 (N_32678,N_31138,N_30662);
xnor U32679 (N_32679,N_30023,N_32388);
and U32680 (N_32680,N_30949,N_31014);
or U32681 (N_32681,N_30799,N_30536);
and U32682 (N_32682,N_31149,N_31172);
and U32683 (N_32683,N_31495,N_31800);
nand U32684 (N_32684,N_32033,N_30192);
nor U32685 (N_32685,N_30596,N_31251);
nand U32686 (N_32686,N_31321,N_31068);
nor U32687 (N_32687,N_30593,N_30848);
or U32688 (N_32688,N_30789,N_32418);
or U32689 (N_32689,N_31351,N_30215);
xor U32690 (N_32690,N_31200,N_30469);
nand U32691 (N_32691,N_30370,N_31437);
nand U32692 (N_32692,N_31083,N_30853);
or U32693 (N_32693,N_31361,N_31156);
nand U32694 (N_32694,N_30911,N_31219);
nand U32695 (N_32695,N_32429,N_32197);
xor U32696 (N_32696,N_31416,N_32180);
nor U32697 (N_32697,N_32025,N_31408);
xor U32698 (N_32698,N_30194,N_30872);
nor U32699 (N_32699,N_31968,N_32127);
or U32700 (N_32700,N_30106,N_31559);
and U32701 (N_32701,N_32145,N_31900);
or U32702 (N_32702,N_31714,N_31412);
nand U32703 (N_32703,N_31288,N_30444);
xor U32704 (N_32704,N_30416,N_30787);
xor U32705 (N_32705,N_30975,N_31122);
xnor U32706 (N_32706,N_32008,N_31587);
xnor U32707 (N_32707,N_32455,N_30824);
xnor U32708 (N_32708,N_30180,N_30272);
and U32709 (N_32709,N_30781,N_31253);
nor U32710 (N_32710,N_31565,N_30618);
nand U32711 (N_32711,N_30560,N_30297);
nand U32712 (N_32712,N_31024,N_31469);
xor U32713 (N_32713,N_32312,N_31338);
nand U32714 (N_32714,N_30762,N_32046);
xor U32715 (N_32715,N_31638,N_31103);
and U32716 (N_32716,N_31732,N_32257);
nand U32717 (N_32717,N_31729,N_31656);
xnor U32718 (N_32718,N_30384,N_30165);
nand U32719 (N_32719,N_30513,N_32132);
nand U32720 (N_32720,N_31074,N_30705);
or U32721 (N_32721,N_32271,N_32488);
xnor U32722 (N_32722,N_32082,N_31636);
xor U32723 (N_32723,N_32050,N_30223);
nor U32724 (N_32724,N_30814,N_32122);
xnor U32725 (N_32725,N_31192,N_30191);
or U32726 (N_32726,N_30526,N_31626);
xnor U32727 (N_32727,N_32364,N_31323);
and U32728 (N_32728,N_30563,N_30753);
or U32729 (N_32729,N_30284,N_30453);
and U32730 (N_32730,N_32128,N_31330);
and U32731 (N_32731,N_30324,N_30005);
and U32732 (N_32732,N_30361,N_31511);
nand U32733 (N_32733,N_32178,N_30979);
nand U32734 (N_32734,N_30196,N_30920);
xor U32735 (N_32735,N_31081,N_30669);
nor U32736 (N_32736,N_31611,N_31308);
nand U32737 (N_32737,N_32112,N_30939);
and U32738 (N_32738,N_31349,N_30932);
xnor U32739 (N_32739,N_31371,N_30549);
nor U32740 (N_32740,N_31981,N_31017);
or U32741 (N_32741,N_32047,N_31500);
and U32742 (N_32742,N_31977,N_31707);
nor U32743 (N_32743,N_30225,N_31622);
and U32744 (N_32744,N_31135,N_31071);
and U32745 (N_32745,N_31833,N_30802);
nand U32746 (N_32746,N_30508,N_31834);
or U32747 (N_32747,N_31206,N_30017);
or U32748 (N_32748,N_31654,N_30721);
xor U32749 (N_32749,N_32331,N_30770);
nand U32750 (N_32750,N_30123,N_31664);
and U32751 (N_32751,N_30689,N_30651);
and U32752 (N_32752,N_30294,N_32039);
xnor U32753 (N_32753,N_32218,N_31811);
xnor U32754 (N_32754,N_32148,N_30521);
or U32755 (N_32755,N_31797,N_32297);
or U32756 (N_32756,N_31842,N_31905);
and U32757 (N_32757,N_30958,N_32332);
nand U32758 (N_32758,N_32425,N_31906);
and U32759 (N_32759,N_31446,N_31169);
xnor U32760 (N_32760,N_30012,N_31547);
or U32761 (N_32761,N_30648,N_31372);
and U32762 (N_32762,N_31198,N_31356);
and U32763 (N_32763,N_31929,N_32109);
or U32764 (N_32764,N_31476,N_31618);
nor U32765 (N_32765,N_31933,N_30700);
and U32766 (N_32766,N_31576,N_31178);
xnor U32767 (N_32767,N_31525,N_30581);
or U32768 (N_32768,N_31730,N_32134);
and U32769 (N_32769,N_31228,N_30424);
nand U32770 (N_32770,N_31215,N_30646);
nor U32771 (N_32771,N_32048,N_30020);
xnor U32772 (N_32772,N_31771,N_30405);
xor U32773 (N_32773,N_32456,N_30585);
and U32774 (N_32774,N_30529,N_32460);
and U32775 (N_32775,N_31804,N_31111);
or U32776 (N_32776,N_32300,N_31316);
nor U32777 (N_32777,N_31144,N_30172);
xnor U32778 (N_32778,N_30778,N_31011);
and U32779 (N_32779,N_31816,N_32130);
or U32780 (N_32780,N_31617,N_31951);
nor U32781 (N_32781,N_30703,N_31233);
and U32782 (N_32782,N_31637,N_32414);
xnor U32783 (N_32783,N_31504,N_30790);
xnor U32784 (N_32784,N_31399,N_31969);
or U32785 (N_32785,N_32049,N_31678);
xor U32786 (N_32786,N_31166,N_31153);
or U32787 (N_32787,N_31946,N_31965);
nand U32788 (N_32788,N_30013,N_31904);
or U32789 (N_32789,N_31837,N_31684);
or U32790 (N_32790,N_31396,N_30210);
nor U32791 (N_32791,N_30976,N_32027);
or U32792 (N_32792,N_31537,N_31991);
and U32793 (N_32793,N_31073,N_31768);
xnor U32794 (N_32794,N_31419,N_31065);
and U32795 (N_32795,N_30782,N_30230);
and U32796 (N_32796,N_32435,N_31443);
and U32797 (N_32797,N_30378,N_30414);
and U32798 (N_32798,N_31868,N_30745);
nand U32799 (N_32799,N_30679,N_31864);
and U32800 (N_32800,N_31791,N_31869);
and U32801 (N_32801,N_31191,N_31086);
and U32802 (N_32802,N_32473,N_30347);
nand U32803 (N_32803,N_31845,N_31176);
nand U32804 (N_32804,N_31613,N_30663);
nand U32805 (N_32805,N_32317,N_30216);
or U32806 (N_32806,N_31049,N_30992);
and U32807 (N_32807,N_30654,N_31080);
and U32808 (N_32808,N_32443,N_31418);
and U32809 (N_32809,N_31325,N_30143);
nand U32810 (N_32810,N_32465,N_31647);
nand U32811 (N_32811,N_30537,N_30959);
or U32812 (N_32812,N_32053,N_31944);
nor U32813 (N_32813,N_32153,N_31533);
xnor U32814 (N_32814,N_32177,N_31846);
and U32815 (N_32815,N_31244,N_30883);
xnor U32816 (N_32816,N_30484,N_31831);
nand U32817 (N_32817,N_30503,N_30661);
xnor U32818 (N_32818,N_30859,N_31194);
xnor U32819 (N_32819,N_30168,N_31789);
nor U32820 (N_32820,N_31018,N_30984);
xor U32821 (N_32821,N_32475,N_32023);
nand U32822 (N_32822,N_31920,N_31827);
or U32823 (N_32823,N_32254,N_30293);
nor U32824 (N_32824,N_30380,N_30164);
nand U32825 (N_32825,N_31874,N_30183);
xor U32826 (N_32826,N_31562,N_30092);
nand U32827 (N_32827,N_31686,N_30058);
and U32828 (N_32828,N_30026,N_30300);
nor U32829 (N_32829,N_30229,N_30760);
nand U32830 (N_32830,N_32436,N_30097);
or U32831 (N_32831,N_31276,N_32335);
xor U32832 (N_32832,N_30610,N_30601);
xnor U32833 (N_32833,N_31197,N_32058);
and U32834 (N_32834,N_32244,N_30224);
nor U32835 (N_32835,N_32171,N_30948);
nand U32836 (N_32836,N_30885,N_31688);
nor U32837 (N_32837,N_31739,N_32412);
xnor U32838 (N_32838,N_31260,N_31569);
nand U32839 (N_32839,N_30674,N_30201);
nand U32840 (N_32840,N_32144,N_31272);
or U32841 (N_32841,N_31004,N_32092);
xnor U32842 (N_32842,N_30819,N_32207);
nand U32843 (N_32843,N_31513,N_30025);
nand U32844 (N_32844,N_31069,N_30010);
or U32845 (N_32845,N_31047,N_31844);
nor U32846 (N_32846,N_31683,N_32370);
or U32847 (N_32847,N_30954,N_30288);
nor U32848 (N_32848,N_31857,N_32494);
or U32849 (N_32849,N_30124,N_31802);
nor U32850 (N_32850,N_30652,N_31340);
nand U32851 (N_32851,N_30989,N_32433);
and U32852 (N_32852,N_31928,N_31903);
xnor U32853 (N_32853,N_32476,N_30685);
xor U32854 (N_32854,N_30792,N_31403);
nor U32855 (N_32855,N_32295,N_32184);
nor U32856 (N_32856,N_30021,N_31107);
or U32857 (N_32857,N_30723,N_30906);
nor U32858 (N_32858,N_31120,N_31404);
xor U32859 (N_32859,N_30346,N_30356);
xnor U32860 (N_32860,N_32227,N_30677);
nand U32861 (N_32861,N_30788,N_30573);
and U32862 (N_32862,N_30772,N_31990);
or U32863 (N_32863,N_31980,N_30009);
nor U32864 (N_32864,N_30323,N_30256);
xor U32865 (N_32865,N_31589,N_31189);
or U32866 (N_32866,N_30667,N_31652);
or U32867 (N_32867,N_30680,N_31865);
nand U32868 (N_32868,N_30886,N_30904);
xor U32869 (N_32869,N_32291,N_31359);
xor U32870 (N_32870,N_31973,N_30517);
and U32871 (N_32871,N_30795,N_30547);
nand U32872 (N_32872,N_31012,N_32131);
or U32873 (N_32873,N_32327,N_32115);
xor U32874 (N_32874,N_30957,N_30402);
nand U32875 (N_32875,N_32040,N_30100);
xnor U32876 (N_32876,N_30446,N_32007);
and U32877 (N_32877,N_32166,N_32438);
nand U32878 (N_32878,N_30511,N_31180);
nand U32879 (N_32879,N_30724,N_32497);
xor U32880 (N_32880,N_30973,N_32398);
xor U32881 (N_32881,N_30931,N_30112);
and U32882 (N_32882,N_32400,N_31556);
and U32883 (N_32883,N_31202,N_30915);
and U32884 (N_32884,N_31719,N_32155);
xor U32885 (N_32885,N_31348,N_32347);
or U32886 (N_32886,N_30457,N_31494);
xor U32887 (N_32887,N_30109,N_31291);
nor U32888 (N_32888,N_30706,N_30566);
xnor U32889 (N_32889,N_30709,N_31456);
xnor U32890 (N_32890,N_31431,N_31383);
or U32891 (N_32891,N_30423,N_31401);
or U32892 (N_32892,N_32483,N_30748);
nand U32893 (N_32893,N_31642,N_30360);
nand U32894 (N_32894,N_31790,N_32448);
xnor U32895 (N_32895,N_30909,N_31118);
nor U32896 (N_32896,N_30086,N_32100);
and U32897 (N_32897,N_31364,N_30339);
or U32898 (N_32898,N_30178,N_31373);
and U32899 (N_32899,N_32098,N_31640);
nand U32900 (N_32900,N_30896,N_30236);
nand U32901 (N_32901,N_32278,N_30632);
xor U32902 (N_32902,N_31209,N_30726);
nand U32903 (N_32903,N_31136,N_31901);
xor U32904 (N_32904,N_30968,N_32350);
nor U32905 (N_32905,N_32225,N_31639);
nor U32906 (N_32906,N_30313,N_31218);
or U32907 (N_32907,N_30683,N_32439);
xnor U32908 (N_32908,N_31092,N_31459);
or U32909 (N_32909,N_32070,N_31574);
xnor U32910 (N_32910,N_31117,N_31932);
and U32911 (N_32911,N_30144,N_32256);
or U32912 (N_32912,N_31058,N_32085);
or U32913 (N_32913,N_32310,N_32243);
xor U32914 (N_32914,N_31784,N_32138);
xnor U32915 (N_32915,N_30714,N_31539);
or U32916 (N_32916,N_30349,N_30090);
and U32917 (N_32917,N_32296,N_31295);
nand U32918 (N_32918,N_31343,N_31898);
and U32919 (N_32919,N_31313,N_30544);
nand U32920 (N_32920,N_31452,N_31745);
or U32921 (N_32921,N_30946,N_31948);
nand U32922 (N_32922,N_30893,N_30412);
or U32923 (N_32923,N_31806,N_30376);
nor U32924 (N_32924,N_32348,N_32251);
xnor U32925 (N_32925,N_30504,N_31566);
nor U32926 (N_32926,N_31884,N_31247);
xnor U32927 (N_32927,N_31822,N_31052);
xor U32928 (N_32928,N_32378,N_30155);
xnor U32929 (N_32929,N_30362,N_30564);
nor U32930 (N_32930,N_30372,N_32176);
nand U32931 (N_32931,N_30757,N_30592);
and U32932 (N_32932,N_30333,N_31173);
nand U32933 (N_32933,N_31516,N_32352);
nand U32934 (N_32934,N_30242,N_31971);
nand U32935 (N_32935,N_31394,N_30327);
nor U32936 (N_32936,N_31447,N_32343);
nand U32937 (N_32937,N_30892,N_30827);
or U32938 (N_32938,N_30950,N_32301);
nor U32939 (N_32939,N_32060,N_30785);
nor U32940 (N_32940,N_30068,N_30019);
or U32941 (N_32941,N_31645,N_30919);
and U32942 (N_32942,N_30273,N_31161);
or U32943 (N_32943,N_30660,N_30087);
nor U32944 (N_32944,N_31016,N_30214);
nand U32945 (N_32945,N_31579,N_31575);
and U32946 (N_32946,N_31685,N_30101);
and U32947 (N_32947,N_31873,N_31248);
nand U32948 (N_32948,N_31557,N_32273);
nor U32949 (N_32949,N_30638,N_32303);
or U32950 (N_32950,N_30040,N_30438);
nor U32951 (N_32951,N_31570,N_31380);
and U32952 (N_32952,N_31387,N_31914);
nor U32953 (N_32953,N_30133,N_30897);
xor U32954 (N_32954,N_32489,N_30157);
nor U32955 (N_32955,N_31155,N_31964);
nand U32956 (N_32956,N_31713,N_31774);
or U32957 (N_32957,N_30594,N_30315);
nor U32958 (N_32958,N_30923,N_30675);
nor U32959 (N_32959,N_31509,N_32140);
nand U32960 (N_32960,N_31098,N_32305);
xor U32961 (N_32961,N_31145,N_30797);
nand U32962 (N_32962,N_32189,N_31183);
nand U32963 (N_32963,N_31097,N_30319);
xor U32964 (N_32964,N_30153,N_30500);
or U32965 (N_32965,N_30239,N_32080);
xnor U32966 (N_32966,N_31182,N_30332);
nor U32967 (N_32967,N_31397,N_31677);
and U32968 (N_32968,N_30903,N_31564);
or U32969 (N_32969,N_31561,N_31283);
or U32970 (N_32970,N_30727,N_30676);
xor U32971 (N_32971,N_31473,N_30890);
nor U32972 (N_32972,N_30631,N_30694);
and U32973 (N_32973,N_31139,N_31852);
nor U32974 (N_32974,N_32013,N_31329);
nor U32975 (N_32975,N_31821,N_30690);
xor U32976 (N_32976,N_30783,N_31490);
nor U32977 (N_32977,N_30921,N_32204);
nor U32978 (N_32978,N_32212,N_31909);
and U32979 (N_32979,N_32107,N_30729);
xor U32980 (N_32980,N_31059,N_32194);
and U32981 (N_32981,N_31324,N_31021);
nand U32982 (N_32982,N_31376,N_31147);
nor U32983 (N_32983,N_31597,N_31548);
or U32984 (N_32984,N_31152,N_31370);
xnor U32985 (N_32985,N_31957,N_30067);
or U32986 (N_32986,N_30656,N_31801);
xnor U32987 (N_32987,N_32419,N_30812);
nand U32988 (N_32988,N_30138,N_32213);
nor U32989 (N_32989,N_31942,N_31384);
nor U32990 (N_32990,N_30364,N_30222);
or U32991 (N_32991,N_32123,N_30540);
nor U32992 (N_32992,N_30924,N_30546);
nor U32993 (N_32993,N_30441,N_31541);
xnor U32994 (N_32994,N_30996,N_32160);
or U32995 (N_32995,N_30119,N_31572);
nand U32996 (N_32996,N_31084,N_30490);
xnor U32997 (N_32997,N_32054,N_32441);
and U32998 (N_32998,N_30449,N_31275);
or U32999 (N_32999,N_30377,N_30158);
and U33000 (N_33000,N_31967,N_30953);
nand U33001 (N_33001,N_31993,N_30572);
or U33002 (N_33002,N_31355,N_31602);
xor U33003 (N_33003,N_31285,N_31440);
or U33004 (N_33004,N_30047,N_31249);
or U33005 (N_33005,N_30041,N_31950);
and U33006 (N_33006,N_32151,N_30514);
or U33007 (N_33007,N_31535,N_32259);
nand U33008 (N_33008,N_31924,N_31696);
or U33009 (N_33009,N_32173,N_30425);
nand U33010 (N_33010,N_30771,N_30003);
and U33011 (N_33011,N_32282,N_32466);
nand U33012 (N_33012,N_30985,N_31508);
or U33013 (N_33013,N_31326,N_31450);
or U33014 (N_33014,N_30379,N_31954);
or U33015 (N_33015,N_30409,N_30352);
xor U33016 (N_33016,N_32404,N_31615);
nand U33017 (N_33017,N_31826,N_31415);
xnor U33018 (N_33018,N_31881,N_30244);
and U33019 (N_33019,N_31381,N_30922);
or U33020 (N_33020,N_32234,N_32361);
nand U33021 (N_33021,N_31764,N_31143);
and U33022 (N_33022,N_30744,N_31493);
nor U33023 (N_33023,N_30382,N_32408);
nand U33024 (N_33024,N_31204,N_30718);
xor U33025 (N_33025,N_30562,N_30348);
nor U33026 (N_33026,N_32156,N_30358);
or U33027 (N_33027,N_31488,N_31553);
nor U33028 (N_33028,N_30485,N_30643);
and U33029 (N_33029,N_31299,N_31862);
or U33030 (N_33030,N_30483,N_31962);
nor U33031 (N_33031,N_31824,N_30877);
nand U33032 (N_33032,N_30681,N_32203);
xnor U33033 (N_33033,N_31038,N_31187);
and U33034 (N_33034,N_32289,N_31132);
nand U33035 (N_33035,N_32351,N_30688);
or U33036 (N_33036,N_32042,N_31045);
or U33037 (N_33037,N_30611,N_30290);
nor U33038 (N_33038,N_30752,N_30813);
or U33039 (N_33039,N_30761,N_30389);
nand U33040 (N_33040,N_31988,N_31742);
nand U33041 (N_33041,N_31506,N_30278);
xnor U33042 (N_33042,N_32270,N_30184);
nor U33043 (N_33043,N_30699,N_30552);
nor U33044 (N_33044,N_32190,N_30553);
or U33045 (N_33045,N_31672,N_30450);
xnor U33046 (N_33046,N_30042,N_32387);
xnor U33047 (N_33047,N_31778,N_31007);
nand U33048 (N_33048,N_30633,N_30386);
nand U33049 (N_33049,N_30967,N_30163);
and U33050 (N_33050,N_30151,N_31769);
nor U33051 (N_33051,N_31532,N_30050);
nor U33052 (N_33052,N_32264,N_30299);
nand U33053 (N_33053,N_30081,N_32093);
xor U33054 (N_33054,N_30755,N_30489);
or U33055 (N_33055,N_32102,N_31478);
nand U33056 (N_33056,N_30644,N_31499);
nor U33057 (N_33057,N_32434,N_31432);
or U33058 (N_33058,N_30861,N_32002);
and U33059 (N_33059,N_32457,N_30079);
xor U33060 (N_33060,N_30245,N_30149);
nand U33061 (N_33061,N_31245,N_30088);
and U33062 (N_33062,N_30863,N_32467);
xor U33063 (N_33063,N_31895,N_30066);
or U33064 (N_33064,N_31051,N_31703);
xor U33065 (N_33065,N_32272,N_30186);
xnor U33066 (N_33066,N_30637,N_31430);
or U33067 (N_33067,N_31830,N_31505);
nor U33068 (N_33068,N_30524,N_30837);
and U33069 (N_33069,N_30227,N_30807);
or U33070 (N_33070,N_31353,N_30055);
xor U33071 (N_33071,N_30137,N_32399);
and U33072 (N_33072,N_31633,N_31650);
nand U33073 (N_33073,N_30658,N_30545);
or U33074 (N_33074,N_30139,N_30117);
xor U33075 (N_33075,N_30046,N_30970);
nand U33076 (N_33076,N_30532,N_30353);
nor U33077 (N_33077,N_31926,N_30832);
or U33078 (N_33078,N_31810,N_31819);
and U33079 (N_33079,N_30276,N_31010);
xnor U33080 (N_33080,N_30664,N_31246);
xor U33081 (N_33081,N_31444,N_32265);
nor U33082 (N_33082,N_32302,N_30966);
and U33083 (N_33083,N_31375,N_32191);
xnor U33084 (N_33084,N_31391,N_32095);
xnor U33085 (N_33085,N_32413,N_30129);
nor U33086 (N_33086,N_30038,N_30103);
nand U33087 (N_33087,N_30995,N_30929);
xnor U33088 (N_33088,N_30775,N_32389);
or U33089 (N_33089,N_31787,N_30322);
nand U33090 (N_33090,N_30304,N_31188);
nand U33091 (N_33091,N_31581,N_31369);
and U33092 (N_33092,N_31216,N_31580);
nand U33093 (N_33093,N_31237,N_30597);
xor U33094 (N_33094,N_32246,N_30247);
xnor U33095 (N_33095,N_31170,N_30670);
and U33096 (N_33096,N_31257,N_30804);
and U33097 (N_33097,N_30821,N_32326);
nand U33098 (N_33098,N_30204,N_30808);
nand U33099 (N_33099,N_30342,N_32375);
and U33100 (N_33100,N_31736,N_32417);
nor U33101 (N_33101,N_30447,N_31518);
or U33102 (N_33102,N_31958,N_30135);
nand U33103 (N_33103,N_32141,N_30431);
and U33104 (N_33104,N_30120,N_32308);
nand U33105 (N_33105,N_32346,N_30616);
nor U33106 (N_33106,N_31592,N_31140);
and U33107 (N_33107,N_31673,N_32119);
nor U33108 (N_33108,N_32306,N_31264);
nand U33109 (N_33109,N_32187,N_31996);
and U33110 (N_33110,N_30875,N_30263);
and U33111 (N_33111,N_32161,N_30873);
nor U33112 (N_33112,N_30187,N_31799);
nand U33113 (N_33113,N_30965,N_31526);
nor U33114 (N_33114,N_31388,N_31099);
nor U33115 (N_33115,N_32149,N_32403);
or U33116 (N_33116,N_31953,N_30754);
or U33117 (N_33117,N_31410,N_30233);
xor U33118 (N_33118,N_30889,N_32238);
nor U33119 (N_33119,N_30127,N_32365);
nor U33120 (N_33120,N_31651,N_31207);
xor U33121 (N_33121,N_30898,N_32208);
and U33122 (N_33122,N_31461,N_31595);
nor U33123 (N_33123,N_32044,N_31885);
or U33124 (N_33124,N_31995,N_31718);
nand U33125 (N_33125,N_30502,N_30270);
and U33126 (N_33126,N_30570,N_31442);
nand U33127 (N_33127,N_30960,N_32220);
xnor U33128 (N_33128,N_31849,N_31502);
xnor U33129 (N_33129,N_31019,N_30285);
nand U33130 (N_33130,N_32334,N_31445);
or U33131 (N_33131,N_30878,N_30043);
and U33132 (N_33132,N_31542,N_30428);
xnor U33133 (N_33133,N_31455,N_30895);
nand U33134 (N_33134,N_30419,N_31105);
or U33135 (N_33135,N_30884,N_32322);
nand U33136 (N_33136,N_30255,N_30525);
nor U33137 (N_33137,N_30867,N_30018);
xor U33138 (N_33138,N_31875,N_31022);
and U33139 (N_33139,N_31630,N_30057);
nor U33140 (N_33140,N_31405,N_32239);
nor U33141 (N_33141,N_30941,N_31832);
nand U33142 (N_33142,N_30015,N_32081);
nand U33143 (N_33143,N_30328,N_31438);
and U33144 (N_33144,N_32250,N_30751);
or U33145 (N_33145,N_30369,N_30833);
and U33146 (N_33146,N_31365,N_30882);
or U33147 (N_33147,N_31619,N_31133);
xor U33148 (N_33148,N_30207,N_31039);
xor U33149 (N_33149,N_31311,N_32099);
xnor U33150 (N_33150,N_32329,N_30107);
nor U33151 (N_33151,N_32096,N_32136);
xnor U33152 (N_33152,N_31614,N_32342);
xnor U33153 (N_33153,N_31982,N_32219);
nand U33154 (N_33154,N_30831,N_30176);
nand U33155 (N_33155,N_30195,N_32360);
and U33156 (N_33156,N_32069,N_30917);
xor U33157 (N_33157,N_31839,N_31082);
nor U33158 (N_33158,N_31880,N_30037);
and U33159 (N_33159,N_30625,N_31690);
and U33160 (N_33160,N_31793,N_31304);
or U33161 (N_33161,N_31050,N_30518);
and U33162 (N_33162,N_32292,N_31417);
and U33163 (N_33163,N_31712,N_31436);
nand U33164 (N_33164,N_30391,N_31992);
and U33165 (N_33165,N_30980,N_30580);
or U33166 (N_33166,N_31658,N_32321);
nand U33167 (N_33167,N_32468,N_31448);
or U33168 (N_33168,N_32083,N_31912);
nor U33169 (N_33169,N_30971,N_31583);
nor U33170 (N_33170,N_30764,N_31231);
or U33171 (N_33171,N_30105,N_31393);
or U33172 (N_33172,N_31031,N_30810);
and U33173 (N_33173,N_32186,N_30118);
xnor U33174 (N_33174,N_30619,N_31130);
and U33175 (N_33175,N_31489,N_30598);
or U33176 (N_33176,N_30238,N_32432);
nor U33177 (N_33177,N_31377,N_31282);
or U33178 (N_33178,N_30188,N_31468);
nand U33179 (N_33179,N_31085,N_30189);
or U33180 (N_33180,N_32126,N_31514);
nand U33181 (N_33181,N_31277,N_31545);
and U33182 (N_33182,N_31307,N_31635);
or U33183 (N_33183,N_32260,N_31167);
or U33184 (N_33184,N_31250,N_32397);
nand U33185 (N_33185,N_32142,N_31843);
nand U33186 (N_33186,N_32110,N_32043);
xor U33187 (N_33187,N_31470,N_32280);
and U33188 (N_33188,N_31036,N_31040);
and U33189 (N_33189,N_31385,N_30612);
and U33190 (N_33190,N_31560,N_32315);
or U33191 (N_33191,N_30161,N_30182);
nor U33192 (N_33192,N_32236,N_30335);
nand U33193 (N_33193,N_31704,N_31861);
or U33194 (N_33194,N_30691,N_30620);
and U33195 (N_33195,N_30154,N_32359);
or U33196 (N_33196,N_32091,N_31700);
nand U33197 (N_33197,N_31866,N_30731);
and U33198 (N_33198,N_30743,N_31414);
nand U33199 (N_33199,N_32175,N_32031);
nor U33200 (N_33200,N_31817,N_31297);
and U33201 (N_33201,N_32195,N_30558);
and U33202 (N_33202,N_32470,N_31876);
nand U33203 (N_33203,N_32420,N_30413);
xnor U33204 (N_33204,N_32163,N_30219);
or U33205 (N_33205,N_30606,N_30028);
xor U33206 (N_33206,N_30952,N_30568);
nor U33207 (N_33207,N_31701,N_32143);
and U33208 (N_33208,N_30584,N_32192);
nand U33209 (N_33209,N_30136,N_30282);
and U33210 (N_33210,N_32041,N_31053);
or U33211 (N_33211,N_30308,N_30829);
nand U33212 (N_33212,N_30397,N_31970);
and U33213 (N_33213,N_31994,N_30759);
and U33214 (N_33214,N_32279,N_31634);
xnor U33215 (N_33215,N_31644,N_31760);
nand U33216 (N_33216,N_31205,N_30497);
or U33217 (N_33217,N_30928,N_31910);
xor U33218 (N_33218,N_30271,N_30857);
or U33219 (N_33219,N_32495,N_30434);
nor U33220 (N_33220,N_31121,N_32150);
xnor U33221 (N_33221,N_31274,N_30539);
or U33222 (N_33222,N_31961,N_30466);
and U33223 (N_33223,N_30515,N_31600);
and U33224 (N_33224,N_31344,N_31649);
or U33225 (N_33225,N_30260,N_32016);
or U33226 (N_33226,N_31854,N_32032);
or U33227 (N_33227,N_31057,N_30576);
and U33228 (N_33228,N_30717,N_32022);
and U33229 (N_33229,N_31350,N_31115);
nand U33230 (N_33230,N_32182,N_32068);
or U33231 (N_33231,N_30150,N_30478);
and U33232 (N_33232,N_30543,N_31550);
nor U33233 (N_33233,N_30266,N_30701);
nor U33234 (N_33234,N_30032,N_32314);
nand U33235 (N_33235,N_30056,N_31503);
nor U33236 (N_33236,N_31923,N_32167);
nand U33237 (N_33237,N_31695,N_30286);
nor U33238 (N_33238,N_30226,N_31867);
nor U33239 (N_33239,N_31657,N_31694);
and U33240 (N_33240,N_31661,N_30209);
xnor U33241 (N_33241,N_31894,N_31314);
and U33242 (N_33242,N_31668,N_31471);
nand U33243 (N_33243,N_30199,N_30988);
and U33244 (N_33244,N_31632,N_30574);
xor U33245 (N_33245,N_31720,N_30063);
nor U33246 (N_33246,N_32076,N_31662);
nor U33247 (N_33247,N_32274,N_32262);
nor U33248 (N_33248,N_32382,N_30728);
xor U33249 (N_33249,N_31236,N_30203);
nand U33250 (N_33250,N_31847,N_31271);
nor U33251 (N_33251,N_31429,N_31232);
or U33252 (N_33252,N_30693,N_30331);
nor U33253 (N_33253,N_32472,N_31983);
nand U33254 (N_33254,N_32062,N_30942);
nor U33255 (N_33255,N_31226,N_31978);
xor U33256 (N_33256,N_31681,N_31241);
and U33257 (N_33257,N_30801,N_31612);
nor U33258 (N_33258,N_32288,N_30647);
nor U33259 (N_33259,N_31104,N_31240);
and U33260 (N_33260,N_30421,N_31346);
nand U33261 (N_33261,N_30854,N_32216);
or U33262 (N_33262,N_31146,N_31788);
nor U33263 (N_33263,N_30531,N_32383);
nor U33264 (N_33264,N_30623,N_30142);
or U33265 (N_33265,N_30064,N_30987);
nor U33266 (N_33266,N_30437,N_31141);
and U33267 (N_33267,N_31339,N_31620);
nand U33268 (N_33268,N_31289,N_31064);
or U33269 (N_33269,N_31002,N_30350);
nand U33270 (N_33270,N_32453,N_31254);
nor U33271 (N_33271,N_31072,N_30556);
nor U33272 (N_33272,N_32372,N_30014);
nand U33273 (N_33273,N_30488,N_31616);
or U33274 (N_33274,N_30211,N_31777);
and U33275 (N_33275,N_32117,N_32353);
nor U33276 (N_33276,N_32478,N_31882);
nand U33277 (N_33277,N_31917,N_32379);
nand U33278 (N_33278,N_32371,N_31534);
nor U33279 (N_33279,N_31794,N_31302);
nand U33280 (N_33280,N_32174,N_30374);
nor U33281 (N_33281,N_30609,N_30075);
and U33282 (N_33282,N_30626,N_30912);
and U33283 (N_33283,N_30213,N_31258);
and U33284 (N_33284,N_30707,N_31268);
and U33285 (N_33285,N_30432,N_30035);
nor U33286 (N_33286,N_31999,N_31949);
xor U33287 (N_33287,N_30825,N_30093);
and U33288 (N_33288,N_30926,N_30604);
nor U33289 (N_33289,N_30471,N_30653);
or U33290 (N_33290,N_31522,N_30141);
xnor U33291 (N_33291,N_31003,N_31214);
xnor U33292 (N_33292,N_30768,N_31142);
nor U33293 (N_33293,N_31689,N_32323);
or U33294 (N_33294,N_30108,N_30341);
and U33295 (N_33295,N_30070,N_30668);
nand U33296 (N_33296,N_31838,N_31485);
nand U33297 (N_33297,N_30280,N_30852);
nand U33298 (N_33298,N_30951,N_31222);
or U33299 (N_33299,N_30682,N_30710);
nor U33300 (N_33300,N_31062,N_31676);
xnor U33301 (N_33301,N_30846,N_30368);
and U33302 (N_33302,N_31731,N_30309);
or U33303 (N_33303,N_30933,N_30687);
xor U33304 (N_33304,N_31915,N_31037);
nor U33305 (N_33305,N_30044,N_32045);
xor U33306 (N_33306,N_31347,N_30793);
xor U33307 (N_33307,N_31598,N_31734);
or U33308 (N_33308,N_30561,N_30371);
nand U33309 (N_33309,N_30452,N_31956);
xor U33310 (N_33310,N_31892,N_31578);
nand U33311 (N_33311,N_32275,N_30870);
and U33312 (N_33312,N_30841,N_31335);
xor U33313 (N_33313,N_31853,N_32354);
or U33314 (N_33314,N_30815,N_30779);
and U33315 (N_33315,N_31124,N_31716);
and U33316 (N_33316,N_32090,N_30480);
or U33317 (N_33317,N_30102,N_30672);
nor U33318 (N_33318,N_32015,N_31773);
xor U33319 (N_33319,N_30298,N_30869);
nand U33320 (N_33320,N_32196,N_32451);
nand U33321 (N_33321,N_31706,N_30408);
xnor U33322 (N_33322,N_30039,N_30363);
nand U33323 (N_33323,N_31536,N_31628);
nand U33324 (N_33324,N_31466,N_31342);
nor U33325 (N_33325,N_30048,N_30880);
or U33326 (N_33326,N_32487,N_30252);
or U33327 (N_33327,N_30758,N_31259);
or U33328 (N_33328,N_31828,N_31738);
nor U33329 (N_33329,N_30404,N_31114);
xor U33330 (N_33330,N_30868,N_31060);
xor U33331 (N_33331,N_30393,N_30258);
or U33332 (N_33332,N_30605,N_31496);
or U33333 (N_33333,N_31859,N_30881);
and U33334 (N_33334,N_31551,N_30253);
and U33335 (N_33335,N_30715,N_30914);
nand U33336 (N_33336,N_30295,N_31733);
nand U33337 (N_33337,N_30736,N_30218);
nor U33338 (N_33338,N_30330,N_30822);
or U33339 (N_33339,N_30134,N_31692);
xnor U33340 (N_33340,N_30673,N_32065);
xor U33341 (N_33341,N_31125,N_31026);
nor U33342 (N_33342,N_30956,N_31697);
or U33343 (N_33343,N_31221,N_32410);
and U33344 (N_33344,N_31938,N_30791);
nand U33345 (N_33345,N_32318,N_32146);
and U33346 (N_33346,N_32035,N_30365);
nand U33347 (N_33347,N_30579,N_32345);
xor U33348 (N_33348,N_32480,N_31201);
nor U33349 (N_33349,N_31320,N_31593);
and U33350 (N_33350,N_30834,N_30257);
and U33351 (N_33351,N_31540,N_30351);
and U33352 (N_33352,N_31520,N_32021);
xnor U33353 (N_33353,N_30190,N_30876);
or U33354 (N_33354,N_31046,N_31997);
xor U33355 (N_33355,N_30990,N_31402);
and U33356 (N_33356,N_31523,N_32409);
nor U33357 (N_33357,N_32014,N_31239);
xor U33358 (N_33358,N_30221,N_30314);
nand U33359 (N_33359,N_31280,N_30463);
nor U33360 (N_33360,N_31273,N_30879);
nand U33361 (N_33361,N_31186,N_31484);
nor U33362 (N_33362,N_30011,N_30542);
or U33363 (N_33363,N_31779,N_32137);
or U33364 (N_33364,N_32169,N_30589);
or U33365 (N_33365,N_31425,N_32423);
nor U33366 (N_33366,N_30805,N_31588);
and U33367 (N_33367,N_31610,N_31196);
nor U33368 (N_33368,N_31945,N_30800);
xor U33369 (N_33369,N_30325,N_31034);
nand U33370 (N_33370,N_31362,N_32258);
or U33371 (N_33371,N_32411,N_32482);
nand U33372 (N_33372,N_30527,N_32052);
or U33373 (N_33373,N_31426,N_31643);
xnor U33374 (N_33374,N_31727,N_32263);
and U33375 (N_33375,N_30918,N_32484);
nor U33376 (N_33376,N_30955,N_30078);
and U33377 (N_33377,N_32320,N_30571);
nand U33378 (N_33378,N_32336,N_32471);
nand U33379 (N_33379,N_30235,N_30465);
xor U33380 (N_33380,N_30555,N_31546);
xnor U33381 (N_33381,N_31428,N_30908);
xor U33382 (N_33382,N_31702,N_30089);
nor U33383 (N_33383,N_30519,N_31812);
nor U33384 (N_33384,N_30004,N_32442);
xnor U33385 (N_33385,N_31803,N_30937);
nor U33386 (N_33386,N_32481,N_30375);
nor U33387 (N_33387,N_30045,N_30641);
xnor U33388 (N_33388,N_32458,N_31212);
xnor U33389 (N_33389,N_31199,N_31491);
xor U33390 (N_33390,N_30481,N_30121);
nor U33391 (N_33391,N_31863,N_30498);
nand U33392 (N_33392,N_32237,N_31737);
and U33393 (N_33393,N_31814,N_31931);
nor U33394 (N_33394,N_31076,N_31744);
and U33395 (N_33395,N_30036,N_31487);
and U33396 (N_33396,N_30072,N_32325);
xnor U33397 (N_33397,N_32188,N_30551);
and U33398 (N_33398,N_30443,N_31918);
xor U33399 (N_33399,N_31030,N_32198);
xor U33400 (N_33400,N_30334,N_32010);
or U33401 (N_33401,N_30359,N_32415);
nor U33402 (N_33402,N_31558,N_31102);
or U33403 (N_33403,N_32444,N_31795);
or U33404 (N_33404,N_30071,N_31337);
nand U33405 (N_33405,N_30845,N_31735);
nor U33406 (N_33406,N_30292,N_31160);
and U33407 (N_33407,N_32055,N_32452);
and U33408 (N_33408,N_30962,N_30243);
xnor U33409 (N_33409,N_31263,N_31252);
and U33410 (N_33410,N_31998,N_30399);
or U33411 (N_33411,N_30994,N_30512);
or U33412 (N_33412,N_31032,N_31041);
or U33413 (N_33413,N_31501,N_32431);
and U33414 (N_33414,N_30355,N_32430);
and U33415 (N_33415,N_32267,N_32061);
xor U33416 (N_33416,N_30776,N_31519);
xnor U33417 (N_33417,N_32214,N_32063);
and U33418 (N_33418,N_30624,N_31129);
or U33419 (N_33419,N_30240,N_30251);
nor U33420 (N_33420,N_31266,N_32168);
or U33421 (N_33421,N_32479,N_32009);
nor U33422 (N_33422,N_31292,N_32356);
nor U33423 (N_33423,N_30455,N_31357);
or U33424 (N_33424,N_31013,N_30398);
nor U33425 (N_33425,N_32057,N_31762);
and U33426 (N_33426,N_30741,N_31483);
nand U33427 (N_33427,N_32018,N_31127);
nand U33428 (N_33428,N_31077,N_30510);
xnor U33429 (N_33429,N_32037,N_31406);
or U33430 (N_33430,N_31893,N_30132);
nor U33431 (N_33431,N_30769,N_31462);
or U33432 (N_33432,N_31128,N_30392);
nand U33433 (N_33433,N_32459,N_31987);
nand U33434 (N_33434,N_32477,N_32385);
nor U33435 (N_33435,N_30467,N_30820);
and U33436 (N_33436,N_30738,N_32124);
and U33437 (N_33437,N_31256,N_30001);
nor U33438 (N_33438,N_30842,N_32384);
and U33439 (N_33439,N_31671,N_31441);
xnor U33440 (N_33440,N_30847,N_32255);
nor U33441 (N_33441,N_31667,N_31230);
nor U33442 (N_33442,N_31919,N_31151);
xnor U33443 (N_33443,N_30642,N_32245);
and U33444 (N_33444,N_31163,N_31300);
nor U33445 (N_33445,N_31911,N_30530);
or U33446 (N_33446,N_32445,N_32103);
nor U33447 (N_33447,N_32120,N_30740);
and U33448 (N_33448,N_30798,N_30410);
or U33449 (N_33449,N_31223,N_30343);
nor U33450 (N_33450,N_32200,N_30575);
nand U33451 (N_33451,N_32496,N_31586);
nor U33452 (N_33452,N_31044,N_32217);
nand U33453 (N_33453,N_32401,N_30274);
nor U33454 (N_33454,N_31048,N_30628);
and U33455 (N_33455,N_31422,N_30034);
xnor U33456 (N_33456,N_31608,N_30704);
nor U33457 (N_33457,N_31748,N_32133);
nor U33458 (N_33458,N_30051,N_31877);
nand U33459 (N_33459,N_31660,N_31984);
and U33460 (N_33460,N_32172,N_30780);
and U33461 (N_33461,N_30016,N_31243);
and U33462 (N_33462,N_30640,N_31935);
nand U33463 (N_33463,N_30174,N_31179);
and U33464 (N_33464,N_31067,N_31623);
and U33465 (N_33465,N_31162,N_32030);
nand U33466 (N_33466,N_31897,N_30231);
xor U33467 (N_33467,N_31460,N_30265);
xnor U33468 (N_33468,N_31211,N_32094);
nand U33469 (N_33469,N_31113,N_30765);
and U33470 (N_33470,N_32101,N_32421);
and U33471 (N_33471,N_31517,N_30725);
nand U33472 (N_33472,N_30116,N_31679);
nor U33473 (N_33473,N_30722,N_30115);
or U33474 (N_33474,N_32125,N_31367);
and U33475 (N_33475,N_31451,N_31989);
and U33476 (N_33476,N_30307,N_30301);
xor U33477 (N_33477,N_31235,N_31543);
xnor U33478 (N_33478,N_30417,N_31467);
and U33479 (N_33479,N_30993,N_30175);
nor U33480 (N_33480,N_30538,N_31322);
xor U33481 (N_33481,N_32159,N_30528);
or U33482 (N_33482,N_30259,N_30850);
nand U33483 (N_33483,N_30179,N_30773);
xor U33484 (N_33484,N_31939,N_30716);
or U33485 (N_33485,N_30366,N_32051);
xnor U33486 (N_33486,N_30160,N_32437);
and U33487 (N_33487,N_30167,N_31109);
nor U33488 (N_33488,N_31818,N_31465);
nor U33489 (N_33489,N_31298,N_32499);
xor U33490 (N_33490,N_32261,N_30999);
nor U33491 (N_33491,N_31497,N_30582);
nor U33492 (N_33492,N_31808,N_31829);
xor U33493 (N_33493,N_30499,N_30650);
nor U33494 (N_33494,N_31055,N_31458);
nor U33495 (N_33495,N_32248,N_31708);
or U33496 (N_33496,N_31723,N_31871);
nor U33497 (N_33497,N_32422,N_31663);
xnor U33498 (N_33498,N_32392,N_31070);
or U33499 (N_33499,N_31492,N_31123);
xnor U33500 (N_33500,N_31020,N_32313);
xnor U33501 (N_33501,N_32330,N_31116);
and U33502 (N_33502,N_32108,N_31262);
nor U33503 (N_33503,N_30445,N_30978);
and U33504 (N_33504,N_30635,N_32020);
or U33505 (N_33505,N_31096,N_32242);
or U33506 (N_33506,N_31358,N_30613);
nor U33507 (N_33507,N_31033,N_30479);
or U33508 (N_33508,N_30337,N_30277);
nand U33509 (N_33509,N_31607,N_30152);
xnor U33510 (N_33510,N_31336,N_30902);
nor U33511 (N_33511,N_30666,N_31411);
and U33512 (N_33512,N_32241,N_32028);
xnor U33513 (N_33513,N_30913,N_30073);
or U33514 (N_33514,N_31963,N_31242);
and U33515 (N_33515,N_31825,N_30049);
or U33516 (N_33516,N_30496,N_31725);
or U33517 (N_33517,N_30823,N_30031);
nand U33518 (N_33518,N_30099,N_30472);
nand U33519 (N_33519,N_32199,N_31281);
xnor U33520 (N_33520,N_32402,N_31889);
nor U33521 (N_33521,N_30983,N_30569);
xnor U33522 (N_33522,N_30145,N_30767);
and U33523 (N_33523,N_32224,N_32165);
and U33524 (N_33524,N_30461,N_31751);
nor U33525 (N_33525,N_30459,N_31354);
or U33526 (N_33526,N_32230,N_31746);
xor U33527 (N_33527,N_32211,N_32427);
xor U33528 (N_33528,N_31168,N_31395);
and U33529 (N_33529,N_31093,N_31382);
and U33530 (N_33530,N_30849,N_30816);
xor U33531 (N_33531,N_31887,N_32304);
nand U33532 (N_33532,N_31786,N_31486);
or U33533 (N_33533,N_30925,N_30794);
nand U33534 (N_33534,N_30456,N_30474);
or U33535 (N_33535,N_30900,N_30548);
and U33536 (N_33536,N_30430,N_31079);
and U33537 (N_33537,N_32349,N_31835);
xnor U33538 (N_33538,N_30720,N_30279);
nand U33539 (N_33539,N_32162,N_31908);
and U33540 (N_33540,N_31699,N_32249);
xnor U33541 (N_33541,N_31409,N_31807);
and U33542 (N_33542,N_30422,N_31174);
nor U33543 (N_33543,N_31682,N_31940);
or U33544 (N_33544,N_31238,N_30622);
nand U33545 (N_33545,N_30166,N_30390);
nor U33546 (N_33546,N_30608,N_30381);
and U33547 (N_33547,N_32339,N_32114);
xor U33548 (N_33548,N_31765,N_31648);
or U33549 (N_33549,N_30318,N_30171);
nand U33550 (N_33550,N_31848,N_30267);
and U33551 (N_33551,N_31227,N_31840);
or U33552 (N_33552,N_32268,N_30338);
nand U33553 (N_33553,N_30940,N_32017);
or U33554 (N_33554,N_31680,N_30501);
nand U33555 (N_33555,N_32498,N_31315);
or U33556 (N_33556,N_30864,N_32366);
and U33557 (N_33557,N_31531,N_30065);
or U33558 (N_33558,N_32416,N_31234);
or U33559 (N_33559,N_31872,N_30305);
nand U33560 (N_33560,N_30427,N_31270);
or U33561 (N_33561,N_32293,N_30599);
nor U33562 (N_33562,N_30111,N_30053);
nand U33563 (N_33563,N_30639,N_31165);
nor U33564 (N_33564,N_31555,N_32056);
nor U33565 (N_33565,N_31331,N_30839);
or U33566 (N_33566,N_30836,N_31296);
nand U33567 (N_33567,N_32084,N_31100);
or U33568 (N_33568,N_31930,N_30426);
nor U33569 (N_33569,N_31599,N_30938);
and U33570 (N_33570,N_31061,N_31665);
nand U33571 (N_33571,N_31319,N_31776);
nor U33572 (N_33572,N_30858,N_31400);
and U33573 (N_33573,N_31255,N_31907);
and U33574 (N_33574,N_32006,N_30345);
nor U33575 (N_33575,N_30269,N_32491);
xnor U33576 (N_33576,N_31698,N_31886);
nor U33577 (N_33577,N_30595,N_32449);
and U33578 (N_33578,N_31110,N_30185);
and U33579 (N_33579,N_30407,N_31890);
nor U33580 (N_33580,N_30655,N_31294);
and U33581 (N_33581,N_31624,N_31042);
nor U33582 (N_33582,N_32253,N_30291);
or U33583 (N_33583,N_31743,N_31345);
nand U33584 (N_33584,N_31766,N_30110);
nand U33585 (N_33585,N_31805,N_30385);
xor U33586 (N_33586,N_30943,N_31278);
xnor U33587 (N_33587,N_30429,N_31392);
nand U33588 (N_33588,N_30934,N_31427);
xor U33589 (N_33589,N_30636,N_30826);
or U33590 (N_33590,N_31750,N_31879);
nand U33591 (N_33591,N_31568,N_30310);
xnor U33592 (N_33592,N_32447,N_32474);
xor U33593 (N_33593,N_30312,N_30535);
or U33594 (N_33594,N_31783,N_30205);
nor U33595 (N_33595,N_31029,N_30126);
and U33596 (N_33596,N_32287,N_31936);
xor U33597 (N_33597,N_32440,N_30094);
xnor U33598 (N_33598,N_32071,N_31043);
or U33599 (N_33599,N_32111,N_30763);
or U33600 (N_33600,N_31001,N_30321);
xnor U33601 (N_33601,N_31027,N_30400);
nand U33602 (N_33602,N_30181,N_32333);
xor U33603 (N_33603,N_31157,N_31360);
or U33604 (N_33604,N_30396,N_31941);
or U33605 (N_33605,N_30733,N_31154);
xor U33606 (N_33606,N_32064,N_32170);
or U33607 (N_33607,N_30586,N_31922);
nor U33608 (N_33608,N_30024,N_32139);
nor U33609 (N_33609,N_30007,N_30317);
and U33610 (N_33610,N_30228,N_31195);
xnor U33611 (N_33611,N_31475,N_31217);
nor U33612 (N_33612,N_30436,N_30098);
and U33613 (N_33613,N_31763,N_31366);
nor U33614 (N_33614,N_32185,N_31921);
and U33615 (N_33615,N_31290,N_30406);
or U33616 (N_33616,N_32357,N_30698);
or U33617 (N_33617,N_31158,N_32362);
xor U33618 (N_33618,N_30507,N_30250);
and U33619 (N_33619,N_31883,N_31573);
or U33620 (N_33620,N_31424,N_31025);
xor U33621 (N_33621,N_30969,N_30083);
nor U33622 (N_33622,N_31054,N_31472);
xnor U33623 (N_33623,N_31666,N_32247);
nor U33624 (N_33624,N_32328,N_31943);
and U33625 (N_33625,N_30354,N_30433);
xnor U33626 (N_33626,N_31870,N_30200);
or U33627 (N_33627,N_30696,N_31567);
and U33628 (N_33628,N_30732,N_30008);
or U33629 (N_33629,N_30146,N_31390);
or U33630 (N_33630,N_30254,N_31481);
and U33631 (N_33631,N_30383,N_30835);
nand U33632 (N_33632,N_30930,N_32086);
xor U33633 (N_33633,N_30494,N_32380);
and U33634 (N_33634,N_30000,N_30482);
nor U33635 (N_33635,N_30756,N_30156);
and U33636 (N_33636,N_31112,N_30475);
and U33637 (N_33637,N_32228,N_31090);
nand U33638 (N_33638,N_30173,N_31753);
or U33639 (N_33639,N_31210,N_30486);
nand U33640 (N_33640,N_30006,N_32233);
nand U33641 (N_33641,N_30888,N_31150);
nor U33642 (N_33642,N_31590,N_30678);
xor U33643 (N_33643,N_30122,N_30289);
nor U33644 (N_33644,N_32088,N_30125);
and U33645 (N_33645,N_30320,N_32340);
nor U33646 (N_33646,N_30336,N_32395);
xor U33647 (N_33647,N_31891,N_31009);
nor U33648 (N_33648,N_31975,N_31301);
and U33649 (N_33649,N_31585,N_30899);
or U33650 (N_33650,N_31813,N_32309);
and U33651 (N_33651,N_32087,N_30734);
or U33652 (N_33652,N_30936,N_30162);
or U33653 (N_33653,N_30746,N_31265);
nand U33654 (N_33654,N_31498,N_32215);
and U33655 (N_33655,N_31269,N_32118);
xnor U33656 (N_33656,N_30862,N_30621);
and U33657 (N_33657,N_32157,N_31423);
xnor U33658 (N_33658,N_30262,N_30344);
xor U33659 (N_33659,N_30945,N_30246);
and U33660 (N_33660,N_30607,N_32026);
nand U33661 (N_33661,N_30600,N_32276);
xor U33662 (N_33662,N_30991,N_31796);
or U33663 (N_33663,N_30972,N_32129);
nand U33664 (N_33664,N_31023,N_31659);
nand U33665 (N_33665,N_32105,N_31549);
and U33666 (N_33666,N_31334,N_31836);
and U33667 (N_33667,N_31966,N_30212);
and U33668 (N_33668,N_30448,N_30828);
nor U33669 (N_33669,N_32462,N_31454);
and U33670 (N_33670,N_31952,N_30844);
and U33671 (N_33671,N_30665,N_31675);
nand U33672 (N_33672,N_32004,N_30891);
and U33673 (N_33673,N_31976,N_31986);
nor U33674 (N_33674,N_30059,N_32446);
and U33675 (N_33675,N_30784,N_31530);
nand U33676 (N_33676,N_32003,N_32183);
nand U33677 (N_33677,N_32024,N_31641);
or U33678 (N_33678,N_31785,N_30522);
xnor U33679 (N_33679,N_31177,N_32285);
nand U33680 (N_33680,N_31229,N_30096);
xor U33681 (N_33681,N_30692,N_31507);
and U33682 (N_33682,N_30027,N_30843);
xnor U33683 (N_33683,N_31088,N_30916);
or U33684 (N_33684,N_32074,N_31979);
nand U33685 (N_33685,N_30401,N_30811);
or U33686 (N_33686,N_30464,N_32493);
or U33687 (N_33687,N_30287,N_31453);
and U33688 (N_33688,N_32377,N_32492);
and U33689 (N_33689,N_31368,N_32072);
and U33690 (N_33690,N_31286,N_30454);
xnor U33691 (N_33691,N_30440,N_32038);
and U33692 (N_33692,N_31740,N_31131);
and U33693 (N_33693,N_31527,N_30074);
xnor U33694 (N_33694,N_31669,N_31193);
nand U33695 (N_33695,N_32210,N_31106);
nor U33696 (N_33696,N_30281,N_30774);
nand U33697 (N_33697,N_31761,N_31724);
nor U33698 (N_33698,N_30590,N_30901);
nor U33699 (N_33699,N_30634,N_31896);
or U33700 (N_33700,N_30232,N_31601);
or U33701 (N_33701,N_31960,N_30964);
nand U33702 (N_33702,N_31609,N_31164);
nand U33703 (N_33703,N_31463,N_30217);
or U33704 (N_33704,N_30615,N_30029);
nand U33705 (N_33705,N_31757,N_30357);
or U33706 (N_33706,N_32341,N_30311);
nand U33707 (N_33707,N_30403,N_30061);
xor U33708 (N_33708,N_31087,N_31782);
xnor U33709 (N_33709,N_30866,N_30766);
xor U33710 (N_33710,N_30415,N_30803);
nor U33711 (N_33711,N_30198,N_31279);
nor U33712 (N_33712,N_30220,N_30961);
xnor U33713 (N_33713,N_32406,N_31759);
and U33714 (N_33714,N_30645,N_30095);
nand U33715 (N_33715,N_31653,N_32266);
xor U33716 (N_33716,N_30509,N_31181);
nand U33717 (N_33717,N_31711,N_32469);
or U33718 (N_33718,N_31913,N_32029);
and U33719 (N_33719,N_31604,N_30477);
or U33720 (N_33720,N_32202,N_31309);
xnor U33721 (N_33721,N_30559,N_32067);
xnor U33722 (N_33722,N_31538,N_30614);
nand U33723 (N_33723,N_30786,N_31449);
nand U33724 (N_33724,N_32393,N_31148);
or U33725 (N_33725,N_32179,N_30458);
nand U33726 (N_33726,N_30565,N_32152);
xor U33727 (N_33727,N_31435,N_31306);
xnor U33728 (N_33728,N_30268,N_30713);
nor U33729 (N_33729,N_31772,N_32386);
nor U33730 (N_33730,N_31078,N_30739);
nor U33731 (N_33731,N_31203,N_32116);
nor U33732 (N_33732,N_30296,N_31332);
xor U33733 (N_33733,N_32390,N_31333);
xnor U33734 (N_33734,N_32376,N_31378);
xor U33735 (N_33735,N_30303,N_31563);
xnor U33736 (N_33736,N_31972,N_32066);
and U33737 (N_33737,N_30777,N_32338);
and U33738 (N_33738,N_31303,N_30856);
or U33739 (N_33739,N_30193,N_32113);
xor U33740 (N_33740,N_31974,N_32426);
or U33741 (N_33741,N_30817,N_30085);
xor U33742 (N_33742,N_32450,N_30874);
xor U33743 (N_33743,N_30871,N_30302);
nor U33744 (N_33744,N_32154,N_31091);
or U33745 (N_33745,N_32363,N_32205);
or U33746 (N_33746,N_31888,N_30935);
xnor U33747 (N_33747,N_31318,N_32231);
nand U33748 (N_33748,N_31715,N_32206);
xor U33749 (N_33749,N_32281,N_32097);
or U33750 (N_33750,N_30605,N_30805);
xnor U33751 (N_33751,N_31652,N_30551);
xnor U33752 (N_33752,N_30388,N_30286);
or U33753 (N_33753,N_30705,N_31237);
or U33754 (N_33754,N_30559,N_32273);
and U33755 (N_33755,N_32329,N_30312);
or U33756 (N_33756,N_30450,N_31797);
nor U33757 (N_33757,N_30913,N_30889);
and U33758 (N_33758,N_31691,N_32471);
nand U33759 (N_33759,N_31086,N_31599);
and U33760 (N_33760,N_31201,N_31125);
or U33761 (N_33761,N_31150,N_31859);
and U33762 (N_33762,N_30639,N_30473);
xnor U33763 (N_33763,N_30899,N_31181);
xnor U33764 (N_33764,N_32034,N_30345);
xnor U33765 (N_33765,N_31106,N_31743);
nor U33766 (N_33766,N_30487,N_30653);
and U33767 (N_33767,N_31778,N_32395);
xor U33768 (N_33768,N_31667,N_31391);
nand U33769 (N_33769,N_31707,N_30056);
nand U33770 (N_33770,N_31864,N_31967);
or U33771 (N_33771,N_32499,N_31250);
xnor U33772 (N_33772,N_31625,N_32435);
nor U33773 (N_33773,N_31295,N_31755);
nor U33774 (N_33774,N_30532,N_30450);
xnor U33775 (N_33775,N_32173,N_30734);
xnor U33776 (N_33776,N_31945,N_31863);
or U33777 (N_33777,N_30574,N_31349);
nor U33778 (N_33778,N_31433,N_30371);
nand U33779 (N_33779,N_32496,N_30534);
nand U33780 (N_33780,N_32264,N_30793);
and U33781 (N_33781,N_30150,N_31091);
xnor U33782 (N_33782,N_31670,N_30247);
xnor U33783 (N_33783,N_31450,N_30003);
and U33784 (N_33784,N_30112,N_31498);
or U33785 (N_33785,N_30967,N_30800);
or U33786 (N_33786,N_31675,N_30936);
and U33787 (N_33787,N_32292,N_32383);
nor U33788 (N_33788,N_32498,N_30244);
and U33789 (N_33789,N_31074,N_30220);
or U33790 (N_33790,N_32022,N_30067);
nand U33791 (N_33791,N_31547,N_30821);
nand U33792 (N_33792,N_31425,N_30880);
xnor U33793 (N_33793,N_31786,N_31341);
xnor U33794 (N_33794,N_32435,N_32172);
nand U33795 (N_33795,N_31068,N_31314);
nor U33796 (N_33796,N_30423,N_31918);
or U33797 (N_33797,N_30578,N_31868);
nand U33798 (N_33798,N_30847,N_30251);
nand U33799 (N_33799,N_31216,N_32098);
nand U33800 (N_33800,N_31599,N_30004);
xnor U33801 (N_33801,N_30104,N_32325);
and U33802 (N_33802,N_31400,N_31825);
xnor U33803 (N_33803,N_32444,N_31379);
xor U33804 (N_33804,N_30400,N_30893);
nand U33805 (N_33805,N_31745,N_32239);
xor U33806 (N_33806,N_31260,N_30522);
nor U33807 (N_33807,N_32138,N_32465);
xnor U33808 (N_33808,N_32366,N_31681);
xor U33809 (N_33809,N_30963,N_32205);
or U33810 (N_33810,N_31715,N_31177);
nand U33811 (N_33811,N_32018,N_31192);
nand U33812 (N_33812,N_30100,N_32298);
and U33813 (N_33813,N_30938,N_32438);
nor U33814 (N_33814,N_30006,N_30493);
nor U33815 (N_33815,N_31064,N_31700);
nor U33816 (N_33816,N_30855,N_31176);
nand U33817 (N_33817,N_31272,N_31646);
xnor U33818 (N_33818,N_31655,N_30553);
xor U33819 (N_33819,N_30252,N_30554);
xnor U33820 (N_33820,N_30720,N_31758);
nor U33821 (N_33821,N_30025,N_32086);
nand U33822 (N_33822,N_32222,N_30317);
and U33823 (N_33823,N_30624,N_31316);
xnor U33824 (N_33824,N_31088,N_31749);
nand U33825 (N_33825,N_32032,N_31608);
or U33826 (N_33826,N_31637,N_30235);
xnor U33827 (N_33827,N_30178,N_31090);
or U33828 (N_33828,N_30016,N_30411);
and U33829 (N_33829,N_31187,N_30127);
nor U33830 (N_33830,N_32225,N_31175);
nand U33831 (N_33831,N_30977,N_30361);
and U33832 (N_33832,N_31912,N_31612);
nand U33833 (N_33833,N_30417,N_31829);
nor U33834 (N_33834,N_32116,N_32130);
and U33835 (N_33835,N_32307,N_31589);
nand U33836 (N_33836,N_32275,N_30515);
or U33837 (N_33837,N_31670,N_30565);
and U33838 (N_33838,N_31346,N_31081);
and U33839 (N_33839,N_30414,N_31562);
nand U33840 (N_33840,N_32238,N_30486);
nand U33841 (N_33841,N_30882,N_31566);
and U33842 (N_33842,N_31013,N_30510);
and U33843 (N_33843,N_30394,N_31044);
nor U33844 (N_33844,N_31395,N_31454);
xor U33845 (N_33845,N_31943,N_30656);
and U33846 (N_33846,N_31139,N_30621);
and U33847 (N_33847,N_31535,N_30854);
nand U33848 (N_33848,N_30179,N_32391);
nand U33849 (N_33849,N_30319,N_31962);
nand U33850 (N_33850,N_31479,N_31777);
or U33851 (N_33851,N_30956,N_30830);
nand U33852 (N_33852,N_30544,N_32267);
nand U33853 (N_33853,N_32116,N_32158);
or U33854 (N_33854,N_32475,N_31092);
or U33855 (N_33855,N_31570,N_30055);
or U33856 (N_33856,N_31946,N_31915);
nor U33857 (N_33857,N_30043,N_31445);
nor U33858 (N_33858,N_31102,N_32269);
nand U33859 (N_33859,N_31250,N_30696);
or U33860 (N_33860,N_32027,N_31927);
or U33861 (N_33861,N_31346,N_31861);
and U33862 (N_33862,N_32358,N_30004);
and U33863 (N_33863,N_32264,N_30492);
and U33864 (N_33864,N_32336,N_31402);
xor U33865 (N_33865,N_30714,N_31179);
nand U33866 (N_33866,N_30376,N_31994);
xnor U33867 (N_33867,N_30326,N_32186);
and U33868 (N_33868,N_30769,N_31267);
nand U33869 (N_33869,N_30240,N_32020);
and U33870 (N_33870,N_31095,N_31444);
xnor U33871 (N_33871,N_30653,N_32173);
and U33872 (N_33872,N_31819,N_31265);
nand U33873 (N_33873,N_30500,N_32311);
or U33874 (N_33874,N_30904,N_31303);
nor U33875 (N_33875,N_32170,N_30572);
xnor U33876 (N_33876,N_30026,N_32201);
nand U33877 (N_33877,N_32113,N_31918);
nor U33878 (N_33878,N_32263,N_31684);
xor U33879 (N_33879,N_31406,N_30964);
or U33880 (N_33880,N_30251,N_30289);
and U33881 (N_33881,N_31598,N_30799);
xor U33882 (N_33882,N_31330,N_30345);
and U33883 (N_33883,N_30815,N_31837);
or U33884 (N_33884,N_31468,N_31889);
or U33885 (N_33885,N_30546,N_30752);
nor U33886 (N_33886,N_30594,N_31102);
nor U33887 (N_33887,N_30806,N_30522);
nand U33888 (N_33888,N_31781,N_31497);
or U33889 (N_33889,N_31842,N_32114);
and U33890 (N_33890,N_31518,N_30600);
and U33891 (N_33891,N_30784,N_32405);
nor U33892 (N_33892,N_30479,N_30185);
or U33893 (N_33893,N_31011,N_32076);
nand U33894 (N_33894,N_31995,N_32107);
and U33895 (N_33895,N_31395,N_31320);
xor U33896 (N_33896,N_30498,N_30712);
xnor U33897 (N_33897,N_30581,N_31541);
nor U33898 (N_33898,N_30038,N_31278);
or U33899 (N_33899,N_32252,N_31231);
and U33900 (N_33900,N_31050,N_30575);
and U33901 (N_33901,N_32414,N_30927);
and U33902 (N_33902,N_31203,N_31800);
nand U33903 (N_33903,N_32262,N_30414);
nor U33904 (N_33904,N_30040,N_31197);
and U33905 (N_33905,N_30993,N_32366);
and U33906 (N_33906,N_31343,N_31557);
nand U33907 (N_33907,N_30065,N_32205);
nand U33908 (N_33908,N_32211,N_31614);
nand U33909 (N_33909,N_31659,N_31010);
or U33910 (N_33910,N_31795,N_31646);
or U33911 (N_33911,N_32018,N_32318);
nand U33912 (N_33912,N_31665,N_30045);
xor U33913 (N_33913,N_30698,N_32018);
and U33914 (N_33914,N_32339,N_31747);
or U33915 (N_33915,N_30526,N_31047);
nor U33916 (N_33916,N_30623,N_32134);
xnor U33917 (N_33917,N_30060,N_31965);
and U33918 (N_33918,N_31965,N_32010);
or U33919 (N_33919,N_30706,N_31741);
xnor U33920 (N_33920,N_31517,N_30097);
and U33921 (N_33921,N_31563,N_30819);
or U33922 (N_33922,N_32175,N_31522);
nand U33923 (N_33923,N_32487,N_31102);
xnor U33924 (N_33924,N_32453,N_31227);
xnor U33925 (N_33925,N_31616,N_30999);
xnor U33926 (N_33926,N_30801,N_31950);
xor U33927 (N_33927,N_31906,N_30381);
nand U33928 (N_33928,N_30497,N_30199);
xnor U33929 (N_33929,N_31842,N_32433);
nor U33930 (N_33930,N_30484,N_32433);
nand U33931 (N_33931,N_31332,N_31861);
nand U33932 (N_33932,N_32032,N_30124);
or U33933 (N_33933,N_32116,N_32234);
nand U33934 (N_33934,N_30774,N_32445);
nand U33935 (N_33935,N_30900,N_30988);
or U33936 (N_33936,N_31686,N_31192);
and U33937 (N_33937,N_31520,N_31712);
or U33938 (N_33938,N_31467,N_31996);
and U33939 (N_33939,N_31927,N_30009);
nand U33940 (N_33940,N_30459,N_30451);
or U33941 (N_33941,N_31236,N_31014);
nand U33942 (N_33942,N_32050,N_30872);
nand U33943 (N_33943,N_31736,N_31872);
and U33944 (N_33944,N_31619,N_31989);
nor U33945 (N_33945,N_31321,N_32145);
and U33946 (N_33946,N_30723,N_31664);
nand U33947 (N_33947,N_30633,N_30597);
nor U33948 (N_33948,N_30558,N_30158);
or U33949 (N_33949,N_30300,N_30008);
or U33950 (N_33950,N_30062,N_30082);
xnor U33951 (N_33951,N_32350,N_32055);
and U33952 (N_33952,N_31279,N_32168);
nand U33953 (N_33953,N_31800,N_30922);
or U33954 (N_33954,N_31255,N_30662);
or U33955 (N_33955,N_31954,N_31792);
and U33956 (N_33956,N_30636,N_30928);
and U33957 (N_33957,N_31617,N_32102);
nand U33958 (N_33958,N_30185,N_31091);
and U33959 (N_33959,N_32044,N_31863);
and U33960 (N_33960,N_31728,N_31962);
and U33961 (N_33961,N_30175,N_31395);
and U33962 (N_33962,N_30021,N_30390);
and U33963 (N_33963,N_31944,N_31980);
xnor U33964 (N_33964,N_31207,N_30978);
xnor U33965 (N_33965,N_32296,N_32376);
or U33966 (N_33966,N_31699,N_31912);
xnor U33967 (N_33967,N_31586,N_31719);
xor U33968 (N_33968,N_31130,N_31303);
nand U33969 (N_33969,N_31308,N_31413);
nand U33970 (N_33970,N_32173,N_32039);
nand U33971 (N_33971,N_32305,N_30050);
xor U33972 (N_33972,N_31132,N_32233);
and U33973 (N_33973,N_31495,N_31258);
nor U33974 (N_33974,N_30305,N_31382);
or U33975 (N_33975,N_30015,N_30232);
xnor U33976 (N_33976,N_30496,N_30407);
nor U33977 (N_33977,N_30824,N_31352);
and U33978 (N_33978,N_32429,N_31932);
xor U33979 (N_33979,N_31735,N_31777);
nand U33980 (N_33980,N_31116,N_30811);
nand U33981 (N_33981,N_31629,N_30705);
nand U33982 (N_33982,N_31822,N_31542);
nand U33983 (N_33983,N_30813,N_31431);
and U33984 (N_33984,N_30447,N_31684);
nand U33985 (N_33985,N_31506,N_31022);
xnor U33986 (N_33986,N_31824,N_30033);
and U33987 (N_33987,N_31426,N_30625);
xnor U33988 (N_33988,N_30131,N_32180);
and U33989 (N_33989,N_30736,N_30689);
nand U33990 (N_33990,N_31140,N_31217);
xor U33991 (N_33991,N_32030,N_32362);
or U33992 (N_33992,N_30849,N_30554);
and U33993 (N_33993,N_31735,N_30476);
nor U33994 (N_33994,N_30388,N_30857);
nand U33995 (N_33995,N_31548,N_31414);
nand U33996 (N_33996,N_32310,N_32109);
and U33997 (N_33997,N_31845,N_30176);
nor U33998 (N_33998,N_31038,N_32021);
nor U33999 (N_33999,N_30825,N_32149);
xnor U34000 (N_34000,N_30902,N_31378);
or U34001 (N_34001,N_31228,N_30756);
or U34002 (N_34002,N_31369,N_30317);
or U34003 (N_34003,N_30832,N_30524);
nor U34004 (N_34004,N_31826,N_31166);
nand U34005 (N_34005,N_30126,N_30909);
nor U34006 (N_34006,N_31644,N_31437);
nor U34007 (N_34007,N_31977,N_31025);
xnor U34008 (N_34008,N_30539,N_30666);
nand U34009 (N_34009,N_30632,N_32434);
nor U34010 (N_34010,N_30329,N_30963);
nand U34011 (N_34011,N_32138,N_31725);
xor U34012 (N_34012,N_30124,N_31137);
xor U34013 (N_34013,N_31553,N_31678);
or U34014 (N_34014,N_32337,N_30946);
nand U34015 (N_34015,N_30704,N_31900);
nand U34016 (N_34016,N_31461,N_30179);
or U34017 (N_34017,N_30603,N_30764);
nand U34018 (N_34018,N_31405,N_30815);
and U34019 (N_34019,N_30927,N_30735);
xor U34020 (N_34020,N_31989,N_31520);
and U34021 (N_34021,N_32286,N_30461);
or U34022 (N_34022,N_30774,N_30891);
xnor U34023 (N_34023,N_31139,N_32218);
xnor U34024 (N_34024,N_30160,N_31561);
xor U34025 (N_34025,N_31674,N_30253);
xnor U34026 (N_34026,N_32246,N_31374);
nand U34027 (N_34027,N_31415,N_32296);
xor U34028 (N_34028,N_30248,N_32113);
and U34029 (N_34029,N_30584,N_31411);
nor U34030 (N_34030,N_32302,N_30963);
xnor U34031 (N_34031,N_32068,N_30937);
nand U34032 (N_34032,N_32263,N_31553);
xnor U34033 (N_34033,N_31687,N_30159);
and U34034 (N_34034,N_32008,N_31869);
nand U34035 (N_34035,N_31481,N_31083);
xnor U34036 (N_34036,N_31991,N_31608);
xnor U34037 (N_34037,N_30218,N_31662);
nand U34038 (N_34038,N_32396,N_30284);
or U34039 (N_34039,N_31588,N_31708);
or U34040 (N_34040,N_32200,N_31241);
or U34041 (N_34041,N_31780,N_30806);
or U34042 (N_34042,N_30100,N_31655);
or U34043 (N_34043,N_31355,N_31050);
and U34044 (N_34044,N_30758,N_30636);
nor U34045 (N_34045,N_30992,N_31670);
nand U34046 (N_34046,N_32079,N_31196);
and U34047 (N_34047,N_30775,N_30764);
or U34048 (N_34048,N_30195,N_32095);
xnor U34049 (N_34049,N_30192,N_31747);
xnor U34050 (N_34050,N_32022,N_31578);
nand U34051 (N_34051,N_30980,N_31985);
or U34052 (N_34052,N_30436,N_30534);
nor U34053 (N_34053,N_30449,N_31217);
nand U34054 (N_34054,N_32167,N_32105);
or U34055 (N_34055,N_31231,N_31985);
xor U34056 (N_34056,N_31419,N_31645);
or U34057 (N_34057,N_30568,N_32447);
and U34058 (N_34058,N_30634,N_30994);
xor U34059 (N_34059,N_32326,N_31803);
nand U34060 (N_34060,N_30815,N_30610);
nand U34061 (N_34061,N_30512,N_30373);
xor U34062 (N_34062,N_32264,N_30083);
xnor U34063 (N_34063,N_30881,N_32357);
and U34064 (N_34064,N_31202,N_31117);
and U34065 (N_34065,N_31683,N_32381);
xor U34066 (N_34066,N_31634,N_31545);
nor U34067 (N_34067,N_30282,N_32301);
and U34068 (N_34068,N_31390,N_31343);
or U34069 (N_34069,N_30431,N_31015);
nand U34070 (N_34070,N_30571,N_31675);
xor U34071 (N_34071,N_31331,N_31381);
or U34072 (N_34072,N_30045,N_31048);
nor U34073 (N_34073,N_30543,N_31869);
xor U34074 (N_34074,N_30605,N_31683);
xor U34075 (N_34075,N_32104,N_30178);
nor U34076 (N_34076,N_31763,N_30202);
xor U34077 (N_34077,N_31644,N_31024);
and U34078 (N_34078,N_30700,N_30514);
or U34079 (N_34079,N_31124,N_31189);
and U34080 (N_34080,N_31273,N_30073);
nand U34081 (N_34081,N_30435,N_31857);
or U34082 (N_34082,N_31882,N_31396);
and U34083 (N_34083,N_30422,N_30942);
and U34084 (N_34084,N_31877,N_31891);
nand U34085 (N_34085,N_31166,N_32240);
nor U34086 (N_34086,N_30437,N_30398);
or U34087 (N_34087,N_30571,N_31079);
xor U34088 (N_34088,N_30863,N_32492);
and U34089 (N_34089,N_30312,N_32018);
nand U34090 (N_34090,N_30104,N_31698);
and U34091 (N_34091,N_30567,N_30245);
nand U34092 (N_34092,N_30708,N_30187);
nand U34093 (N_34093,N_30103,N_31335);
nand U34094 (N_34094,N_30486,N_30517);
nand U34095 (N_34095,N_30138,N_30881);
xnor U34096 (N_34096,N_32087,N_30944);
xnor U34097 (N_34097,N_30039,N_31417);
xnor U34098 (N_34098,N_31093,N_30718);
xor U34099 (N_34099,N_30185,N_31904);
and U34100 (N_34100,N_31741,N_32225);
and U34101 (N_34101,N_32149,N_31604);
and U34102 (N_34102,N_30667,N_31827);
nor U34103 (N_34103,N_31072,N_30152);
nand U34104 (N_34104,N_30760,N_31977);
nor U34105 (N_34105,N_31155,N_30306);
xnor U34106 (N_34106,N_30919,N_32389);
or U34107 (N_34107,N_31138,N_31091);
or U34108 (N_34108,N_32436,N_31734);
nand U34109 (N_34109,N_30537,N_30497);
nand U34110 (N_34110,N_30123,N_32286);
nor U34111 (N_34111,N_30757,N_30210);
and U34112 (N_34112,N_30825,N_30861);
or U34113 (N_34113,N_31451,N_30557);
and U34114 (N_34114,N_30347,N_32396);
xnor U34115 (N_34115,N_31942,N_31403);
xnor U34116 (N_34116,N_30862,N_30980);
or U34117 (N_34117,N_31179,N_30496);
nor U34118 (N_34118,N_30733,N_31759);
or U34119 (N_34119,N_32412,N_30594);
xnor U34120 (N_34120,N_32082,N_31788);
and U34121 (N_34121,N_31891,N_31234);
or U34122 (N_34122,N_30977,N_32111);
xor U34123 (N_34123,N_31898,N_30446);
and U34124 (N_34124,N_31227,N_30941);
nand U34125 (N_34125,N_31642,N_31324);
nor U34126 (N_34126,N_30722,N_32358);
and U34127 (N_34127,N_32449,N_32263);
nand U34128 (N_34128,N_32237,N_30931);
or U34129 (N_34129,N_30057,N_31585);
nand U34130 (N_34130,N_31134,N_32433);
nand U34131 (N_34131,N_30436,N_30317);
xor U34132 (N_34132,N_32139,N_32380);
xnor U34133 (N_34133,N_31287,N_30059);
nand U34134 (N_34134,N_32487,N_30550);
nand U34135 (N_34135,N_30433,N_31949);
nand U34136 (N_34136,N_31568,N_30861);
nand U34137 (N_34137,N_32153,N_30552);
xor U34138 (N_34138,N_31496,N_30479);
nor U34139 (N_34139,N_30695,N_30488);
xor U34140 (N_34140,N_32368,N_31820);
nor U34141 (N_34141,N_32321,N_30109);
xor U34142 (N_34142,N_30013,N_31495);
and U34143 (N_34143,N_30940,N_30306);
nor U34144 (N_34144,N_30340,N_30121);
nor U34145 (N_34145,N_31895,N_31325);
nand U34146 (N_34146,N_31644,N_31907);
nand U34147 (N_34147,N_30968,N_31745);
or U34148 (N_34148,N_31094,N_30139);
or U34149 (N_34149,N_30549,N_31207);
nand U34150 (N_34150,N_30573,N_31363);
nand U34151 (N_34151,N_30659,N_30189);
or U34152 (N_34152,N_30015,N_31327);
xnor U34153 (N_34153,N_31213,N_30581);
and U34154 (N_34154,N_31155,N_32498);
xor U34155 (N_34155,N_30271,N_32217);
xor U34156 (N_34156,N_31574,N_30419);
or U34157 (N_34157,N_30454,N_31322);
or U34158 (N_34158,N_30630,N_31655);
and U34159 (N_34159,N_31167,N_30627);
or U34160 (N_34160,N_32010,N_30872);
nand U34161 (N_34161,N_30408,N_32432);
and U34162 (N_34162,N_31030,N_30113);
nand U34163 (N_34163,N_32355,N_30372);
or U34164 (N_34164,N_30547,N_30448);
xnor U34165 (N_34165,N_32367,N_30179);
nor U34166 (N_34166,N_30835,N_30669);
nor U34167 (N_34167,N_30057,N_30091);
and U34168 (N_34168,N_31453,N_31801);
xor U34169 (N_34169,N_30845,N_32430);
or U34170 (N_34170,N_31825,N_32341);
nand U34171 (N_34171,N_30527,N_32329);
xnor U34172 (N_34172,N_32198,N_31485);
and U34173 (N_34173,N_32342,N_32379);
nor U34174 (N_34174,N_30211,N_31798);
xnor U34175 (N_34175,N_32278,N_32178);
nand U34176 (N_34176,N_30454,N_31303);
xnor U34177 (N_34177,N_31449,N_32028);
nand U34178 (N_34178,N_30888,N_31008);
xnor U34179 (N_34179,N_30041,N_30760);
nand U34180 (N_34180,N_31186,N_32262);
and U34181 (N_34181,N_31478,N_30938);
nor U34182 (N_34182,N_32015,N_31691);
nand U34183 (N_34183,N_30315,N_30010);
nand U34184 (N_34184,N_32346,N_30456);
or U34185 (N_34185,N_31150,N_31052);
xor U34186 (N_34186,N_32344,N_30123);
nand U34187 (N_34187,N_30548,N_31218);
or U34188 (N_34188,N_32002,N_32375);
xor U34189 (N_34189,N_30781,N_30384);
or U34190 (N_34190,N_30397,N_31397);
or U34191 (N_34191,N_32167,N_30669);
xor U34192 (N_34192,N_30022,N_30990);
nand U34193 (N_34193,N_32389,N_31755);
nor U34194 (N_34194,N_31289,N_32234);
nor U34195 (N_34195,N_31579,N_30641);
nor U34196 (N_34196,N_31940,N_31730);
nand U34197 (N_34197,N_32044,N_31670);
and U34198 (N_34198,N_31757,N_30435);
nor U34199 (N_34199,N_30414,N_31051);
xnor U34200 (N_34200,N_31534,N_30755);
and U34201 (N_34201,N_31226,N_30176);
nand U34202 (N_34202,N_31809,N_32023);
or U34203 (N_34203,N_32051,N_31010);
or U34204 (N_34204,N_31939,N_31247);
xnor U34205 (N_34205,N_31178,N_30387);
and U34206 (N_34206,N_30276,N_32466);
nand U34207 (N_34207,N_32461,N_31839);
nand U34208 (N_34208,N_32020,N_32320);
or U34209 (N_34209,N_32492,N_32128);
xor U34210 (N_34210,N_32108,N_30565);
nor U34211 (N_34211,N_30582,N_30904);
or U34212 (N_34212,N_30902,N_32404);
and U34213 (N_34213,N_32323,N_30743);
and U34214 (N_34214,N_31212,N_31189);
nand U34215 (N_34215,N_31775,N_32264);
or U34216 (N_34216,N_30294,N_31447);
and U34217 (N_34217,N_31540,N_31876);
xor U34218 (N_34218,N_32060,N_31917);
or U34219 (N_34219,N_32180,N_32085);
or U34220 (N_34220,N_30022,N_31552);
xnor U34221 (N_34221,N_30844,N_30754);
xnor U34222 (N_34222,N_32422,N_30958);
or U34223 (N_34223,N_32248,N_31673);
nand U34224 (N_34224,N_30977,N_31099);
and U34225 (N_34225,N_32447,N_31895);
or U34226 (N_34226,N_30950,N_30177);
and U34227 (N_34227,N_32334,N_30241);
xor U34228 (N_34228,N_31198,N_32009);
and U34229 (N_34229,N_30580,N_30585);
nor U34230 (N_34230,N_32262,N_31801);
nor U34231 (N_34231,N_32369,N_31749);
and U34232 (N_34232,N_30082,N_31919);
nor U34233 (N_34233,N_30216,N_30986);
xor U34234 (N_34234,N_31422,N_31521);
nand U34235 (N_34235,N_30129,N_31500);
xor U34236 (N_34236,N_31172,N_30523);
or U34237 (N_34237,N_32347,N_30688);
nand U34238 (N_34238,N_30716,N_31675);
nor U34239 (N_34239,N_30362,N_31319);
xor U34240 (N_34240,N_30842,N_31664);
xnor U34241 (N_34241,N_31135,N_30687);
xor U34242 (N_34242,N_30106,N_30637);
or U34243 (N_34243,N_30361,N_32460);
and U34244 (N_34244,N_32284,N_31378);
or U34245 (N_34245,N_31006,N_32382);
nand U34246 (N_34246,N_31319,N_30839);
xor U34247 (N_34247,N_30926,N_30163);
nand U34248 (N_34248,N_31616,N_30824);
nor U34249 (N_34249,N_30313,N_30789);
nor U34250 (N_34250,N_31251,N_31613);
nor U34251 (N_34251,N_32241,N_30951);
xor U34252 (N_34252,N_31423,N_30926);
xor U34253 (N_34253,N_32212,N_30525);
nor U34254 (N_34254,N_32432,N_30997);
or U34255 (N_34255,N_32252,N_30614);
xnor U34256 (N_34256,N_31907,N_30339);
xnor U34257 (N_34257,N_31062,N_30119);
and U34258 (N_34258,N_32022,N_30539);
or U34259 (N_34259,N_30658,N_31118);
and U34260 (N_34260,N_31686,N_30367);
xor U34261 (N_34261,N_31494,N_31182);
nand U34262 (N_34262,N_31273,N_32409);
and U34263 (N_34263,N_31880,N_31381);
or U34264 (N_34264,N_32269,N_32121);
or U34265 (N_34265,N_31305,N_31671);
and U34266 (N_34266,N_30472,N_31798);
nand U34267 (N_34267,N_32309,N_31311);
xor U34268 (N_34268,N_30564,N_31275);
and U34269 (N_34269,N_31275,N_31827);
nand U34270 (N_34270,N_30560,N_32323);
or U34271 (N_34271,N_31217,N_30969);
and U34272 (N_34272,N_31575,N_30868);
xor U34273 (N_34273,N_31374,N_30919);
and U34274 (N_34274,N_32026,N_31020);
or U34275 (N_34275,N_32289,N_32430);
or U34276 (N_34276,N_31067,N_31941);
nor U34277 (N_34277,N_30684,N_31661);
nand U34278 (N_34278,N_31263,N_30037);
nand U34279 (N_34279,N_31977,N_32372);
nor U34280 (N_34280,N_30623,N_31356);
nand U34281 (N_34281,N_31307,N_31629);
nand U34282 (N_34282,N_30748,N_30181);
nand U34283 (N_34283,N_32064,N_30234);
nand U34284 (N_34284,N_31625,N_32441);
nor U34285 (N_34285,N_30324,N_30994);
or U34286 (N_34286,N_31660,N_30295);
or U34287 (N_34287,N_30311,N_32466);
nand U34288 (N_34288,N_32325,N_31071);
xor U34289 (N_34289,N_31854,N_32430);
or U34290 (N_34290,N_30719,N_31122);
xor U34291 (N_34291,N_31260,N_30880);
nand U34292 (N_34292,N_32317,N_32060);
nand U34293 (N_34293,N_31370,N_30753);
xnor U34294 (N_34294,N_30426,N_31964);
xor U34295 (N_34295,N_32240,N_31075);
xnor U34296 (N_34296,N_30776,N_31201);
nor U34297 (N_34297,N_31693,N_31929);
and U34298 (N_34298,N_31593,N_32175);
xnor U34299 (N_34299,N_31382,N_31314);
nand U34300 (N_34300,N_31638,N_32364);
and U34301 (N_34301,N_31134,N_32445);
and U34302 (N_34302,N_32204,N_31659);
xnor U34303 (N_34303,N_31580,N_31537);
and U34304 (N_34304,N_32345,N_30989);
nand U34305 (N_34305,N_31165,N_30207);
nor U34306 (N_34306,N_30439,N_30969);
nor U34307 (N_34307,N_31964,N_31205);
nand U34308 (N_34308,N_30412,N_30233);
or U34309 (N_34309,N_31688,N_32472);
xor U34310 (N_34310,N_31186,N_32040);
nand U34311 (N_34311,N_31921,N_30420);
or U34312 (N_34312,N_30282,N_32348);
nand U34313 (N_34313,N_30090,N_31677);
xnor U34314 (N_34314,N_30381,N_31545);
xnor U34315 (N_34315,N_30913,N_31336);
and U34316 (N_34316,N_30201,N_30627);
nand U34317 (N_34317,N_31692,N_31124);
nor U34318 (N_34318,N_30456,N_30788);
nor U34319 (N_34319,N_31079,N_31126);
and U34320 (N_34320,N_32137,N_30147);
xor U34321 (N_34321,N_32247,N_31655);
or U34322 (N_34322,N_31905,N_31059);
nand U34323 (N_34323,N_32347,N_31917);
or U34324 (N_34324,N_30657,N_31998);
xnor U34325 (N_34325,N_30698,N_32069);
xnor U34326 (N_34326,N_31200,N_31896);
xor U34327 (N_34327,N_30963,N_30298);
nand U34328 (N_34328,N_30517,N_30903);
xor U34329 (N_34329,N_31521,N_31779);
and U34330 (N_34330,N_31623,N_32497);
and U34331 (N_34331,N_30937,N_30412);
or U34332 (N_34332,N_32204,N_31825);
nand U34333 (N_34333,N_30262,N_30196);
and U34334 (N_34334,N_32242,N_31810);
and U34335 (N_34335,N_31502,N_32428);
nor U34336 (N_34336,N_31856,N_31464);
and U34337 (N_34337,N_30206,N_30391);
and U34338 (N_34338,N_30920,N_30736);
nor U34339 (N_34339,N_30179,N_30883);
and U34340 (N_34340,N_32164,N_30125);
nand U34341 (N_34341,N_32328,N_32214);
nand U34342 (N_34342,N_30475,N_31396);
and U34343 (N_34343,N_32212,N_30458);
nor U34344 (N_34344,N_30323,N_32323);
nand U34345 (N_34345,N_32375,N_31306);
nand U34346 (N_34346,N_31567,N_31447);
nand U34347 (N_34347,N_30592,N_30816);
xnor U34348 (N_34348,N_31668,N_32063);
or U34349 (N_34349,N_30671,N_30311);
nand U34350 (N_34350,N_31966,N_32377);
nand U34351 (N_34351,N_32330,N_30424);
nor U34352 (N_34352,N_30167,N_31207);
nand U34353 (N_34353,N_31793,N_32399);
nand U34354 (N_34354,N_32473,N_31200);
xor U34355 (N_34355,N_30047,N_30045);
nand U34356 (N_34356,N_31308,N_31682);
or U34357 (N_34357,N_31477,N_32177);
and U34358 (N_34358,N_30932,N_30513);
xnor U34359 (N_34359,N_31285,N_31355);
nand U34360 (N_34360,N_32333,N_31147);
nor U34361 (N_34361,N_30792,N_32434);
and U34362 (N_34362,N_31827,N_31034);
nand U34363 (N_34363,N_31907,N_30897);
xnor U34364 (N_34364,N_31120,N_31677);
and U34365 (N_34365,N_30569,N_31407);
xnor U34366 (N_34366,N_32089,N_31484);
nor U34367 (N_34367,N_30428,N_31301);
xor U34368 (N_34368,N_30263,N_30337);
or U34369 (N_34369,N_30005,N_31152);
and U34370 (N_34370,N_30909,N_30124);
and U34371 (N_34371,N_30886,N_30056);
or U34372 (N_34372,N_30675,N_31777);
nand U34373 (N_34373,N_31100,N_30075);
and U34374 (N_34374,N_30939,N_30578);
or U34375 (N_34375,N_31612,N_30777);
or U34376 (N_34376,N_30732,N_32182);
nand U34377 (N_34377,N_30608,N_31271);
and U34378 (N_34378,N_30085,N_31779);
xnor U34379 (N_34379,N_31423,N_31403);
and U34380 (N_34380,N_31922,N_31966);
and U34381 (N_34381,N_30418,N_30174);
xor U34382 (N_34382,N_30769,N_31271);
or U34383 (N_34383,N_30989,N_31578);
or U34384 (N_34384,N_30112,N_30650);
nor U34385 (N_34385,N_31407,N_30989);
or U34386 (N_34386,N_31944,N_31926);
or U34387 (N_34387,N_31426,N_32251);
nand U34388 (N_34388,N_31433,N_31080);
or U34389 (N_34389,N_31242,N_31152);
nand U34390 (N_34390,N_30125,N_32040);
xor U34391 (N_34391,N_31768,N_31964);
nor U34392 (N_34392,N_31260,N_31061);
nand U34393 (N_34393,N_32493,N_30233);
nor U34394 (N_34394,N_30548,N_31921);
or U34395 (N_34395,N_30994,N_30570);
xor U34396 (N_34396,N_32222,N_31912);
nand U34397 (N_34397,N_30964,N_32488);
xor U34398 (N_34398,N_31920,N_30369);
and U34399 (N_34399,N_32004,N_30020);
or U34400 (N_34400,N_31425,N_31666);
xnor U34401 (N_34401,N_30981,N_31247);
nand U34402 (N_34402,N_30371,N_31021);
or U34403 (N_34403,N_30488,N_31744);
or U34404 (N_34404,N_31068,N_31051);
nand U34405 (N_34405,N_30330,N_31892);
and U34406 (N_34406,N_31349,N_31262);
nor U34407 (N_34407,N_31683,N_30523);
nor U34408 (N_34408,N_30537,N_31551);
xnor U34409 (N_34409,N_32312,N_31347);
nor U34410 (N_34410,N_31941,N_31358);
xnor U34411 (N_34411,N_31803,N_31031);
and U34412 (N_34412,N_31136,N_30859);
and U34413 (N_34413,N_30450,N_31227);
nor U34414 (N_34414,N_31346,N_31151);
or U34415 (N_34415,N_32291,N_31609);
nor U34416 (N_34416,N_31622,N_31501);
and U34417 (N_34417,N_30230,N_30797);
nand U34418 (N_34418,N_30412,N_31693);
nand U34419 (N_34419,N_32310,N_30497);
nor U34420 (N_34420,N_31172,N_31131);
or U34421 (N_34421,N_32423,N_31979);
and U34422 (N_34422,N_31147,N_31797);
nor U34423 (N_34423,N_30241,N_30911);
or U34424 (N_34424,N_31174,N_31652);
xor U34425 (N_34425,N_31958,N_30724);
nand U34426 (N_34426,N_32337,N_31316);
nor U34427 (N_34427,N_30778,N_31405);
and U34428 (N_34428,N_31413,N_30108);
xor U34429 (N_34429,N_32083,N_31565);
xor U34430 (N_34430,N_30974,N_30955);
xor U34431 (N_34431,N_30925,N_30753);
nand U34432 (N_34432,N_32211,N_30588);
or U34433 (N_34433,N_31638,N_30466);
nor U34434 (N_34434,N_31158,N_31398);
nor U34435 (N_34435,N_32260,N_32487);
nor U34436 (N_34436,N_30016,N_31738);
nand U34437 (N_34437,N_32317,N_30907);
and U34438 (N_34438,N_31726,N_30311);
nand U34439 (N_34439,N_31763,N_31814);
and U34440 (N_34440,N_31410,N_30871);
or U34441 (N_34441,N_30532,N_32315);
and U34442 (N_34442,N_30194,N_30004);
nor U34443 (N_34443,N_30898,N_32357);
xor U34444 (N_34444,N_30044,N_31266);
and U34445 (N_34445,N_30144,N_31174);
nor U34446 (N_34446,N_30751,N_30857);
xor U34447 (N_34447,N_30826,N_30104);
xor U34448 (N_34448,N_30014,N_31956);
xor U34449 (N_34449,N_30488,N_31379);
nand U34450 (N_34450,N_30433,N_30079);
or U34451 (N_34451,N_31188,N_32457);
and U34452 (N_34452,N_31378,N_32267);
xor U34453 (N_34453,N_32073,N_31800);
or U34454 (N_34454,N_30070,N_30280);
nor U34455 (N_34455,N_30116,N_31759);
xor U34456 (N_34456,N_31202,N_31363);
nor U34457 (N_34457,N_31398,N_32313);
nor U34458 (N_34458,N_30340,N_31796);
nor U34459 (N_34459,N_31159,N_31864);
nor U34460 (N_34460,N_31119,N_30334);
nand U34461 (N_34461,N_31722,N_31691);
and U34462 (N_34462,N_31343,N_30693);
xnor U34463 (N_34463,N_31351,N_30925);
nor U34464 (N_34464,N_30698,N_31149);
and U34465 (N_34465,N_31707,N_31913);
xor U34466 (N_34466,N_32242,N_30575);
nor U34467 (N_34467,N_30064,N_30430);
xor U34468 (N_34468,N_31073,N_30600);
xnor U34469 (N_34469,N_31415,N_32324);
or U34470 (N_34470,N_30993,N_30644);
nand U34471 (N_34471,N_30927,N_32010);
nor U34472 (N_34472,N_30335,N_30632);
and U34473 (N_34473,N_31520,N_32272);
xnor U34474 (N_34474,N_31360,N_32403);
nor U34475 (N_34475,N_31793,N_30712);
xor U34476 (N_34476,N_32059,N_32218);
xor U34477 (N_34477,N_30583,N_30111);
nor U34478 (N_34478,N_31318,N_32458);
nand U34479 (N_34479,N_31551,N_32460);
nor U34480 (N_34480,N_31670,N_31411);
nand U34481 (N_34481,N_30042,N_32099);
or U34482 (N_34482,N_32354,N_31897);
xnor U34483 (N_34483,N_31077,N_32409);
or U34484 (N_34484,N_31839,N_32027);
nor U34485 (N_34485,N_31524,N_31762);
or U34486 (N_34486,N_30642,N_32093);
and U34487 (N_34487,N_31592,N_30469);
and U34488 (N_34488,N_31943,N_32357);
nor U34489 (N_34489,N_30302,N_31630);
nor U34490 (N_34490,N_31691,N_31559);
nand U34491 (N_34491,N_32068,N_30292);
xnor U34492 (N_34492,N_31337,N_31446);
nand U34493 (N_34493,N_32337,N_31567);
xnor U34494 (N_34494,N_30419,N_30644);
xor U34495 (N_34495,N_30622,N_31583);
xor U34496 (N_34496,N_31876,N_30733);
or U34497 (N_34497,N_30853,N_30609);
nor U34498 (N_34498,N_32421,N_32010);
nor U34499 (N_34499,N_31010,N_32299);
nand U34500 (N_34500,N_31953,N_30350);
xor U34501 (N_34501,N_30149,N_32477);
and U34502 (N_34502,N_32420,N_31750);
xor U34503 (N_34503,N_30759,N_31064);
xor U34504 (N_34504,N_30742,N_31858);
or U34505 (N_34505,N_30531,N_31526);
xnor U34506 (N_34506,N_30556,N_31613);
nand U34507 (N_34507,N_31072,N_30475);
nor U34508 (N_34508,N_32483,N_31211);
xor U34509 (N_34509,N_32406,N_30375);
xor U34510 (N_34510,N_32111,N_30530);
or U34511 (N_34511,N_31133,N_32288);
and U34512 (N_34512,N_30350,N_31424);
xnor U34513 (N_34513,N_30609,N_30033);
nand U34514 (N_34514,N_31677,N_31179);
nor U34515 (N_34515,N_31824,N_31222);
nand U34516 (N_34516,N_30821,N_31981);
nand U34517 (N_34517,N_30268,N_30400);
nand U34518 (N_34518,N_32044,N_32420);
and U34519 (N_34519,N_30570,N_31119);
nor U34520 (N_34520,N_31641,N_30372);
nor U34521 (N_34521,N_31048,N_31370);
xnor U34522 (N_34522,N_30418,N_31115);
or U34523 (N_34523,N_30956,N_31369);
xor U34524 (N_34524,N_30710,N_30647);
nand U34525 (N_34525,N_30111,N_32292);
nand U34526 (N_34526,N_31061,N_31704);
nand U34527 (N_34527,N_32449,N_30517);
nor U34528 (N_34528,N_31655,N_31825);
nor U34529 (N_34529,N_31052,N_31125);
xnor U34530 (N_34530,N_31672,N_31005);
or U34531 (N_34531,N_30109,N_30551);
nor U34532 (N_34532,N_30405,N_31465);
xor U34533 (N_34533,N_30069,N_30142);
or U34534 (N_34534,N_31479,N_30508);
or U34535 (N_34535,N_31229,N_32351);
or U34536 (N_34536,N_31756,N_32487);
xnor U34537 (N_34537,N_30109,N_31590);
xor U34538 (N_34538,N_32375,N_30203);
xnor U34539 (N_34539,N_30221,N_30509);
xnor U34540 (N_34540,N_32062,N_30538);
xnor U34541 (N_34541,N_31851,N_30571);
nor U34542 (N_34542,N_30873,N_32273);
xnor U34543 (N_34543,N_30986,N_30104);
xor U34544 (N_34544,N_32276,N_30255);
nor U34545 (N_34545,N_31971,N_32086);
or U34546 (N_34546,N_32354,N_32038);
xor U34547 (N_34547,N_32089,N_31811);
xor U34548 (N_34548,N_31008,N_30509);
xor U34549 (N_34549,N_30404,N_30984);
nor U34550 (N_34550,N_30847,N_31027);
and U34551 (N_34551,N_31734,N_32353);
or U34552 (N_34552,N_31093,N_32101);
nor U34553 (N_34553,N_31763,N_30027);
xnor U34554 (N_34554,N_31887,N_32057);
nand U34555 (N_34555,N_31672,N_30105);
and U34556 (N_34556,N_30943,N_32065);
and U34557 (N_34557,N_31815,N_32291);
and U34558 (N_34558,N_30287,N_32188);
nor U34559 (N_34559,N_32081,N_31606);
or U34560 (N_34560,N_31052,N_32334);
nor U34561 (N_34561,N_30129,N_30046);
nand U34562 (N_34562,N_30849,N_30430);
and U34563 (N_34563,N_30589,N_31647);
and U34564 (N_34564,N_32397,N_30665);
xor U34565 (N_34565,N_30622,N_30673);
nand U34566 (N_34566,N_32391,N_30270);
nor U34567 (N_34567,N_30655,N_30053);
xnor U34568 (N_34568,N_32040,N_30600);
and U34569 (N_34569,N_30246,N_31768);
nand U34570 (N_34570,N_30440,N_31636);
or U34571 (N_34571,N_32255,N_30546);
nor U34572 (N_34572,N_31210,N_31608);
xor U34573 (N_34573,N_31737,N_30642);
nor U34574 (N_34574,N_31853,N_31816);
or U34575 (N_34575,N_30031,N_31631);
nand U34576 (N_34576,N_31372,N_30297);
and U34577 (N_34577,N_30654,N_31732);
xnor U34578 (N_34578,N_30412,N_31706);
xor U34579 (N_34579,N_30004,N_31504);
and U34580 (N_34580,N_31275,N_31183);
and U34581 (N_34581,N_30787,N_30989);
nor U34582 (N_34582,N_32226,N_30091);
nor U34583 (N_34583,N_32186,N_30252);
nand U34584 (N_34584,N_30974,N_31280);
nand U34585 (N_34585,N_31230,N_31307);
nand U34586 (N_34586,N_31649,N_32071);
xnor U34587 (N_34587,N_31653,N_30449);
nand U34588 (N_34588,N_30940,N_30117);
nand U34589 (N_34589,N_30859,N_32471);
and U34590 (N_34590,N_30183,N_30665);
nor U34591 (N_34591,N_31309,N_30164);
xnor U34592 (N_34592,N_31906,N_31128);
or U34593 (N_34593,N_31211,N_32337);
xnor U34594 (N_34594,N_31432,N_30325);
nor U34595 (N_34595,N_31891,N_32051);
nand U34596 (N_34596,N_30130,N_32135);
and U34597 (N_34597,N_31783,N_31301);
and U34598 (N_34598,N_31730,N_31679);
and U34599 (N_34599,N_30712,N_30442);
or U34600 (N_34600,N_30676,N_32216);
and U34601 (N_34601,N_31557,N_31354);
nand U34602 (N_34602,N_30606,N_31534);
nor U34603 (N_34603,N_30598,N_31862);
and U34604 (N_34604,N_32322,N_31501);
and U34605 (N_34605,N_30906,N_31997);
xnor U34606 (N_34606,N_31333,N_30446);
nor U34607 (N_34607,N_31238,N_30083);
or U34608 (N_34608,N_30901,N_30900);
and U34609 (N_34609,N_30286,N_30129);
and U34610 (N_34610,N_31364,N_31203);
or U34611 (N_34611,N_30205,N_31682);
nor U34612 (N_34612,N_31267,N_31309);
nor U34613 (N_34613,N_30579,N_32186);
or U34614 (N_34614,N_32372,N_30716);
xor U34615 (N_34615,N_30945,N_30224);
nand U34616 (N_34616,N_31001,N_31519);
xnor U34617 (N_34617,N_30720,N_31112);
nand U34618 (N_34618,N_30863,N_31265);
and U34619 (N_34619,N_30567,N_30388);
nand U34620 (N_34620,N_30915,N_30663);
nand U34621 (N_34621,N_30847,N_31270);
and U34622 (N_34622,N_31164,N_31599);
and U34623 (N_34623,N_30355,N_30160);
and U34624 (N_34624,N_31920,N_31268);
or U34625 (N_34625,N_32386,N_30939);
or U34626 (N_34626,N_31985,N_30771);
or U34627 (N_34627,N_31672,N_31170);
xnor U34628 (N_34628,N_30575,N_32170);
nand U34629 (N_34629,N_31919,N_31576);
and U34630 (N_34630,N_32454,N_30406);
or U34631 (N_34631,N_30477,N_30192);
and U34632 (N_34632,N_30307,N_31299);
nor U34633 (N_34633,N_30019,N_30144);
xor U34634 (N_34634,N_32463,N_31552);
xnor U34635 (N_34635,N_30823,N_31461);
nor U34636 (N_34636,N_30851,N_30534);
or U34637 (N_34637,N_32405,N_31922);
or U34638 (N_34638,N_31073,N_31050);
or U34639 (N_34639,N_30196,N_31517);
and U34640 (N_34640,N_32264,N_30281);
nand U34641 (N_34641,N_31039,N_32318);
xor U34642 (N_34642,N_32466,N_32202);
nand U34643 (N_34643,N_30356,N_31275);
nand U34644 (N_34644,N_31481,N_31393);
or U34645 (N_34645,N_30579,N_30860);
or U34646 (N_34646,N_30142,N_30641);
nand U34647 (N_34647,N_31096,N_31848);
xnor U34648 (N_34648,N_32349,N_31192);
nor U34649 (N_34649,N_30770,N_30558);
and U34650 (N_34650,N_31409,N_32339);
nor U34651 (N_34651,N_31655,N_32285);
nor U34652 (N_34652,N_31076,N_30660);
xnor U34653 (N_34653,N_30783,N_31836);
and U34654 (N_34654,N_32178,N_30272);
or U34655 (N_34655,N_30541,N_31805);
or U34656 (N_34656,N_30958,N_31169);
xnor U34657 (N_34657,N_31215,N_32279);
and U34658 (N_34658,N_30645,N_31342);
nand U34659 (N_34659,N_31955,N_30663);
nand U34660 (N_34660,N_31867,N_31301);
and U34661 (N_34661,N_30808,N_31633);
nor U34662 (N_34662,N_31273,N_31924);
or U34663 (N_34663,N_31242,N_32393);
or U34664 (N_34664,N_31285,N_32365);
or U34665 (N_34665,N_30244,N_32267);
nor U34666 (N_34666,N_30848,N_30855);
and U34667 (N_34667,N_32276,N_31961);
nand U34668 (N_34668,N_30863,N_30759);
and U34669 (N_34669,N_31131,N_32297);
and U34670 (N_34670,N_30382,N_30116);
nand U34671 (N_34671,N_31432,N_30560);
nor U34672 (N_34672,N_31437,N_32123);
nand U34673 (N_34673,N_31913,N_31781);
and U34674 (N_34674,N_31523,N_30893);
xor U34675 (N_34675,N_32066,N_30490);
or U34676 (N_34676,N_30559,N_31394);
nand U34677 (N_34677,N_30049,N_31983);
xnor U34678 (N_34678,N_31442,N_30320);
nand U34679 (N_34679,N_31842,N_31442);
nor U34680 (N_34680,N_32153,N_31608);
or U34681 (N_34681,N_30781,N_30585);
or U34682 (N_34682,N_31087,N_30473);
or U34683 (N_34683,N_32199,N_32242);
and U34684 (N_34684,N_30824,N_32348);
xnor U34685 (N_34685,N_30066,N_30266);
xor U34686 (N_34686,N_30937,N_30618);
nand U34687 (N_34687,N_31096,N_30892);
or U34688 (N_34688,N_31062,N_30734);
xnor U34689 (N_34689,N_30101,N_31517);
nor U34690 (N_34690,N_31832,N_31595);
and U34691 (N_34691,N_32068,N_32430);
xnor U34692 (N_34692,N_30973,N_30384);
nor U34693 (N_34693,N_31007,N_32394);
or U34694 (N_34694,N_30579,N_30516);
nor U34695 (N_34695,N_30810,N_30528);
xor U34696 (N_34696,N_32190,N_31478);
nor U34697 (N_34697,N_31984,N_32283);
nand U34698 (N_34698,N_30876,N_30182);
nor U34699 (N_34699,N_30116,N_31325);
nand U34700 (N_34700,N_32282,N_31940);
nand U34701 (N_34701,N_30840,N_30100);
and U34702 (N_34702,N_31261,N_30525);
xnor U34703 (N_34703,N_30084,N_31617);
and U34704 (N_34704,N_32232,N_30591);
or U34705 (N_34705,N_30581,N_30984);
nor U34706 (N_34706,N_31189,N_30397);
or U34707 (N_34707,N_32202,N_32237);
xnor U34708 (N_34708,N_30683,N_30216);
or U34709 (N_34709,N_31006,N_31957);
and U34710 (N_34710,N_32005,N_30377);
or U34711 (N_34711,N_31765,N_32225);
and U34712 (N_34712,N_30184,N_31487);
nand U34713 (N_34713,N_30839,N_30833);
and U34714 (N_34714,N_32388,N_32068);
xor U34715 (N_34715,N_31107,N_31332);
nand U34716 (N_34716,N_32489,N_30343);
nand U34717 (N_34717,N_32283,N_30831);
or U34718 (N_34718,N_30551,N_30613);
or U34719 (N_34719,N_30011,N_30489);
xor U34720 (N_34720,N_31983,N_31847);
and U34721 (N_34721,N_31752,N_31305);
and U34722 (N_34722,N_31962,N_31775);
and U34723 (N_34723,N_30955,N_32307);
nand U34724 (N_34724,N_30726,N_32018);
and U34725 (N_34725,N_32107,N_31436);
xnor U34726 (N_34726,N_31169,N_30307);
nand U34727 (N_34727,N_30454,N_30298);
and U34728 (N_34728,N_30293,N_30878);
nor U34729 (N_34729,N_31890,N_30217);
nand U34730 (N_34730,N_30669,N_30920);
nand U34731 (N_34731,N_32181,N_31471);
nand U34732 (N_34732,N_32048,N_30762);
xnor U34733 (N_34733,N_30361,N_30910);
or U34734 (N_34734,N_31153,N_30157);
and U34735 (N_34735,N_30171,N_30323);
xnor U34736 (N_34736,N_30954,N_30910);
nand U34737 (N_34737,N_30257,N_30163);
or U34738 (N_34738,N_31557,N_31357);
nand U34739 (N_34739,N_31242,N_32399);
nor U34740 (N_34740,N_32264,N_32370);
nor U34741 (N_34741,N_30136,N_30766);
nor U34742 (N_34742,N_31200,N_31106);
nand U34743 (N_34743,N_30746,N_32160);
xnor U34744 (N_34744,N_31102,N_31126);
nor U34745 (N_34745,N_31205,N_30428);
nor U34746 (N_34746,N_30521,N_30943);
or U34747 (N_34747,N_30380,N_30669);
xnor U34748 (N_34748,N_30171,N_31303);
or U34749 (N_34749,N_30896,N_31553);
nor U34750 (N_34750,N_30588,N_30901);
nand U34751 (N_34751,N_30182,N_32214);
xnor U34752 (N_34752,N_31356,N_30462);
or U34753 (N_34753,N_31600,N_31456);
xor U34754 (N_34754,N_30556,N_30653);
and U34755 (N_34755,N_30081,N_32001);
nor U34756 (N_34756,N_30407,N_32274);
or U34757 (N_34757,N_32129,N_32448);
nor U34758 (N_34758,N_32052,N_31938);
and U34759 (N_34759,N_30282,N_32032);
nor U34760 (N_34760,N_31797,N_30402);
xnor U34761 (N_34761,N_30460,N_31946);
xnor U34762 (N_34762,N_30832,N_30342);
and U34763 (N_34763,N_31554,N_31697);
and U34764 (N_34764,N_31551,N_30598);
xnor U34765 (N_34765,N_31833,N_31386);
and U34766 (N_34766,N_30472,N_31713);
and U34767 (N_34767,N_31496,N_30696);
and U34768 (N_34768,N_31374,N_32446);
or U34769 (N_34769,N_31779,N_31561);
xor U34770 (N_34770,N_31563,N_31721);
or U34771 (N_34771,N_32219,N_32058);
xnor U34772 (N_34772,N_31182,N_30120);
and U34773 (N_34773,N_30189,N_32331);
or U34774 (N_34774,N_30612,N_30853);
or U34775 (N_34775,N_30529,N_32155);
and U34776 (N_34776,N_32235,N_32060);
nor U34777 (N_34777,N_30048,N_31438);
and U34778 (N_34778,N_31950,N_30290);
xnor U34779 (N_34779,N_32052,N_30502);
or U34780 (N_34780,N_31241,N_31272);
xor U34781 (N_34781,N_32371,N_30208);
or U34782 (N_34782,N_32401,N_32450);
xnor U34783 (N_34783,N_32285,N_32104);
or U34784 (N_34784,N_32445,N_30486);
nand U34785 (N_34785,N_31843,N_30451);
xnor U34786 (N_34786,N_32331,N_32486);
and U34787 (N_34787,N_30117,N_31706);
or U34788 (N_34788,N_30574,N_31013);
or U34789 (N_34789,N_32185,N_30361);
nor U34790 (N_34790,N_31604,N_32181);
or U34791 (N_34791,N_31370,N_31591);
xor U34792 (N_34792,N_31128,N_30620);
nor U34793 (N_34793,N_32164,N_31294);
nand U34794 (N_34794,N_30794,N_30965);
nor U34795 (N_34795,N_31594,N_30059);
nand U34796 (N_34796,N_30090,N_32005);
nor U34797 (N_34797,N_30469,N_31307);
nor U34798 (N_34798,N_30266,N_30018);
or U34799 (N_34799,N_31346,N_31134);
and U34800 (N_34800,N_30092,N_31331);
xor U34801 (N_34801,N_31297,N_30245);
nand U34802 (N_34802,N_31273,N_30937);
nor U34803 (N_34803,N_31320,N_30923);
nor U34804 (N_34804,N_30751,N_30845);
and U34805 (N_34805,N_30084,N_31411);
xnor U34806 (N_34806,N_30616,N_30943);
or U34807 (N_34807,N_30700,N_31708);
xor U34808 (N_34808,N_30874,N_31371);
or U34809 (N_34809,N_30677,N_32246);
xor U34810 (N_34810,N_30812,N_32372);
xnor U34811 (N_34811,N_31324,N_31419);
nand U34812 (N_34812,N_31466,N_30859);
or U34813 (N_34813,N_30632,N_31378);
nand U34814 (N_34814,N_31976,N_32138);
nor U34815 (N_34815,N_30952,N_32368);
nor U34816 (N_34816,N_30216,N_30078);
or U34817 (N_34817,N_31471,N_32031);
nand U34818 (N_34818,N_30458,N_31240);
xor U34819 (N_34819,N_31201,N_30332);
and U34820 (N_34820,N_31089,N_30828);
xnor U34821 (N_34821,N_30267,N_32261);
nand U34822 (N_34822,N_32088,N_30158);
or U34823 (N_34823,N_31649,N_30838);
nand U34824 (N_34824,N_30204,N_32152);
and U34825 (N_34825,N_31144,N_30642);
and U34826 (N_34826,N_32415,N_30144);
nor U34827 (N_34827,N_31778,N_31924);
nand U34828 (N_34828,N_31541,N_31940);
or U34829 (N_34829,N_31820,N_32254);
nor U34830 (N_34830,N_30822,N_31779);
nand U34831 (N_34831,N_30722,N_30893);
and U34832 (N_34832,N_30562,N_30118);
nand U34833 (N_34833,N_31142,N_31157);
and U34834 (N_34834,N_31782,N_30692);
nor U34835 (N_34835,N_32230,N_30267);
and U34836 (N_34836,N_31492,N_30670);
xnor U34837 (N_34837,N_31162,N_30795);
or U34838 (N_34838,N_32297,N_32378);
and U34839 (N_34839,N_32278,N_31492);
xnor U34840 (N_34840,N_32120,N_32473);
and U34841 (N_34841,N_30851,N_32015);
xor U34842 (N_34842,N_31487,N_31271);
and U34843 (N_34843,N_32011,N_30282);
xor U34844 (N_34844,N_30887,N_30614);
xor U34845 (N_34845,N_32357,N_31919);
xnor U34846 (N_34846,N_31592,N_30374);
nand U34847 (N_34847,N_32173,N_31468);
or U34848 (N_34848,N_30583,N_31692);
xor U34849 (N_34849,N_30093,N_30930);
nor U34850 (N_34850,N_31201,N_30777);
nor U34851 (N_34851,N_30809,N_31312);
or U34852 (N_34852,N_30146,N_32323);
nand U34853 (N_34853,N_30493,N_31542);
or U34854 (N_34854,N_30482,N_32116);
nor U34855 (N_34855,N_31125,N_31852);
or U34856 (N_34856,N_31301,N_30669);
nand U34857 (N_34857,N_30699,N_31194);
xnor U34858 (N_34858,N_30619,N_31178);
nand U34859 (N_34859,N_30506,N_30596);
xor U34860 (N_34860,N_31650,N_30200);
or U34861 (N_34861,N_30537,N_30733);
or U34862 (N_34862,N_30300,N_31484);
and U34863 (N_34863,N_30484,N_32149);
and U34864 (N_34864,N_30417,N_30763);
nor U34865 (N_34865,N_31076,N_30656);
and U34866 (N_34866,N_31213,N_30252);
nor U34867 (N_34867,N_31091,N_31213);
nor U34868 (N_34868,N_31380,N_30466);
or U34869 (N_34869,N_30068,N_30552);
nand U34870 (N_34870,N_31622,N_31678);
nor U34871 (N_34871,N_31656,N_30307);
nor U34872 (N_34872,N_30737,N_30654);
nor U34873 (N_34873,N_31979,N_30468);
xnor U34874 (N_34874,N_30308,N_31542);
and U34875 (N_34875,N_31846,N_31169);
xnor U34876 (N_34876,N_31421,N_32347);
xor U34877 (N_34877,N_30947,N_31292);
xor U34878 (N_34878,N_31756,N_31006);
or U34879 (N_34879,N_31424,N_32294);
xnor U34880 (N_34880,N_31262,N_31303);
and U34881 (N_34881,N_31402,N_32475);
nor U34882 (N_34882,N_30285,N_30028);
xor U34883 (N_34883,N_30845,N_30335);
nand U34884 (N_34884,N_32171,N_32206);
and U34885 (N_34885,N_32327,N_30901);
nor U34886 (N_34886,N_32137,N_31848);
or U34887 (N_34887,N_31116,N_30336);
xnor U34888 (N_34888,N_30714,N_31803);
xor U34889 (N_34889,N_31958,N_31372);
nand U34890 (N_34890,N_32005,N_30137);
or U34891 (N_34891,N_31932,N_32472);
nand U34892 (N_34892,N_30232,N_32443);
nand U34893 (N_34893,N_31863,N_30539);
and U34894 (N_34894,N_31980,N_31642);
nand U34895 (N_34895,N_30409,N_30191);
nor U34896 (N_34896,N_32206,N_31419);
nor U34897 (N_34897,N_31623,N_30234);
nor U34898 (N_34898,N_31036,N_30319);
nor U34899 (N_34899,N_31706,N_31393);
nor U34900 (N_34900,N_32173,N_30957);
xnor U34901 (N_34901,N_30933,N_31686);
nand U34902 (N_34902,N_30389,N_32267);
nor U34903 (N_34903,N_31457,N_31119);
and U34904 (N_34904,N_30551,N_31999);
xnor U34905 (N_34905,N_30506,N_32057);
nor U34906 (N_34906,N_31457,N_30049);
xor U34907 (N_34907,N_30148,N_32270);
or U34908 (N_34908,N_30052,N_30797);
xnor U34909 (N_34909,N_32081,N_31320);
xnor U34910 (N_34910,N_30277,N_30158);
or U34911 (N_34911,N_32041,N_32018);
nor U34912 (N_34912,N_31560,N_31807);
or U34913 (N_34913,N_32247,N_31624);
or U34914 (N_34914,N_32024,N_30749);
and U34915 (N_34915,N_30961,N_32023);
and U34916 (N_34916,N_31370,N_32397);
or U34917 (N_34917,N_31210,N_31888);
nor U34918 (N_34918,N_30861,N_32138);
nor U34919 (N_34919,N_32449,N_31458);
and U34920 (N_34920,N_32299,N_30042);
xnor U34921 (N_34921,N_31280,N_31445);
or U34922 (N_34922,N_31996,N_32454);
nor U34923 (N_34923,N_30731,N_31062);
nor U34924 (N_34924,N_31993,N_30373);
xnor U34925 (N_34925,N_30472,N_31570);
nor U34926 (N_34926,N_31459,N_30361);
xnor U34927 (N_34927,N_30292,N_32107);
nor U34928 (N_34928,N_31417,N_32254);
nor U34929 (N_34929,N_32352,N_31035);
nor U34930 (N_34930,N_31947,N_31945);
xor U34931 (N_34931,N_30161,N_31900);
and U34932 (N_34932,N_30816,N_31751);
or U34933 (N_34933,N_30644,N_31756);
nand U34934 (N_34934,N_31386,N_31413);
and U34935 (N_34935,N_31969,N_32063);
and U34936 (N_34936,N_30166,N_32116);
and U34937 (N_34937,N_32226,N_30349);
nor U34938 (N_34938,N_31254,N_30523);
nand U34939 (N_34939,N_30330,N_32023);
nor U34940 (N_34940,N_30273,N_31931);
nand U34941 (N_34941,N_30752,N_32381);
nor U34942 (N_34942,N_30140,N_32141);
nor U34943 (N_34943,N_32146,N_30691);
and U34944 (N_34944,N_31418,N_31635);
or U34945 (N_34945,N_32470,N_30047);
and U34946 (N_34946,N_32100,N_31768);
xor U34947 (N_34947,N_30756,N_31585);
and U34948 (N_34948,N_30464,N_31916);
nand U34949 (N_34949,N_31719,N_32442);
and U34950 (N_34950,N_30035,N_32070);
nand U34951 (N_34951,N_31595,N_31588);
nor U34952 (N_34952,N_30643,N_30211);
nand U34953 (N_34953,N_30259,N_31167);
nor U34954 (N_34954,N_30879,N_31666);
xor U34955 (N_34955,N_30337,N_32198);
nand U34956 (N_34956,N_30710,N_32227);
or U34957 (N_34957,N_31782,N_31187);
nor U34958 (N_34958,N_32435,N_30409);
nor U34959 (N_34959,N_32255,N_30729);
nand U34960 (N_34960,N_31368,N_30192);
or U34961 (N_34961,N_32344,N_32490);
and U34962 (N_34962,N_31587,N_32001);
nor U34963 (N_34963,N_31400,N_31823);
xor U34964 (N_34964,N_31712,N_32252);
xnor U34965 (N_34965,N_31424,N_30896);
xnor U34966 (N_34966,N_30426,N_30043);
nand U34967 (N_34967,N_32176,N_30239);
or U34968 (N_34968,N_31913,N_30923);
nand U34969 (N_34969,N_30974,N_31114);
xor U34970 (N_34970,N_32427,N_31858);
xor U34971 (N_34971,N_31833,N_30993);
or U34972 (N_34972,N_32290,N_30007);
xnor U34973 (N_34973,N_30688,N_31935);
nand U34974 (N_34974,N_31531,N_30930);
nand U34975 (N_34975,N_31986,N_31872);
and U34976 (N_34976,N_31593,N_30666);
xor U34977 (N_34977,N_31738,N_31195);
and U34978 (N_34978,N_31745,N_32326);
nand U34979 (N_34979,N_31766,N_30772);
xnor U34980 (N_34980,N_31555,N_30752);
nor U34981 (N_34981,N_31768,N_32475);
and U34982 (N_34982,N_31902,N_31581);
nor U34983 (N_34983,N_31390,N_32489);
nand U34984 (N_34984,N_30525,N_31293);
or U34985 (N_34985,N_30426,N_32267);
xor U34986 (N_34986,N_30520,N_31768);
nor U34987 (N_34987,N_30702,N_30779);
nand U34988 (N_34988,N_31427,N_30047);
nor U34989 (N_34989,N_30502,N_31501);
nor U34990 (N_34990,N_31753,N_31636);
xor U34991 (N_34991,N_30286,N_32371);
and U34992 (N_34992,N_31333,N_30619);
or U34993 (N_34993,N_30308,N_30230);
nor U34994 (N_34994,N_32186,N_31397);
nand U34995 (N_34995,N_30187,N_31460);
nand U34996 (N_34996,N_30390,N_31163);
nor U34997 (N_34997,N_31994,N_30638);
xor U34998 (N_34998,N_31809,N_31211);
and U34999 (N_34999,N_31588,N_30571);
xnor U35000 (N_35000,N_34448,N_34313);
and U35001 (N_35001,N_34523,N_34743);
and U35002 (N_35002,N_34581,N_33321);
or U35003 (N_35003,N_34425,N_33579);
nor U35004 (N_35004,N_33815,N_34783);
nand U35005 (N_35005,N_34476,N_32833);
nand U35006 (N_35006,N_34121,N_33340);
xnor U35007 (N_35007,N_33115,N_33374);
nor U35008 (N_35008,N_33810,N_34629);
xor U35009 (N_35009,N_34284,N_32899);
nand U35010 (N_35010,N_33848,N_32936);
and U35011 (N_35011,N_32914,N_34498);
and U35012 (N_35012,N_33934,N_34630);
and U35013 (N_35013,N_33492,N_32657);
or U35014 (N_35014,N_34037,N_33763);
nand U35015 (N_35015,N_34496,N_33314);
nand U35016 (N_35016,N_34068,N_34748);
nor U35017 (N_35017,N_33277,N_32993);
and U35018 (N_35018,N_32977,N_33935);
and U35019 (N_35019,N_34534,N_33705);
or U35020 (N_35020,N_33610,N_34938);
or U35021 (N_35021,N_34773,N_33731);
nor U35022 (N_35022,N_32901,N_34461);
and U35023 (N_35023,N_32644,N_34031);
nor U35024 (N_35024,N_33615,N_32837);
xnor U35025 (N_35025,N_33226,N_32806);
nor U35026 (N_35026,N_33104,N_33920);
xor U35027 (N_35027,N_34598,N_33549);
xnor U35028 (N_35028,N_33659,N_34660);
nand U35029 (N_35029,N_33852,N_34149);
nand U35030 (N_35030,N_33976,N_33926);
and U35031 (N_35031,N_34157,N_34678);
nor U35032 (N_35032,N_33708,N_34557);
nand U35033 (N_35033,N_34456,N_33042);
nor U35034 (N_35034,N_34004,N_33525);
or U35035 (N_35035,N_33805,N_33380);
and U35036 (N_35036,N_33213,N_32858);
and U35037 (N_35037,N_33139,N_34823);
or U35038 (N_35038,N_33790,N_33968);
and U35039 (N_35039,N_33393,N_34764);
or U35040 (N_35040,N_32821,N_33023);
nand U35041 (N_35041,N_33496,N_33202);
or U35042 (N_35042,N_33727,N_33644);
and U35043 (N_35043,N_33126,N_34306);
xor U35044 (N_35044,N_34072,N_33361);
and U35045 (N_35045,N_33105,N_33590);
or U35046 (N_35046,N_33501,N_34751);
and U35047 (N_35047,N_33983,N_34971);
or U35048 (N_35048,N_32687,N_34712);
nand U35049 (N_35049,N_33099,N_32947);
xor U35050 (N_35050,N_33307,N_32618);
nand U35051 (N_35051,N_34670,N_33047);
nor U35052 (N_35052,N_34744,N_33979);
nor U35053 (N_35053,N_33252,N_34277);
or U35054 (N_35054,N_33468,N_32729);
nor U35055 (N_35055,N_34194,N_33284);
or U35056 (N_35056,N_34305,N_33187);
and U35057 (N_35057,N_34835,N_32684);
or U35058 (N_35058,N_33214,N_32773);
nand U35059 (N_35059,N_32725,N_33089);
xor U35060 (N_35060,N_33000,N_34188);
nand U35061 (N_35061,N_33925,N_32791);
nand U35062 (N_35062,N_32873,N_33118);
nand U35063 (N_35063,N_34836,N_32979);
xor U35064 (N_35064,N_34969,N_33158);
xnor U35065 (N_35065,N_33565,N_32962);
or U35066 (N_35066,N_33973,N_34538);
and U35067 (N_35067,N_34303,N_34292);
nor U35068 (N_35068,N_33583,N_33410);
xnor U35069 (N_35069,N_33866,N_34316);
nor U35070 (N_35070,N_34260,N_33632);
xnor U35071 (N_35071,N_33399,N_33235);
xnor U35072 (N_35072,N_34834,N_33677);
or U35073 (N_35073,N_33312,N_33211);
or U35074 (N_35074,N_34162,N_34071);
nand U35075 (N_35075,N_34919,N_33945);
xnor U35076 (N_35076,N_32996,N_34936);
nand U35077 (N_35077,N_33617,N_33998);
and U35078 (N_35078,N_33980,N_34325);
nor U35079 (N_35079,N_34333,N_33512);
xnor U35080 (N_35080,N_32578,N_34424);
and U35081 (N_35081,N_34252,N_34628);
nor U35082 (N_35082,N_34694,N_34552);
nor U35083 (N_35083,N_33043,N_34457);
and U35084 (N_35084,N_33928,N_33210);
nand U35085 (N_35085,N_33335,N_33142);
and U35086 (N_35086,N_33624,N_33529);
nand U35087 (N_35087,N_33337,N_34626);
nor U35088 (N_35088,N_33379,N_34645);
nand U35089 (N_35089,N_34963,N_32814);
or U35090 (N_35090,N_34625,N_34524);
or U35091 (N_35091,N_34654,N_34433);
nand U35092 (N_35092,N_33301,N_33884);
xor U35093 (N_35093,N_33939,N_34314);
or U35094 (N_35094,N_34308,N_33865);
or U35095 (N_35095,N_34088,N_33627);
nor U35096 (N_35096,N_33030,N_33164);
nand U35097 (N_35097,N_33288,N_34736);
or U35098 (N_35098,N_32940,N_33206);
or U35099 (N_35099,N_34503,N_32963);
nor U35100 (N_35100,N_34055,N_32712);
nand U35101 (N_35101,N_34061,N_33630);
nand U35102 (N_35102,N_33290,N_34439);
nor U35103 (N_35103,N_33720,N_34792);
nor U35104 (N_35104,N_32988,N_33351);
xnor U35105 (N_35105,N_32860,N_34639);
and U35106 (N_35106,N_34819,N_32994);
nor U35107 (N_35107,N_33902,N_32722);
nand U35108 (N_35108,N_34803,N_33199);
or U35109 (N_35109,N_34817,N_33191);
nor U35110 (N_35110,N_34758,N_33446);
or U35111 (N_35111,N_33432,N_32894);
nor U35112 (N_35112,N_32749,N_33100);
or U35113 (N_35113,N_34018,N_34231);
and U35114 (N_35114,N_34367,N_34417);
nand U35115 (N_35115,N_34052,N_32561);
nor U35116 (N_35116,N_33083,N_34652);
nand U35117 (N_35117,N_33806,N_34992);
or U35118 (N_35118,N_34890,N_33192);
or U35119 (N_35119,N_33108,N_33480);
nor U35120 (N_35120,N_33362,N_34315);
and U35121 (N_35121,N_33128,N_34985);
xor U35122 (N_35122,N_33258,N_33072);
nand U35123 (N_35123,N_33029,N_34827);
and U35124 (N_35124,N_33656,N_34297);
xor U35125 (N_35125,N_32674,N_33596);
and U35126 (N_35126,N_34786,N_34454);
and U35127 (N_35127,N_33510,N_33240);
nor U35128 (N_35128,N_34261,N_33456);
xnor U35129 (N_35129,N_32699,N_34339);
or U35130 (N_35130,N_33531,N_34102);
xor U35131 (N_35131,N_34545,N_32670);
and U35132 (N_35132,N_34504,N_33260);
and U35133 (N_35133,N_33401,N_33227);
nor U35134 (N_35134,N_34691,N_34894);
xnor U35135 (N_35135,N_33909,N_33354);
nor U35136 (N_35136,N_32810,N_34093);
and U35137 (N_35137,N_34599,N_34832);
xnor U35138 (N_35138,N_32523,N_33500);
and U35139 (N_35139,N_32949,N_33699);
and U35140 (N_35140,N_34362,N_33882);
and U35141 (N_35141,N_33576,N_34405);
xnor U35142 (N_35142,N_33960,N_33355);
nor U35143 (N_35143,N_33435,N_34353);
and U35144 (N_35144,N_34531,N_33154);
nor U35145 (N_35145,N_32768,N_34126);
and U35146 (N_35146,N_32842,N_33800);
nand U35147 (N_35147,N_32807,N_33444);
nor U35148 (N_35148,N_33068,N_34506);
nand U35149 (N_35149,N_33838,N_34499);
and U35150 (N_35150,N_34582,N_32874);
xor U35151 (N_35151,N_34606,N_34595);
nor U35152 (N_35152,N_32642,N_33103);
or U35153 (N_35153,N_34198,N_34702);
xnor U35154 (N_35154,N_32702,N_33484);
nand U35155 (N_35155,N_32911,N_33259);
or U35156 (N_35156,N_33692,N_33863);
or U35157 (N_35157,N_33328,N_33864);
or U35158 (N_35158,N_32967,N_32841);
and U35159 (N_35159,N_34667,N_33660);
xnor U35160 (N_35160,N_34382,N_33333);
or U35161 (N_35161,N_33229,N_33106);
nor U35162 (N_35162,N_33704,N_33737);
nor U35163 (N_35163,N_34608,N_34212);
or U35164 (N_35164,N_34515,N_32844);
nor U35165 (N_35165,N_34885,N_32809);
or U35166 (N_35166,N_33069,N_32598);
xor U35167 (N_35167,N_33324,N_34273);
xor U35168 (N_35168,N_33276,N_33170);
nand U35169 (N_35169,N_32944,N_33777);
xnor U35170 (N_35170,N_33548,N_34972);
or U35171 (N_35171,N_32905,N_32533);
nor U35172 (N_35172,N_33051,N_34804);
and U35173 (N_35173,N_33709,N_34211);
nand U35174 (N_35174,N_32728,N_33534);
or U35175 (N_35175,N_34455,N_34167);
nand U35176 (N_35176,N_34214,N_32960);
nor U35177 (N_35177,N_34087,N_33070);
and U35178 (N_35178,N_33652,N_33987);
or U35179 (N_35179,N_33894,N_34540);
nor U35180 (N_35180,N_33918,N_33936);
nor U35181 (N_35181,N_32827,N_33901);
nand U35182 (N_35182,N_32673,N_32521);
nor U35183 (N_35183,N_32585,N_32703);
xnor U35184 (N_35184,N_33948,N_34653);
nand U35185 (N_35185,N_34183,N_32504);
nor U35186 (N_35186,N_32694,N_33578);
xor U35187 (N_35187,N_34267,N_34726);
nor U35188 (N_35188,N_33491,N_33642);
and U35189 (N_35189,N_34006,N_33015);
nor U35190 (N_35190,N_32720,N_32715);
nand U35191 (N_35191,N_33411,N_32519);
nand U35192 (N_35192,N_33779,N_33670);
nand U35193 (N_35193,N_32916,N_32678);
or U35194 (N_35194,N_33268,N_33001);
or U35195 (N_35195,N_32972,N_33765);
and U35196 (N_35196,N_34798,N_34710);
xor U35197 (N_35197,N_34255,N_32711);
nand U35198 (N_35198,N_34911,N_32737);
xor U35199 (N_35199,N_33651,N_33357);
nor U35200 (N_35200,N_33829,N_32924);
or U35201 (N_35201,N_34522,N_32835);
and U35202 (N_35202,N_33378,N_34650);
and U35203 (N_35203,N_34579,N_32600);
and U35204 (N_35204,N_34427,N_34727);
xnor U35205 (N_35205,N_34283,N_34254);
nand U35206 (N_35206,N_34684,N_32796);
nor U35207 (N_35207,N_32650,N_34191);
nor U35208 (N_35208,N_33041,N_33772);
or U35209 (N_35209,N_32958,N_32552);
xnor U35210 (N_35210,N_34793,N_33915);
nand U35211 (N_35211,N_32632,N_34415);
nand U35212 (N_35212,N_32772,N_33917);
and U35213 (N_35213,N_32939,N_34663);
nand U35214 (N_35214,N_34551,N_34820);
and U35215 (N_35215,N_34091,N_32760);
and U35216 (N_35216,N_33239,N_34867);
and U35217 (N_35217,N_33178,N_33978);
nor U35218 (N_35218,N_33466,N_34022);
nor U35219 (N_35219,N_32647,N_33967);
nor U35220 (N_35220,N_34500,N_33336);
xnor U35221 (N_35221,N_32777,N_33021);
nor U35222 (N_35222,N_33817,N_33353);
xor U35223 (N_35223,N_33143,N_33940);
and U35224 (N_35224,N_34416,N_34081);
or U35225 (N_35225,N_34622,N_33782);
and U35226 (N_35226,N_33875,N_32513);
xnor U35227 (N_35227,N_34511,N_33587);
and U35228 (N_35228,N_33295,N_33825);
or U35229 (N_35229,N_34884,N_33741);
nand U35230 (N_35230,N_33219,N_32690);
nor U35231 (N_35231,N_34049,N_32630);
nor U35232 (N_35232,N_34145,N_34999);
xor U35233 (N_35233,N_33217,N_32525);
xnor U35234 (N_35234,N_33959,N_34830);
or U35235 (N_35235,N_33009,N_32984);
nor U35236 (N_35236,N_34891,N_34854);
nand U35237 (N_35237,N_33039,N_33962);
nor U35238 (N_35238,N_32654,N_33322);
xor U35239 (N_35239,N_32981,N_34734);
xor U35240 (N_35240,N_34860,N_34723);
nor U35241 (N_35241,N_32567,N_32802);
and U35242 (N_35242,N_34053,N_33236);
xnor U35243 (N_35243,N_34258,N_32652);
or U35244 (N_35244,N_33954,N_34208);
nand U35245 (N_35245,N_34100,N_33007);
xnor U35246 (N_35246,N_32787,N_33033);
xnor U35247 (N_35247,N_34458,N_34588);
nand U35248 (N_35248,N_32907,N_33752);
xnor U35249 (N_35249,N_33593,N_33345);
or U35250 (N_35250,N_34064,N_34440);
nand U35251 (N_35251,N_33700,N_34510);
nand U35252 (N_35252,N_33653,N_34253);
nor U35253 (N_35253,N_33136,N_34131);
nor U35254 (N_35254,N_34863,N_33847);
nor U35255 (N_35255,N_33286,N_33204);
and U35256 (N_35256,N_34327,N_33562);
xor U35257 (N_35257,N_33249,N_34352);
and U35258 (N_35258,N_34329,N_33231);
xor U35259 (N_35259,N_33332,N_32653);
or U35260 (N_35260,N_34442,N_33524);
nand U35261 (N_35261,N_32869,N_34922);
nand U35262 (N_35262,N_34613,N_34990);
nand U35263 (N_35263,N_33611,N_34568);
nand U35264 (N_35264,N_33119,N_32676);
xor U35265 (N_35265,N_32903,N_33110);
or U35266 (N_35266,N_32961,N_34943);
nand U35267 (N_35267,N_34815,N_33430);
and U35268 (N_35268,N_34393,N_32571);
nand U35269 (N_35269,N_32512,N_34430);
xor U35270 (N_35270,N_34173,N_33330);
nand U35271 (N_35271,N_33554,N_34507);
or U35272 (N_35272,N_34029,N_33405);
nor U35273 (N_35273,N_33996,N_33732);
and U35274 (N_35274,N_34226,N_34493);
and U35275 (N_35275,N_34828,N_34561);
nand U35276 (N_35276,N_33543,N_34364);
or U35277 (N_35277,N_33313,N_33963);
xor U35278 (N_35278,N_34624,N_34343);
xnor U35279 (N_35279,N_34365,N_33400);
and U35280 (N_35280,N_34806,N_34731);
nand U35281 (N_35281,N_34392,N_34024);
and U35282 (N_35282,N_34187,N_33190);
and U35283 (N_35283,N_34341,N_33280);
or U35284 (N_35284,N_34097,N_33366);
xnor U35285 (N_35285,N_33724,N_32782);
nand U35286 (N_35286,N_33818,N_33842);
and U35287 (N_35287,N_34346,N_33589);
or U35288 (N_35288,N_34218,N_34658);
or U35289 (N_35289,N_34117,N_34707);
or U35290 (N_35290,N_32534,N_34945);
and U35291 (N_35291,N_34428,N_33050);
nand U35292 (N_35292,N_34395,N_33076);
or U35293 (N_35293,N_34334,N_32691);
nor U35294 (N_35294,N_33426,N_34378);
and U35295 (N_35295,N_33470,N_33483);
and U35296 (N_35296,N_33157,N_32524);
nand U35297 (N_35297,N_34805,N_32861);
nor U35298 (N_35298,N_32774,N_32880);
nand U35299 (N_35299,N_32664,N_34620);
or U35300 (N_35300,N_32889,N_33547);
or U35301 (N_35301,N_32884,N_33486);
nor U35302 (N_35302,N_33747,N_34359);
or U35303 (N_35303,N_34192,N_33246);
and U35304 (N_35304,N_34889,N_34381);
and U35305 (N_35305,N_33306,N_34878);
xnor U35306 (N_35306,N_32666,N_34237);
nand U35307 (N_35307,N_33311,N_33661);
or U35308 (N_35308,N_34866,N_34368);
nand U35309 (N_35309,N_32502,N_32550);
and U35310 (N_35310,N_34175,N_34697);
xor U35311 (N_35311,N_32742,N_34408);
or U35312 (N_35312,N_33016,N_34358);
and U35313 (N_35313,N_32992,N_33442);
and U35314 (N_35314,N_33478,N_33497);
nor U35315 (N_35315,N_33580,N_34947);
nand U35316 (N_35316,N_34853,N_32727);
nand U35317 (N_35317,N_34310,N_34497);
and U35318 (N_35318,N_34057,N_34669);
or U35319 (N_35319,N_34577,N_33795);
nor U35320 (N_35320,N_34824,N_32544);
xor U35321 (N_35321,N_33880,N_33289);
xnor U35322 (N_35322,N_34763,N_32709);
nand U35323 (N_35323,N_33389,N_34997);
nor U35324 (N_35324,N_32932,N_33695);
and U35325 (N_35325,N_32815,N_33232);
and U35326 (N_35326,N_32843,N_34536);
and U35327 (N_35327,N_34423,N_34893);
nand U35328 (N_35328,N_34554,N_32797);
or U35329 (N_35329,N_32954,N_32516);
and U35330 (N_35330,N_34228,N_33930);
or U35331 (N_35331,N_34881,N_32770);
xor U35332 (N_35332,N_33261,N_34438);
xnor U35333 (N_35333,N_34281,N_33792);
and U35334 (N_35334,N_34956,N_33294);
xor U35335 (N_35335,N_32734,N_34485);
nor U35336 (N_35336,N_33436,N_32671);
or U35337 (N_35337,N_33155,N_33542);
or U35338 (N_35338,N_34528,N_34151);
and U35339 (N_35339,N_33734,N_33857);
and U35340 (N_35340,N_34459,N_33796);
nand U35341 (N_35341,N_32510,N_33736);
nand U35342 (N_35342,N_34583,N_34787);
or U35343 (N_35343,N_32917,N_32601);
nand U35344 (N_35344,N_34375,N_34099);
nor U35345 (N_35345,N_34908,N_33171);
xor U35346 (N_35346,N_34299,N_33844);
nor U35347 (N_35347,N_32568,N_34435);
nor U35348 (N_35348,N_34095,N_32934);
and U35349 (N_35349,N_34903,N_33092);
nor U35350 (N_35350,N_33783,N_34373);
nand U35351 (N_35351,N_32863,N_32978);
or U35352 (N_35352,N_34553,N_32877);
nor U35353 (N_35353,N_33101,N_34016);
xor U35354 (N_35354,N_34904,N_32898);
nand U35355 (N_35355,N_34342,N_34348);
nor U35356 (N_35356,N_34689,N_34322);
nor U35357 (N_35357,N_34671,N_33515);
and U35358 (N_35358,N_32915,N_33808);
or U35359 (N_35359,N_33740,N_32596);
nand U35360 (N_35360,N_33152,N_32970);
nor U35361 (N_35361,N_33640,N_34537);
nor U35362 (N_35362,N_32595,N_32526);
nor U35363 (N_35363,N_32562,N_33251);
nor U35364 (N_35364,N_33738,N_33600);
nor U35365 (N_35365,N_32704,N_33985);
nor U35366 (N_35366,N_33262,N_34794);
and U35367 (N_35367,N_34215,N_34789);
nor U35368 (N_35368,N_34711,N_34372);
nor U35369 (N_35369,N_34201,N_33384);
or U35370 (N_35370,N_34270,N_33801);
nand U35371 (N_35371,N_33561,N_33879);
xnor U35372 (N_35372,N_33612,N_34705);
nor U35373 (N_35373,N_34009,N_32738);
xor U35374 (N_35374,N_34810,N_34034);
and U35375 (N_35375,N_33634,N_33506);
and U35376 (N_35376,N_34740,N_32919);
nand U35377 (N_35377,N_34585,N_34739);
xnor U35378 (N_35378,N_32941,N_33212);
xnor U35379 (N_35379,N_33933,N_33304);
nor U35380 (N_35380,N_34855,N_34642);
nand U35381 (N_35381,N_32558,N_32681);
or U35382 (N_35382,N_34951,N_33176);
xnor U35383 (N_35383,N_34632,N_33673);
or U35384 (N_35384,N_33225,N_33165);
and U35385 (N_35385,N_33837,N_33823);
nand U35386 (N_35386,N_34140,N_33595);
nor U35387 (N_35387,N_34357,N_34054);
nor U35388 (N_35388,N_33356,N_33943);
nand U35389 (N_35389,N_33528,N_33216);
or U35390 (N_35390,N_33493,N_32823);
and U35391 (N_35391,N_33012,N_34488);
xor U35392 (N_35392,N_33602,N_34337);
xnor U35393 (N_35393,N_34513,N_33748);
nand U35394 (N_35394,N_34570,N_34478);
and U35395 (N_35395,N_34356,N_33994);
nand U35396 (N_35396,N_34470,N_33567);
nor U35397 (N_35397,N_33938,N_32689);
nor U35398 (N_35398,N_33876,N_33856);
or U35399 (N_35399,N_33148,N_34431);
nand U35400 (N_35400,N_33044,N_33490);
nor U35401 (N_35401,N_34877,N_34977);
and U35402 (N_35402,N_33413,N_34092);
and U35403 (N_35403,N_33745,N_33761);
nand U35404 (N_35404,N_33594,N_33953);
and U35405 (N_35405,N_32937,N_33417);
nand U35406 (N_35406,N_34244,N_33751);
nand U35407 (N_35407,N_33683,N_33889);
xnor U35408 (N_35408,N_33424,N_33318);
and U35409 (N_35409,N_34133,N_34136);
nor U35410 (N_35410,N_33887,N_33680);
nor U35411 (N_35411,N_34045,N_34900);
xnor U35412 (N_35412,N_32990,N_32918);
nand U35413 (N_35413,N_34812,N_34563);
nand U35414 (N_35414,N_33707,N_34238);
and U35415 (N_35415,N_34895,N_32549);
or U35416 (N_35416,N_34120,N_32626);
nor U35417 (N_35417,N_34482,N_32695);
nor U35418 (N_35418,N_34328,N_33387);
xor U35419 (N_35419,N_34135,N_34839);
xor U35420 (N_35420,N_33766,N_32518);
nand U35421 (N_35421,N_33568,N_34401);
and U35422 (N_35422,N_33907,N_34112);
nor U35423 (N_35423,N_34014,N_33180);
nand U35424 (N_35424,N_34869,N_33675);
nand U35425 (N_35425,N_34562,N_32622);
nand U35426 (N_35426,N_34926,N_33559);
nor U35427 (N_35427,N_32680,N_33981);
xnor U35428 (N_35428,N_33151,N_33555);
or U35429 (N_35429,N_34453,N_33767);
nand U35430 (N_35430,N_34268,N_34355);
nand U35431 (N_35431,N_34409,N_32538);
and U35432 (N_35432,N_32623,N_33693);
xor U35433 (N_35433,N_34287,N_34398);
xnor U35434 (N_35434,N_33317,N_32555);
nand U35435 (N_35435,N_33215,N_34086);
nand U35436 (N_35436,N_34648,N_33096);
and U35437 (N_35437,N_33545,N_32784);
xor U35438 (N_35438,N_34550,N_33722);
and U35439 (N_35439,N_33367,N_33679);
xnor U35440 (N_35440,N_34508,N_34760);
xor U35441 (N_35441,N_34130,N_33826);
nand U35442 (N_35442,N_34124,N_34021);
nand U35443 (N_35443,N_34814,N_33095);
nor U35444 (N_35444,N_33712,N_32638);
xnor U35445 (N_35445,N_32885,N_34471);
or U35446 (N_35446,N_33584,N_33034);
xnor U35447 (N_35447,N_34407,N_32926);
or U35448 (N_35448,N_33475,N_33682);
xnor U35449 (N_35449,N_33088,N_34330);
xor U35450 (N_35450,N_32672,N_34033);
nand U35451 (N_35451,N_33750,N_33167);
xnor U35452 (N_35452,N_33331,N_34206);
and U35453 (N_35453,N_32912,N_34125);
and U35454 (N_35454,N_32845,N_33438);
nand U35455 (N_35455,N_34605,N_34539);
nand U35456 (N_35456,N_34114,N_34616);
and U35457 (N_35457,N_33971,N_32635);
and U35458 (N_35458,N_34007,N_32879);
and U35459 (N_35459,N_34580,N_34347);
xor U35460 (N_35460,N_34360,N_33688);
or U35461 (N_35461,N_33363,N_34040);
xnor U35462 (N_35462,N_34477,N_32636);
or U35463 (N_35463,N_32648,N_34638);
nor U35464 (N_35464,N_34755,N_33418);
or U35465 (N_35465,N_34715,N_34901);
nor U35466 (N_35466,N_33858,N_33040);
xor U35467 (N_35467,N_32779,N_33522);
or U35468 (N_35468,N_33886,N_33035);
and U35469 (N_35469,N_32581,N_34189);
xor U35470 (N_35470,N_33485,N_33173);
and U35471 (N_35471,N_34321,N_34390);
and U35472 (N_35472,N_33282,N_34842);
nor U35473 (N_35473,N_34841,N_34469);
or U35474 (N_35474,N_32500,N_34899);
nor U35475 (N_35475,N_34171,N_32566);
nand U35476 (N_35476,N_34000,N_32862);
xnor U35477 (N_35477,N_33308,N_34176);
xor U35478 (N_35478,N_33819,N_34935);
or U35479 (N_35479,N_34032,N_33824);
and U35480 (N_35480,N_34934,N_34647);
nor U35481 (N_35481,N_34202,N_34002);
nor U35482 (N_35482,N_32882,N_34856);
nand U35483 (N_35483,N_33382,N_32640);
and U35484 (N_35484,N_34958,N_33121);
xnor U35485 (N_35485,N_33265,N_34600);
nand U35486 (N_35486,N_34116,N_33658);
nor U35487 (N_35487,N_34933,N_34023);
xnor U35488 (N_35488,N_33063,N_34491);
xor U35489 (N_35489,N_32649,N_34150);
xnor U35490 (N_35490,N_33460,N_32535);
nor U35491 (N_35491,N_33182,N_33017);
nand U35492 (N_35492,N_33992,N_33717);
or U35493 (N_35493,N_34475,N_32953);
or U35494 (N_35494,N_33686,N_33581);
and U35495 (N_35495,N_34155,N_33832);
xnor U35496 (N_35496,N_34084,N_33788);
or U35497 (N_35497,N_33274,N_34559);
nor U35498 (N_35498,N_34962,N_34396);
or U35499 (N_35499,N_33278,N_34419);
or U35500 (N_35500,N_32998,N_33133);
nor U35501 (N_35501,N_32783,N_33643);
and U35502 (N_35502,N_32700,N_33342);
nor U35503 (N_35503,N_33910,N_34222);
nor U35504 (N_35504,N_32875,N_34701);
nor U35505 (N_35505,N_34486,N_34278);
xnor U35506 (N_35506,N_33031,N_34833);
nand U35507 (N_35507,N_32706,N_32741);
nor U35508 (N_35508,N_33586,N_32633);
xor U35509 (N_35509,N_33323,N_34436);
nor U35510 (N_35510,N_32767,N_32769);
nand U35511 (N_35511,N_34722,N_33224);
xnor U35512 (N_35512,N_33377,N_34808);
nor U35513 (N_35513,N_32831,N_34627);
nor U35514 (N_35514,N_32748,N_34111);
nor U35515 (N_35515,N_34959,N_34777);
xor U35516 (N_35516,N_33997,N_33408);
or U35517 (N_35517,N_33368,N_32964);
xor U35518 (N_35518,N_33820,N_34008);
nand U35519 (N_35519,N_34849,N_34041);
and U35520 (N_35520,N_33955,N_34335);
nor U35521 (N_35521,N_34179,N_33447);
xnor U35522 (N_35522,N_32805,N_32923);
nor U35523 (N_35523,N_34324,N_34269);
nand U35524 (N_35524,N_34541,N_32560);
nor U35525 (N_35525,N_32505,N_34158);
nor U35526 (N_35526,N_34153,N_32982);
nor U35527 (N_35527,N_33637,N_33575);
nand U35528 (N_35528,N_34902,N_34251);
nor U35529 (N_35529,N_33409,N_33185);
xnor U35530 (N_35530,N_34509,N_34621);
nand U35531 (N_35531,N_34249,N_33625);
nand U35532 (N_35532,N_33455,N_34526);
or U35533 (N_35533,N_33947,N_33364);
or U35534 (N_35534,N_34818,N_32811);
xnor U35535 (N_35535,N_33538,N_34043);
nor U35536 (N_35536,N_33461,N_32818);
nor U35537 (N_35537,N_34848,N_32718);
and U35538 (N_35538,N_34400,N_32965);
nand U35539 (N_35539,N_33786,N_32620);
and U35540 (N_35540,N_33974,N_34949);
and U35541 (N_35541,N_33871,N_34354);
and U35542 (N_35542,N_32582,N_34429);
xor U35543 (N_35543,N_34615,N_34132);
nor U35544 (N_35544,N_34421,N_32624);
and U35545 (N_35545,N_32825,N_33293);
and U35546 (N_35546,N_32755,N_34593);
nand U35547 (N_35547,N_34730,N_33097);
nor U35548 (N_35548,N_33885,N_33450);
nor U35549 (N_35549,N_32857,N_33551);
nor U35550 (N_35550,N_34800,N_32832);
or U35551 (N_35551,N_34771,N_34144);
nor U35552 (N_35552,N_34858,N_33853);
and U35553 (N_35553,N_33846,N_34300);
nor U35554 (N_35554,N_33297,N_33729);
or U35555 (N_35555,N_33305,N_33471);
or U35556 (N_35556,N_32864,N_32929);
xnor U35557 (N_35557,N_34665,N_34484);
nor U35558 (N_35558,N_33020,N_34466);
and U35559 (N_35559,N_33757,N_32606);
nand U35560 (N_35560,N_34657,N_34385);
xor U35561 (N_35561,N_32865,N_33631);
and U35562 (N_35562,N_33991,N_32890);
nand U35563 (N_35563,N_34403,N_33903);
nand U35564 (N_35564,N_33609,N_32881);
nand U35565 (N_35565,N_33710,N_34161);
xor U35566 (N_35566,N_32628,N_33177);
nor U35567 (N_35567,N_34307,N_32599);
xor U35568 (N_35568,N_33591,N_32570);
nor U35569 (N_35569,N_33742,N_33681);
and U35570 (N_35570,N_33623,N_33055);
or U35571 (N_35571,N_33391,N_34750);
and U35572 (N_35572,N_34336,N_32829);
nor U35573 (N_35573,N_33124,N_33309);
or U35574 (N_35574,N_33776,N_32781);
and U35575 (N_35575,N_34123,N_33221);
or U35576 (N_35576,N_32780,N_34413);
xor U35577 (N_35577,N_34290,N_34474);
or U35578 (N_35578,N_33018,N_33739);
nand U35579 (N_35579,N_33343,N_34791);
xor U35580 (N_35580,N_34811,N_33385);
nor U35581 (N_35581,N_34449,N_34695);
or U35582 (N_35582,N_32580,N_32540);
nor U35583 (N_35583,N_33648,N_33546);
xor U35584 (N_35584,N_34274,N_33144);
xnor U35585 (N_35585,N_32589,N_33898);
nand U35586 (N_35586,N_33507,N_34604);
xor U35587 (N_35587,N_32789,N_33714);
and U35588 (N_35588,N_34070,N_32794);
nor U35589 (N_35589,N_32959,N_32995);
and U35590 (N_35590,N_33065,N_32710);
and U35591 (N_35591,N_33647,N_34432);
nand U35592 (N_35592,N_33621,N_34674);
xnor U35593 (N_35593,N_33395,N_34716);
or U35594 (N_35594,N_34871,N_32631);
nor U35595 (N_35595,N_34163,N_33560);
or U35596 (N_35596,N_34825,N_34746);
nand U35597 (N_35597,N_33431,N_33775);
nand U35598 (N_35598,N_34896,N_33462);
xor U35599 (N_35599,N_33989,N_34769);
nand U35600 (N_35600,N_34338,N_33785);
nand U35601 (N_35601,N_32745,N_34391);
nor U35602 (N_35602,N_33129,N_32515);
or U35603 (N_35603,N_34259,N_34193);
nand U35604 (N_35604,N_33616,N_34224);
and U35605 (N_35605,N_33607,N_33025);
xor U35606 (N_35606,N_33137,N_33965);
xor U35607 (N_35607,N_34344,N_33376);
or U35608 (N_35608,N_33420,N_33530);
xor U35609 (N_35609,N_34248,N_33827);
and U35610 (N_35610,N_33895,N_34350);
or U35611 (N_35611,N_32661,N_33622);
xor U35612 (N_35612,N_33196,N_32951);
nor U35613 (N_35613,N_34062,N_33912);
and U35614 (N_35614,N_34967,N_34184);
xor U35615 (N_35615,N_32529,N_34655);
and U35616 (N_35616,N_32514,N_33398);
and U35617 (N_35617,N_34756,N_32611);
nor U35618 (N_35618,N_34295,N_33564);
nor U35619 (N_35619,N_33753,N_33027);
nand U35620 (N_35620,N_33758,N_32507);
or U35621 (N_35621,N_33728,N_33339);
or U35622 (N_35622,N_34845,N_34565);
nor U35623 (N_35623,N_33762,N_34675);
or U35624 (N_35624,N_33476,N_32665);
nand U35625 (N_35625,N_33140,N_32655);
or U35626 (N_35626,N_33502,N_34098);
nand U35627 (N_35627,N_33181,N_34502);
nand U35628 (N_35628,N_33448,N_34569);
xor U35629 (N_35629,N_34318,N_33950);
nor U35630 (N_35630,N_33702,N_32563);
nand U35631 (N_35631,N_34857,N_33905);
nor U35632 (N_35632,N_34721,N_34177);
nor U35633 (N_35633,N_32634,N_34930);
or U35634 (N_35634,N_33526,N_33013);
and U35635 (N_35635,N_33924,N_34809);
nor U35636 (N_35636,N_32617,N_32743);
and U35637 (N_35637,N_33381,N_34351);
nand U35638 (N_35638,N_34544,N_33508);
or U35639 (N_35639,N_33156,N_33498);
and U35640 (N_35640,N_32747,N_34229);
nand U35641 (N_35641,N_33544,N_33371);
or U35642 (N_35642,N_33791,N_33888);
nor U35643 (N_35643,N_34148,N_34923);
xnor U35644 (N_35644,N_34137,N_32933);
and U35645 (N_35645,N_34380,N_34319);
or U35646 (N_35646,N_34205,N_32766);
nor U35647 (N_35647,N_33407,N_34242);
nor U35648 (N_35648,N_34075,N_33535);
nand U35649 (N_35649,N_33666,N_33678);
and U35650 (N_35650,N_32997,N_32731);
or U35651 (N_35651,N_33620,N_34916);
and U35652 (N_35652,N_32697,N_33834);
and U35653 (N_35653,N_34576,N_33325);
nor U35654 (N_35654,N_34699,N_33822);
xor U35655 (N_35655,N_33285,N_33893);
and U35656 (N_35656,N_33646,N_33588);
or U35657 (N_35657,N_32803,N_33883);
nor U35658 (N_35658,N_32974,N_34532);
and U35659 (N_35659,N_33457,N_32646);
xor U35660 (N_35660,N_34331,N_34566);
nand U35661 (N_35661,N_32786,N_33861);
or U35662 (N_35662,N_33599,N_34636);
xnor U35663 (N_35663,N_34452,N_33802);
or U35664 (N_35664,N_34957,N_32851);
nor U35665 (N_35665,N_32920,N_33107);
nand U35666 (N_35666,N_33797,N_33582);
nand U35667 (N_35667,N_33255,N_34236);
xnor U35668 (N_35668,N_32893,N_34005);
nand U35669 (N_35669,N_33166,N_34003);
nor U35670 (N_35670,N_34840,N_34914);
or U35671 (N_35671,N_33477,N_32651);
xor U35672 (N_35672,N_34056,N_34905);
nor U35673 (N_35673,N_34862,N_33756);
xor U35674 (N_35674,N_33862,N_34912);
nor U35675 (N_35675,N_34245,N_34924);
and U35676 (N_35676,N_34312,N_32572);
xor U35677 (N_35677,N_32956,N_33037);
xnor U35678 (N_35678,N_33603,N_32973);
and U35679 (N_35679,N_32577,N_34641);
nand U35680 (N_35680,N_32927,N_33669);
and U35681 (N_35681,N_34745,N_34596);
nor U35682 (N_35682,N_32547,N_34759);
or U35683 (N_35683,N_33566,N_32619);
nand U35684 (N_35684,N_32771,N_34156);
nand U35685 (N_35685,N_32928,N_34799);
nand U35686 (N_35686,N_34291,N_33084);
nand U35687 (N_35687,N_32641,N_34134);
xor U35688 (N_35688,N_34048,N_32759);
nor U35689 (N_35689,N_34386,N_32913);
and U35690 (N_35690,N_33906,N_34941);
and U35691 (N_35691,N_34272,N_33472);
xnor U35692 (N_35692,N_34463,N_34696);
nor U35693 (N_35693,N_33049,N_33764);
or U35694 (N_35694,N_32614,N_34781);
or U35695 (N_35695,N_34113,N_34406);
xor U35696 (N_35696,N_32537,N_33557);
nand U35697 (N_35697,N_33003,N_33302);
or U35698 (N_35698,N_32724,N_34426);
nand U35699 (N_35699,N_34573,N_33053);
nand U35700 (N_35700,N_34250,N_32853);
or U35701 (N_35701,N_33949,N_32985);
and U35702 (N_35702,N_33841,N_34241);
or U35703 (N_35703,N_33816,N_33505);
nand U35704 (N_35704,N_33189,N_33172);
or U35705 (N_35705,N_34742,N_33038);
xor U35706 (N_35706,N_33188,N_33969);
nand U35707 (N_35707,N_34185,N_34996);
nand U35708 (N_35708,N_32686,N_33944);
xor U35709 (N_35709,N_34897,N_34038);
or U35710 (N_35710,N_32946,N_33814);
nand U35711 (N_35711,N_33394,N_33234);
and U35712 (N_35712,N_33080,N_34944);
xor U35713 (N_35713,N_33071,N_34975);
xnor U35714 (N_35714,N_34837,N_34282);
and U35715 (N_35715,N_34059,N_34887);
or U35716 (N_35716,N_33111,N_33533);
and U35717 (N_35717,N_32902,N_34679);
and U35718 (N_35718,N_33706,N_32795);
and U35719 (N_35719,N_34169,N_32717);
xnor U35720 (N_35720,N_32758,N_34795);
and U35721 (N_35721,N_34402,N_34128);
nand U35722 (N_35722,N_33597,N_33558);
or U35723 (N_35723,N_33689,N_32945);
nor U35724 (N_35724,N_33629,N_34298);
or U35725 (N_35725,N_34235,N_32746);
xor U35726 (N_35726,N_34517,N_32804);
nor U35727 (N_35727,N_33984,N_34525);
or U35728 (N_35728,N_32682,N_33499);
or U35729 (N_35729,N_33014,N_33716);
nand U35730 (N_35730,N_34546,N_32931);
or U35731 (N_35731,N_34995,N_33798);
and U35732 (N_35732,N_34685,N_32817);
xnor U35733 (N_35733,N_33223,N_34529);
xor U35734 (N_35734,N_32888,N_34219);
or U35735 (N_35735,N_34389,N_33606);
nor U35736 (N_35736,N_34784,N_32586);
nand U35737 (N_35737,N_32859,N_33134);
nand U35738 (N_35738,N_33454,N_34190);
xnor U35739 (N_35739,N_33633,N_34414);
or U35740 (N_35740,N_33937,N_33877);
nor U35741 (N_35741,N_33059,N_32658);
xnor U35742 (N_35742,N_33671,N_34692);
and U35743 (N_35743,N_34578,N_34221);
nand U35744 (N_35744,N_33329,N_34547);
xnor U35745 (N_35745,N_34309,N_33123);
or U35746 (N_35746,N_34276,N_33334);
or U35747 (N_35747,N_33443,N_32757);
and U35748 (N_35748,N_32663,N_34141);
nand U35749 (N_35749,N_34607,N_33207);
or U35750 (N_35750,N_34079,N_34010);
nand U35751 (N_35751,N_32592,N_33197);
nor U35752 (N_35752,N_32612,N_34065);
xnor U35753 (N_35753,N_32904,N_33375);
and U35754 (N_35754,N_33093,N_33445);
or U35755 (N_35755,N_33032,N_34807);
or U35756 (N_35756,N_33469,N_32667);
nand U35757 (N_35757,N_34704,N_33760);
nor U35758 (N_35758,N_34479,N_32812);
nand U35759 (N_35759,N_33645,N_32613);
xor U35760 (N_35760,N_33010,N_32751);
xor U35761 (N_35761,N_34256,N_34637);
nor U35762 (N_35762,N_32506,N_34729);
xor U35763 (N_35763,N_34768,N_33464);
nor U35764 (N_35764,N_34618,N_34234);
and U35765 (N_35765,N_34662,N_33237);
xnor U35766 (N_35766,N_33439,N_34984);
nand U35767 (N_35767,N_33434,N_33899);
or U35768 (N_35768,N_34882,N_34910);
nand U35769 (N_35769,N_32527,N_33459);
xor U35770 (N_35770,N_33563,N_34932);
nor U35771 (N_35771,N_34770,N_34586);
nand U35772 (N_35772,N_33718,N_32813);
xnor U35773 (N_35773,N_33613,N_33977);
xnor U35774 (N_35774,N_33664,N_33452);
or U35775 (N_35775,N_34418,N_33098);
xnor U35776 (N_35776,N_34349,N_34886);
xor U35777 (N_35777,N_34286,N_33657);
nand U35778 (N_35778,N_34774,N_34672);
and U35779 (N_35779,N_33350,N_33701);
xnor U35780 (N_35780,N_34105,N_34266);
nand U35781 (N_35781,N_33303,N_34230);
nand U35782 (N_35782,N_34719,N_34673);
xor U35783 (N_35783,N_34993,N_34384);
xor U35784 (N_35784,N_34915,N_33573);
nand U35785 (N_35785,N_34974,N_34089);
nand U35786 (N_35786,N_33694,N_32713);
and U35787 (N_35787,N_32925,N_33536);
and U35788 (N_35788,N_32602,N_33744);
nor U35789 (N_35789,N_33403,N_33789);
and U35790 (N_35790,N_32616,N_33585);
xnor U35791 (N_35791,N_34634,N_34700);
or U35792 (N_35792,N_34994,N_33986);
xnor U35793 (N_35793,N_32501,N_33650);
or U35794 (N_35794,N_34542,N_32546);
nand U35795 (N_35795,N_34294,N_33222);
nand U35796 (N_35796,N_33230,N_34168);
xor U35797 (N_35797,N_34765,N_32520);
xor U35798 (N_35798,N_34913,N_34661);
and U35799 (N_35799,N_32639,N_34028);
nand U35800 (N_35800,N_33022,N_33125);
and U35801 (N_35801,N_33872,N_34960);
and U35802 (N_35802,N_33873,N_34483);
nand U35803 (N_35803,N_33067,N_34296);
or U35804 (N_35804,N_33243,N_34101);
and U35805 (N_35805,N_32800,N_33900);
and U35806 (N_35806,N_34521,N_33298);
or U35807 (N_35807,N_33254,N_34986);
and U35808 (N_35808,N_33075,N_34909);
nand U35809 (N_35809,N_34883,N_33614);
or U35810 (N_35810,N_34852,N_34533);
or U35811 (N_35811,N_34376,N_32938);
nor U35812 (N_35812,N_32705,N_34535);
or U35813 (N_35813,N_34146,N_34213);
nor U35814 (N_35814,N_33839,N_34527);
nand U35815 (N_35815,N_34159,N_34640);
nor U35816 (N_35816,N_34964,N_33932);
xor U35817 (N_35817,N_33415,N_32716);
nand U35818 (N_35818,N_33338,N_33754);
xnor U35819 (N_35819,N_33482,N_32878);
nor U35820 (N_35820,N_34978,N_32922);
or U35821 (N_35821,N_34998,N_33521);
nor U35822 (N_35822,N_33869,N_33060);
xnor U35823 (N_35823,N_33778,N_34107);
xnor U35824 (N_35824,N_34285,N_33636);
or U35825 (N_35825,N_34142,N_32594);
and U35826 (N_35826,N_32999,N_33299);
or U35827 (N_35827,N_33828,N_32871);
xnor U35828 (N_35828,N_33881,N_34572);
nand U35829 (N_35829,N_33275,N_34077);
or U35830 (N_35830,N_34688,N_33066);
nor U35831 (N_35831,N_34968,N_34954);
or U35832 (N_35832,N_34767,N_34646);
and U35833 (N_35833,N_34399,N_33203);
xnor U35834 (N_35834,N_34154,N_34437);
xor U35835 (N_35835,N_34831,N_34464);
xor U35836 (N_35836,N_34779,N_34044);
xnor U35837 (N_35837,N_33341,N_33799);
nand U35838 (N_35838,N_33966,N_32645);
nor U35839 (N_35839,N_34080,N_34085);
and U35840 (N_35840,N_33972,N_32530);
or U35841 (N_35841,N_34571,N_33982);
xnor U35842 (N_35842,N_33713,N_34377);
and U35843 (N_35843,N_34681,N_34802);
or U35844 (N_35844,N_34762,N_34988);
nor U35845 (N_35845,N_32528,N_34165);
nand U35846 (N_35846,N_32693,N_34443);
nand U35847 (N_35847,N_33292,N_34042);
or U35848 (N_35848,N_34821,N_34575);
nand U35849 (N_35849,N_33257,N_33927);
and U35850 (N_35850,N_32989,N_33999);
xor U35851 (N_35851,N_33941,N_34374);
xor U35852 (N_35852,N_34927,N_34659);
nand U35853 (N_35853,N_33423,N_34614);
nand U35854 (N_35854,N_33057,N_33131);
or U35855 (N_35855,N_34361,N_34797);
nor U35856 (N_35856,N_34843,N_32542);
nand U35857 (N_35857,N_34737,N_34718);
nor U35858 (N_35858,N_33780,N_32840);
nor U35859 (N_35859,N_32866,N_33270);
nor U35860 (N_35860,N_34872,N_32625);
nand U35861 (N_35861,N_34850,N_33419);
and U35862 (N_35862,N_33540,N_33467);
nor U35863 (N_35863,N_32867,N_32588);
nor U35864 (N_35864,N_32669,N_34874);
nor U35865 (N_35865,N_34020,N_33056);
and U35866 (N_35866,N_33511,N_32587);
and U35867 (N_35867,N_33193,N_34160);
nor U35868 (N_35868,N_32943,N_33687);
or U35869 (N_35869,N_33273,N_34441);
nor U35870 (N_35870,N_33735,N_32799);
nor U35871 (N_35871,N_34199,N_34058);
xnor U35872 (N_35872,N_34204,N_33153);
nor U35873 (N_35873,N_33315,N_34703);
xor U35874 (N_35874,N_32788,N_33697);
and U35875 (N_35875,N_34633,N_33916);
and U35876 (N_35876,N_34846,N_33665);
xnor U35877 (N_35877,N_33896,N_32895);
nand U35878 (N_35878,N_33250,N_34209);
or U35879 (N_35879,N_32798,N_32950);
nor U35880 (N_35880,N_34738,N_33256);
xor U35881 (N_35881,N_32698,N_34844);
xnor U35882 (N_35882,N_34447,N_32660);
or U35883 (N_35883,N_34025,N_33964);
nand U35884 (N_35884,N_33897,N_32590);
nor U35885 (N_35885,N_32597,N_33488);
and U35886 (N_35886,N_33696,N_34516);
or U35887 (N_35887,N_34288,N_34217);
nor U35888 (N_35888,N_32987,N_33649);
and U35889 (N_35889,N_34492,N_32838);
or U35890 (N_35890,N_33061,N_33537);
nand U35891 (N_35891,N_34494,N_34051);
xnor U35892 (N_35892,N_34129,N_33160);
nor U35893 (N_35893,N_34422,N_32733);
and U35894 (N_35894,N_32629,N_34979);
xor U35895 (N_35895,N_32872,N_32906);
nand U35896 (N_35896,N_34078,N_34567);
or U35897 (N_35897,N_34240,N_34603);
xor U35898 (N_35898,N_33833,N_34983);
nand U35899 (N_35899,N_34982,N_32908);
nor U35900 (N_35900,N_33319,N_32991);
xnor U35901 (N_35901,N_33922,N_34987);
nand U35902 (N_35902,N_34444,N_34210);
nor U35903 (N_35903,N_33162,N_33347);
or U35904 (N_35904,N_33019,N_33358);
nor U35905 (N_35905,N_33141,N_34505);
xnor U35906 (N_35906,N_33958,N_33360);
and U35907 (N_35907,N_34859,N_33390);
nand U35908 (N_35908,N_34706,N_32508);
and U35909 (N_35909,N_33749,N_34271);
or U35910 (N_35910,N_34186,N_32683);
nand U35911 (N_35911,N_32819,N_34772);
nor U35912 (N_35912,N_33369,N_34445);
xor U35913 (N_35913,N_32721,N_34644);
and U35914 (N_35914,N_34518,N_33392);
or U35915 (N_35915,N_33052,N_34082);
or U35916 (N_35916,N_33626,N_32677);
or U35917 (N_35917,N_32935,N_33914);
and U35918 (N_35918,N_33264,N_33296);
and U35919 (N_35919,N_32554,N_33803);
nand U35920 (N_35920,N_34619,N_33113);
or U35921 (N_35921,N_33890,N_32883);
or U35922 (N_35922,N_34279,N_33835);
or U35923 (N_35923,N_34970,N_34289);
nand U35924 (N_35924,N_34649,N_34543);
nor U35925 (N_35925,N_33248,N_34876);
xnor U35926 (N_35926,N_32604,N_33326);
nand U35927 (N_35927,N_34232,N_33102);
nand U35928 (N_35928,N_33247,N_33674);
nor U35929 (N_35929,N_33552,N_34668);
nand U35930 (N_35930,N_33208,N_33509);
or U35931 (N_35931,N_33619,N_34753);
and U35932 (N_35932,N_34584,N_34594);
nand U35933 (N_35933,N_32593,N_34724);
nor U35934 (N_35934,N_34371,N_32662);
and U35935 (N_35935,N_34780,N_32876);
and U35936 (N_35936,N_34063,N_34473);
and U35937 (N_35937,N_34495,N_34468);
nand U35938 (N_35938,N_34489,N_34677);
nand U35939 (N_35939,N_32778,N_33209);
and U35940 (N_35940,N_33465,N_34766);
and U35941 (N_35941,N_33730,N_33891);
or U35942 (N_35942,N_32752,N_32532);
and U35943 (N_35943,N_34046,N_34946);
nand U35944 (N_35944,N_32548,N_34601);
xnor U35945 (N_35945,N_33715,N_34265);
and U35946 (N_35946,N_33011,N_33281);
nor U35947 (N_35947,N_34397,N_32891);
xnor U35948 (N_35948,N_33242,N_33961);
nand U35949 (N_35949,N_33703,N_34709);
or U35950 (N_35950,N_33769,N_33479);
and U35951 (N_35951,N_33919,N_34181);
and U35952 (N_35952,N_34754,N_33773);
or U35953 (N_35953,N_32627,N_33970);
and U35954 (N_35954,N_33359,N_33245);
xor U35955 (N_35955,N_33676,N_33759);
xnor U35956 (N_35956,N_32643,N_33807);
nor U35957 (N_35957,N_34143,N_32957);
nand U35958 (N_35958,N_33316,N_32607);
or U35959 (N_35959,N_33327,N_33238);
or U35960 (N_35960,N_33639,N_33771);
xor U35961 (N_35961,N_32531,N_33517);
and U35962 (N_35962,N_34017,N_33604);
xnor U35963 (N_35963,N_32509,N_32824);
nor U35964 (N_35964,N_34420,N_34015);
nand U35965 (N_35965,N_33348,N_34394);
nor U35966 (N_35966,N_32830,N_32921);
nand U35967 (N_35967,N_33279,N_34683);
nand U35968 (N_35968,N_32900,N_32735);
and U35969 (N_35969,N_34197,N_33291);
and U35970 (N_35970,N_33449,N_34686);
xor U35971 (N_35971,N_32826,N_32579);
nor U35972 (N_35972,N_34664,N_33241);
xor U35973 (N_35973,N_33913,N_33539);
nand U35974 (N_35974,N_34138,N_34404);
nand U35975 (N_35975,N_33388,N_33830);
nand U35976 (N_35976,N_33195,N_34966);
nor U35977 (N_35977,N_34920,N_34166);
or U35978 (N_35978,N_33006,N_34304);
and U35979 (N_35979,N_32801,N_34263);
nand U35980 (N_35980,N_33283,N_33048);
nand U35981 (N_35981,N_33269,N_33147);
nand U35982 (N_35982,N_34411,N_33079);
nor U35983 (N_35983,N_34139,N_33698);
nor U35984 (N_35984,N_34708,N_33608);
xnor U35985 (N_35985,N_34490,N_34955);
and U35986 (N_35986,N_33489,N_34880);
xor U35987 (N_35987,N_33161,N_34870);
nor U35988 (N_35988,N_33046,N_34196);
nand U35989 (N_35989,N_32868,N_34069);
xor U35990 (N_35990,N_33036,N_33929);
nor U35991 (N_35991,N_33159,N_34379);
and U35992 (N_35992,N_33122,N_34311);
nor U35993 (N_35993,N_34066,N_32846);
nor U35994 (N_35994,N_34929,N_33168);
and U35995 (N_35995,N_33770,N_33868);
and U35996 (N_35996,N_34280,N_32775);
nor U35997 (N_35997,N_33386,N_33028);
xnor U35998 (N_35998,N_32792,N_34555);
or U35999 (N_35999,N_33266,N_32765);
xor U36000 (N_36000,N_33553,N_33244);
nand U36001 (N_36001,N_33691,N_32511);
nor U36002 (N_36002,N_33956,N_32701);
and U36003 (N_36003,N_34965,N_34602);
or U36004 (N_36004,N_32708,N_32565);
or U36005 (N_36005,N_34147,N_33618);
nor U36006 (N_36006,N_33519,N_32719);
nand U36007 (N_36007,N_33781,N_33975);
and U36008 (N_36008,N_34035,N_33074);
nor U36009 (N_36009,N_34302,N_33843);
and U36010 (N_36010,N_34519,N_34693);
nand U36011 (N_36011,N_34720,N_34907);
nor U36012 (N_36012,N_34195,N_32952);
nor U36013 (N_36013,N_32615,N_32574);
xnor U36014 (N_36014,N_34450,N_34012);
or U36015 (N_36015,N_33725,N_34460);
nand U36016 (N_36016,N_34060,N_33993);
nor U36017 (N_36017,N_33794,N_34838);
xnor U36018 (N_36018,N_34549,N_33711);
xnor U36019 (N_36019,N_34651,N_33437);
or U36020 (N_36020,N_32761,N_33908);
nand U36021 (N_36021,N_33127,N_34178);
xor U36022 (N_36022,N_32576,N_33921);
xnor U36023 (N_36023,N_32828,N_33574);
xnor U36024 (N_36024,N_32707,N_33091);
nor U36025 (N_36025,N_32942,N_33402);
nor U36026 (N_36026,N_33094,N_34917);
nand U36027 (N_36027,N_33628,N_34981);
nor U36028 (N_36028,N_33952,N_32816);
nor U36029 (N_36029,N_32886,N_33850);
and U36030 (N_36030,N_33518,N_33481);
nand U36031 (N_36031,N_34047,N_33346);
or U36032 (N_36032,N_33690,N_34363);
nor U36033 (N_36033,N_34467,N_33349);
and U36034 (N_36034,N_34119,N_34480);
nand U36035 (N_36035,N_34676,N_32714);
nand U36036 (N_36036,N_34939,N_34036);
or U36037 (N_36037,N_34050,N_34714);
and U36038 (N_36038,N_33344,N_33002);
xor U36039 (N_36039,N_33946,N_34950);
nand U36040 (N_36040,N_32685,N_32793);
xor U36041 (N_36041,N_34026,N_32850);
nor U36042 (N_36042,N_33163,N_33310);
and U36043 (N_36043,N_33570,N_32668);
nand U36044 (N_36044,N_34383,N_33541);
xor U36045 (N_36045,N_33495,N_33073);
xor U36046 (N_36046,N_34790,N_32583);
xor U36047 (N_36047,N_34067,N_33923);
or U36048 (N_36048,N_34164,N_32539);
nor U36049 (N_36049,N_34170,N_32688);
nor U36050 (N_36050,N_34952,N_33635);
nor U36051 (N_36051,N_34735,N_32744);
and U36052 (N_36052,N_32834,N_33253);
xnor U36053 (N_36053,N_33267,N_34976);
or U36054 (N_36054,N_34239,N_34472);
nand U36055 (N_36055,N_32675,N_34785);
and U36056 (N_36056,N_34370,N_32753);
xor U36057 (N_36057,N_32762,N_34556);
and U36058 (N_36058,N_34918,N_32971);
xor U36059 (N_36059,N_32656,N_34412);
nand U36060 (N_36060,N_33904,N_33641);
xnor U36061 (N_36061,N_34152,N_34680);
xor U36062 (N_36062,N_33109,N_34257);
or U36063 (N_36063,N_32551,N_34320);
xor U36064 (N_36064,N_32573,N_34749);
or U36065 (N_36065,N_32839,N_33746);
xor U36066 (N_36066,N_32754,N_34530);
xor U36067 (N_36067,N_33523,N_33397);
and U36068 (N_36068,N_33116,N_32966);
nand U36069 (N_36069,N_34590,N_34953);
or U36070 (N_36070,N_33821,N_33085);
xnor U36071 (N_36071,N_32930,N_32559);
xnor U36072 (N_36072,N_34813,N_33520);
and U36073 (N_36073,N_33685,N_34888);
xor U36074 (N_36074,N_34906,N_33026);
nor U36075 (N_36075,N_33406,N_34548);
and U36076 (N_36076,N_32849,N_34174);
or U36077 (N_36077,N_34925,N_33931);
and U36078 (N_36078,N_34451,N_32679);
nand U36079 (N_36079,N_33186,N_33201);
xnor U36080 (N_36080,N_33078,N_34108);
nand U36081 (N_36081,N_32808,N_33263);
xnor U36082 (N_36082,N_32584,N_34733);
nand U36083 (N_36083,N_34074,N_33845);
xnor U36084 (N_36084,N_32730,N_33569);
xnor U36085 (N_36085,N_32896,N_34937);
xor U36086 (N_36086,N_33425,N_32892);
and U36087 (N_36087,N_32756,N_33150);
or U36088 (N_36088,N_33733,N_34410);
nand U36089 (N_36089,N_34801,N_32541);
nand U36090 (N_36090,N_32764,N_32696);
nor U36091 (N_36091,N_34822,N_33370);
or U36092 (N_36092,N_32732,N_33383);
nor U36093 (N_36093,N_34564,N_34717);
nand U36094 (N_36094,N_34747,N_32983);
nor U36095 (N_36095,N_33667,N_33090);
nor U36096 (N_36096,N_33668,N_33672);
and U36097 (N_36097,N_34118,N_34829);
nor U36098 (N_36098,N_33811,N_34301);
and U36099 (N_36099,N_33433,N_33320);
nand U36100 (N_36100,N_33831,N_34589);
and U36101 (N_36101,N_34796,N_33081);
xor U36102 (N_36102,N_33487,N_34462);
nor U36103 (N_36103,N_33809,N_32591);
nand U36104 (N_36104,N_33440,N_33995);
or U36105 (N_36105,N_33550,N_34980);
and U36106 (N_36106,N_34520,N_34741);
nand U36107 (N_36107,N_34207,N_34083);
xnor U36108 (N_36108,N_32986,N_34690);
nor U36109 (N_36109,N_32785,N_34728);
nand U36110 (N_36110,N_34115,N_34942);
and U36111 (N_36111,N_34687,N_34635);
or U36112 (N_36112,N_33169,N_33784);
xnor U36113 (N_36113,N_34481,N_34073);
nand U36114 (N_36114,N_33412,N_33087);
nand U36115 (N_36115,N_34203,N_34446);
and U36116 (N_36116,N_34643,N_32522);
and U36117 (N_36117,N_34434,N_34172);
or U36118 (N_36118,N_33205,N_32955);
xor U36119 (N_36119,N_34104,N_32556);
nor U36120 (N_36120,N_32856,N_34225);
and U36121 (N_36121,N_33024,N_34223);
nand U36122 (N_36122,N_34227,N_32603);
xor U36123 (N_36123,N_34898,N_34233);
nand U36124 (N_36124,N_32637,N_34076);
or U36125 (N_36125,N_33228,N_32536);
and U36126 (N_36126,N_33062,N_33458);
and U36127 (N_36127,N_34243,N_33404);
and U36128 (N_36128,N_34597,N_33422);
nand U36129 (N_36129,N_32692,N_34861);
nand U36130 (N_36130,N_33849,N_33726);
xnor U36131 (N_36131,N_33373,N_33086);
and U36132 (N_36132,N_32575,N_32847);
or U36133 (N_36133,N_33516,N_33951);
nand U36134 (N_36134,N_34512,N_33429);
xnor U36135 (N_36135,N_32790,N_34039);
or U36136 (N_36136,N_34847,N_34216);
xnor U36137 (N_36137,N_33813,N_33556);
nand U36138 (N_36138,N_34782,N_33743);
or U36139 (N_36139,N_34778,N_33138);
xnor U36140 (N_36140,N_34011,N_32870);
xor U36141 (N_36141,N_33045,N_34631);
and U36142 (N_36142,N_33175,N_34775);
and U36143 (N_36143,N_34326,N_34574);
nand U36144 (N_36144,N_32610,N_33870);
and U36145 (N_36145,N_32897,N_32909);
or U36146 (N_36146,N_32822,N_34096);
xor U36147 (N_36147,N_33768,N_33058);
or U36148 (N_36148,N_32852,N_32855);
or U36149 (N_36149,N_34612,N_33855);
nand U36150 (N_36150,N_33474,N_34864);
and U36151 (N_36151,N_33571,N_32608);
nor U36152 (N_36152,N_34019,N_33874);
nor U36153 (N_36153,N_34275,N_33859);
xor U36154 (N_36154,N_34610,N_33812);
or U36155 (N_36155,N_34609,N_33723);
or U36156 (N_36156,N_33416,N_34264);
nor U36157 (N_36157,N_34868,N_33663);
nor U36158 (N_36158,N_34001,N_34752);
nor U36159 (N_36159,N_34013,N_33287);
xor U36160 (N_36160,N_33414,N_33942);
nor U36161 (N_36161,N_34940,N_33755);
xnor U36162 (N_36162,N_33719,N_33494);
xnor U36163 (N_36163,N_33149,N_33988);
nor U36164 (N_36164,N_33774,N_33577);
xor U36165 (N_36165,N_33194,N_34879);
nor U36166 (N_36166,N_34247,N_33503);
and U36167 (N_36167,N_33504,N_33473);
nand U36168 (N_36168,N_33451,N_34698);
or U36169 (N_36169,N_32740,N_33300);
nand U36170 (N_36170,N_34948,N_32887);
or U36171 (N_36171,N_34122,N_33200);
and U36172 (N_36172,N_32750,N_33135);
nor U36173 (N_36173,N_34106,N_34973);
xor U36174 (N_36174,N_33684,N_34732);
or U36175 (N_36175,N_34340,N_32543);
nand U36176 (N_36176,N_34682,N_34345);
nand U36177 (N_36177,N_33990,N_33428);
and U36178 (N_36178,N_33220,N_34611);
nor U36179 (N_36179,N_32739,N_34931);
or U36180 (N_36180,N_33878,N_32969);
and U36181 (N_36181,N_33114,N_33145);
or U36182 (N_36182,N_33272,N_34323);
or U36183 (N_36183,N_33514,N_33793);
nand U36184 (N_36184,N_34587,N_33064);
and U36185 (N_36185,N_32569,N_32659);
nand U36186 (N_36186,N_34369,N_34816);
xnor U36187 (N_36187,N_34873,N_32854);
xnor U36188 (N_36188,N_33601,N_33179);
nor U36189 (N_36189,N_33527,N_32848);
xnor U36190 (N_36190,N_34501,N_34558);
nand U36191 (N_36191,N_33130,N_33638);
and U36192 (N_36192,N_33598,N_32975);
nand U36193 (N_36193,N_33352,N_33860);
nor U36194 (N_36194,N_34182,N_34776);
or U36195 (N_36195,N_34875,N_33132);
and U36196 (N_36196,N_34617,N_34725);
nor U36197 (N_36197,N_34094,N_32553);
and U36198 (N_36198,N_33271,N_33721);
xnor U36199 (N_36199,N_34262,N_32763);
and U36200 (N_36200,N_34246,N_34851);
and U36201 (N_36201,N_34666,N_32723);
nand U36202 (N_36202,N_33077,N_34826);
nand U36203 (N_36203,N_33218,N_33184);
nor U36204 (N_36204,N_34961,N_34465);
or U36205 (N_36205,N_34788,N_32605);
or U36206 (N_36206,N_33453,N_34110);
xor U36207 (N_36207,N_32609,N_34921);
and U36208 (N_36208,N_34623,N_34387);
nand U36209 (N_36209,N_34487,N_33892);
and U36210 (N_36210,N_33957,N_33233);
nor U36211 (N_36211,N_32910,N_34713);
nor U36212 (N_36212,N_34592,N_34030);
xor U36213 (N_36213,N_34293,N_32726);
xnor U36214 (N_36214,N_34366,N_33365);
and U36215 (N_36215,N_34109,N_34865);
nand U36216 (N_36216,N_33441,N_34761);
nor U36217 (N_36217,N_34656,N_33840);
nand U36218 (N_36218,N_34200,N_33654);
xor U36219 (N_36219,N_33662,N_33532);
xnor U36220 (N_36220,N_32836,N_33005);
xor U36221 (N_36221,N_34892,N_34991);
nand U36222 (N_36222,N_33867,N_34560);
or U36223 (N_36223,N_33854,N_33117);
or U36224 (N_36224,N_33082,N_33120);
nand U36225 (N_36225,N_34989,N_34591);
or U36226 (N_36226,N_33421,N_33836);
or U36227 (N_36227,N_33804,N_33655);
or U36228 (N_36228,N_34103,N_34317);
or U36229 (N_36229,N_33427,N_34757);
or U36230 (N_36230,N_34090,N_33572);
or U36231 (N_36231,N_33174,N_32948);
nor U36232 (N_36232,N_33054,N_32820);
and U36233 (N_36233,N_33463,N_34514);
and U36234 (N_36234,N_33004,N_33372);
nor U36235 (N_36235,N_34332,N_32557);
xor U36236 (N_36236,N_33911,N_33396);
xnor U36237 (N_36237,N_33513,N_34180);
nor U36238 (N_36238,N_33605,N_34928);
xor U36239 (N_36239,N_32776,N_33851);
nor U36240 (N_36240,N_33112,N_32736);
nand U36241 (N_36241,N_34388,N_33008);
or U36242 (N_36242,N_32980,N_32503);
or U36243 (N_36243,N_32621,N_34220);
xnor U36244 (N_36244,N_34027,N_34127);
nand U36245 (N_36245,N_32968,N_33146);
xor U36246 (N_36246,N_32545,N_33198);
and U36247 (N_36247,N_32976,N_33787);
or U36248 (N_36248,N_33592,N_33183);
xnor U36249 (N_36249,N_32564,N_32517);
nand U36250 (N_36250,N_33733,N_33033);
and U36251 (N_36251,N_34760,N_32552);
nor U36252 (N_36252,N_34396,N_33415);
xnor U36253 (N_36253,N_34900,N_33388);
xor U36254 (N_36254,N_32919,N_33554);
and U36255 (N_36255,N_34943,N_32918);
or U36256 (N_36256,N_33767,N_32842);
or U36257 (N_36257,N_34296,N_33384);
nand U36258 (N_36258,N_33658,N_32929);
xor U36259 (N_36259,N_33576,N_34189);
or U36260 (N_36260,N_33832,N_32719);
nand U36261 (N_36261,N_32774,N_34868);
xor U36262 (N_36262,N_34093,N_33807);
nor U36263 (N_36263,N_34694,N_33967);
xnor U36264 (N_36264,N_34835,N_32623);
xor U36265 (N_36265,N_34455,N_34734);
and U36266 (N_36266,N_32581,N_34168);
and U36267 (N_36267,N_32774,N_34197);
or U36268 (N_36268,N_34925,N_33836);
and U36269 (N_36269,N_32514,N_34336);
nand U36270 (N_36270,N_34524,N_33370);
or U36271 (N_36271,N_33626,N_34268);
xor U36272 (N_36272,N_33648,N_33095);
nand U36273 (N_36273,N_33274,N_34761);
nand U36274 (N_36274,N_34555,N_33906);
and U36275 (N_36275,N_33871,N_33417);
nor U36276 (N_36276,N_33220,N_32715);
xnor U36277 (N_36277,N_33130,N_33886);
nor U36278 (N_36278,N_33141,N_33581);
nor U36279 (N_36279,N_32702,N_33443);
nor U36280 (N_36280,N_33878,N_33874);
nor U36281 (N_36281,N_34037,N_32502);
and U36282 (N_36282,N_34630,N_33240);
nand U36283 (N_36283,N_32571,N_34904);
nor U36284 (N_36284,N_34401,N_34442);
nand U36285 (N_36285,N_34015,N_32971);
xor U36286 (N_36286,N_33421,N_34459);
xor U36287 (N_36287,N_32964,N_34938);
nand U36288 (N_36288,N_33170,N_34521);
and U36289 (N_36289,N_32878,N_34805);
or U36290 (N_36290,N_32764,N_32875);
nor U36291 (N_36291,N_32629,N_34811);
nor U36292 (N_36292,N_34789,N_32773);
nand U36293 (N_36293,N_34700,N_34156);
or U36294 (N_36294,N_34466,N_33630);
or U36295 (N_36295,N_32850,N_32600);
xor U36296 (N_36296,N_33459,N_32675);
nor U36297 (N_36297,N_33326,N_33576);
nand U36298 (N_36298,N_34610,N_34140);
nand U36299 (N_36299,N_33720,N_33761);
nor U36300 (N_36300,N_34984,N_34790);
and U36301 (N_36301,N_34637,N_34650);
xor U36302 (N_36302,N_34691,N_32955);
nor U36303 (N_36303,N_34896,N_34747);
or U36304 (N_36304,N_33946,N_34932);
or U36305 (N_36305,N_33528,N_33960);
nor U36306 (N_36306,N_33668,N_33435);
and U36307 (N_36307,N_33478,N_34348);
and U36308 (N_36308,N_34495,N_34711);
or U36309 (N_36309,N_33436,N_33726);
xnor U36310 (N_36310,N_34504,N_33505);
nor U36311 (N_36311,N_34805,N_33998);
nor U36312 (N_36312,N_32781,N_33511);
and U36313 (N_36313,N_32911,N_33074);
or U36314 (N_36314,N_33594,N_33429);
nor U36315 (N_36315,N_34468,N_34146);
nand U36316 (N_36316,N_33235,N_34103);
xnor U36317 (N_36317,N_34157,N_33272);
or U36318 (N_36318,N_34922,N_32571);
xnor U36319 (N_36319,N_33350,N_33669);
nand U36320 (N_36320,N_33149,N_34693);
and U36321 (N_36321,N_33240,N_32683);
and U36322 (N_36322,N_34516,N_33300);
nand U36323 (N_36323,N_34967,N_34038);
and U36324 (N_36324,N_33547,N_33326);
nand U36325 (N_36325,N_34490,N_32843);
nor U36326 (N_36326,N_33844,N_33808);
and U36327 (N_36327,N_33167,N_34333);
or U36328 (N_36328,N_34231,N_33888);
nand U36329 (N_36329,N_33311,N_32613);
and U36330 (N_36330,N_32936,N_33039);
nand U36331 (N_36331,N_34697,N_33528);
xnor U36332 (N_36332,N_34280,N_34009);
nor U36333 (N_36333,N_34873,N_33113);
xnor U36334 (N_36334,N_33478,N_34550);
or U36335 (N_36335,N_34523,N_34189);
or U36336 (N_36336,N_33705,N_33624);
and U36337 (N_36337,N_32993,N_34474);
xor U36338 (N_36338,N_32710,N_34486);
nor U36339 (N_36339,N_34022,N_34957);
and U36340 (N_36340,N_34968,N_33811);
xnor U36341 (N_36341,N_33216,N_34971);
and U36342 (N_36342,N_33995,N_34459);
or U36343 (N_36343,N_34739,N_34211);
nand U36344 (N_36344,N_33984,N_34512);
or U36345 (N_36345,N_33812,N_32562);
xnor U36346 (N_36346,N_33424,N_34132);
or U36347 (N_36347,N_32662,N_33405);
nor U36348 (N_36348,N_34874,N_32726);
nand U36349 (N_36349,N_33945,N_34844);
or U36350 (N_36350,N_34324,N_32624);
xor U36351 (N_36351,N_33103,N_33569);
or U36352 (N_36352,N_34704,N_34785);
and U36353 (N_36353,N_34293,N_33870);
xnor U36354 (N_36354,N_34443,N_33922);
xnor U36355 (N_36355,N_34271,N_33689);
and U36356 (N_36356,N_33928,N_34740);
nand U36357 (N_36357,N_34016,N_33568);
xor U36358 (N_36358,N_33154,N_33445);
nand U36359 (N_36359,N_32666,N_33527);
nor U36360 (N_36360,N_34263,N_34944);
xnor U36361 (N_36361,N_33076,N_32506);
and U36362 (N_36362,N_33581,N_33212);
nor U36363 (N_36363,N_33078,N_34888);
nand U36364 (N_36364,N_32659,N_33076);
xnor U36365 (N_36365,N_32892,N_33013);
or U36366 (N_36366,N_32824,N_33012);
or U36367 (N_36367,N_32698,N_33505);
or U36368 (N_36368,N_33197,N_33050);
or U36369 (N_36369,N_33690,N_33110);
xor U36370 (N_36370,N_32909,N_33031);
nor U36371 (N_36371,N_34190,N_32546);
or U36372 (N_36372,N_32969,N_32884);
nand U36373 (N_36373,N_33926,N_34080);
and U36374 (N_36374,N_32926,N_34626);
nor U36375 (N_36375,N_33342,N_32835);
xnor U36376 (N_36376,N_32523,N_34130);
nand U36377 (N_36377,N_32754,N_32799);
or U36378 (N_36378,N_33816,N_34945);
xnor U36379 (N_36379,N_34273,N_34173);
or U36380 (N_36380,N_34928,N_34484);
nand U36381 (N_36381,N_33519,N_32998);
nor U36382 (N_36382,N_34893,N_32770);
and U36383 (N_36383,N_32612,N_33479);
and U36384 (N_36384,N_33622,N_32900);
nor U36385 (N_36385,N_32933,N_34123);
or U36386 (N_36386,N_34722,N_32535);
or U36387 (N_36387,N_34866,N_32891);
or U36388 (N_36388,N_33538,N_32946);
nand U36389 (N_36389,N_34876,N_32899);
nand U36390 (N_36390,N_33004,N_33657);
xnor U36391 (N_36391,N_33151,N_34461);
nor U36392 (N_36392,N_33212,N_34678);
nor U36393 (N_36393,N_33924,N_33667);
nand U36394 (N_36394,N_33152,N_34372);
xnor U36395 (N_36395,N_33707,N_32565);
and U36396 (N_36396,N_32881,N_34733);
xnor U36397 (N_36397,N_34540,N_34063);
nor U36398 (N_36398,N_32515,N_32530);
or U36399 (N_36399,N_32572,N_33112);
nor U36400 (N_36400,N_34966,N_33740);
or U36401 (N_36401,N_34067,N_34948);
or U36402 (N_36402,N_33905,N_33862);
nand U36403 (N_36403,N_34749,N_32742);
nand U36404 (N_36404,N_33335,N_33837);
xnor U36405 (N_36405,N_33515,N_33129);
and U36406 (N_36406,N_33886,N_34990);
xor U36407 (N_36407,N_34869,N_34247);
and U36408 (N_36408,N_34415,N_32984);
xnor U36409 (N_36409,N_34959,N_33998);
and U36410 (N_36410,N_33777,N_33250);
nand U36411 (N_36411,N_34595,N_33737);
and U36412 (N_36412,N_33149,N_33579);
nor U36413 (N_36413,N_34215,N_33751);
and U36414 (N_36414,N_34809,N_34407);
nor U36415 (N_36415,N_33034,N_34217);
nor U36416 (N_36416,N_33799,N_34063);
xor U36417 (N_36417,N_34139,N_32797);
nand U36418 (N_36418,N_34098,N_33673);
nand U36419 (N_36419,N_34884,N_33502);
nor U36420 (N_36420,N_34124,N_32784);
or U36421 (N_36421,N_32905,N_33098);
nor U36422 (N_36422,N_33074,N_33002);
nor U36423 (N_36423,N_32521,N_33095);
or U36424 (N_36424,N_33106,N_33952);
or U36425 (N_36425,N_34464,N_33287);
nor U36426 (N_36426,N_34324,N_32585);
and U36427 (N_36427,N_34864,N_33297);
xnor U36428 (N_36428,N_32840,N_33685);
and U36429 (N_36429,N_33283,N_34804);
or U36430 (N_36430,N_34957,N_33033);
or U36431 (N_36431,N_33550,N_34308);
or U36432 (N_36432,N_32741,N_32754);
xor U36433 (N_36433,N_34945,N_33323);
nor U36434 (N_36434,N_32658,N_34874);
nand U36435 (N_36435,N_32868,N_34477);
nor U36436 (N_36436,N_34918,N_33200);
and U36437 (N_36437,N_33803,N_34252);
xnor U36438 (N_36438,N_33666,N_34346);
and U36439 (N_36439,N_32500,N_34711);
nor U36440 (N_36440,N_33354,N_34311);
or U36441 (N_36441,N_33702,N_32775);
or U36442 (N_36442,N_33015,N_34723);
nor U36443 (N_36443,N_34219,N_34315);
or U36444 (N_36444,N_32809,N_33853);
nor U36445 (N_36445,N_34722,N_33560);
nand U36446 (N_36446,N_33861,N_32906);
nand U36447 (N_36447,N_34341,N_34893);
or U36448 (N_36448,N_34756,N_33806);
and U36449 (N_36449,N_34492,N_34102);
and U36450 (N_36450,N_34834,N_32702);
and U36451 (N_36451,N_33336,N_33407);
nand U36452 (N_36452,N_33591,N_34541);
nand U36453 (N_36453,N_34685,N_33098);
and U36454 (N_36454,N_34791,N_34269);
and U36455 (N_36455,N_34760,N_33507);
and U36456 (N_36456,N_33547,N_33671);
and U36457 (N_36457,N_34642,N_34569);
or U36458 (N_36458,N_34035,N_32774);
or U36459 (N_36459,N_33569,N_34086);
nor U36460 (N_36460,N_32719,N_34158);
nand U36461 (N_36461,N_34410,N_32993);
nand U36462 (N_36462,N_33124,N_33322);
xor U36463 (N_36463,N_34050,N_34637);
and U36464 (N_36464,N_32974,N_34981);
nor U36465 (N_36465,N_32952,N_33040);
nor U36466 (N_36466,N_34325,N_33264);
xnor U36467 (N_36467,N_32778,N_34435);
xnor U36468 (N_36468,N_33466,N_33791);
or U36469 (N_36469,N_34068,N_33129);
nor U36470 (N_36470,N_34478,N_33903);
xnor U36471 (N_36471,N_33193,N_33782);
or U36472 (N_36472,N_34794,N_34839);
nand U36473 (N_36473,N_34907,N_34690);
xor U36474 (N_36474,N_32519,N_34236);
xor U36475 (N_36475,N_33318,N_33174);
nor U36476 (N_36476,N_33725,N_33355);
nor U36477 (N_36477,N_34554,N_33499);
nand U36478 (N_36478,N_32811,N_33890);
nor U36479 (N_36479,N_33042,N_34025);
and U36480 (N_36480,N_32671,N_32629);
xor U36481 (N_36481,N_33863,N_34358);
nand U36482 (N_36482,N_33413,N_33804);
nor U36483 (N_36483,N_32683,N_32700);
nor U36484 (N_36484,N_34272,N_33417);
nor U36485 (N_36485,N_34767,N_34955);
or U36486 (N_36486,N_33049,N_33316);
xnor U36487 (N_36487,N_32504,N_34396);
or U36488 (N_36488,N_34892,N_33763);
nor U36489 (N_36489,N_33226,N_34436);
nor U36490 (N_36490,N_32997,N_33316);
xnor U36491 (N_36491,N_34812,N_32686);
xnor U36492 (N_36492,N_33187,N_33870);
nand U36493 (N_36493,N_32799,N_33689);
nor U36494 (N_36494,N_33051,N_33510);
and U36495 (N_36495,N_34097,N_34553);
nand U36496 (N_36496,N_34712,N_34539);
or U36497 (N_36497,N_34810,N_34802);
xnor U36498 (N_36498,N_32735,N_34260);
or U36499 (N_36499,N_34040,N_34961);
or U36500 (N_36500,N_33274,N_33470);
xnor U36501 (N_36501,N_34196,N_34867);
or U36502 (N_36502,N_33109,N_33319);
or U36503 (N_36503,N_32673,N_34938);
xnor U36504 (N_36504,N_32539,N_33514);
or U36505 (N_36505,N_33993,N_33689);
xnor U36506 (N_36506,N_34797,N_34272);
or U36507 (N_36507,N_34701,N_33763);
xor U36508 (N_36508,N_34481,N_32996);
or U36509 (N_36509,N_33423,N_34127);
xnor U36510 (N_36510,N_32971,N_33924);
and U36511 (N_36511,N_33700,N_33419);
nand U36512 (N_36512,N_33445,N_32864);
and U36513 (N_36513,N_33302,N_33876);
nor U36514 (N_36514,N_33382,N_33213);
nor U36515 (N_36515,N_34933,N_33773);
or U36516 (N_36516,N_34259,N_33122);
nand U36517 (N_36517,N_34176,N_34373);
and U36518 (N_36518,N_32613,N_32961);
or U36519 (N_36519,N_34930,N_34583);
nand U36520 (N_36520,N_33790,N_33076);
nor U36521 (N_36521,N_34923,N_33967);
and U36522 (N_36522,N_34718,N_33845);
xnor U36523 (N_36523,N_34792,N_32927);
nand U36524 (N_36524,N_32731,N_34959);
nor U36525 (N_36525,N_32693,N_34188);
and U36526 (N_36526,N_34231,N_32832);
and U36527 (N_36527,N_34521,N_34544);
or U36528 (N_36528,N_33449,N_33863);
nand U36529 (N_36529,N_33344,N_33090);
nor U36530 (N_36530,N_34676,N_32630);
nor U36531 (N_36531,N_33057,N_32704);
nor U36532 (N_36532,N_34994,N_34314);
or U36533 (N_36533,N_34171,N_34433);
or U36534 (N_36534,N_32809,N_32505);
nor U36535 (N_36535,N_34861,N_34709);
nand U36536 (N_36536,N_33609,N_34159);
or U36537 (N_36537,N_32832,N_34842);
and U36538 (N_36538,N_32717,N_34114);
nand U36539 (N_36539,N_33362,N_33963);
xnor U36540 (N_36540,N_34304,N_32694);
or U36541 (N_36541,N_34337,N_33302);
xor U36542 (N_36542,N_34820,N_33468);
or U36543 (N_36543,N_34834,N_34351);
or U36544 (N_36544,N_34801,N_33469);
or U36545 (N_36545,N_34789,N_33024);
nand U36546 (N_36546,N_33409,N_34655);
nor U36547 (N_36547,N_33163,N_32581);
and U36548 (N_36548,N_33648,N_34440);
xnor U36549 (N_36549,N_34902,N_34418);
and U36550 (N_36550,N_34661,N_32718);
and U36551 (N_36551,N_32542,N_33062);
nor U36552 (N_36552,N_32688,N_34066);
nand U36553 (N_36553,N_32961,N_33593);
or U36554 (N_36554,N_34711,N_33883);
or U36555 (N_36555,N_32656,N_33657);
or U36556 (N_36556,N_33810,N_34087);
nor U36557 (N_36557,N_34161,N_34692);
and U36558 (N_36558,N_34445,N_33103);
xnor U36559 (N_36559,N_34923,N_34919);
xnor U36560 (N_36560,N_34497,N_32565);
or U36561 (N_36561,N_34916,N_33763);
xor U36562 (N_36562,N_34001,N_33977);
nor U36563 (N_36563,N_34733,N_34683);
nor U36564 (N_36564,N_33863,N_34874);
or U36565 (N_36565,N_32837,N_33937);
or U36566 (N_36566,N_33312,N_34552);
or U36567 (N_36567,N_32697,N_34543);
nand U36568 (N_36568,N_34744,N_32946);
nor U36569 (N_36569,N_33253,N_33950);
or U36570 (N_36570,N_34013,N_32813);
or U36571 (N_36571,N_34525,N_34791);
nand U36572 (N_36572,N_32656,N_32645);
xnor U36573 (N_36573,N_34392,N_33005);
or U36574 (N_36574,N_34727,N_33901);
nor U36575 (N_36575,N_32807,N_34680);
or U36576 (N_36576,N_34100,N_32517);
nor U36577 (N_36577,N_34867,N_33523);
xnor U36578 (N_36578,N_33682,N_32519);
nand U36579 (N_36579,N_32749,N_34490);
or U36580 (N_36580,N_33113,N_34616);
nor U36581 (N_36581,N_33862,N_34828);
nand U36582 (N_36582,N_32794,N_32637);
nor U36583 (N_36583,N_33676,N_33070);
or U36584 (N_36584,N_33311,N_33854);
xor U36585 (N_36585,N_34582,N_33427);
nor U36586 (N_36586,N_34008,N_33743);
xor U36587 (N_36587,N_32935,N_33188);
nand U36588 (N_36588,N_33096,N_33212);
and U36589 (N_36589,N_34312,N_32815);
nor U36590 (N_36590,N_34291,N_33526);
nor U36591 (N_36591,N_34822,N_33971);
nor U36592 (N_36592,N_34023,N_34869);
xnor U36593 (N_36593,N_34453,N_34617);
and U36594 (N_36594,N_33634,N_34385);
xor U36595 (N_36595,N_34891,N_34729);
xnor U36596 (N_36596,N_34175,N_34141);
nand U36597 (N_36597,N_33070,N_34897);
nand U36598 (N_36598,N_34868,N_34201);
or U36599 (N_36599,N_33619,N_34573);
and U36600 (N_36600,N_34629,N_33143);
and U36601 (N_36601,N_32793,N_32701);
nor U36602 (N_36602,N_33593,N_34703);
or U36603 (N_36603,N_33252,N_34653);
nor U36604 (N_36604,N_34554,N_32986);
and U36605 (N_36605,N_34962,N_33771);
xnor U36606 (N_36606,N_34762,N_32966);
and U36607 (N_36607,N_33003,N_32732);
xor U36608 (N_36608,N_33345,N_34068);
or U36609 (N_36609,N_32929,N_32548);
nand U36610 (N_36610,N_33747,N_34599);
or U36611 (N_36611,N_33055,N_32978);
nor U36612 (N_36612,N_34137,N_32591);
nand U36613 (N_36613,N_34070,N_33613);
nor U36614 (N_36614,N_34691,N_34078);
nor U36615 (N_36615,N_34926,N_34738);
nor U36616 (N_36616,N_32609,N_33777);
nor U36617 (N_36617,N_33486,N_34377);
nor U36618 (N_36618,N_33658,N_34527);
xor U36619 (N_36619,N_33033,N_34877);
and U36620 (N_36620,N_33849,N_34466);
xor U36621 (N_36621,N_32616,N_33082);
xnor U36622 (N_36622,N_32930,N_34078);
or U36623 (N_36623,N_33329,N_33245);
or U36624 (N_36624,N_34156,N_34347);
or U36625 (N_36625,N_32527,N_33460);
nor U36626 (N_36626,N_32841,N_32763);
nand U36627 (N_36627,N_33121,N_34317);
nand U36628 (N_36628,N_34579,N_34352);
or U36629 (N_36629,N_33913,N_34364);
xor U36630 (N_36630,N_34450,N_32877);
and U36631 (N_36631,N_33178,N_34493);
nor U36632 (N_36632,N_33521,N_33128);
nand U36633 (N_36633,N_34862,N_34579);
xor U36634 (N_36634,N_34094,N_32802);
and U36635 (N_36635,N_33739,N_34357);
nand U36636 (N_36636,N_34243,N_33457);
nor U36637 (N_36637,N_32657,N_34321);
nand U36638 (N_36638,N_33978,N_32873);
xor U36639 (N_36639,N_34186,N_34398);
or U36640 (N_36640,N_33021,N_33617);
and U36641 (N_36641,N_33064,N_33436);
or U36642 (N_36642,N_34938,N_33661);
nand U36643 (N_36643,N_32718,N_32932);
and U36644 (N_36644,N_33141,N_33858);
and U36645 (N_36645,N_32896,N_33949);
or U36646 (N_36646,N_32560,N_33999);
or U36647 (N_36647,N_34734,N_32501);
or U36648 (N_36648,N_33663,N_33752);
and U36649 (N_36649,N_33118,N_34869);
or U36650 (N_36650,N_34664,N_33489);
nor U36651 (N_36651,N_32888,N_33215);
nand U36652 (N_36652,N_33898,N_33472);
nand U36653 (N_36653,N_32631,N_32609);
or U36654 (N_36654,N_32520,N_32655);
and U36655 (N_36655,N_34385,N_34166);
xor U36656 (N_36656,N_32790,N_32883);
or U36657 (N_36657,N_34789,N_32985);
and U36658 (N_36658,N_34352,N_34730);
and U36659 (N_36659,N_34582,N_34338);
xor U36660 (N_36660,N_33650,N_33426);
nand U36661 (N_36661,N_34368,N_34047);
xor U36662 (N_36662,N_32862,N_32857);
nor U36663 (N_36663,N_34678,N_33742);
nor U36664 (N_36664,N_33155,N_34566);
xnor U36665 (N_36665,N_34895,N_33739);
and U36666 (N_36666,N_33824,N_32742);
xor U36667 (N_36667,N_34751,N_32784);
and U36668 (N_36668,N_32855,N_32635);
nor U36669 (N_36669,N_34579,N_33699);
or U36670 (N_36670,N_34215,N_34273);
and U36671 (N_36671,N_33536,N_34762);
or U36672 (N_36672,N_34329,N_33648);
nand U36673 (N_36673,N_33716,N_32627);
xor U36674 (N_36674,N_32873,N_32761);
xor U36675 (N_36675,N_32631,N_34530);
nand U36676 (N_36676,N_32998,N_32838);
or U36677 (N_36677,N_33088,N_34077);
nand U36678 (N_36678,N_32659,N_32916);
xnor U36679 (N_36679,N_33392,N_32892);
xor U36680 (N_36680,N_34977,N_33410);
or U36681 (N_36681,N_33807,N_33473);
or U36682 (N_36682,N_34965,N_33406);
and U36683 (N_36683,N_33376,N_32600);
nor U36684 (N_36684,N_34846,N_32707);
and U36685 (N_36685,N_33493,N_33604);
xor U36686 (N_36686,N_33434,N_32925);
nand U36687 (N_36687,N_34839,N_34155);
xor U36688 (N_36688,N_33031,N_32927);
nand U36689 (N_36689,N_32760,N_34250);
xor U36690 (N_36690,N_34346,N_33118);
nand U36691 (N_36691,N_34644,N_32799);
or U36692 (N_36692,N_32713,N_34691);
nand U36693 (N_36693,N_32542,N_34371);
nand U36694 (N_36694,N_34161,N_33680);
nor U36695 (N_36695,N_33787,N_33065);
nor U36696 (N_36696,N_33148,N_33228);
nor U36697 (N_36697,N_34018,N_33940);
or U36698 (N_36698,N_33674,N_32733);
nor U36699 (N_36699,N_32677,N_33962);
nand U36700 (N_36700,N_32529,N_33991);
xnor U36701 (N_36701,N_34846,N_33699);
nand U36702 (N_36702,N_33773,N_34328);
or U36703 (N_36703,N_34849,N_34118);
nor U36704 (N_36704,N_33796,N_33067);
nand U36705 (N_36705,N_33534,N_32663);
nor U36706 (N_36706,N_34412,N_34213);
nor U36707 (N_36707,N_33198,N_33554);
or U36708 (N_36708,N_33269,N_33704);
nand U36709 (N_36709,N_33909,N_33139);
and U36710 (N_36710,N_33436,N_34200);
nand U36711 (N_36711,N_32746,N_34022);
or U36712 (N_36712,N_34781,N_34816);
and U36713 (N_36713,N_33595,N_33945);
and U36714 (N_36714,N_33257,N_34133);
xor U36715 (N_36715,N_34322,N_33627);
xnor U36716 (N_36716,N_33185,N_34913);
nand U36717 (N_36717,N_34588,N_34524);
or U36718 (N_36718,N_34898,N_33983);
nand U36719 (N_36719,N_33995,N_34007);
nand U36720 (N_36720,N_34454,N_34129);
nor U36721 (N_36721,N_33155,N_34730);
nor U36722 (N_36722,N_34688,N_33831);
nor U36723 (N_36723,N_34202,N_33420);
and U36724 (N_36724,N_34430,N_33514);
xnor U36725 (N_36725,N_32783,N_32812);
xor U36726 (N_36726,N_33437,N_33199);
or U36727 (N_36727,N_32825,N_33677);
nor U36728 (N_36728,N_32996,N_34763);
nor U36729 (N_36729,N_33936,N_33464);
nor U36730 (N_36730,N_34042,N_34938);
and U36731 (N_36731,N_34876,N_33352);
nor U36732 (N_36732,N_33373,N_32891);
xnor U36733 (N_36733,N_34533,N_33363);
and U36734 (N_36734,N_34007,N_33440);
nand U36735 (N_36735,N_33705,N_34483);
xnor U36736 (N_36736,N_33243,N_34860);
nand U36737 (N_36737,N_34194,N_34311);
xnor U36738 (N_36738,N_33187,N_34442);
nand U36739 (N_36739,N_32833,N_34895);
and U36740 (N_36740,N_32910,N_33059);
and U36741 (N_36741,N_33766,N_33099);
nand U36742 (N_36742,N_33160,N_32524);
nand U36743 (N_36743,N_34057,N_34264);
or U36744 (N_36744,N_32971,N_32569);
xor U36745 (N_36745,N_34312,N_33609);
xnor U36746 (N_36746,N_33562,N_33034);
xnor U36747 (N_36747,N_32759,N_33824);
and U36748 (N_36748,N_34691,N_34528);
nor U36749 (N_36749,N_33372,N_33743);
and U36750 (N_36750,N_32644,N_34182);
nor U36751 (N_36751,N_34397,N_34228);
nand U36752 (N_36752,N_34116,N_32703);
or U36753 (N_36753,N_34110,N_34869);
nand U36754 (N_36754,N_34313,N_33602);
nor U36755 (N_36755,N_34125,N_34220);
nor U36756 (N_36756,N_34552,N_33593);
xnor U36757 (N_36757,N_33951,N_33232);
nand U36758 (N_36758,N_33610,N_34227);
nand U36759 (N_36759,N_33032,N_33799);
and U36760 (N_36760,N_33504,N_32636);
nand U36761 (N_36761,N_33371,N_34645);
nand U36762 (N_36762,N_32942,N_34775);
nand U36763 (N_36763,N_32911,N_32632);
and U36764 (N_36764,N_33904,N_34443);
nand U36765 (N_36765,N_32726,N_33978);
or U36766 (N_36766,N_34931,N_34475);
or U36767 (N_36767,N_34755,N_34507);
nand U36768 (N_36768,N_32858,N_34436);
or U36769 (N_36769,N_34341,N_33467);
nor U36770 (N_36770,N_32893,N_33974);
or U36771 (N_36771,N_34154,N_33665);
xnor U36772 (N_36772,N_34976,N_34564);
nor U36773 (N_36773,N_32633,N_33689);
nand U36774 (N_36774,N_33524,N_33277);
nor U36775 (N_36775,N_33506,N_34812);
xor U36776 (N_36776,N_33039,N_33756);
or U36777 (N_36777,N_34310,N_33642);
nand U36778 (N_36778,N_32760,N_33443);
nand U36779 (N_36779,N_33368,N_34867);
or U36780 (N_36780,N_32657,N_33327);
and U36781 (N_36781,N_33898,N_34323);
and U36782 (N_36782,N_33650,N_34829);
xnor U36783 (N_36783,N_32523,N_33753);
or U36784 (N_36784,N_33476,N_34166);
xnor U36785 (N_36785,N_33839,N_34364);
nor U36786 (N_36786,N_34510,N_34673);
and U36787 (N_36787,N_34212,N_33004);
xor U36788 (N_36788,N_34668,N_33541);
and U36789 (N_36789,N_34468,N_34306);
and U36790 (N_36790,N_33359,N_33945);
and U36791 (N_36791,N_33985,N_32518);
nand U36792 (N_36792,N_34020,N_32741);
nor U36793 (N_36793,N_32613,N_33004);
and U36794 (N_36794,N_33736,N_33567);
nand U36795 (N_36795,N_34264,N_33144);
and U36796 (N_36796,N_32843,N_32942);
nand U36797 (N_36797,N_34204,N_33093);
and U36798 (N_36798,N_32925,N_33942);
nor U36799 (N_36799,N_32632,N_34909);
or U36800 (N_36800,N_34381,N_32723);
and U36801 (N_36801,N_32688,N_33759);
xnor U36802 (N_36802,N_32945,N_32850);
nor U36803 (N_36803,N_34449,N_32523);
and U36804 (N_36804,N_33048,N_33396);
nor U36805 (N_36805,N_33734,N_34764);
nor U36806 (N_36806,N_34668,N_32533);
nand U36807 (N_36807,N_34493,N_33513);
and U36808 (N_36808,N_34206,N_33230);
or U36809 (N_36809,N_33144,N_33885);
xor U36810 (N_36810,N_34033,N_32732);
nand U36811 (N_36811,N_33174,N_33268);
or U36812 (N_36812,N_34626,N_34373);
and U36813 (N_36813,N_33430,N_33675);
xnor U36814 (N_36814,N_33339,N_34239);
xor U36815 (N_36815,N_33119,N_33646);
and U36816 (N_36816,N_34166,N_34097);
nand U36817 (N_36817,N_34770,N_32987);
and U36818 (N_36818,N_33523,N_34077);
nand U36819 (N_36819,N_34641,N_34403);
or U36820 (N_36820,N_34166,N_34514);
xnor U36821 (N_36821,N_33345,N_33031);
nor U36822 (N_36822,N_33981,N_32719);
xor U36823 (N_36823,N_34973,N_34261);
and U36824 (N_36824,N_33976,N_32894);
and U36825 (N_36825,N_33003,N_34980);
xor U36826 (N_36826,N_33668,N_33179);
or U36827 (N_36827,N_33417,N_32794);
nand U36828 (N_36828,N_32998,N_33144);
nand U36829 (N_36829,N_32745,N_34971);
nand U36830 (N_36830,N_34365,N_34598);
and U36831 (N_36831,N_33466,N_33270);
xnor U36832 (N_36832,N_34551,N_34437);
and U36833 (N_36833,N_34176,N_34899);
nand U36834 (N_36834,N_33662,N_33939);
nor U36835 (N_36835,N_33485,N_33204);
xnor U36836 (N_36836,N_34570,N_33641);
nand U36837 (N_36837,N_33985,N_34052);
nor U36838 (N_36838,N_32601,N_34777);
xor U36839 (N_36839,N_32561,N_33377);
nor U36840 (N_36840,N_34549,N_32535);
or U36841 (N_36841,N_33537,N_32971);
nand U36842 (N_36842,N_32688,N_34053);
nand U36843 (N_36843,N_33927,N_32698);
nor U36844 (N_36844,N_33821,N_34317);
xor U36845 (N_36845,N_33234,N_34038);
xor U36846 (N_36846,N_33706,N_32739);
nand U36847 (N_36847,N_33640,N_33936);
or U36848 (N_36848,N_32562,N_33350);
and U36849 (N_36849,N_33133,N_34221);
nor U36850 (N_36850,N_33514,N_32953);
nand U36851 (N_36851,N_34999,N_32505);
and U36852 (N_36852,N_33770,N_33378);
or U36853 (N_36853,N_33266,N_34253);
nor U36854 (N_36854,N_33487,N_33062);
and U36855 (N_36855,N_33273,N_33246);
nor U36856 (N_36856,N_33209,N_34293);
or U36857 (N_36857,N_33414,N_34001);
and U36858 (N_36858,N_33416,N_34692);
nand U36859 (N_36859,N_33835,N_34430);
nand U36860 (N_36860,N_34070,N_32905);
and U36861 (N_36861,N_33177,N_33922);
or U36862 (N_36862,N_34460,N_34038);
nor U36863 (N_36863,N_33166,N_34090);
or U36864 (N_36864,N_34975,N_33511);
and U36865 (N_36865,N_33706,N_33114);
nand U36866 (N_36866,N_33097,N_32617);
xor U36867 (N_36867,N_33011,N_34976);
xnor U36868 (N_36868,N_34744,N_34973);
nand U36869 (N_36869,N_32881,N_34358);
and U36870 (N_36870,N_32789,N_34803);
nand U36871 (N_36871,N_33074,N_34911);
nand U36872 (N_36872,N_34455,N_34303);
and U36873 (N_36873,N_33999,N_33897);
and U36874 (N_36874,N_33338,N_32811);
nor U36875 (N_36875,N_33186,N_34164);
and U36876 (N_36876,N_33898,N_34821);
nand U36877 (N_36877,N_34401,N_33565);
nand U36878 (N_36878,N_33484,N_33666);
nor U36879 (N_36879,N_33615,N_33470);
nor U36880 (N_36880,N_34807,N_34704);
nand U36881 (N_36881,N_34033,N_33385);
and U36882 (N_36882,N_32620,N_33639);
xnor U36883 (N_36883,N_34337,N_32580);
xnor U36884 (N_36884,N_32822,N_34023);
or U36885 (N_36885,N_33951,N_34484);
and U36886 (N_36886,N_33655,N_34536);
and U36887 (N_36887,N_33426,N_33559);
xor U36888 (N_36888,N_33348,N_32512);
xor U36889 (N_36889,N_33892,N_33020);
xnor U36890 (N_36890,N_33691,N_32969);
or U36891 (N_36891,N_32801,N_33381);
nor U36892 (N_36892,N_32566,N_32908);
nand U36893 (N_36893,N_33724,N_32770);
xnor U36894 (N_36894,N_33726,N_33997);
nand U36895 (N_36895,N_33762,N_32942);
nor U36896 (N_36896,N_33475,N_34156);
nand U36897 (N_36897,N_33420,N_32730);
xnor U36898 (N_36898,N_33316,N_32611);
nand U36899 (N_36899,N_34531,N_34321);
or U36900 (N_36900,N_34347,N_33689);
nand U36901 (N_36901,N_32933,N_33373);
nand U36902 (N_36902,N_34139,N_33356);
nand U36903 (N_36903,N_34377,N_33421);
nand U36904 (N_36904,N_32869,N_32519);
and U36905 (N_36905,N_34502,N_34457);
nand U36906 (N_36906,N_34079,N_34828);
or U36907 (N_36907,N_33344,N_33264);
and U36908 (N_36908,N_34265,N_34554);
nor U36909 (N_36909,N_34187,N_32570);
xnor U36910 (N_36910,N_34870,N_33611);
and U36911 (N_36911,N_34131,N_33333);
nand U36912 (N_36912,N_33612,N_33158);
xor U36913 (N_36913,N_34222,N_33270);
nor U36914 (N_36914,N_34292,N_34731);
nor U36915 (N_36915,N_32681,N_34158);
and U36916 (N_36916,N_34703,N_34804);
xor U36917 (N_36917,N_34682,N_34174);
nand U36918 (N_36918,N_34865,N_33249);
or U36919 (N_36919,N_34572,N_33094);
and U36920 (N_36920,N_32947,N_33236);
or U36921 (N_36921,N_34843,N_33389);
xnor U36922 (N_36922,N_34016,N_33039);
xnor U36923 (N_36923,N_32854,N_32776);
xor U36924 (N_36924,N_32675,N_32589);
nand U36925 (N_36925,N_32788,N_32941);
xor U36926 (N_36926,N_34033,N_33462);
nand U36927 (N_36927,N_34164,N_34685);
xnor U36928 (N_36928,N_33550,N_34421);
or U36929 (N_36929,N_32524,N_34977);
nor U36930 (N_36930,N_34425,N_33806);
nand U36931 (N_36931,N_33514,N_33797);
and U36932 (N_36932,N_34093,N_32921);
nor U36933 (N_36933,N_34897,N_32613);
xnor U36934 (N_36934,N_33417,N_34770);
xnor U36935 (N_36935,N_33882,N_34117);
nor U36936 (N_36936,N_32601,N_33918);
xnor U36937 (N_36937,N_34006,N_32566);
nor U36938 (N_36938,N_34010,N_34606);
xnor U36939 (N_36939,N_33873,N_34688);
or U36940 (N_36940,N_33607,N_34509);
xnor U36941 (N_36941,N_32716,N_34486);
and U36942 (N_36942,N_32612,N_33043);
or U36943 (N_36943,N_32698,N_33624);
and U36944 (N_36944,N_32972,N_32746);
nand U36945 (N_36945,N_34134,N_34192);
and U36946 (N_36946,N_33109,N_33108);
or U36947 (N_36947,N_32764,N_32599);
nand U36948 (N_36948,N_32893,N_32860);
and U36949 (N_36949,N_33822,N_32570);
nand U36950 (N_36950,N_32577,N_34826);
or U36951 (N_36951,N_34107,N_33137);
xnor U36952 (N_36952,N_34613,N_34309);
nand U36953 (N_36953,N_34034,N_33884);
nand U36954 (N_36954,N_32615,N_32736);
and U36955 (N_36955,N_33600,N_33490);
nor U36956 (N_36956,N_33802,N_33285);
and U36957 (N_36957,N_34286,N_33435);
nand U36958 (N_36958,N_33569,N_34538);
xor U36959 (N_36959,N_34803,N_34782);
nand U36960 (N_36960,N_32672,N_34592);
nand U36961 (N_36961,N_33623,N_34578);
xor U36962 (N_36962,N_34925,N_33390);
or U36963 (N_36963,N_32994,N_33973);
and U36964 (N_36964,N_34978,N_32924);
xor U36965 (N_36965,N_32711,N_33040);
or U36966 (N_36966,N_34744,N_33545);
xor U36967 (N_36967,N_33038,N_33442);
or U36968 (N_36968,N_34293,N_32750);
and U36969 (N_36969,N_34371,N_34322);
and U36970 (N_36970,N_33429,N_34244);
xnor U36971 (N_36971,N_32830,N_34737);
nand U36972 (N_36972,N_33422,N_33863);
xnor U36973 (N_36973,N_33078,N_34491);
xnor U36974 (N_36974,N_34394,N_33540);
nand U36975 (N_36975,N_33290,N_33453);
xnor U36976 (N_36976,N_32998,N_33430);
nor U36977 (N_36977,N_32690,N_33514);
xnor U36978 (N_36978,N_34717,N_32569);
nand U36979 (N_36979,N_34582,N_34365);
and U36980 (N_36980,N_32922,N_33637);
and U36981 (N_36981,N_33474,N_34904);
or U36982 (N_36982,N_33819,N_34861);
and U36983 (N_36983,N_33395,N_33700);
or U36984 (N_36984,N_34154,N_33264);
and U36985 (N_36985,N_34373,N_33542);
nor U36986 (N_36986,N_33734,N_34821);
or U36987 (N_36987,N_33407,N_34370);
and U36988 (N_36988,N_34261,N_34563);
or U36989 (N_36989,N_33277,N_32859);
or U36990 (N_36990,N_33862,N_32590);
xor U36991 (N_36991,N_34914,N_33373);
and U36992 (N_36992,N_33612,N_33397);
nand U36993 (N_36993,N_32778,N_33960);
nand U36994 (N_36994,N_32759,N_34040);
xor U36995 (N_36995,N_32624,N_34929);
or U36996 (N_36996,N_33438,N_33758);
nand U36997 (N_36997,N_34022,N_34001);
and U36998 (N_36998,N_33364,N_33136);
nand U36999 (N_36999,N_33871,N_34712);
nand U37000 (N_37000,N_34801,N_34547);
nor U37001 (N_37001,N_32687,N_33193);
nand U37002 (N_37002,N_32686,N_34855);
xnor U37003 (N_37003,N_33076,N_34290);
xnor U37004 (N_37004,N_33492,N_33395);
xnor U37005 (N_37005,N_34459,N_34715);
and U37006 (N_37006,N_33784,N_33715);
or U37007 (N_37007,N_33061,N_34512);
xor U37008 (N_37008,N_34447,N_33676);
or U37009 (N_37009,N_33683,N_33151);
and U37010 (N_37010,N_33628,N_33319);
or U37011 (N_37011,N_34160,N_34505);
xor U37012 (N_37012,N_32610,N_33026);
or U37013 (N_37013,N_33720,N_33183);
nor U37014 (N_37014,N_34122,N_32716);
xor U37015 (N_37015,N_33351,N_32916);
and U37016 (N_37016,N_33143,N_33914);
nor U37017 (N_37017,N_33368,N_34618);
or U37018 (N_37018,N_33212,N_32598);
or U37019 (N_37019,N_34039,N_33118);
nand U37020 (N_37020,N_32831,N_32816);
xor U37021 (N_37021,N_33141,N_33704);
xor U37022 (N_37022,N_34192,N_34952);
and U37023 (N_37023,N_33914,N_33672);
nand U37024 (N_37024,N_34635,N_32561);
nand U37025 (N_37025,N_33610,N_34484);
and U37026 (N_37026,N_34180,N_32945);
nor U37027 (N_37027,N_32937,N_34107);
and U37028 (N_37028,N_34434,N_33995);
nor U37029 (N_37029,N_32699,N_33157);
xor U37030 (N_37030,N_34291,N_32958);
nand U37031 (N_37031,N_34829,N_34804);
xor U37032 (N_37032,N_33149,N_33327);
xnor U37033 (N_37033,N_33314,N_32812);
nand U37034 (N_37034,N_34605,N_34382);
or U37035 (N_37035,N_34030,N_33826);
nand U37036 (N_37036,N_32819,N_34305);
nor U37037 (N_37037,N_33554,N_33435);
or U37038 (N_37038,N_34811,N_32643);
and U37039 (N_37039,N_34015,N_33745);
xnor U37040 (N_37040,N_34372,N_34048);
nand U37041 (N_37041,N_34701,N_32990);
or U37042 (N_37042,N_34239,N_34714);
or U37043 (N_37043,N_32913,N_34532);
xor U37044 (N_37044,N_34422,N_34035);
nor U37045 (N_37045,N_34888,N_32967);
and U37046 (N_37046,N_34179,N_34064);
or U37047 (N_37047,N_32842,N_33802);
xor U37048 (N_37048,N_33000,N_33088);
nand U37049 (N_37049,N_33592,N_34721);
xor U37050 (N_37050,N_34550,N_33314);
and U37051 (N_37051,N_32508,N_34671);
nor U37052 (N_37052,N_34999,N_33709);
nand U37053 (N_37053,N_33392,N_33521);
or U37054 (N_37054,N_33339,N_33399);
and U37055 (N_37055,N_33987,N_33635);
nor U37056 (N_37056,N_34902,N_34662);
nor U37057 (N_37057,N_34386,N_34296);
or U37058 (N_37058,N_33821,N_33006);
nand U37059 (N_37059,N_33781,N_32738);
or U37060 (N_37060,N_33829,N_32599);
or U37061 (N_37061,N_33894,N_32824);
xor U37062 (N_37062,N_34572,N_34345);
nand U37063 (N_37063,N_34551,N_33833);
or U37064 (N_37064,N_33639,N_32649);
nand U37065 (N_37065,N_34916,N_34712);
and U37066 (N_37066,N_34345,N_34364);
or U37067 (N_37067,N_33839,N_34140);
nand U37068 (N_37068,N_33539,N_34312);
or U37069 (N_37069,N_33319,N_34894);
nor U37070 (N_37070,N_32620,N_32946);
nand U37071 (N_37071,N_33327,N_33525);
and U37072 (N_37072,N_33907,N_34401);
xor U37073 (N_37073,N_34013,N_33532);
nor U37074 (N_37074,N_32545,N_34416);
nor U37075 (N_37075,N_33373,N_34644);
nand U37076 (N_37076,N_32905,N_32773);
xor U37077 (N_37077,N_34548,N_32529);
xor U37078 (N_37078,N_33651,N_34369);
xor U37079 (N_37079,N_34655,N_34992);
and U37080 (N_37080,N_33851,N_33703);
xor U37081 (N_37081,N_34767,N_33657);
nand U37082 (N_37082,N_34091,N_34214);
xor U37083 (N_37083,N_32781,N_32508);
and U37084 (N_37084,N_34305,N_34012);
nor U37085 (N_37085,N_34408,N_32671);
xnor U37086 (N_37086,N_34392,N_33208);
or U37087 (N_37087,N_33630,N_34667);
nor U37088 (N_37088,N_34836,N_33034);
or U37089 (N_37089,N_34246,N_33007);
or U37090 (N_37090,N_34702,N_34154);
nor U37091 (N_37091,N_33839,N_33515);
or U37092 (N_37092,N_32865,N_33703);
or U37093 (N_37093,N_33427,N_32955);
xnor U37094 (N_37094,N_34130,N_34990);
nand U37095 (N_37095,N_32995,N_34432);
or U37096 (N_37096,N_34490,N_33632);
and U37097 (N_37097,N_33829,N_32511);
nand U37098 (N_37098,N_34423,N_34085);
nor U37099 (N_37099,N_32818,N_32799);
or U37100 (N_37100,N_33238,N_34453);
nor U37101 (N_37101,N_33547,N_34116);
or U37102 (N_37102,N_34709,N_32824);
and U37103 (N_37103,N_34361,N_34360);
xor U37104 (N_37104,N_34737,N_34677);
or U37105 (N_37105,N_33641,N_34720);
xnor U37106 (N_37106,N_33170,N_32810);
xor U37107 (N_37107,N_33793,N_32910);
xnor U37108 (N_37108,N_33021,N_33964);
nor U37109 (N_37109,N_33317,N_34071);
and U37110 (N_37110,N_32817,N_34702);
nand U37111 (N_37111,N_33091,N_32659);
xnor U37112 (N_37112,N_34445,N_34747);
xnor U37113 (N_37113,N_33226,N_33148);
xor U37114 (N_37114,N_33084,N_34086);
nand U37115 (N_37115,N_33855,N_32631);
nor U37116 (N_37116,N_33000,N_33023);
nand U37117 (N_37117,N_33643,N_33513);
xnor U37118 (N_37118,N_33443,N_34510);
nand U37119 (N_37119,N_33911,N_33224);
or U37120 (N_37120,N_34682,N_34430);
xor U37121 (N_37121,N_33429,N_33148);
and U37122 (N_37122,N_34718,N_34666);
nand U37123 (N_37123,N_33289,N_34316);
nand U37124 (N_37124,N_33106,N_33934);
or U37125 (N_37125,N_32895,N_34867);
xnor U37126 (N_37126,N_34722,N_34617);
xnor U37127 (N_37127,N_34435,N_32906);
nor U37128 (N_37128,N_33457,N_34576);
nor U37129 (N_37129,N_33391,N_33810);
and U37130 (N_37130,N_34612,N_32740);
or U37131 (N_37131,N_33953,N_34392);
nand U37132 (N_37132,N_32805,N_32900);
nor U37133 (N_37133,N_34962,N_33097);
or U37134 (N_37134,N_33646,N_33662);
xor U37135 (N_37135,N_32827,N_34514);
nand U37136 (N_37136,N_34907,N_32663);
nor U37137 (N_37137,N_34513,N_33068);
xor U37138 (N_37138,N_34068,N_33945);
or U37139 (N_37139,N_34034,N_34578);
nor U37140 (N_37140,N_33873,N_34229);
or U37141 (N_37141,N_34024,N_33298);
xor U37142 (N_37142,N_34422,N_32863);
nand U37143 (N_37143,N_33155,N_32578);
nand U37144 (N_37144,N_34819,N_33152);
or U37145 (N_37145,N_34334,N_34473);
xor U37146 (N_37146,N_33140,N_33751);
and U37147 (N_37147,N_33822,N_33933);
nor U37148 (N_37148,N_34449,N_32588);
xor U37149 (N_37149,N_34020,N_34514);
nor U37150 (N_37150,N_32706,N_34087);
and U37151 (N_37151,N_33096,N_33502);
and U37152 (N_37152,N_34596,N_34826);
nand U37153 (N_37153,N_34079,N_33875);
xor U37154 (N_37154,N_34391,N_32643);
nand U37155 (N_37155,N_34321,N_33745);
xor U37156 (N_37156,N_32538,N_33431);
nor U37157 (N_37157,N_32934,N_32886);
nor U37158 (N_37158,N_32511,N_33544);
or U37159 (N_37159,N_33437,N_33284);
nand U37160 (N_37160,N_33943,N_34604);
and U37161 (N_37161,N_34190,N_34171);
or U37162 (N_37162,N_32744,N_33928);
nor U37163 (N_37163,N_33665,N_33186);
xnor U37164 (N_37164,N_32510,N_34017);
or U37165 (N_37165,N_33976,N_33535);
or U37166 (N_37166,N_33504,N_33563);
nand U37167 (N_37167,N_34434,N_33797);
and U37168 (N_37168,N_33109,N_33313);
nor U37169 (N_37169,N_32790,N_34804);
xor U37170 (N_37170,N_33105,N_33607);
nor U37171 (N_37171,N_33431,N_34821);
and U37172 (N_37172,N_34594,N_33428);
nor U37173 (N_37173,N_32658,N_34178);
nand U37174 (N_37174,N_33471,N_34969);
nand U37175 (N_37175,N_32692,N_34330);
nor U37176 (N_37176,N_34725,N_34865);
and U37177 (N_37177,N_33510,N_32867);
xor U37178 (N_37178,N_34949,N_34511);
and U37179 (N_37179,N_34723,N_32664);
or U37180 (N_37180,N_33639,N_34699);
nand U37181 (N_37181,N_34357,N_33191);
xor U37182 (N_37182,N_34138,N_33499);
and U37183 (N_37183,N_33095,N_34695);
and U37184 (N_37184,N_32917,N_32724);
and U37185 (N_37185,N_33902,N_33203);
nand U37186 (N_37186,N_32589,N_33729);
and U37187 (N_37187,N_32694,N_34838);
nor U37188 (N_37188,N_34948,N_33452);
nand U37189 (N_37189,N_34607,N_34208);
nor U37190 (N_37190,N_33795,N_33427);
or U37191 (N_37191,N_32689,N_33001);
nand U37192 (N_37192,N_33477,N_33361);
xnor U37193 (N_37193,N_33874,N_34070);
xnor U37194 (N_37194,N_33615,N_34823);
nand U37195 (N_37195,N_33401,N_33427);
nand U37196 (N_37196,N_33569,N_34528);
or U37197 (N_37197,N_32603,N_33079);
xnor U37198 (N_37198,N_33863,N_34402);
nor U37199 (N_37199,N_33272,N_33832);
nand U37200 (N_37200,N_32874,N_32536);
nor U37201 (N_37201,N_33811,N_33747);
and U37202 (N_37202,N_33652,N_34612);
or U37203 (N_37203,N_33102,N_32519);
or U37204 (N_37204,N_33178,N_32853);
xnor U37205 (N_37205,N_32508,N_32813);
or U37206 (N_37206,N_34596,N_33282);
and U37207 (N_37207,N_33801,N_32813);
or U37208 (N_37208,N_33706,N_32581);
xor U37209 (N_37209,N_33019,N_32588);
or U37210 (N_37210,N_32978,N_33057);
and U37211 (N_37211,N_34638,N_32978);
xor U37212 (N_37212,N_34272,N_34610);
xor U37213 (N_37213,N_32996,N_33932);
and U37214 (N_37214,N_34824,N_34700);
or U37215 (N_37215,N_32830,N_32858);
or U37216 (N_37216,N_32827,N_34040);
and U37217 (N_37217,N_34344,N_34458);
or U37218 (N_37218,N_33658,N_33317);
and U37219 (N_37219,N_34847,N_34808);
xnor U37220 (N_37220,N_33302,N_34552);
nand U37221 (N_37221,N_34152,N_33725);
or U37222 (N_37222,N_32936,N_33364);
xor U37223 (N_37223,N_34434,N_32838);
nand U37224 (N_37224,N_33625,N_32597);
nand U37225 (N_37225,N_32791,N_33893);
or U37226 (N_37226,N_32897,N_33016);
or U37227 (N_37227,N_33676,N_33917);
or U37228 (N_37228,N_34599,N_34571);
xnor U37229 (N_37229,N_32802,N_32844);
nand U37230 (N_37230,N_34918,N_33071);
xor U37231 (N_37231,N_34143,N_32682);
nor U37232 (N_37232,N_34789,N_34026);
xnor U37233 (N_37233,N_32588,N_32749);
xnor U37234 (N_37234,N_34638,N_33786);
nand U37235 (N_37235,N_32671,N_33645);
and U37236 (N_37236,N_34796,N_34206);
nand U37237 (N_37237,N_33790,N_34835);
or U37238 (N_37238,N_34296,N_32990);
and U37239 (N_37239,N_32753,N_34235);
and U37240 (N_37240,N_34964,N_33827);
and U37241 (N_37241,N_34555,N_32610);
and U37242 (N_37242,N_34766,N_33718);
or U37243 (N_37243,N_33970,N_33821);
nor U37244 (N_37244,N_33747,N_33690);
and U37245 (N_37245,N_32840,N_33168);
xor U37246 (N_37246,N_34624,N_33584);
and U37247 (N_37247,N_33037,N_33613);
or U37248 (N_37248,N_33064,N_34226);
xor U37249 (N_37249,N_34117,N_34239);
or U37250 (N_37250,N_33779,N_34588);
or U37251 (N_37251,N_32999,N_32846);
or U37252 (N_37252,N_32638,N_33583);
and U37253 (N_37253,N_33326,N_34185);
and U37254 (N_37254,N_34638,N_33160);
or U37255 (N_37255,N_32868,N_34372);
or U37256 (N_37256,N_34688,N_34504);
xnor U37257 (N_37257,N_32708,N_32614);
or U37258 (N_37258,N_32797,N_34907);
xor U37259 (N_37259,N_32640,N_32597);
and U37260 (N_37260,N_34649,N_32677);
nand U37261 (N_37261,N_32608,N_33147);
xor U37262 (N_37262,N_33947,N_32668);
nor U37263 (N_37263,N_33899,N_34891);
and U37264 (N_37264,N_32911,N_34682);
nor U37265 (N_37265,N_33328,N_34234);
nor U37266 (N_37266,N_34242,N_32773);
and U37267 (N_37267,N_33896,N_34268);
xor U37268 (N_37268,N_33198,N_34939);
nand U37269 (N_37269,N_32709,N_33776);
or U37270 (N_37270,N_33037,N_34131);
nor U37271 (N_37271,N_34885,N_32681);
and U37272 (N_37272,N_34297,N_34900);
nor U37273 (N_37273,N_34390,N_32705);
nand U37274 (N_37274,N_34991,N_33100);
and U37275 (N_37275,N_34269,N_32892);
nor U37276 (N_37276,N_33464,N_32831);
nand U37277 (N_37277,N_34770,N_34476);
nor U37278 (N_37278,N_34861,N_34883);
nand U37279 (N_37279,N_32847,N_32943);
and U37280 (N_37280,N_33049,N_34786);
or U37281 (N_37281,N_32982,N_34460);
xnor U37282 (N_37282,N_32710,N_34865);
and U37283 (N_37283,N_33961,N_32580);
nand U37284 (N_37284,N_33674,N_32585);
nor U37285 (N_37285,N_34727,N_34370);
or U37286 (N_37286,N_34354,N_34296);
nor U37287 (N_37287,N_33376,N_32688);
xnor U37288 (N_37288,N_34320,N_32714);
nor U37289 (N_37289,N_33150,N_34885);
and U37290 (N_37290,N_34928,N_33194);
nor U37291 (N_37291,N_34071,N_33993);
nand U37292 (N_37292,N_33004,N_34530);
nand U37293 (N_37293,N_33972,N_33467);
xor U37294 (N_37294,N_33920,N_34506);
or U37295 (N_37295,N_34161,N_32633);
or U37296 (N_37296,N_34600,N_33176);
and U37297 (N_37297,N_34657,N_33876);
or U37298 (N_37298,N_33597,N_32587);
xor U37299 (N_37299,N_34283,N_33520);
or U37300 (N_37300,N_33188,N_34458);
nor U37301 (N_37301,N_32969,N_33554);
or U37302 (N_37302,N_32865,N_34444);
and U37303 (N_37303,N_34837,N_33228);
nor U37304 (N_37304,N_33005,N_32555);
or U37305 (N_37305,N_32802,N_34962);
nand U37306 (N_37306,N_33769,N_34500);
nand U37307 (N_37307,N_34663,N_33813);
or U37308 (N_37308,N_34175,N_32939);
and U37309 (N_37309,N_34871,N_34647);
and U37310 (N_37310,N_32999,N_32883);
nor U37311 (N_37311,N_33439,N_34622);
nor U37312 (N_37312,N_34502,N_34405);
nand U37313 (N_37313,N_32514,N_34325);
nand U37314 (N_37314,N_33974,N_34400);
xor U37315 (N_37315,N_33522,N_34058);
nand U37316 (N_37316,N_34872,N_34899);
nor U37317 (N_37317,N_32816,N_34739);
or U37318 (N_37318,N_33211,N_32532);
xor U37319 (N_37319,N_32618,N_34421);
or U37320 (N_37320,N_33714,N_34623);
and U37321 (N_37321,N_34605,N_34793);
nand U37322 (N_37322,N_34056,N_34755);
xor U37323 (N_37323,N_32573,N_33565);
nor U37324 (N_37324,N_33042,N_33216);
nor U37325 (N_37325,N_34580,N_34735);
and U37326 (N_37326,N_33791,N_33990);
nor U37327 (N_37327,N_34829,N_33415);
and U37328 (N_37328,N_32573,N_34810);
nor U37329 (N_37329,N_34519,N_33514);
nor U37330 (N_37330,N_34865,N_34903);
xnor U37331 (N_37331,N_34065,N_33232);
or U37332 (N_37332,N_32565,N_34267);
nand U37333 (N_37333,N_33095,N_34615);
nand U37334 (N_37334,N_34795,N_33022);
xnor U37335 (N_37335,N_32944,N_33210);
nor U37336 (N_37336,N_34553,N_33643);
xnor U37337 (N_37337,N_33986,N_33904);
nor U37338 (N_37338,N_34095,N_34345);
nand U37339 (N_37339,N_33952,N_34414);
nand U37340 (N_37340,N_34301,N_33373);
nand U37341 (N_37341,N_33600,N_32630);
xnor U37342 (N_37342,N_32741,N_34453);
nand U37343 (N_37343,N_33188,N_32744);
xnor U37344 (N_37344,N_32541,N_34081);
or U37345 (N_37345,N_33038,N_33978);
nand U37346 (N_37346,N_34085,N_34813);
or U37347 (N_37347,N_33487,N_33324);
nor U37348 (N_37348,N_32937,N_32523);
or U37349 (N_37349,N_34201,N_33255);
nand U37350 (N_37350,N_33589,N_33528);
nor U37351 (N_37351,N_32623,N_33119);
xor U37352 (N_37352,N_34190,N_33171);
xnor U37353 (N_37353,N_32997,N_32521);
xor U37354 (N_37354,N_33757,N_33112);
and U37355 (N_37355,N_33283,N_34229);
and U37356 (N_37356,N_32581,N_33329);
and U37357 (N_37357,N_33521,N_34053);
or U37358 (N_37358,N_34204,N_32616);
or U37359 (N_37359,N_34559,N_34253);
xnor U37360 (N_37360,N_34039,N_33874);
and U37361 (N_37361,N_34505,N_34150);
or U37362 (N_37362,N_32543,N_34341);
xor U37363 (N_37363,N_33097,N_34933);
nand U37364 (N_37364,N_32850,N_32520);
or U37365 (N_37365,N_32535,N_32992);
xor U37366 (N_37366,N_34392,N_34534);
xnor U37367 (N_37367,N_32620,N_33633);
nand U37368 (N_37368,N_33615,N_33246);
or U37369 (N_37369,N_33774,N_32751);
nor U37370 (N_37370,N_33096,N_33690);
xor U37371 (N_37371,N_33733,N_32809);
and U37372 (N_37372,N_34255,N_34636);
nor U37373 (N_37373,N_34862,N_33314);
xnor U37374 (N_37374,N_32714,N_33409);
nand U37375 (N_37375,N_34297,N_32662);
nand U37376 (N_37376,N_33649,N_33505);
or U37377 (N_37377,N_33073,N_34669);
or U37378 (N_37378,N_34106,N_33151);
and U37379 (N_37379,N_33353,N_33292);
nor U37380 (N_37380,N_32789,N_33817);
and U37381 (N_37381,N_32650,N_34028);
nor U37382 (N_37382,N_32847,N_33241);
and U37383 (N_37383,N_33631,N_32981);
nor U37384 (N_37384,N_34708,N_33966);
or U37385 (N_37385,N_34890,N_32712);
and U37386 (N_37386,N_34739,N_34907);
nor U37387 (N_37387,N_34754,N_33258);
nor U37388 (N_37388,N_32575,N_32828);
xnor U37389 (N_37389,N_33406,N_32808);
xnor U37390 (N_37390,N_32565,N_34428);
nand U37391 (N_37391,N_34837,N_33768);
nor U37392 (N_37392,N_34359,N_32831);
nand U37393 (N_37393,N_33036,N_34422);
nor U37394 (N_37394,N_33417,N_32918);
and U37395 (N_37395,N_33963,N_33399);
and U37396 (N_37396,N_33090,N_34640);
xnor U37397 (N_37397,N_32878,N_34595);
and U37398 (N_37398,N_34156,N_33413);
nand U37399 (N_37399,N_33783,N_34317);
or U37400 (N_37400,N_33312,N_32817);
nor U37401 (N_37401,N_32547,N_34252);
nor U37402 (N_37402,N_34313,N_34624);
and U37403 (N_37403,N_34223,N_33242);
xor U37404 (N_37404,N_32879,N_34402);
or U37405 (N_37405,N_33733,N_32915);
or U37406 (N_37406,N_32851,N_33558);
and U37407 (N_37407,N_33803,N_33150);
nor U37408 (N_37408,N_34797,N_33342);
or U37409 (N_37409,N_32756,N_33625);
xnor U37410 (N_37410,N_34376,N_34781);
nor U37411 (N_37411,N_32980,N_33043);
xnor U37412 (N_37412,N_34502,N_34963);
and U37413 (N_37413,N_32631,N_33507);
or U37414 (N_37414,N_33651,N_32564);
xor U37415 (N_37415,N_34932,N_33634);
nor U37416 (N_37416,N_34162,N_34519);
nand U37417 (N_37417,N_34337,N_32890);
or U37418 (N_37418,N_33420,N_34504);
xor U37419 (N_37419,N_34461,N_34033);
nand U37420 (N_37420,N_33674,N_34785);
xnor U37421 (N_37421,N_33254,N_34969);
xnor U37422 (N_37422,N_34460,N_34402);
and U37423 (N_37423,N_33507,N_33007);
nand U37424 (N_37424,N_34533,N_32550);
and U37425 (N_37425,N_32530,N_33963);
or U37426 (N_37426,N_34660,N_34273);
or U37427 (N_37427,N_33951,N_34840);
nor U37428 (N_37428,N_34645,N_33868);
or U37429 (N_37429,N_32508,N_33333);
xnor U37430 (N_37430,N_33988,N_34616);
and U37431 (N_37431,N_33933,N_33366);
nor U37432 (N_37432,N_34202,N_32723);
nor U37433 (N_37433,N_34802,N_32767);
or U37434 (N_37434,N_34956,N_33322);
nand U37435 (N_37435,N_34850,N_32664);
and U37436 (N_37436,N_34539,N_33572);
or U37437 (N_37437,N_33907,N_34216);
and U37438 (N_37438,N_33050,N_33609);
and U37439 (N_37439,N_33598,N_32624);
nor U37440 (N_37440,N_34493,N_33128);
and U37441 (N_37441,N_33860,N_34555);
and U37442 (N_37442,N_34166,N_33394);
or U37443 (N_37443,N_34124,N_33381);
or U37444 (N_37444,N_32759,N_32772);
nand U37445 (N_37445,N_34541,N_34434);
or U37446 (N_37446,N_33076,N_34905);
and U37447 (N_37447,N_33745,N_33288);
or U37448 (N_37448,N_34809,N_32739);
nor U37449 (N_37449,N_34558,N_33599);
or U37450 (N_37450,N_34504,N_34496);
nand U37451 (N_37451,N_32765,N_34534);
nor U37452 (N_37452,N_33145,N_34573);
and U37453 (N_37453,N_34846,N_34032);
nand U37454 (N_37454,N_34823,N_34897);
nand U37455 (N_37455,N_33235,N_34725);
and U37456 (N_37456,N_34850,N_32501);
nor U37457 (N_37457,N_34693,N_34026);
nand U37458 (N_37458,N_33797,N_33268);
xnor U37459 (N_37459,N_32540,N_34840);
or U37460 (N_37460,N_32663,N_32598);
xor U37461 (N_37461,N_34127,N_33038);
and U37462 (N_37462,N_32671,N_32901);
nor U37463 (N_37463,N_34231,N_33410);
nor U37464 (N_37464,N_34147,N_34812);
nand U37465 (N_37465,N_33029,N_33776);
nor U37466 (N_37466,N_34579,N_33934);
and U37467 (N_37467,N_34532,N_34157);
and U37468 (N_37468,N_33605,N_33497);
or U37469 (N_37469,N_33385,N_32619);
xor U37470 (N_37470,N_32723,N_33729);
nor U37471 (N_37471,N_34233,N_33515);
xor U37472 (N_37472,N_33500,N_34239);
nor U37473 (N_37473,N_34826,N_33678);
nor U37474 (N_37474,N_34809,N_33057);
and U37475 (N_37475,N_34771,N_33282);
and U37476 (N_37476,N_32624,N_32576);
xor U37477 (N_37477,N_32743,N_32996);
nand U37478 (N_37478,N_34766,N_33805);
nor U37479 (N_37479,N_33634,N_34470);
xnor U37480 (N_37480,N_32682,N_34415);
xnor U37481 (N_37481,N_34775,N_34294);
or U37482 (N_37482,N_33638,N_34202);
nor U37483 (N_37483,N_32595,N_32589);
or U37484 (N_37484,N_33498,N_32908);
nor U37485 (N_37485,N_33710,N_32651);
or U37486 (N_37486,N_33823,N_33932);
nor U37487 (N_37487,N_34530,N_34215);
and U37488 (N_37488,N_32723,N_34157);
xor U37489 (N_37489,N_34694,N_34288);
or U37490 (N_37490,N_34320,N_34883);
nor U37491 (N_37491,N_32812,N_32509);
and U37492 (N_37492,N_32837,N_34673);
or U37493 (N_37493,N_32746,N_33394);
and U37494 (N_37494,N_33741,N_33940);
or U37495 (N_37495,N_33964,N_32629);
xnor U37496 (N_37496,N_32844,N_33460);
nand U37497 (N_37497,N_33784,N_34436);
nor U37498 (N_37498,N_33331,N_33804);
nor U37499 (N_37499,N_34454,N_34728);
xnor U37500 (N_37500,N_36524,N_36424);
or U37501 (N_37501,N_36333,N_37071);
nor U37502 (N_37502,N_37485,N_35024);
or U37503 (N_37503,N_36943,N_37182);
nor U37504 (N_37504,N_37322,N_36355);
and U37505 (N_37505,N_35250,N_35271);
and U37506 (N_37506,N_35722,N_35035);
xnor U37507 (N_37507,N_37378,N_36398);
nor U37508 (N_37508,N_36701,N_36986);
and U37509 (N_37509,N_36338,N_35437);
or U37510 (N_37510,N_37460,N_37133);
or U37511 (N_37511,N_37302,N_36092);
or U37512 (N_37512,N_35167,N_37035);
nand U37513 (N_37513,N_35404,N_37254);
nand U37514 (N_37514,N_35081,N_35071);
nor U37515 (N_37515,N_36453,N_35925);
xor U37516 (N_37516,N_35462,N_36569);
nor U37517 (N_37517,N_36924,N_35236);
and U37518 (N_37518,N_35832,N_37179);
nand U37519 (N_37519,N_36987,N_36893);
nor U37520 (N_37520,N_36726,N_37354);
and U37521 (N_37521,N_36533,N_36527);
xnor U37522 (N_37522,N_36509,N_35149);
xor U37523 (N_37523,N_35066,N_35018);
or U37524 (N_37524,N_35456,N_35284);
or U37525 (N_37525,N_35879,N_35045);
or U37526 (N_37526,N_36684,N_35325);
nand U37527 (N_37527,N_35418,N_36538);
or U37528 (N_37528,N_36362,N_37134);
and U37529 (N_37529,N_37203,N_35472);
or U37530 (N_37530,N_35356,N_37454);
and U37531 (N_37531,N_37358,N_37443);
xnor U37532 (N_37532,N_36948,N_37205);
and U37533 (N_37533,N_37076,N_35906);
nand U37534 (N_37534,N_37039,N_36175);
xor U37535 (N_37535,N_36310,N_37029);
and U37536 (N_37536,N_36865,N_35312);
nand U37537 (N_37537,N_36216,N_36014);
and U37538 (N_37538,N_35085,N_37256);
nand U37539 (N_37539,N_36096,N_35015);
and U37540 (N_37540,N_36226,N_35428);
nand U37541 (N_37541,N_35429,N_37157);
nor U37542 (N_37542,N_36196,N_35545);
or U37543 (N_37543,N_37193,N_36162);
nand U37544 (N_37544,N_36003,N_36033);
and U37545 (N_37545,N_36159,N_35176);
and U37546 (N_37546,N_37216,N_36472);
and U37547 (N_37547,N_35354,N_36897);
nor U37548 (N_37548,N_35308,N_36781);
nor U37549 (N_37549,N_36093,N_35178);
or U37550 (N_37550,N_36268,N_35978);
or U37551 (N_37551,N_37158,N_35638);
nor U37552 (N_37552,N_36493,N_37468);
nand U37553 (N_37553,N_37279,N_35280);
nor U37554 (N_37554,N_36690,N_37237);
or U37555 (N_37555,N_35665,N_35927);
xnor U37556 (N_37556,N_37094,N_36755);
xnor U37557 (N_37557,N_36507,N_35020);
nor U37558 (N_37558,N_35949,N_36151);
xnor U37559 (N_37559,N_37127,N_36473);
or U37560 (N_37560,N_36469,N_37299);
and U37561 (N_37561,N_36676,N_36140);
nand U37562 (N_37562,N_37457,N_36366);
nand U37563 (N_37563,N_36702,N_35387);
nor U37564 (N_37564,N_36132,N_37480);
and U37565 (N_37565,N_36077,N_36441);
or U37566 (N_37566,N_36013,N_35068);
xnor U37567 (N_37567,N_35723,N_35923);
or U37568 (N_37568,N_37424,N_36642);
and U37569 (N_37569,N_36724,N_35503);
xnor U37570 (N_37570,N_37130,N_35302);
nor U37571 (N_37571,N_37431,N_35724);
and U37572 (N_37572,N_37275,N_35481);
and U37573 (N_37573,N_35643,N_36011);
nor U37574 (N_37574,N_35448,N_36756);
xnor U37575 (N_37575,N_35818,N_37447);
or U37576 (N_37576,N_37318,N_36904);
xnor U37577 (N_37577,N_35351,N_35861);
xor U37578 (N_37578,N_36858,N_35410);
nor U37579 (N_37579,N_37079,N_35238);
nor U37580 (N_37580,N_37408,N_35393);
nand U37581 (N_37581,N_37102,N_36364);
and U37582 (N_37582,N_36063,N_35430);
or U37583 (N_37583,N_36225,N_35529);
or U37584 (N_37584,N_37272,N_36766);
and U37585 (N_37585,N_37415,N_35594);
or U37586 (N_37586,N_35575,N_35726);
or U37587 (N_37587,N_35884,N_36435);
or U37588 (N_37588,N_35050,N_36452);
nand U37589 (N_37589,N_37494,N_35847);
and U37590 (N_37590,N_35101,N_36431);
or U37591 (N_37591,N_35341,N_36311);
nor U37592 (N_37592,N_35496,N_37381);
xnor U37593 (N_37593,N_36059,N_35819);
xor U37594 (N_37594,N_35548,N_36902);
xor U37595 (N_37595,N_37033,N_36546);
nand U37596 (N_37596,N_36542,N_35403);
or U37597 (N_37597,N_35713,N_36387);
or U37598 (N_37598,N_35672,N_36451);
xor U37599 (N_37599,N_37263,N_35439);
or U37600 (N_37600,N_36985,N_35577);
or U37601 (N_37601,N_35014,N_35477);
nand U37602 (N_37602,N_35019,N_35752);
nor U37603 (N_37603,N_35597,N_36518);
xnor U37604 (N_37604,N_35603,N_36977);
nor U37605 (N_37605,N_35182,N_35118);
or U37606 (N_37606,N_36401,N_35533);
or U37607 (N_37607,N_36845,N_35322);
xor U37608 (N_37608,N_35260,N_36868);
and U37609 (N_37609,N_36298,N_35595);
nand U37610 (N_37610,N_35979,N_37394);
or U37611 (N_37611,N_36358,N_36982);
or U37612 (N_37612,N_36091,N_37296);
nand U37613 (N_37613,N_36625,N_35930);
or U37614 (N_37614,N_36609,N_36791);
nor U37615 (N_37615,N_35968,N_35854);
xnor U37616 (N_37616,N_36848,N_36534);
nor U37617 (N_37617,N_36859,N_37086);
xnor U37618 (N_37618,N_36880,N_36984);
and U37619 (N_37619,N_36267,N_35109);
nor U37620 (N_37620,N_35309,N_35757);
or U37621 (N_37621,N_35041,N_37348);
and U37622 (N_37622,N_35576,N_36434);
xnor U37623 (N_37623,N_37377,N_36694);
xnor U37624 (N_37624,N_36686,N_35796);
or U37625 (N_37625,N_36969,N_35685);
xnor U37626 (N_37626,N_35328,N_36342);
or U37627 (N_37627,N_36009,N_36309);
nand U37628 (N_37628,N_35069,N_37373);
or U37629 (N_37629,N_35324,N_37233);
nand U37630 (N_37630,N_36630,N_36255);
xor U37631 (N_37631,N_37174,N_35047);
and U37632 (N_37632,N_36496,N_36754);
nor U37633 (N_37633,N_36936,N_35358);
nand U37634 (N_37634,N_35692,N_37015);
nor U37635 (N_37635,N_36956,N_36057);
and U37636 (N_37636,N_35952,N_35781);
and U37637 (N_37637,N_36371,N_36891);
nand U37638 (N_37638,N_37006,N_35307);
or U37639 (N_37639,N_36032,N_35834);
and U37640 (N_37640,N_37479,N_35891);
xor U37641 (N_37641,N_35855,N_35886);
or U37642 (N_37642,N_37199,N_35487);
xor U37643 (N_37643,N_36055,N_35426);
and U37644 (N_37644,N_36976,N_36753);
nor U37645 (N_37645,N_36047,N_37321);
and U37646 (N_37646,N_37442,N_37068);
nand U37647 (N_37647,N_37271,N_37308);
xnor U37648 (N_37648,N_35252,N_35580);
or U37649 (N_37649,N_37289,N_36747);
nand U37650 (N_37650,N_36909,N_36651);
nand U37651 (N_37651,N_36039,N_37387);
and U37652 (N_37652,N_35684,N_35158);
xor U37653 (N_37653,N_36210,N_35231);
nand U37654 (N_37654,N_37359,N_37230);
and U37655 (N_37655,N_36591,N_36847);
nand U37656 (N_37656,N_35230,N_35763);
and U37657 (N_37657,N_35080,N_36248);
and U37658 (N_37658,N_37218,N_35212);
nor U37659 (N_37659,N_36922,N_36385);
and U37660 (N_37660,N_36321,N_37267);
and U37661 (N_37661,N_35626,N_36413);
or U37662 (N_37662,N_36919,N_35229);
or U37663 (N_37663,N_35601,N_37420);
and U37664 (N_37664,N_35579,N_35352);
xnor U37665 (N_37665,N_35720,N_36565);
nor U37666 (N_37666,N_37007,N_35918);
nand U37667 (N_37667,N_37148,N_35772);
or U37668 (N_37668,N_35877,N_36719);
xor U37669 (N_37669,N_35895,N_35004);
or U37670 (N_37670,N_37389,N_36634);
and U37671 (N_37671,N_36138,N_37103);
xor U37672 (N_37672,N_36751,N_36894);
and U37673 (N_37673,N_36103,N_35534);
and U37674 (N_37674,N_35520,N_35999);
nor U37675 (N_37675,N_37100,N_35645);
nand U37676 (N_37676,N_35950,N_36721);
or U37677 (N_37677,N_36388,N_35259);
nand U37678 (N_37678,N_36863,N_36040);
or U37679 (N_37679,N_36838,N_35394);
xnor U37680 (N_37680,N_36307,N_36635);
xnor U37681 (N_37681,N_36372,N_37278);
or U37682 (N_37682,N_35868,N_37138);
or U37683 (N_37683,N_37131,N_35216);
nor U37684 (N_37684,N_35138,N_35857);
or U37685 (N_37685,N_35388,N_37057);
nand U37686 (N_37686,N_36019,N_36742);
or U37687 (N_37687,N_35513,N_36641);
nor U37688 (N_37688,N_35465,N_35370);
or U37689 (N_37689,N_36604,N_35803);
nand U37690 (N_37690,N_35632,N_35851);
nand U37691 (N_37691,N_35179,N_36184);
nand U37692 (N_37692,N_36677,N_37108);
and U37693 (N_37693,N_36376,N_35668);
and U37694 (N_37694,N_35186,N_35738);
nor U37695 (N_37695,N_36078,N_35790);
and U37696 (N_37696,N_35026,N_36736);
or U37697 (N_37697,N_36367,N_35215);
and U37698 (N_37698,N_37324,N_36145);
nor U37699 (N_37699,N_35820,N_37433);
or U37700 (N_37700,N_37453,N_36082);
nand U37701 (N_37701,N_35390,N_37327);
or U37702 (N_37702,N_36996,N_37117);
nand U37703 (N_37703,N_35326,N_37334);
or U37704 (N_37704,N_35299,N_35223);
or U37705 (N_37705,N_35960,N_36537);
nand U37706 (N_37706,N_37087,N_37478);
and U37707 (N_37707,N_37211,N_35147);
nand U37708 (N_37708,N_35521,N_35644);
nor U37709 (N_37709,N_37353,N_37341);
and U37710 (N_37710,N_36664,N_36100);
nand U37711 (N_37711,N_35546,N_35381);
nand U37712 (N_37712,N_36560,N_36708);
or U37713 (N_37713,N_37037,N_36645);
nand U37714 (N_37714,N_35082,N_36220);
nor U37715 (N_37715,N_36878,N_36959);
nand U37716 (N_37716,N_35409,N_35800);
xnor U37717 (N_37717,N_35982,N_36275);
and U37718 (N_37718,N_37294,N_35453);
and U37719 (N_37719,N_36025,N_35746);
and U37720 (N_37720,N_36028,N_35469);
or U37721 (N_37721,N_36657,N_36612);
nor U37722 (N_37722,N_35689,N_35075);
or U37723 (N_37723,N_35728,N_36809);
or U37724 (N_37724,N_35366,N_35770);
nand U37725 (N_37725,N_36841,N_36592);
nand U37726 (N_37726,N_37115,N_35170);
nor U37727 (N_37727,N_36076,N_37099);
nor U37728 (N_37728,N_37264,N_37255);
nand U37729 (N_37729,N_35987,N_35831);
and U37730 (N_37730,N_35249,N_35301);
nor U37731 (N_37731,N_35733,N_36354);
or U37732 (N_37732,N_36038,N_37180);
or U37733 (N_37733,N_36839,N_35707);
xnor U37734 (N_37734,N_36883,N_37195);
nand U37735 (N_37735,N_37034,N_36257);
nand U37736 (N_37736,N_35051,N_37482);
and U37737 (N_37737,N_35330,N_35188);
or U37738 (N_37738,N_35994,N_35120);
and U37739 (N_37739,N_35584,N_36946);
xnor U37740 (N_37740,N_35293,N_35272);
nand U37741 (N_37741,N_36829,N_35125);
xnor U37742 (N_37742,N_37463,N_36615);
and U37743 (N_37743,N_35807,N_36213);
nor U37744 (N_37744,N_35571,N_37104);
nor U37745 (N_37745,N_36500,N_35115);
nor U37746 (N_37746,N_35676,N_36583);
and U37747 (N_37747,N_37124,N_35773);
xor U37748 (N_37748,N_36222,N_36823);
or U37749 (N_37749,N_37292,N_36420);
and U37750 (N_37750,N_36195,N_35697);
or U37751 (N_37751,N_36990,N_36284);
and U37752 (N_37752,N_36306,N_36085);
or U37753 (N_37753,N_35269,N_35140);
nor U37754 (N_37754,N_37449,N_35150);
nand U37755 (N_37755,N_35031,N_35531);
and U37756 (N_37756,N_35136,N_36429);
nand U37757 (N_37757,N_35849,N_36483);
nor U37758 (N_37758,N_37499,N_35460);
and U37759 (N_37759,N_35265,N_35205);
or U37760 (N_37760,N_37498,N_36317);
nand U37761 (N_37761,N_36397,N_37222);
and U37762 (N_37762,N_36286,N_36329);
nand U37763 (N_37763,N_36037,N_35700);
nand U37764 (N_37764,N_36541,N_35466);
nand U37765 (N_37765,N_35553,N_35817);
nand U37766 (N_37766,N_36789,N_36734);
and U37767 (N_37767,N_36813,N_37444);
and U37768 (N_37768,N_35910,N_36042);
xor U37769 (N_37769,N_36617,N_35134);
or U37770 (N_37770,N_37097,N_37247);
nand U37771 (N_37771,N_36044,N_35667);
or U37772 (N_37772,N_36336,N_35289);
xor U37773 (N_37773,N_36763,N_36646);
nand U37774 (N_37774,N_37301,N_35996);
and U37775 (N_37775,N_35113,N_35701);
xnor U37776 (N_37776,N_35542,N_35392);
and U37777 (N_37777,N_35515,N_37270);
nand U37778 (N_37778,N_36274,N_35633);
or U37779 (N_37779,N_36206,N_35507);
xor U37780 (N_37780,N_36410,N_37364);
nor U37781 (N_37781,N_36532,N_37466);
and U37782 (N_37782,N_36827,N_35596);
xnor U37783 (N_37783,N_36021,N_37372);
or U37784 (N_37784,N_35905,N_36670);
nor U37785 (N_37785,N_35609,N_37151);
and U37786 (N_37786,N_37305,N_36402);
or U37787 (N_37787,N_35199,N_36672);
xor U37788 (N_37788,N_35245,N_36292);
nor U37789 (N_37789,N_36027,N_37239);
xnor U37790 (N_37790,N_35489,N_36631);
xnor U37791 (N_37791,N_36191,N_36474);
or U37792 (N_37792,N_36266,N_36816);
nand U37793 (N_37793,N_36983,N_36488);
xnor U37794 (N_37794,N_37352,N_35578);
nand U37795 (N_37795,N_36460,N_35153);
and U37796 (N_37796,N_35840,N_36819);
or U37797 (N_37797,N_36992,N_37345);
xnor U37798 (N_37798,N_36414,N_36898);
nor U37799 (N_37799,N_36046,N_35630);
and U37800 (N_37800,N_35433,N_35743);
nand U37801 (N_37801,N_36593,N_36189);
or U37802 (N_37802,N_36219,N_36957);
xor U37803 (N_37803,N_35776,N_36283);
xor U37804 (N_37804,N_36475,N_36211);
nand U37805 (N_37805,N_37045,N_37388);
xnor U37806 (N_37806,N_36157,N_37046);
nand U37807 (N_37807,N_35490,N_36130);
nand U37808 (N_37808,N_36826,N_35267);
or U37809 (N_37809,N_37176,N_36947);
nand U37810 (N_37810,N_36901,N_35655);
nor U37811 (N_37811,N_35621,N_35291);
or U37812 (N_37812,N_37277,N_36914);
or U37813 (N_37813,N_37075,N_36938);
xor U37814 (N_37814,N_36554,N_35373);
nor U37815 (N_37815,N_36862,N_37186);
xnor U37816 (N_37816,N_36411,N_36716);
nand U37817 (N_37817,N_35843,N_36034);
xnor U37818 (N_37818,N_36667,N_35344);
xor U37819 (N_37819,N_35094,N_35517);
and U37820 (N_37820,N_35907,N_36844);
nor U37821 (N_37821,N_36115,N_35880);
nor U37822 (N_37822,N_37259,N_36405);
and U37823 (N_37823,N_36728,N_36780);
nor U37824 (N_37824,N_35736,N_36740);
nand U37825 (N_37825,N_36895,N_36589);
nor U37826 (N_37826,N_36064,N_35364);
or U37827 (N_37827,N_35005,N_37067);
nand U37828 (N_37828,N_35040,N_35193);
or U37829 (N_37829,N_35320,N_36558);
xor U37830 (N_37830,N_36950,N_37481);
nor U37831 (N_37831,N_37450,N_37220);
or U37832 (N_37832,N_36205,N_37145);
nand U37833 (N_37833,N_35591,N_36815);
xor U37834 (N_37834,N_37336,N_36575);
and U37835 (N_37835,N_35001,N_35924);
nor U37836 (N_37836,N_36339,N_36192);
and U37837 (N_37837,N_35449,N_35247);
nand U37838 (N_37838,N_35866,N_36910);
nor U37839 (N_37839,N_35076,N_36998);
nor U37840 (N_37840,N_35967,N_36523);
nor U37841 (N_37841,N_35053,N_35336);
nand U37842 (N_37842,N_35262,N_37098);
or U37843 (N_37843,N_36389,N_36663);
or U37844 (N_37844,N_37391,N_35213);
and U37845 (N_37845,N_36611,N_36539);
or U37846 (N_37846,N_35435,N_36466);
nor U37847 (N_37847,N_36679,N_35098);
and U37848 (N_37848,N_35604,N_37200);
xor U37849 (N_37849,N_36571,N_36515);
nor U37850 (N_37850,N_36525,N_36198);
xor U37851 (N_37851,N_35117,N_36409);
nor U37852 (N_37852,N_36836,N_36871);
nand U37853 (N_37853,N_35953,N_36293);
and U37854 (N_37854,N_37116,N_36422);
and U37855 (N_37855,N_36758,N_37392);
nand U37856 (N_37856,N_35493,N_37137);
nor U37857 (N_37857,N_35497,N_35780);
nand U37858 (N_37858,N_35057,N_36098);
xnor U37859 (N_37859,N_35530,N_37465);
nand U37860 (N_37860,N_36842,N_37089);
xor U37861 (N_37861,N_36797,N_35421);
and U37862 (N_37862,N_36720,N_37021);
nand U37863 (N_37863,N_36102,N_35343);
and U37864 (N_37864,N_35942,N_36737);
nand U37865 (N_37865,N_36018,N_36104);
xor U37866 (N_37866,N_36359,N_35876);
nor U37867 (N_37867,N_36335,N_36079);
and U37868 (N_37868,N_35105,N_35391);
and U37869 (N_37869,N_35708,N_35902);
nor U37870 (N_37870,N_37234,N_37112);
or U37871 (N_37871,N_36529,N_36399);
or U37872 (N_37872,N_36622,N_37400);
xnor U37873 (N_37873,N_37063,N_36303);
and U37874 (N_37874,N_37056,N_36712);
xor U37875 (N_37875,N_35363,N_37312);
or U37876 (N_37876,N_36711,N_35956);
and U37877 (N_37877,N_35152,N_37258);
xor U37878 (N_37878,N_36428,N_37446);
nand U37879 (N_37879,N_35878,N_36408);
or U37880 (N_37880,N_35455,N_35275);
nand U37881 (N_37881,N_36105,N_37282);
and U37882 (N_37882,N_35036,N_36927);
and U37883 (N_37883,N_36278,N_36407);
or U37884 (N_37884,N_35812,N_37208);
or U37885 (N_37885,N_37224,N_35498);
nor U37886 (N_37886,N_35875,N_35240);
nor U37887 (N_37887,N_36223,N_36857);
or U37888 (N_37888,N_36066,N_36680);
nand U37889 (N_37889,N_35059,N_35268);
nor U37890 (N_37890,N_36920,N_35184);
nand U37891 (N_37891,N_36973,N_37078);
xnor U37892 (N_37892,N_35402,N_37265);
or U37893 (N_37893,N_36832,N_37448);
or U37894 (N_37894,N_36294,N_37248);
xnor U37895 (N_37895,N_36786,N_35835);
and U37896 (N_37896,N_37207,N_35845);
xor U37897 (N_37897,N_35901,N_37360);
nand U37898 (N_37898,N_36094,N_35771);
nand U37899 (N_37899,N_35470,N_35397);
nand U37900 (N_37900,N_37347,N_36252);
or U37901 (N_37901,N_36940,N_36099);
xnor U37902 (N_37902,N_36276,N_36967);
nor U37903 (N_37903,N_35463,N_37004);
nor U37904 (N_37904,N_36377,N_36723);
xor U37905 (N_37905,N_36134,N_37171);
or U37906 (N_37906,N_37003,N_37191);
or U37907 (N_37907,N_35151,N_35306);
or U37908 (N_37908,N_37083,N_36295);
xor U37909 (N_37909,N_37366,N_36775);
xor U37910 (N_37910,N_36981,N_36553);
or U37911 (N_37911,N_36650,N_37050);
nand U37912 (N_37912,N_35973,N_36512);
or U37913 (N_37913,N_36545,N_35587);
nor U37914 (N_37914,N_35395,N_36665);
nor U37915 (N_37915,N_35756,N_36465);
nand U37916 (N_37916,N_35505,N_35423);
or U37917 (N_37917,N_36696,N_35635);
and U37918 (N_37918,N_36877,N_36052);
xnor U37919 (N_37919,N_37316,N_37060);
nand U37920 (N_37920,N_36655,N_35173);
xor U37921 (N_37921,N_35916,N_35552);
or U37922 (N_37922,N_37118,N_35919);
and U37923 (N_37923,N_37091,N_37418);
nor U37924 (N_37924,N_37344,N_35224);
xor U37925 (N_37925,N_36116,N_35810);
nor U37926 (N_37926,N_36563,N_37475);
or U37927 (N_37927,N_35417,N_35822);
and U37928 (N_37928,N_36831,N_35030);
nand U37929 (N_37929,N_37121,N_36029);
or U37930 (N_37930,N_35127,N_35922);
nor U37931 (N_37931,N_36406,N_35908);
xor U37932 (N_37932,N_35983,N_36261);
nor U37933 (N_37933,N_35480,N_35331);
xnor U37934 (N_37934,N_35420,N_35618);
nor U37935 (N_37935,N_35185,N_36979);
nand U37936 (N_37936,N_35624,N_36521);
nor U37937 (N_37937,N_36993,N_35142);
xor U37938 (N_37938,N_35376,N_35204);
nand U37939 (N_37939,N_36127,N_35642);
or U37940 (N_37940,N_37088,N_35714);
nand U37941 (N_37941,N_37362,N_37043);
or U37942 (N_37942,N_35934,N_36290);
xor U37943 (N_37943,N_36476,N_37404);
nor U37944 (N_37944,N_35010,N_35547);
and U37945 (N_37945,N_37196,N_37160);
and U37946 (N_37946,N_35725,N_36653);
nand U37947 (N_37947,N_36061,N_35869);
xnor U37948 (N_37948,N_37014,N_36698);
nor U37949 (N_37949,N_35750,N_35677);
xnor U37950 (N_37950,N_36351,N_36089);
xor U37951 (N_37951,N_36621,N_37261);
and U37952 (N_37952,N_35365,N_36444);
or U37953 (N_37953,N_36971,N_37235);
and U37954 (N_37954,N_35887,N_36925);
nand U37955 (N_37955,N_36505,N_36380);
xnor U37956 (N_37956,N_35457,N_36260);
nor U37957 (N_37957,N_37262,N_36254);
or U37958 (N_37958,N_36771,N_36854);
and U37959 (N_37959,N_37152,N_35788);
nor U37960 (N_37960,N_35683,N_35941);
xor U37961 (N_37961,N_37315,N_36830);
and U37962 (N_37962,N_36156,N_35248);
or U37963 (N_37963,N_37325,N_35998);
nor U37964 (N_37964,N_35270,N_35829);
and U37965 (N_37965,N_35957,N_37147);
xor U37966 (N_37966,N_35300,N_35933);
and U37967 (N_37967,N_37030,N_35648);
nor U37968 (N_37968,N_35741,N_35129);
or U37969 (N_37969,N_37390,N_36263);
nor U37970 (N_37970,N_35454,N_36494);
xor U37971 (N_37971,N_35037,N_35558);
or U37972 (N_37972,N_36824,N_35589);
nand U37973 (N_37973,N_35445,N_35898);
xnor U37974 (N_37974,N_35532,N_35342);
xor U37975 (N_37975,N_36872,N_35966);
or U37976 (N_37976,N_36229,N_35110);
nor U37977 (N_37977,N_36045,N_37298);
xnor U37978 (N_37978,N_35640,N_37363);
nand U37979 (N_37979,N_36808,N_36688);
nor U37980 (N_37980,N_35029,N_35681);
or U37981 (N_37981,N_36442,N_35296);
and U37982 (N_37982,N_35244,N_35639);
and U37983 (N_37983,N_35073,N_37101);
nor U37984 (N_37984,N_36403,N_35610);
nor U37985 (N_37985,N_37379,N_36489);
nor U37986 (N_37986,N_36911,N_35605);
or U37987 (N_37987,N_35657,N_37242);
and U37988 (N_37988,N_36889,N_36587);
nand U37989 (N_37989,N_35860,N_36709);
and U37990 (N_37990,N_36852,N_35844);
nand U37991 (N_37991,N_37452,N_37253);
nor U37992 (N_37992,N_35755,N_36875);
xnor U37993 (N_37993,N_36150,N_36508);
nand U37994 (N_37994,N_36051,N_36133);
or U37995 (N_37995,N_37062,N_37048);
nor U37996 (N_37996,N_36360,N_35789);
nor U37997 (N_37997,N_35917,N_36256);
nand U37998 (N_37998,N_35442,N_36790);
nor U37999 (N_37999,N_37053,N_36574);
nor U38000 (N_38000,N_36536,N_37339);
nand U38001 (N_38001,N_35039,N_35637);
nand U38002 (N_38002,N_36165,N_35912);
nor U38003 (N_38003,N_35961,N_35705);
nor U38004 (N_38004,N_35634,N_35382);
xor U38005 (N_38005,N_37074,N_35815);
or U38006 (N_38006,N_37064,N_35232);
and U38007 (N_38007,N_35243,N_35375);
xor U38008 (N_38008,N_37192,N_35201);
nand U38009 (N_38009,N_36168,N_37393);
nor U38010 (N_38010,N_35279,N_35126);
or U38011 (N_38011,N_36695,N_36580);
nor U38012 (N_38012,N_37212,N_36114);
nor U38013 (N_38013,N_37436,N_35964);
or U38014 (N_38014,N_36008,N_35258);
and U38015 (N_38015,N_35981,N_36770);
or U38016 (N_38016,N_35305,N_37080);
xnor U38017 (N_38017,N_36289,N_35468);
xor U38018 (N_38018,N_36968,N_35485);
xnor U38019 (N_38019,N_36937,N_36485);
nand U38020 (N_38020,N_35623,N_36492);
nor U38021 (N_38021,N_35864,N_36171);
or U38022 (N_38022,N_36777,N_35011);
xnor U38023 (N_38023,N_36666,N_36597);
nand U38024 (N_38024,N_36426,N_36110);
nand U38025 (N_38025,N_35288,N_36470);
nor U38026 (N_38026,N_37132,N_36733);
nor U38027 (N_38027,N_36520,N_36764);
nor U38028 (N_38028,N_36112,N_35737);
xnor U38029 (N_38029,N_35144,N_35814);
and U38030 (N_38030,N_35241,N_36903);
nand U38031 (N_38031,N_35239,N_35846);
xor U38032 (N_38032,N_36067,N_36855);
nand U38033 (N_38033,N_36608,N_36975);
xnor U38034 (N_38034,N_35135,N_36744);
and U38035 (N_38035,N_36022,N_37268);
xnor U38036 (N_38036,N_37441,N_36337);
xnor U38037 (N_38037,N_35298,N_37423);
or U38038 (N_38038,N_36461,N_35091);
xor U38039 (N_38039,N_35911,N_37395);
nand U38040 (N_38040,N_36228,N_37295);
or U38041 (N_38041,N_35896,N_35237);
nand U38042 (N_38042,N_36095,N_36185);
or U38043 (N_38043,N_35959,N_35518);
xor U38044 (N_38044,N_36436,N_35067);
nand U38045 (N_38045,N_36869,N_36419);
nand U38046 (N_38046,N_37141,N_36707);
xor U38047 (N_38047,N_36448,N_35797);
nor U38048 (N_38048,N_36459,N_37069);
nand U38049 (N_38049,N_36368,N_37291);
nor U38050 (N_38050,N_36396,N_35656);
nand U38051 (N_38051,N_36879,N_36482);
and U38052 (N_38052,N_36590,N_35581);
or U38053 (N_38053,N_37406,N_36020);
or U38054 (N_38054,N_35883,N_37107);
or U38055 (N_38055,N_35602,N_36212);
and U38056 (N_38056,N_36450,N_35446);
or U38057 (N_38057,N_37001,N_36714);
nor U38058 (N_38058,N_36330,N_37461);
nand U38059 (N_38059,N_35122,N_35483);
and U38060 (N_38060,N_35281,N_37153);
and U38061 (N_38061,N_35346,N_35164);
and U38062 (N_38062,N_35206,N_35499);
nor U38063 (N_38063,N_35706,N_35338);
xnor U38064 (N_38064,N_36250,N_35765);
xor U38065 (N_38065,N_36564,N_35203);
xnor U38066 (N_38066,N_35962,N_37187);
or U38067 (N_38067,N_37483,N_36349);
nand U38068 (N_38068,N_36319,N_35318);
and U38069 (N_38069,N_35913,N_35888);
nor U38070 (N_38070,N_36447,N_35625);
nor U38071 (N_38071,N_36739,N_35551);
or U38072 (N_38072,N_35192,N_36187);
nor U38073 (N_38073,N_36350,N_35823);
and U38074 (N_38074,N_37473,N_35416);
nor U38075 (N_38075,N_36643,N_36562);
nand U38076 (N_38076,N_36487,N_35347);
xor U38077 (N_38077,N_36490,N_36190);
nand U38078 (N_38078,N_36030,N_37059);
or U38079 (N_38079,N_37486,N_36896);
xnor U38080 (N_38080,N_35220,N_35873);
nand U38081 (N_38081,N_37243,N_36599);
xor U38082 (N_38082,N_37399,N_36023);
xor U38083 (N_38083,N_36917,N_35181);
or U38084 (N_38084,N_35254,N_37320);
and U38085 (N_38085,N_36083,N_35096);
nor U38086 (N_38086,N_35653,N_35691);
xnor U38087 (N_38087,N_35168,N_37085);
nor U38088 (N_38088,N_35761,N_35311);
or U38089 (N_38089,N_36683,N_37206);
nor U38090 (N_38090,N_35321,N_36543);
or U38091 (N_38091,N_36531,N_35811);
or U38092 (N_38092,N_37346,N_36787);
and U38093 (N_38093,N_35915,N_36750);
and U38094 (N_38094,N_36070,N_37273);
and U38095 (N_38095,N_35102,N_36193);
and U38096 (N_38096,N_36633,N_35148);
xor U38097 (N_38097,N_35508,N_36113);
nor U38098 (N_38098,N_36353,N_36892);
xor U38099 (N_38099,N_35674,N_36907);
xnor U38100 (N_38100,N_37113,N_37170);
or U38101 (N_38101,N_36752,N_36549);
and U38102 (N_38102,N_35963,N_37349);
and U38103 (N_38103,N_37311,N_35695);
or U38104 (N_38104,N_36656,N_35974);
nor U38105 (N_38105,N_35687,N_37011);
xor U38106 (N_38106,N_36258,N_36671);
nand U38107 (N_38107,N_37142,N_37013);
xnor U38108 (N_38108,N_37340,N_36821);
and U38109 (N_38109,N_35786,N_36588);
and U38110 (N_38110,N_35512,N_37169);
xor U38111 (N_38111,N_37313,N_36443);
xnor U38112 (N_38112,N_36860,N_35486);
or U38113 (N_38113,N_36139,N_36296);
and U38114 (N_38114,N_35690,N_36491);
nor U38115 (N_38115,N_35475,N_37042);
and U38116 (N_38116,N_36681,N_37065);
or U38117 (N_38117,N_35143,N_37283);
nor U38118 (N_38118,N_36551,N_36194);
or U38119 (N_38119,N_37084,N_37432);
nor U38120 (N_38120,N_35294,N_35833);
and U38121 (N_38121,N_36506,N_35233);
or U38122 (N_38122,N_37038,N_37031);
nand U38123 (N_38123,N_36001,N_35012);
and U38124 (N_38124,N_35389,N_35436);
or U38125 (N_38125,N_36259,N_35495);
nand U38126 (N_38126,N_35985,N_35361);
nor U38127 (N_38127,N_36795,N_37209);
nand U38128 (N_38128,N_36908,N_36675);
nand U38129 (N_38129,N_36129,N_35827);
nor U38130 (N_38130,N_36050,N_35124);
xnor U38131 (N_38131,N_35734,N_37350);
and U38132 (N_38132,N_36245,N_36999);
or U38133 (N_38133,N_35836,N_35995);
nor U38134 (N_38134,N_36556,N_36264);
nor U38135 (N_38135,N_37111,N_35937);
nand U38136 (N_38136,N_35972,N_36288);
xnor U38137 (N_38137,N_36867,N_36160);
xnor U38138 (N_38138,N_37051,N_35928);
or U38139 (N_38139,N_35006,N_36109);
nand U38140 (N_38140,N_35471,N_35092);
and U38141 (N_38141,N_36861,N_35903);
or U38142 (N_38142,N_37410,N_36423);
nand U38143 (N_38143,N_35694,N_36432);
nand U38144 (N_38144,N_35177,N_36144);
and U38145 (N_38145,N_37434,N_35398);
nand U38146 (N_38146,N_35993,N_36535);
and U38147 (N_38147,N_35662,N_35693);
or U38148 (N_38148,N_35900,N_35593);
nor U38149 (N_38149,N_35938,N_36135);
nand U38150 (N_38150,N_37106,N_37023);
and U38151 (N_38151,N_37326,N_35452);
nor U38152 (N_38152,N_37204,N_35759);
and U38153 (N_38153,N_37333,N_36997);
nor U38154 (N_38154,N_37251,N_36960);
xnor U38155 (N_38155,N_37018,N_36224);
nor U38156 (N_38156,N_36949,N_37110);
nand U38157 (N_38157,N_36179,N_36363);
xnor U38158 (N_38158,N_35494,N_35660);
nor U38159 (N_38159,N_36888,N_36323);
xnor U38160 (N_38160,N_36010,N_35315);
or U38161 (N_38161,N_35856,N_35538);
nor U38162 (N_38162,N_37055,N_37041);
nand U38163 (N_38163,N_35367,N_36594);
xnor U38164 (N_38164,N_36794,N_35550);
xor U38165 (N_38165,N_35500,N_36926);
nor U38166 (N_38166,N_35732,N_35742);
and U38167 (N_38167,N_36056,N_36530);
or U38168 (N_38168,N_35313,N_36548);
nand U38169 (N_38169,N_36239,N_36090);
or U38170 (N_38170,N_36966,N_36610);
nand U38171 (N_38171,N_36626,N_37397);
xor U38172 (N_38172,N_36073,N_36921);
nand U38173 (N_38173,N_35615,N_35286);
or U38174 (N_38174,N_36328,N_37309);
xnor U38175 (N_38175,N_37168,N_37185);
nor U38176 (N_38176,N_36834,N_37337);
or U38177 (N_38177,N_35980,N_36961);
nand U38178 (N_38178,N_35044,N_37081);
and U38179 (N_38179,N_36300,N_37225);
and U38180 (N_38180,N_35567,N_35560);
nand U38181 (N_38181,N_36214,N_37245);
nor U38182 (N_38182,N_36075,N_35329);
xnor U38183 (N_38183,N_36801,N_35717);
nand U38184 (N_38184,N_36265,N_35025);
or U38185 (N_38185,N_35565,N_37459);
xor U38186 (N_38186,N_36304,N_36203);
nor U38187 (N_38187,N_37109,N_37439);
nor U38188 (N_38188,N_35592,N_35958);
nand U38189 (N_38189,N_37425,N_36000);
and U38190 (N_38190,N_37156,N_36291);
or U38191 (N_38191,N_35865,N_35986);
nor U38192 (N_38192,N_36713,N_36743);
or U38193 (N_38193,N_35202,N_35951);
nor U38194 (N_38194,N_36729,N_36566);
or U38195 (N_38195,N_36811,N_37375);
and U38196 (N_38196,N_35943,N_35509);
xnor U38197 (N_38197,N_35132,N_37005);
nand U38198 (N_38198,N_36935,N_36238);
nand U38199 (N_38199,N_36570,N_35696);
or U38200 (N_38200,N_37092,N_35541);
or U38201 (N_38201,N_35778,N_35432);
and U38202 (N_38202,N_36757,N_35106);
and U38203 (N_38203,N_36087,N_36793);
nor U38204 (N_38204,N_35214,N_35337);
nor U38205 (N_38205,N_37032,N_36627);
or U38206 (N_38206,N_35611,N_35710);
or U38207 (N_38207,N_37329,N_35702);
and U38208 (N_38208,N_36899,N_35622);
xnor U38209 (N_38209,N_35062,N_37260);
or U38210 (N_38210,N_37323,N_36202);
or U38211 (N_38211,N_35798,N_36404);
nor U38212 (N_38212,N_36814,N_35097);
nand U38213 (N_38213,N_36273,N_35378);
xnor U38214 (N_38214,N_37496,N_35362);
and U38215 (N_38215,N_35791,N_35909);
nor U38216 (N_38216,N_35264,N_36567);
nor U38217 (N_38217,N_35555,N_36438);
nor U38218 (N_38218,N_35228,N_37129);
nand U38219 (N_38219,N_35678,N_36746);
or U38220 (N_38220,N_35606,N_36803);
or U38221 (N_38221,N_36586,N_36944);
nand U38222 (N_38222,N_35133,N_35476);
or U38223 (N_38223,N_36885,N_36479);
xor U38224 (N_38224,N_35516,N_36644);
xor U38225 (N_38225,N_36624,N_36272);
xnor U38226 (N_38226,N_36463,N_35598);
nand U38227 (N_38227,N_36149,N_36305);
and U38228 (N_38228,N_36715,N_35540);
or U38229 (N_38229,N_36941,N_37250);
nand U38230 (N_38230,N_35799,N_35826);
or U38231 (N_38231,N_36439,N_37020);
and U38232 (N_38232,N_36172,N_36352);
nor U38233 (N_38233,N_36890,N_35825);
nand U38234 (N_38234,N_36201,N_36015);
nor U38235 (N_38235,N_35821,N_37300);
xnor U38236 (N_38236,N_36934,N_35327);
and U38237 (N_38237,N_37286,N_35501);
nand U38238 (N_38238,N_36674,N_36881);
xor U38239 (N_38239,N_36783,N_35795);
and U38240 (N_38240,N_37422,N_36123);
xnor U38241 (N_38241,N_36774,N_35712);
and U38242 (N_38242,N_36727,N_37172);
nor U38243 (N_38243,N_36965,N_35686);
and U38244 (N_38244,N_37044,N_36963);
and U38245 (N_38245,N_37314,N_35948);
and U38246 (N_38246,N_35511,N_35251);
or U38247 (N_38247,N_35839,N_36218);
and U38248 (N_38248,N_37070,N_36572);
nor U38249 (N_38249,N_36253,N_35740);
nand U38250 (N_38250,N_35673,N_36913);
or U38251 (N_38251,N_37269,N_37066);
or U38252 (N_38252,N_35600,N_36478);
xor U38253 (N_38253,N_35016,N_35897);
nor U38254 (N_38254,N_37307,N_35100);
or U38255 (N_38255,N_36421,N_35090);
or U38256 (N_38256,N_37244,N_36384);
or U38257 (N_38257,N_36503,N_37365);
nand U38258 (N_38258,N_36978,N_35443);
nand U38259 (N_38259,N_35474,N_35401);
nor U38260 (N_38260,N_36240,N_36718);
or U38261 (N_38261,N_36955,N_36471);
nor U38262 (N_38262,N_37416,N_37231);
nand U38263 (N_38263,N_35121,N_36687);
nand U38264 (N_38264,N_36163,N_35585);
nand U38265 (N_38265,N_37214,N_35641);
xnor U38266 (N_38266,N_35157,N_36710);
xor U38267 (N_38267,N_35619,N_35089);
and U38268 (N_38268,N_37414,N_35242);
xor U38269 (N_38269,N_36153,N_36662);
or U38270 (N_38270,N_37487,N_35479);
xnor U38271 (N_38271,N_35721,N_36953);
or U38272 (N_38272,N_35467,N_37120);
and U38273 (N_38273,N_35473,N_35141);
xnor U38274 (N_38274,N_36762,N_35451);
nand U38275 (N_38275,N_36241,N_36146);
nor U38276 (N_38276,N_36706,N_35282);
or U38277 (N_38277,N_35360,N_36741);
and U38278 (N_38278,N_36697,N_37163);
or U38279 (N_38279,N_35590,N_36299);
and U38280 (N_38280,N_37123,N_35688);
xnor U38281 (N_38281,N_36320,N_36118);
nor U38282 (N_38282,N_36629,N_36041);
and U38283 (N_38283,N_35412,N_35380);
nand U38284 (N_38284,N_36602,N_37287);
or U38285 (N_38285,N_35234,N_36584);
nand U38286 (N_38286,N_36601,N_35568);
xnor U38287 (N_38287,N_35719,N_37143);
and U38288 (N_38288,N_37246,N_36345);
and U38289 (N_38289,N_35128,N_36779);
or U38290 (N_38290,N_36126,N_37213);
xnor U38291 (N_38291,N_35627,N_36178);
and U38292 (N_38292,N_36208,N_36623);
and U38293 (N_38293,N_35021,N_36800);
xor U38294 (N_38294,N_35658,N_36945);
xor U38295 (N_38295,N_37492,N_35892);
nand U38296 (N_38296,N_35425,N_36689);
xor U38297 (N_38297,N_35614,N_36326);
nor U38298 (N_38298,N_35939,N_36928);
and U38299 (N_38299,N_37016,N_35936);
and U38300 (N_38300,N_35303,N_36923);
xnor U38301 (N_38301,N_36552,N_35458);
xor U38302 (N_38302,N_36555,N_35769);
nand U38303 (N_38303,N_36346,N_36017);
nand U38304 (N_38304,N_35054,N_36585);
xor U38305 (N_38305,N_36595,N_36484);
and U38306 (N_38306,N_35731,N_35255);
nor U38307 (N_38307,N_36691,N_35478);
nor U38308 (N_38308,N_37190,N_36540);
and U38309 (N_38309,N_36933,N_37061);
and U38310 (N_38310,N_37464,N_37497);
xor U38311 (N_38311,N_36235,N_35669);
xnor U38312 (N_38312,N_35146,N_36952);
nand U38313 (N_38313,N_36170,N_36246);
xnor U38314 (N_38314,N_36559,N_36340);
or U38315 (N_38315,N_35261,N_37403);
nor U38316 (N_38316,N_36799,N_36394);
xor U38317 (N_38317,N_36131,N_36918);
or U38318 (N_38318,N_36199,N_36874);
or U38319 (N_38319,N_35616,N_35093);
nand U38320 (N_38320,N_37343,N_35256);
nor U38321 (N_38321,N_37367,N_37280);
xnor U38322 (N_38322,N_36071,N_35988);
or U38323 (N_38323,N_37426,N_36722);
nand U38324 (N_38324,N_35165,N_35652);
nand U38325 (N_38325,N_36152,N_36164);
or U38326 (N_38326,N_35649,N_35043);
or U38327 (N_38327,N_36605,N_35049);
nand U38328 (N_38328,N_37266,N_35762);
or U38329 (N_38329,N_36954,N_36200);
and U38330 (N_38330,N_36480,N_35095);
and U38331 (N_38331,N_36361,N_36761);
nor U38332 (N_38332,N_37166,N_36356);
nor U38333 (N_38333,N_36481,N_36703);
xnor U38334 (N_38334,N_35607,N_36457);
xor U38335 (N_38335,N_35659,N_37419);
nor U38336 (N_38336,N_36522,N_37405);
xor U38337 (N_38337,N_35277,N_35116);
and U38338 (N_38338,N_36324,N_36856);
and U38339 (N_38339,N_36468,N_35863);
nor U38340 (N_38340,N_36280,N_37351);
nand U38341 (N_38341,N_36804,N_36828);
nor U38342 (N_38342,N_37238,N_35647);
or U38343 (N_38343,N_35310,N_36620);
nand U38344 (N_38344,N_35748,N_36467);
nor U38345 (N_38345,N_36932,N_36598);
nor U38346 (N_38346,N_35582,N_35976);
or U38347 (N_38347,N_35984,N_36886);
or U38348 (N_38348,N_36147,N_35675);
nand U38349 (N_38349,N_35107,N_36850);
or U38350 (N_38350,N_36822,N_35405);
xnor U38351 (N_38351,N_35768,N_36327);
or U38352 (N_38352,N_36390,N_35379);
nor U38353 (N_38353,N_35070,N_35211);
or U38354 (N_38354,N_35008,N_36313);
nand U38355 (N_38355,N_36391,N_35613);
and U38356 (N_38356,N_37228,N_36344);
xor U38357 (N_38357,N_35779,N_37409);
nor U38358 (N_38358,N_37173,N_37240);
and U38359 (N_38359,N_37241,N_36693);
nor U38360 (N_38360,N_36312,N_35348);
or U38361 (N_38361,N_36504,N_36049);
or U38362 (N_38362,N_37024,N_36765);
or U38363 (N_38363,N_36418,N_37495);
xnor U38364 (N_38364,N_36108,N_36876);
or U38365 (N_38365,N_36792,N_37355);
or U38366 (N_38366,N_37119,N_36704);
xnor U38367 (N_38367,N_35536,N_36730);
xor U38368 (N_38368,N_35061,N_36400);
xnor U38369 (N_38369,N_35083,N_36561);
nand U38370 (N_38370,N_36269,N_37249);
xnor U38371 (N_38371,N_36513,N_37165);
nand U38372 (N_38372,N_36233,N_36154);
nand U38373 (N_38373,N_36433,N_35899);
xnor U38374 (N_38374,N_35427,N_35932);
and U38375 (N_38375,N_37058,N_35078);
xor U38376 (N_38376,N_37219,N_36124);
nand U38377 (N_38377,N_35599,N_36725);
nand U38378 (N_38378,N_35028,N_37028);
or U38379 (N_38379,N_36692,N_35217);
and U38380 (N_38380,N_35156,N_37188);
nand U38381 (N_38381,N_36882,N_35730);
or U38382 (N_38382,N_35620,N_35137);
nor U38383 (N_38383,N_35112,N_36632);
and U38384 (N_38384,N_36652,N_36314);
nand U38385 (N_38385,N_35852,N_36528);
and U38386 (N_38386,N_36640,N_35931);
nand U38387 (N_38387,N_37440,N_35084);
or U38388 (N_38388,N_36768,N_36088);
and U38389 (N_38389,N_35808,N_36392);
nor U38390 (N_38390,N_35805,N_36084);
nor U38391 (N_38391,N_36207,N_36315);
xor U38392 (N_38392,N_37429,N_36805);
xnor U38393 (N_38393,N_35086,N_37140);
xor U38394 (N_38394,N_36951,N_35774);
xnor U38395 (N_38395,N_37181,N_37090);
xnor U38396 (N_38396,N_36174,N_36301);
nor U38397 (N_38397,N_35871,N_35629);
xnor U38398 (N_38398,N_36991,N_37229);
nor U38399 (N_38399,N_37022,N_36177);
or U38400 (N_38400,N_37474,N_37009);
xor U38401 (N_38401,N_37317,N_37178);
nor U38402 (N_38402,N_36767,N_35527);
nor U38403 (N_38403,N_36004,N_37398);
and U38404 (N_38404,N_37293,N_35422);
nand U38405 (N_38405,N_36748,N_35297);
or U38406 (N_38406,N_37428,N_35729);
or U38407 (N_38407,N_36636,N_35046);
nor U38408 (N_38408,N_35459,N_37493);
or U38409 (N_38409,N_36519,N_37197);
nor U38410 (N_38410,N_36884,N_36576);
or U38411 (N_38411,N_37136,N_35349);
nor U38412 (N_38412,N_36060,N_36437);
xor U38413 (N_38413,N_35716,N_37072);
nor U38414 (N_38414,N_35954,N_35573);
nor U38415 (N_38415,N_36173,N_35850);
or U38416 (N_38416,N_36930,N_36188);
nor U38417 (N_38417,N_35890,N_36341);
xor U38418 (N_38418,N_35103,N_35914);
or U38419 (N_38419,N_37000,N_35461);
xor U38420 (N_38420,N_35940,N_35502);
nand U38421 (N_38421,N_35191,N_36912);
nand U38422 (N_38422,N_36782,N_36669);
nand U38423 (N_38423,N_36738,N_35314);
nor U38424 (N_38424,N_36271,N_37184);
nor U38425 (N_38425,N_36121,N_35566);
nor U38426 (N_38426,N_37019,N_35159);
nor U38427 (N_38427,N_36242,N_36582);
and U38428 (N_38428,N_37427,N_35218);
nor U38429 (N_38429,N_36760,N_36784);
and U38430 (N_38430,N_35990,N_35007);
or U38431 (N_38431,N_36430,N_36318);
or U38432 (N_38432,N_36378,N_36843);
nand U38433 (N_38433,N_36072,N_36717);
xnor U38434 (N_38434,N_35563,N_35920);
nor U38435 (N_38435,N_37382,N_35543);
and U38436 (N_38436,N_35504,N_36155);
nand U38437 (N_38437,N_36182,N_37017);
xor U38438 (N_38438,N_35782,N_35965);
or U38439 (N_38439,N_36215,N_35775);
xnor U38440 (N_38440,N_36251,N_35383);
or U38441 (N_38441,N_36416,N_35333);
nand U38442 (N_38442,N_35227,N_35000);
and U38443 (N_38443,N_36024,N_37306);
and U38444 (N_38444,N_35345,N_37149);
or U38445 (N_38445,N_35785,N_35175);
xor U38446 (N_38446,N_36972,N_36649);
or U38447 (N_38447,N_35570,N_35519);
and U38448 (N_38448,N_36458,N_36143);
xnor U38449 (N_38449,N_36381,N_36887);
nand U38450 (N_38450,N_35323,N_36820);
and U38451 (N_38451,N_36048,N_37469);
or U38452 (N_38452,N_36106,N_35650);
or U38453 (N_38453,N_35858,N_35921);
nor U38454 (N_38454,N_37371,N_36853);
or U38455 (N_38455,N_35130,N_35077);
or U38456 (N_38456,N_37369,N_35802);
xnor U38457 (N_38457,N_36616,N_37162);
nor U38458 (N_38458,N_35699,N_35524);
or U38459 (N_38459,N_37194,N_37036);
nor U38460 (N_38460,N_37407,N_35027);
xnor U38461 (N_38461,N_37096,N_35816);
nor U38462 (N_38462,N_36383,N_37025);
nor U38463 (N_38463,N_35440,N_35372);
or U38464 (N_38464,N_36802,N_35079);
or U38465 (N_38465,N_36158,N_36279);
and U38466 (N_38466,N_35209,N_36136);
or U38467 (N_38467,N_36002,N_37421);
nor U38468 (N_38468,N_36142,N_37161);
or U38469 (N_38469,N_37135,N_35764);
nand U38470 (N_38470,N_35319,N_37139);
xnor U38471 (N_38471,N_35334,N_36550);
nor U38472 (N_38472,N_36573,N_36994);
and U38473 (N_38473,N_35946,N_37396);
or U38474 (N_38474,N_35715,N_35374);
xnor U38475 (N_38475,N_36005,N_36270);
and U38476 (N_38476,N_36825,N_35198);
xnor U38477 (N_38477,N_37276,N_36778);
or U38478 (N_38478,N_36647,N_35564);
and U38479 (N_38479,N_36648,N_37338);
or U38480 (N_38480,N_35651,N_36204);
xor U38481 (N_38481,N_36395,N_35257);
xor U38482 (N_38482,N_35145,N_35169);
and U38483 (N_38483,N_37328,N_36379);
and U38484 (N_38484,N_36974,N_36807);
nand U38485 (N_38485,N_36581,N_35087);
xor U38486 (N_38486,N_35210,N_35208);
nor U38487 (N_38487,N_36557,N_36454);
nand U38488 (N_38488,N_35104,N_36732);
xnor U38489 (N_38489,N_36081,N_35867);
nand U38490 (N_38490,N_36244,N_35065);
xor U38491 (N_38491,N_35491,N_37412);
nand U38492 (N_38492,N_37183,N_36980);
nand U38493 (N_38493,N_35441,N_35703);
xor U38494 (N_38494,N_36915,N_35488);
and U38495 (N_38495,N_35032,N_36180);
and U38496 (N_38496,N_35009,N_35682);
or U38497 (N_38497,N_36332,N_37332);
or U38498 (N_38498,N_37077,N_36514);
and U38499 (N_38499,N_36989,N_37370);
or U38500 (N_38500,N_35357,N_36618);
nand U38501 (N_38501,N_36281,N_35386);
or U38502 (N_38502,N_35537,N_35661);
xnor U38503 (N_38503,N_36176,N_36678);
nand U38504 (N_38504,N_35287,N_36117);
nor U38505 (N_38505,N_36517,N_36101);
xor U38506 (N_38506,N_36511,N_37201);
nor U38507 (N_38507,N_36905,N_36970);
nor U38508 (N_38508,N_36866,N_37217);
xnor U38509 (N_38509,N_36705,N_36054);
xor U38510 (N_38510,N_36325,N_35842);
and U38511 (N_38511,N_37210,N_35523);
nand U38512 (N_38512,N_35434,N_35767);
nand U38513 (N_38513,N_35792,N_35806);
nand U38514 (N_38514,N_37049,N_35893);
xor U38515 (N_38515,N_35464,N_37284);
nor U38516 (N_38516,N_35588,N_37008);
or U38517 (N_38517,N_37281,N_35219);
or U38518 (N_38518,N_35783,N_37458);
nand U38519 (N_38519,N_35853,N_36209);
nand U38520 (N_38520,N_36906,N_35222);
or U38521 (N_38521,N_35283,N_35295);
nor U38522 (N_38522,N_35549,N_37164);
nand U38523 (N_38523,N_36369,N_36249);
and U38524 (N_38524,N_35447,N_37376);
or U38525 (N_38525,N_35945,N_36277);
nor U38526 (N_38526,N_37488,N_35285);
and U38527 (N_38527,N_35801,N_37189);
or U38528 (N_38528,N_35377,N_36840);
xor U38529 (N_38529,N_35670,N_35424);
nor U38530 (N_38530,N_35522,N_35190);
nand U38531 (N_38531,N_36654,N_35970);
and U38532 (N_38532,N_36058,N_37437);
and U38533 (N_38533,N_36348,N_36230);
nor U38534 (N_38534,N_36148,N_35777);
nor U38535 (N_38535,N_37126,N_37159);
nand U38536 (N_38536,N_37331,N_36316);
nand U38537 (N_38537,N_35997,N_37490);
nand U38538 (N_38538,N_35556,N_36477);
xor U38539 (N_38539,N_35274,N_35131);
nand U38540 (N_38540,N_36769,N_35992);
xor U38541 (N_38541,N_36759,N_35745);
nor U38542 (N_38542,N_36370,N_37361);
or U38543 (N_38543,N_35889,N_35074);
and U38544 (N_38544,N_36818,N_36606);
xor U38545 (N_38545,N_37285,N_36122);
or U38546 (N_38546,N_36462,N_37402);
and U38547 (N_38547,N_36988,N_35557);
and U38548 (N_38548,N_35304,N_37386);
and U38549 (N_38549,N_36607,N_37274);
or U38550 (N_38550,N_36637,N_35163);
nor U38551 (N_38551,N_35166,N_36639);
and U38552 (N_38552,N_36939,N_36417);
or U38553 (N_38553,N_36069,N_36234);
and U38554 (N_38554,N_35514,N_36699);
and U38555 (N_38555,N_35340,N_36600);
xor U38556 (N_38556,N_37052,N_36186);
nor U38557 (N_38557,N_35353,N_36544);
nand U38558 (N_38558,N_37175,N_36628);
nor U38559 (N_38559,N_35704,N_35872);
nor U38560 (N_38560,N_36137,N_37202);
nand U38561 (N_38561,N_36107,N_35060);
nor U38562 (N_38562,N_36788,N_35114);
or U38563 (N_38563,N_35196,N_35171);
and U38564 (N_38564,N_36817,N_36619);
or U38565 (N_38565,N_35450,N_35235);
or U38566 (N_38566,N_37417,N_35048);
nand U38567 (N_38567,N_36183,N_35787);
nand U38568 (N_38568,N_37445,N_36455);
nand U38569 (N_38569,N_36749,N_35444);
and U38570 (N_38570,N_37073,N_35187);
nand U38571 (N_38571,N_37368,N_35399);
or U38572 (N_38572,N_36285,N_37385);
or U38573 (N_38573,N_37047,N_37122);
xor U38574 (N_38574,N_36334,N_37356);
nor U38575 (N_38575,N_36357,N_35881);
nand U38576 (N_38576,N_36297,N_35022);
xnor U38577 (N_38577,N_35316,N_37114);
or U38578 (N_38578,N_35263,N_36486);
xnor U38579 (N_38579,N_35290,N_36772);
nand U38580 (N_38580,N_36995,N_36849);
nand U38581 (N_38581,N_37236,N_36343);
and U38582 (N_38582,N_37040,N_37027);
nor U38583 (N_38583,N_37144,N_36016);
or U38584 (N_38584,N_36931,N_36125);
nand U38585 (N_38585,N_35809,N_36227);
xnor U38586 (N_38586,N_35038,N_36386);
nand U38587 (N_38587,N_36958,N_37054);
nor U38588 (N_38588,N_35484,N_35195);
and U38589 (N_38589,N_36700,N_37226);
and U38590 (N_38590,N_36425,N_35506);
or U38591 (N_38591,N_35414,N_37125);
and U38592 (N_38592,N_35559,N_36499);
or U38593 (N_38593,N_36365,N_35617);
nand U38594 (N_38594,N_35926,N_37221);
xor U38595 (N_38595,N_35058,N_36833);
and U38596 (N_38596,N_35088,N_36668);
nand U38597 (N_38597,N_36231,N_36007);
xor U38598 (N_38598,N_35226,N_35407);
xor U38599 (N_38599,N_35033,N_35569);
nand U38600 (N_38600,N_36578,N_37384);
nand U38601 (N_38601,N_36347,N_36846);
or U38602 (N_38602,N_35760,N_36012);
nand U38603 (N_38603,N_36086,N_37257);
and U38604 (N_38604,N_37380,N_36916);
nor U38605 (N_38605,N_35828,N_35332);
nor U38606 (N_38606,N_37093,N_36673);
nand U38607 (N_38607,N_35894,N_37252);
nand U38608 (N_38608,N_37150,N_36446);
xnor U38609 (N_38609,N_35525,N_35492);
or U38610 (N_38610,N_35017,N_36043);
nand U38611 (N_38611,N_35528,N_37413);
and U38612 (N_38612,N_36036,N_37438);
xnor U38613 (N_38613,N_37484,N_36236);
and U38614 (N_38614,N_35636,N_35359);
nand U38615 (N_38615,N_36873,N_35064);
xnor U38616 (N_38616,N_35419,N_36776);
or U38617 (N_38617,N_36031,N_37310);
nand U38618 (N_38618,N_36440,N_36660);
nand U38619 (N_38619,N_36613,N_35711);
or U38620 (N_38620,N_36929,N_36900);
or U38621 (N_38621,N_36614,N_36870);
nor U38622 (N_38622,N_35413,N_35848);
nor U38623 (N_38623,N_36026,N_35099);
nand U38624 (N_38624,N_37095,N_35794);
or U38625 (N_38625,N_35335,N_35052);
and U38626 (N_38626,N_35111,N_35292);
xnor U38627 (N_38627,N_36308,N_37435);
nand U38628 (N_38628,N_36393,N_35350);
xnor U38629 (N_38629,N_37456,N_35989);
nor U38630 (N_38630,N_35384,N_35947);
nand U38631 (N_38631,N_36373,N_36141);
and U38632 (N_38632,N_37215,N_37319);
xor U38633 (N_38633,N_36579,N_37128);
nand U38634 (N_38634,N_36806,N_36685);
xor U38635 (N_38635,N_37411,N_36464);
nand U38636 (N_38636,N_36526,N_35882);
xnor U38637 (N_38637,N_35221,N_36812);
nand U38638 (N_38638,N_35561,N_35574);
xnor U38639 (N_38639,N_36080,N_36302);
nand U38640 (N_38640,N_35744,N_36375);
and U38641 (N_38641,N_36785,N_36964);
or U38642 (N_38642,N_35991,N_35628);
nor U38643 (N_38643,N_36495,N_35013);
nor U38644 (N_38644,N_37330,N_37290);
xnor U38645 (N_38645,N_36287,N_37470);
xnor U38646 (N_38646,N_36851,N_35838);
xor U38647 (N_38647,N_35608,N_36068);
nor U38648 (N_38648,N_35747,N_35154);
nand U38649 (N_38649,N_36516,N_35371);
or U38650 (N_38650,N_35804,N_37167);
nand U38651 (N_38651,N_35904,N_35003);
nor U38652 (N_38652,N_35162,N_37467);
nor U38653 (N_38653,N_36221,N_37491);
xnor U38654 (N_38654,N_36237,N_37342);
nand U38655 (N_38655,N_35572,N_35709);
or U38656 (N_38656,N_35885,N_36942);
or U38657 (N_38657,N_35400,N_35200);
and U38658 (N_38658,N_36731,N_35753);
or U38659 (N_38659,N_36181,N_35935);
or U38660 (N_38660,N_37472,N_36661);
nor U38661 (N_38661,N_36547,N_35751);
xor U38662 (N_38662,N_35793,N_35253);
nand U38663 (N_38663,N_35654,N_35072);
and U38664 (N_38664,N_35535,N_37288);
and U38665 (N_38665,N_35539,N_36243);
and U38666 (N_38666,N_35207,N_36837);
or U38667 (N_38667,N_35837,N_35758);
nand U38668 (N_38668,N_37374,N_35174);
and U38669 (N_38669,N_36074,N_37304);
or U38670 (N_38670,N_35431,N_37146);
nor U38671 (N_38671,N_36282,N_37476);
and U38672 (N_38672,N_36217,N_35612);
or U38673 (N_38673,N_37471,N_35969);
xor U38674 (N_38674,N_35870,N_35406);
xnor U38675 (N_38675,N_35739,N_35735);
nand U38676 (N_38676,N_37489,N_37383);
or U38677 (N_38677,N_35355,N_36773);
nand U38678 (N_38678,N_35754,N_37154);
xnor U38679 (N_38679,N_35955,N_35042);
nand U38680 (N_38680,N_35841,N_35510);
xnor U38681 (N_38681,N_35063,N_37105);
or U38682 (N_38682,N_35663,N_35189);
xor U38683 (N_38683,N_36119,N_37357);
nand U38684 (N_38684,N_36331,N_36247);
nand U38685 (N_38685,N_37223,N_36427);
nand U38686 (N_38686,N_36498,N_35562);
nor U38687 (N_38687,N_35977,N_36111);
xnor U38688 (N_38688,N_35023,N_35971);
xnor U38689 (N_38689,N_35225,N_37462);
and U38690 (N_38690,N_35718,N_35161);
and U38691 (N_38691,N_35859,N_36745);
and U38692 (N_38692,N_35055,N_36798);
nor U38693 (N_38693,N_36603,N_36864);
nor U38694 (N_38694,N_36501,N_36120);
xor U38695 (N_38695,N_35246,N_36062);
or U38696 (N_38696,N_36197,N_36415);
xnor U38697 (N_38697,N_35646,N_36445);
and U38698 (N_38698,N_35339,N_36638);
xnor U38699 (N_38699,N_35975,N_35671);
nor U38700 (N_38700,N_35438,N_35766);
and U38701 (N_38701,N_35698,N_35276);
or U38702 (N_38702,N_35727,N_35586);
or U38703 (N_38703,N_36596,N_36412);
and U38704 (N_38704,N_36796,N_37012);
nor U38705 (N_38705,N_35664,N_35317);
nand U38706 (N_38706,N_36835,N_36006);
or U38707 (N_38707,N_37335,N_37477);
xor U38708 (N_38708,N_36497,N_36502);
or U38709 (N_38709,N_37198,N_37232);
nand U38710 (N_38710,N_35396,N_35631);
or U38711 (N_38711,N_35273,N_35155);
nand U38712 (N_38712,N_35183,N_35526);
nand U38713 (N_38713,N_36658,N_36577);
or U38714 (N_38714,N_35056,N_37297);
or U38715 (N_38715,N_35034,N_36735);
and U38716 (N_38716,N_37401,N_35194);
or U38717 (N_38717,N_36382,N_36659);
xnor U38718 (N_38718,N_35411,N_37430);
nor U38719 (N_38719,N_36097,N_36166);
or U38720 (N_38720,N_35944,N_36322);
nor U38721 (N_38721,N_36232,N_36128);
and U38722 (N_38722,N_35139,N_36374);
and U38723 (N_38723,N_35108,N_35929);
nand U38724 (N_38724,N_35749,N_36810);
nand U38725 (N_38725,N_37026,N_35160);
and U38726 (N_38726,N_37002,N_37177);
nand U38727 (N_38727,N_35266,N_35824);
xor U38728 (N_38728,N_35666,N_36449);
and U38729 (N_38729,N_35554,N_36682);
and U38730 (N_38730,N_35119,N_35415);
nor U38731 (N_38731,N_37451,N_36456);
nor U38732 (N_38732,N_36962,N_37155);
xnor U38733 (N_38733,N_36035,N_35002);
nand U38734 (N_38734,N_37455,N_37010);
nand U38735 (N_38735,N_36065,N_37303);
or U38736 (N_38736,N_35197,N_35813);
nor U38737 (N_38737,N_35172,N_35680);
xor U38738 (N_38738,N_35544,N_36053);
and U38739 (N_38739,N_35784,N_36510);
xor U38740 (N_38740,N_35368,N_36161);
and U38741 (N_38741,N_36169,N_35123);
or U38742 (N_38742,N_37227,N_35180);
and U38743 (N_38743,N_35583,N_35278);
nand U38744 (N_38744,N_36262,N_35862);
xnor U38745 (N_38745,N_35482,N_35830);
or U38746 (N_38746,N_37082,N_35874);
nor U38747 (N_38747,N_35408,N_36167);
xnor U38748 (N_38748,N_35369,N_35385);
nand U38749 (N_38749,N_35679,N_36568);
or U38750 (N_38750,N_35201,N_35893);
and U38751 (N_38751,N_36897,N_35633);
and U38752 (N_38752,N_36730,N_36126);
and U38753 (N_38753,N_35159,N_35493);
xnor U38754 (N_38754,N_36997,N_35042);
and U38755 (N_38755,N_36913,N_35189);
or U38756 (N_38756,N_35546,N_36467);
nand U38757 (N_38757,N_35778,N_35985);
xor U38758 (N_38758,N_35333,N_35736);
xnor U38759 (N_38759,N_35300,N_35745);
nor U38760 (N_38760,N_36679,N_37257);
and U38761 (N_38761,N_37351,N_37254);
and U38762 (N_38762,N_36372,N_35267);
nand U38763 (N_38763,N_36409,N_36246);
xor U38764 (N_38764,N_37243,N_35694);
nand U38765 (N_38765,N_36689,N_37003);
nand U38766 (N_38766,N_36140,N_36725);
nand U38767 (N_38767,N_36838,N_36956);
or U38768 (N_38768,N_35423,N_35504);
nor U38769 (N_38769,N_37177,N_36243);
xnor U38770 (N_38770,N_36545,N_36112);
xnor U38771 (N_38771,N_35539,N_35932);
or U38772 (N_38772,N_36257,N_36806);
nor U38773 (N_38773,N_35660,N_36259);
xnor U38774 (N_38774,N_35090,N_37165);
nand U38775 (N_38775,N_36303,N_36038);
nand U38776 (N_38776,N_37107,N_36607);
nor U38777 (N_38777,N_36666,N_36512);
nand U38778 (N_38778,N_37314,N_36832);
xor U38779 (N_38779,N_36447,N_36516);
xor U38780 (N_38780,N_36422,N_36921);
nor U38781 (N_38781,N_36161,N_35728);
xnor U38782 (N_38782,N_35300,N_37118);
nor U38783 (N_38783,N_36838,N_36443);
or U38784 (N_38784,N_36140,N_35810);
nand U38785 (N_38785,N_36553,N_37096);
nor U38786 (N_38786,N_35944,N_37419);
nand U38787 (N_38787,N_36877,N_36830);
nand U38788 (N_38788,N_36709,N_36919);
nand U38789 (N_38789,N_36254,N_35913);
or U38790 (N_38790,N_36137,N_36656);
nor U38791 (N_38791,N_36654,N_37293);
nor U38792 (N_38792,N_36840,N_37021);
xor U38793 (N_38793,N_36802,N_35305);
xnor U38794 (N_38794,N_36493,N_37303);
or U38795 (N_38795,N_36846,N_35547);
or U38796 (N_38796,N_35102,N_36035);
or U38797 (N_38797,N_37166,N_35962);
xnor U38798 (N_38798,N_36620,N_35952);
or U38799 (N_38799,N_36998,N_36815);
xor U38800 (N_38800,N_36785,N_36095);
nor U38801 (N_38801,N_36090,N_36650);
nand U38802 (N_38802,N_36047,N_37097);
xnor U38803 (N_38803,N_36019,N_35894);
or U38804 (N_38804,N_36724,N_37330);
or U38805 (N_38805,N_37087,N_35642);
nor U38806 (N_38806,N_36043,N_36480);
xnor U38807 (N_38807,N_37395,N_36966);
nor U38808 (N_38808,N_36034,N_36742);
xor U38809 (N_38809,N_35415,N_35571);
xnor U38810 (N_38810,N_36860,N_36174);
nand U38811 (N_38811,N_36737,N_35335);
nand U38812 (N_38812,N_36148,N_35491);
and U38813 (N_38813,N_37242,N_37138);
xor U38814 (N_38814,N_36158,N_37274);
or U38815 (N_38815,N_36825,N_36534);
and U38816 (N_38816,N_35998,N_37313);
and U38817 (N_38817,N_35745,N_36441);
and U38818 (N_38818,N_35116,N_36577);
nor U38819 (N_38819,N_36774,N_36343);
or U38820 (N_38820,N_37085,N_36477);
or U38821 (N_38821,N_36514,N_36779);
or U38822 (N_38822,N_35785,N_37198);
nand U38823 (N_38823,N_36748,N_36210);
nand U38824 (N_38824,N_35048,N_35798);
nand U38825 (N_38825,N_36803,N_36375);
or U38826 (N_38826,N_36099,N_37370);
and U38827 (N_38827,N_36624,N_35995);
xor U38828 (N_38828,N_35164,N_36601);
and U38829 (N_38829,N_35796,N_35216);
nand U38830 (N_38830,N_36384,N_37379);
nor U38831 (N_38831,N_35330,N_35558);
nor U38832 (N_38832,N_35354,N_35010);
nand U38833 (N_38833,N_36270,N_36739);
and U38834 (N_38834,N_35830,N_35576);
and U38835 (N_38835,N_37391,N_36276);
xnor U38836 (N_38836,N_36739,N_35338);
nor U38837 (N_38837,N_37018,N_36201);
nor U38838 (N_38838,N_37487,N_36064);
nand U38839 (N_38839,N_36363,N_37421);
nand U38840 (N_38840,N_35364,N_36238);
or U38841 (N_38841,N_37090,N_36067);
xor U38842 (N_38842,N_35703,N_36071);
xnor U38843 (N_38843,N_35959,N_37030);
xor U38844 (N_38844,N_37036,N_36250);
nor U38845 (N_38845,N_35410,N_36432);
nor U38846 (N_38846,N_35150,N_36592);
nand U38847 (N_38847,N_35789,N_36441);
or U38848 (N_38848,N_36894,N_36725);
nor U38849 (N_38849,N_35371,N_35897);
or U38850 (N_38850,N_36784,N_36487);
or U38851 (N_38851,N_37151,N_36871);
nor U38852 (N_38852,N_35018,N_37266);
or U38853 (N_38853,N_36468,N_35629);
xnor U38854 (N_38854,N_36687,N_35186);
nor U38855 (N_38855,N_36402,N_36824);
or U38856 (N_38856,N_36028,N_36274);
nor U38857 (N_38857,N_36215,N_36963);
xor U38858 (N_38858,N_37004,N_35887);
or U38859 (N_38859,N_36865,N_36752);
and U38860 (N_38860,N_36792,N_37229);
nor U38861 (N_38861,N_35214,N_36950);
nor U38862 (N_38862,N_35191,N_35714);
or U38863 (N_38863,N_36725,N_35712);
nor U38864 (N_38864,N_35788,N_35848);
and U38865 (N_38865,N_35524,N_35780);
nor U38866 (N_38866,N_37156,N_35510);
xnor U38867 (N_38867,N_35471,N_36027);
or U38868 (N_38868,N_36033,N_35716);
and U38869 (N_38869,N_36795,N_36501);
and U38870 (N_38870,N_35852,N_36139);
or U38871 (N_38871,N_35630,N_37397);
and U38872 (N_38872,N_36308,N_35442);
xnor U38873 (N_38873,N_36217,N_36816);
and U38874 (N_38874,N_37163,N_36490);
nand U38875 (N_38875,N_36129,N_36204);
or U38876 (N_38876,N_35982,N_36036);
and U38877 (N_38877,N_35414,N_36393);
xor U38878 (N_38878,N_35981,N_35456);
and U38879 (N_38879,N_35491,N_36007);
and U38880 (N_38880,N_35185,N_36140);
and U38881 (N_38881,N_35254,N_35342);
nand U38882 (N_38882,N_35750,N_36490);
nand U38883 (N_38883,N_35616,N_35737);
nand U38884 (N_38884,N_36304,N_35685);
or U38885 (N_38885,N_36478,N_37498);
xor U38886 (N_38886,N_35504,N_35419);
and U38887 (N_38887,N_35516,N_37444);
nand U38888 (N_38888,N_35145,N_36524);
and U38889 (N_38889,N_35325,N_35987);
xor U38890 (N_38890,N_37123,N_35037);
xor U38891 (N_38891,N_35325,N_35135);
nor U38892 (N_38892,N_35218,N_37262);
nor U38893 (N_38893,N_37079,N_37086);
nand U38894 (N_38894,N_36132,N_36948);
nand U38895 (N_38895,N_37128,N_35142);
nand U38896 (N_38896,N_37093,N_36718);
nand U38897 (N_38897,N_35366,N_36895);
or U38898 (N_38898,N_35443,N_36528);
nand U38899 (N_38899,N_36109,N_36869);
xor U38900 (N_38900,N_35758,N_36494);
nor U38901 (N_38901,N_36312,N_35328);
nand U38902 (N_38902,N_35780,N_36367);
or U38903 (N_38903,N_35354,N_36919);
nor U38904 (N_38904,N_35840,N_37067);
or U38905 (N_38905,N_36447,N_35382);
or U38906 (N_38906,N_36578,N_36825);
or U38907 (N_38907,N_35467,N_35434);
nor U38908 (N_38908,N_36461,N_35971);
nor U38909 (N_38909,N_35406,N_36020);
xor U38910 (N_38910,N_35477,N_35353);
nor U38911 (N_38911,N_36726,N_36323);
xnor U38912 (N_38912,N_35993,N_35875);
nand U38913 (N_38913,N_37057,N_36517);
xnor U38914 (N_38914,N_35701,N_37457);
nor U38915 (N_38915,N_35006,N_36309);
nor U38916 (N_38916,N_36536,N_35635);
xnor U38917 (N_38917,N_36888,N_35022);
nand U38918 (N_38918,N_36917,N_36860);
or U38919 (N_38919,N_37430,N_36190);
xor U38920 (N_38920,N_36661,N_35195);
and U38921 (N_38921,N_35324,N_37239);
and U38922 (N_38922,N_35615,N_36903);
nor U38923 (N_38923,N_36070,N_36785);
nand U38924 (N_38924,N_36109,N_36384);
nand U38925 (N_38925,N_35021,N_35396);
nor U38926 (N_38926,N_36485,N_36316);
nand U38927 (N_38927,N_36679,N_35107);
nor U38928 (N_38928,N_35379,N_35794);
or U38929 (N_38929,N_37203,N_37402);
and U38930 (N_38930,N_35709,N_35120);
nor U38931 (N_38931,N_35939,N_35947);
or U38932 (N_38932,N_35209,N_35151);
nor U38933 (N_38933,N_35141,N_37446);
xor U38934 (N_38934,N_35770,N_36703);
xnor U38935 (N_38935,N_35787,N_35135);
nor U38936 (N_38936,N_35923,N_35398);
nand U38937 (N_38937,N_36967,N_36800);
nor U38938 (N_38938,N_35373,N_35055);
nor U38939 (N_38939,N_35380,N_36934);
xor U38940 (N_38940,N_36810,N_36265);
and U38941 (N_38941,N_36103,N_37328);
and U38942 (N_38942,N_35570,N_36054);
or U38943 (N_38943,N_35880,N_35715);
and U38944 (N_38944,N_37425,N_35209);
nor U38945 (N_38945,N_36345,N_36255);
or U38946 (N_38946,N_36912,N_37171);
nand U38947 (N_38947,N_37366,N_37398);
nand U38948 (N_38948,N_35575,N_37442);
and U38949 (N_38949,N_35257,N_35949);
or U38950 (N_38950,N_36167,N_36352);
nor U38951 (N_38951,N_35884,N_35123);
nor U38952 (N_38952,N_37455,N_35816);
xnor U38953 (N_38953,N_36669,N_36123);
nand U38954 (N_38954,N_35277,N_35702);
or U38955 (N_38955,N_37247,N_36399);
and U38956 (N_38956,N_35551,N_36329);
or U38957 (N_38957,N_35988,N_37139);
xnor U38958 (N_38958,N_35912,N_37202);
nand U38959 (N_38959,N_36378,N_35313);
or U38960 (N_38960,N_36038,N_36603);
nand U38961 (N_38961,N_36001,N_35565);
and U38962 (N_38962,N_36858,N_35938);
nand U38963 (N_38963,N_35384,N_35470);
and U38964 (N_38964,N_35997,N_36020);
nor U38965 (N_38965,N_35866,N_37098);
and U38966 (N_38966,N_37421,N_37484);
xor U38967 (N_38967,N_37486,N_36462);
and U38968 (N_38968,N_36191,N_37283);
and U38969 (N_38969,N_35076,N_36071);
xor U38970 (N_38970,N_37038,N_35622);
or U38971 (N_38971,N_36772,N_35495);
xnor U38972 (N_38972,N_35042,N_36756);
and U38973 (N_38973,N_35174,N_35457);
xnor U38974 (N_38974,N_36619,N_37302);
xnor U38975 (N_38975,N_37172,N_36638);
xor U38976 (N_38976,N_35953,N_37169);
nand U38977 (N_38977,N_36406,N_36104);
xnor U38978 (N_38978,N_35554,N_36506);
nor U38979 (N_38979,N_37009,N_36452);
xor U38980 (N_38980,N_35526,N_35696);
nor U38981 (N_38981,N_36615,N_36025);
or U38982 (N_38982,N_37443,N_35249);
and U38983 (N_38983,N_36973,N_36839);
nand U38984 (N_38984,N_35451,N_35863);
nor U38985 (N_38985,N_36169,N_35975);
nor U38986 (N_38986,N_36277,N_35620);
or U38987 (N_38987,N_35787,N_36452);
and U38988 (N_38988,N_36579,N_37466);
nand U38989 (N_38989,N_36508,N_36366);
nand U38990 (N_38990,N_37112,N_36307);
and U38991 (N_38991,N_35951,N_36763);
and U38992 (N_38992,N_37305,N_36504);
nand U38993 (N_38993,N_35330,N_35511);
xnor U38994 (N_38994,N_36890,N_36898);
or U38995 (N_38995,N_35671,N_35745);
or U38996 (N_38996,N_35553,N_35104);
nor U38997 (N_38997,N_35458,N_36844);
and U38998 (N_38998,N_35552,N_36922);
or U38999 (N_38999,N_35790,N_36835);
nand U39000 (N_39000,N_36488,N_36461);
and U39001 (N_39001,N_35431,N_36959);
nand U39002 (N_39002,N_36266,N_36214);
nor U39003 (N_39003,N_36522,N_35833);
nor U39004 (N_39004,N_37474,N_35305);
xor U39005 (N_39005,N_36300,N_36634);
nand U39006 (N_39006,N_35963,N_37127);
or U39007 (N_39007,N_36367,N_35061);
or U39008 (N_39008,N_35871,N_36496);
xor U39009 (N_39009,N_36703,N_36132);
xor U39010 (N_39010,N_36774,N_35557);
nand U39011 (N_39011,N_37369,N_36827);
and U39012 (N_39012,N_37117,N_36009);
nor U39013 (N_39013,N_37273,N_37030);
nand U39014 (N_39014,N_35583,N_36788);
or U39015 (N_39015,N_36763,N_36040);
and U39016 (N_39016,N_37265,N_35109);
xor U39017 (N_39017,N_36068,N_36458);
or U39018 (N_39018,N_35800,N_37000);
or U39019 (N_39019,N_36488,N_35928);
nand U39020 (N_39020,N_35303,N_36921);
xnor U39021 (N_39021,N_35861,N_36868);
xnor U39022 (N_39022,N_36654,N_36623);
nor U39023 (N_39023,N_36570,N_36070);
and U39024 (N_39024,N_36451,N_36584);
nor U39025 (N_39025,N_35539,N_35185);
nand U39026 (N_39026,N_35469,N_36555);
and U39027 (N_39027,N_37199,N_37211);
nand U39028 (N_39028,N_36732,N_37162);
nor U39029 (N_39029,N_36059,N_35764);
or U39030 (N_39030,N_36354,N_36069);
xnor U39031 (N_39031,N_36021,N_36352);
and U39032 (N_39032,N_36576,N_36113);
xor U39033 (N_39033,N_37045,N_35470);
nor U39034 (N_39034,N_35671,N_36542);
xnor U39035 (N_39035,N_36389,N_36906);
xnor U39036 (N_39036,N_37428,N_36078);
nor U39037 (N_39037,N_35572,N_35688);
and U39038 (N_39038,N_37388,N_36561);
nand U39039 (N_39039,N_35615,N_36104);
xnor U39040 (N_39040,N_37049,N_37291);
nor U39041 (N_39041,N_37344,N_36459);
or U39042 (N_39042,N_35735,N_35883);
and U39043 (N_39043,N_35700,N_36221);
xnor U39044 (N_39044,N_37303,N_35603);
nor U39045 (N_39045,N_37411,N_36672);
or U39046 (N_39046,N_35664,N_37409);
and U39047 (N_39047,N_35851,N_36030);
or U39048 (N_39048,N_35519,N_35855);
xor U39049 (N_39049,N_37150,N_36541);
xor U39050 (N_39050,N_36017,N_36695);
and U39051 (N_39051,N_35573,N_36932);
nor U39052 (N_39052,N_37372,N_35736);
nor U39053 (N_39053,N_35818,N_35858);
xnor U39054 (N_39054,N_37106,N_35748);
xor U39055 (N_39055,N_35326,N_36348);
and U39056 (N_39056,N_36545,N_36040);
nor U39057 (N_39057,N_35179,N_35074);
or U39058 (N_39058,N_37320,N_36920);
nand U39059 (N_39059,N_36935,N_36373);
nor U39060 (N_39060,N_37038,N_36062);
nand U39061 (N_39061,N_35073,N_35380);
nand U39062 (N_39062,N_36741,N_35308);
and U39063 (N_39063,N_36931,N_37469);
nand U39064 (N_39064,N_35105,N_35235);
nand U39065 (N_39065,N_36401,N_35640);
nand U39066 (N_39066,N_37256,N_35749);
or U39067 (N_39067,N_36273,N_36044);
nand U39068 (N_39068,N_36459,N_36467);
xor U39069 (N_39069,N_35778,N_35084);
nor U39070 (N_39070,N_36948,N_36088);
nand U39071 (N_39071,N_36194,N_37202);
and U39072 (N_39072,N_36034,N_36555);
nand U39073 (N_39073,N_37006,N_36719);
nand U39074 (N_39074,N_36202,N_35522);
xnor U39075 (N_39075,N_35126,N_35470);
or U39076 (N_39076,N_36989,N_35451);
and U39077 (N_39077,N_36129,N_36201);
xnor U39078 (N_39078,N_36036,N_35851);
or U39079 (N_39079,N_36394,N_36188);
nor U39080 (N_39080,N_36307,N_35093);
nand U39081 (N_39081,N_36696,N_36605);
nand U39082 (N_39082,N_35634,N_35573);
nand U39083 (N_39083,N_35235,N_36127);
and U39084 (N_39084,N_35687,N_36374);
or U39085 (N_39085,N_35239,N_36049);
and U39086 (N_39086,N_35129,N_36376);
nand U39087 (N_39087,N_35631,N_35910);
or U39088 (N_39088,N_36808,N_35660);
and U39089 (N_39089,N_35680,N_35527);
nand U39090 (N_39090,N_36470,N_35122);
xor U39091 (N_39091,N_37021,N_37151);
xor U39092 (N_39092,N_36392,N_35960);
or U39093 (N_39093,N_37038,N_37440);
or U39094 (N_39094,N_36366,N_37189);
or U39095 (N_39095,N_36133,N_36987);
nor U39096 (N_39096,N_36726,N_36626);
nand U39097 (N_39097,N_36701,N_36876);
or U39098 (N_39098,N_35208,N_36589);
nand U39099 (N_39099,N_36823,N_37393);
nor U39100 (N_39100,N_35496,N_36959);
nor U39101 (N_39101,N_37240,N_36083);
nand U39102 (N_39102,N_35666,N_35576);
nand U39103 (N_39103,N_35699,N_36953);
or U39104 (N_39104,N_35047,N_35432);
xor U39105 (N_39105,N_36151,N_35432);
nor U39106 (N_39106,N_35247,N_35659);
and U39107 (N_39107,N_36748,N_36088);
nor U39108 (N_39108,N_36076,N_36024);
nor U39109 (N_39109,N_35222,N_35156);
or U39110 (N_39110,N_37441,N_37049);
or U39111 (N_39111,N_36620,N_35213);
nor U39112 (N_39112,N_35836,N_35384);
or U39113 (N_39113,N_35107,N_35820);
xor U39114 (N_39114,N_35891,N_37470);
or U39115 (N_39115,N_36685,N_36656);
nor U39116 (N_39116,N_35090,N_37370);
or U39117 (N_39117,N_35611,N_37304);
nand U39118 (N_39118,N_35987,N_35252);
nand U39119 (N_39119,N_35739,N_36940);
nor U39120 (N_39120,N_35477,N_35234);
nor U39121 (N_39121,N_35578,N_37456);
xnor U39122 (N_39122,N_36603,N_36396);
and U39123 (N_39123,N_36618,N_36146);
xnor U39124 (N_39124,N_35466,N_35094);
xnor U39125 (N_39125,N_36640,N_35726);
nand U39126 (N_39126,N_36305,N_35250);
and U39127 (N_39127,N_37479,N_35555);
nor U39128 (N_39128,N_37135,N_36729);
xnor U39129 (N_39129,N_35147,N_37233);
nand U39130 (N_39130,N_36950,N_36051);
and U39131 (N_39131,N_36650,N_35100);
nor U39132 (N_39132,N_35938,N_36231);
or U39133 (N_39133,N_37448,N_36226);
xnor U39134 (N_39134,N_36209,N_37034);
nor U39135 (N_39135,N_36574,N_35593);
nand U39136 (N_39136,N_36843,N_36462);
and U39137 (N_39137,N_37234,N_36383);
or U39138 (N_39138,N_36861,N_37041);
nand U39139 (N_39139,N_36926,N_37466);
xor U39140 (N_39140,N_36604,N_35950);
xnor U39141 (N_39141,N_36351,N_37308);
or U39142 (N_39142,N_35331,N_35830);
or U39143 (N_39143,N_35234,N_35213);
nand U39144 (N_39144,N_36167,N_35717);
xnor U39145 (N_39145,N_35260,N_35913);
nor U39146 (N_39146,N_37336,N_35988);
or U39147 (N_39147,N_36625,N_36881);
nand U39148 (N_39148,N_36837,N_35820);
and U39149 (N_39149,N_37032,N_36796);
or U39150 (N_39150,N_36037,N_37002);
or U39151 (N_39151,N_37338,N_36290);
nor U39152 (N_39152,N_35807,N_36884);
nor U39153 (N_39153,N_35562,N_36592);
nand U39154 (N_39154,N_36558,N_37238);
xnor U39155 (N_39155,N_36279,N_35166);
and U39156 (N_39156,N_37206,N_35966);
and U39157 (N_39157,N_36383,N_35013);
nor U39158 (N_39158,N_35638,N_36626);
xor U39159 (N_39159,N_37226,N_37315);
xnor U39160 (N_39160,N_37011,N_37092);
nand U39161 (N_39161,N_35011,N_36015);
and U39162 (N_39162,N_35989,N_35477);
nand U39163 (N_39163,N_35468,N_35494);
nor U39164 (N_39164,N_37130,N_37253);
xor U39165 (N_39165,N_36772,N_35106);
nand U39166 (N_39166,N_36700,N_36877);
nor U39167 (N_39167,N_37073,N_35756);
or U39168 (N_39168,N_36386,N_35270);
nor U39169 (N_39169,N_35420,N_37213);
and U39170 (N_39170,N_37346,N_35814);
and U39171 (N_39171,N_37287,N_35010);
nor U39172 (N_39172,N_35523,N_35391);
nand U39173 (N_39173,N_36447,N_36285);
nor U39174 (N_39174,N_36046,N_36105);
xnor U39175 (N_39175,N_35810,N_35850);
nand U39176 (N_39176,N_36903,N_35835);
nand U39177 (N_39177,N_35148,N_37327);
nand U39178 (N_39178,N_36364,N_37358);
or U39179 (N_39179,N_36506,N_35090);
xnor U39180 (N_39180,N_35835,N_36266);
and U39181 (N_39181,N_36921,N_36472);
and U39182 (N_39182,N_35169,N_35061);
or U39183 (N_39183,N_37337,N_36323);
nand U39184 (N_39184,N_35631,N_36075);
nand U39185 (N_39185,N_36428,N_37199);
or U39186 (N_39186,N_36327,N_35702);
nand U39187 (N_39187,N_36177,N_36995);
xor U39188 (N_39188,N_35732,N_36927);
nand U39189 (N_39189,N_37030,N_35015);
nor U39190 (N_39190,N_35725,N_35705);
xnor U39191 (N_39191,N_36398,N_36671);
nor U39192 (N_39192,N_37340,N_37376);
nor U39193 (N_39193,N_36662,N_35030);
nor U39194 (N_39194,N_35829,N_36928);
nor U39195 (N_39195,N_35327,N_36251);
and U39196 (N_39196,N_37423,N_35223);
nor U39197 (N_39197,N_35197,N_36644);
nand U39198 (N_39198,N_37356,N_36080);
or U39199 (N_39199,N_36100,N_36261);
xor U39200 (N_39200,N_35893,N_35623);
or U39201 (N_39201,N_37453,N_35126);
or U39202 (N_39202,N_35835,N_35028);
and U39203 (N_39203,N_36334,N_36716);
or U39204 (N_39204,N_37246,N_36335);
nor U39205 (N_39205,N_35174,N_36591);
xor U39206 (N_39206,N_35974,N_36622);
nor U39207 (N_39207,N_37030,N_36773);
or U39208 (N_39208,N_35397,N_36944);
or U39209 (N_39209,N_35335,N_36150);
and U39210 (N_39210,N_35450,N_37286);
and U39211 (N_39211,N_36179,N_36776);
and U39212 (N_39212,N_37490,N_35796);
and U39213 (N_39213,N_35271,N_35196);
nand U39214 (N_39214,N_36701,N_35935);
or U39215 (N_39215,N_35472,N_37389);
or U39216 (N_39216,N_35091,N_37224);
nand U39217 (N_39217,N_36212,N_36951);
and U39218 (N_39218,N_36896,N_35483);
and U39219 (N_39219,N_36154,N_35935);
nand U39220 (N_39220,N_37096,N_35843);
xnor U39221 (N_39221,N_36176,N_36114);
nand U39222 (N_39222,N_36192,N_36265);
nor U39223 (N_39223,N_35752,N_35404);
xnor U39224 (N_39224,N_35922,N_36514);
xnor U39225 (N_39225,N_35258,N_35555);
nand U39226 (N_39226,N_36845,N_35727);
nor U39227 (N_39227,N_37472,N_37320);
or U39228 (N_39228,N_35394,N_36466);
or U39229 (N_39229,N_37355,N_35158);
and U39230 (N_39230,N_36206,N_36811);
and U39231 (N_39231,N_36547,N_37092);
or U39232 (N_39232,N_35875,N_35408);
nand U39233 (N_39233,N_36405,N_35843);
nand U39234 (N_39234,N_35687,N_35807);
xor U39235 (N_39235,N_35176,N_36322);
xnor U39236 (N_39236,N_35730,N_35849);
nand U39237 (N_39237,N_35143,N_37167);
and U39238 (N_39238,N_36184,N_36910);
xor U39239 (N_39239,N_36526,N_37194);
nor U39240 (N_39240,N_35525,N_35326);
or U39241 (N_39241,N_36143,N_35083);
nand U39242 (N_39242,N_35612,N_35816);
or U39243 (N_39243,N_36730,N_35283);
xor U39244 (N_39244,N_37432,N_35591);
nor U39245 (N_39245,N_35013,N_36798);
nand U39246 (N_39246,N_37345,N_35452);
xor U39247 (N_39247,N_36631,N_35254);
nand U39248 (N_39248,N_36834,N_36217);
or U39249 (N_39249,N_37032,N_37474);
nand U39250 (N_39250,N_37139,N_35611);
or U39251 (N_39251,N_35649,N_35224);
or U39252 (N_39252,N_35022,N_36687);
or U39253 (N_39253,N_37251,N_35912);
nor U39254 (N_39254,N_35559,N_37088);
or U39255 (N_39255,N_35764,N_37310);
nor U39256 (N_39256,N_35309,N_36655);
or U39257 (N_39257,N_35800,N_37416);
and U39258 (N_39258,N_35879,N_36920);
or U39259 (N_39259,N_36012,N_36610);
nor U39260 (N_39260,N_35542,N_37031);
or U39261 (N_39261,N_35053,N_36044);
xor U39262 (N_39262,N_36676,N_35327);
xnor U39263 (N_39263,N_35958,N_36599);
nand U39264 (N_39264,N_35617,N_35975);
xor U39265 (N_39265,N_37478,N_35834);
nand U39266 (N_39266,N_36589,N_36149);
and U39267 (N_39267,N_35789,N_35019);
nor U39268 (N_39268,N_36023,N_36571);
and U39269 (N_39269,N_35219,N_35716);
nor U39270 (N_39270,N_36614,N_35524);
and U39271 (N_39271,N_35619,N_36910);
or U39272 (N_39272,N_36926,N_35004);
nand U39273 (N_39273,N_37447,N_36961);
nand U39274 (N_39274,N_36222,N_36196);
xnor U39275 (N_39275,N_37268,N_35725);
xnor U39276 (N_39276,N_35218,N_35320);
nand U39277 (N_39277,N_35060,N_36245);
nand U39278 (N_39278,N_35234,N_35873);
nor U39279 (N_39279,N_35641,N_36429);
nor U39280 (N_39280,N_36978,N_35146);
and U39281 (N_39281,N_36784,N_37095);
nor U39282 (N_39282,N_37393,N_35209);
or U39283 (N_39283,N_36756,N_37136);
and U39284 (N_39284,N_35192,N_35847);
xnor U39285 (N_39285,N_35973,N_35544);
nor U39286 (N_39286,N_35478,N_36400);
or U39287 (N_39287,N_36509,N_37137);
or U39288 (N_39288,N_36664,N_35436);
nand U39289 (N_39289,N_35785,N_35633);
xnor U39290 (N_39290,N_35335,N_36173);
nor U39291 (N_39291,N_36529,N_36456);
nor U39292 (N_39292,N_36562,N_35762);
or U39293 (N_39293,N_37341,N_37497);
nor U39294 (N_39294,N_36265,N_36250);
nor U39295 (N_39295,N_36068,N_36461);
nand U39296 (N_39296,N_37175,N_37319);
and U39297 (N_39297,N_35597,N_36130);
or U39298 (N_39298,N_35380,N_36222);
nor U39299 (N_39299,N_35348,N_36763);
nand U39300 (N_39300,N_36661,N_35865);
or U39301 (N_39301,N_35012,N_37407);
and U39302 (N_39302,N_36850,N_36544);
nor U39303 (N_39303,N_35908,N_35889);
and U39304 (N_39304,N_37434,N_36734);
or U39305 (N_39305,N_36569,N_37391);
or U39306 (N_39306,N_37394,N_35051);
and U39307 (N_39307,N_36333,N_35058);
nor U39308 (N_39308,N_35384,N_37462);
and U39309 (N_39309,N_36429,N_36596);
nand U39310 (N_39310,N_36718,N_36402);
xor U39311 (N_39311,N_37002,N_36704);
or U39312 (N_39312,N_36076,N_37168);
xnor U39313 (N_39313,N_36892,N_35081);
or U39314 (N_39314,N_35522,N_36939);
xnor U39315 (N_39315,N_35345,N_35441);
xnor U39316 (N_39316,N_35771,N_35830);
xor U39317 (N_39317,N_35198,N_35795);
xnor U39318 (N_39318,N_35476,N_35901);
xor U39319 (N_39319,N_36857,N_35013);
nand U39320 (N_39320,N_36346,N_35698);
nor U39321 (N_39321,N_35748,N_36317);
nand U39322 (N_39322,N_37082,N_36452);
and U39323 (N_39323,N_35862,N_36749);
and U39324 (N_39324,N_35356,N_36144);
and U39325 (N_39325,N_36278,N_36910);
and U39326 (N_39326,N_37212,N_35001);
or U39327 (N_39327,N_35008,N_35931);
or U39328 (N_39328,N_35453,N_35414);
and U39329 (N_39329,N_35920,N_36864);
nand U39330 (N_39330,N_35214,N_35439);
xor U39331 (N_39331,N_35415,N_35872);
nor U39332 (N_39332,N_37367,N_35496);
or U39333 (N_39333,N_35914,N_37048);
nand U39334 (N_39334,N_35904,N_36487);
nor U39335 (N_39335,N_35273,N_36489);
nand U39336 (N_39336,N_37265,N_36085);
nand U39337 (N_39337,N_35066,N_36408);
nand U39338 (N_39338,N_35499,N_37424);
and U39339 (N_39339,N_36248,N_35344);
nor U39340 (N_39340,N_35551,N_36041);
nand U39341 (N_39341,N_36424,N_36756);
or U39342 (N_39342,N_37397,N_35092);
xor U39343 (N_39343,N_35618,N_37214);
xor U39344 (N_39344,N_36099,N_35654);
or U39345 (N_39345,N_35438,N_35580);
and U39346 (N_39346,N_35813,N_36531);
xor U39347 (N_39347,N_36031,N_36473);
xor U39348 (N_39348,N_35060,N_36074);
nand U39349 (N_39349,N_36153,N_37254);
nand U39350 (N_39350,N_36541,N_35389);
or U39351 (N_39351,N_35295,N_37479);
nor U39352 (N_39352,N_37304,N_36315);
nor U39353 (N_39353,N_36875,N_36395);
nand U39354 (N_39354,N_35875,N_37435);
nand U39355 (N_39355,N_35626,N_36801);
nand U39356 (N_39356,N_37356,N_37428);
xnor U39357 (N_39357,N_35292,N_35821);
nand U39358 (N_39358,N_35241,N_37074);
nand U39359 (N_39359,N_36674,N_36561);
nand U39360 (N_39360,N_36088,N_36619);
nand U39361 (N_39361,N_35950,N_37423);
and U39362 (N_39362,N_35494,N_36766);
nor U39363 (N_39363,N_35450,N_35667);
nor U39364 (N_39364,N_36233,N_35849);
or U39365 (N_39365,N_35047,N_35857);
and U39366 (N_39366,N_36469,N_35634);
and U39367 (N_39367,N_35833,N_37236);
and U39368 (N_39368,N_37339,N_37286);
nand U39369 (N_39369,N_37244,N_35899);
nor U39370 (N_39370,N_37212,N_35641);
and U39371 (N_39371,N_36622,N_36767);
or U39372 (N_39372,N_37373,N_36118);
and U39373 (N_39373,N_37179,N_37370);
xnor U39374 (N_39374,N_35826,N_35925);
or U39375 (N_39375,N_35857,N_37182);
or U39376 (N_39376,N_35205,N_35061);
nor U39377 (N_39377,N_36491,N_35420);
nand U39378 (N_39378,N_36247,N_36040);
or U39379 (N_39379,N_36845,N_35564);
or U39380 (N_39380,N_35200,N_35165);
xnor U39381 (N_39381,N_36690,N_35394);
and U39382 (N_39382,N_36220,N_35247);
and U39383 (N_39383,N_36025,N_36369);
xnor U39384 (N_39384,N_36078,N_35413);
and U39385 (N_39385,N_35865,N_35082);
nor U39386 (N_39386,N_37473,N_35884);
or U39387 (N_39387,N_35184,N_36336);
or U39388 (N_39388,N_36077,N_37344);
or U39389 (N_39389,N_37023,N_37011);
and U39390 (N_39390,N_36610,N_36565);
or U39391 (N_39391,N_35775,N_36796);
nor U39392 (N_39392,N_37462,N_36287);
or U39393 (N_39393,N_35537,N_36168);
nand U39394 (N_39394,N_37361,N_37051);
and U39395 (N_39395,N_36466,N_35763);
and U39396 (N_39396,N_36191,N_36367);
and U39397 (N_39397,N_37324,N_35716);
and U39398 (N_39398,N_36654,N_36847);
nand U39399 (N_39399,N_35769,N_36966);
nand U39400 (N_39400,N_36980,N_35815);
nand U39401 (N_39401,N_37247,N_35304);
and U39402 (N_39402,N_36830,N_36815);
or U39403 (N_39403,N_35381,N_35208);
and U39404 (N_39404,N_37112,N_35393);
or U39405 (N_39405,N_35238,N_37090);
nor U39406 (N_39406,N_35409,N_37220);
or U39407 (N_39407,N_37312,N_36037);
nor U39408 (N_39408,N_36392,N_35481);
and U39409 (N_39409,N_35862,N_36359);
xnor U39410 (N_39410,N_36373,N_35716);
xor U39411 (N_39411,N_35625,N_36481);
xnor U39412 (N_39412,N_35575,N_36724);
or U39413 (N_39413,N_36613,N_35408);
or U39414 (N_39414,N_35611,N_36148);
nor U39415 (N_39415,N_37230,N_36013);
xor U39416 (N_39416,N_35657,N_37096);
or U39417 (N_39417,N_37374,N_35583);
nor U39418 (N_39418,N_36060,N_35817);
or U39419 (N_39419,N_35866,N_36612);
xnor U39420 (N_39420,N_37001,N_35033);
and U39421 (N_39421,N_35699,N_35463);
xor U39422 (N_39422,N_37340,N_35045);
and U39423 (N_39423,N_35705,N_36033);
or U39424 (N_39424,N_36522,N_37399);
nor U39425 (N_39425,N_37182,N_36702);
and U39426 (N_39426,N_35145,N_35055);
xor U39427 (N_39427,N_36671,N_35592);
and U39428 (N_39428,N_35258,N_36690);
nor U39429 (N_39429,N_37366,N_35632);
xnor U39430 (N_39430,N_37131,N_37211);
nor U39431 (N_39431,N_35404,N_35430);
or U39432 (N_39432,N_35753,N_37326);
nor U39433 (N_39433,N_35987,N_35106);
nand U39434 (N_39434,N_36553,N_37148);
and U39435 (N_39435,N_35949,N_35259);
and U39436 (N_39436,N_36199,N_36701);
nand U39437 (N_39437,N_35017,N_37216);
or U39438 (N_39438,N_36098,N_35673);
xnor U39439 (N_39439,N_35408,N_36937);
and U39440 (N_39440,N_37451,N_36999);
or U39441 (N_39441,N_35552,N_36989);
xnor U39442 (N_39442,N_36218,N_35359);
and U39443 (N_39443,N_37330,N_36767);
nor U39444 (N_39444,N_37260,N_35578);
nor U39445 (N_39445,N_35000,N_37139);
nand U39446 (N_39446,N_37089,N_37231);
nor U39447 (N_39447,N_37226,N_35457);
nor U39448 (N_39448,N_37409,N_35116);
and U39449 (N_39449,N_35282,N_35745);
xor U39450 (N_39450,N_37145,N_35761);
or U39451 (N_39451,N_35325,N_36438);
or U39452 (N_39452,N_36649,N_37259);
xnor U39453 (N_39453,N_35097,N_35465);
xnor U39454 (N_39454,N_36282,N_37429);
nand U39455 (N_39455,N_37291,N_35779);
and U39456 (N_39456,N_37256,N_35497);
xnor U39457 (N_39457,N_36735,N_35885);
or U39458 (N_39458,N_36668,N_35265);
nor U39459 (N_39459,N_35620,N_35995);
xnor U39460 (N_39460,N_36026,N_37255);
xnor U39461 (N_39461,N_35069,N_36224);
xor U39462 (N_39462,N_37039,N_37143);
and U39463 (N_39463,N_36990,N_36328);
nand U39464 (N_39464,N_35324,N_35145);
nand U39465 (N_39465,N_37280,N_37001);
nor U39466 (N_39466,N_35322,N_36832);
and U39467 (N_39467,N_35958,N_37316);
and U39468 (N_39468,N_37326,N_36261);
nand U39469 (N_39469,N_37152,N_36562);
xor U39470 (N_39470,N_36619,N_35118);
nor U39471 (N_39471,N_36111,N_36267);
and U39472 (N_39472,N_36507,N_36712);
nor U39473 (N_39473,N_36824,N_36653);
nor U39474 (N_39474,N_35276,N_37114);
and U39475 (N_39475,N_37372,N_36573);
nand U39476 (N_39476,N_35057,N_36428);
xor U39477 (N_39477,N_36803,N_35777);
or U39478 (N_39478,N_35074,N_35932);
and U39479 (N_39479,N_36835,N_36245);
nand U39480 (N_39480,N_35150,N_36927);
nand U39481 (N_39481,N_36757,N_36080);
nor U39482 (N_39482,N_37060,N_36050);
nor U39483 (N_39483,N_36818,N_35846);
xor U39484 (N_39484,N_35578,N_36157);
and U39485 (N_39485,N_35279,N_36134);
nand U39486 (N_39486,N_37445,N_37300);
or U39487 (N_39487,N_35864,N_37299);
and U39488 (N_39488,N_35547,N_35491);
xnor U39489 (N_39489,N_35878,N_35946);
xor U39490 (N_39490,N_37214,N_37409);
or U39491 (N_39491,N_37124,N_36030);
or U39492 (N_39492,N_35867,N_35915);
and U39493 (N_39493,N_37392,N_37366);
and U39494 (N_39494,N_37272,N_35298);
xor U39495 (N_39495,N_37187,N_37326);
nand U39496 (N_39496,N_35355,N_37182);
and U39497 (N_39497,N_36900,N_35003);
and U39498 (N_39498,N_35139,N_35603);
xor U39499 (N_39499,N_36654,N_37461);
and U39500 (N_39500,N_36538,N_36724);
or U39501 (N_39501,N_37191,N_37134);
xnor U39502 (N_39502,N_37328,N_36880);
and U39503 (N_39503,N_36163,N_36286);
and U39504 (N_39504,N_36824,N_35371);
nor U39505 (N_39505,N_36506,N_36521);
or U39506 (N_39506,N_37194,N_36765);
xor U39507 (N_39507,N_35499,N_35593);
nand U39508 (N_39508,N_37441,N_35094);
xor U39509 (N_39509,N_36679,N_37156);
nand U39510 (N_39510,N_36868,N_35289);
xor U39511 (N_39511,N_35185,N_35449);
nor U39512 (N_39512,N_35803,N_37474);
or U39513 (N_39513,N_36702,N_35504);
and U39514 (N_39514,N_35693,N_36023);
nor U39515 (N_39515,N_35289,N_37150);
nand U39516 (N_39516,N_35999,N_36877);
and U39517 (N_39517,N_35476,N_36246);
nor U39518 (N_39518,N_37259,N_35177);
xor U39519 (N_39519,N_35622,N_35232);
or U39520 (N_39520,N_35909,N_35208);
xnor U39521 (N_39521,N_35275,N_35736);
and U39522 (N_39522,N_35445,N_35986);
nor U39523 (N_39523,N_36042,N_35760);
or U39524 (N_39524,N_37439,N_36744);
xnor U39525 (N_39525,N_37421,N_36415);
nor U39526 (N_39526,N_36214,N_35677);
or U39527 (N_39527,N_35565,N_36402);
or U39528 (N_39528,N_35172,N_37433);
nor U39529 (N_39529,N_35360,N_36895);
and U39530 (N_39530,N_37451,N_35754);
and U39531 (N_39531,N_35192,N_35077);
xnor U39532 (N_39532,N_35993,N_35193);
nand U39533 (N_39533,N_37253,N_35130);
nor U39534 (N_39534,N_35440,N_36373);
nor U39535 (N_39535,N_37203,N_35576);
nor U39536 (N_39536,N_37250,N_36899);
nor U39537 (N_39537,N_36651,N_36248);
and U39538 (N_39538,N_36356,N_35455);
xor U39539 (N_39539,N_37326,N_35021);
xor U39540 (N_39540,N_35145,N_35744);
or U39541 (N_39541,N_36531,N_36722);
xnor U39542 (N_39542,N_35585,N_37448);
nor U39543 (N_39543,N_35887,N_36635);
xnor U39544 (N_39544,N_36349,N_36378);
nor U39545 (N_39545,N_35082,N_35587);
nor U39546 (N_39546,N_35952,N_37265);
or U39547 (N_39547,N_36046,N_36442);
and U39548 (N_39548,N_35834,N_37463);
and U39549 (N_39549,N_36007,N_36162);
nand U39550 (N_39550,N_36673,N_35491);
nand U39551 (N_39551,N_36046,N_35836);
nand U39552 (N_39552,N_35885,N_36867);
or U39553 (N_39553,N_36444,N_36134);
nand U39554 (N_39554,N_36457,N_35044);
nor U39555 (N_39555,N_36476,N_36284);
and U39556 (N_39556,N_35566,N_36931);
or U39557 (N_39557,N_36780,N_35388);
or U39558 (N_39558,N_36911,N_35984);
nor U39559 (N_39559,N_37256,N_36030);
xor U39560 (N_39560,N_35563,N_36223);
nand U39561 (N_39561,N_36906,N_36253);
xor U39562 (N_39562,N_36207,N_37002);
or U39563 (N_39563,N_36352,N_35804);
xnor U39564 (N_39564,N_36315,N_36370);
nand U39565 (N_39565,N_36593,N_37423);
nand U39566 (N_39566,N_37297,N_35006);
nand U39567 (N_39567,N_35943,N_36980);
or U39568 (N_39568,N_36512,N_35389);
xnor U39569 (N_39569,N_36446,N_35142);
xor U39570 (N_39570,N_35330,N_36582);
or U39571 (N_39571,N_35688,N_35414);
xnor U39572 (N_39572,N_36034,N_35588);
or U39573 (N_39573,N_35677,N_35933);
nor U39574 (N_39574,N_35314,N_37153);
or U39575 (N_39575,N_35373,N_36267);
or U39576 (N_39576,N_35144,N_37248);
or U39577 (N_39577,N_36204,N_36041);
nor U39578 (N_39578,N_36116,N_37355);
or U39579 (N_39579,N_37188,N_35664);
or U39580 (N_39580,N_36683,N_37080);
or U39581 (N_39581,N_35657,N_37035);
and U39582 (N_39582,N_36883,N_36927);
xnor U39583 (N_39583,N_36954,N_36519);
xor U39584 (N_39584,N_35036,N_36572);
or U39585 (N_39585,N_35820,N_35502);
and U39586 (N_39586,N_37355,N_36162);
nor U39587 (N_39587,N_35929,N_36315);
nand U39588 (N_39588,N_37375,N_35055);
nor U39589 (N_39589,N_36058,N_37089);
or U39590 (N_39590,N_37215,N_35590);
nand U39591 (N_39591,N_35246,N_36061);
nor U39592 (N_39592,N_35056,N_37376);
and U39593 (N_39593,N_35730,N_36396);
nor U39594 (N_39594,N_35761,N_37496);
xor U39595 (N_39595,N_35644,N_37346);
nor U39596 (N_39596,N_36444,N_36105);
xor U39597 (N_39597,N_35008,N_37444);
or U39598 (N_39598,N_36827,N_36133);
or U39599 (N_39599,N_36519,N_35043);
nor U39600 (N_39600,N_35772,N_35487);
and U39601 (N_39601,N_36898,N_36595);
xor U39602 (N_39602,N_35697,N_36528);
and U39603 (N_39603,N_35287,N_35460);
xnor U39604 (N_39604,N_35390,N_35708);
and U39605 (N_39605,N_37151,N_37475);
nand U39606 (N_39606,N_37474,N_36732);
and U39607 (N_39607,N_36104,N_35650);
xnor U39608 (N_39608,N_35478,N_35560);
and U39609 (N_39609,N_36218,N_36738);
and U39610 (N_39610,N_36414,N_37473);
or U39611 (N_39611,N_37171,N_35166);
or U39612 (N_39612,N_36796,N_36412);
nor U39613 (N_39613,N_36791,N_35063);
xor U39614 (N_39614,N_37427,N_36916);
nor U39615 (N_39615,N_37183,N_35316);
and U39616 (N_39616,N_36284,N_36718);
nor U39617 (N_39617,N_35248,N_36175);
xnor U39618 (N_39618,N_36573,N_35541);
nand U39619 (N_39619,N_37265,N_36402);
or U39620 (N_39620,N_35854,N_37055);
xor U39621 (N_39621,N_36342,N_35546);
and U39622 (N_39622,N_37044,N_37496);
nor U39623 (N_39623,N_37498,N_37309);
or U39624 (N_39624,N_36556,N_37309);
and U39625 (N_39625,N_37042,N_35711);
or U39626 (N_39626,N_35148,N_37485);
nand U39627 (N_39627,N_35170,N_37447);
nor U39628 (N_39628,N_35351,N_36135);
nand U39629 (N_39629,N_37058,N_37200);
and U39630 (N_39630,N_35070,N_35442);
nor U39631 (N_39631,N_36041,N_35324);
and U39632 (N_39632,N_35412,N_35672);
nor U39633 (N_39633,N_36896,N_35355);
nand U39634 (N_39634,N_36928,N_36124);
or U39635 (N_39635,N_36417,N_37058);
xnor U39636 (N_39636,N_36405,N_37008);
and U39637 (N_39637,N_35498,N_35250);
nand U39638 (N_39638,N_37099,N_36269);
or U39639 (N_39639,N_37205,N_35642);
nand U39640 (N_39640,N_36618,N_37265);
or U39641 (N_39641,N_36889,N_36853);
xor U39642 (N_39642,N_36014,N_35001);
and U39643 (N_39643,N_36722,N_37207);
nand U39644 (N_39644,N_36387,N_37025);
nand U39645 (N_39645,N_35885,N_36153);
nor U39646 (N_39646,N_37346,N_36736);
nand U39647 (N_39647,N_35364,N_36182);
and U39648 (N_39648,N_35420,N_36329);
or U39649 (N_39649,N_36557,N_36343);
and U39650 (N_39650,N_36249,N_36239);
nor U39651 (N_39651,N_35062,N_36353);
nor U39652 (N_39652,N_35593,N_35649);
or U39653 (N_39653,N_35461,N_36269);
nand U39654 (N_39654,N_36140,N_35209);
or U39655 (N_39655,N_35886,N_37049);
and U39656 (N_39656,N_35053,N_35395);
xor U39657 (N_39657,N_37323,N_36497);
or U39658 (N_39658,N_37327,N_35510);
or U39659 (N_39659,N_36585,N_35077);
nor U39660 (N_39660,N_35631,N_35680);
and U39661 (N_39661,N_35909,N_35698);
nand U39662 (N_39662,N_37348,N_35103);
nand U39663 (N_39663,N_36224,N_35318);
and U39664 (N_39664,N_37354,N_37142);
and U39665 (N_39665,N_36997,N_35856);
xor U39666 (N_39666,N_36448,N_36951);
xnor U39667 (N_39667,N_35449,N_37036);
or U39668 (N_39668,N_35079,N_36943);
nand U39669 (N_39669,N_36409,N_36543);
and U39670 (N_39670,N_36430,N_36521);
nand U39671 (N_39671,N_37158,N_36544);
nor U39672 (N_39672,N_36026,N_35240);
nand U39673 (N_39673,N_36031,N_36054);
or U39674 (N_39674,N_37238,N_35508);
nand U39675 (N_39675,N_36640,N_36544);
and U39676 (N_39676,N_36559,N_36259);
or U39677 (N_39677,N_36440,N_35922);
xor U39678 (N_39678,N_35365,N_36277);
nand U39679 (N_39679,N_36888,N_35850);
nor U39680 (N_39680,N_36510,N_36799);
or U39681 (N_39681,N_37422,N_36987);
xnor U39682 (N_39682,N_36990,N_36358);
xnor U39683 (N_39683,N_35786,N_37345);
nand U39684 (N_39684,N_36461,N_36958);
nand U39685 (N_39685,N_37320,N_35045);
nor U39686 (N_39686,N_35515,N_35897);
nor U39687 (N_39687,N_35039,N_36080);
nand U39688 (N_39688,N_36323,N_35449);
xor U39689 (N_39689,N_35596,N_35167);
and U39690 (N_39690,N_35932,N_35838);
xor U39691 (N_39691,N_37132,N_36261);
or U39692 (N_39692,N_35154,N_37119);
nand U39693 (N_39693,N_35183,N_35959);
xor U39694 (N_39694,N_37119,N_35799);
nand U39695 (N_39695,N_35354,N_35462);
xor U39696 (N_39696,N_37077,N_36016);
and U39697 (N_39697,N_35784,N_37058);
xor U39698 (N_39698,N_35708,N_35589);
or U39699 (N_39699,N_37263,N_36192);
xnor U39700 (N_39700,N_35253,N_36342);
nor U39701 (N_39701,N_36654,N_37382);
nor U39702 (N_39702,N_35249,N_35860);
nor U39703 (N_39703,N_35681,N_35234);
nor U39704 (N_39704,N_36277,N_35593);
nand U39705 (N_39705,N_36233,N_37317);
and U39706 (N_39706,N_35431,N_36438);
and U39707 (N_39707,N_35112,N_36121);
and U39708 (N_39708,N_35197,N_35710);
xor U39709 (N_39709,N_35361,N_36122);
and U39710 (N_39710,N_36072,N_35907);
xnor U39711 (N_39711,N_35422,N_36480);
or U39712 (N_39712,N_36323,N_35368);
or U39713 (N_39713,N_36888,N_35432);
nand U39714 (N_39714,N_35861,N_36552);
and U39715 (N_39715,N_35428,N_36531);
and U39716 (N_39716,N_35336,N_36207);
nor U39717 (N_39717,N_35104,N_36906);
or U39718 (N_39718,N_35089,N_36105);
and U39719 (N_39719,N_35099,N_35708);
and U39720 (N_39720,N_37070,N_35041);
and U39721 (N_39721,N_35624,N_36068);
nor U39722 (N_39722,N_36439,N_37061);
nor U39723 (N_39723,N_36447,N_36425);
and U39724 (N_39724,N_35318,N_37472);
nor U39725 (N_39725,N_36612,N_37173);
xor U39726 (N_39726,N_35869,N_37251);
nor U39727 (N_39727,N_36963,N_36510);
nand U39728 (N_39728,N_36866,N_36734);
nor U39729 (N_39729,N_35311,N_35528);
and U39730 (N_39730,N_36053,N_35516);
or U39731 (N_39731,N_36659,N_37024);
nand U39732 (N_39732,N_35178,N_36366);
or U39733 (N_39733,N_36663,N_36080);
nand U39734 (N_39734,N_35986,N_36492);
nor U39735 (N_39735,N_36168,N_36016);
or U39736 (N_39736,N_35687,N_35204);
nand U39737 (N_39737,N_35085,N_36048);
nor U39738 (N_39738,N_35622,N_35549);
nor U39739 (N_39739,N_35378,N_37431);
nor U39740 (N_39740,N_37430,N_36133);
nand U39741 (N_39741,N_35980,N_35667);
nor U39742 (N_39742,N_35391,N_36082);
or U39743 (N_39743,N_36858,N_35710);
xor U39744 (N_39744,N_35079,N_37175);
or U39745 (N_39745,N_36707,N_36038);
and U39746 (N_39746,N_36884,N_35018);
or U39747 (N_39747,N_37130,N_36981);
and U39748 (N_39748,N_36779,N_37359);
nor U39749 (N_39749,N_36273,N_35705);
nor U39750 (N_39750,N_36308,N_35635);
nand U39751 (N_39751,N_35519,N_36254);
or U39752 (N_39752,N_35588,N_35137);
or U39753 (N_39753,N_36049,N_36603);
nand U39754 (N_39754,N_37488,N_36626);
xor U39755 (N_39755,N_35033,N_36497);
nand U39756 (N_39756,N_36883,N_35959);
xnor U39757 (N_39757,N_35166,N_35842);
xor U39758 (N_39758,N_35866,N_36136);
and U39759 (N_39759,N_36434,N_36823);
nor U39760 (N_39760,N_35298,N_36875);
or U39761 (N_39761,N_36253,N_36285);
nand U39762 (N_39762,N_36776,N_35243);
nor U39763 (N_39763,N_37097,N_36916);
nand U39764 (N_39764,N_36178,N_35953);
or U39765 (N_39765,N_35684,N_36400);
and U39766 (N_39766,N_35216,N_36446);
nor U39767 (N_39767,N_35640,N_35598);
nor U39768 (N_39768,N_35983,N_36396);
nor U39769 (N_39769,N_36701,N_36089);
nor U39770 (N_39770,N_36913,N_35222);
xnor U39771 (N_39771,N_36795,N_35123);
and U39772 (N_39772,N_36890,N_35717);
or U39773 (N_39773,N_35312,N_36779);
or U39774 (N_39774,N_37411,N_36269);
xor U39775 (N_39775,N_35505,N_35223);
nand U39776 (N_39776,N_37126,N_36586);
xnor U39777 (N_39777,N_36864,N_35206);
nand U39778 (N_39778,N_35852,N_35699);
nor U39779 (N_39779,N_37288,N_35335);
nand U39780 (N_39780,N_37298,N_36161);
nor U39781 (N_39781,N_35635,N_35197);
and U39782 (N_39782,N_35707,N_35954);
nand U39783 (N_39783,N_35506,N_36344);
and U39784 (N_39784,N_36758,N_35587);
and U39785 (N_39785,N_35086,N_36217);
nor U39786 (N_39786,N_35803,N_36539);
nor U39787 (N_39787,N_37416,N_35328);
or U39788 (N_39788,N_35021,N_37195);
nand U39789 (N_39789,N_37466,N_36750);
nor U39790 (N_39790,N_36960,N_36142);
nand U39791 (N_39791,N_36610,N_36507);
xnor U39792 (N_39792,N_35922,N_37092);
or U39793 (N_39793,N_35892,N_35281);
and U39794 (N_39794,N_37201,N_37473);
and U39795 (N_39795,N_37185,N_35941);
and U39796 (N_39796,N_37127,N_36583);
nor U39797 (N_39797,N_36385,N_37375);
nand U39798 (N_39798,N_36647,N_36855);
or U39799 (N_39799,N_36188,N_35904);
and U39800 (N_39800,N_35012,N_35480);
or U39801 (N_39801,N_36437,N_37431);
nor U39802 (N_39802,N_35877,N_35376);
and U39803 (N_39803,N_35235,N_35518);
nor U39804 (N_39804,N_36217,N_36015);
or U39805 (N_39805,N_35338,N_36334);
nor U39806 (N_39806,N_36095,N_35057);
and U39807 (N_39807,N_37241,N_35520);
or U39808 (N_39808,N_37254,N_35950);
nand U39809 (N_39809,N_36896,N_35334);
nand U39810 (N_39810,N_35669,N_36091);
nor U39811 (N_39811,N_35385,N_36658);
xnor U39812 (N_39812,N_35179,N_37129);
and U39813 (N_39813,N_37285,N_36244);
and U39814 (N_39814,N_36995,N_36853);
nand U39815 (N_39815,N_35919,N_35413);
xnor U39816 (N_39816,N_36931,N_35532);
and U39817 (N_39817,N_35606,N_36522);
xnor U39818 (N_39818,N_35055,N_36070);
nor U39819 (N_39819,N_37277,N_37140);
nor U39820 (N_39820,N_35437,N_35392);
and U39821 (N_39821,N_37295,N_36000);
nor U39822 (N_39822,N_35457,N_37241);
nand U39823 (N_39823,N_36410,N_37168);
and U39824 (N_39824,N_36109,N_35898);
xor U39825 (N_39825,N_37269,N_35762);
xnor U39826 (N_39826,N_37158,N_35534);
or U39827 (N_39827,N_35539,N_37069);
and U39828 (N_39828,N_36610,N_35064);
nand U39829 (N_39829,N_36693,N_36305);
nor U39830 (N_39830,N_35796,N_36667);
or U39831 (N_39831,N_35002,N_36687);
nand U39832 (N_39832,N_36461,N_36664);
nand U39833 (N_39833,N_36863,N_36709);
or U39834 (N_39834,N_36579,N_35826);
nor U39835 (N_39835,N_36137,N_35302);
nand U39836 (N_39836,N_36915,N_36247);
nor U39837 (N_39837,N_36484,N_35125);
xor U39838 (N_39838,N_35467,N_36368);
or U39839 (N_39839,N_36604,N_36408);
nand U39840 (N_39840,N_36299,N_35837);
nor U39841 (N_39841,N_36778,N_36512);
nand U39842 (N_39842,N_35272,N_35373);
nor U39843 (N_39843,N_36801,N_37163);
nand U39844 (N_39844,N_35760,N_36544);
nor U39845 (N_39845,N_35845,N_35252);
nand U39846 (N_39846,N_35476,N_36366);
or U39847 (N_39847,N_37063,N_36345);
or U39848 (N_39848,N_36073,N_35716);
nor U39849 (N_39849,N_35580,N_37147);
nand U39850 (N_39850,N_36099,N_36862);
nor U39851 (N_39851,N_35458,N_37470);
and U39852 (N_39852,N_36890,N_35294);
nor U39853 (N_39853,N_36060,N_35028);
nand U39854 (N_39854,N_36845,N_35803);
or U39855 (N_39855,N_36380,N_35727);
nand U39856 (N_39856,N_37313,N_36415);
nand U39857 (N_39857,N_37374,N_36071);
and U39858 (N_39858,N_35144,N_35767);
xor U39859 (N_39859,N_35658,N_37134);
and U39860 (N_39860,N_36253,N_36149);
nor U39861 (N_39861,N_35199,N_36992);
xor U39862 (N_39862,N_36834,N_36040);
or U39863 (N_39863,N_35990,N_37168);
and U39864 (N_39864,N_37351,N_36850);
nand U39865 (N_39865,N_36235,N_35247);
or U39866 (N_39866,N_36875,N_35261);
or U39867 (N_39867,N_36533,N_36110);
nor U39868 (N_39868,N_36262,N_35857);
xnor U39869 (N_39869,N_37278,N_36160);
nor U39870 (N_39870,N_35267,N_37347);
nor U39871 (N_39871,N_36056,N_36597);
nand U39872 (N_39872,N_36121,N_36449);
or U39873 (N_39873,N_36100,N_37016);
or U39874 (N_39874,N_37415,N_35062);
nor U39875 (N_39875,N_36517,N_36838);
xor U39876 (N_39876,N_36131,N_37006);
xor U39877 (N_39877,N_35482,N_36566);
xnor U39878 (N_39878,N_35203,N_35519);
nor U39879 (N_39879,N_35651,N_36710);
nand U39880 (N_39880,N_35419,N_37286);
or U39881 (N_39881,N_35868,N_36892);
and U39882 (N_39882,N_37315,N_35227);
or U39883 (N_39883,N_35767,N_37134);
nand U39884 (N_39884,N_35582,N_37029);
or U39885 (N_39885,N_36981,N_36267);
and U39886 (N_39886,N_36712,N_36730);
or U39887 (N_39887,N_35164,N_35409);
or U39888 (N_39888,N_35148,N_36950);
or U39889 (N_39889,N_35914,N_36763);
xor U39890 (N_39890,N_35979,N_35225);
nand U39891 (N_39891,N_35256,N_36179);
and U39892 (N_39892,N_36475,N_35795);
nand U39893 (N_39893,N_35483,N_35923);
nor U39894 (N_39894,N_35915,N_37012);
nand U39895 (N_39895,N_36723,N_36768);
or U39896 (N_39896,N_36338,N_35284);
or U39897 (N_39897,N_35368,N_35017);
nand U39898 (N_39898,N_37013,N_36376);
xor U39899 (N_39899,N_35904,N_36709);
nand U39900 (N_39900,N_35850,N_35096);
xnor U39901 (N_39901,N_37203,N_35173);
or U39902 (N_39902,N_36104,N_36658);
nand U39903 (N_39903,N_35302,N_37408);
or U39904 (N_39904,N_36396,N_36781);
nand U39905 (N_39905,N_36964,N_35398);
or U39906 (N_39906,N_36407,N_37180);
and U39907 (N_39907,N_37242,N_36304);
nor U39908 (N_39908,N_35274,N_37289);
nor U39909 (N_39909,N_36438,N_35511);
or U39910 (N_39910,N_35676,N_35036);
or U39911 (N_39911,N_35470,N_35507);
xor U39912 (N_39912,N_35054,N_35978);
or U39913 (N_39913,N_36904,N_37473);
xnor U39914 (N_39914,N_35147,N_37498);
nand U39915 (N_39915,N_35829,N_36549);
xor U39916 (N_39916,N_37141,N_35717);
nand U39917 (N_39917,N_35814,N_36265);
and U39918 (N_39918,N_36171,N_36967);
xor U39919 (N_39919,N_36306,N_36026);
nor U39920 (N_39920,N_37319,N_37300);
or U39921 (N_39921,N_36736,N_36777);
nand U39922 (N_39922,N_36015,N_35783);
and U39923 (N_39923,N_36621,N_35158);
and U39924 (N_39924,N_35438,N_37390);
or U39925 (N_39925,N_36876,N_36809);
and U39926 (N_39926,N_35823,N_36210);
nand U39927 (N_39927,N_37228,N_35697);
nand U39928 (N_39928,N_35454,N_36377);
or U39929 (N_39929,N_37266,N_35177);
xnor U39930 (N_39930,N_35159,N_36016);
nor U39931 (N_39931,N_36008,N_35067);
and U39932 (N_39932,N_35478,N_36610);
or U39933 (N_39933,N_35031,N_35790);
nand U39934 (N_39934,N_37407,N_35106);
or U39935 (N_39935,N_35324,N_35389);
or U39936 (N_39936,N_35893,N_36220);
nand U39937 (N_39937,N_36485,N_35433);
and U39938 (N_39938,N_35370,N_35013);
nand U39939 (N_39939,N_35295,N_37364);
nor U39940 (N_39940,N_36450,N_37294);
xor U39941 (N_39941,N_36416,N_36532);
nand U39942 (N_39942,N_35405,N_35275);
or U39943 (N_39943,N_36191,N_35451);
nor U39944 (N_39944,N_36980,N_35300);
nand U39945 (N_39945,N_36625,N_37456);
and U39946 (N_39946,N_37133,N_36647);
xnor U39947 (N_39947,N_36985,N_37127);
xor U39948 (N_39948,N_35976,N_35431);
and U39949 (N_39949,N_37146,N_35770);
and U39950 (N_39950,N_35864,N_36663);
nor U39951 (N_39951,N_35400,N_36910);
and U39952 (N_39952,N_35876,N_35253);
nor U39953 (N_39953,N_36737,N_35228);
xnor U39954 (N_39954,N_35041,N_35634);
and U39955 (N_39955,N_37197,N_35526);
nand U39956 (N_39956,N_36119,N_35677);
or U39957 (N_39957,N_36998,N_36592);
nor U39958 (N_39958,N_36537,N_35893);
or U39959 (N_39959,N_36151,N_35813);
xor U39960 (N_39960,N_35945,N_37195);
nor U39961 (N_39961,N_35192,N_35383);
or U39962 (N_39962,N_35883,N_35376);
nor U39963 (N_39963,N_35380,N_35207);
or U39964 (N_39964,N_35501,N_35925);
nand U39965 (N_39965,N_37148,N_36138);
xor U39966 (N_39966,N_36881,N_36970);
or U39967 (N_39967,N_35155,N_36234);
xnor U39968 (N_39968,N_36800,N_35040);
xor U39969 (N_39969,N_35170,N_36147);
xor U39970 (N_39970,N_37035,N_35414);
xor U39971 (N_39971,N_35084,N_36690);
or U39972 (N_39972,N_36650,N_37048);
nor U39973 (N_39973,N_35868,N_37480);
and U39974 (N_39974,N_35293,N_37118);
or U39975 (N_39975,N_36720,N_35434);
nand U39976 (N_39976,N_35723,N_35458);
xnor U39977 (N_39977,N_37235,N_37421);
nor U39978 (N_39978,N_36652,N_36471);
and U39979 (N_39979,N_37124,N_36941);
nor U39980 (N_39980,N_37226,N_36707);
xnor U39981 (N_39981,N_35467,N_35103);
nor U39982 (N_39982,N_37238,N_36712);
or U39983 (N_39983,N_35721,N_37125);
xnor U39984 (N_39984,N_36908,N_35248);
xnor U39985 (N_39985,N_37044,N_35544);
and U39986 (N_39986,N_36707,N_36407);
nor U39987 (N_39987,N_35305,N_37399);
and U39988 (N_39988,N_36817,N_35756);
nor U39989 (N_39989,N_35946,N_36547);
and U39990 (N_39990,N_35515,N_35417);
xnor U39991 (N_39991,N_36427,N_35785);
nand U39992 (N_39992,N_36936,N_36508);
and U39993 (N_39993,N_35227,N_35967);
xor U39994 (N_39994,N_37192,N_35454);
xnor U39995 (N_39995,N_36463,N_36397);
xnor U39996 (N_39996,N_36582,N_35556);
and U39997 (N_39997,N_36611,N_35234);
or U39998 (N_39998,N_35930,N_36309);
nand U39999 (N_39999,N_36766,N_35686);
nor U40000 (N_40000,N_38408,N_38865);
xnor U40001 (N_40001,N_38213,N_39324);
and U40002 (N_40002,N_38382,N_37800);
and U40003 (N_40003,N_38592,N_39712);
nand U40004 (N_40004,N_38914,N_38240);
xnor U40005 (N_40005,N_38902,N_37845);
nor U40006 (N_40006,N_37639,N_39305);
or U40007 (N_40007,N_37673,N_38156);
or U40008 (N_40008,N_37681,N_37608);
or U40009 (N_40009,N_38053,N_38999);
xor U40010 (N_40010,N_38314,N_39379);
nor U40011 (N_40011,N_38151,N_37878);
nand U40012 (N_40012,N_38602,N_39396);
and U40013 (N_40013,N_38386,N_38623);
and U40014 (N_40014,N_38438,N_38540);
or U40015 (N_40015,N_37983,N_38395);
and U40016 (N_40016,N_39401,N_38858);
xor U40017 (N_40017,N_37719,N_38588);
and U40018 (N_40018,N_39467,N_37892);
xnor U40019 (N_40019,N_38308,N_38742);
nand U40020 (N_40020,N_38167,N_39373);
and U40021 (N_40021,N_37834,N_37505);
and U40022 (N_40022,N_39386,N_39322);
and U40023 (N_40023,N_39795,N_39351);
nand U40024 (N_40024,N_37678,N_38854);
xnor U40025 (N_40025,N_39514,N_39819);
and U40026 (N_40026,N_38568,N_39357);
xnor U40027 (N_40027,N_39275,N_38991);
and U40028 (N_40028,N_38951,N_39016);
or U40029 (N_40029,N_38823,N_37944);
or U40030 (N_40030,N_39135,N_37709);
nand U40031 (N_40031,N_38440,N_38948);
nand U40032 (N_40032,N_39944,N_38917);
or U40033 (N_40033,N_39958,N_38507);
nand U40034 (N_40034,N_39165,N_38866);
xor U40035 (N_40035,N_38725,N_38277);
nor U40036 (N_40036,N_38757,N_39519);
nand U40037 (N_40037,N_39445,N_38882);
nand U40038 (N_40038,N_39708,N_38223);
nand U40039 (N_40039,N_37605,N_39633);
xnor U40040 (N_40040,N_37975,N_39179);
nand U40041 (N_40041,N_37818,N_38543);
nand U40042 (N_40042,N_39659,N_38590);
and U40043 (N_40043,N_38895,N_39508);
nor U40044 (N_40044,N_39882,N_38424);
xor U40045 (N_40045,N_39950,N_38913);
nand U40046 (N_40046,N_39364,N_38700);
nor U40047 (N_40047,N_38899,N_39991);
or U40048 (N_40048,N_39718,N_39833);
xnor U40049 (N_40049,N_37597,N_38388);
or U40050 (N_40050,N_38585,N_39033);
nor U40051 (N_40051,N_37692,N_38406);
nand U40052 (N_40052,N_38580,N_37882);
xor U40053 (N_40053,N_39417,N_37787);
and U40054 (N_40054,N_37573,N_38934);
xor U40055 (N_40055,N_37943,N_39735);
nand U40056 (N_40056,N_39737,N_38530);
or U40057 (N_40057,N_38557,N_38840);
and U40058 (N_40058,N_39687,N_39136);
nor U40059 (N_40059,N_38443,N_39640);
nor U40060 (N_40060,N_37508,N_37902);
xnor U40061 (N_40061,N_37657,N_39931);
and U40062 (N_40062,N_37691,N_38337);
nand U40063 (N_40063,N_37520,N_38176);
or U40064 (N_40064,N_38367,N_39554);
xnor U40065 (N_40065,N_39465,N_39487);
nor U40066 (N_40066,N_39030,N_38643);
nor U40067 (N_40067,N_37895,N_39667);
nand U40068 (N_40068,N_37519,N_37796);
and U40069 (N_40069,N_39437,N_39488);
nor U40070 (N_40070,N_38068,N_39891);
xnor U40071 (N_40071,N_38679,N_38041);
or U40072 (N_40072,N_38433,N_38920);
xor U40073 (N_40073,N_37526,N_38509);
and U40074 (N_40074,N_39630,N_39060);
nand U40075 (N_40075,N_38606,N_38409);
or U40076 (N_40076,N_39404,N_39564);
nand U40077 (N_40077,N_38446,N_39252);
or U40078 (N_40078,N_37633,N_39051);
or U40079 (N_40079,N_39068,N_38564);
and U40080 (N_40080,N_37851,N_38555);
xor U40081 (N_40081,N_37821,N_38935);
nor U40082 (N_40082,N_38239,N_39538);
and U40083 (N_40083,N_39064,N_39578);
nand U40084 (N_40084,N_39828,N_39800);
nor U40085 (N_40085,N_37516,N_39682);
or U40086 (N_40086,N_39518,N_39907);
nand U40087 (N_40087,N_38937,N_38259);
nor U40088 (N_40088,N_38230,N_38879);
nor U40089 (N_40089,N_38181,N_37789);
and U40090 (N_40090,N_37718,N_39365);
xor U40091 (N_40091,N_38010,N_39694);
xor U40092 (N_40092,N_39367,N_38856);
or U40093 (N_40093,N_39425,N_37893);
nand U40094 (N_40094,N_39428,N_39658);
and U40095 (N_40095,N_39317,N_38921);
or U40096 (N_40096,N_38488,N_38610);
and U40097 (N_40097,N_38779,N_38207);
or U40098 (N_40098,N_38510,N_39112);
and U40099 (N_40099,N_39778,N_39957);
or U40100 (N_40100,N_38476,N_39414);
xnor U40101 (N_40101,N_38248,N_39599);
nor U40102 (N_40102,N_37914,N_37799);
xnor U40103 (N_40103,N_37768,N_39710);
and U40104 (N_40104,N_38430,N_38561);
nor U40105 (N_40105,N_39638,N_39174);
nand U40106 (N_40106,N_38302,N_38467);
nor U40107 (N_40107,N_38579,N_39119);
and U40108 (N_40108,N_39966,N_38023);
nand U40109 (N_40109,N_39495,N_38817);
or U40110 (N_40110,N_39688,N_39183);
or U40111 (N_40111,N_37534,N_37643);
nor U40112 (N_40112,N_39701,N_39143);
xnor U40113 (N_40113,N_39159,N_38925);
nor U40114 (N_40114,N_38855,N_38318);
nand U40115 (N_40115,N_38361,N_39360);
and U40116 (N_40116,N_39486,N_37765);
nand U40117 (N_40117,N_38738,N_38296);
or U40118 (N_40118,N_37886,N_39949);
nand U40119 (N_40119,N_39935,N_38799);
or U40120 (N_40120,N_37953,N_39766);
and U40121 (N_40121,N_38743,N_39539);
and U40122 (N_40122,N_37791,N_37770);
nor U40123 (N_40123,N_38164,N_38997);
and U40124 (N_40124,N_39526,N_37815);
or U40125 (N_40125,N_38607,N_39319);
and U40126 (N_40126,N_39607,N_39644);
or U40127 (N_40127,N_39408,N_39499);
nor U40128 (N_40128,N_39559,N_39310);
or U40129 (N_40129,N_38881,N_39483);
nand U40130 (N_40130,N_38576,N_38560);
or U40131 (N_40131,N_39240,N_38050);
nand U40132 (N_40132,N_39296,N_39382);
and U40133 (N_40133,N_39468,N_38215);
nor U40134 (N_40134,N_38208,N_38319);
xor U40135 (N_40135,N_38864,N_37781);
nand U40136 (N_40136,N_39103,N_38535);
xor U40137 (N_40137,N_39995,N_38279);
xor U40138 (N_40138,N_39190,N_38158);
nand U40139 (N_40139,N_37969,N_39042);
nand U40140 (N_40140,N_37972,N_39561);
and U40141 (N_40141,N_38235,N_39723);
nor U40142 (N_40142,N_39522,N_38619);
nor U40143 (N_40143,N_39491,N_39091);
nand U40144 (N_40144,N_39510,N_39978);
xnor U40145 (N_40145,N_37826,N_38227);
and U40146 (N_40146,N_39615,N_39237);
or U40147 (N_40147,N_39147,N_38170);
and U40148 (N_40148,N_39243,N_38403);
nor U40149 (N_40149,N_39482,N_39655);
and U40150 (N_40150,N_39082,N_38187);
xor U40151 (N_40151,N_39732,N_38718);
or U40152 (N_40152,N_38454,N_38286);
nand U40153 (N_40153,N_39196,N_38995);
or U40154 (N_40154,N_37712,N_39044);
nand U40155 (N_40155,N_39129,N_39527);
xnor U40156 (N_40156,N_38791,N_38265);
xnor U40157 (N_40157,N_38055,N_37501);
or U40158 (N_40158,N_39820,N_38062);
xor U40159 (N_40159,N_37568,N_37683);
or U40160 (N_40160,N_37711,N_39493);
and U40161 (N_40161,N_39881,N_37662);
nor U40162 (N_40162,N_39444,N_39844);
xor U40163 (N_40163,N_38599,N_39755);
nor U40164 (N_40164,N_39283,N_37959);
nand U40165 (N_40165,N_39650,N_37872);
xnor U40166 (N_40166,N_38830,N_37612);
or U40167 (N_40167,N_39320,N_37804);
nor U40168 (N_40168,N_38275,N_39794);
and U40169 (N_40169,N_39123,N_38922);
nor U40170 (N_40170,N_38089,N_38548);
nand U40171 (N_40171,N_37729,N_39853);
or U40172 (N_40172,N_39854,N_39062);
nor U40173 (N_40173,N_37701,N_38106);
xnor U40174 (N_40174,N_38168,N_39864);
nand U40175 (N_40175,N_37772,N_39228);
nor U40176 (N_40176,N_39739,N_38013);
xnor U40177 (N_40177,N_37962,N_38414);
xnor U40178 (N_40178,N_37951,N_39779);
and U40179 (N_40179,N_37922,N_38480);
nor U40180 (N_40180,N_37580,N_39328);
or U40181 (N_40181,N_38005,N_37952);
xnor U40182 (N_40182,N_38877,N_38150);
and U40183 (N_40183,N_39805,N_39069);
nand U40184 (N_40184,N_39842,N_38975);
xnor U40185 (N_40185,N_39341,N_39241);
nand U40186 (N_40186,N_38002,N_38003);
nand U40187 (N_40187,N_37535,N_39646);
xor U40188 (N_40188,N_37682,N_39504);
nor U40189 (N_40189,N_38924,N_39156);
nor U40190 (N_40190,N_39740,N_38056);
and U40191 (N_40191,N_38836,N_37559);
xnor U40192 (N_40192,N_39450,N_38824);
or U40193 (N_40193,N_39680,N_38832);
and U40194 (N_40194,N_39497,N_39407);
or U40195 (N_40195,N_39734,N_37672);
nand U40196 (N_40196,N_37599,N_37801);
and U40197 (N_40197,N_38985,N_38411);
xnor U40198 (N_40198,N_39756,N_39541);
xor U40199 (N_40199,N_39372,N_39690);
xor U40200 (N_40200,N_37561,N_38959);
xor U40201 (N_40201,N_39791,N_38664);
xnor U40202 (N_40202,N_38040,N_38853);
xnor U40203 (N_40203,N_38165,N_39822);
nand U40204 (N_40204,N_38380,N_38456);
xnor U40205 (N_40205,N_38701,N_38867);
or U40206 (N_40206,N_39329,N_38415);
or U40207 (N_40207,N_39188,N_38805);
or U40208 (N_40208,N_39919,N_38465);
nand U40209 (N_40209,N_39339,N_38061);
xor U40210 (N_40210,N_39413,N_39035);
or U40211 (N_40211,N_39577,N_37925);
xor U40212 (N_40212,N_37758,N_39323);
nand U40213 (N_40213,N_37993,N_38511);
nor U40214 (N_40214,N_37610,N_39337);
nand U40215 (N_40215,N_38578,N_37745);
xor U40216 (N_40216,N_37759,N_39567);
and U40217 (N_40217,N_37536,N_39021);
nor U40218 (N_40218,N_39751,N_37531);
and U40219 (N_40219,N_38255,N_39804);
or U40220 (N_40220,N_39203,N_38519);
or U40221 (N_40221,N_39420,N_38283);
nor U40222 (N_40222,N_38980,N_38027);
and U40223 (N_40223,N_39045,N_39879);
nand U40224 (N_40224,N_39975,N_37858);
and U40225 (N_40225,N_39273,N_37644);
xor U40226 (N_40226,N_38608,N_39993);
nand U40227 (N_40227,N_38596,N_38137);
nor U40228 (N_40228,N_37660,N_39586);
nand U40229 (N_40229,N_38039,N_39370);
xnor U40230 (N_40230,N_38604,N_38807);
nor U40231 (N_40231,N_38004,N_38886);
or U40232 (N_40232,N_38368,N_38897);
nand U40233 (N_40233,N_39847,N_38225);
or U40234 (N_40234,N_39209,N_39169);
nor U40235 (N_40235,N_37553,N_37912);
xnor U40236 (N_40236,N_39485,N_39478);
or U40237 (N_40237,N_39392,N_38401);
xnor U40238 (N_40238,N_37564,N_37947);
and U40239 (N_40239,N_39581,N_37847);
or U40240 (N_40240,N_38735,N_38697);
and U40241 (N_40241,N_37806,N_37589);
xor U40242 (N_40242,N_38307,N_37549);
or U40243 (N_40243,N_38378,N_39344);
xor U40244 (N_40244,N_39703,N_38007);
and U40245 (N_40245,N_37514,N_39972);
xor U40246 (N_40246,N_38503,N_38715);
nand U40247 (N_40247,N_38675,N_38315);
nor U40248 (N_40248,N_39525,N_37769);
nor U40249 (N_40249,N_38801,N_39609);
xnor U40250 (N_40250,N_39571,N_38976);
and U40251 (N_40251,N_39848,N_39587);
nand U40252 (N_40252,N_38819,N_39124);
xor U40253 (N_40253,N_39551,N_39956);
nand U40254 (N_40254,N_39385,N_37511);
xnor U40255 (N_40255,N_38605,N_39532);
or U40256 (N_40256,N_38138,N_37704);
nand U40257 (N_40257,N_37970,N_38891);
nand U40258 (N_40258,N_37849,N_38998);
and U40259 (N_40259,N_39231,N_39639);
nand U40260 (N_40260,N_39632,N_37773);
nor U40261 (N_40261,N_38345,N_38583);
and U40262 (N_40262,N_38067,N_39851);
xnor U40263 (N_40263,N_38110,N_39890);
nand U40264 (N_40264,N_39276,N_39137);
or U40265 (N_40265,N_38703,N_38927);
and U40266 (N_40266,N_38827,N_38375);
and U40267 (N_40267,N_38441,N_38483);
or U40268 (N_40268,N_37824,N_38086);
or U40269 (N_40269,N_39164,N_37618);
nand U40270 (N_40270,N_38698,N_39888);
and U40271 (N_40271,N_37632,N_38571);
or U40272 (N_40272,N_37786,N_38473);
nor U40273 (N_40273,N_38276,N_38767);
or U40274 (N_40274,N_38667,N_37737);
and U40275 (N_40275,N_39874,N_39318);
or U40276 (N_40276,N_38019,N_38774);
and U40277 (N_40277,N_39388,N_38224);
and U40278 (N_40278,N_39185,N_38874);
nor U40279 (N_40279,N_37687,N_39764);
nand U40280 (N_40280,N_38332,N_39007);
and U40281 (N_40281,N_37888,N_39783);
or U40282 (N_40282,N_38575,N_39754);
nor U40283 (N_40283,N_39004,N_39942);
or U40284 (N_40284,N_38828,N_38662);
xor U40285 (N_40285,N_39566,N_39178);
or U40286 (N_40286,N_39789,N_38246);
and U40287 (N_40287,N_38525,N_38748);
or U40288 (N_40288,N_39937,N_37569);
xnor U40289 (N_40289,N_37503,N_37584);
nor U40290 (N_40290,N_37819,N_37583);
nor U40291 (N_40291,N_38582,N_38981);
and U40292 (N_40292,N_37811,N_39479);
or U40293 (N_40293,N_39358,N_38155);
nor U40294 (N_40294,N_37909,N_39434);
xnor U40295 (N_40295,N_38966,N_39979);
and U40296 (N_40296,N_38945,N_38033);
and U40297 (N_40297,N_38124,N_39221);
xnor U40298 (N_40298,N_38074,N_38898);
and U40299 (N_40299,N_39162,N_37680);
nand U40300 (N_40300,N_39161,N_39948);
or U40301 (N_40301,N_39049,N_38638);
nor U40302 (N_40302,N_39788,N_37901);
and U40303 (N_40303,N_38105,N_38944);
and U40304 (N_40304,N_38732,N_37864);
and U40305 (N_40305,N_39821,N_37546);
nand U40306 (N_40306,N_38731,N_39114);
xnor U40307 (N_40307,N_39065,N_37714);
xor U40308 (N_40308,N_38189,N_37986);
and U40309 (N_40309,N_37782,N_39301);
and U40310 (N_40310,N_39748,N_37848);
nor U40311 (N_40311,N_38344,N_38264);
and U40312 (N_40312,N_38673,N_38694);
or U40313 (N_40313,N_39025,N_39459);
and U40314 (N_40314,N_38090,N_38025);
nand U40315 (N_40315,N_38835,N_38531);
nor U40316 (N_40316,N_39175,N_38093);
xnor U40317 (N_40317,N_38706,N_37860);
nor U40318 (N_40318,N_38437,N_38135);
and U40319 (N_40319,N_39464,N_39715);
and U40320 (N_40320,N_38299,N_39523);
xor U40321 (N_40321,N_38569,N_39052);
or U40322 (N_40322,N_39120,N_39335);
xnor U40323 (N_40323,N_38195,N_39006);
nand U40324 (N_40324,N_39731,N_39573);
xnor U40325 (N_40325,N_39439,N_37996);
nand U40326 (N_40326,N_39053,N_39440);
or U40327 (N_40327,N_39387,N_38237);
or U40328 (N_40328,N_39097,N_39997);
xor U40329 (N_40329,N_39697,N_38736);
and U40330 (N_40330,N_39102,N_38630);
or U40331 (N_40331,N_39160,N_37948);
xnor U40332 (N_40332,N_39670,N_38071);
nand U40333 (N_40333,N_37507,N_39291);
or U40334 (N_40334,N_37626,N_38120);
and U40335 (N_40335,N_38979,N_38589);
and U40336 (N_40336,N_39889,N_39570);
nor U40337 (N_40337,N_37852,N_39066);
or U40338 (N_40338,N_37794,N_39803);
and U40339 (N_40339,N_38479,N_38085);
or U40340 (N_40340,N_37931,N_37923);
and U40341 (N_40341,N_39969,N_39238);
nand U40342 (N_40342,N_38047,N_38955);
xor U40343 (N_40343,N_38946,N_39782);
or U40344 (N_40344,N_37707,N_39177);
and U40345 (N_40345,N_38633,N_38770);
and U40346 (N_40346,N_37928,N_38097);
or U40347 (N_40347,N_38175,N_39260);
and U40348 (N_40348,N_39503,N_39953);
or U40349 (N_40349,N_37686,N_37844);
nand U40350 (N_40350,N_37788,N_37596);
nand U40351 (N_40351,N_37699,N_37907);
and U40352 (N_40352,N_38804,N_39806);
nand U40353 (N_40353,N_39197,N_38219);
xnor U40354 (N_40354,N_38100,N_39256);
and U40355 (N_40355,N_38676,N_39515);
and U40356 (N_40356,N_37763,N_38313);
nor U40357 (N_40357,N_38044,N_38566);
nand U40358 (N_40358,N_37945,N_39691);
nor U40359 (N_40359,N_39709,N_38983);
or U40360 (N_40360,N_39664,N_37968);
or U40361 (N_40361,N_37631,N_39208);
and U40362 (N_40362,N_38968,N_38193);
xor U40363 (N_40363,N_39597,N_38938);
and U40364 (N_40364,N_39166,N_39880);
nor U40365 (N_40365,N_39032,N_37880);
nor U40366 (N_40366,N_38058,N_38232);
or U40367 (N_40367,N_38852,N_38372);
or U40368 (N_40368,N_39222,N_38421);
xnor U40369 (N_40369,N_39974,N_38896);
nor U40370 (N_40370,N_38764,N_38449);
xnor U40371 (N_40371,N_37883,N_39151);
nand U40372 (N_40372,N_39608,N_37991);
nor U40373 (N_40373,N_38627,N_39116);
or U40374 (N_40374,N_38696,N_37924);
or U40375 (N_40375,N_38123,N_39696);
nor U40376 (N_40376,N_38941,N_39768);
xnor U40377 (N_40377,N_38932,N_39430);
xor U40378 (N_40378,N_38300,N_38108);
nor U40379 (N_40379,N_39282,N_39113);
or U40380 (N_40380,N_39476,N_38661);
nand U40381 (N_40381,N_38690,N_37735);
nor U40382 (N_40382,N_37839,N_38992);
xor U40383 (N_40383,N_39406,N_38659);
xor U40384 (N_40384,N_39543,N_39517);
or U40385 (N_40385,N_38103,N_38876);
and U40386 (N_40386,N_37904,N_37598);
or U40387 (N_40387,N_38140,N_38185);
or U40388 (N_40388,N_39122,N_39770);
nand U40389 (N_40389,N_38842,N_39451);
or U40390 (N_40390,N_38459,N_38741);
or U40391 (N_40391,N_37509,N_37600);
xnor U40392 (N_40392,N_39574,N_39247);
or U40393 (N_40393,N_39153,N_39878);
xor U40394 (N_40394,N_38048,N_38839);
xor U40395 (N_40395,N_38177,N_38052);
xnor U40396 (N_40396,N_39786,N_39433);
nand U40397 (N_40397,N_39355,N_38851);
xor U40398 (N_40398,N_38143,N_39898);
nor U40399 (N_40399,N_38129,N_37675);
and U40400 (N_40400,N_38733,N_39227);
and U40401 (N_40401,N_38258,N_38280);
or U40402 (N_40402,N_39498,N_39870);
and U40403 (N_40403,N_38113,N_39613);
nand U40404 (N_40404,N_38884,N_38015);
xor U40405 (N_40405,N_39552,N_39193);
nand U40406 (N_40406,N_38171,N_38260);
nor U40407 (N_40407,N_37710,N_38445);
and U40408 (N_40408,N_39968,N_37767);
nor U40409 (N_40409,N_39810,N_37679);
or U40410 (N_40410,N_39921,N_38148);
nor U40411 (N_40411,N_38719,N_38420);
nor U40412 (N_40412,N_38594,N_39915);
nor U40413 (N_40413,N_37690,N_38651);
nor U40414 (N_40414,N_39895,N_38848);
xnor U40415 (N_40415,N_39584,N_38844);
and U40416 (N_40416,N_39563,N_38648);
and U40417 (N_40417,N_38760,N_39947);
xnor U40418 (N_40418,N_38758,N_39389);
or U40419 (N_40419,N_38046,N_38098);
nor U40420 (N_40420,N_37930,N_39126);
nor U40421 (N_40421,N_38849,N_37853);
xor U40422 (N_40422,N_39668,N_38190);
xor U40423 (N_40423,N_37656,N_38136);
xor U40424 (N_40424,N_39704,N_39908);
nand U40425 (N_40425,N_38154,N_39824);
and U40426 (N_40426,N_37971,N_39375);
and U40427 (N_40427,N_39366,N_39125);
and U40428 (N_40428,N_38771,N_39206);
nand U40429 (N_40429,N_37578,N_38262);
xnor U40430 (N_40430,N_39652,N_39999);
nand U40431 (N_40431,N_39628,N_38726);
nand U40432 (N_40432,N_38474,N_38036);
nor U40433 (N_40433,N_37581,N_38978);
nor U40434 (N_40434,N_38365,N_38335);
and U40435 (N_40435,N_38458,N_39376);
or U40436 (N_40436,N_37798,N_39941);
xor U40437 (N_40437,N_39651,N_38766);
xnor U40438 (N_40438,N_38699,N_39105);
xor U40439 (N_40439,N_38524,N_37877);
xor U40440 (N_40440,N_39588,N_39077);
and U40441 (N_40441,N_39904,N_38947);
or U40442 (N_40442,N_37870,N_37905);
and U40443 (N_40443,N_37558,N_37539);
and U40444 (N_40444,N_38618,N_38180);
or U40445 (N_40445,N_37997,N_37793);
nor U40446 (N_40446,N_39402,N_39505);
xnor U40447 (N_40447,N_38915,N_37903);
or U40448 (N_40448,N_38523,N_39758);
or U40449 (N_40449,N_38534,N_38763);
xnor U40450 (N_40450,N_39281,N_39471);
and U40451 (N_40451,N_39424,N_39446);
and U40452 (N_40452,N_38567,N_39167);
nand U40453 (N_40453,N_38486,N_39780);
xor U40454 (N_40454,N_38873,N_39549);
xor U40455 (N_40455,N_38965,N_38631);
or U40456 (N_40456,N_39534,N_38722);
and U40457 (N_40457,N_38883,N_38014);
or U40458 (N_40458,N_38723,N_39678);
and U40459 (N_40459,N_38472,N_38006);
xnor U40460 (N_40460,N_38383,N_39677);
and U40461 (N_40461,N_39531,N_39391);
xnor U40462 (N_40462,N_37929,N_39099);
or U40463 (N_40463,N_37621,N_39753);
nand U40464 (N_40464,N_39716,N_38250);
xnor U40465 (N_40465,N_39802,N_39987);
and U40466 (N_40466,N_39168,N_38077);
or U40467 (N_40467,N_39138,N_39757);
nand U40468 (N_40468,N_38778,N_37667);
and U40469 (N_40469,N_38847,N_38145);
and U40470 (N_40470,N_38721,N_39321);
and U40471 (N_40471,N_38954,N_39332);
and U40472 (N_40472,N_39246,N_38655);
nor U40473 (N_40473,N_38029,N_37841);
nor U40474 (N_40474,N_39769,N_38125);
and U40475 (N_40475,N_37960,N_38892);
nand U40476 (N_40476,N_38744,N_39244);
nor U40477 (N_40477,N_38418,N_38179);
or U40478 (N_40478,N_38261,N_39290);
nand U40479 (N_40479,N_38903,N_37795);
nand U40480 (N_40480,N_37627,N_39343);
and U40481 (N_40481,N_38521,N_39614);
xor U40482 (N_40482,N_38172,N_39191);
or U40483 (N_40483,N_38402,N_39015);
nor U40484 (N_40484,N_38485,N_39046);
nor U40485 (N_40485,N_39250,N_38496);
or U40486 (N_40486,N_39259,N_39264);
xor U40487 (N_40487,N_38786,N_39455);
nor U40488 (N_40488,N_37694,N_37830);
or U40489 (N_40489,N_39918,N_38815);
or U40490 (N_40490,N_39520,N_37708);
nand U40491 (N_40491,N_39965,N_38747);
nor U40492 (N_40492,N_37606,N_38427);
nor U40493 (N_40493,N_39832,N_39666);
and U40494 (N_40494,N_37720,N_39325);
xnor U40495 (N_40495,N_38072,N_39249);
xnor U40496 (N_40496,N_38912,N_39954);
xnor U40497 (N_40497,N_39108,N_38812);
xnor U40498 (N_40498,N_37832,N_38829);
nor U40499 (N_40499,N_38196,N_38457);
or U40500 (N_40500,N_37650,N_38413);
or U40501 (N_40501,N_38439,N_38009);
and U40502 (N_40502,N_39906,N_37855);
nand U40503 (N_40503,N_37868,N_37748);
nor U40504 (N_40504,N_38958,N_37994);
nand U40505 (N_40505,N_39580,N_39189);
xor U40506 (N_40506,N_39299,N_38984);
or U40507 (N_40507,N_39187,N_37956);
nand U40508 (N_40508,N_37776,N_38501);
nand U40509 (N_40509,N_38419,N_38628);
xnor U40510 (N_40510,N_38267,N_37829);
nand U40511 (N_40511,N_39925,N_38789);
xor U40512 (N_40512,N_39749,N_37889);
and U40513 (N_40513,N_39058,N_39812);
nand U40514 (N_40514,N_38026,N_37554);
or U40515 (N_40515,N_39378,N_39171);
nand U40516 (N_40516,N_39263,N_39500);
nand U40517 (N_40517,N_38102,N_38359);
or U40518 (N_40518,N_39726,N_38349);
nand U40519 (N_40519,N_39436,N_38652);
or U40520 (N_40520,N_38289,N_38159);
nand U40521 (N_40521,N_37805,N_38964);
nor U40522 (N_40522,N_39985,N_39717);
and U40523 (N_40523,N_37935,N_39901);
or U40524 (N_40524,N_39182,N_38730);
and U40525 (N_40525,N_37676,N_38777);
nand U40526 (N_40526,N_38518,N_39115);
and U40527 (N_40527,N_39265,N_39873);
or U40528 (N_40528,N_38092,N_38448);
and U40529 (N_40529,N_38312,N_37512);
nand U40530 (N_40530,N_38182,N_38814);
nor U40531 (N_40531,N_38245,N_39314);
nand U40532 (N_40532,N_38890,N_39130);
nor U40533 (N_40533,N_39288,N_39825);
and U40534 (N_40534,N_39315,N_38512);
nor U40535 (N_40535,N_39477,N_39826);
and U40536 (N_40536,N_38251,N_37642);
xor U40537 (N_40537,N_37736,N_39683);
and U40538 (N_40538,N_39807,N_38268);
or U40539 (N_40539,N_38134,N_37827);
and U40540 (N_40540,N_38668,N_39040);
xnor U40541 (N_40541,N_39811,N_39635);
or U40542 (N_40542,N_39910,N_38432);
nand U40543 (N_40543,N_37777,N_37881);
nand U40544 (N_40544,N_37571,N_37808);
nor U40545 (N_40545,N_38183,N_39217);
or U40546 (N_40546,N_37835,N_37649);
nand U40547 (N_40547,N_39596,N_37560);
or U40548 (N_40548,N_39435,N_39106);
nand U40549 (N_40549,N_39923,N_38609);
nand U40550 (N_40550,N_38205,N_37529);
nand U40551 (N_40551,N_39371,N_37999);
nand U40552 (N_40552,N_38271,N_39381);
or U40553 (N_40553,N_38504,N_39932);
or U40554 (N_40554,N_39792,N_39695);
or U40555 (N_40555,N_37695,N_39349);
or U40556 (N_40556,N_37728,N_39239);
xnor U40557 (N_40557,N_38869,N_38099);
nor U40558 (N_40558,N_39547,N_38339);
nand U40559 (N_40559,N_38505,N_37607);
nand U40560 (N_40560,N_39516,N_37950);
xnor U40561 (N_40561,N_38933,N_39741);
or U40562 (N_40562,N_38907,N_38537);
nand U40563 (N_40563,N_37664,N_37822);
xor U40564 (N_40564,N_39591,N_38317);
nor U40565 (N_40565,N_38341,N_38775);
nand U40566 (N_40566,N_39837,N_39198);
or U40567 (N_40567,N_38549,N_38773);
or U40568 (N_40568,N_38209,N_39213);
or U40569 (N_40569,N_37937,N_38768);
xnor U40570 (N_40570,N_37920,N_39605);
or U40571 (N_40571,N_37785,N_39180);
nor U40572 (N_40572,N_39509,N_37843);
nor U40573 (N_40573,N_38366,N_39257);
nand U40574 (N_40574,N_39297,N_39867);
xor U40575 (N_40575,N_37521,N_39261);
nand U40576 (N_40576,N_38597,N_39777);
and U40577 (N_40577,N_39730,N_38256);
xnor U40578 (N_40578,N_37563,N_39154);
nor U40579 (N_40579,N_38541,N_38682);
xor U40580 (N_40580,N_37982,N_39951);
nor U40581 (N_40581,N_39070,N_38451);
or U40582 (N_40582,N_39254,N_39063);
or U40583 (N_40583,N_37731,N_38544);
nor U40584 (N_40584,N_39767,N_39393);
and U40585 (N_40585,N_38574,N_39469);
or U40586 (N_40586,N_39347,N_38634);
nor U40587 (N_40587,N_38199,N_37715);
nor U40588 (N_40588,N_39916,N_39745);
xnor U40589 (N_40589,N_39617,N_37661);
or U40590 (N_40590,N_39940,N_37645);
nand U40591 (N_40591,N_39096,N_37622);
xnor U40592 (N_40592,N_39269,N_38516);
nand U40593 (N_40593,N_38547,N_38970);
xor U40594 (N_40594,N_37706,N_37619);
nor U40595 (N_40595,N_38573,N_39462);
nor U40596 (N_40596,N_38042,N_37863);
and U40597 (N_40597,N_38515,N_38893);
xor U40598 (N_40598,N_38384,N_37658);
nor U40599 (N_40599,N_39170,N_39374);
nand U40600 (N_40600,N_39416,N_37575);
nor U40601 (N_40601,N_37916,N_37754);
nor U40602 (N_40602,N_38845,N_38803);
or U40603 (N_40603,N_37502,N_38563);
xor U40604 (N_40604,N_39223,N_39456);
nand U40605 (N_40605,N_38772,N_37638);
nand U40606 (N_40606,N_39251,N_39280);
or U40607 (N_40607,N_38011,N_38243);
and U40608 (N_40608,N_39146,N_39403);
or U40609 (N_40609,N_38214,N_38810);
nor U40610 (N_40610,N_37885,N_39606);
nor U40611 (N_40611,N_39194,N_39286);
nor U40612 (N_40612,N_37544,N_39308);
and U40613 (N_40613,N_37884,N_39234);
or U40614 (N_40614,N_39218,N_38083);
nor U40615 (N_40615,N_37648,N_39742);
nor U40616 (N_40616,N_39302,N_38043);
or U40617 (N_40617,N_39142,N_37774);
xor U40618 (N_40618,N_38115,N_39738);
and U40619 (N_40619,N_38186,N_38529);
xor U40620 (N_40620,N_39913,N_38021);
or U40621 (N_40621,N_37530,N_39797);
xor U40622 (N_40622,N_39988,N_39657);
nor U40623 (N_40623,N_39936,N_37775);
nand U40624 (N_40624,N_38422,N_38233);
nor U40625 (N_40625,N_38257,N_39970);
or U40626 (N_40626,N_39899,N_37703);
nor U40627 (N_40627,N_37913,N_39431);
xor U40628 (N_40628,N_39662,N_38894);
nand U40629 (N_40629,N_38231,N_38707);
xor U40630 (N_40630,N_38202,N_38054);
and U40631 (N_40631,N_38931,N_38127);
xnor U40632 (N_40632,N_39307,N_37674);
nand U40633 (N_40633,N_37854,N_38716);
nand U40634 (N_40634,N_39660,N_38929);
xor U40635 (N_40635,N_37725,N_39986);
xor U40636 (N_40636,N_37857,N_38943);
nand U40637 (N_40637,N_39955,N_37603);
xor U40638 (N_40638,N_38498,N_38740);
or U40639 (N_40639,N_38621,N_39946);
nor U40640 (N_40640,N_38806,N_39029);
nor U40641 (N_40641,N_38989,N_38916);
nand U40642 (N_40642,N_39340,N_39472);
nand U40643 (N_40643,N_37936,N_38550);
nand U40644 (N_40644,N_37752,N_37611);
nand U40645 (N_40645,N_38994,N_38900);
xnor U40646 (N_40646,N_38645,N_39207);
and U40647 (N_40647,N_37570,N_37572);
nor U40648 (N_40648,N_37590,N_39542);
or U40649 (N_40649,N_38570,N_38338);
or U40650 (N_40650,N_39109,N_38163);
nor U40651 (N_40651,N_38669,N_37602);
and U40652 (N_40652,N_38442,N_39279);
and U40653 (N_40653,N_39298,N_39595);
nor U40654 (N_40654,N_39869,N_39248);
and U40655 (N_40655,N_38392,N_39368);
or U40656 (N_40656,N_38666,N_38971);
and U40657 (N_40657,N_38918,N_39815);
nor U40658 (N_40658,N_38252,N_39056);
nor U40659 (N_40659,N_37543,N_39380);
xnor U40660 (N_40660,N_37987,N_37696);
nor U40661 (N_40661,N_37957,N_38565);
xor U40662 (N_40662,N_37540,N_38436);
nor U40663 (N_40663,N_39028,N_38428);
nand U40664 (N_40664,N_38377,N_39557);
or U40665 (N_40665,N_37537,N_37663);
or U40666 (N_40666,N_39176,N_38494);
nand U40667 (N_40667,N_37555,N_39560);
or U40668 (N_40668,N_38051,N_37973);
and U40669 (N_40669,N_39400,N_37734);
xor U40670 (N_40670,N_37523,N_37641);
nor U40671 (N_40671,N_38577,N_37946);
nand U40672 (N_40672,N_38923,N_39054);
nor U40673 (N_40673,N_37942,N_39494);
and U40674 (N_40674,N_39686,N_38360);
and U40675 (N_40675,N_37918,N_37875);
nor U40676 (N_40676,N_39513,N_38389);
and U40677 (N_40677,N_39300,N_38405);
nand U40678 (N_40678,N_39868,N_39155);
or U40679 (N_40679,N_38184,N_38687);
xnor U40680 (N_40680,N_37746,N_37749);
or U40681 (N_40681,N_38974,N_38693);
nand U40682 (N_40682,N_38952,N_37921);
nor U40683 (N_40683,N_38909,N_37616);
and U40684 (N_40684,N_39598,N_37846);
xnor U40685 (N_40685,N_39023,N_39216);
nand U40686 (N_40686,N_39685,N_39507);
nor U40687 (N_40687,N_39134,N_39418);
or U40688 (N_40688,N_38489,N_39994);
and U40689 (N_40689,N_38532,N_38228);
or U40690 (N_40690,N_39866,N_38826);
or U40691 (N_40691,N_38904,N_39480);
nor U40692 (N_40692,N_39841,N_38794);
nand U40693 (N_40693,N_38362,N_39454);
xnor U40694 (N_40694,N_38084,N_39843);
or U40695 (N_40695,N_37528,N_37552);
xnor U40696 (N_40696,N_39857,N_37807);
or U40697 (N_40697,N_37640,N_38713);
or U40698 (N_40698,N_38328,N_38491);
nand U40699 (N_40699,N_37965,N_38091);
xor U40700 (N_40700,N_37577,N_39511);
nor U40701 (N_40701,N_37550,N_39037);
or U40702 (N_40702,N_38453,N_39001);
or U40703 (N_40703,N_38800,N_38455);
or U40704 (N_40704,N_37723,N_38686);
nand U40705 (N_40705,N_37504,N_39359);
nand U40706 (N_40706,N_37614,N_37979);
nor U40707 (N_40707,N_39733,N_38790);
xor U40708 (N_40708,N_39415,N_39293);
or U40709 (N_40709,N_39622,N_38174);
or U40710 (N_40710,N_39002,N_39041);
or U40711 (N_40711,N_39000,N_39038);
or U40712 (N_40712,N_39158,N_39992);
and U40713 (N_40713,N_37792,N_39289);
and U40714 (N_40714,N_38431,N_39012);
nor U40715 (N_40715,N_39647,N_39061);
nor U40716 (N_40716,N_39353,N_38028);
nand U40717 (N_40717,N_38755,N_38087);
nand U40718 (N_40718,N_37634,N_39760);
xor U40719 (N_40719,N_38320,N_38957);
xor U40720 (N_40720,N_39681,N_37601);
or U40721 (N_40721,N_39896,N_39871);
xor U40722 (N_40722,N_39369,N_38132);
and U40723 (N_40723,N_39761,N_39653);
xnor U40724 (N_40724,N_38095,N_37817);
and U40725 (N_40725,N_38689,N_39872);
and U40726 (N_40726,N_37862,N_37859);
or U40727 (N_40727,N_38825,N_39453);
and U40728 (N_40728,N_38354,N_39625);
and U40729 (N_40729,N_38506,N_39752);
nand U40730 (N_40730,N_38254,N_39090);
nand U40731 (N_40731,N_39903,N_38502);
nand U40732 (N_40732,N_39977,N_38121);
and U40733 (N_40733,N_39095,N_38355);
or U40734 (N_40734,N_39423,N_38684);
xor U40735 (N_40735,N_39031,N_39793);
xnor U40736 (N_40736,N_39781,N_37628);
xor U40737 (N_40737,N_37716,N_38562);
and U40738 (N_40738,N_39084,N_39858);
or U40739 (N_40739,N_39914,N_38426);
or U40740 (N_40740,N_38393,N_37820);
or U40741 (N_40741,N_38756,N_39724);
nor U40742 (N_40742,N_37803,N_37582);
or U40743 (N_40743,N_38635,N_38324);
xnor U40744 (N_40744,N_37506,N_37828);
nor U40745 (N_40745,N_38461,N_38220);
nand U40746 (N_40746,N_37867,N_39814);
and U40747 (N_40747,N_37780,N_38769);
xor U40748 (N_40748,N_38032,N_38273);
nor U40749 (N_40749,N_39849,N_38369);
and U40750 (N_40750,N_39980,N_39473);
xor U40751 (N_40751,N_38119,N_39934);
nor U40752 (N_40752,N_38323,N_37685);
xor U40753 (N_40753,N_38200,N_39528);
and U40754 (N_40754,N_38517,N_39714);
xnor U40755 (N_40755,N_39924,N_37964);
nor U40756 (N_40756,N_39665,N_38281);
and U40757 (N_40757,N_38990,N_38330);
and U40758 (N_40758,N_38820,N_39157);
xor U40759 (N_40759,N_37747,N_39863);
or U40760 (N_40760,N_37995,N_37542);
nor U40761 (N_40761,N_39303,N_38963);
nor U40762 (N_40762,N_39771,N_37980);
nand U40763 (N_40763,N_38434,N_39003);
nand U40764 (N_40764,N_38728,N_37966);
nand U40765 (N_40765,N_37739,N_38466);
and U40766 (N_40766,N_37961,N_38834);
xnor U40767 (N_40767,N_39285,N_37992);
or U40768 (N_40768,N_39845,N_38162);
xor U40769 (N_40769,N_39277,N_37814);
nand U40770 (N_40770,N_39558,N_39593);
xor U40771 (N_40771,N_38860,N_37587);
and U40772 (N_40772,N_37566,N_39861);
and U40773 (N_40773,N_37556,N_38301);
or U40774 (N_40774,N_38038,N_39111);
nand U40775 (N_40775,N_37873,N_39850);
nor U40776 (N_40776,N_38452,N_38688);
nand U40777 (N_40777,N_39550,N_38236);
and U40778 (N_40778,N_38288,N_39074);
xnor U40779 (N_40779,N_39117,N_38711);
xnor U40780 (N_40780,N_39700,N_37981);
nand U40781 (N_40781,N_39104,N_39998);
xnor U40782 (N_40782,N_39073,N_39836);
and U40783 (N_40783,N_39211,N_38475);
and U40784 (N_40784,N_37927,N_38987);
xnor U40785 (N_40785,N_37762,N_39312);
nor U40786 (N_40786,N_39173,N_39506);
and U40787 (N_40787,N_38650,N_37698);
nor U40788 (N_40788,N_38065,N_38045);
nand U40789 (N_40789,N_37866,N_39361);
xor U40790 (N_40790,N_37740,N_39594);
and U40791 (N_40791,N_39327,N_38739);
xnor U40792 (N_40792,N_38212,N_39132);
or U40793 (N_40793,N_39398,N_37778);
xnor U40794 (N_40794,N_39059,N_37790);
nor U40795 (N_40795,N_38714,N_38292);
and U40796 (N_40796,N_39929,N_39081);
nor U40797 (N_40797,N_38782,N_39585);
or U40798 (N_40798,N_39967,N_37911);
and U40799 (N_40799,N_39692,N_39075);
and U40800 (N_40800,N_38285,N_38298);
nand U40801 (N_40801,N_39705,N_39399);
nor U40802 (N_40802,N_37545,N_38130);
xor U40803 (N_40803,N_38996,N_38057);
or U40804 (N_40804,N_37551,N_38166);
xor U40805 (N_40805,N_39110,N_38203);
nand U40806 (N_40806,N_38720,N_39088);
and U40807 (N_40807,N_37697,N_39626);
xor U40808 (N_40808,N_39627,N_38637);
or U40809 (N_40809,N_39774,N_39922);
xor U40810 (N_40810,N_39675,N_39618);
nor U40811 (N_40811,N_38928,N_38226);
nand U40812 (N_40812,N_38263,N_38147);
nor U40813 (N_40813,N_38206,N_37717);
nand U40814 (N_40814,N_39540,N_38468);
nor U40815 (N_40815,N_38905,N_38822);
xor U40816 (N_40816,N_39887,N_38674);
nand U40817 (N_40817,N_37688,N_39900);
nor U40818 (N_40818,N_39311,N_38333);
or U40819 (N_40819,N_38704,N_38906);
nand U40820 (N_40820,N_38846,N_38114);
or U40821 (N_40821,N_38327,N_38734);
nand U40822 (N_40822,N_38070,N_38204);
nor U40823 (N_40823,N_38161,N_37812);
or U40824 (N_40824,N_38107,N_39267);
and U40825 (N_40825,N_38234,N_37977);
xor U40826 (N_40826,N_38781,N_38653);
and U40827 (N_40827,N_39927,N_38746);
or U40828 (N_40828,N_38539,N_38216);
and U40829 (N_40829,N_37861,N_38144);
and U40830 (N_40830,N_38930,N_39270);
nor U40831 (N_40831,N_38888,N_39746);
nand U40832 (N_40832,N_38191,N_38069);
and U40833 (N_40833,N_37910,N_38598);
nor U40834 (N_40834,N_38837,N_39020);
xnor U40835 (N_40835,N_37730,N_38001);
or U40836 (N_40836,N_39649,N_39034);
and U40837 (N_40837,N_38871,N_39438);
xor U40838 (N_40838,N_37525,N_37955);
or U40839 (N_40839,N_38526,N_39645);
nand U40840 (N_40840,N_38538,N_39055);
or U40841 (N_40841,N_39024,N_37624);
and U40842 (N_40842,N_38499,N_39195);
nor U40843 (N_40843,N_38500,N_39763);
nor U40844 (N_40844,N_39817,N_39463);
nor U40845 (N_40845,N_38031,N_38911);
and U40846 (N_40846,N_39885,N_39530);
xnor U40847 (N_40847,N_38616,N_37665);
or U40848 (N_40848,N_39233,N_37651);
xnor U40849 (N_40849,N_39306,N_39458);
nand U40850 (N_40850,N_38950,N_39449);
xor U40851 (N_40851,N_38717,N_39048);
and U40852 (N_40852,N_38075,N_38765);
nor U40853 (N_40853,N_37836,N_38647);
nand U40854 (N_40854,N_39629,N_37779);
nand U40855 (N_40855,N_37513,N_37908);
nand U40856 (N_40856,N_39656,N_38595);
or U40857 (N_40857,N_39011,N_39799);
nor U40858 (N_40858,N_39911,N_39546);
and U40859 (N_40859,N_39611,N_39982);
xnor U40860 (N_40860,N_39838,N_39362);
or U40861 (N_40861,N_37900,N_39725);
nand U40862 (N_40862,N_37755,N_39569);
nor U40863 (N_40863,N_39984,N_37684);
xnor U40864 (N_40864,N_38311,N_39669);
and U40865 (N_40865,N_39621,N_38112);
or U40866 (N_40866,N_39535,N_38508);
nor U40867 (N_40867,N_37756,N_39905);
nor U40868 (N_40868,N_38649,N_39253);
nor U40869 (N_40869,N_38484,N_37940);
nand U40870 (N_40870,N_37833,N_37547);
or U40871 (N_40871,N_39834,N_38622);
xnor U40872 (N_40872,N_37988,N_39562);
and U40873 (N_40873,N_38615,N_38859);
or U40874 (N_40874,N_38342,N_39089);
xnor U40875 (N_40875,N_39642,N_37533);
nand U40876 (N_40876,N_39230,N_39076);
nor U40877 (N_40877,N_39582,N_38788);
or U40878 (N_40878,N_38394,N_39713);
nand U40879 (N_40879,N_37974,N_38961);
nand U40880 (N_40880,N_39590,N_37750);
and U40881 (N_40881,N_39294,N_39796);
nor U40882 (N_40882,N_39214,N_38244);
nor U40883 (N_40883,N_39427,N_39390);
xor U40884 (N_40884,N_38910,N_37976);
or U40885 (N_40885,N_38613,N_39926);
xnor U40886 (N_40886,N_38513,N_37637);
xor U40887 (N_40887,N_38270,N_38364);
nor U40888 (N_40888,N_38391,N_37978);
or U40889 (N_40889,N_39501,N_38435);
and U40890 (N_40890,N_39674,N_38076);
xor U40891 (N_40891,N_39461,N_38020);
nand U40892 (N_40892,N_39897,N_38482);
nand U40893 (N_40893,N_38000,N_38982);
nor U40894 (N_40894,N_39938,N_38657);
or U40895 (N_40895,N_38593,N_37934);
nor U40896 (N_40896,N_38064,N_38060);
xor U40897 (N_40897,N_38101,N_38287);
nand U40898 (N_40898,N_39728,N_37594);
and U40899 (N_40899,N_37515,N_39865);
and U40900 (N_40900,N_37856,N_37869);
nor U40901 (N_40901,N_38624,N_39536);
or U40902 (N_40902,N_38663,N_39663);
and U40903 (N_40903,N_38646,N_39579);
or U40904 (N_40904,N_39684,N_38644);
and U40905 (N_40905,N_38536,N_38708);
nand U40906 (N_40906,N_37527,N_38141);
nand U40907 (N_40907,N_37802,N_38880);
nand U40908 (N_40908,N_39600,N_37917);
xor U40909 (N_40909,N_39830,N_37653);
xor U40910 (N_40910,N_39859,N_38821);
xnor U40911 (N_40911,N_39548,N_39971);
and U40912 (N_40912,N_38625,N_39466);
nor U40913 (N_40913,N_38552,N_37896);
and U40914 (N_40914,N_39447,N_39983);
xnor U40915 (N_40915,N_39776,N_38861);
nand U40916 (N_40916,N_38626,N_38811);
xor U40917 (N_40917,N_39457,N_37891);
nand U40918 (N_40918,N_39902,N_37823);
nor U40919 (N_40919,N_39823,N_39693);
nor U40920 (N_40920,N_38217,N_37518);
xor U40921 (N_40921,N_39790,N_39698);
nand U40922 (N_40922,N_37850,N_37871);
xor U40923 (N_40923,N_38729,N_38863);
xor U40924 (N_40924,N_38221,N_39699);
or U40925 (N_40925,N_38385,N_39711);
and U40926 (N_40926,N_38400,N_37574);
nand U40927 (N_40927,N_37766,N_39232);
xnor U40928 (N_40928,N_37963,N_38022);
and U40929 (N_40929,N_39039,N_39643);
or U40930 (N_40930,N_39098,N_38049);
xor U40931 (N_40931,N_39989,N_37702);
or U40932 (N_40932,N_38356,N_38153);
or U40933 (N_40933,N_38358,N_39118);
xor U40934 (N_40934,N_38792,N_38350);
xnor U40935 (N_40935,N_39127,N_37879);
or U40936 (N_40936,N_38949,N_37958);
and U40937 (N_40937,N_38665,N_37876);
nor U40938 (N_40938,N_37722,N_39204);
nor U40939 (N_40939,N_39448,N_38885);
and U40940 (N_40940,N_38629,N_37693);
xor U40941 (N_40941,N_39619,N_39592);
and U40942 (N_40942,N_39545,N_39676);
nand U40943 (N_40943,N_39671,N_37713);
or U40944 (N_40944,N_38642,N_38802);
and U40945 (N_40945,N_39121,N_39384);
or U40946 (N_40946,N_39397,N_39295);
nand U40947 (N_40947,N_38034,N_39274);
nor U40948 (N_40948,N_38387,N_37887);
and U40949 (N_40949,N_38094,N_38709);
nand U40950 (N_40950,N_39287,N_39172);
nor U40951 (N_40951,N_38940,N_38305);
nand U40952 (N_40952,N_38346,N_38553);
or U40953 (N_40953,N_37985,N_37751);
and U40954 (N_40954,N_39145,N_38724);
xor U40955 (N_40955,N_38784,N_37604);
and U40956 (N_40956,N_38681,N_37647);
or U40957 (N_40957,N_38363,N_38210);
or U40958 (N_40958,N_37842,N_39350);
or U40959 (N_40959,N_39474,N_38993);
and U40960 (N_40960,N_39813,N_38600);
nor U40961 (N_40961,N_39489,N_39152);
and U40962 (N_40962,N_39702,N_39086);
nor U40963 (N_40963,N_37666,N_38581);
xor U40964 (N_40964,N_38080,N_37757);
nand U40965 (N_40965,N_38201,N_39225);
nor U40966 (N_40966,N_39087,N_39345);
xor U40967 (N_40967,N_37635,N_38793);
xor U40968 (N_40968,N_39354,N_39419);
or U40969 (N_40969,N_38357,N_37810);
nand U40970 (N_40970,N_38329,N_39148);
nor U40971 (N_40971,N_38988,N_37753);
nand U40972 (N_40972,N_39637,N_39529);
nor U40973 (N_40973,N_39144,N_38919);
and U40974 (N_40974,N_39405,N_39266);
nand U40975 (N_40975,N_39959,N_38660);
nor U40976 (N_40976,N_38018,N_38218);
or U40977 (N_40977,N_38417,N_38303);
and U40978 (N_40978,N_38639,N_38833);
xnor U40979 (N_40979,N_38586,N_39743);
nor U40980 (N_40980,N_37615,N_38762);
xnor U40981 (N_40981,N_38798,N_39604);
nor U40982 (N_40982,N_38816,N_37939);
and U40983 (N_40983,N_39917,N_38783);
and U40984 (N_40984,N_39631,N_38073);
nor U40985 (N_40985,N_39772,N_39930);
and U40986 (N_40986,N_39107,N_39565);
and U40987 (N_40987,N_39330,N_38702);
or U40988 (N_40988,N_37990,N_39005);
nand U40989 (N_40989,N_39920,N_37609);
and U40990 (N_40990,N_37593,N_38390);
nand U40991 (N_40991,N_39809,N_38347);
and U40992 (N_40992,N_38878,N_38211);
and U40993 (N_40993,N_39043,N_38291);
nand U40994 (N_40994,N_39411,N_38149);
and U40995 (N_40995,N_39326,N_39610);
nor U40996 (N_40996,N_39572,N_38887);
nand U40997 (N_40997,N_38477,N_38297);
xnor U40998 (N_40998,N_39336,N_38274);
or U40999 (N_40999,N_39047,N_39624);
and U41000 (N_41000,N_37576,N_38404);
nand U41001 (N_41001,N_38416,N_38116);
and U41002 (N_41002,N_39292,N_38785);
xor U41003 (N_41003,N_39333,N_38813);
nor U41004 (N_41004,N_38527,N_39331);
nand U41005 (N_41005,N_37579,N_37761);
or U41006 (N_41006,N_39133,N_38587);
xnor U41007 (N_41007,N_39014,N_39765);
xor U41008 (N_41008,N_39346,N_38617);
xnor U41009 (N_41009,N_39224,N_39205);
xnor U41010 (N_41010,N_39960,N_37742);
xor U41011 (N_41011,N_38397,N_39304);
nand U41012 (N_41012,N_39181,N_38759);
nand U41013 (N_41013,N_38620,N_38692);
nor U41014 (N_41014,N_39201,N_39964);
nand U41015 (N_41015,N_38059,N_39636);
and U41016 (N_41016,N_38712,N_38242);
nand U41017 (N_41017,N_38310,N_37915);
nand U41018 (N_41018,N_37613,N_37894);
nor U41019 (N_41019,N_39149,N_39338);
nand U41020 (N_41020,N_39943,N_38797);
and U41021 (N_41021,N_39502,N_37565);
or U41022 (N_41022,N_37655,N_37938);
xnor U41023 (N_41023,N_39481,N_39342);
or U41024 (N_41024,N_37625,N_38533);
and U41025 (N_41025,N_38109,N_39883);
and U41026 (N_41026,N_38737,N_38381);
and U41027 (N_41027,N_38131,N_38373);
nand U41028 (N_41028,N_38122,N_38967);
and U41029 (N_41029,N_39212,N_39672);
xor U41030 (N_41030,N_39441,N_39210);
xor U41031 (N_41031,N_37865,N_39620);
or U41032 (N_41032,N_39008,N_38754);
or U41033 (N_41033,N_39616,N_37541);
or U41034 (N_41034,N_39831,N_38253);
and U41035 (N_41035,N_39775,N_37738);
or U41036 (N_41036,N_39242,N_38841);
xor U41037 (N_41037,N_39348,N_38096);
nand U41038 (N_41038,N_38572,N_39072);
and U41039 (N_41039,N_38352,N_38611);
and U41040 (N_41040,N_38238,N_39093);
nor U41041 (N_41041,N_39762,N_38889);
nor U41042 (N_41042,N_39271,N_38066);
or U41043 (N_41043,N_39284,N_38658);
or U41044 (N_41044,N_37967,N_39019);
xnor U41045 (N_41045,N_38471,N_38680);
nand U41046 (N_41046,N_39818,N_38178);
xor U41047 (N_41047,N_38481,N_39722);
or U41048 (N_41048,N_37623,N_39583);
xor U41049 (N_41049,N_38340,N_37592);
nand U41050 (N_41050,N_38194,N_38514);
and U41051 (N_41051,N_38795,N_39602);
xor U41052 (N_41052,N_39744,N_38469);
and U41053 (N_41053,N_37562,N_38685);
nand U41054 (N_41054,N_38750,N_37654);
xor U41055 (N_41055,N_39673,N_39192);
nor U41056 (N_41056,N_37838,N_38396);
or U41057 (N_41057,N_38321,N_39747);
nand U41058 (N_41058,N_37984,N_38374);
or U41059 (N_41059,N_38614,N_37630);
and U41060 (N_41060,N_38247,N_39893);
or U41061 (N_41061,N_38554,N_37670);
nand U41062 (N_41062,N_39973,N_38926);
xor U41063 (N_41063,N_39840,N_39689);
or U41064 (N_41064,N_38370,N_39512);
nor U41065 (N_41065,N_39026,N_38284);
nor U41066 (N_41066,N_39229,N_37897);
or U41067 (N_41067,N_37532,N_38407);
nor U41068 (N_41068,N_39679,N_37595);
nand U41069 (N_41069,N_39912,N_37677);
nand U41070 (N_41070,N_38082,N_39071);
nand U41071 (N_41071,N_37524,N_38294);
xor U41072 (N_41072,N_39727,N_39067);
and U41073 (N_41073,N_38470,N_38809);
or U41074 (N_41074,N_38133,N_38584);
xnor U41075 (N_41075,N_39961,N_37954);
and U41076 (N_41076,N_39394,N_38017);
or U41077 (N_41077,N_37890,N_39236);
or U41078 (N_41078,N_39484,N_39421);
or U41079 (N_41079,N_38012,N_38462);
nor U41080 (N_41080,N_39410,N_37874);
nor U41081 (N_41081,N_38463,N_38088);
nand U41082 (N_41082,N_38953,N_39537);
and U41083 (N_41083,N_38117,N_38343);
nand U41084 (N_41084,N_38325,N_39186);
nand U41085 (N_41085,N_37669,N_37989);
or U41086 (N_41086,N_38558,N_38126);
nand U41087 (N_41087,N_37837,N_38241);
nand U41088 (N_41088,N_39352,N_39443);
nor U41089 (N_41089,N_38522,N_39140);
nand U41090 (N_41090,N_38671,N_38351);
or U41091 (N_41091,N_38229,N_38497);
nor U41092 (N_41092,N_39017,N_37813);
xor U41093 (N_41093,N_39009,N_38331);
nand U41094 (N_41094,N_38969,N_38152);
and U41095 (N_41095,N_39884,N_38376);
and U41096 (N_41096,N_37668,N_39576);
or U41097 (N_41097,N_37760,N_38677);
or U41098 (N_41098,N_38412,N_39442);
or U41099 (N_41099,N_38379,N_38353);
or U41100 (N_41100,N_38545,N_39601);
nor U41101 (N_41101,N_39835,N_38956);
nand U41102 (N_41102,N_37816,N_39080);
xor U41103 (N_41103,N_38556,N_37705);
nor U41104 (N_41104,N_38818,N_38831);
xor U41105 (N_41105,N_39981,N_39706);
xnor U41106 (N_41106,N_39852,N_37557);
nand U41107 (N_41107,N_38752,N_38081);
or U41108 (N_41108,N_39490,N_38749);
xor U41109 (N_41109,N_39309,N_39875);
or U41110 (N_41110,N_38528,N_39432);
nor U41111 (N_41111,N_39078,N_39022);
and U41112 (N_41112,N_37899,N_38640);
xor U41113 (N_41113,N_39085,N_39719);
nand U41114 (N_41114,N_38495,N_39533);
or U41115 (N_41115,N_39363,N_39623);
xnor U41116 (N_41116,N_39429,N_38410);
and U41117 (N_41117,N_37784,N_39235);
or U41118 (N_41118,N_39555,N_38450);
or U41119 (N_41119,N_38146,N_38977);
or U41120 (N_41120,N_39720,N_38316);
nand U41121 (N_41121,N_38293,N_39150);
xnor U41122 (N_41122,N_39736,N_39939);
xor U41123 (N_41123,N_37517,N_37724);
nor U41124 (N_41124,N_39272,N_38973);
or U41125 (N_41125,N_38862,N_38780);
xor U41126 (N_41126,N_38037,N_39092);
xnor U41127 (N_41127,N_37743,N_38857);
nor U41128 (N_41128,N_39226,N_38078);
nor U41129 (N_41129,N_37941,N_37932);
or U41130 (N_41130,N_39356,N_39892);
nor U41131 (N_41131,N_38139,N_37926);
or U41132 (N_41132,N_38654,N_38104);
nand U41133 (N_41133,N_39846,N_38542);
nor U41134 (N_41134,N_38672,N_39909);
nor U41135 (N_41135,N_38192,N_39094);
xnor U41136 (N_41136,N_38348,N_39654);
or U41137 (N_41137,N_38295,N_38157);
nor U41138 (N_41138,N_39750,N_37825);
nand U41139 (N_41139,N_39801,N_38487);
xnor U41140 (N_41140,N_38591,N_38942);
xor U41141 (N_41141,N_39377,N_39334);
and U41142 (N_41142,N_37689,N_37783);
nand U41143 (N_41143,N_37906,N_39648);
or U41144 (N_41144,N_38304,N_38678);
nand U41145 (N_41145,N_38492,N_39575);
nand U41146 (N_41146,N_38872,N_39603);
or U41147 (N_41147,N_38939,N_39036);
nor U41148 (N_41148,N_38868,N_39409);
nand U41149 (N_41149,N_37510,N_38761);
nand U41150 (N_41150,N_38278,N_37949);
nand U41151 (N_41151,N_37646,N_38972);
nand U41152 (N_41152,N_37744,N_39010);
and U41153 (N_41153,N_37591,N_37726);
nand U41154 (N_41154,N_39202,N_39219);
xnor U41155 (N_41155,N_39141,N_38776);
nand U41156 (N_41156,N_38128,N_38546);
nand U41157 (N_41157,N_39100,N_37898);
or U41158 (N_41158,N_39894,N_38656);
nand U41159 (N_41159,N_39215,N_37617);
xor U41160 (N_41160,N_39589,N_39050);
and U41161 (N_41161,N_37585,N_38160);
xnor U41162 (N_41162,N_37797,N_39018);
or U41163 (N_41163,N_39933,N_38551);
and U41164 (N_41164,N_38272,N_38111);
xor U41165 (N_41165,N_38188,N_39886);
xnor U41166 (N_41166,N_37671,N_39721);
and U41167 (N_41167,N_39816,N_38843);
xnor U41168 (N_41168,N_38460,N_39524);
or U41169 (N_41169,N_38612,N_39556);
nor U41170 (N_41170,N_37721,N_39996);
nor U41171 (N_41171,N_38960,N_38398);
or U41172 (N_41172,N_39928,N_37586);
nor U41173 (N_41173,N_37933,N_39553);
or U41174 (N_41174,N_39962,N_37500);
and U41175 (N_41175,N_38169,N_37831);
nor U41176 (N_41176,N_39976,N_39952);
xnor U41177 (N_41177,N_38444,N_38962);
nor U41178 (N_41178,N_39773,N_39383);
nor U41179 (N_41179,N_39808,N_38118);
nor U41180 (N_41180,N_39426,N_37809);
nand U41181 (N_41181,N_39395,N_38249);
or U41182 (N_41182,N_38753,N_37567);
nand U41183 (N_41183,N_39787,N_39829);
nand U41184 (N_41184,N_39839,N_38601);
nand U41185 (N_41185,N_38322,N_38632);
nand U41186 (N_41186,N_39568,N_37919);
nor U41187 (N_41187,N_39027,N_39784);
nor U41188 (N_41188,N_39128,N_38636);
nor U41189 (N_41189,N_39661,N_39496);
nand U41190 (N_41190,N_37732,N_38787);
nor U41191 (N_41191,N_39013,N_38603);
nand U41192 (N_41192,N_37998,N_38870);
nor U41193 (N_41193,N_38282,N_39785);
xnor U41194 (N_41194,N_39163,N_38198);
nand U41195 (N_41195,N_39245,N_39945);
nand U41196 (N_41196,N_38269,N_38559);
nand U41197 (N_41197,N_38490,N_38309);
nor U41198 (N_41198,N_38035,N_38751);
xor U41199 (N_41199,N_39278,N_38986);
nand U41200 (N_41200,N_39855,N_37840);
xnor U41201 (N_41201,N_39860,N_37741);
nand U41202 (N_41202,N_38326,N_38641);
or U41203 (N_41203,N_38429,N_39057);
or U41204 (N_41204,N_39422,N_38850);
and U41205 (N_41205,N_39759,N_38423);
nor U41206 (N_41206,N_38173,N_39634);
nand U41207 (N_41207,N_38222,N_38336);
or U41208 (N_41208,N_39641,N_39492);
xor U41209 (N_41209,N_39612,N_39990);
nor U41210 (N_41210,N_37522,N_38683);
and U41211 (N_41211,N_39452,N_38306);
xnor U41212 (N_41212,N_38710,N_39200);
nor U41213 (N_41213,N_37733,N_37764);
nand U41214 (N_41214,N_38334,N_39139);
and U41215 (N_41215,N_39475,N_39544);
xor U41216 (N_41216,N_39707,N_38425);
or U41217 (N_41217,N_39313,N_38266);
and U41218 (N_41218,N_39460,N_39412);
and U41219 (N_41219,N_39255,N_39199);
xnor U41220 (N_41220,N_39316,N_37727);
xor U41221 (N_41221,N_38796,N_38371);
xor U41222 (N_41222,N_39258,N_38447);
nor U41223 (N_41223,N_39876,N_39079);
nand U41224 (N_41224,N_38705,N_37700);
nand U41225 (N_41225,N_38493,N_39862);
xnor U41226 (N_41226,N_38875,N_37620);
nor U41227 (N_41227,N_39877,N_38808);
nand U41228 (N_41228,N_38016,N_38399);
nand U41229 (N_41229,N_37652,N_37659);
nor U41230 (N_41230,N_38030,N_38908);
xor U41231 (N_41231,N_37771,N_39184);
nor U41232 (N_41232,N_38695,N_38936);
nor U41233 (N_41233,N_38838,N_39470);
nor U41234 (N_41234,N_39220,N_38520);
nor U41235 (N_41235,N_38008,N_38142);
or U41236 (N_41236,N_37629,N_37548);
nor U41237 (N_41237,N_37636,N_39268);
and U41238 (N_41238,N_39262,N_38670);
nand U41239 (N_41239,N_37538,N_38197);
nor U41240 (N_41240,N_38901,N_39798);
nand U41241 (N_41241,N_39101,N_39827);
or U41242 (N_41242,N_39729,N_38464);
nand U41243 (N_41243,N_39131,N_38691);
or U41244 (N_41244,N_38290,N_39083);
and U41245 (N_41245,N_38024,N_38478);
nor U41246 (N_41246,N_39521,N_39856);
or U41247 (N_41247,N_38079,N_38727);
xnor U41248 (N_41248,N_39963,N_38745);
xnor U41249 (N_41249,N_37588,N_38063);
xor U41250 (N_41250,N_39806,N_38119);
and U41251 (N_41251,N_39507,N_39407);
or U41252 (N_41252,N_37818,N_38330);
and U41253 (N_41253,N_37518,N_38032);
nor U41254 (N_41254,N_39332,N_38939);
nor U41255 (N_41255,N_38686,N_39017);
nor U41256 (N_41256,N_38081,N_37838);
and U41257 (N_41257,N_38306,N_38062);
or U41258 (N_41258,N_39686,N_38719);
xor U41259 (N_41259,N_39526,N_39479);
nand U41260 (N_41260,N_37740,N_39772);
nor U41261 (N_41261,N_39664,N_37504);
xor U41262 (N_41262,N_39542,N_37856);
nand U41263 (N_41263,N_37921,N_39478);
nand U41264 (N_41264,N_39152,N_38305);
nor U41265 (N_41265,N_39806,N_38251);
xnor U41266 (N_41266,N_39813,N_37768);
or U41267 (N_41267,N_38314,N_38745);
nor U41268 (N_41268,N_37689,N_39027);
or U41269 (N_41269,N_37748,N_39163);
and U41270 (N_41270,N_39321,N_37623);
xnor U41271 (N_41271,N_39212,N_38736);
nand U41272 (N_41272,N_38165,N_37917);
and U41273 (N_41273,N_39148,N_38263);
and U41274 (N_41274,N_38841,N_37782);
or U41275 (N_41275,N_37850,N_37516);
and U41276 (N_41276,N_39479,N_39618);
or U41277 (N_41277,N_38082,N_38526);
or U41278 (N_41278,N_39224,N_37666);
xnor U41279 (N_41279,N_39101,N_38684);
and U41280 (N_41280,N_37933,N_37640);
or U41281 (N_41281,N_38395,N_38566);
xor U41282 (N_41282,N_38581,N_39994);
and U41283 (N_41283,N_39326,N_39679);
and U41284 (N_41284,N_39893,N_39992);
or U41285 (N_41285,N_39259,N_38755);
xor U41286 (N_41286,N_38070,N_39866);
nand U41287 (N_41287,N_38621,N_38236);
nor U41288 (N_41288,N_39792,N_39331);
nand U41289 (N_41289,N_38908,N_37765);
xor U41290 (N_41290,N_38912,N_38693);
nor U41291 (N_41291,N_37543,N_39665);
nand U41292 (N_41292,N_38459,N_39969);
nor U41293 (N_41293,N_37828,N_38750);
or U41294 (N_41294,N_39355,N_39983);
nor U41295 (N_41295,N_38911,N_38421);
and U41296 (N_41296,N_38156,N_38636);
xnor U41297 (N_41297,N_39463,N_37877);
and U41298 (N_41298,N_39628,N_39027);
and U41299 (N_41299,N_37665,N_37696);
nor U41300 (N_41300,N_38721,N_38039);
nor U41301 (N_41301,N_38450,N_39086);
nand U41302 (N_41302,N_38759,N_38364);
or U41303 (N_41303,N_39525,N_37861);
and U41304 (N_41304,N_37618,N_39272);
and U41305 (N_41305,N_38064,N_38549);
nand U41306 (N_41306,N_39824,N_39589);
and U41307 (N_41307,N_39555,N_37863);
and U41308 (N_41308,N_38216,N_37662);
or U41309 (N_41309,N_38339,N_39843);
xnor U41310 (N_41310,N_39811,N_37785);
xor U41311 (N_41311,N_38712,N_39004);
and U41312 (N_41312,N_39803,N_38958);
nor U41313 (N_41313,N_38411,N_38634);
nand U41314 (N_41314,N_38555,N_39904);
or U41315 (N_41315,N_39882,N_37863);
and U41316 (N_41316,N_39182,N_39159);
or U41317 (N_41317,N_38838,N_39612);
nor U41318 (N_41318,N_39252,N_39799);
nor U41319 (N_41319,N_39177,N_38774);
and U41320 (N_41320,N_37957,N_37960);
or U41321 (N_41321,N_39648,N_38805);
or U41322 (N_41322,N_38094,N_38301);
or U41323 (N_41323,N_39774,N_38955);
nand U41324 (N_41324,N_39554,N_38312);
xnor U41325 (N_41325,N_37930,N_38658);
nand U41326 (N_41326,N_39938,N_39476);
and U41327 (N_41327,N_37926,N_39879);
xnor U41328 (N_41328,N_39744,N_39353);
xnor U41329 (N_41329,N_37674,N_39410);
nor U41330 (N_41330,N_38419,N_38933);
xnor U41331 (N_41331,N_39828,N_39231);
nand U41332 (N_41332,N_38233,N_39185);
nand U41333 (N_41333,N_38073,N_38856);
xnor U41334 (N_41334,N_37728,N_39306);
nand U41335 (N_41335,N_39601,N_38809);
or U41336 (N_41336,N_37637,N_38838);
nor U41337 (N_41337,N_39057,N_37691);
or U41338 (N_41338,N_37881,N_38823);
and U41339 (N_41339,N_39796,N_39110);
nor U41340 (N_41340,N_37720,N_39735);
nand U41341 (N_41341,N_37766,N_38975);
nand U41342 (N_41342,N_39354,N_39340);
nor U41343 (N_41343,N_39299,N_38695);
nor U41344 (N_41344,N_38439,N_39775);
or U41345 (N_41345,N_39074,N_38222);
nor U41346 (N_41346,N_39358,N_38291);
or U41347 (N_41347,N_38355,N_37868);
xor U41348 (N_41348,N_39772,N_38654);
xnor U41349 (N_41349,N_38205,N_38928);
nor U41350 (N_41350,N_39416,N_39797);
and U41351 (N_41351,N_37893,N_39732);
nand U41352 (N_41352,N_38722,N_39055);
or U41353 (N_41353,N_39035,N_39683);
nor U41354 (N_41354,N_38746,N_39541);
nor U41355 (N_41355,N_39544,N_39899);
xnor U41356 (N_41356,N_38896,N_38789);
xor U41357 (N_41357,N_38704,N_38020);
or U41358 (N_41358,N_38814,N_37558);
or U41359 (N_41359,N_39469,N_38418);
nand U41360 (N_41360,N_38626,N_38693);
nor U41361 (N_41361,N_37863,N_39572);
xor U41362 (N_41362,N_38508,N_37916);
or U41363 (N_41363,N_38982,N_39213);
xnor U41364 (N_41364,N_39314,N_38311);
xor U41365 (N_41365,N_39440,N_37787);
xnor U41366 (N_41366,N_38055,N_37529);
nor U41367 (N_41367,N_39377,N_39575);
nand U41368 (N_41368,N_37892,N_38886);
xnor U41369 (N_41369,N_39490,N_39384);
or U41370 (N_41370,N_39193,N_39933);
nand U41371 (N_41371,N_38192,N_38125);
nand U41372 (N_41372,N_39235,N_37586);
nor U41373 (N_41373,N_37780,N_38390);
and U41374 (N_41374,N_39840,N_39705);
or U41375 (N_41375,N_39589,N_39933);
nor U41376 (N_41376,N_38114,N_38297);
nor U41377 (N_41377,N_39899,N_39761);
nand U41378 (N_41378,N_39196,N_38994);
or U41379 (N_41379,N_37548,N_38992);
xor U41380 (N_41380,N_39013,N_37756);
xor U41381 (N_41381,N_39173,N_38930);
nand U41382 (N_41382,N_37534,N_38799);
nand U41383 (N_41383,N_37889,N_38306);
and U41384 (N_41384,N_39776,N_39679);
nor U41385 (N_41385,N_38708,N_39763);
nor U41386 (N_41386,N_37793,N_39498);
and U41387 (N_41387,N_39218,N_37972);
xnor U41388 (N_41388,N_39128,N_39809);
nand U41389 (N_41389,N_37517,N_38427);
nand U41390 (N_41390,N_39524,N_38975);
xor U41391 (N_41391,N_39194,N_37523);
xor U41392 (N_41392,N_37509,N_38522);
xor U41393 (N_41393,N_37873,N_37877);
xnor U41394 (N_41394,N_38795,N_38547);
nor U41395 (N_41395,N_38502,N_39329);
and U41396 (N_41396,N_38876,N_38029);
and U41397 (N_41397,N_39956,N_38316);
or U41398 (N_41398,N_38281,N_38678);
and U41399 (N_41399,N_39662,N_39245);
and U41400 (N_41400,N_38902,N_39514);
or U41401 (N_41401,N_38729,N_38925);
nor U41402 (N_41402,N_38082,N_39308);
and U41403 (N_41403,N_38384,N_39095);
nand U41404 (N_41404,N_39159,N_38186);
xnor U41405 (N_41405,N_38144,N_38228);
nor U41406 (N_41406,N_38093,N_39948);
xor U41407 (N_41407,N_39875,N_39638);
xnor U41408 (N_41408,N_37533,N_38875);
nand U41409 (N_41409,N_39203,N_38227);
or U41410 (N_41410,N_39112,N_39943);
xnor U41411 (N_41411,N_38169,N_39559);
and U41412 (N_41412,N_37845,N_38101);
and U41413 (N_41413,N_39035,N_39173);
or U41414 (N_41414,N_38288,N_38305);
and U41415 (N_41415,N_38529,N_38747);
and U41416 (N_41416,N_38201,N_39107);
nor U41417 (N_41417,N_39756,N_37845);
and U41418 (N_41418,N_39584,N_39830);
xor U41419 (N_41419,N_37874,N_39741);
nor U41420 (N_41420,N_38505,N_37828);
xnor U41421 (N_41421,N_37534,N_38748);
and U41422 (N_41422,N_39013,N_39402);
xor U41423 (N_41423,N_37731,N_39600);
xor U41424 (N_41424,N_37858,N_39594);
xor U41425 (N_41425,N_39823,N_39630);
xnor U41426 (N_41426,N_37915,N_39037);
or U41427 (N_41427,N_38107,N_39790);
or U41428 (N_41428,N_38122,N_39934);
nor U41429 (N_41429,N_38589,N_38834);
and U41430 (N_41430,N_38909,N_39549);
nand U41431 (N_41431,N_37943,N_37851);
xnor U41432 (N_41432,N_37891,N_39038);
nand U41433 (N_41433,N_39510,N_39686);
nand U41434 (N_41434,N_39917,N_37637);
nor U41435 (N_41435,N_39263,N_38483);
and U41436 (N_41436,N_38903,N_38465);
nand U41437 (N_41437,N_37890,N_38069);
nor U41438 (N_41438,N_39448,N_38781);
nand U41439 (N_41439,N_38407,N_39325);
or U41440 (N_41440,N_39124,N_39845);
nand U41441 (N_41441,N_39095,N_39995);
and U41442 (N_41442,N_39721,N_38907);
xor U41443 (N_41443,N_37505,N_37702);
and U41444 (N_41444,N_38843,N_37724);
nand U41445 (N_41445,N_37812,N_37505);
or U41446 (N_41446,N_38548,N_38975);
xor U41447 (N_41447,N_37850,N_39070);
or U41448 (N_41448,N_38728,N_39503);
nand U41449 (N_41449,N_38202,N_38946);
or U41450 (N_41450,N_38680,N_39905);
or U41451 (N_41451,N_39706,N_39138);
nand U41452 (N_41452,N_39039,N_39863);
and U41453 (N_41453,N_39428,N_38761);
xnor U41454 (N_41454,N_37532,N_38801);
nor U41455 (N_41455,N_37591,N_37921);
or U41456 (N_41456,N_37558,N_39262);
nor U41457 (N_41457,N_38925,N_37574);
xor U41458 (N_41458,N_39641,N_38539);
nor U41459 (N_41459,N_39617,N_39157);
or U41460 (N_41460,N_39261,N_38906);
or U41461 (N_41461,N_39727,N_38234);
and U41462 (N_41462,N_39100,N_39983);
nor U41463 (N_41463,N_37553,N_39635);
nand U41464 (N_41464,N_39390,N_38267);
nor U41465 (N_41465,N_38961,N_38340);
and U41466 (N_41466,N_38569,N_38539);
xor U41467 (N_41467,N_38616,N_39608);
or U41468 (N_41468,N_39440,N_39768);
nor U41469 (N_41469,N_38117,N_37790);
nand U41470 (N_41470,N_38293,N_39782);
nand U41471 (N_41471,N_39138,N_39616);
or U41472 (N_41472,N_37721,N_37509);
or U41473 (N_41473,N_38346,N_39249);
nor U41474 (N_41474,N_39983,N_39960);
and U41475 (N_41475,N_38529,N_39904);
nor U41476 (N_41476,N_39406,N_38409);
nand U41477 (N_41477,N_38790,N_37982);
xor U41478 (N_41478,N_38258,N_38362);
or U41479 (N_41479,N_38261,N_38276);
nand U41480 (N_41480,N_39353,N_38718);
or U41481 (N_41481,N_38429,N_38695);
nor U41482 (N_41482,N_39649,N_39580);
nor U41483 (N_41483,N_38898,N_38224);
and U41484 (N_41484,N_38739,N_39453);
or U41485 (N_41485,N_39184,N_37501);
or U41486 (N_41486,N_38501,N_38242);
xnor U41487 (N_41487,N_38465,N_38428);
nor U41488 (N_41488,N_37948,N_39598);
nor U41489 (N_41489,N_39058,N_38840);
nand U41490 (N_41490,N_39766,N_37606);
nand U41491 (N_41491,N_39385,N_39267);
xor U41492 (N_41492,N_38385,N_39707);
nor U41493 (N_41493,N_37547,N_38557);
or U41494 (N_41494,N_38296,N_38014);
nor U41495 (N_41495,N_39516,N_39222);
or U41496 (N_41496,N_38611,N_37867);
and U41497 (N_41497,N_38827,N_39545);
or U41498 (N_41498,N_38607,N_38782);
or U41499 (N_41499,N_39426,N_39035);
nand U41500 (N_41500,N_38810,N_39112);
nor U41501 (N_41501,N_38000,N_39638);
xor U41502 (N_41502,N_39481,N_38873);
or U41503 (N_41503,N_39872,N_39034);
and U41504 (N_41504,N_39713,N_37644);
nor U41505 (N_41505,N_39965,N_37509);
nor U41506 (N_41506,N_39985,N_37903);
or U41507 (N_41507,N_38113,N_37598);
and U41508 (N_41508,N_39161,N_39208);
xor U41509 (N_41509,N_38072,N_38117);
or U41510 (N_41510,N_38078,N_37865);
nor U41511 (N_41511,N_39942,N_37747);
or U41512 (N_41512,N_37658,N_39848);
and U41513 (N_41513,N_38669,N_37946);
nand U41514 (N_41514,N_39698,N_38580);
nor U41515 (N_41515,N_38970,N_38473);
or U41516 (N_41516,N_38442,N_38099);
nand U41517 (N_41517,N_38830,N_38767);
xor U41518 (N_41518,N_39197,N_39270);
nand U41519 (N_41519,N_38798,N_38916);
xnor U41520 (N_41520,N_38488,N_38219);
nand U41521 (N_41521,N_38275,N_38547);
and U41522 (N_41522,N_38844,N_38279);
xor U41523 (N_41523,N_38739,N_37703);
xnor U41524 (N_41524,N_39934,N_39945);
and U41525 (N_41525,N_39125,N_39724);
nor U41526 (N_41526,N_37802,N_37698);
nor U41527 (N_41527,N_39093,N_38048);
and U41528 (N_41528,N_38617,N_39011);
xor U41529 (N_41529,N_39407,N_38280);
or U41530 (N_41530,N_39429,N_38230);
nand U41531 (N_41531,N_38303,N_39011);
or U41532 (N_41532,N_39707,N_39857);
nand U41533 (N_41533,N_38807,N_37690);
nand U41534 (N_41534,N_38929,N_39076);
xor U41535 (N_41535,N_39602,N_39569);
or U41536 (N_41536,N_38821,N_39064);
and U41537 (N_41537,N_37985,N_38742);
xor U41538 (N_41538,N_39705,N_38530);
and U41539 (N_41539,N_37852,N_39027);
and U41540 (N_41540,N_39079,N_39617);
or U41541 (N_41541,N_38136,N_37784);
nand U41542 (N_41542,N_39512,N_38426);
or U41543 (N_41543,N_39487,N_38852);
xnor U41544 (N_41544,N_39443,N_38645);
and U41545 (N_41545,N_38193,N_37689);
and U41546 (N_41546,N_39418,N_38797);
nand U41547 (N_41547,N_39274,N_38801);
nor U41548 (N_41548,N_38700,N_39640);
or U41549 (N_41549,N_39383,N_39349);
or U41550 (N_41550,N_39066,N_38408);
or U41551 (N_41551,N_39095,N_39563);
xor U41552 (N_41552,N_39464,N_39606);
xnor U41553 (N_41553,N_39844,N_39739);
nand U41554 (N_41554,N_38224,N_37993);
and U41555 (N_41555,N_38393,N_39702);
nand U41556 (N_41556,N_38765,N_38215);
nand U41557 (N_41557,N_38276,N_38829);
or U41558 (N_41558,N_38552,N_39536);
xnor U41559 (N_41559,N_39358,N_39914);
xnor U41560 (N_41560,N_39427,N_37667);
nand U41561 (N_41561,N_37532,N_37850);
and U41562 (N_41562,N_38948,N_38525);
and U41563 (N_41563,N_39040,N_37639);
nor U41564 (N_41564,N_38704,N_38334);
and U41565 (N_41565,N_38669,N_38363);
nand U41566 (N_41566,N_38543,N_38736);
xor U41567 (N_41567,N_39062,N_38532);
nor U41568 (N_41568,N_38337,N_39646);
nor U41569 (N_41569,N_38665,N_39434);
nor U41570 (N_41570,N_37669,N_39522);
and U41571 (N_41571,N_39740,N_39264);
and U41572 (N_41572,N_37994,N_39680);
nand U41573 (N_41573,N_37986,N_38642);
or U41574 (N_41574,N_37675,N_38495);
or U41575 (N_41575,N_37544,N_39624);
nor U41576 (N_41576,N_39429,N_37583);
or U41577 (N_41577,N_37961,N_38129);
and U41578 (N_41578,N_39505,N_39332);
or U41579 (N_41579,N_38942,N_37941);
xor U41580 (N_41580,N_39475,N_37944);
or U41581 (N_41581,N_39796,N_39712);
nor U41582 (N_41582,N_38986,N_39641);
and U41583 (N_41583,N_38079,N_39478);
or U41584 (N_41584,N_37930,N_39690);
nor U41585 (N_41585,N_39099,N_38744);
nand U41586 (N_41586,N_37937,N_38946);
nor U41587 (N_41587,N_37656,N_38930);
and U41588 (N_41588,N_39496,N_37851);
nor U41589 (N_41589,N_39365,N_38241);
or U41590 (N_41590,N_38314,N_38107);
or U41591 (N_41591,N_39769,N_39775);
nor U41592 (N_41592,N_39522,N_38772);
or U41593 (N_41593,N_37847,N_38087);
xnor U41594 (N_41594,N_38033,N_38660);
xor U41595 (N_41595,N_38299,N_38683);
xor U41596 (N_41596,N_39758,N_38824);
nor U41597 (N_41597,N_38719,N_39708);
nor U41598 (N_41598,N_37960,N_38996);
nand U41599 (N_41599,N_38790,N_38718);
nor U41600 (N_41600,N_38262,N_39646);
and U41601 (N_41601,N_39652,N_38411);
xnor U41602 (N_41602,N_38934,N_39420);
and U41603 (N_41603,N_39032,N_37801);
xor U41604 (N_41604,N_38221,N_37784);
nor U41605 (N_41605,N_38219,N_39746);
and U41606 (N_41606,N_39654,N_39295);
nor U41607 (N_41607,N_37937,N_39505);
nor U41608 (N_41608,N_38722,N_37584);
or U41609 (N_41609,N_38821,N_38897);
nor U41610 (N_41610,N_38711,N_38882);
nor U41611 (N_41611,N_39608,N_39451);
nor U41612 (N_41612,N_39312,N_38405);
xor U41613 (N_41613,N_39342,N_38766);
xor U41614 (N_41614,N_39514,N_39850);
nand U41615 (N_41615,N_38061,N_39206);
nor U41616 (N_41616,N_39032,N_38828);
nor U41617 (N_41617,N_37917,N_39328);
nor U41618 (N_41618,N_37608,N_38688);
and U41619 (N_41619,N_38600,N_38878);
or U41620 (N_41620,N_38860,N_37953);
nor U41621 (N_41621,N_39283,N_37643);
and U41622 (N_41622,N_37818,N_38342);
xor U41623 (N_41623,N_39928,N_38106);
xnor U41624 (N_41624,N_39732,N_38512);
xnor U41625 (N_41625,N_39780,N_39700);
and U41626 (N_41626,N_37558,N_39977);
and U41627 (N_41627,N_38577,N_37984);
and U41628 (N_41628,N_37711,N_38582);
or U41629 (N_41629,N_38369,N_39475);
and U41630 (N_41630,N_39237,N_38774);
nor U41631 (N_41631,N_39558,N_38172);
or U41632 (N_41632,N_37535,N_37938);
xor U41633 (N_41633,N_38484,N_37785);
nand U41634 (N_41634,N_37966,N_38288);
and U41635 (N_41635,N_39726,N_37807);
xnor U41636 (N_41636,N_37757,N_39841);
nor U41637 (N_41637,N_38698,N_37975);
nor U41638 (N_41638,N_39614,N_38440);
or U41639 (N_41639,N_39660,N_39970);
and U41640 (N_41640,N_37867,N_39725);
nand U41641 (N_41641,N_38230,N_38208);
and U41642 (N_41642,N_38000,N_39817);
or U41643 (N_41643,N_39876,N_39603);
and U41644 (N_41644,N_37615,N_37707);
and U41645 (N_41645,N_37910,N_38400);
nand U41646 (N_41646,N_39326,N_37884);
xor U41647 (N_41647,N_39898,N_38460);
nor U41648 (N_41648,N_39438,N_38990);
and U41649 (N_41649,N_39269,N_38659);
xnor U41650 (N_41650,N_39193,N_39917);
nand U41651 (N_41651,N_38974,N_37945);
and U41652 (N_41652,N_39503,N_38066);
xnor U41653 (N_41653,N_39730,N_38962);
nor U41654 (N_41654,N_39734,N_37703);
and U41655 (N_41655,N_38825,N_39740);
or U41656 (N_41656,N_38882,N_39540);
xor U41657 (N_41657,N_38714,N_39214);
or U41658 (N_41658,N_39738,N_37764);
and U41659 (N_41659,N_38856,N_39651);
nand U41660 (N_41660,N_39159,N_38759);
or U41661 (N_41661,N_39558,N_39653);
nand U41662 (N_41662,N_38211,N_37961);
nor U41663 (N_41663,N_37700,N_38761);
and U41664 (N_41664,N_39566,N_38102);
nand U41665 (N_41665,N_37680,N_38221);
or U41666 (N_41666,N_39724,N_39421);
nor U41667 (N_41667,N_38117,N_37702);
nor U41668 (N_41668,N_38640,N_39047);
nor U41669 (N_41669,N_38663,N_37521);
and U41670 (N_41670,N_38144,N_39214);
nor U41671 (N_41671,N_38319,N_39396);
and U41672 (N_41672,N_37646,N_37995);
and U41673 (N_41673,N_39435,N_39876);
or U41674 (N_41674,N_38454,N_39112);
nand U41675 (N_41675,N_39210,N_38422);
xor U41676 (N_41676,N_39203,N_39950);
nor U41677 (N_41677,N_38918,N_38793);
nand U41678 (N_41678,N_38823,N_37530);
nand U41679 (N_41679,N_38527,N_37528);
xnor U41680 (N_41680,N_39238,N_38766);
xnor U41681 (N_41681,N_37815,N_38003);
nor U41682 (N_41682,N_39984,N_37753);
nand U41683 (N_41683,N_39761,N_38632);
and U41684 (N_41684,N_39475,N_39891);
nand U41685 (N_41685,N_38721,N_39232);
nand U41686 (N_41686,N_38730,N_39860);
xor U41687 (N_41687,N_38997,N_39539);
nor U41688 (N_41688,N_38783,N_38866);
and U41689 (N_41689,N_39838,N_39179);
or U41690 (N_41690,N_37787,N_38082);
or U41691 (N_41691,N_39663,N_39152);
nor U41692 (N_41692,N_39461,N_38718);
nor U41693 (N_41693,N_39526,N_39120);
nor U41694 (N_41694,N_39538,N_39410);
nor U41695 (N_41695,N_37953,N_38098);
and U41696 (N_41696,N_39813,N_39649);
or U41697 (N_41697,N_37796,N_38590);
nor U41698 (N_41698,N_39280,N_39913);
or U41699 (N_41699,N_37759,N_38158);
or U41700 (N_41700,N_38839,N_38192);
xor U41701 (N_41701,N_37894,N_38744);
nand U41702 (N_41702,N_38458,N_37821);
nand U41703 (N_41703,N_37636,N_39839);
nand U41704 (N_41704,N_38765,N_37859);
nor U41705 (N_41705,N_38335,N_39571);
xor U41706 (N_41706,N_39775,N_39997);
and U41707 (N_41707,N_38903,N_39740);
or U41708 (N_41708,N_38717,N_39250);
and U41709 (N_41709,N_38148,N_37552);
nand U41710 (N_41710,N_37966,N_38678);
or U41711 (N_41711,N_37505,N_39939);
or U41712 (N_41712,N_38790,N_39839);
or U41713 (N_41713,N_38558,N_38926);
nor U41714 (N_41714,N_38018,N_39258);
xor U41715 (N_41715,N_39440,N_38611);
xor U41716 (N_41716,N_39595,N_38415);
nor U41717 (N_41717,N_39078,N_39648);
nor U41718 (N_41718,N_38509,N_38137);
xnor U41719 (N_41719,N_37867,N_39026);
or U41720 (N_41720,N_38939,N_38509);
nor U41721 (N_41721,N_39414,N_38344);
nand U41722 (N_41722,N_37923,N_38647);
xor U41723 (N_41723,N_37515,N_38604);
or U41724 (N_41724,N_37962,N_37523);
nor U41725 (N_41725,N_37695,N_39722);
xor U41726 (N_41726,N_37599,N_38725);
or U41727 (N_41727,N_39645,N_38445);
xor U41728 (N_41728,N_39292,N_37587);
nor U41729 (N_41729,N_37793,N_38256);
and U41730 (N_41730,N_38304,N_39671);
and U41731 (N_41731,N_38454,N_37805);
nor U41732 (N_41732,N_37660,N_39931);
or U41733 (N_41733,N_37560,N_37718);
and U41734 (N_41734,N_37823,N_38153);
nand U41735 (N_41735,N_38693,N_39819);
or U41736 (N_41736,N_39400,N_38700);
and U41737 (N_41737,N_38953,N_38830);
or U41738 (N_41738,N_38019,N_38603);
nand U41739 (N_41739,N_38038,N_39992);
or U41740 (N_41740,N_37689,N_39099);
or U41741 (N_41741,N_39311,N_39920);
nand U41742 (N_41742,N_38390,N_38550);
nand U41743 (N_41743,N_38895,N_37852);
nor U41744 (N_41744,N_38307,N_38663);
nor U41745 (N_41745,N_38189,N_37602);
nor U41746 (N_41746,N_38427,N_37631);
or U41747 (N_41747,N_39464,N_39378);
or U41748 (N_41748,N_37870,N_39878);
or U41749 (N_41749,N_37636,N_39874);
and U41750 (N_41750,N_39234,N_38576);
xor U41751 (N_41751,N_37707,N_37825);
nand U41752 (N_41752,N_37819,N_37769);
or U41753 (N_41753,N_39243,N_37642);
xnor U41754 (N_41754,N_38906,N_38475);
or U41755 (N_41755,N_39174,N_39663);
and U41756 (N_41756,N_39472,N_37503);
nor U41757 (N_41757,N_37909,N_39830);
nor U41758 (N_41758,N_37721,N_39621);
xor U41759 (N_41759,N_38892,N_39777);
or U41760 (N_41760,N_38608,N_39444);
nor U41761 (N_41761,N_39737,N_38491);
xnor U41762 (N_41762,N_37607,N_37594);
nor U41763 (N_41763,N_38605,N_37968);
nor U41764 (N_41764,N_37518,N_37724);
xor U41765 (N_41765,N_39938,N_39260);
nor U41766 (N_41766,N_38723,N_39807);
nor U41767 (N_41767,N_37749,N_38694);
xor U41768 (N_41768,N_39828,N_38625);
nand U41769 (N_41769,N_38410,N_39119);
or U41770 (N_41770,N_39279,N_39440);
or U41771 (N_41771,N_38202,N_38874);
or U41772 (N_41772,N_37974,N_39361);
nand U41773 (N_41773,N_39587,N_38038);
nor U41774 (N_41774,N_39512,N_39349);
nand U41775 (N_41775,N_38780,N_39190);
xnor U41776 (N_41776,N_39467,N_37831);
xor U41777 (N_41777,N_39811,N_39123);
xor U41778 (N_41778,N_39285,N_39139);
or U41779 (N_41779,N_38314,N_37511);
and U41780 (N_41780,N_39800,N_37922);
xnor U41781 (N_41781,N_38699,N_37547);
nand U41782 (N_41782,N_37607,N_38792);
xor U41783 (N_41783,N_38626,N_38563);
nand U41784 (N_41784,N_39791,N_39390);
and U41785 (N_41785,N_38765,N_37851);
xnor U41786 (N_41786,N_38244,N_37928);
nor U41787 (N_41787,N_38176,N_37680);
and U41788 (N_41788,N_39205,N_37768);
or U41789 (N_41789,N_39154,N_38365);
and U41790 (N_41790,N_37522,N_38193);
xnor U41791 (N_41791,N_38797,N_38911);
or U41792 (N_41792,N_39346,N_38684);
nand U41793 (N_41793,N_38028,N_39932);
or U41794 (N_41794,N_38351,N_39201);
or U41795 (N_41795,N_38911,N_39385);
nand U41796 (N_41796,N_39482,N_38575);
nand U41797 (N_41797,N_39248,N_38209);
xor U41798 (N_41798,N_38604,N_38265);
xnor U41799 (N_41799,N_39612,N_38971);
and U41800 (N_41800,N_39859,N_38785);
nor U41801 (N_41801,N_38301,N_38372);
nor U41802 (N_41802,N_38666,N_39006);
xnor U41803 (N_41803,N_37637,N_39980);
or U41804 (N_41804,N_38983,N_38845);
or U41805 (N_41805,N_39938,N_38268);
nand U41806 (N_41806,N_38389,N_38893);
xor U41807 (N_41807,N_39558,N_38354);
and U41808 (N_41808,N_38726,N_39848);
or U41809 (N_41809,N_39005,N_38675);
nor U41810 (N_41810,N_39817,N_38344);
or U41811 (N_41811,N_37974,N_37903);
nor U41812 (N_41812,N_37940,N_38370);
and U41813 (N_41813,N_39619,N_38018);
nor U41814 (N_41814,N_38983,N_38284);
nor U41815 (N_41815,N_37950,N_39950);
nor U41816 (N_41816,N_37548,N_37724);
nor U41817 (N_41817,N_37834,N_38282);
nor U41818 (N_41818,N_38619,N_39765);
or U41819 (N_41819,N_37919,N_38728);
or U41820 (N_41820,N_39471,N_38771);
nand U41821 (N_41821,N_38005,N_39000);
or U41822 (N_41822,N_39730,N_37780);
xor U41823 (N_41823,N_37539,N_39089);
and U41824 (N_41824,N_39680,N_37657);
and U41825 (N_41825,N_38513,N_39834);
nand U41826 (N_41826,N_39195,N_39503);
xnor U41827 (N_41827,N_37759,N_37700);
nor U41828 (N_41828,N_39568,N_39449);
nand U41829 (N_41829,N_38142,N_39460);
xnor U41830 (N_41830,N_39263,N_38697);
and U41831 (N_41831,N_38920,N_38011);
nand U41832 (N_41832,N_37644,N_37509);
xnor U41833 (N_41833,N_38840,N_39620);
or U41834 (N_41834,N_39940,N_38871);
and U41835 (N_41835,N_39943,N_38154);
or U41836 (N_41836,N_38561,N_38120);
nor U41837 (N_41837,N_38374,N_39896);
nor U41838 (N_41838,N_39784,N_39440);
nand U41839 (N_41839,N_39365,N_39179);
or U41840 (N_41840,N_39478,N_39243);
or U41841 (N_41841,N_39665,N_38038);
and U41842 (N_41842,N_38655,N_39422);
and U41843 (N_41843,N_38129,N_37510);
or U41844 (N_41844,N_38230,N_38552);
nor U41845 (N_41845,N_38149,N_39754);
xnor U41846 (N_41846,N_39414,N_39365);
or U41847 (N_41847,N_38158,N_39439);
and U41848 (N_41848,N_37730,N_37549);
nor U41849 (N_41849,N_39138,N_38545);
or U41850 (N_41850,N_38308,N_39133);
or U41851 (N_41851,N_37835,N_38955);
nor U41852 (N_41852,N_37578,N_37648);
nand U41853 (N_41853,N_39538,N_38391);
and U41854 (N_41854,N_39287,N_38684);
or U41855 (N_41855,N_37911,N_37794);
nor U41856 (N_41856,N_37845,N_39870);
or U41857 (N_41857,N_39172,N_39557);
nor U41858 (N_41858,N_38971,N_39574);
or U41859 (N_41859,N_38286,N_39577);
xor U41860 (N_41860,N_37536,N_38725);
xnor U41861 (N_41861,N_39075,N_38924);
or U41862 (N_41862,N_39165,N_39237);
and U41863 (N_41863,N_39077,N_37639);
xnor U41864 (N_41864,N_38110,N_38619);
nor U41865 (N_41865,N_37644,N_37524);
nand U41866 (N_41866,N_38416,N_38731);
xnor U41867 (N_41867,N_38753,N_38681);
nand U41868 (N_41868,N_39679,N_38023);
nand U41869 (N_41869,N_37960,N_38930);
xor U41870 (N_41870,N_38686,N_39934);
or U41871 (N_41871,N_38524,N_39392);
xor U41872 (N_41872,N_39501,N_39955);
nand U41873 (N_41873,N_38590,N_39095);
nor U41874 (N_41874,N_39631,N_38281);
and U41875 (N_41875,N_38928,N_38713);
and U41876 (N_41876,N_39786,N_39294);
xnor U41877 (N_41877,N_38499,N_39796);
nand U41878 (N_41878,N_38350,N_38471);
nand U41879 (N_41879,N_38666,N_39683);
nand U41880 (N_41880,N_38799,N_38564);
nand U41881 (N_41881,N_38016,N_38817);
xor U41882 (N_41882,N_38700,N_37823);
and U41883 (N_41883,N_39324,N_39613);
nand U41884 (N_41884,N_38018,N_38638);
xor U41885 (N_41885,N_38232,N_38945);
or U41886 (N_41886,N_39560,N_39856);
nor U41887 (N_41887,N_39382,N_37838);
nor U41888 (N_41888,N_39042,N_38614);
and U41889 (N_41889,N_37550,N_38304);
nand U41890 (N_41890,N_37673,N_38208);
nor U41891 (N_41891,N_38602,N_39868);
nand U41892 (N_41892,N_37855,N_38075);
and U41893 (N_41893,N_37562,N_39025);
and U41894 (N_41894,N_39641,N_38863);
nand U41895 (N_41895,N_39181,N_38966);
or U41896 (N_41896,N_39832,N_39631);
nand U41897 (N_41897,N_39576,N_38403);
nor U41898 (N_41898,N_38501,N_39526);
xnor U41899 (N_41899,N_39102,N_37836);
and U41900 (N_41900,N_39580,N_39955);
nand U41901 (N_41901,N_39987,N_39103);
nand U41902 (N_41902,N_37539,N_39307);
xor U41903 (N_41903,N_38809,N_39322);
and U41904 (N_41904,N_39688,N_38517);
and U41905 (N_41905,N_39481,N_38366);
nand U41906 (N_41906,N_37975,N_39103);
or U41907 (N_41907,N_37976,N_38454);
xnor U41908 (N_41908,N_37672,N_38593);
and U41909 (N_41909,N_38628,N_37678);
xnor U41910 (N_41910,N_38894,N_38880);
and U41911 (N_41911,N_38884,N_38583);
nand U41912 (N_41912,N_39269,N_39723);
nand U41913 (N_41913,N_38576,N_38895);
and U41914 (N_41914,N_38213,N_39138);
xor U41915 (N_41915,N_38013,N_38043);
nor U41916 (N_41916,N_39580,N_39651);
nand U41917 (N_41917,N_39947,N_38793);
nor U41918 (N_41918,N_38042,N_39744);
or U41919 (N_41919,N_37605,N_37883);
and U41920 (N_41920,N_38952,N_38652);
nor U41921 (N_41921,N_37943,N_38564);
nand U41922 (N_41922,N_38652,N_39971);
nor U41923 (N_41923,N_37783,N_39304);
and U41924 (N_41924,N_39583,N_38855);
or U41925 (N_41925,N_38007,N_38362);
and U41926 (N_41926,N_38528,N_37738);
nand U41927 (N_41927,N_37670,N_38003);
and U41928 (N_41928,N_39155,N_38067);
nor U41929 (N_41929,N_39976,N_38725);
or U41930 (N_41930,N_39793,N_39173);
nor U41931 (N_41931,N_37564,N_38529);
and U41932 (N_41932,N_39580,N_39738);
and U41933 (N_41933,N_39858,N_39334);
nand U41934 (N_41934,N_37629,N_38579);
nand U41935 (N_41935,N_38461,N_39754);
nor U41936 (N_41936,N_39444,N_39484);
xor U41937 (N_41937,N_39691,N_39411);
or U41938 (N_41938,N_38294,N_38207);
nand U41939 (N_41939,N_39108,N_39180);
or U41940 (N_41940,N_39240,N_37777);
or U41941 (N_41941,N_39406,N_39565);
nand U41942 (N_41942,N_39794,N_37934);
xor U41943 (N_41943,N_39752,N_39905);
nand U41944 (N_41944,N_37564,N_38818);
nand U41945 (N_41945,N_38083,N_37632);
nor U41946 (N_41946,N_39554,N_37516);
nor U41947 (N_41947,N_37590,N_37706);
or U41948 (N_41948,N_39268,N_39130);
nor U41949 (N_41949,N_37550,N_39526);
xnor U41950 (N_41950,N_37579,N_38922);
xor U41951 (N_41951,N_38842,N_39417);
xor U41952 (N_41952,N_39200,N_38943);
nand U41953 (N_41953,N_39828,N_38572);
or U41954 (N_41954,N_38076,N_39259);
nor U41955 (N_41955,N_38304,N_37627);
xnor U41956 (N_41956,N_37701,N_37837);
nand U41957 (N_41957,N_39450,N_38078);
nor U41958 (N_41958,N_37564,N_39472);
or U41959 (N_41959,N_39196,N_38654);
xnor U41960 (N_41960,N_38723,N_39189);
nor U41961 (N_41961,N_39012,N_39782);
and U41962 (N_41962,N_38384,N_37802);
nor U41963 (N_41963,N_38970,N_37615);
and U41964 (N_41964,N_39916,N_39133);
or U41965 (N_41965,N_38246,N_39143);
or U41966 (N_41966,N_39080,N_39014);
nand U41967 (N_41967,N_38272,N_38206);
nor U41968 (N_41968,N_38531,N_39369);
nand U41969 (N_41969,N_39154,N_38469);
and U41970 (N_41970,N_39605,N_38304);
xnor U41971 (N_41971,N_38581,N_38656);
nand U41972 (N_41972,N_38723,N_38647);
xnor U41973 (N_41973,N_39093,N_38274);
nor U41974 (N_41974,N_37863,N_39713);
nand U41975 (N_41975,N_37690,N_39928);
xnor U41976 (N_41976,N_38256,N_39276);
xnor U41977 (N_41977,N_38307,N_38491);
and U41978 (N_41978,N_39023,N_39602);
nor U41979 (N_41979,N_38963,N_39868);
nand U41980 (N_41980,N_38650,N_39946);
and U41981 (N_41981,N_38583,N_39176);
nand U41982 (N_41982,N_38170,N_37510);
or U41983 (N_41983,N_37514,N_39150);
xnor U41984 (N_41984,N_39107,N_39487);
xnor U41985 (N_41985,N_37845,N_38943);
or U41986 (N_41986,N_37846,N_37775);
xor U41987 (N_41987,N_39070,N_37934);
nand U41988 (N_41988,N_37827,N_38289);
xnor U41989 (N_41989,N_39161,N_37667);
nor U41990 (N_41990,N_38690,N_37984);
or U41991 (N_41991,N_39625,N_37804);
nand U41992 (N_41992,N_38188,N_39922);
or U41993 (N_41993,N_39400,N_38729);
and U41994 (N_41994,N_38079,N_37554);
or U41995 (N_41995,N_37559,N_39886);
and U41996 (N_41996,N_38332,N_37638);
and U41997 (N_41997,N_37574,N_38405);
nor U41998 (N_41998,N_38417,N_39903);
or U41999 (N_41999,N_37587,N_38661);
or U42000 (N_42000,N_39291,N_38706);
nor U42001 (N_42001,N_38207,N_38165);
and U42002 (N_42002,N_38651,N_38722);
and U42003 (N_42003,N_38520,N_39467);
and U42004 (N_42004,N_39592,N_39389);
or U42005 (N_42005,N_39007,N_39443);
and U42006 (N_42006,N_39366,N_38974);
nand U42007 (N_42007,N_38610,N_38900);
nand U42008 (N_42008,N_39509,N_37898);
xor U42009 (N_42009,N_38550,N_38883);
xor U42010 (N_42010,N_39230,N_38283);
xor U42011 (N_42011,N_38646,N_38235);
and U42012 (N_42012,N_39362,N_38870);
nor U42013 (N_42013,N_38139,N_37541);
xnor U42014 (N_42014,N_38758,N_38384);
or U42015 (N_42015,N_37729,N_39325);
xor U42016 (N_42016,N_38158,N_38683);
nand U42017 (N_42017,N_37624,N_38414);
and U42018 (N_42018,N_38966,N_39660);
nor U42019 (N_42019,N_38201,N_37948);
nor U42020 (N_42020,N_37542,N_38685);
and U42021 (N_42021,N_39286,N_39815);
nand U42022 (N_42022,N_39263,N_38996);
nor U42023 (N_42023,N_38042,N_38117);
xnor U42024 (N_42024,N_38855,N_39304);
xnor U42025 (N_42025,N_39213,N_39670);
nor U42026 (N_42026,N_39282,N_39218);
nand U42027 (N_42027,N_39090,N_38067);
and U42028 (N_42028,N_39967,N_39784);
or U42029 (N_42029,N_38958,N_37564);
nand U42030 (N_42030,N_38840,N_38334);
and U42031 (N_42031,N_37862,N_39864);
or U42032 (N_42032,N_39765,N_37994);
or U42033 (N_42033,N_39655,N_37815);
nand U42034 (N_42034,N_39628,N_38107);
nor U42035 (N_42035,N_39519,N_39778);
xnor U42036 (N_42036,N_39369,N_38229);
xor U42037 (N_42037,N_39633,N_38538);
nand U42038 (N_42038,N_38785,N_38268);
nor U42039 (N_42039,N_37855,N_38569);
nand U42040 (N_42040,N_38474,N_38238);
nor U42041 (N_42041,N_39788,N_39470);
nand U42042 (N_42042,N_39304,N_38697);
and U42043 (N_42043,N_38783,N_39276);
or U42044 (N_42044,N_37737,N_38144);
and U42045 (N_42045,N_38221,N_39167);
or U42046 (N_42046,N_38955,N_39449);
nor U42047 (N_42047,N_37823,N_39510);
nand U42048 (N_42048,N_38709,N_39109);
nor U42049 (N_42049,N_37655,N_39702);
xnor U42050 (N_42050,N_39246,N_37739);
xor U42051 (N_42051,N_39207,N_39205);
nand U42052 (N_42052,N_38499,N_39555);
xnor U42053 (N_42053,N_38590,N_37946);
or U42054 (N_42054,N_37750,N_37859);
or U42055 (N_42055,N_38838,N_38735);
nand U42056 (N_42056,N_39090,N_37682);
and U42057 (N_42057,N_38345,N_39350);
nand U42058 (N_42058,N_39437,N_39649);
and U42059 (N_42059,N_38553,N_38409);
xor U42060 (N_42060,N_37625,N_38447);
nor U42061 (N_42061,N_38850,N_38213);
and U42062 (N_42062,N_39165,N_38895);
nor U42063 (N_42063,N_38220,N_39224);
nand U42064 (N_42064,N_38425,N_39725);
or U42065 (N_42065,N_37576,N_38150);
and U42066 (N_42066,N_38423,N_37881);
nand U42067 (N_42067,N_38095,N_39465);
or U42068 (N_42068,N_37581,N_39834);
nor U42069 (N_42069,N_37910,N_38054);
xor U42070 (N_42070,N_38974,N_38939);
and U42071 (N_42071,N_39645,N_38257);
nor U42072 (N_42072,N_39885,N_38367);
nand U42073 (N_42073,N_37816,N_38385);
xnor U42074 (N_42074,N_39474,N_39982);
and U42075 (N_42075,N_38726,N_39475);
nand U42076 (N_42076,N_38566,N_39889);
nand U42077 (N_42077,N_38877,N_38322);
nor U42078 (N_42078,N_37932,N_37653);
and U42079 (N_42079,N_38764,N_38000);
and U42080 (N_42080,N_38853,N_37844);
nand U42081 (N_42081,N_38506,N_37798);
xnor U42082 (N_42082,N_38344,N_38566);
or U42083 (N_42083,N_37691,N_38410);
nor U42084 (N_42084,N_39763,N_39298);
or U42085 (N_42085,N_38407,N_38831);
or U42086 (N_42086,N_39253,N_38961);
and U42087 (N_42087,N_39428,N_38304);
or U42088 (N_42088,N_38313,N_39074);
or U42089 (N_42089,N_38659,N_37524);
xor U42090 (N_42090,N_38561,N_39203);
xnor U42091 (N_42091,N_38183,N_39690);
and U42092 (N_42092,N_37666,N_39858);
and U42093 (N_42093,N_38602,N_37948);
xor U42094 (N_42094,N_37752,N_37885);
nor U42095 (N_42095,N_37859,N_37659);
and U42096 (N_42096,N_39183,N_37689);
nor U42097 (N_42097,N_39853,N_38913);
or U42098 (N_42098,N_39862,N_39279);
and U42099 (N_42099,N_38664,N_37680);
nand U42100 (N_42100,N_38458,N_37671);
nand U42101 (N_42101,N_37973,N_39070);
and U42102 (N_42102,N_38092,N_38486);
nor U42103 (N_42103,N_38625,N_39975);
nand U42104 (N_42104,N_37733,N_38484);
nand U42105 (N_42105,N_39557,N_39507);
and U42106 (N_42106,N_38207,N_39313);
xor U42107 (N_42107,N_39062,N_38558);
or U42108 (N_42108,N_38716,N_37524);
nand U42109 (N_42109,N_37796,N_39879);
and U42110 (N_42110,N_37528,N_37546);
xor U42111 (N_42111,N_38301,N_38154);
and U42112 (N_42112,N_38940,N_37926);
xor U42113 (N_42113,N_39179,N_38626);
xor U42114 (N_42114,N_38141,N_38772);
and U42115 (N_42115,N_38645,N_39263);
xnor U42116 (N_42116,N_39957,N_39473);
nor U42117 (N_42117,N_38691,N_39037);
nor U42118 (N_42118,N_37779,N_37661);
nor U42119 (N_42119,N_38400,N_38122);
nor U42120 (N_42120,N_38726,N_37504);
nor U42121 (N_42121,N_39778,N_39560);
xor U42122 (N_42122,N_39889,N_39395);
nor U42123 (N_42123,N_39369,N_38917);
nor U42124 (N_42124,N_38970,N_37877);
xnor U42125 (N_42125,N_39909,N_38655);
nor U42126 (N_42126,N_38110,N_38350);
or U42127 (N_42127,N_39427,N_39776);
or U42128 (N_42128,N_37648,N_37555);
or U42129 (N_42129,N_39810,N_38799);
nor U42130 (N_42130,N_38464,N_39388);
xor U42131 (N_42131,N_38174,N_38388);
nor U42132 (N_42132,N_39889,N_39717);
or U42133 (N_42133,N_39377,N_38879);
xnor U42134 (N_42134,N_37971,N_37722);
or U42135 (N_42135,N_38166,N_39151);
and U42136 (N_42136,N_39501,N_38537);
and U42137 (N_42137,N_37812,N_38762);
xor U42138 (N_42138,N_39251,N_37936);
and U42139 (N_42139,N_38721,N_39649);
nor U42140 (N_42140,N_38154,N_39931);
nor U42141 (N_42141,N_39894,N_39390);
xor U42142 (N_42142,N_38089,N_39991);
nor U42143 (N_42143,N_39240,N_38525);
or U42144 (N_42144,N_38558,N_38372);
and U42145 (N_42145,N_37891,N_38968);
xor U42146 (N_42146,N_37737,N_38109);
xor U42147 (N_42147,N_39396,N_38499);
and U42148 (N_42148,N_37696,N_37973);
nand U42149 (N_42149,N_37867,N_39710);
and U42150 (N_42150,N_38513,N_38787);
or U42151 (N_42151,N_39286,N_39460);
nor U42152 (N_42152,N_39484,N_39058);
nor U42153 (N_42153,N_38998,N_39721);
and U42154 (N_42154,N_37753,N_39009);
or U42155 (N_42155,N_37564,N_37862);
and U42156 (N_42156,N_39531,N_39403);
nor U42157 (N_42157,N_38010,N_38828);
and U42158 (N_42158,N_39404,N_38505);
or U42159 (N_42159,N_38414,N_38875);
nand U42160 (N_42160,N_38943,N_39998);
xnor U42161 (N_42161,N_39927,N_38987);
nand U42162 (N_42162,N_39864,N_38604);
nand U42163 (N_42163,N_38557,N_37980);
or U42164 (N_42164,N_38793,N_38547);
nor U42165 (N_42165,N_39839,N_38538);
and U42166 (N_42166,N_39722,N_37648);
nor U42167 (N_42167,N_39766,N_39015);
or U42168 (N_42168,N_37983,N_39745);
nor U42169 (N_42169,N_37849,N_38986);
nand U42170 (N_42170,N_39949,N_39061);
xnor U42171 (N_42171,N_38661,N_38123);
nor U42172 (N_42172,N_39401,N_38803);
or U42173 (N_42173,N_38657,N_39281);
nand U42174 (N_42174,N_37527,N_39343);
nor U42175 (N_42175,N_39614,N_38367);
xnor U42176 (N_42176,N_39234,N_37554);
nor U42177 (N_42177,N_37920,N_39809);
or U42178 (N_42178,N_37550,N_39478);
xor U42179 (N_42179,N_39823,N_39607);
and U42180 (N_42180,N_39796,N_37561);
xor U42181 (N_42181,N_38958,N_39309);
or U42182 (N_42182,N_38782,N_37527);
xnor U42183 (N_42183,N_38466,N_38321);
nor U42184 (N_42184,N_39490,N_39082);
nor U42185 (N_42185,N_37635,N_37820);
and U42186 (N_42186,N_39006,N_38948);
xnor U42187 (N_42187,N_39501,N_39480);
xor U42188 (N_42188,N_38857,N_38901);
or U42189 (N_42189,N_39372,N_39623);
xnor U42190 (N_42190,N_39885,N_38474);
nand U42191 (N_42191,N_39835,N_38873);
nor U42192 (N_42192,N_37865,N_38207);
xnor U42193 (N_42193,N_39414,N_39429);
xnor U42194 (N_42194,N_39561,N_39427);
and U42195 (N_42195,N_39559,N_38508);
xor U42196 (N_42196,N_38968,N_38777);
nand U42197 (N_42197,N_38970,N_38602);
and U42198 (N_42198,N_39108,N_39364);
nor U42199 (N_42199,N_39099,N_37515);
xor U42200 (N_42200,N_39942,N_38805);
nand U42201 (N_42201,N_38396,N_38099);
nor U42202 (N_42202,N_38467,N_38289);
or U42203 (N_42203,N_38518,N_39162);
nand U42204 (N_42204,N_37696,N_38535);
xnor U42205 (N_42205,N_38421,N_38197);
nand U42206 (N_42206,N_37509,N_39281);
nor U42207 (N_42207,N_39451,N_38611);
xor U42208 (N_42208,N_38955,N_39400);
or U42209 (N_42209,N_39408,N_39061);
nor U42210 (N_42210,N_38728,N_37743);
and U42211 (N_42211,N_39632,N_39545);
nor U42212 (N_42212,N_37533,N_39215);
nand U42213 (N_42213,N_38453,N_39678);
nand U42214 (N_42214,N_39496,N_37501);
and U42215 (N_42215,N_38870,N_38997);
nand U42216 (N_42216,N_38927,N_39563);
nand U42217 (N_42217,N_38473,N_38094);
nor U42218 (N_42218,N_37966,N_38850);
xnor U42219 (N_42219,N_39241,N_39868);
xor U42220 (N_42220,N_39380,N_37957);
or U42221 (N_42221,N_39269,N_39594);
or U42222 (N_42222,N_38827,N_39172);
nand U42223 (N_42223,N_37619,N_37861);
nand U42224 (N_42224,N_38456,N_38053);
nand U42225 (N_42225,N_39834,N_38915);
or U42226 (N_42226,N_38105,N_38644);
or U42227 (N_42227,N_39556,N_39318);
or U42228 (N_42228,N_39319,N_37685);
or U42229 (N_42229,N_38662,N_38083);
nor U42230 (N_42230,N_37520,N_38583);
and U42231 (N_42231,N_39703,N_39868);
and U42232 (N_42232,N_38350,N_38029);
or U42233 (N_42233,N_38923,N_38749);
nand U42234 (N_42234,N_38282,N_38355);
and U42235 (N_42235,N_39028,N_37646);
nor U42236 (N_42236,N_39775,N_39945);
nand U42237 (N_42237,N_37949,N_37931);
or U42238 (N_42238,N_39630,N_38876);
and U42239 (N_42239,N_38468,N_39827);
nand U42240 (N_42240,N_39224,N_38840);
nor U42241 (N_42241,N_39780,N_37872);
nor U42242 (N_42242,N_39889,N_39779);
nor U42243 (N_42243,N_39216,N_37596);
nand U42244 (N_42244,N_37823,N_37893);
xnor U42245 (N_42245,N_38429,N_38580);
and U42246 (N_42246,N_38664,N_37744);
nand U42247 (N_42247,N_37617,N_38946);
or U42248 (N_42248,N_38622,N_39132);
xor U42249 (N_42249,N_39049,N_39831);
and U42250 (N_42250,N_37761,N_39482);
or U42251 (N_42251,N_39382,N_38343);
nor U42252 (N_42252,N_37532,N_38154);
or U42253 (N_42253,N_39390,N_38945);
nand U42254 (N_42254,N_37893,N_39869);
nand U42255 (N_42255,N_37770,N_39479);
or U42256 (N_42256,N_37711,N_38474);
nor U42257 (N_42257,N_38108,N_38024);
xnor U42258 (N_42258,N_39773,N_37939);
nand U42259 (N_42259,N_39993,N_38313);
xor U42260 (N_42260,N_38547,N_38872);
nor U42261 (N_42261,N_37989,N_38490);
xor U42262 (N_42262,N_38239,N_38229);
or U42263 (N_42263,N_39061,N_39486);
or U42264 (N_42264,N_39685,N_37524);
nand U42265 (N_42265,N_39497,N_38482);
xnor U42266 (N_42266,N_37580,N_37617);
nand U42267 (N_42267,N_39366,N_38454);
nor U42268 (N_42268,N_38069,N_38449);
nand U42269 (N_42269,N_38784,N_39782);
or U42270 (N_42270,N_38238,N_39611);
xor U42271 (N_42271,N_38653,N_39350);
xnor U42272 (N_42272,N_37557,N_38388);
nor U42273 (N_42273,N_37605,N_37805);
or U42274 (N_42274,N_37591,N_38653);
nor U42275 (N_42275,N_37961,N_37670);
nand U42276 (N_42276,N_38309,N_37609);
or U42277 (N_42277,N_39193,N_38384);
nand U42278 (N_42278,N_38948,N_38638);
or U42279 (N_42279,N_37527,N_38157);
nor U42280 (N_42280,N_39090,N_39079);
nor U42281 (N_42281,N_37786,N_39570);
nand U42282 (N_42282,N_39394,N_38307);
nand U42283 (N_42283,N_38892,N_38528);
nor U42284 (N_42284,N_38347,N_38576);
nand U42285 (N_42285,N_39627,N_37894);
and U42286 (N_42286,N_39761,N_39333);
and U42287 (N_42287,N_38392,N_39050);
and U42288 (N_42288,N_38384,N_38470);
and U42289 (N_42289,N_39317,N_38094);
and U42290 (N_42290,N_39037,N_39910);
or U42291 (N_42291,N_39302,N_38170);
and U42292 (N_42292,N_37983,N_38966);
and U42293 (N_42293,N_39186,N_39317);
nand U42294 (N_42294,N_38105,N_39641);
nor U42295 (N_42295,N_38855,N_39284);
nand U42296 (N_42296,N_39729,N_38755);
or U42297 (N_42297,N_37622,N_39687);
and U42298 (N_42298,N_38045,N_38839);
xnor U42299 (N_42299,N_38043,N_38388);
or U42300 (N_42300,N_39603,N_39855);
nor U42301 (N_42301,N_39854,N_38164);
xor U42302 (N_42302,N_37677,N_37608);
xor U42303 (N_42303,N_38187,N_37811);
xnor U42304 (N_42304,N_39314,N_38316);
nor U42305 (N_42305,N_38841,N_39814);
nand U42306 (N_42306,N_38081,N_39556);
nand U42307 (N_42307,N_38362,N_39623);
xor U42308 (N_42308,N_37832,N_38282);
nor U42309 (N_42309,N_39982,N_38747);
xnor U42310 (N_42310,N_39395,N_39210);
nor U42311 (N_42311,N_37563,N_39088);
and U42312 (N_42312,N_39405,N_37994);
and U42313 (N_42313,N_39178,N_38414);
or U42314 (N_42314,N_39495,N_39819);
and U42315 (N_42315,N_38548,N_38360);
xor U42316 (N_42316,N_39996,N_39524);
and U42317 (N_42317,N_38931,N_38508);
nand U42318 (N_42318,N_38456,N_38181);
xor U42319 (N_42319,N_38640,N_38118);
nor U42320 (N_42320,N_39218,N_37712);
and U42321 (N_42321,N_38700,N_38126);
nor U42322 (N_42322,N_39530,N_38541);
nand U42323 (N_42323,N_38946,N_38373);
nand U42324 (N_42324,N_39188,N_38834);
nor U42325 (N_42325,N_37557,N_37919);
xnor U42326 (N_42326,N_37598,N_37968);
and U42327 (N_42327,N_38589,N_39681);
xnor U42328 (N_42328,N_38026,N_38380);
nand U42329 (N_42329,N_39518,N_39541);
nand U42330 (N_42330,N_39428,N_38552);
or U42331 (N_42331,N_37905,N_37729);
xnor U42332 (N_42332,N_38463,N_37632);
nor U42333 (N_42333,N_37889,N_38090);
nand U42334 (N_42334,N_39757,N_39992);
xnor U42335 (N_42335,N_37833,N_38750);
and U42336 (N_42336,N_38085,N_38684);
or U42337 (N_42337,N_39093,N_38589);
xnor U42338 (N_42338,N_37669,N_39940);
and U42339 (N_42339,N_38136,N_38456);
nor U42340 (N_42340,N_38039,N_39372);
xor U42341 (N_42341,N_39599,N_39042);
or U42342 (N_42342,N_39295,N_39071);
and U42343 (N_42343,N_39580,N_38662);
nor U42344 (N_42344,N_39695,N_38089);
and U42345 (N_42345,N_37722,N_38940);
nor U42346 (N_42346,N_39394,N_39959);
nor U42347 (N_42347,N_37680,N_38477);
xnor U42348 (N_42348,N_37550,N_39827);
nor U42349 (N_42349,N_38161,N_38540);
and U42350 (N_42350,N_38129,N_37697);
nor U42351 (N_42351,N_39114,N_37810);
xor U42352 (N_42352,N_38706,N_39201);
and U42353 (N_42353,N_39627,N_39962);
and U42354 (N_42354,N_38777,N_39893);
or U42355 (N_42355,N_37978,N_38224);
xor U42356 (N_42356,N_39131,N_37879);
and U42357 (N_42357,N_37549,N_37916);
nor U42358 (N_42358,N_37910,N_39786);
xnor U42359 (N_42359,N_39184,N_39041);
or U42360 (N_42360,N_38342,N_38514);
or U42361 (N_42361,N_37672,N_37857);
nand U42362 (N_42362,N_39028,N_38119);
nor U42363 (N_42363,N_39777,N_37768);
nand U42364 (N_42364,N_39387,N_38160);
nand U42365 (N_42365,N_39403,N_39514);
nand U42366 (N_42366,N_39003,N_39654);
and U42367 (N_42367,N_38418,N_38178);
nor U42368 (N_42368,N_38075,N_39358);
and U42369 (N_42369,N_39580,N_38589);
nand U42370 (N_42370,N_37792,N_38676);
or U42371 (N_42371,N_38246,N_38510);
xor U42372 (N_42372,N_38702,N_37871);
nand U42373 (N_42373,N_39038,N_39438);
nand U42374 (N_42374,N_39803,N_39411);
xnor U42375 (N_42375,N_39373,N_38752);
or U42376 (N_42376,N_38194,N_37535);
or U42377 (N_42377,N_39432,N_39671);
nor U42378 (N_42378,N_38640,N_39923);
and U42379 (N_42379,N_39238,N_37918);
and U42380 (N_42380,N_39905,N_37841);
nand U42381 (N_42381,N_39999,N_39995);
and U42382 (N_42382,N_38016,N_38096);
or U42383 (N_42383,N_38884,N_39739);
nand U42384 (N_42384,N_39906,N_39375);
nand U42385 (N_42385,N_39020,N_37864);
xnor U42386 (N_42386,N_38081,N_37984);
or U42387 (N_42387,N_39140,N_39726);
or U42388 (N_42388,N_39356,N_37877);
and U42389 (N_42389,N_38338,N_39514);
nand U42390 (N_42390,N_39587,N_38268);
nor U42391 (N_42391,N_37837,N_39331);
nand U42392 (N_42392,N_39672,N_38116);
and U42393 (N_42393,N_39884,N_38332);
nand U42394 (N_42394,N_37519,N_37550);
or U42395 (N_42395,N_39799,N_39694);
xor U42396 (N_42396,N_38483,N_38030);
and U42397 (N_42397,N_37549,N_38007);
xor U42398 (N_42398,N_37710,N_39210);
xnor U42399 (N_42399,N_38324,N_38147);
and U42400 (N_42400,N_38779,N_39179);
xnor U42401 (N_42401,N_38116,N_39858);
nor U42402 (N_42402,N_37622,N_37787);
and U42403 (N_42403,N_39432,N_39998);
and U42404 (N_42404,N_39194,N_38605);
nand U42405 (N_42405,N_37797,N_37668);
xnor U42406 (N_42406,N_39361,N_37920);
or U42407 (N_42407,N_39046,N_38003);
or U42408 (N_42408,N_37798,N_39001);
xnor U42409 (N_42409,N_37754,N_39624);
nand U42410 (N_42410,N_38550,N_39769);
or U42411 (N_42411,N_38153,N_37769);
or U42412 (N_42412,N_39230,N_39305);
nor U42413 (N_42413,N_37575,N_38754);
and U42414 (N_42414,N_39924,N_39697);
nand U42415 (N_42415,N_38209,N_38049);
xor U42416 (N_42416,N_38093,N_38553);
xor U42417 (N_42417,N_38185,N_39755);
xnor U42418 (N_42418,N_39149,N_39047);
nand U42419 (N_42419,N_37854,N_37783);
nor U42420 (N_42420,N_39579,N_39758);
xor U42421 (N_42421,N_37683,N_39178);
or U42422 (N_42422,N_38250,N_39748);
xor U42423 (N_42423,N_39143,N_37713);
nor U42424 (N_42424,N_38424,N_38396);
or U42425 (N_42425,N_37585,N_37995);
nor U42426 (N_42426,N_37835,N_39932);
xor U42427 (N_42427,N_38541,N_37970);
nand U42428 (N_42428,N_39595,N_37899);
nand U42429 (N_42429,N_38390,N_38431);
and U42430 (N_42430,N_39834,N_39458);
xnor U42431 (N_42431,N_39126,N_39404);
nand U42432 (N_42432,N_39080,N_38775);
nor U42433 (N_42433,N_38438,N_37790);
nand U42434 (N_42434,N_38029,N_39459);
nand U42435 (N_42435,N_39324,N_39729);
and U42436 (N_42436,N_38429,N_38691);
nor U42437 (N_42437,N_39963,N_38927);
nor U42438 (N_42438,N_38818,N_38485);
or U42439 (N_42439,N_39499,N_38634);
nand U42440 (N_42440,N_39259,N_38353);
and U42441 (N_42441,N_37874,N_38017);
nor U42442 (N_42442,N_38770,N_38296);
and U42443 (N_42443,N_38574,N_39943);
nor U42444 (N_42444,N_38992,N_37707);
nor U42445 (N_42445,N_38239,N_38963);
and U42446 (N_42446,N_38187,N_37595);
xor U42447 (N_42447,N_38825,N_37991);
xor U42448 (N_42448,N_39885,N_38258);
nor U42449 (N_42449,N_38967,N_38116);
or U42450 (N_42450,N_39460,N_38225);
xnor U42451 (N_42451,N_38037,N_38184);
or U42452 (N_42452,N_39142,N_38450);
xor U42453 (N_42453,N_37843,N_39027);
and U42454 (N_42454,N_38530,N_38053);
and U42455 (N_42455,N_38932,N_37903);
or U42456 (N_42456,N_38773,N_39927);
nor U42457 (N_42457,N_38466,N_39699);
or U42458 (N_42458,N_37855,N_38497);
nor U42459 (N_42459,N_38058,N_37997);
nand U42460 (N_42460,N_39609,N_38204);
and U42461 (N_42461,N_39184,N_37658);
or U42462 (N_42462,N_39281,N_37579);
and U42463 (N_42463,N_38489,N_38642);
and U42464 (N_42464,N_39081,N_38449);
nor U42465 (N_42465,N_38907,N_37548);
and U42466 (N_42466,N_39119,N_37869);
or U42467 (N_42467,N_39048,N_37603);
or U42468 (N_42468,N_37552,N_38969);
and U42469 (N_42469,N_39187,N_37835);
xnor U42470 (N_42470,N_39072,N_39260);
and U42471 (N_42471,N_38103,N_37580);
and U42472 (N_42472,N_37788,N_38441);
xnor U42473 (N_42473,N_39036,N_37733);
nor U42474 (N_42474,N_38574,N_38203);
xnor U42475 (N_42475,N_38587,N_39850);
xnor U42476 (N_42476,N_38038,N_39509);
or U42477 (N_42477,N_39887,N_39687);
nand U42478 (N_42478,N_39397,N_38359);
nor U42479 (N_42479,N_39228,N_38780);
nand U42480 (N_42480,N_37861,N_37638);
nand U42481 (N_42481,N_38760,N_39492);
nor U42482 (N_42482,N_38131,N_38542);
xnor U42483 (N_42483,N_38951,N_39528);
nand U42484 (N_42484,N_38363,N_39929);
nor U42485 (N_42485,N_39935,N_39230);
and U42486 (N_42486,N_37655,N_38269);
or U42487 (N_42487,N_38122,N_38176);
nand U42488 (N_42488,N_39597,N_37533);
or U42489 (N_42489,N_38959,N_39090);
nor U42490 (N_42490,N_39974,N_38927);
nor U42491 (N_42491,N_38147,N_38830);
nand U42492 (N_42492,N_38940,N_39133);
and U42493 (N_42493,N_39630,N_39977);
or U42494 (N_42494,N_39502,N_39625);
nand U42495 (N_42495,N_38843,N_38585);
nor U42496 (N_42496,N_37980,N_39804);
nor U42497 (N_42497,N_39982,N_38516);
and U42498 (N_42498,N_38580,N_38416);
nand U42499 (N_42499,N_38552,N_39245);
xnor U42500 (N_42500,N_42079,N_41988);
nand U42501 (N_42501,N_42024,N_40866);
and U42502 (N_42502,N_41587,N_41721);
nand U42503 (N_42503,N_41920,N_40144);
nor U42504 (N_42504,N_40595,N_41555);
and U42505 (N_42505,N_42311,N_41450);
and U42506 (N_42506,N_41709,N_42017);
xor U42507 (N_42507,N_41663,N_41342);
xnor U42508 (N_42508,N_40607,N_41614);
nor U42509 (N_42509,N_40703,N_40585);
and U42510 (N_42510,N_41627,N_42211);
xnor U42511 (N_42511,N_42253,N_41959);
xor U42512 (N_42512,N_41950,N_40831);
nor U42513 (N_42513,N_40734,N_40430);
nand U42514 (N_42514,N_41640,N_42153);
nor U42515 (N_42515,N_40971,N_41675);
or U42516 (N_42516,N_40209,N_41298);
nand U42517 (N_42517,N_42318,N_40551);
nor U42518 (N_42518,N_41641,N_41708);
xnor U42519 (N_42519,N_40077,N_40255);
and U42520 (N_42520,N_41690,N_41304);
xor U42521 (N_42521,N_42159,N_40745);
xnor U42522 (N_42522,N_42063,N_41102);
and U42523 (N_42523,N_40974,N_41666);
or U42524 (N_42524,N_42165,N_41412);
xnor U42525 (N_42525,N_42258,N_40966);
or U42526 (N_42526,N_41455,N_41445);
and U42527 (N_42527,N_42012,N_41389);
nand U42528 (N_42528,N_40402,N_40446);
nand U42529 (N_42529,N_42321,N_40435);
nand U42530 (N_42530,N_41140,N_41009);
xnor U42531 (N_42531,N_41317,N_40489);
nand U42532 (N_42532,N_40601,N_40915);
nand U42533 (N_42533,N_41846,N_40958);
xnor U42534 (N_42534,N_41778,N_40976);
xor U42535 (N_42535,N_42499,N_40955);
and U42536 (N_42536,N_41919,N_40740);
or U42537 (N_42537,N_40823,N_40818);
and U42538 (N_42538,N_41998,N_41377);
xnor U42539 (N_42539,N_41732,N_40796);
nor U42540 (N_42540,N_41073,N_40942);
and U42541 (N_42541,N_41507,N_40065);
nor U42542 (N_42542,N_41154,N_42131);
nand U42543 (N_42543,N_41972,N_40340);
nor U42544 (N_42544,N_40137,N_41814);
and U42545 (N_42545,N_40004,N_40512);
xnor U42546 (N_42546,N_42198,N_40559);
or U42547 (N_42547,N_41239,N_40706);
or U42548 (N_42548,N_41457,N_40509);
nor U42549 (N_42549,N_41247,N_41479);
nand U42550 (N_42550,N_40284,N_41250);
xor U42551 (N_42551,N_40968,N_40134);
xnor U42552 (N_42552,N_40461,N_42491);
nand U42553 (N_42553,N_41837,N_40550);
and U42554 (N_42554,N_40961,N_42465);
xor U42555 (N_42555,N_41206,N_41536);
nor U42556 (N_42556,N_40672,N_41053);
nand U42557 (N_42557,N_40313,N_41547);
nand U42558 (N_42558,N_41001,N_40462);
or U42559 (N_42559,N_42289,N_40693);
nand U42560 (N_42560,N_42046,N_40821);
xnor U42561 (N_42561,N_41993,N_42252);
or U42562 (N_42562,N_40241,N_40235);
nand U42563 (N_42563,N_41598,N_42039);
xnor U42564 (N_42564,N_41884,N_40094);
or U42565 (N_42565,N_40754,N_40609);
nor U42566 (N_42566,N_42002,N_41227);
nand U42567 (N_42567,N_40404,N_41753);
xor U42568 (N_42568,N_40376,N_42383);
and U42569 (N_42569,N_42105,N_41111);
or U42570 (N_42570,N_40702,N_41806);
nand U42571 (N_42571,N_40040,N_41222);
xnor U42572 (N_42572,N_41725,N_40309);
xor U42573 (N_42573,N_42379,N_41965);
or U42574 (N_42574,N_41251,N_41544);
and U42575 (N_42575,N_41231,N_40890);
and U42576 (N_42576,N_40417,N_42082);
nand U42577 (N_42577,N_41207,N_41116);
xnor U42578 (N_42578,N_40088,N_40036);
and U42579 (N_42579,N_41881,N_41918);
nor U42580 (N_42580,N_42224,N_41002);
nor U42581 (N_42581,N_42229,N_40501);
and U42582 (N_42582,N_40405,N_40939);
and U42583 (N_42583,N_40883,N_41411);
and U42584 (N_42584,N_40524,N_41233);
xor U42585 (N_42585,N_41015,N_40730);
nand U42586 (N_42586,N_41456,N_41962);
or U42587 (N_42587,N_40289,N_41296);
nor U42588 (N_42588,N_40649,N_40732);
and U42589 (N_42589,N_41785,N_40078);
nand U42590 (N_42590,N_41888,N_40247);
or U42591 (N_42591,N_40494,N_42120);
and U42592 (N_42592,N_42097,N_40673);
nand U42593 (N_42593,N_41451,N_40764);
nor U42594 (N_42594,N_40837,N_42133);
or U42595 (N_42595,N_41608,N_41285);
and U42596 (N_42596,N_41391,N_41243);
and U42597 (N_42597,N_41754,N_42042);
and U42598 (N_42598,N_42410,N_41063);
nand U42599 (N_42599,N_40026,N_42295);
nor U42600 (N_42600,N_41548,N_41356);
and U42601 (N_42601,N_40936,N_41392);
nor U42602 (N_42602,N_41973,N_42437);
or U42603 (N_42603,N_41804,N_40534);
xnor U42604 (N_42604,N_41299,N_40843);
or U42605 (N_42605,N_42006,N_40492);
xnor U42606 (N_42606,N_40502,N_41875);
xnor U42607 (N_42607,N_41664,N_41705);
nand U42608 (N_42608,N_40445,N_40024);
or U42609 (N_42609,N_41399,N_41008);
or U42610 (N_42610,N_40046,N_41007);
or U42611 (N_42611,N_42354,N_41513);
xor U42612 (N_42612,N_42325,N_42487);
or U42613 (N_42613,N_42247,N_40786);
or U42614 (N_42614,N_42449,N_40700);
and U42615 (N_42615,N_41030,N_41883);
nand U42616 (N_42616,N_41802,N_40272);
nand U42617 (N_42617,N_41596,N_41910);
nand U42618 (N_42618,N_41272,N_40119);
nand U42619 (N_42619,N_40620,N_41012);
xor U42620 (N_42620,N_40262,N_41280);
or U42621 (N_42621,N_40259,N_41812);
nor U42622 (N_42622,N_41937,N_40811);
or U42623 (N_42623,N_40029,N_42376);
and U42624 (N_42624,N_40989,N_42496);
nor U42625 (N_42625,N_42266,N_41694);
nor U42626 (N_42626,N_40467,N_41024);
xnor U42627 (N_42627,N_42186,N_42317);
and U42628 (N_42628,N_41398,N_41338);
xnor U42629 (N_42629,N_41543,N_42190);
and U42630 (N_42630,N_40882,N_41135);
nand U42631 (N_42631,N_41306,N_41620);
and U42632 (N_42632,N_41158,N_40816);
nand U42633 (N_42633,N_42112,N_42389);
xor U42634 (N_42634,N_40903,N_40741);
xnor U42635 (N_42635,N_41057,N_41617);
and U42636 (N_42636,N_41021,N_40378);
nor U42637 (N_42637,N_41677,N_41215);
nor U42638 (N_42638,N_41795,N_42044);
nand U42639 (N_42639,N_40973,N_40675);
or U42640 (N_42640,N_41890,N_42277);
nand U42641 (N_42641,N_41365,N_40248);
nor U42642 (N_42642,N_40617,N_40396);
nand U42643 (N_42643,N_42092,N_41773);
and U42644 (N_42644,N_40510,N_40229);
and U42645 (N_42645,N_42302,N_42430);
xnor U42646 (N_42646,N_40034,N_42156);
and U42647 (N_42647,N_40329,N_41626);
and U42648 (N_42648,N_41843,N_40047);
nor U42649 (N_42649,N_41560,N_41330);
or U42650 (N_42650,N_40710,N_42108);
nor U42651 (N_42651,N_41343,N_40564);
xnor U42652 (N_42652,N_41963,N_40577);
and U42653 (N_42653,N_42096,N_41538);
and U42654 (N_42654,N_40951,N_40182);
or U42655 (N_42655,N_41208,N_40932);
xnor U42656 (N_42656,N_40893,N_40493);
xor U42657 (N_42657,N_40170,N_40367);
and U42658 (N_42658,N_41047,N_42250);
xor U42659 (N_42659,N_42228,N_41006);
or U42660 (N_42660,N_41223,N_42132);
nand U42661 (N_42661,N_41136,N_42322);
and U42662 (N_42662,N_41258,N_40214);
or U42663 (N_42663,N_42148,N_40561);
nand U42664 (N_42664,N_42206,N_40257);
or U42665 (N_42665,N_40233,N_40850);
nor U42666 (N_42666,N_41145,N_40689);
and U42667 (N_42667,N_42005,N_42265);
or U42668 (N_42668,N_41696,N_40621);
or U42669 (N_42669,N_42257,N_42439);
or U42670 (N_42670,N_40148,N_42174);
nand U42671 (N_42671,N_41005,N_41246);
xnor U42672 (N_42672,N_40232,N_42427);
or U42673 (N_42673,N_41750,N_41410);
and U42674 (N_42674,N_40061,N_41681);
or U42675 (N_42675,N_40717,N_42492);
nor U42676 (N_42676,N_41000,N_41066);
and U42677 (N_42677,N_41686,N_40762);
or U42678 (N_42678,N_41613,N_40991);
and U42679 (N_42679,N_41413,N_41070);
nand U42680 (N_42680,N_42248,N_40436);
xor U42681 (N_42681,N_40071,N_41799);
and U42682 (N_42682,N_41662,N_42194);
nand U42683 (N_42683,N_40814,N_41147);
and U42684 (N_42684,N_41395,N_42087);
or U42685 (N_42685,N_41635,N_42320);
nand U42686 (N_42686,N_40964,N_41822);
or U42687 (N_42687,N_41935,N_41465);
nand U42688 (N_42688,N_41764,N_42454);
or U42689 (N_42689,N_40372,N_41446);
xnor U42690 (N_42690,N_40133,N_40881);
and U42691 (N_42691,N_40539,N_40149);
xnor U42692 (N_42692,N_41186,N_40569);
and U42693 (N_42693,N_40504,N_42388);
and U42694 (N_42694,N_40102,N_42184);
nor U42695 (N_42695,N_40031,N_40185);
nor U42696 (N_42696,N_41939,N_41194);
nand U42697 (N_42697,N_42381,N_41089);
xor U42698 (N_42698,N_40878,N_40836);
or U42699 (N_42699,N_42422,N_41037);
or U42700 (N_42700,N_40498,N_42009);
nor U42701 (N_42701,N_41228,N_40444);
nand U42702 (N_42702,N_42155,N_41311);
xor U42703 (N_42703,N_41344,N_42490);
and U42704 (N_42704,N_42141,N_41992);
nor U42705 (N_42705,N_40742,N_41575);
nor U42706 (N_42706,N_41895,N_41520);
nand U42707 (N_42707,N_42064,N_41847);
nand U42708 (N_42708,N_40195,N_40990);
xor U42709 (N_42709,N_40473,N_40200);
nand U42710 (N_42710,N_41436,N_41960);
or U42711 (N_42711,N_41758,N_40806);
xor U42712 (N_42712,N_40325,N_41362);
or U42713 (N_42713,N_42452,N_41909);
or U42714 (N_42714,N_40793,N_42134);
nor U42715 (N_42715,N_40364,N_41175);
or U42716 (N_42716,N_41531,N_41166);
or U42717 (N_42717,N_41320,N_40800);
and U42718 (N_42718,N_41373,N_41099);
or U42719 (N_42719,N_40797,N_42345);
nand U42720 (N_42720,N_40736,N_40535);
nand U42721 (N_42721,N_40937,N_42021);
nand U42722 (N_42722,N_41401,N_40483);
and U42723 (N_42723,N_42106,N_41284);
nor U42724 (N_42724,N_40008,N_40227);
xor U42725 (N_42725,N_41276,N_41938);
and U42726 (N_42726,N_40335,N_42406);
nand U42727 (N_42727,N_40027,N_40877);
and U42728 (N_42728,N_42426,N_40669);
xor U42729 (N_42729,N_42428,N_40645);
and U42730 (N_42730,N_40610,N_40129);
nor U42731 (N_42731,N_42489,N_42008);
xnor U42732 (N_42732,N_42110,N_41290);
xor U42733 (N_42733,N_42144,N_40900);
or U42734 (N_42734,N_42051,N_41076);
xnor U42735 (N_42735,N_42358,N_42371);
xnor U42736 (N_42736,N_40819,N_41271);
and U42737 (N_42737,N_42101,N_41085);
nand U42738 (N_42738,N_41218,N_42460);
nor U42739 (N_42739,N_41489,N_41984);
nand U42740 (N_42740,N_41482,N_40723);
and U42741 (N_42741,N_40316,N_42129);
and U42742 (N_42742,N_42209,N_41829);
nand U42743 (N_42743,N_40028,N_41490);
xnor U42744 (N_42744,N_40377,N_42204);
nand U42745 (N_42745,N_42037,N_40884);
xnor U42746 (N_42746,N_41660,N_41858);
and U42747 (N_42747,N_41093,N_41610);
nand U42748 (N_42748,N_41332,N_41865);
nor U42749 (N_42749,N_42377,N_41638);
or U42750 (N_42750,N_40727,N_41034);
and U42751 (N_42751,N_41232,N_41402);
nand U42752 (N_42752,N_41431,N_41683);
nor U42753 (N_42753,N_41331,N_40472);
and U42754 (N_42754,N_41882,N_41183);
nor U42755 (N_42755,N_40411,N_40712);
or U42756 (N_42756,N_42260,N_40676);
nor U42757 (N_42757,N_41958,N_41086);
nor U42758 (N_42758,N_40231,N_42226);
xor U42759 (N_42759,N_41711,N_41534);
or U42760 (N_42760,N_40537,N_41056);
and U42761 (N_42761,N_41966,N_40753);
xor U42762 (N_42762,N_40776,N_40245);
xnor U42763 (N_42763,N_40766,N_41226);
xor U42764 (N_42764,N_40326,N_41335);
nand U42765 (N_42765,N_41651,N_41771);
nand U42766 (N_42766,N_42275,N_42220);
nand U42767 (N_42767,N_41496,N_41794);
nor U42768 (N_42768,N_41872,N_40516);
nor U42769 (N_42769,N_41493,N_42058);
and U42770 (N_42770,N_41674,N_42059);
and U42771 (N_42771,N_40508,N_40923);
nand U42772 (N_42772,N_42154,N_41976);
xnor U42773 (N_42773,N_42472,N_40997);
and U42774 (N_42774,N_42035,N_42308);
xnor U42775 (N_42775,N_42337,N_41917);
nor U42776 (N_42776,N_40566,N_40197);
nor U42777 (N_42777,N_41607,N_42494);
nand U42778 (N_42778,N_40844,N_42103);
nand U42779 (N_42779,N_40117,N_40924);
nor U42780 (N_42780,N_41573,N_41191);
xor U42781 (N_42781,N_42353,N_40729);
nand U42782 (N_42782,N_40389,N_41355);
or U42783 (N_42783,N_40012,N_41945);
nand U42784 (N_42784,N_40708,N_40548);
nand U42785 (N_42785,N_42298,N_41472);
nor U42786 (N_42786,N_40292,N_41720);
xnor U42787 (N_42787,N_40327,N_40464);
nor U42788 (N_42788,N_41704,N_40875);
nand U42789 (N_42789,N_40661,N_42338);
nor U42790 (N_42790,N_40815,N_41670);
nor U42791 (N_42791,N_41813,N_42115);
or U42792 (N_42792,N_40021,N_41500);
xor U42793 (N_42793,N_41830,N_41975);
or U42794 (N_42794,N_40352,N_40168);
nand U42795 (N_42795,N_42399,N_41584);
nand U42796 (N_42796,N_40192,N_41484);
nand U42797 (N_42797,N_42125,N_42161);
nand U42798 (N_42798,N_42135,N_41755);
and U42799 (N_42799,N_42164,N_40637);
xnor U42800 (N_42800,N_41903,N_40523);
xor U42801 (N_42801,N_41114,N_40670);
xor U42802 (N_42802,N_41634,N_41551);
nand U42803 (N_42803,N_41756,N_41252);
and U42804 (N_42804,N_42301,N_41899);
xor U42805 (N_42805,N_41698,N_42196);
nor U42806 (N_42806,N_41418,N_40422);
nor U42807 (N_42807,N_40013,N_40840);
or U42808 (N_42808,N_41098,N_41078);
or U42809 (N_42809,N_41152,N_41556);
nor U42810 (N_42810,N_41928,N_40604);
nand U42811 (N_42811,N_40152,N_40159);
nor U42812 (N_42812,N_40629,N_41112);
or U42813 (N_42813,N_40089,N_41011);
or U42814 (N_42814,N_40981,N_41368);
xnor U42815 (N_42815,N_40290,N_42312);
nor U42816 (N_42816,N_41309,N_41458);
nor U42817 (N_42817,N_41644,N_40304);
xnor U42818 (N_42818,N_42294,N_42343);
xor U42819 (N_42819,N_40306,N_41775);
nor U42820 (N_42820,N_40506,N_40879);
nor U42821 (N_42821,N_42233,N_41748);
nor U42822 (N_42822,N_40362,N_41997);
and U42823 (N_42823,N_42384,N_40543);
or U42824 (N_42824,N_40400,N_40947);
and U42825 (N_42825,N_41557,N_40663);
xnor U42826 (N_42826,N_40401,N_41386);
and U42827 (N_42827,N_41502,N_41323);
nor U42828 (N_42828,N_41163,N_40808);
nand U42829 (N_42829,N_41321,N_41559);
nand U42830 (N_42830,N_42117,N_42483);
nand U42831 (N_42831,N_41808,N_42062);
nand U42832 (N_42832,N_42116,N_41160);
nand U42833 (N_42833,N_40346,N_40655);
or U42834 (N_42834,N_41891,N_41372);
xnor U42835 (N_42835,N_41853,N_42292);
xnor U42836 (N_42836,N_40941,N_41067);
or U42837 (N_42837,N_41254,N_40220);
nand U42838 (N_42838,N_40674,N_41943);
nor U42839 (N_42839,N_41390,N_40910);
nand U42840 (N_42840,N_42173,N_40748);
nand U42841 (N_42841,N_42176,N_42239);
nor U42842 (N_42842,N_40416,N_40563);
xnor U42843 (N_42843,N_40558,N_41653);
and U42844 (N_42844,N_42382,N_41952);
xnor U42845 (N_42845,N_40860,N_41027);
xor U42846 (N_42846,N_40511,N_40765);
and U42847 (N_42847,N_41878,N_40686);
nand U42848 (N_42848,N_42393,N_41054);
and U42849 (N_42849,N_40238,N_42394);
nand U42850 (N_42850,N_41713,N_40091);
or U42851 (N_42851,N_41549,N_41103);
xnor U42852 (N_42852,N_40781,N_41733);
and U42853 (N_42853,N_41915,N_41170);
or U42854 (N_42854,N_40809,N_42441);
and U42855 (N_42855,N_40758,N_41961);
nand U42856 (N_42856,N_41328,N_40145);
nand U42857 (N_42857,N_41026,N_40599);
and U42858 (N_42858,N_42149,N_42072);
nand U42859 (N_42859,N_41565,N_40805);
nor U42860 (N_42860,N_41369,N_40338);
nor U42861 (N_42861,N_41761,N_42109);
or U42862 (N_42862,N_40902,N_41521);
nand U42863 (N_42863,N_40279,N_40640);
xnor U42864 (N_42864,N_40442,N_40565);
nand U42865 (N_42865,N_42126,N_40994);
nand U42866 (N_42866,N_42438,N_40162);
or U42867 (N_42867,N_41022,N_42180);
nand U42868 (N_42868,N_40588,N_41550);
or U42869 (N_42869,N_41481,N_41768);
or U42870 (N_42870,N_40849,N_40050);
nand U42871 (N_42871,N_40798,N_40124);
nand U42872 (N_42872,N_41739,N_40591);
or U42873 (N_42873,N_40804,N_40186);
and U42874 (N_42874,N_41714,N_41319);
nand U42875 (N_42875,N_42231,N_40651);
nor U42876 (N_42876,N_41359,N_41429);
nor U42877 (N_42877,N_41759,N_41318);
nor U42878 (N_42878,N_41509,N_41564);
or U42879 (N_42879,N_41475,N_40810);
xnor U42880 (N_42880,N_40963,N_40048);
nor U42881 (N_42881,N_42130,N_40438);
xor U42882 (N_42882,N_41478,N_40908);
xor U42883 (N_42883,N_41715,N_42111);
xnor U42884 (N_42884,N_40383,N_40839);
nand U42885 (N_42885,N_40240,N_41762);
nor U42886 (N_42886,N_41236,N_41312);
xnor U42887 (N_42887,N_41927,N_42296);
nor U42888 (N_42888,N_41907,N_40449);
nor U42889 (N_42889,N_42171,N_40180);
or U42890 (N_42890,N_42276,N_40682);
xor U42891 (N_42891,N_41679,N_40488);
nor U42892 (N_42892,N_40190,N_41168);
or U42893 (N_42893,N_40600,N_42340);
or U42894 (N_42894,N_41645,N_42434);
nor U42895 (N_42895,N_42263,N_40847);
xnor U42896 (N_42896,N_41498,N_42205);
or U42897 (N_42897,N_40300,N_41454);
nand U42898 (N_42898,N_40332,N_41852);
nand U42899 (N_42899,N_40751,N_41108);
nor U42900 (N_42900,N_42259,N_42417);
nand U42901 (N_42901,N_40324,N_40905);
and U42902 (N_42902,N_41483,N_42177);
xor U42903 (N_42903,N_40965,N_40253);
and U42904 (N_42904,N_41642,N_41894);
xnor U42905 (N_42905,N_40533,N_40037);
nand U42906 (N_42906,N_40116,N_40140);
and U42907 (N_42907,N_40992,N_40624);
or U42908 (N_42908,N_41185,N_40169);
nor U42909 (N_42909,N_40618,N_40813);
nor U42910 (N_42910,N_40178,N_40330);
and U42911 (N_42911,N_40475,N_40101);
nand U42912 (N_42912,N_41126,N_42145);
or U42913 (N_42913,N_40746,N_40665);
xor U42914 (N_42914,N_42477,N_40474);
or U42915 (N_42915,N_41408,N_41581);
nand U42916 (N_42916,N_41810,N_42278);
nand U42917 (N_42917,N_40928,N_40086);
xnor U42918 (N_42918,N_40653,N_40221);
xor U42919 (N_42919,N_41876,N_41659);
xor U42920 (N_42920,N_40275,N_41133);
nand U42921 (N_42921,N_41148,N_41582);
or U42922 (N_42922,N_42251,N_41261);
xnor U42923 (N_42923,N_42331,N_41530);
nor U42924 (N_42924,N_41926,N_42307);
nand U42925 (N_42925,N_41908,N_42305);
or U42926 (N_42926,N_41120,N_41225);
xnor U42927 (N_42927,N_40421,N_41469);
nor U42928 (N_42928,N_41177,N_40977);
nand U42929 (N_42929,N_40782,N_42372);
nor U42930 (N_42930,N_42279,N_40580);
or U42931 (N_42931,N_40589,N_40288);
xnor U42932 (N_42932,N_42412,N_40911);
nor U42933 (N_42933,N_42081,N_41187);
nand U42934 (N_42934,N_41707,N_41791);
xor U42935 (N_42935,N_40542,N_41731);
xor U42936 (N_42936,N_42335,N_41691);
nor U42937 (N_42937,N_40830,N_41602);
and U42938 (N_42938,N_42241,N_42235);
nor U42939 (N_42939,N_41453,N_40590);
xor U42940 (N_42940,N_41699,N_41134);
nor U42941 (N_42941,N_42473,N_41374);
and U42942 (N_42942,N_40373,N_42032);
or U42943 (N_42943,N_40045,N_40722);
xor U42944 (N_42944,N_40778,N_40298);
or U42945 (N_42945,N_40656,N_40592);
xnor U42946 (N_42946,N_40154,N_41447);
or U42947 (N_42947,N_40032,N_42172);
xor U42948 (N_42948,N_40864,N_40230);
or U42949 (N_42949,N_42215,N_42359);
nand U42950 (N_42950,N_42055,N_41375);
nand U42951 (N_42951,N_42380,N_41801);
and U42952 (N_42952,N_41259,N_40070);
nand U42953 (N_42953,N_40455,N_41407);
nor U42954 (N_42954,N_42232,N_41379);
nor U42955 (N_42955,N_40581,N_41850);
or U42956 (N_42956,N_42398,N_40254);
nand U42957 (N_42957,N_40876,N_41836);
nor U42958 (N_42958,N_41864,N_41184);
or U42959 (N_42959,N_40852,N_41886);
xnor U42960 (N_42960,N_42004,N_40576);
nand U42961 (N_42961,N_41990,N_42498);
and U42962 (N_42962,N_40606,N_42027);
xnor U42963 (N_42963,N_40728,N_40153);
nor U42964 (N_42964,N_41511,N_41717);
or U42965 (N_42965,N_42396,N_40783);
or U42966 (N_42966,N_41036,N_41774);
and U42967 (N_42967,N_41578,N_42089);
and U42968 (N_42968,N_41572,N_42168);
and U42969 (N_42969,N_41084,N_41848);
or U42970 (N_42970,N_42182,N_40657);
nor U42971 (N_42971,N_40983,N_41081);
and U42972 (N_42972,N_42075,N_41562);
nor U42973 (N_42973,N_40978,N_40519);
nor U42974 (N_42974,N_42485,N_41570);
xor U42975 (N_42975,N_40268,N_40016);
or U42976 (N_42976,N_42467,N_41173);
xor U42977 (N_42977,N_41874,N_42474);
or U42978 (N_42978,N_42187,N_42351);
nand U42979 (N_42979,N_40068,N_40480);
nor U42980 (N_42980,N_42118,N_40419);
xnor U42981 (N_42981,N_40339,N_42071);
and U42982 (N_42982,N_42271,N_42476);
nor U42983 (N_42983,N_40586,N_41994);
nor U42984 (N_42984,N_40768,N_40820);
xor U42985 (N_42985,N_42214,N_41117);
nand U42986 (N_42986,N_41149,N_41817);
and U42987 (N_42987,N_40587,N_41090);
and U42988 (N_42988,N_40271,N_41786);
nor U42989 (N_42989,N_40921,N_41833);
nor U42990 (N_42990,N_40387,N_40451);
or U42991 (N_42991,N_42378,N_41612);
xor U42992 (N_42992,N_41912,N_40056);
xnor U42993 (N_42993,N_40320,N_41042);
and U42994 (N_42994,N_41684,N_40369);
or U42995 (N_42995,N_40395,N_40812);
nand U42996 (N_42996,N_40160,N_40156);
nand U42997 (N_42997,N_41180,N_40633);
or U42998 (N_42998,N_41189,N_40760);
or U42999 (N_42999,N_40536,N_40570);
and U43000 (N_43000,N_40613,N_40459);
or U43001 (N_43001,N_40164,N_42189);
and U43002 (N_43002,N_42234,N_40603);
or U43003 (N_43003,N_41256,N_41712);
xnor U43004 (N_43004,N_42053,N_41055);
and U43005 (N_43005,N_41658,N_41383);
xnor U43006 (N_43006,N_42392,N_40944);
nand U43007 (N_43007,N_41504,N_42025);
and U43008 (N_43008,N_40626,N_41657);
and U43009 (N_43009,N_41156,N_41887);
nor U43010 (N_43010,N_40064,N_41655);
or U43011 (N_43011,N_40052,N_41893);
and U43012 (N_43012,N_42256,N_42342);
or U43013 (N_43013,N_40943,N_41949);
nand U43014 (N_43014,N_41906,N_41260);
xnor U43015 (N_43015,N_42090,N_42185);
and U43016 (N_43016,N_41533,N_40215);
xnor U43017 (N_43017,N_40468,N_40582);
or U43018 (N_43018,N_40485,N_40496);
nor U43019 (N_43019,N_42033,N_42423);
or U43020 (N_43020,N_41980,N_42349);
nor U43021 (N_43021,N_41821,N_42113);
xor U43022 (N_43022,N_40769,N_40869);
and U43023 (N_43023,N_40948,N_41849);
or U43024 (N_43024,N_40891,N_42188);
nand U43025 (N_43025,N_41669,N_40108);
xnor U43026 (N_43026,N_40381,N_41800);
nor U43027 (N_43027,N_41028,N_41334);
nand U43028 (N_43028,N_40666,N_40286);
or U43029 (N_43029,N_40863,N_40406);
xnor U43030 (N_43030,N_42020,N_41703);
xor U43031 (N_43031,N_41201,N_40458);
and U43032 (N_43032,N_40249,N_41477);
xor U43033 (N_43033,N_41188,N_42362);
and U43034 (N_43034,N_42080,N_40022);
nand U43035 (N_43035,N_42245,N_41898);
or U43036 (N_43036,N_41671,N_42078);
or U43037 (N_43037,N_40956,N_40750);
nor U43038 (N_43038,N_42313,N_40246);
or U43039 (N_43039,N_40375,N_40683);
nor U43040 (N_43040,N_41097,N_41234);
nor U43041 (N_43041,N_41746,N_41956);
nand U43042 (N_43042,N_40774,N_40701);
and U43043 (N_43043,N_41196,N_41378);
nand U43044 (N_43044,N_40478,N_41491);
and U43045 (N_43045,N_41676,N_40125);
nor U43046 (N_43046,N_40322,N_41623);
xnor U43047 (N_43047,N_42076,N_41545);
xor U43048 (N_43048,N_41933,N_40092);
nand U43049 (N_43049,N_42334,N_41741);
or U43050 (N_43050,N_40625,N_41510);
xor U43051 (N_43051,N_40775,N_41592);
nand U43052 (N_43052,N_41648,N_42481);
nor U43053 (N_43053,N_40386,N_41265);
or U43054 (N_43054,N_42040,N_40738);
nand U43055 (N_43055,N_40889,N_41101);
nor U43056 (N_43056,N_41463,N_40393);
nor U43057 (N_43057,N_42385,N_40314);
and U43058 (N_43058,N_41245,N_40873);
and U43059 (N_43059,N_42453,N_41438);
nor U43060 (N_43060,N_40130,N_41032);
or U43061 (N_43061,N_41300,N_41591);
nand U43062 (N_43062,N_41440,N_40213);
xnor U43063 (N_43063,N_40846,N_41172);
xnor U43064 (N_43064,N_40010,N_41274);
or U43065 (N_43065,N_41724,N_40370);
nand U43066 (N_43066,N_41673,N_40042);
nand U43067 (N_43067,N_40055,N_41827);
nand U43068 (N_43068,N_41512,N_42143);
and U43069 (N_43069,N_41605,N_40526);
nand U43070 (N_43070,N_41722,N_41841);
nor U43071 (N_43071,N_40038,N_41210);
and U43072 (N_43072,N_42146,N_42306);
nor U43073 (N_43073,N_40243,N_40555);
nor U43074 (N_43074,N_40410,N_40407);
nand U43075 (N_43075,N_40895,N_42065);
nand U43076 (N_43076,N_41688,N_42218);
xor U43077 (N_43077,N_41122,N_42074);
or U43078 (N_43078,N_40447,N_41685);
and U43079 (N_43079,N_40053,N_42367);
xnor U43080 (N_43080,N_41710,N_40194);
xnor U43081 (N_43081,N_41946,N_40529);
nand U43082 (N_43082,N_40000,N_41080);
nand U43083 (N_43083,N_40960,N_41253);
nor U43084 (N_43084,N_42470,N_41151);
or U43085 (N_43085,N_42395,N_41182);
nor U43086 (N_43086,N_41485,N_42478);
xor U43087 (N_43087,N_40312,N_41464);
xnor U43088 (N_43088,N_41062,N_40639);
or U43089 (N_43089,N_42435,N_41835);
and U43090 (N_43090,N_41257,N_41220);
or U43091 (N_43091,N_41382,N_41922);
nor U43092 (N_43092,N_41460,N_40500);
xnor U43093 (N_43093,N_41048,N_42028);
and U43094 (N_43094,N_41217,N_41553);
or U43095 (N_43095,N_40677,N_40120);
xor U43096 (N_43096,N_40515,N_40142);
or U43097 (N_43097,N_40718,N_42119);
xnor U43098 (N_43098,N_40434,N_41035);
nor U43099 (N_43099,N_42069,N_41769);
or U43100 (N_43100,N_41293,N_40636);
and U43101 (N_43101,N_41576,N_42013);
nand U43102 (N_43102,N_42375,N_40291);
and U43103 (N_43103,N_41441,N_42199);
nor U43104 (N_43104,N_42243,N_40658);
xnor U43105 (N_43105,N_40183,N_40069);
and U43106 (N_43106,N_40574,N_40499);
xnor U43107 (N_43107,N_40871,N_42030);
nand U43108 (N_43108,N_40196,N_42444);
nand U43109 (N_43109,N_41574,N_41861);
nor U43110 (N_43110,N_40263,N_40874);
xor U43111 (N_43111,N_42036,N_41405);
or U43112 (N_43112,N_41700,N_42212);
nand U43113 (N_43113,N_41105,N_40030);
xnor U43114 (N_43114,N_40103,N_40634);
or U43115 (N_43115,N_40638,N_40007);
xor U43116 (N_43116,N_40173,N_41593);
and U43117 (N_43117,N_42152,N_40979);
nor U43118 (N_43118,N_41291,N_40167);
xor U43119 (N_43119,N_42203,N_40163);
or U43120 (N_43120,N_40265,N_42056);
nor U43121 (N_43121,N_41552,N_42293);
or U43122 (N_43122,N_41083,N_42272);
or U43123 (N_43123,N_42254,N_42195);
xnor U43124 (N_43124,N_42330,N_40719);
nand U43125 (N_43125,N_40486,N_40017);
and U43126 (N_43126,N_40694,N_40440);
nor U43127 (N_43127,N_42142,N_42475);
or U43128 (N_43128,N_41929,N_40110);
nand U43129 (N_43129,N_42370,N_40726);
or U43130 (N_43130,N_40453,N_42240);
and U43131 (N_43131,N_41425,N_41424);
xnor U43132 (N_43132,N_41123,N_40897);
nor U43133 (N_43133,N_42207,N_42297);
nand U43134 (N_43134,N_41855,N_40773);
xnor U43135 (N_43135,N_40179,N_41396);
nand U43136 (N_43136,N_40790,N_40394);
nand U43137 (N_43137,N_40733,N_41743);
nor U43138 (N_43138,N_41740,N_40073);
nor U43139 (N_43139,N_41970,N_42390);
xnor U43140 (N_43140,N_42282,N_41796);
xor U43141 (N_43141,N_41068,N_41313);
xnor U43142 (N_43142,N_41580,N_40756);
xor U43143 (N_43143,N_42464,N_40074);
nor U43144 (N_43144,N_40342,N_41567);
xor U43145 (N_43145,N_40822,N_40998);
nor U43146 (N_43146,N_40361,N_41248);
or U43147 (N_43147,N_40771,N_40759);
nand U43148 (N_43148,N_40151,N_40009);
nand U43149 (N_43149,N_40350,N_41130);
xnor U43150 (N_43150,N_41197,N_40950);
nor U43151 (N_43151,N_42099,N_42050);
or U43152 (N_43152,N_40336,N_40772);
or U43153 (N_43153,N_41824,N_40199);
nand U43154 (N_43154,N_41702,N_40520);
nand U43155 (N_43155,N_40984,N_42236);
nand U43156 (N_43156,N_40938,N_40390);
nand U43157 (N_43157,N_40105,N_41204);
xor U43158 (N_43158,N_40743,N_41967);
nor U43159 (N_43159,N_40547,N_41088);
nand U43160 (N_43160,N_40223,N_41745);
and U43161 (N_43161,N_41242,N_41826);
and U43162 (N_43162,N_42365,N_41706);
or U43163 (N_43163,N_40926,N_40437);
and U43164 (N_43164,N_42238,N_40039);
and U43165 (N_43165,N_41870,N_41726);
or U43166 (N_43166,N_41840,N_40909);
and U43167 (N_43167,N_41264,N_40345);
and U43168 (N_43168,N_41678,N_40631);
nand U43169 (N_43169,N_41643,N_40755);
or U43170 (N_43170,N_40371,N_42077);
nor U43171 (N_43171,N_42429,N_40384);
nor U43172 (N_43172,N_41286,N_41924);
or U43173 (N_43173,N_41075,N_40059);
or U43174 (N_43174,N_41380,N_41828);
xnor U43175 (N_43175,N_42128,N_41324);
nand U43176 (N_43176,N_40205,N_41190);
nand U43177 (N_43177,N_42014,N_40331);
and U43178 (N_43178,N_41905,N_40833);
and U43179 (N_43179,N_40696,N_40260);
xor U43180 (N_43180,N_41143,N_40632);
nand U43181 (N_43181,N_40270,N_40767);
nor U43182 (N_43182,N_40513,N_42222);
or U43183 (N_43183,N_41273,N_41045);
and U43184 (N_43184,N_40293,N_41381);
or U43185 (N_43185,N_41780,N_40917);
nor U43186 (N_43186,N_41654,N_41569);
and U43187 (N_43187,N_40920,N_40107);
or U43188 (N_43188,N_41235,N_41942);
xnor U43189 (N_43189,N_40019,N_41107);
nand U43190 (N_43190,N_41241,N_42034);
nor U43191 (N_43191,N_40295,N_42421);
nand U43192 (N_43192,N_41069,N_41625);
nand U43193 (N_43193,N_41609,N_41792);
or U43194 (N_43194,N_41776,N_42360);
xor U43195 (N_43195,N_42281,N_40157);
or U43196 (N_43196,N_40470,N_41867);
or U43197 (N_43197,N_42397,N_42167);
nor U43198 (N_43198,N_41586,N_40041);
and U43199 (N_43199,N_40100,N_41583);
nor U43200 (N_43200,N_41283,N_41985);
and U43201 (N_43201,N_41568,N_40466);
nor U43202 (N_43202,N_41652,N_41092);
and U43203 (N_43203,N_42373,N_40842);
xor U43204 (N_43204,N_41124,N_40622);
xor U43205 (N_43205,N_42344,N_40015);
nand U43206 (N_43206,N_40479,N_41019);
or U43207 (N_43207,N_40827,N_40668);
nand U43208 (N_43208,N_41765,N_40365);
and U43209 (N_43209,N_40518,N_41981);
nor U43210 (N_43210,N_40784,N_40379);
xor U43211 (N_43211,N_41516,N_42329);
nor U43212 (N_43212,N_40681,N_40980);
nand U43213 (N_43213,N_42332,N_41665);
and U43214 (N_43214,N_40423,N_42401);
nor U43215 (N_43215,N_40217,N_40063);
nor U43216 (N_43216,N_42070,N_42244);
and U43217 (N_43217,N_40749,N_40415);
xor U43218 (N_43218,N_41880,N_40612);
or U43219 (N_43219,N_41996,N_40212);
xor U43220 (N_43220,N_40165,N_40349);
nand U43221 (N_43221,N_40680,N_42347);
xnor U43222 (N_43222,N_41467,N_41003);
nand U43223 (N_43223,N_40081,N_40481);
nand U43224 (N_43224,N_41656,N_40261);
nand U43225 (N_43225,N_41059,N_41018);
and U43226 (N_43226,N_40228,N_41630);
xor U43227 (N_43227,N_40828,N_40868);
and U43228 (N_43228,N_42175,N_40573);
nand U43229 (N_43229,N_40420,N_41316);
xor U43230 (N_43230,N_41951,N_40299);
nand U43231 (N_43231,N_41471,N_41303);
nand U43232 (N_43232,N_41421,N_40351);
xnor U43233 (N_43233,N_41606,N_40439);
and U43234 (N_43234,N_41157,N_41216);
nor U43235 (N_43235,N_41539,N_41132);
and U43236 (N_43236,N_42100,N_41119);
nand U43237 (N_43237,N_40906,N_41701);
nand U43238 (N_43238,N_41159,N_40360);
nand U43239 (N_43239,N_42448,N_41416);
nor U43240 (N_43240,N_42085,N_41348);
or U43241 (N_43241,N_42093,N_41842);
nor U43242 (N_43242,N_41628,N_40294);
nor U43243 (N_43243,N_40654,N_41305);
nand U43244 (N_43244,N_40602,N_40664);
xnor U43245 (N_43245,N_40918,N_41155);
nor U43246 (N_43246,N_41816,N_41221);
nor U43247 (N_43247,N_40567,N_41767);
and U43248 (N_43248,N_41488,N_41459);
nor U43249 (N_43249,N_40131,N_42193);
or U43250 (N_43250,N_42136,N_42262);
or U43251 (N_43251,N_42346,N_41470);
nor U43252 (N_43252,N_40385,N_41844);
and U43253 (N_43253,N_40175,N_41807);
xor U43254 (N_43254,N_42230,N_40647);
and U43255 (N_43255,N_41476,N_41747);
and U43256 (N_43256,N_40744,N_41589);
and U43257 (N_43257,N_41532,N_41461);
nor U43258 (N_43258,N_40049,N_41499);
or U43259 (N_43259,N_40572,N_40158);
or U43260 (N_43260,N_41811,N_41366);
or U43261 (N_43261,N_41370,N_40033);
or U43262 (N_43262,N_41921,N_41433);
or U43263 (N_43263,N_40066,N_40763);
or U43264 (N_43264,N_40794,N_40619);
and U43265 (N_43265,N_41384,N_41289);
or U43266 (N_43266,N_41333,N_41809);
nor U43267 (N_43267,N_41480,N_42197);
and U43268 (N_43268,N_40605,N_42057);
nand U43269 (N_43269,N_41622,N_42374);
or U43270 (N_43270,N_41672,N_41473);
nor U43271 (N_43271,N_40801,N_40448);
and U43272 (N_43272,N_40020,N_42471);
xnor U43273 (N_43273,N_41831,N_40691);
nand U43274 (N_43274,N_41505,N_42045);
or U43275 (N_43275,N_41506,N_40450);
nand U43276 (N_43276,N_41211,N_41310);
nand U43277 (N_43277,N_40704,N_41162);
xnor U43278 (N_43278,N_40678,N_40366);
nand U43279 (N_43279,N_41517,N_41834);
or U43280 (N_43280,N_40181,N_41427);
xnor U43281 (N_43281,N_42217,N_42280);
nand U43282 (N_43282,N_40104,N_41629);
nor U43283 (N_43283,N_40252,N_41072);
and U43284 (N_43284,N_41437,N_41601);
nand U43285 (N_43285,N_42402,N_42242);
or U43286 (N_43286,N_40935,N_40925);
xor U43287 (N_43287,N_40126,N_42041);
xor U43288 (N_43288,N_41077,N_40497);
or U43289 (N_43289,N_40913,N_40456);
and U43290 (N_43290,N_41044,N_41016);
nand U43291 (N_43291,N_42451,N_42486);
and U43292 (N_43292,N_40930,N_42400);
nor U43293 (N_43293,N_41528,N_40747);
nand U43294 (N_43294,N_42095,N_42352);
and U43295 (N_43295,N_41200,N_40457);
nand U43296 (N_43296,N_40954,N_40826);
nand U43297 (N_43297,N_42088,N_40662);
xor U43298 (N_43298,N_40348,N_40429);
or U43299 (N_43299,N_40514,N_40269);
xor U43300 (N_43300,N_40648,N_40428);
nand U43301 (N_43301,N_40690,N_40002);
nor U43302 (N_43302,N_40460,N_40835);
nor U43303 (N_43303,N_40115,N_42011);
and U43304 (N_43304,N_41901,N_40899);
nand U43305 (N_43305,N_42267,N_41501);
nor U43306 (N_43306,N_40218,N_41353);
xnor U43307 (N_43307,N_40174,N_42202);
xnor U43308 (N_43308,N_40355,N_40111);
and U43309 (N_43309,N_41668,N_40391);
and U43310 (N_43310,N_41859,N_42391);
xor U43311 (N_43311,N_41879,N_40477);
or U43312 (N_43312,N_42366,N_40082);
and U43313 (N_43313,N_41329,N_41695);
or U43314 (N_43314,N_40357,N_41350);
xor U43315 (N_43315,N_42285,N_42310);
and U43316 (N_43316,N_41013,N_41346);
nand U43317 (N_43317,N_40888,N_41094);
nand U43318 (N_43318,N_40044,N_40652);
nand U43319 (N_43319,N_40528,N_42291);
or U43320 (N_43320,N_40043,N_42420);
nor U43321 (N_43321,N_42482,N_41885);
or U43322 (N_43322,N_41650,N_40721);
and U43323 (N_43323,N_42049,N_40285);
xor U43324 (N_43324,N_41444,N_41363);
xnor U43325 (N_43325,N_41934,N_40611);
or U43326 (N_43326,N_40356,N_40959);
xor U43327 (N_43327,N_41198,N_41931);
and U43328 (N_43328,N_40465,N_41360);
or U43329 (N_43329,N_41851,N_40770);
xor U43330 (N_43330,N_42356,N_41219);
or U43331 (N_43331,N_42466,N_40080);
or U43332 (N_43332,N_41783,N_41165);
or U43333 (N_43333,N_40323,N_41983);
nor U43334 (N_43334,N_41932,N_41295);
and U43335 (N_43335,N_41270,N_41730);
nand U43336 (N_43336,N_40136,N_41315);
and U43337 (N_43337,N_40014,N_40273);
or U43338 (N_43338,N_40171,N_40886);
nor U43339 (N_43339,N_41142,N_41387);
nand U43340 (N_43340,N_41029,N_41989);
xnor U43341 (N_43341,N_41193,N_40578);
xor U43342 (N_43342,N_41604,N_41327);
nand U43343 (N_43343,N_41354,N_42061);
and U43344 (N_43344,N_40121,N_42350);
nor U43345 (N_43345,N_41515,N_42237);
and U43346 (N_43346,N_41541,N_41268);
xnor U43347 (N_43347,N_40687,N_40817);
nand U43348 (N_43348,N_40005,N_40671);
nor U43349 (N_43349,N_40714,N_40549);
xor U43350 (N_43350,N_40242,N_41352);
xnor U43351 (N_43351,N_40688,N_40067);
nand U43352 (N_43352,N_41043,N_40713);
nor U43353 (N_43353,N_41588,N_41038);
or U43354 (N_43354,N_42031,N_42462);
and U43355 (N_43355,N_40358,N_40172);
nand U43356 (N_43356,N_42408,N_40278);
and U43357 (N_43357,N_41065,N_41823);
nand U43358 (N_43358,N_41930,N_42328);
and U43359 (N_43359,N_41760,N_41742);
xnor U43360 (N_43360,N_40087,N_41689);
nand U43361 (N_43361,N_40933,N_40283);
and U43362 (N_43362,N_42270,N_41734);
nand U43363 (N_43363,N_41523,N_41141);
nand U43364 (N_43364,N_42415,N_42029);
nand U43365 (N_43365,N_41205,N_41982);
nand U43366 (N_43366,N_40296,N_40731);
nand U43367 (N_43367,N_42403,N_41964);
nand U43368 (N_43368,N_40398,N_41563);
nor U43369 (N_43369,N_40659,N_42015);
or U43370 (N_43370,N_40568,N_40146);
and U43371 (N_43371,N_40953,N_40845);
or U43372 (N_43372,N_41079,N_41462);
and U43373 (N_43373,N_42432,N_40642);
or U43374 (N_43374,N_41508,N_40857);
nor U43375 (N_43375,N_40341,N_40737);
nand U43376 (N_43376,N_40579,N_40319);
nor U43377 (N_43377,N_40058,N_40431);
nand U43378 (N_43378,N_40970,N_42026);
nor U43379 (N_43379,N_40517,N_42138);
and U43380 (N_43380,N_42436,N_40627);
nor U43381 (N_43381,N_42166,N_41301);
or U43382 (N_43382,N_40025,N_41109);
nor U43383 (N_43383,N_42386,N_41832);
nor U43384 (N_43384,N_41125,N_42369);
nand U43385 (N_43385,N_40851,N_40443);
nand U43386 (N_43386,N_41326,N_41978);
or U43387 (N_43387,N_40219,N_41986);
xor U43388 (N_43388,N_42140,N_42455);
and U43389 (N_43389,N_40650,N_42179);
xor U43390 (N_43390,N_41716,N_42458);
and U43391 (N_43391,N_41449,N_41738);
or U43392 (N_43392,N_41118,N_42364);
and U43393 (N_43393,N_40503,N_41209);
nand U43394 (N_43394,N_40711,N_41889);
and U43395 (N_43395,N_40206,N_41171);
xnor U43396 (N_43396,N_40571,N_40628);
nor U43397 (N_43397,N_41288,N_41394);
nor U43398 (N_43398,N_41452,N_40256);
or U43399 (N_43399,N_41106,N_41863);
xor U43400 (N_43400,N_42083,N_41585);
nand U43401 (N_43401,N_40427,N_40198);
and U43402 (N_43402,N_41633,N_41337);
nand U43403 (N_43403,N_41428,N_41139);
and U43404 (N_43404,N_41579,N_41540);
and U43405 (N_43405,N_41213,N_41287);
and U43406 (N_43406,N_41868,N_41873);
and U43407 (N_43407,N_41176,N_42054);
xnor U43408 (N_43408,N_40343,N_40305);
nand U43409 (N_43409,N_42158,N_40484);
nor U43410 (N_43410,N_40985,N_40226);
or U43411 (N_43411,N_42303,N_41178);
nand U43412 (N_43412,N_41667,N_40277);
and U43413 (N_43413,N_41624,N_42127);
and U43414 (N_43414,N_40596,N_41071);
or U43415 (N_43415,N_41214,N_40344);
nor U43416 (N_43416,N_40311,N_41820);
nand U43417 (N_43417,N_40308,N_41292);
or U43418 (N_43418,N_41752,N_42048);
nor U43419 (N_43419,N_42170,N_41199);
nand U43420 (N_43420,N_42066,N_41779);
or U43421 (N_43421,N_42479,N_40337);
nand U43422 (N_43422,N_42447,N_40922);
nand U43423 (N_43423,N_40684,N_41789);
xor U43424 (N_43424,N_40425,N_42052);
nand U43425 (N_43425,N_40699,N_40003);
nor U43426 (N_43426,N_40608,N_40297);
or U43427 (N_43427,N_40403,N_40216);
xor U43428 (N_43428,N_41095,N_41279);
xnor U43429 (N_43429,N_40317,N_41603);
or U43430 (N_43430,N_41594,N_42067);
and U43431 (N_43431,N_40554,N_40685);
nand U43432 (N_43432,N_40412,N_41266);
xnor U43433 (N_43433,N_41202,N_41367);
nor U43434 (N_43434,N_40799,N_40949);
and U43435 (N_43435,N_42414,N_40739);
and U43436 (N_43436,N_41341,N_40679);
xor U43437 (N_43437,N_40854,N_40807);
nor U43438 (N_43438,N_41838,N_41571);
xor U43439 (N_43439,N_41968,N_42341);
nor U43440 (N_43440,N_40872,N_41349);
and U43441 (N_43441,N_40354,N_41925);
nand U43442 (N_43442,N_40161,N_40904);
nand U43443 (N_43443,N_40720,N_40051);
nor U43444 (N_43444,N_40789,N_40562);
or U43445 (N_43445,N_40128,N_41877);
nand U43446 (N_43446,N_42003,N_40266);
or U43447 (N_43447,N_40698,N_40802);
and U43448 (N_43448,N_41435,N_40593);
xor U43449 (N_43449,N_42010,N_40546);
or U43450 (N_43450,N_40795,N_42139);
nand U43451 (N_43451,N_40531,N_40072);
xor U43452 (N_43452,N_40575,N_41788);
nor U43453 (N_43453,N_40201,N_40203);
nand U43454 (N_43454,N_41519,N_42264);
xnor U43455 (N_43455,N_41522,N_42018);
or U43456 (N_43456,N_42261,N_42122);
nor U43457 (N_43457,N_41728,N_41595);
or U43458 (N_43458,N_42223,N_40193);
or U43459 (N_43459,N_41104,N_40660);
and U43460 (N_43460,N_40207,N_41599);
xnor U43461 (N_43461,N_41376,N_40644);
nand U43462 (N_43462,N_42124,N_41957);
or U43463 (N_43463,N_41238,N_40150);
nor U43464 (N_43464,N_41944,N_41777);
nand U43465 (N_43465,N_41388,N_42361);
nand U43466 (N_43466,N_41535,N_40995);
or U43467 (N_43467,N_40090,N_41466);
xnor U43468 (N_43468,N_40527,N_42405);
nor U43469 (N_43469,N_42357,N_42488);
and U43470 (N_43470,N_41082,N_40280);
xnor U43471 (N_43471,N_40545,N_40099);
nand U43472 (N_43472,N_41503,N_41051);
and U43473 (N_43473,N_41023,N_40532);
or U43474 (N_43474,N_40752,N_40892);
nand U43475 (N_43475,N_41854,N_42246);
nand U43476 (N_43476,N_42463,N_42459);
nor U43477 (N_43477,N_41417,N_40359);
nand U43478 (N_43478,N_40083,N_42416);
nand U43479 (N_43479,N_41953,N_40792);
or U43480 (N_43480,N_41736,N_42404);
or U43481 (N_43481,N_40957,N_41031);
and U43482 (N_43482,N_40023,N_42290);
xnor U43483 (N_43483,N_40147,N_40224);
and U43484 (N_43484,N_40188,N_42314);
or U43485 (N_43485,N_42425,N_40239);
or U43486 (N_43486,N_42323,N_41347);
or U43487 (N_43487,N_42413,N_40490);
or U43488 (N_43488,N_41014,N_40735);
nor U43489 (N_43489,N_40276,N_42160);
or U43490 (N_43490,N_40267,N_41979);
or U43491 (N_43491,N_41611,N_40967);
xnor U43492 (N_43492,N_42137,N_40452);
xnor U43493 (N_43493,N_40018,N_40969);
xnor U43494 (N_43494,N_41546,N_41339);
xor U43495 (N_43495,N_40757,N_40521);
nand U43496 (N_43496,N_41487,N_40006);
nor U43497 (N_43497,N_40353,N_40552);
and U43498 (N_43498,N_42162,N_41040);
xnor U43499 (N_43499,N_40716,N_40084);
nor U43500 (N_43500,N_42269,N_40085);
and U43501 (N_43501,N_41181,N_40281);
xor U43502 (N_43502,N_40413,N_42213);
nor U43503 (N_43503,N_40725,N_41430);
nor U43504 (N_43504,N_40060,N_40934);
nor U43505 (N_43505,N_40318,N_41941);
and U43506 (N_43506,N_41314,N_40709);
nor U43507 (N_43507,N_41336,N_42210);
nand U43508 (N_43508,N_40779,N_42123);
and U43509 (N_43509,N_42001,N_42221);
nor U43510 (N_43510,N_40113,N_41987);
nand U43511 (N_43511,N_41096,N_41913);
xor U43512 (N_43512,N_41262,N_41744);
or U43513 (N_43513,N_41977,N_42023);
nor U43514 (N_43514,N_41897,N_42457);
and U43515 (N_43515,N_40507,N_42440);
or U43516 (N_43516,N_40143,N_41693);
xnor U43517 (N_43517,N_41025,N_40867);
and U43518 (N_43518,N_41561,N_41969);
xor U43519 (N_43519,N_41230,N_41064);
xor U43520 (N_43520,N_41443,N_41039);
or U43521 (N_43521,N_42268,N_41948);
xnor U43522 (N_43522,N_42098,N_41839);
nand U43523 (N_43523,N_42319,N_42286);
nand U43524 (N_43524,N_41818,N_40476);
or U43525 (N_43525,N_42363,N_42163);
nor U43526 (N_43526,N_40643,N_41406);
and U43527 (N_43527,N_41409,N_41127);
nand U43528 (N_43528,N_40962,N_41646);
or U43529 (N_43529,N_40282,N_40495);
and U43530 (N_43530,N_42208,N_41351);
nor U43531 (N_43531,N_42468,N_42326);
or U43532 (N_43532,N_40635,N_40641);
nor U43533 (N_43533,N_40374,N_41866);
nand U43534 (N_43534,N_41403,N_40630);
nand U43535 (N_43535,N_40392,N_40222);
xor U43536 (N_43536,N_40075,N_40095);
xor U43537 (N_43537,N_41616,N_41825);
and U43538 (N_43538,N_41719,N_40945);
xnor U43539 (N_43539,N_41680,N_40785);
nor U43540 (N_43540,N_41524,N_40408);
xor U43541 (N_43541,N_40715,N_41150);
xor U43542 (N_43542,N_41325,N_41518);
and U43543 (N_43543,N_40418,N_42327);
nand U43544 (N_43544,N_41914,N_41400);
or U43545 (N_43545,N_40079,N_41058);
xor U43546 (N_43546,N_42450,N_40096);
xor U43547 (N_43547,N_42445,N_41647);
nor U43548 (N_43548,N_40139,N_41781);
nor U43549 (N_43549,N_42339,N_42219);
nor U43550 (N_43550,N_42288,N_40880);
nand U43551 (N_43551,N_42493,N_41790);
nor U43552 (N_43552,N_41896,N_41439);
nor U43553 (N_43553,N_41558,N_41751);
xor U43554 (N_43554,N_42424,N_40505);
nor U43555 (N_43555,N_40187,N_40287);
and U43556 (N_43556,N_40885,N_41527);
nor U43557 (N_43557,N_42016,N_42418);
nand U43558 (N_43558,N_40829,N_41947);
or U43559 (N_43559,N_40825,N_42169);
or U43560 (N_43560,N_41999,N_41636);
nand U43561 (N_43561,N_40491,N_40594);
nand U43562 (N_43562,N_40258,N_40097);
nor U43563 (N_43563,N_40824,N_41415);
nand U43564 (N_43564,N_41682,N_41263);
or U43565 (N_43565,N_41203,N_42192);
xnor U43566 (N_43566,N_40583,N_41146);
nand U43567 (N_43567,N_40855,N_42316);
and U43568 (N_43568,N_41419,N_41167);
nand U43569 (N_43569,N_41423,N_40993);
and U43570 (N_43570,N_41639,N_42324);
xnor U43571 (N_43571,N_41229,N_42183);
nand U43572 (N_43572,N_40388,N_40380);
xnor U43573 (N_43573,N_40098,N_42181);
nor U43574 (N_43574,N_41871,N_40553);
nor U43575 (N_43575,N_42387,N_41577);
xor U43576 (N_43576,N_41278,N_41249);
or U43577 (N_43577,N_40236,N_42007);
nand U43578 (N_43578,N_41169,N_41631);
xor U43579 (N_43579,N_42407,N_40862);
nor U43580 (N_43580,N_40237,N_42368);
nand U43581 (N_43581,N_40062,N_41974);
nand U43582 (N_43582,N_42255,N_41017);
xnor U43583 (N_43583,N_41597,N_40487);
xor U43584 (N_43584,N_40328,N_42107);
and U43585 (N_43585,N_41128,N_40463);
nand U43586 (N_43586,N_40204,N_41422);
xnor U43587 (N_43587,N_40832,N_41121);
or U43588 (N_43588,N_40598,N_41649);
xnor U43589 (N_43589,N_41345,N_40525);
xor U43590 (N_43590,N_40861,N_40931);
xnor U43591 (N_43591,N_40803,N_40210);
nand U43592 (N_43592,N_40912,N_42333);
xnor U43593 (N_43593,N_40901,N_40914);
or U43594 (N_43594,N_41050,N_41129);
nor U43595 (N_43595,N_40853,N_41302);
xnor U43596 (N_43596,N_40697,N_41110);
and U43597 (N_43597,N_41737,N_42178);
and U43598 (N_43598,N_40887,N_42315);
nor U43599 (N_43599,N_41434,N_40054);
or U43600 (N_43600,N_42073,N_41033);
nor U43601 (N_43601,N_42084,N_40321);
or U43602 (N_43602,N_42022,N_40996);
nand U43603 (N_43603,N_41923,N_40838);
or U43604 (N_43604,N_40556,N_41164);
nor U43605 (N_43605,N_42060,N_40368);
and U43606 (N_43606,N_40191,N_41294);
nand U43607 (N_43607,N_40986,N_42000);
nor U43608 (N_43608,N_41637,N_41297);
nor U43609 (N_43609,N_40972,N_40940);
nand U43610 (N_43610,N_41900,N_41137);
xnor U43611 (N_43611,N_40894,N_40646);
or U43612 (N_43612,N_40865,N_42104);
nor U43613 (N_43613,N_40426,N_41240);
nand U43614 (N_43614,N_42495,N_40244);
nor U43615 (N_43615,N_41904,N_41161);
nor U43616 (N_43616,N_40441,N_40787);
and U43617 (N_43617,N_41537,N_41995);
xnor U43618 (N_43618,N_42201,N_40399);
xnor U43619 (N_43619,N_41397,N_40560);
nor U43620 (N_43620,N_42147,N_41308);
nand U43621 (N_43621,N_41529,N_41212);
nand U43622 (N_43622,N_41955,N_41803);
or U43623 (N_43623,N_41474,N_40177);
and U43624 (N_43624,N_41426,N_40896);
nor U43625 (N_43625,N_41340,N_41525);
nor U43626 (N_43626,N_41195,N_40988);
nor U43627 (N_43627,N_42433,N_40093);
nand U43628 (N_43628,N_40234,N_40975);
and U43629 (N_43629,N_40856,N_42094);
or U43630 (N_43630,N_41991,N_40987);
and U43631 (N_43631,N_41010,N_41554);
xor U43632 (N_43632,N_40122,N_41385);
and U43633 (N_43633,N_41361,N_40616);
xor U43634 (N_43634,N_41237,N_41267);
nand U43635 (N_43635,N_41468,N_40667);
nor U43636 (N_43636,N_41420,N_41255);
xnor U43637 (N_43637,N_40301,N_40001);
and U43638 (N_43638,N_42216,N_42409);
xor U43639 (N_43639,N_40614,N_41322);
or U43640 (N_43640,N_42304,N_42249);
nand U43641 (N_43641,N_41486,N_41492);
nand U43642 (N_43642,N_40315,N_41448);
nand U43643 (N_43643,N_41784,N_41797);
or U43644 (N_43644,N_41113,N_41869);
xor U43645 (N_43645,N_41857,N_40898);
or U43646 (N_43646,N_40184,N_40076);
or U43647 (N_43647,N_41307,N_40274);
and U43648 (N_43648,N_40432,N_42102);
xnor U43649 (N_43649,N_42287,N_41514);
and U43650 (N_43650,N_41046,N_42121);
nor U43651 (N_43651,N_40834,N_41692);
and U43652 (N_43652,N_41757,N_40409);
nor U43653 (N_43653,N_41138,N_42456);
nand U43654 (N_43654,N_41819,N_40208);
xnor U43655 (N_43655,N_41144,N_40106);
or U43656 (N_43656,N_41661,N_41566);
nor U43657 (N_43657,N_41414,N_40303);
nand U43658 (N_43658,N_40471,N_42300);
nand U43659 (N_43659,N_40557,N_41131);
or U43660 (N_43660,N_40907,N_41049);
nand U43661 (N_43661,N_40544,N_40454);
or U43662 (N_43662,N_41782,N_41087);
nand U43663 (N_43663,N_41497,N_41729);
nor U43664 (N_43664,N_41060,N_41004);
xnor U43665 (N_43665,N_41269,N_40424);
or U43666 (N_43666,N_42151,N_42497);
and U43667 (N_43667,N_41940,N_40225);
nand U43668 (N_43668,N_40522,N_40397);
nor U43669 (N_43669,N_41244,N_40264);
xor U43670 (N_43670,N_41393,N_40433);
nand U43671 (N_43671,N_40538,N_40695);
nor U43672 (N_43672,N_40540,N_41697);
or U43673 (N_43673,N_40777,N_40946);
nand U43674 (N_43674,N_40623,N_41404);
or U43675 (N_43675,N_40333,N_42431);
xnor U43676 (N_43676,N_42019,N_40155);
nand U43677 (N_43677,N_41153,N_40469);
xor U43678 (N_43678,N_41277,N_41224);
nand U43679 (N_43679,N_40347,N_40916);
or U43680 (N_43680,N_42225,N_41936);
xor U43681 (N_43681,N_40761,N_41041);
nor U43682 (N_43682,N_41275,N_40858);
xor U43683 (N_43683,N_41600,N_41621);
nor U43684 (N_43684,N_41892,N_41590);
or U43685 (N_43685,N_41971,N_40138);
and U43686 (N_43686,N_41954,N_40123);
or U43687 (N_43687,N_40705,N_40109);
and U43688 (N_43688,N_40202,N_42114);
nand U43689 (N_43689,N_40251,N_41526);
and U43690 (N_43690,N_42274,N_40541);
and U43691 (N_43691,N_41735,N_42191);
and U43692 (N_43692,N_42443,N_42091);
or U43693 (N_43693,N_40841,N_42480);
or U43694 (N_43694,N_42336,N_41020);
nand U43695 (N_43695,N_41845,N_40057);
and U43696 (N_43696,N_41052,N_42348);
nor U43697 (N_43697,N_41766,N_41805);
nand U43698 (N_43698,N_40859,N_42157);
xnor U43699 (N_43699,N_41192,N_42200);
nand U43700 (N_43700,N_40035,N_40011);
nor U43701 (N_43701,N_42150,N_40189);
nand U43702 (N_43702,N_42411,N_40414);
nor U43703 (N_43703,N_41618,N_41061);
and U43704 (N_43704,N_41798,N_41619);
nor U43705 (N_43705,N_41357,N_40692);
nand U43706 (N_43706,N_41179,N_40848);
or U43707 (N_43707,N_40141,N_40707);
or U43708 (N_43708,N_40929,N_40166);
xor U43709 (N_43709,N_41174,N_42442);
and U43710 (N_43710,N_40114,N_41687);
nand U43711 (N_43711,N_40919,N_41494);
nand U43712 (N_43712,N_40132,N_40780);
nand U43713 (N_43713,N_40118,N_40927);
nand U43714 (N_43714,N_40870,N_41542);
nor U43715 (N_43715,N_40135,N_42043);
or U43716 (N_43716,N_41282,N_41358);
nand U43717 (N_43717,N_41074,N_40615);
and U43718 (N_43718,N_41115,N_42299);
and U43719 (N_43719,N_42484,N_40310);
nor U43720 (N_43720,N_41371,N_41442);
and U43721 (N_43721,N_40482,N_40982);
nor U43722 (N_43722,N_41632,N_40127);
or U43723 (N_43723,N_42419,N_41615);
or U43724 (N_43724,N_41860,N_40791);
xor U43725 (N_43725,N_42068,N_40112);
xor U43726 (N_43726,N_41091,N_40999);
xor U43727 (N_43727,N_40952,N_41749);
and U43728 (N_43728,N_40724,N_42309);
or U43729 (N_43729,N_41862,N_40302);
or U43730 (N_43730,N_42273,N_41432);
xor U43731 (N_43731,N_41763,N_42047);
and U43732 (N_43732,N_40334,N_40530);
and U43733 (N_43733,N_40363,N_41916);
xnor U43734 (N_43734,N_41911,N_42284);
nand U43735 (N_43735,N_41856,N_40307);
xor U43736 (N_43736,N_41364,N_40788);
and U43737 (N_43737,N_41770,N_41723);
and U43738 (N_43738,N_42283,N_41793);
nand U43739 (N_43739,N_42469,N_40211);
nand U43740 (N_43740,N_41787,N_41495);
or U43741 (N_43741,N_41100,N_42038);
nand U43742 (N_43742,N_42446,N_41815);
xnor U43743 (N_43743,N_41718,N_41772);
nand U43744 (N_43744,N_40176,N_41281);
or U43745 (N_43745,N_40584,N_42227);
or U43746 (N_43746,N_41727,N_42086);
or U43747 (N_43747,N_42461,N_41902);
and U43748 (N_43748,N_40250,N_40382);
xnor U43749 (N_43749,N_40597,N_42355);
nor U43750 (N_43750,N_41030,N_42417);
and U43751 (N_43751,N_42149,N_42056);
xor U43752 (N_43752,N_41662,N_40914);
xnor U43753 (N_43753,N_41137,N_40774);
or U43754 (N_43754,N_42156,N_40118);
nand U43755 (N_43755,N_41684,N_40682);
xnor U43756 (N_43756,N_41261,N_40986);
or U43757 (N_43757,N_41322,N_41292);
and U43758 (N_43758,N_40200,N_41491);
xor U43759 (N_43759,N_40723,N_41245);
and U43760 (N_43760,N_42227,N_42118);
nand U43761 (N_43761,N_40838,N_41254);
or U43762 (N_43762,N_41239,N_41176);
or U43763 (N_43763,N_41531,N_41709);
nand U43764 (N_43764,N_40770,N_42304);
xnor U43765 (N_43765,N_42083,N_40485);
and U43766 (N_43766,N_41658,N_40570);
or U43767 (N_43767,N_40507,N_42079);
and U43768 (N_43768,N_40553,N_41551);
nand U43769 (N_43769,N_41122,N_42418);
nand U43770 (N_43770,N_40284,N_40138);
nand U43771 (N_43771,N_41576,N_41782);
xor U43772 (N_43772,N_40144,N_41961);
nand U43773 (N_43773,N_40093,N_42233);
nand U43774 (N_43774,N_41559,N_41888);
and U43775 (N_43775,N_41917,N_40084);
xnor U43776 (N_43776,N_42491,N_40432);
or U43777 (N_43777,N_41294,N_40065);
and U43778 (N_43778,N_41717,N_40157);
nor U43779 (N_43779,N_41508,N_40636);
nand U43780 (N_43780,N_40918,N_42497);
nor U43781 (N_43781,N_40219,N_40500);
nand U43782 (N_43782,N_41733,N_40676);
or U43783 (N_43783,N_41451,N_42268);
or U43784 (N_43784,N_40444,N_40496);
nand U43785 (N_43785,N_40536,N_41612);
nand U43786 (N_43786,N_40959,N_40921);
nor U43787 (N_43787,N_40661,N_40061);
xnor U43788 (N_43788,N_41527,N_41294);
nand U43789 (N_43789,N_40717,N_40613);
nand U43790 (N_43790,N_42048,N_40864);
and U43791 (N_43791,N_40757,N_40948);
nor U43792 (N_43792,N_42454,N_41049);
xnor U43793 (N_43793,N_40178,N_42043);
nand U43794 (N_43794,N_42264,N_42450);
and U43795 (N_43795,N_40650,N_40531);
or U43796 (N_43796,N_40666,N_40731);
nor U43797 (N_43797,N_40620,N_41826);
and U43798 (N_43798,N_40624,N_40096);
xnor U43799 (N_43799,N_40559,N_42085);
nand U43800 (N_43800,N_41634,N_40680);
nand U43801 (N_43801,N_40766,N_42286);
nand U43802 (N_43802,N_40091,N_40680);
xnor U43803 (N_43803,N_40858,N_41051);
or U43804 (N_43804,N_40552,N_42063);
and U43805 (N_43805,N_40434,N_41286);
and U43806 (N_43806,N_41742,N_40907);
and U43807 (N_43807,N_40651,N_42335);
and U43808 (N_43808,N_40639,N_40822);
nor U43809 (N_43809,N_42187,N_41231);
nand U43810 (N_43810,N_41915,N_40661);
nor U43811 (N_43811,N_41207,N_40016);
or U43812 (N_43812,N_41332,N_41988);
nor U43813 (N_43813,N_42274,N_41124);
and U43814 (N_43814,N_41144,N_40065);
nand U43815 (N_43815,N_42442,N_41955);
and U43816 (N_43816,N_41973,N_41756);
nand U43817 (N_43817,N_40475,N_41099);
and U43818 (N_43818,N_41862,N_42431);
xor U43819 (N_43819,N_41311,N_41395);
nor U43820 (N_43820,N_42400,N_40005);
nand U43821 (N_43821,N_40926,N_40616);
nor U43822 (N_43822,N_41696,N_40702);
and U43823 (N_43823,N_40819,N_40822);
and U43824 (N_43824,N_41071,N_41722);
and U43825 (N_43825,N_40626,N_41066);
or U43826 (N_43826,N_40467,N_40390);
nor U43827 (N_43827,N_41857,N_42177);
and U43828 (N_43828,N_41520,N_42253);
nor U43829 (N_43829,N_40395,N_42194);
and U43830 (N_43830,N_41337,N_41252);
nor U43831 (N_43831,N_40480,N_42269);
and U43832 (N_43832,N_40628,N_41287);
xnor U43833 (N_43833,N_42008,N_41264);
nor U43834 (N_43834,N_42057,N_42378);
nand U43835 (N_43835,N_41219,N_40419);
nor U43836 (N_43836,N_40951,N_40969);
nor U43837 (N_43837,N_40658,N_40560);
nor U43838 (N_43838,N_42041,N_41571);
xnor U43839 (N_43839,N_40802,N_41057);
nand U43840 (N_43840,N_42338,N_40197);
and U43841 (N_43841,N_41763,N_42153);
nand U43842 (N_43842,N_40049,N_40690);
or U43843 (N_43843,N_41180,N_40073);
nor U43844 (N_43844,N_41014,N_40718);
nor U43845 (N_43845,N_41435,N_41325);
or U43846 (N_43846,N_41690,N_40911);
xnor U43847 (N_43847,N_41478,N_41885);
and U43848 (N_43848,N_40006,N_40912);
or U43849 (N_43849,N_41160,N_40252);
nor U43850 (N_43850,N_41388,N_41328);
nor U43851 (N_43851,N_40366,N_41891);
and U43852 (N_43852,N_41933,N_42083);
xor U43853 (N_43853,N_40738,N_40633);
xnor U43854 (N_43854,N_40262,N_41189);
nand U43855 (N_43855,N_40935,N_40791);
xnor U43856 (N_43856,N_40640,N_40844);
or U43857 (N_43857,N_41986,N_40309);
or U43858 (N_43858,N_40820,N_41888);
nand U43859 (N_43859,N_40954,N_41685);
and U43860 (N_43860,N_40597,N_41271);
nand U43861 (N_43861,N_41032,N_42218);
xnor U43862 (N_43862,N_40656,N_40468);
or U43863 (N_43863,N_41124,N_40474);
nand U43864 (N_43864,N_41719,N_42402);
and U43865 (N_43865,N_41829,N_41419);
and U43866 (N_43866,N_40660,N_41876);
or U43867 (N_43867,N_42470,N_41028);
xnor U43868 (N_43868,N_41996,N_40637);
and U43869 (N_43869,N_40007,N_40600);
xnor U43870 (N_43870,N_40467,N_41124);
nand U43871 (N_43871,N_42241,N_41278);
or U43872 (N_43872,N_41818,N_41833);
and U43873 (N_43873,N_40581,N_41804);
xnor U43874 (N_43874,N_42020,N_40150);
nor U43875 (N_43875,N_42281,N_41610);
xor U43876 (N_43876,N_41596,N_41432);
or U43877 (N_43877,N_40940,N_41209);
nand U43878 (N_43878,N_40552,N_41238);
and U43879 (N_43879,N_41649,N_42156);
xor U43880 (N_43880,N_42260,N_42432);
and U43881 (N_43881,N_40016,N_40725);
xnor U43882 (N_43882,N_41632,N_41942);
xor U43883 (N_43883,N_41407,N_42409);
nand U43884 (N_43884,N_41604,N_41681);
nand U43885 (N_43885,N_40782,N_40021);
nor U43886 (N_43886,N_42181,N_41142);
nor U43887 (N_43887,N_41044,N_41472);
nand U43888 (N_43888,N_42029,N_42047);
nand U43889 (N_43889,N_41291,N_41663);
xnor U43890 (N_43890,N_40862,N_40608);
nand U43891 (N_43891,N_40465,N_40409);
and U43892 (N_43892,N_40072,N_40730);
nand U43893 (N_43893,N_41102,N_40781);
xnor U43894 (N_43894,N_41179,N_41262);
and U43895 (N_43895,N_40942,N_42088);
xor U43896 (N_43896,N_41160,N_41852);
nand U43897 (N_43897,N_41548,N_40375);
xor U43898 (N_43898,N_41768,N_40328);
and U43899 (N_43899,N_41519,N_40154);
and U43900 (N_43900,N_41127,N_41310);
nor U43901 (N_43901,N_40408,N_41276);
nor U43902 (N_43902,N_42417,N_41906);
nor U43903 (N_43903,N_40478,N_42303);
nand U43904 (N_43904,N_40729,N_42168);
xnor U43905 (N_43905,N_40807,N_40292);
nand U43906 (N_43906,N_42322,N_41383);
and U43907 (N_43907,N_41934,N_42028);
and U43908 (N_43908,N_40867,N_40313);
or U43909 (N_43909,N_41360,N_42434);
xnor U43910 (N_43910,N_40665,N_41098);
or U43911 (N_43911,N_40039,N_41409);
or U43912 (N_43912,N_40783,N_42325);
xnor U43913 (N_43913,N_41182,N_40200);
nand U43914 (N_43914,N_41706,N_41592);
and U43915 (N_43915,N_40805,N_41832);
and U43916 (N_43916,N_41709,N_40686);
xnor U43917 (N_43917,N_40761,N_40279);
xnor U43918 (N_43918,N_42198,N_42259);
and U43919 (N_43919,N_42033,N_41143);
nor U43920 (N_43920,N_41242,N_41245);
nand U43921 (N_43921,N_41371,N_42164);
nand U43922 (N_43922,N_42258,N_40782);
and U43923 (N_43923,N_40337,N_40565);
and U43924 (N_43924,N_40343,N_42426);
and U43925 (N_43925,N_41664,N_41010);
xnor U43926 (N_43926,N_42221,N_41593);
nand U43927 (N_43927,N_41072,N_40171);
nor U43928 (N_43928,N_40531,N_40649);
or U43929 (N_43929,N_41897,N_40004);
and U43930 (N_43930,N_41833,N_41343);
nand U43931 (N_43931,N_40761,N_40466);
and U43932 (N_43932,N_40101,N_42196);
nand U43933 (N_43933,N_41093,N_42306);
xor U43934 (N_43934,N_40566,N_41785);
and U43935 (N_43935,N_40462,N_41663);
nor U43936 (N_43936,N_40887,N_42067);
or U43937 (N_43937,N_40392,N_40685);
nand U43938 (N_43938,N_40909,N_41391);
or U43939 (N_43939,N_40319,N_42070);
or U43940 (N_43940,N_41546,N_40932);
nand U43941 (N_43941,N_41108,N_41900);
nor U43942 (N_43942,N_40845,N_41257);
nor U43943 (N_43943,N_41807,N_40696);
and U43944 (N_43944,N_40615,N_41066);
or U43945 (N_43945,N_40061,N_41150);
and U43946 (N_43946,N_40584,N_41321);
and U43947 (N_43947,N_42133,N_41607);
and U43948 (N_43948,N_42116,N_41254);
and U43949 (N_43949,N_41180,N_40168);
nand U43950 (N_43950,N_42058,N_41018);
nand U43951 (N_43951,N_40809,N_41906);
xor U43952 (N_43952,N_40546,N_40083);
nor U43953 (N_43953,N_41499,N_41399);
and U43954 (N_43954,N_40549,N_42032);
nand U43955 (N_43955,N_40949,N_42435);
and U43956 (N_43956,N_42282,N_40090);
xor U43957 (N_43957,N_41198,N_41582);
xor U43958 (N_43958,N_41879,N_40731);
nor U43959 (N_43959,N_42017,N_41358);
or U43960 (N_43960,N_42087,N_41101);
xor U43961 (N_43961,N_42232,N_42046);
nand U43962 (N_43962,N_41621,N_40586);
xor U43963 (N_43963,N_41205,N_41820);
nor U43964 (N_43964,N_41453,N_41339);
nand U43965 (N_43965,N_41314,N_40765);
xor U43966 (N_43966,N_40706,N_41882);
nand U43967 (N_43967,N_40268,N_40369);
xor U43968 (N_43968,N_42363,N_41894);
nand U43969 (N_43969,N_40246,N_41153);
and U43970 (N_43970,N_41142,N_40205);
nand U43971 (N_43971,N_41224,N_40949);
and U43972 (N_43972,N_41585,N_41363);
or U43973 (N_43973,N_41945,N_40486);
and U43974 (N_43974,N_41322,N_41473);
nor U43975 (N_43975,N_40227,N_41122);
or U43976 (N_43976,N_41640,N_41003);
nand U43977 (N_43977,N_41696,N_41779);
xor U43978 (N_43978,N_41701,N_42116);
nor U43979 (N_43979,N_42147,N_41328);
nand U43980 (N_43980,N_42020,N_41879);
or U43981 (N_43981,N_40973,N_42164);
xor U43982 (N_43982,N_42297,N_42360);
nor U43983 (N_43983,N_40539,N_40032);
nor U43984 (N_43984,N_40528,N_40214);
xor U43985 (N_43985,N_42222,N_41569);
nor U43986 (N_43986,N_40154,N_41755);
nand U43987 (N_43987,N_41753,N_41121);
or U43988 (N_43988,N_41842,N_41670);
nor U43989 (N_43989,N_41471,N_41813);
nor U43990 (N_43990,N_40887,N_40059);
nand U43991 (N_43991,N_42229,N_40755);
and U43992 (N_43992,N_41863,N_40567);
or U43993 (N_43993,N_42317,N_42447);
nor U43994 (N_43994,N_41279,N_40077);
nand U43995 (N_43995,N_40118,N_42242);
and U43996 (N_43996,N_40971,N_41604);
and U43997 (N_43997,N_41859,N_40505);
and U43998 (N_43998,N_42161,N_41317);
nand U43999 (N_43999,N_41809,N_41605);
nand U44000 (N_44000,N_41092,N_40669);
xor U44001 (N_44001,N_41250,N_41866);
nor U44002 (N_44002,N_40189,N_40843);
or U44003 (N_44003,N_40172,N_42277);
nand U44004 (N_44004,N_40686,N_40972);
xor U44005 (N_44005,N_40910,N_40561);
xnor U44006 (N_44006,N_40070,N_41769);
xor U44007 (N_44007,N_41489,N_41874);
xor U44008 (N_44008,N_41740,N_40259);
xnor U44009 (N_44009,N_40099,N_40410);
and U44010 (N_44010,N_40723,N_42142);
and U44011 (N_44011,N_41069,N_40999);
or U44012 (N_44012,N_42203,N_41955);
nand U44013 (N_44013,N_42499,N_41430);
xor U44014 (N_44014,N_42280,N_40686);
nor U44015 (N_44015,N_42029,N_42473);
xor U44016 (N_44016,N_41722,N_40258);
nand U44017 (N_44017,N_41796,N_40532);
or U44018 (N_44018,N_40851,N_41516);
nand U44019 (N_44019,N_40461,N_40694);
and U44020 (N_44020,N_41668,N_42475);
or U44021 (N_44021,N_41733,N_41700);
nor U44022 (N_44022,N_41056,N_41441);
nand U44023 (N_44023,N_41592,N_42352);
or U44024 (N_44024,N_41136,N_40101);
nor U44025 (N_44025,N_40227,N_40337);
or U44026 (N_44026,N_41663,N_41865);
nand U44027 (N_44027,N_41981,N_42432);
xor U44028 (N_44028,N_41993,N_40193);
or U44029 (N_44029,N_40908,N_40316);
or U44030 (N_44030,N_41307,N_41715);
nand U44031 (N_44031,N_41475,N_40203);
xnor U44032 (N_44032,N_40453,N_40682);
nand U44033 (N_44033,N_42474,N_40422);
or U44034 (N_44034,N_40841,N_41834);
and U44035 (N_44035,N_40997,N_40870);
nor U44036 (N_44036,N_40277,N_41978);
nor U44037 (N_44037,N_42213,N_41971);
nor U44038 (N_44038,N_41504,N_40140);
or U44039 (N_44039,N_41185,N_40328);
or U44040 (N_44040,N_41757,N_40297);
xnor U44041 (N_44041,N_41814,N_41129);
or U44042 (N_44042,N_40829,N_40514);
or U44043 (N_44043,N_41131,N_40117);
xnor U44044 (N_44044,N_41484,N_40368);
xor U44045 (N_44045,N_42259,N_40386);
nand U44046 (N_44046,N_40074,N_41537);
xor U44047 (N_44047,N_40927,N_40829);
nand U44048 (N_44048,N_42136,N_41204);
nor U44049 (N_44049,N_41026,N_40551);
nor U44050 (N_44050,N_42048,N_40318);
or U44051 (N_44051,N_40011,N_41088);
and U44052 (N_44052,N_41184,N_40613);
xor U44053 (N_44053,N_42113,N_40597);
and U44054 (N_44054,N_42126,N_40603);
or U44055 (N_44055,N_41581,N_41954);
nand U44056 (N_44056,N_42079,N_42461);
nand U44057 (N_44057,N_40810,N_41599);
nand U44058 (N_44058,N_41002,N_40425);
xnor U44059 (N_44059,N_40923,N_40141);
nor U44060 (N_44060,N_40078,N_42049);
and U44061 (N_44061,N_40393,N_41263);
xor U44062 (N_44062,N_41026,N_40371);
nand U44063 (N_44063,N_41085,N_42292);
xnor U44064 (N_44064,N_41884,N_42439);
nor U44065 (N_44065,N_42040,N_41987);
nor U44066 (N_44066,N_42212,N_41205);
nor U44067 (N_44067,N_40347,N_41288);
nor U44068 (N_44068,N_41670,N_41655);
nand U44069 (N_44069,N_41545,N_40198);
or U44070 (N_44070,N_40783,N_41050);
xor U44071 (N_44071,N_41292,N_40385);
or U44072 (N_44072,N_42029,N_42399);
and U44073 (N_44073,N_40488,N_41436);
xor U44074 (N_44074,N_40979,N_40467);
and U44075 (N_44075,N_40527,N_40798);
and U44076 (N_44076,N_42154,N_41985);
and U44077 (N_44077,N_41399,N_40700);
and U44078 (N_44078,N_42192,N_40786);
or U44079 (N_44079,N_40943,N_40318);
nand U44080 (N_44080,N_40233,N_41053);
and U44081 (N_44081,N_41986,N_42343);
or U44082 (N_44082,N_40306,N_40142);
nor U44083 (N_44083,N_40169,N_41590);
xnor U44084 (N_44084,N_41161,N_40679);
and U44085 (N_44085,N_40407,N_40447);
nor U44086 (N_44086,N_40888,N_40889);
and U44087 (N_44087,N_40389,N_41323);
and U44088 (N_44088,N_41988,N_40886);
xnor U44089 (N_44089,N_41924,N_40833);
nand U44090 (N_44090,N_40971,N_41312);
nand U44091 (N_44091,N_40164,N_41751);
or U44092 (N_44092,N_40882,N_40286);
and U44093 (N_44093,N_42182,N_42210);
and U44094 (N_44094,N_41828,N_41690);
xor U44095 (N_44095,N_40374,N_40185);
and U44096 (N_44096,N_41837,N_41375);
nor U44097 (N_44097,N_40422,N_40903);
or U44098 (N_44098,N_41299,N_42388);
or U44099 (N_44099,N_41763,N_41766);
xnor U44100 (N_44100,N_40969,N_41808);
or U44101 (N_44101,N_41592,N_40601);
xnor U44102 (N_44102,N_42098,N_42168);
or U44103 (N_44103,N_40876,N_41354);
nor U44104 (N_44104,N_41113,N_41083);
xnor U44105 (N_44105,N_41893,N_41710);
and U44106 (N_44106,N_41709,N_41834);
nand U44107 (N_44107,N_41036,N_40518);
nand U44108 (N_44108,N_42336,N_40760);
nor U44109 (N_44109,N_41710,N_41610);
nand U44110 (N_44110,N_41339,N_40163);
xor U44111 (N_44111,N_40174,N_40059);
and U44112 (N_44112,N_41444,N_41445);
xnor U44113 (N_44113,N_42282,N_40314);
nand U44114 (N_44114,N_41897,N_41514);
nand U44115 (N_44115,N_41263,N_40719);
xor U44116 (N_44116,N_40338,N_40582);
nor U44117 (N_44117,N_40909,N_41580);
and U44118 (N_44118,N_41470,N_41800);
xor U44119 (N_44119,N_41392,N_40929);
nor U44120 (N_44120,N_41322,N_42103);
nand U44121 (N_44121,N_40377,N_40953);
and U44122 (N_44122,N_41997,N_40774);
or U44123 (N_44123,N_41060,N_41219);
nor U44124 (N_44124,N_41947,N_40920);
xor U44125 (N_44125,N_41717,N_40554);
or U44126 (N_44126,N_42155,N_40245);
nand U44127 (N_44127,N_40117,N_40512);
and U44128 (N_44128,N_40926,N_41788);
and U44129 (N_44129,N_41284,N_41929);
and U44130 (N_44130,N_41469,N_42208);
nand U44131 (N_44131,N_40290,N_42328);
nand U44132 (N_44132,N_40522,N_42217);
and U44133 (N_44133,N_41821,N_40083);
nand U44134 (N_44134,N_40413,N_42149);
xor U44135 (N_44135,N_41367,N_40718);
xor U44136 (N_44136,N_41948,N_40450);
nor U44137 (N_44137,N_42260,N_40025);
nor U44138 (N_44138,N_41768,N_40543);
nand U44139 (N_44139,N_40606,N_40931);
and U44140 (N_44140,N_41854,N_40775);
or U44141 (N_44141,N_40051,N_42017);
xnor U44142 (N_44142,N_40919,N_42395);
and U44143 (N_44143,N_41582,N_40184);
or U44144 (N_44144,N_40361,N_41600);
xor U44145 (N_44145,N_40701,N_41212);
nand U44146 (N_44146,N_42198,N_41604);
nor U44147 (N_44147,N_42368,N_40193);
or U44148 (N_44148,N_40703,N_40876);
nand U44149 (N_44149,N_42443,N_40296);
or U44150 (N_44150,N_42357,N_42016);
nand U44151 (N_44151,N_41989,N_40717);
and U44152 (N_44152,N_41297,N_40858);
and U44153 (N_44153,N_40829,N_40467);
and U44154 (N_44154,N_40816,N_41950);
nand U44155 (N_44155,N_42091,N_42172);
nand U44156 (N_44156,N_41584,N_41090);
and U44157 (N_44157,N_40109,N_40479);
xor U44158 (N_44158,N_40690,N_40275);
or U44159 (N_44159,N_40874,N_40854);
nor U44160 (N_44160,N_41602,N_41430);
nand U44161 (N_44161,N_41459,N_40918);
xnor U44162 (N_44162,N_41709,N_41350);
nor U44163 (N_44163,N_42282,N_40242);
or U44164 (N_44164,N_41653,N_41661);
xnor U44165 (N_44165,N_40704,N_41385);
or U44166 (N_44166,N_41210,N_41678);
nor U44167 (N_44167,N_40890,N_41898);
nor U44168 (N_44168,N_42044,N_40598);
and U44169 (N_44169,N_41747,N_42439);
xor U44170 (N_44170,N_42139,N_41052);
nor U44171 (N_44171,N_40249,N_41968);
and U44172 (N_44172,N_42463,N_42272);
nand U44173 (N_44173,N_41755,N_40666);
xnor U44174 (N_44174,N_40447,N_41589);
or U44175 (N_44175,N_42048,N_41022);
or U44176 (N_44176,N_41473,N_41695);
or U44177 (N_44177,N_42467,N_41871);
or U44178 (N_44178,N_42398,N_42326);
xnor U44179 (N_44179,N_42003,N_41892);
xnor U44180 (N_44180,N_41800,N_41510);
nand U44181 (N_44181,N_40722,N_40041);
or U44182 (N_44182,N_42203,N_42132);
and U44183 (N_44183,N_42397,N_41405);
nand U44184 (N_44184,N_42193,N_40407);
or U44185 (N_44185,N_41026,N_40571);
xor U44186 (N_44186,N_41418,N_42008);
nand U44187 (N_44187,N_42399,N_42160);
or U44188 (N_44188,N_40359,N_40739);
nand U44189 (N_44189,N_42475,N_40092);
or U44190 (N_44190,N_40760,N_40332);
or U44191 (N_44191,N_41059,N_42340);
or U44192 (N_44192,N_42166,N_41471);
or U44193 (N_44193,N_41389,N_41415);
or U44194 (N_44194,N_41764,N_42050);
and U44195 (N_44195,N_40171,N_40002);
nor U44196 (N_44196,N_40903,N_42102);
nand U44197 (N_44197,N_41901,N_41374);
nor U44198 (N_44198,N_41662,N_40882);
nor U44199 (N_44199,N_41989,N_41942);
or U44200 (N_44200,N_42372,N_40250);
nand U44201 (N_44201,N_42385,N_40009);
xnor U44202 (N_44202,N_40967,N_40233);
nor U44203 (N_44203,N_40732,N_41800);
nor U44204 (N_44204,N_40932,N_40394);
nand U44205 (N_44205,N_41111,N_41043);
nor U44206 (N_44206,N_40856,N_40268);
xnor U44207 (N_44207,N_40729,N_40574);
or U44208 (N_44208,N_41068,N_41065);
nor U44209 (N_44209,N_40734,N_40049);
nor U44210 (N_44210,N_41612,N_41866);
or U44211 (N_44211,N_40426,N_42286);
nor U44212 (N_44212,N_40895,N_41630);
nor U44213 (N_44213,N_40701,N_40097);
xor U44214 (N_44214,N_40880,N_42242);
or U44215 (N_44215,N_42013,N_42220);
and U44216 (N_44216,N_40474,N_41732);
and U44217 (N_44217,N_41791,N_40547);
nor U44218 (N_44218,N_40936,N_42132);
xor U44219 (N_44219,N_41892,N_41157);
xor U44220 (N_44220,N_41060,N_42125);
or U44221 (N_44221,N_40960,N_40549);
nand U44222 (N_44222,N_41635,N_42007);
nor U44223 (N_44223,N_41965,N_40657);
and U44224 (N_44224,N_42298,N_40204);
nand U44225 (N_44225,N_42123,N_40870);
nor U44226 (N_44226,N_40359,N_40517);
xor U44227 (N_44227,N_42029,N_42129);
xnor U44228 (N_44228,N_42484,N_41146);
nand U44229 (N_44229,N_40510,N_42044);
nand U44230 (N_44230,N_41329,N_41884);
or U44231 (N_44231,N_41382,N_42241);
nand U44232 (N_44232,N_40017,N_40532);
and U44233 (N_44233,N_41920,N_40998);
and U44234 (N_44234,N_40780,N_42441);
nor U44235 (N_44235,N_42086,N_40043);
nor U44236 (N_44236,N_41540,N_40697);
nor U44237 (N_44237,N_40909,N_41877);
nor U44238 (N_44238,N_41961,N_40663);
and U44239 (N_44239,N_40377,N_40882);
and U44240 (N_44240,N_42129,N_42058);
xor U44241 (N_44241,N_40871,N_41153);
and U44242 (N_44242,N_40247,N_40444);
xnor U44243 (N_44243,N_42231,N_42489);
nand U44244 (N_44244,N_40615,N_41525);
and U44245 (N_44245,N_41907,N_40664);
or U44246 (N_44246,N_41189,N_41797);
or U44247 (N_44247,N_40240,N_40382);
xnor U44248 (N_44248,N_41944,N_41037);
and U44249 (N_44249,N_41226,N_40641);
and U44250 (N_44250,N_40522,N_41088);
nand U44251 (N_44251,N_41783,N_42452);
and U44252 (N_44252,N_40260,N_41012);
or U44253 (N_44253,N_42323,N_41057);
nand U44254 (N_44254,N_40076,N_40737);
nand U44255 (N_44255,N_42264,N_40222);
nand U44256 (N_44256,N_40244,N_40634);
and U44257 (N_44257,N_42188,N_41216);
and U44258 (N_44258,N_41260,N_42334);
nor U44259 (N_44259,N_40331,N_40749);
nand U44260 (N_44260,N_41456,N_41171);
nor U44261 (N_44261,N_41378,N_42014);
xnor U44262 (N_44262,N_40133,N_40273);
and U44263 (N_44263,N_40062,N_41757);
nand U44264 (N_44264,N_41391,N_41469);
nand U44265 (N_44265,N_41237,N_41629);
xnor U44266 (N_44266,N_40884,N_41097);
or U44267 (N_44267,N_40419,N_40855);
or U44268 (N_44268,N_40296,N_42381);
nand U44269 (N_44269,N_42156,N_40835);
and U44270 (N_44270,N_42107,N_42111);
or U44271 (N_44271,N_40676,N_42067);
or U44272 (N_44272,N_42064,N_41734);
and U44273 (N_44273,N_42047,N_40343);
xor U44274 (N_44274,N_40888,N_40473);
nand U44275 (N_44275,N_40904,N_40917);
nor U44276 (N_44276,N_41928,N_40312);
and U44277 (N_44277,N_41043,N_41824);
or U44278 (N_44278,N_41174,N_40428);
and U44279 (N_44279,N_41889,N_41171);
and U44280 (N_44280,N_41045,N_40374);
nand U44281 (N_44281,N_40841,N_40376);
or U44282 (N_44282,N_42457,N_41868);
or U44283 (N_44283,N_41648,N_41437);
and U44284 (N_44284,N_40547,N_40390);
nand U44285 (N_44285,N_40815,N_40795);
nor U44286 (N_44286,N_40544,N_40975);
or U44287 (N_44287,N_41611,N_40978);
nor U44288 (N_44288,N_41555,N_42279);
nor U44289 (N_44289,N_41783,N_40481);
or U44290 (N_44290,N_40132,N_40253);
xor U44291 (N_44291,N_41682,N_41293);
or U44292 (N_44292,N_41217,N_41301);
nand U44293 (N_44293,N_41754,N_40972);
or U44294 (N_44294,N_40989,N_40795);
nor U44295 (N_44295,N_41678,N_40345);
xor U44296 (N_44296,N_40658,N_40924);
or U44297 (N_44297,N_42314,N_40515);
and U44298 (N_44298,N_41768,N_42449);
xnor U44299 (N_44299,N_41894,N_40802);
nand U44300 (N_44300,N_41366,N_40534);
or U44301 (N_44301,N_40147,N_41173);
or U44302 (N_44302,N_40742,N_41727);
and U44303 (N_44303,N_41626,N_40913);
and U44304 (N_44304,N_41679,N_41177);
nand U44305 (N_44305,N_40244,N_40795);
and U44306 (N_44306,N_40374,N_42493);
xnor U44307 (N_44307,N_40638,N_40709);
nor U44308 (N_44308,N_41608,N_40013);
nor U44309 (N_44309,N_40573,N_41095);
or U44310 (N_44310,N_41177,N_40477);
nor U44311 (N_44311,N_41027,N_40207);
and U44312 (N_44312,N_41228,N_42198);
xor U44313 (N_44313,N_41347,N_41623);
nand U44314 (N_44314,N_40612,N_40155);
xor U44315 (N_44315,N_41098,N_40557);
nand U44316 (N_44316,N_40926,N_40267);
and U44317 (N_44317,N_40340,N_41855);
and U44318 (N_44318,N_41082,N_41808);
xnor U44319 (N_44319,N_42287,N_42213);
nand U44320 (N_44320,N_41585,N_40642);
nand U44321 (N_44321,N_40847,N_40414);
nor U44322 (N_44322,N_41444,N_40161);
nor U44323 (N_44323,N_41167,N_41550);
xor U44324 (N_44324,N_41737,N_42321);
and U44325 (N_44325,N_40948,N_42434);
or U44326 (N_44326,N_40253,N_41448);
xor U44327 (N_44327,N_41566,N_41348);
xor U44328 (N_44328,N_42434,N_40001);
xor U44329 (N_44329,N_40521,N_41972);
nor U44330 (N_44330,N_40638,N_40590);
nor U44331 (N_44331,N_41504,N_40324);
or U44332 (N_44332,N_41202,N_42027);
nand U44333 (N_44333,N_40545,N_42223);
and U44334 (N_44334,N_40936,N_40310);
nor U44335 (N_44335,N_40333,N_41456);
xor U44336 (N_44336,N_41816,N_40689);
nand U44337 (N_44337,N_42006,N_40770);
xnor U44338 (N_44338,N_41110,N_41823);
nor U44339 (N_44339,N_40824,N_41336);
xnor U44340 (N_44340,N_41297,N_40402);
or U44341 (N_44341,N_40556,N_42301);
or U44342 (N_44342,N_40071,N_42389);
xor U44343 (N_44343,N_40515,N_40193);
nand U44344 (N_44344,N_40141,N_42131);
nand U44345 (N_44345,N_40991,N_41160);
and U44346 (N_44346,N_42249,N_40999);
xnor U44347 (N_44347,N_40443,N_40803);
or U44348 (N_44348,N_42192,N_42196);
nand U44349 (N_44349,N_41145,N_41044);
nand U44350 (N_44350,N_42085,N_41890);
nand U44351 (N_44351,N_40956,N_41776);
xnor U44352 (N_44352,N_41265,N_40062);
nand U44353 (N_44353,N_42210,N_40123);
nor U44354 (N_44354,N_40917,N_40019);
or U44355 (N_44355,N_42165,N_40676);
or U44356 (N_44356,N_41766,N_41157);
and U44357 (N_44357,N_42357,N_40919);
nand U44358 (N_44358,N_41984,N_40081);
xnor U44359 (N_44359,N_41579,N_40861);
nor U44360 (N_44360,N_40610,N_42282);
xor U44361 (N_44361,N_40514,N_40436);
xnor U44362 (N_44362,N_40712,N_42122);
and U44363 (N_44363,N_41164,N_41022);
or U44364 (N_44364,N_41711,N_40194);
nor U44365 (N_44365,N_40722,N_41840);
xnor U44366 (N_44366,N_40238,N_40688);
and U44367 (N_44367,N_41793,N_41532);
and U44368 (N_44368,N_41778,N_41422);
nor U44369 (N_44369,N_42227,N_40625);
or U44370 (N_44370,N_40790,N_40736);
nand U44371 (N_44371,N_40586,N_41437);
nor U44372 (N_44372,N_40967,N_40068);
xnor U44373 (N_44373,N_40274,N_41311);
nand U44374 (N_44374,N_42052,N_42202);
or U44375 (N_44375,N_40172,N_40060);
nor U44376 (N_44376,N_41989,N_40802);
and U44377 (N_44377,N_40100,N_41927);
nor U44378 (N_44378,N_40998,N_42200);
nor U44379 (N_44379,N_41388,N_41218);
nand U44380 (N_44380,N_41756,N_40087);
xnor U44381 (N_44381,N_41788,N_42372);
nand U44382 (N_44382,N_42101,N_42283);
nor U44383 (N_44383,N_41474,N_41242);
nand U44384 (N_44384,N_40721,N_42239);
nor U44385 (N_44385,N_40978,N_41551);
nor U44386 (N_44386,N_40657,N_40096);
and U44387 (N_44387,N_40511,N_42125);
or U44388 (N_44388,N_42187,N_40388);
and U44389 (N_44389,N_42022,N_42149);
nor U44390 (N_44390,N_40654,N_40340);
nand U44391 (N_44391,N_41167,N_41293);
nor U44392 (N_44392,N_42184,N_40995);
nor U44393 (N_44393,N_41665,N_40863);
and U44394 (N_44394,N_42144,N_41940);
nor U44395 (N_44395,N_42362,N_42297);
and U44396 (N_44396,N_40520,N_41231);
nand U44397 (N_44397,N_42108,N_40148);
or U44398 (N_44398,N_41916,N_40149);
nand U44399 (N_44399,N_40837,N_41246);
xor U44400 (N_44400,N_41808,N_40167);
xnor U44401 (N_44401,N_42347,N_40958);
nor U44402 (N_44402,N_40158,N_40558);
or U44403 (N_44403,N_42239,N_41972);
and U44404 (N_44404,N_41907,N_42089);
xor U44405 (N_44405,N_40567,N_40019);
nand U44406 (N_44406,N_41895,N_41983);
nand U44407 (N_44407,N_41484,N_40054);
or U44408 (N_44408,N_41011,N_41488);
or U44409 (N_44409,N_40333,N_42334);
nand U44410 (N_44410,N_42000,N_41514);
or U44411 (N_44411,N_42122,N_41466);
or U44412 (N_44412,N_40627,N_41143);
xor U44413 (N_44413,N_40738,N_41890);
or U44414 (N_44414,N_40456,N_40807);
nand U44415 (N_44415,N_40601,N_41052);
and U44416 (N_44416,N_41972,N_42163);
xnor U44417 (N_44417,N_40755,N_40041);
nor U44418 (N_44418,N_41255,N_41026);
nor U44419 (N_44419,N_42043,N_41750);
nor U44420 (N_44420,N_40020,N_40678);
or U44421 (N_44421,N_42100,N_40309);
nor U44422 (N_44422,N_40948,N_40137);
and U44423 (N_44423,N_41457,N_42175);
or U44424 (N_44424,N_41034,N_41257);
nor U44425 (N_44425,N_41324,N_41332);
and U44426 (N_44426,N_41810,N_41556);
nand U44427 (N_44427,N_40834,N_41429);
xnor U44428 (N_44428,N_40336,N_42211);
or U44429 (N_44429,N_41993,N_41783);
or U44430 (N_44430,N_41156,N_42135);
nand U44431 (N_44431,N_40302,N_41654);
nand U44432 (N_44432,N_41735,N_42104);
xnor U44433 (N_44433,N_42036,N_40378);
nor U44434 (N_44434,N_40663,N_42051);
nand U44435 (N_44435,N_41608,N_41703);
and U44436 (N_44436,N_41672,N_40243);
and U44437 (N_44437,N_41310,N_40767);
nand U44438 (N_44438,N_42012,N_42394);
or U44439 (N_44439,N_40948,N_40914);
xnor U44440 (N_44440,N_40772,N_41387);
or U44441 (N_44441,N_41328,N_40489);
nand U44442 (N_44442,N_41715,N_41096);
or U44443 (N_44443,N_40931,N_40123);
xor U44444 (N_44444,N_41686,N_41771);
nor U44445 (N_44445,N_41305,N_41578);
xor U44446 (N_44446,N_41303,N_40726);
and U44447 (N_44447,N_41631,N_40637);
nor U44448 (N_44448,N_42005,N_42498);
nand U44449 (N_44449,N_42326,N_41050);
xnor U44450 (N_44450,N_41341,N_42450);
or U44451 (N_44451,N_42470,N_40279);
nor U44452 (N_44452,N_41303,N_41516);
and U44453 (N_44453,N_41310,N_42266);
or U44454 (N_44454,N_41635,N_40044);
or U44455 (N_44455,N_40090,N_40224);
and U44456 (N_44456,N_41028,N_41378);
and U44457 (N_44457,N_40128,N_41004);
or U44458 (N_44458,N_40103,N_41813);
xnor U44459 (N_44459,N_40736,N_40279);
and U44460 (N_44460,N_40678,N_41231);
and U44461 (N_44461,N_40233,N_40088);
or U44462 (N_44462,N_40966,N_42482);
or U44463 (N_44463,N_40601,N_40023);
or U44464 (N_44464,N_42003,N_40318);
nand U44465 (N_44465,N_42319,N_41960);
nor U44466 (N_44466,N_41620,N_41638);
xnor U44467 (N_44467,N_41200,N_40255);
or U44468 (N_44468,N_40761,N_41787);
or U44469 (N_44469,N_41437,N_41986);
xor U44470 (N_44470,N_41620,N_42490);
xor U44471 (N_44471,N_40919,N_41335);
xnor U44472 (N_44472,N_40616,N_40244);
nor U44473 (N_44473,N_40515,N_40893);
nand U44474 (N_44474,N_41539,N_40937);
nor U44475 (N_44475,N_40383,N_41795);
nor U44476 (N_44476,N_41675,N_40557);
and U44477 (N_44477,N_40417,N_41501);
nand U44478 (N_44478,N_41051,N_41248);
or U44479 (N_44479,N_42494,N_40279);
nor U44480 (N_44480,N_41263,N_40063);
or U44481 (N_44481,N_40842,N_41924);
nand U44482 (N_44482,N_40465,N_40265);
and U44483 (N_44483,N_42273,N_41978);
nor U44484 (N_44484,N_42210,N_41747);
nor U44485 (N_44485,N_41455,N_40610);
xor U44486 (N_44486,N_40606,N_41816);
xnor U44487 (N_44487,N_40805,N_40978);
nand U44488 (N_44488,N_40342,N_42002);
nor U44489 (N_44489,N_41025,N_41991);
nor U44490 (N_44490,N_41579,N_41202);
nand U44491 (N_44491,N_41859,N_42338);
or U44492 (N_44492,N_41157,N_40665);
nand U44493 (N_44493,N_41850,N_41059);
and U44494 (N_44494,N_41091,N_40770);
or U44495 (N_44495,N_40407,N_41870);
and U44496 (N_44496,N_40892,N_40203);
xor U44497 (N_44497,N_42286,N_41673);
nand U44498 (N_44498,N_40623,N_40257);
and U44499 (N_44499,N_40276,N_41727);
xor U44500 (N_44500,N_41396,N_41710);
and U44501 (N_44501,N_40127,N_40769);
nand U44502 (N_44502,N_40203,N_41854);
nand U44503 (N_44503,N_41991,N_40541);
nand U44504 (N_44504,N_41175,N_40692);
xnor U44505 (N_44505,N_42150,N_41365);
xor U44506 (N_44506,N_41819,N_40769);
xor U44507 (N_44507,N_41565,N_41668);
or U44508 (N_44508,N_42077,N_41340);
nand U44509 (N_44509,N_40813,N_40047);
nor U44510 (N_44510,N_42004,N_40995);
xnor U44511 (N_44511,N_42027,N_40328);
xor U44512 (N_44512,N_41587,N_41995);
nor U44513 (N_44513,N_41323,N_41847);
nand U44514 (N_44514,N_42078,N_40844);
and U44515 (N_44515,N_42138,N_40445);
xor U44516 (N_44516,N_42050,N_41779);
and U44517 (N_44517,N_41607,N_40701);
or U44518 (N_44518,N_41736,N_41041);
and U44519 (N_44519,N_41434,N_40190);
nand U44520 (N_44520,N_40174,N_41528);
xnor U44521 (N_44521,N_40741,N_40336);
or U44522 (N_44522,N_41295,N_41663);
xor U44523 (N_44523,N_41553,N_40259);
nand U44524 (N_44524,N_41680,N_40440);
nor U44525 (N_44525,N_40656,N_42318);
or U44526 (N_44526,N_40796,N_40214);
xnor U44527 (N_44527,N_42383,N_41979);
or U44528 (N_44528,N_40262,N_41919);
and U44529 (N_44529,N_42062,N_41734);
nor U44530 (N_44530,N_42303,N_41952);
and U44531 (N_44531,N_41507,N_41543);
nor U44532 (N_44532,N_40350,N_40712);
xnor U44533 (N_44533,N_41585,N_40220);
xnor U44534 (N_44534,N_40183,N_40961);
xor U44535 (N_44535,N_41280,N_41175);
xnor U44536 (N_44536,N_40426,N_42445);
xnor U44537 (N_44537,N_41258,N_42479);
or U44538 (N_44538,N_40623,N_40645);
xor U44539 (N_44539,N_42385,N_40369);
and U44540 (N_44540,N_41457,N_42341);
xor U44541 (N_44541,N_41021,N_40340);
or U44542 (N_44542,N_40234,N_41828);
and U44543 (N_44543,N_40199,N_42368);
or U44544 (N_44544,N_40992,N_40342);
or U44545 (N_44545,N_40221,N_40777);
xor U44546 (N_44546,N_41349,N_40780);
nand U44547 (N_44547,N_40329,N_41573);
and U44548 (N_44548,N_40823,N_42339);
nand U44549 (N_44549,N_40289,N_40967);
or U44550 (N_44550,N_41606,N_42057);
nor U44551 (N_44551,N_41561,N_40599);
and U44552 (N_44552,N_41874,N_41720);
nor U44553 (N_44553,N_41738,N_42119);
or U44554 (N_44554,N_40686,N_42240);
xor U44555 (N_44555,N_42416,N_41454);
nand U44556 (N_44556,N_41467,N_40790);
nor U44557 (N_44557,N_41270,N_40290);
nor U44558 (N_44558,N_40329,N_42248);
xnor U44559 (N_44559,N_40703,N_41923);
nand U44560 (N_44560,N_41927,N_41060);
or U44561 (N_44561,N_40687,N_40740);
nand U44562 (N_44562,N_41884,N_41005);
and U44563 (N_44563,N_42489,N_40194);
and U44564 (N_44564,N_42361,N_42416);
or U44565 (N_44565,N_40414,N_40261);
and U44566 (N_44566,N_40123,N_41583);
or U44567 (N_44567,N_42063,N_41434);
nor U44568 (N_44568,N_41199,N_40798);
xor U44569 (N_44569,N_40984,N_40061);
and U44570 (N_44570,N_40181,N_42001);
and U44571 (N_44571,N_40247,N_41985);
xnor U44572 (N_44572,N_42440,N_41698);
nand U44573 (N_44573,N_40806,N_41906);
or U44574 (N_44574,N_40215,N_40744);
nand U44575 (N_44575,N_42040,N_40246);
and U44576 (N_44576,N_41403,N_40510);
nor U44577 (N_44577,N_41019,N_40706);
nand U44578 (N_44578,N_40197,N_42253);
or U44579 (N_44579,N_40153,N_41356);
and U44580 (N_44580,N_40346,N_42060);
nor U44581 (N_44581,N_41775,N_41478);
xnor U44582 (N_44582,N_41362,N_42216);
or U44583 (N_44583,N_40245,N_42331);
nor U44584 (N_44584,N_41430,N_40032);
nor U44585 (N_44585,N_42104,N_40243);
and U44586 (N_44586,N_40647,N_40726);
or U44587 (N_44587,N_40483,N_40577);
or U44588 (N_44588,N_41928,N_40885);
nor U44589 (N_44589,N_42147,N_40587);
nand U44590 (N_44590,N_41513,N_42216);
or U44591 (N_44591,N_42166,N_40603);
or U44592 (N_44592,N_40960,N_40668);
xor U44593 (N_44593,N_40130,N_41335);
nand U44594 (N_44594,N_40323,N_41598);
nand U44595 (N_44595,N_40811,N_40631);
nand U44596 (N_44596,N_41626,N_41517);
xor U44597 (N_44597,N_41636,N_41037);
or U44598 (N_44598,N_41366,N_41099);
nor U44599 (N_44599,N_42393,N_40124);
nor U44600 (N_44600,N_42435,N_40469);
nor U44601 (N_44601,N_40314,N_40814);
nand U44602 (N_44602,N_40581,N_40555);
or U44603 (N_44603,N_40434,N_41161);
xnor U44604 (N_44604,N_40882,N_41315);
xor U44605 (N_44605,N_40820,N_41916);
nand U44606 (N_44606,N_40525,N_40549);
nor U44607 (N_44607,N_40614,N_40915);
xnor U44608 (N_44608,N_40662,N_41674);
nand U44609 (N_44609,N_41335,N_40629);
nor U44610 (N_44610,N_41165,N_40578);
nand U44611 (N_44611,N_42251,N_41515);
nor U44612 (N_44612,N_40491,N_40882);
nand U44613 (N_44613,N_41731,N_42215);
and U44614 (N_44614,N_41596,N_41328);
xor U44615 (N_44615,N_40442,N_41408);
xor U44616 (N_44616,N_42007,N_41397);
and U44617 (N_44617,N_40311,N_41795);
nand U44618 (N_44618,N_40008,N_42285);
xor U44619 (N_44619,N_42350,N_40435);
xor U44620 (N_44620,N_41455,N_40971);
and U44621 (N_44621,N_40687,N_40647);
or U44622 (N_44622,N_40485,N_40709);
or U44623 (N_44623,N_40970,N_40769);
xnor U44624 (N_44624,N_41527,N_41158);
nor U44625 (N_44625,N_42184,N_40830);
nand U44626 (N_44626,N_40193,N_41778);
nor U44627 (N_44627,N_40190,N_40222);
xor U44628 (N_44628,N_41765,N_41410);
xnor U44629 (N_44629,N_41795,N_40006);
xor U44630 (N_44630,N_42041,N_41898);
nor U44631 (N_44631,N_41847,N_42326);
xnor U44632 (N_44632,N_40491,N_41540);
xor U44633 (N_44633,N_40329,N_41796);
and U44634 (N_44634,N_41807,N_40806);
or U44635 (N_44635,N_40766,N_40750);
nand U44636 (N_44636,N_41357,N_40263);
xnor U44637 (N_44637,N_41916,N_41288);
xor U44638 (N_44638,N_41686,N_40696);
and U44639 (N_44639,N_41191,N_40758);
nand U44640 (N_44640,N_42419,N_42248);
nor U44641 (N_44641,N_41239,N_40340);
xnor U44642 (N_44642,N_40041,N_41702);
or U44643 (N_44643,N_40653,N_40041);
or U44644 (N_44644,N_42391,N_42160);
xnor U44645 (N_44645,N_42408,N_41506);
or U44646 (N_44646,N_41572,N_42200);
or U44647 (N_44647,N_42460,N_40482);
nand U44648 (N_44648,N_42104,N_41365);
xnor U44649 (N_44649,N_40495,N_40411);
nor U44650 (N_44650,N_40359,N_41271);
and U44651 (N_44651,N_40489,N_41567);
or U44652 (N_44652,N_40665,N_40148);
or U44653 (N_44653,N_40066,N_41784);
or U44654 (N_44654,N_40936,N_40222);
nor U44655 (N_44655,N_40669,N_40906);
nor U44656 (N_44656,N_41685,N_41954);
or U44657 (N_44657,N_40281,N_42119);
nand U44658 (N_44658,N_41451,N_40374);
nor U44659 (N_44659,N_40696,N_41837);
nand U44660 (N_44660,N_40678,N_42397);
or U44661 (N_44661,N_41862,N_41770);
nor U44662 (N_44662,N_41258,N_40405);
nand U44663 (N_44663,N_40575,N_40032);
nand U44664 (N_44664,N_42110,N_40992);
and U44665 (N_44665,N_41601,N_42104);
and U44666 (N_44666,N_40238,N_42269);
nand U44667 (N_44667,N_42388,N_41251);
and U44668 (N_44668,N_41443,N_40070);
nand U44669 (N_44669,N_40677,N_40306);
nand U44670 (N_44670,N_41940,N_41846);
xnor U44671 (N_44671,N_40941,N_41306);
nor U44672 (N_44672,N_40927,N_42420);
nand U44673 (N_44673,N_42193,N_42084);
nor U44674 (N_44674,N_40195,N_41946);
xnor U44675 (N_44675,N_40553,N_41001);
nor U44676 (N_44676,N_40885,N_40042);
or U44677 (N_44677,N_40627,N_41151);
nand U44678 (N_44678,N_40389,N_42440);
or U44679 (N_44679,N_41560,N_42301);
xor U44680 (N_44680,N_42012,N_41104);
nor U44681 (N_44681,N_42453,N_40406);
nor U44682 (N_44682,N_40126,N_41705);
nand U44683 (N_44683,N_41423,N_40009);
nand U44684 (N_44684,N_41231,N_42146);
nand U44685 (N_44685,N_41611,N_40840);
xor U44686 (N_44686,N_40479,N_41080);
nor U44687 (N_44687,N_41501,N_41585);
nor U44688 (N_44688,N_41752,N_40671);
or U44689 (N_44689,N_40735,N_42161);
nand U44690 (N_44690,N_41584,N_41326);
nand U44691 (N_44691,N_40108,N_41160);
xnor U44692 (N_44692,N_40366,N_41555);
and U44693 (N_44693,N_40364,N_40269);
or U44694 (N_44694,N_40717,N_41464);
nor U44695 (N_44695,N_41180,N_40116);
or U44696 (N_44696,N_40727,N_40058);
and U44697 (N_44697,N_40786,N_41972);
nor U44698 (N_44698,N_40429,N_40043);
nor U44699 (N_44699,N_40400,N_41171);
nor U44700 (N_44700,N_40796,N_41774);
and U44701 (N_44701,N_40073,N_41329);
and U44702 (N_44702,N_40617,N_41717);
and U44703 (N_44703,N_42445,N_41061);
nor U44704 (N_44704,N_40413,N_42050);
or U44705 (N_44705,N_41805,N_42393);
nor U44706 (N_44706,N_40163,N_41288);
and U44707 (N_44707,N_41391,N_41579);
nand U44708 (N_44708,N_40167,N_40127);
or U44709 (N_44709,N_41719,N_41422);
nor U44710 (N_44710,N_42032,N_40559);
or U44711 (N_44711,N_42062,N_40253);
and U44712 (N_44712,N_41651,N_40870);
and U44713 (N_44713,N_41058,N_40907);
or U44714 (N_44714,N_42088,N_41923);
xor U44715 (N_44715,N_41379,N_40239);
nor U44716 (N_44716,N_40184,N_41668);
and U44717 (N_44717,N_40730,N_40814);
or U44718 (N_44718,N_40102,N_40734);
xor U44719 (N_44719,N_41014,N_40825);
or U44720 (N_44720,N_42280,N_40147);
nor U44721 (N_44721,N_41712,N_40828);
or U44722 (N_44722,N_41018,N_41266);
nand U44723 (N_44723,N_41208,N_40735);
and U44724 (N_44724,N_41443,N_40942);
nor U44725 (N_44725,N_40081,N_42352);
xnor U44726 (N_44726,N_42272,N_42497);
and U44727 (N_44727,N_40796,N_40070);
nor U44728 (N_44728,N_40730,N_41931);
nor U44729 (N_44729,N_40636,N_40757);
xor U44730 (N_44730,N_42016,N_40182);
and U44731 (N_44731,N_40824,N_40096);
nand U44732 (N_44732,N_41414,N_40520);
xor U44733 (N_44733,N_41626,N_42018);
nand U44734 (N_44734,N_41523,N_40405);
nand U44735 (N_44735,N_41374,N_41345);
nand U44736 (N_44736,N_41914,N_40061);
nand U44737 (N_44737,N_41174,N_41644);
or U44738 (N_44738,N_40918,N_40465);
nor U44739 (N_44739,N_41427,N_41435);
nor U44740 (N_44740,N_40779,N_41776);
xnor U44741 (N_44741,N_40452,N_41806);
or U44742 (N_44742,N_41042,N_42334);
and U44743 (N_44743,N_40074,N_41663);
and U44744 (N_44744,N_40878,N_41381);
xor U44745 (N_44745,N_41387,N_40429);
nor U44746 (N_44746,N_42083,N_40476);
or U44747 (N_44747,N_40852,N_40276);
nand U44748 (N_44748,N_40294,N_41833);
and U44749 (N_44749,N_40743,N_40334);
or U44750 (N_44750,N_40893,N_41011);
nand U44751 (N_44751,N_40198,N_40206);
nand U44752 (N_44752,N_41412,N_40235);
and U44753 (N_44753,N_41373,N_42433);
nor U44754 (N_44754,N_40019,N_41698);
xnor U44755 (N_44755,N_40706,N_40785);
nor U44756 (N_44756,N_41957,N_42240);
or U44757 (N_44757,N_41183,N_40778);
xnor U44758 (N_44758,N_41112,N_41402);
or U44759 (N_44759,N_41177,N_42097);
nand U44760 (N_44760,N_40877,N_40282);
xor U44761 (N_44761,N_42451,N_40604);
nand U44762 (N_44762,N_41204,N_41758);
nor U44763 (N_44763,N_40366,N_40333);
and U44764 (N_44764,N_42258,N_40806);
xnor U44765 (N_44765,N_40401,N_41802);
xor U44766 (N_44766,N_42118,N_42430);
and U44767 (N_44767,N_42460,N_41375);
nand U44768 (N_44768,N_40204,N_41522);
nor U44769 (N_44769,N_40824,N_42350);
nor U44770 (N_44770,N_42431,N_40249);
and U44771 (N_44771,N_40933,N_41379);
nand U44772 (N_44772,N_40526,N_41962);
or U44773 (N_44773,N_41438,N_41624);
nor U44774 (N_44774,N_42176,N_40323);
nand U44775 (N_44775,N_42080,N_40343);
nor U44776 (N_44776,N_41424,N_41220);
nand U44777 (N_44777,N_41546,N_42347);
or U44778 (N_44778,N_40243,N_40155);
nand U44779 (N_44779,N_40251,N_41730);
xnor U44780 (N_44780,N_42333,N_40197);
nand U44781 (N_44781,N_41761,N_41170);
nor U44782 (N_44782,N_41297,N_41010);
nor U44783 (N_44783,N_41697,N_41604);
and U44784 (N_44784,N_40699,N_40102);
nor U44785 (N_44785,N_40972,N_40041);
nand U44786 (N_44786,N_41192,N_40311);
xor U44787 (N_44787,N_41651,N_42383);
and U44788 (N_44788,N_41114,N_42419);
nor U44789 (N_44789,N_41631,N_40230);
and U44790 (N_44790,N_41121,N_41439);
and U44791 (N_44791,N_40095,N_40961);
and U44792 (N_44792,N_42174,N_41904);
nor U44793 (N_44793,N_41967,N_42319);
nor U44794 (N_44794,N_40334,N_40643);
nor U44795 (N_44795,N_41849,N_42049);
xnor U44796 (N_44796,N_42117,N_42255);
nor U44797 (N_44797,N_40838,N_40887);
and U44798 (N_44798,N_41995,N_41570);
xor U44799 (N_44799,N_41537,N_42119);
or U44800 (N_44800,N_42152,N_40676);
nor U44801 (N_44801,N_40731,N_40013);
xnor U44802 (N_44802,N_42005,N_40931);
nand U44803 (N_44803,N_41006,N_41112);
nand U44804 (N_44804,N_40870,N_40208);
nand U44805 (N_44805,N_40980,N_42194);
and U44806 (N_44806,N_41147,N_41839);
nand U44807 (N_44807,N_40818,N_40392);
nor U44808 (N_44808,N_40201,N_40425);
xor U44809 (N_44809,N_41470,N_42167);
and U44810 (N_44810,N_41834,N_41904);
xor U44811 (N_44811,N_41213,N_41154);
xor U44812 (N_44812,N_41811,N_41337);
nor U44813 (N_44813,N_42328,N_41149);
xor U44814 (N_44814,N_40031,N_41398);
and U44815 (N_44815,N_42268,N_41999);
and U44816 (N_44816,N_40188,N_41315);
xor U44817 (N_44817,N_41759,N_41795);
nand U44818 (N_44818,N_40873,N_41196);
or U44819 (N_44819,N_40359,N_40586);
nor U44820 (N_44820,N_42308,N_42374);
nand U44821 (N_44821,N_42265,N_40796);
or U44822 (N_44822,N_40323,N_40238);
xor U44823 (N_44823,N_42355,N_41097);
xnor U44824 (N_44824,N_40771,N_40074);
and U44825 (N_44825,N_41293,N_40904);
nand U44826 (N_44826,N_40113,N_41723);
and U44827 (N_44827,N_41178,N_40645);
and U44828 (N_44828,N_42038,N_41251);
nand U44829 (N_44829,N_40672,N_40841);
nand U44830 (N_44830,N_40889,N_42195);
and U44831 (N_44831,N_40727,N_41815);
and U44832 (N_44832,N_41425,N_40127);
xnor U44833 (N_44833,N_40168,N_41848);
or U44834 (N_44834,N_41437,N_40388);
nor U44835 (N_44835,N_40705,N_41650);
and U44836 (N_44836,N_41640,N_42291);
and U44837 (N_44837,N_40525,N_42017);
nand U44838 (N_44838,N_41496,N_41875);
or U44839 (N_44839,N_42083,N_42306);
and U44840 (N_44840,N_40457,N_41235);
or U44841 (N_44841,N_40145,N_41984);
or U44842 (N_44842,N_41614,N_40186);
or U44843 (N_44843,N_41426,N_41846);
xnor U44844 (N_44844,N_41858,N_41815);
xnor U44845 (N_44845,N_41574,N_42420);
nand U44846 (N_44846,N_40232,N_41161);
xnor U44847 (N_44847,N_41743,N_40156);
xnor U44848 (N_44848,N_41074,N_41415);
nor U44849 (N_44849,N_42378,N_42146);
and U44850 (N_44850,N_42349,N_40271);
nor U44851 (N_44851,N_41868,N_41500);
nor U44852 (N_44852,N_40087,N_40971);
or U44853 (N_44853,N_41672,N_42258);
and U44854 (N_44854,N_41442,N_40877);
xnor U44855 (N_44855,N_41414,N_41946);
xnor U44856 (N_44856,N_41644,N_41120);
xor U44857 (N_44857,N_41047,N_40841);
nor U44858 (N_44858,N_40872,N_40467);
nor U44859 (N_44859,N_41227,N_42249);
nand U44860 (N_44860,N_41376,N_42468);
xnor U44861 (N_44861,N_42303,N_40481);
and U44862 (N_44862,N_40391,N_41896);
nand U44863 (N_44863,N_40351,N_41956);
nand U44864 (N_44864,N_40849,N_41053);
and U44865 (N_44865,N_41702,N_40383);
nor U44866 (N_44866,N_40912,N_41187);
xor U44867 (N_44867,N_42447,N_40675);
and U44868 (N_44868,N_41279,N_41352);
nor U44869 (N_44869,N_41418,N_41597);
xor U44870 (N_44870,N_41761,N_41676);
nand U44871 (N_44871,N_40111,N_40485);
nor U44872 (N_44872,N_41451,N_42019);
nand U44873 (N_44873,N_42431,N_41969);
xnor U44874 (N_44874,N_40627,N_41395);
or U44875 (N_44875,N_40439,N_40583);
and U44876 (N_44876,N_40477,N_40732);
or U44877 (N_44877,N_41660,N_41052);
nand U44878 (N_44878,N_41706,N_40212);
nor U44879 (N_44879,N_40647,N_40505);
or U44880 (N_44880,N_41393,N_40400);
xor U44881 (N_44881,N_40750,N_40638);
nor U44882 (N_44882,N_41739,N_41315);
and U44883 (N_44883,N_40708,N_40918);
xor U44884 (N_44884,N_41787,N_41192);
nand U44885 (N_44885,N_41391,N_41528);
nor U44886 (N_44886,N_40281,N_41392);
or U44887 (N_44887,N_41872,N_42254);
nor U44888 (N_44888,N_41638,N_40961);
nand U44889 (N_44889,N_42263,N_40821);
xor U44890 (N_44890,N_42184,N_41030);
or U44891 (N_44891,N_41044,N_40702);
or U44892 (N_44892,N_42404,N_42164);
or U44893 (N_44893,N_40744,N_40797);
or U44894 (N_44894,N_40908,N_42163);
and U44895 (N_44895,N_40006,N_41090);
or U44896 (N_44896,N_42003,N_40826);
nand U44897 (N_44897,N_41081,N_42209);
or U44898 (N_44898,N_41272,N_41068);
and U44899 (N_44899,N_42447,N_42231);
nand U44900 (N_44900,N_40960,N_40810);
nor U44901 (N_44901,N_41577,N_41574);
nor U44902 (N_44902,N_42079,N_40822);
nor U44903 (N_44903,N_40274,N_41896);
and U44904 (N_44904,N_40769,N_41806);
or U44905 (N_44905,N_40107,N_40401);
and U44906 (N_44906,N_42308,N_41874);
xor U44907 (N_44907,N_41879,N_42313);
nand U44908 (N_44908,N_40639,N_40790);
nor U44909 (N_44909,N_41355,N_40519);
nor U44910 (N_44910,N_41759,N_40850);
xnor U44911 (N_44911,N_41195,N_40242);
and U44912 (N_44912,N_40717,N_41746);
nand U44913 (N_44913,N_40010,N_42486);
or U44914 (N_44914,N_41678,N_42269);
xor U44915 (N_44915,N_41936,N_42152);
xor U44916 (N_44916,N_40504,N_41420);
or U44917 (N_44917,N_41293,N_42163);
nand U44918 (N_44918,N_42106,N_42065);
nand U44919 (N_44919,N_40413,N_40688);
nor U44920 (N_44920,N_40918,N_40442);
and U44921 (N_44921,N_40955,N_41558);
xnor U44922 (N_44922,N_40344,N_40867);
and U44923 (N_44923,N_40573,N_40192);
nor U44924 (N_44924,N_40627,N_41717);
xnor U44925 (N_44925,N_41664,N_40562);
nor U44926 (N_44926,N_40977,N_41209);
and U44927 (N_44927,N_42373,N_40501);
nand U44928 (N_44928,N_41916,N_42210);
nand U44929 (N_44929,N_40248,N_40112);
xor U44930 (N_44930,N_42109,N_41767);
nand U44931 (N_44931,N_40011,N_41111);
nand U44932 (N_44932,N_41049,N_40405);
nand U44933 (N_44933,N_41628,N_40470);
nand U44934 (N_44934,N_40256,N_41450);
xnor U44935 (N_44935,N_40858,N_41237);
or U44936 (N_44936,N_40680,N_41567);
or U44937 (N_44937,N_41570,N_40812);
nor U44938 (N_44938,N_40418,N_40861);
nand U44939 (N_44939,N_41524,N_42329);
or U44940 (N_44940,N_41994,N_42422);
xor U44941 (N_44941,N_41923,N_41776);
and U44942 (N_44942,N_41780,N_42096);
nor U44943 (N_44943,N_40907,N_41878);
xor U44944 (N_44944,N_40963,N_42206);
and U44945 (N_44945,N_40494,N_41564);
and U44946 (N_44946,N_41513,N_42351);
xor U44947 (N_44947,N_41333,N_41449);
nand U44948 (N_44948,N_41780,N_42073);
nand U44949 (N_44949,N_40422,N_40596);
xor U44950 (N_44950,N_40772,N_42113);
nand U44951 (N_44951,N_40973,N_40521);
nand U44952 (N_44952,N_40971,N_41307);
nand U44953 (N_44953,N_42226,N_40952);
xnor U44954 (N_44954,N_41040,N_41669);
nand U44955 (N_44955,N_41662,N_41038);
and U44956 (N_44956,N_41403,N_42235);
nand U44957 (N_44957,N_41352,N_40139);
nand U44958 (N_44958,N_40966,N_41536);
nor U44959 (N_44959,N_42272,N_40949);
nor U44960 (N_44960,N_41073,N_41837);
or U44961 (N_44961,N_40003,N_41817);
or U44962 (N_44962,N_40152,N_42395);
and U44963 (N_44963,N_41049,N_40929);
nand U44964 (N_44964,N_40282,N_41293);
nand U44965 (N_44965,N_41711,N_41167);
and U44966 (N_44966,N_40875,N_42051);
or U44967 (N_44967,N_40940,N_42054);
and U44968 (N_44968,N_40350,N_42051);
or U44969 (N_44969,N_41002,N_41852);
nor U44970 (N_44970,N_42077,N_41297);
nor U44971 (N_44971,N_41317,N_41921);
and U44972 (N_44972,N_41982,N_40423);
or U44973 (N_44973,N_41297,N_42401);
xnor U44974 (N_44974,N_41486,N_40701);
nand U44975 (N_44975,N_41738,N_40512);
nand U44976 (N_44976,N_41294,N_40925);
or U44977 (N_44977,N_42125,N_42024);
or U44978 (N_44978,N_41261,N_42282);
nor U44979 (N_44979,N_41342,N_41421);
and U44980 (N_44980,N_42485,N_40179);
and U44981 (N_44981,N_42492,N_41988);
nor U44982 (N_44982,N_42298,N_40373);
nand U44983 (N_44983,N_40880,N_40090);
nor U44984 (N_44984,N_40252,N_41102);
and U44985 (N_44985,N_41005,N_41977);
xnor U44986 (N_44986,N_40939,N_41440);
or U44987 (N_44987,N_42347,N_42278);
nand U44988 (N_44988,N_42170,N_41059);
and U44989 (N_44989,N_41087,N_40811);
and U44990 (N_44990,N_40062,N_41453);
and U44991 (N_44991,N_40756,N_41475);
nor U44992 (N_44992,N_41174,N_42309);
nor U44993 (N_44993,N_40376,N_40250);
nand U44994 (N_44994,N_42103,N_40739);
and U44995 (N_44995,N_41880,N_41448);
or U44996 (N_44996,N_40645,N_40413);
or U44997 (N_44997,N_40754,N_41192);
and U44998 (N_44998,N_40104,N_41750);
nand U44999 (N_44999,N_41994,N_40091);
xor U45000 (N_45000,N_43743,N_43642);
xor U45001 (N_45001,N_44638,N_42528);
and U45002 (N_45002,N_42888,N_42684);
and U45003 (N_45003,N_44708,N_44559);
nand U45004 (N_45004,N_42617,N_43682);
and U45005 (N_45005,N_44733,N_44839);
and U45006 (N_45006,N_43805,N_43134);
nor U45007 (N_45007,N_43321,N_42542);
and U45008 (N_45008,N_44918,N_42850);
nand U45009 (N_45009,N_43222,N_43725);
xnor U45010 (N_45010,N_44676,N_44779);
and U45011 (N_45011,N_44109,N_44623);
xnor U45012 (N_45012,N_43639,N_42966);
nor U45013 (N_45013,N_44387,N_43951);
xnor U45014 (N_45014,N_44157,N_43427);
nand U45015 (N_45015,N_43877,N_44028);
or U45016 (N_45016,N_43962,N_44443);
nand U45017 (N_45017,N_42769,N_44322);
and U45018 (N_45018,N_43989,N_44403);
xnor U45019 (N_45019,N_43934,N_42578);
nor U45020 (N_45020,N_42556,N_42603);
nor U45021 (N_45021,N_44139,N_44657);
nor U45022 (N_45022,N_42593,N_42673);
and U45023 (N_45023,N_43358,N_43498);
nand U45024 (N_45024,N_44613,N_43481);
nor U45025 (N_45025,N_43188,N_44801);
nor U45026 (N_45026,N_44499,N_44743);
xor U45027 (N_45027,N_43325,N_43607);
nand U45028 (N_45028,N_44633,N_43640);
or U45029 (N_45029,N_44718,N_44594);
or U45030 (N_45030,N_43115,N_44212);
nand U45031 (N_45031,N_43081,N_44977);
nand U45032 (N_45032,N_44902,N_42747);
xnor U45033 (N_45033,N_44866,N_43402);
nor U45034 (N_45034,N_43127,N_43944);
or U45035 (N_45035,N_42707,N_43233);
nor U45036 (N_45036,N_43087,N_44531);
xnor U45037 (N_45037,N_43982,N_43373);
or U45038 (N_45038,N_44588,N_44787);
and U45039 (N_45039,N_43330,N_43273);
or U45040 (N_45040,N_42517,N_43089);
or U45041 (N_45041,N_44999,N_42989);
nor U45042 (N_45042,N_43935,N_42735);
and U45043 (N_45043,N_44347,N_42822);
and U45044 (N_45044,N_44105,N_42509);
and U45045 (N_45045,N_43447,N_44686);
nand U45046 (N_45046,N_43984,N_43199);
nor U45047 (N_45047,N_42997,N_42574);
or U45048 (N_45048,N_43119,N_44027);
and U45049 (N_45049,N_43326,N_44989);
and U45050 (N_45050,N_43423,N_42959);
nor U45051 (N_45051,N_42702,N_43223);
nand U45052 (N_45052,N_43336,N_44750);
or U45053 (N_45053,N_42543,N_43974);
xor U45054 (N_45054,N_44771,N_43290);
xor U45055 (N_45055,N_43256,N_44389);
and U45056 (N_45056,N_43605,N_44712);
and U45057 (N_45057,N_44515,N_42787);
nand U45058 (N_45058,N_43202,N_44058);
nand U45059 (N_45059,N_44493,N_44512);
and U45060 (N_45060,N_44348,N_43039);
xnor U45061 (N_45061,N_43339,N_42653);
or U45062 (N_45062,N_43849,N_43883);
nor U45063 (N_45063,N_44184,N_44042);
xnor U45064 (N_45064,N_43026,N_43872);
nand U45065 (N_45065,N_43917,N_42937);
and U45066 (N_45066,N_44381,N_43896);
nor U45067 (N_45067,N_43296,N_44240);
and U45068 (N_45068,N_43588,N_42764);
nor U45069 (N_45069,N_44268,N_43651);
nand U45070 (N_45070,N_43502,N_44262);
or U45071 (N_45071,N_42753,N_42786);
or U45072 (N_45072,N_44907,N_43949);
nor U45073 (N_45073,N_42931,N_44821);
nand U45074 (N_45074,N_43307,N_43299);
and U45075 (N_45075,N_43028,N_44417);
nor U45076 (N_45076,N_44796,N_43845);
or U45077 (N_45077,N_44774,N_44746);
xor U45078 (N_45078,N_44501,N_42527);
xor U45079 (N_45079,N_44649,N_42685);
and U45080 (N_45080,N_44220,N_43577);
nand U45081 (N_45081,N_43455,N_42876);
and U45082 (N_45082,N_44552,N_44336);
xor U45083 (N_45083,N_42559,N_42536);
xor U45084 (N_45084,N_43322,N_44441);
nor U45085 (N_45085,N_43758,N_43298);
nor U45086 (N_45086,N_44452,N_44702);
and U45087 (N_45087,N_44186,N_43141);
nor U45088 (N_45088,N_42810,N_43527);
nand U45089 (N_45089,N_42902,N_44674);
nand U45090 (N_45090,N_42908,N_43611);
xor U45091 (N_45091,N_44057,N_44843);
nor U45092 (N_45092,N_44993,N_43467);
xnor U45093 (N_45093,N_44147,N_43704);
or U45094 (N_45094,N_43305,N_43397);
and U45095 (N_45095,N_44786,N_42643);
and U45096 (N_45096,N_43629,N_42526);
nor U45097 (N_45097,N_43647,N_43338);
nand U45098 (N_45098,N_43323,N_44824);
nor U45099 (N_45099,N_42667,N_43614);
and U45100 (N_45100,N_42602,N_43796);
nor U45101 (N_45101,N_43107,N_42636);
xor U45102 (N_45102,N_43462,N_43094);
nand U45103 (N_45103,N_44126,N_43943);
nor U45104 (N_45104,N_43988,N_44880);
nor U45105 (N_45105,N_43329,N_43245);
nor U45106 (N_45106,N_42855,N_43987);
nor U45107 (N_45107,N_43986,N_44954);
nor U45108 (N_45108,N_44433,N_43058);
nor U45109 (N_45109,N_43038,N_42831);
nand U45110 (N_45110,N_44430,N_43822);
or U45111 (N_45111,N_43341,N_42640);
nor U45112 (N_45112,N_42698,N_42979);
xor U45113 (N_45113,N_43473,N_43565);
nor U45114 (N_45114,N_43976,N_44680);
nand U45115 (N_45115,N_44263,N_44216);
nor U45116 (N_45116,N_43215,N_42631);
or U45117 (N_45117,N_43709,N_42942);
nor U45118 (N_45118,N_42915,N_42838);
xnor U45119 (N_45119,N_42955,N_44914);
and U45120 (N_45120,N_44251,N_44491);
nand U45121 (N_45121,N_42866,N_42918);
and U45122 (N_45122,N_43546,N_42803);
or U45123 (N_45123,N_44812,N_42940);
or U45124 (N_45124,N_42569,N_43711);
nor U45125 (N_45125,N_44530,N_43983);
or U45126 (N_45126,N_42875,N_44995);
and U45127 (N_45127,N_43224,N_44445);
nor U45128 (N_45128,N_42862,N_43610);
or U45129 (N_45129,N_42727,N_42991);
xnor U45130 (N_45130,N_44912,N_44078);
or U45131 (N_45131,N_43412,N_44621);
nor U45132 (N_45132,N_42911,N_44951);
nand U45133 (N_45133,N_44713,N_43626);
xnor U45134 (N_45134,N_43411,N_43545);
and U45135 (N_45135,N_44700,N_44352);
and U45136 (N_45136,N_43770,N_43755);
and U45137 (N_45137,N_44000,N_44190);
nand U45138 (N_45138,N_44324,N_42919);
nor U45139 (N_45139,N_43240,N_43733);
nor U45140 (N_45140,N_43852,N_43308);
or U45141 (N_45141,N_44315,N_44500);
nand U45142 (N_45142,N_44580,N_43333);
xor U45143 (N_45143,N_44972,N_44557);
nor U45144 (N_45144,N_43203,N_42880);
xnor U45145 (N_45145,N_43576,N_44304);
and U45146 (N_45146,N_43117,N_44549);
or U45147 (N_45147,N_43049,N_44419);
or U45148 (N_45148,N_44083,N_43732);
nor U45149 (N_45149,N_43419,N_44947);
and U45150 (N_45150,N_43609,N_42515);
nand U45151 (N_45151,N_44023,N_42534);
nand U45152 (N_45152,N_44505,N_44950);
nor U45153 (N_45153,N_42823,N_44992);
and U45154 (N_45154,N_42645,N_44143);
nand U45155 (N_45155,N_44049,N_43621);
nand U45156 (N_45156,N_43372,N_43169);
xor U45157 (N_45157,N_44041,N_43549);
nand U45158 (N_45158,N_42552,N_44583);
xnor U45159 (N_45159,N_44291,N_44660);
or U45160 (N_45160,N_43698,N_42516);
xor U45161 (N_45161,N_42843,N_43820);
or U45162 (N_45162,N_43275,N_44111);
or U45163 (N_45163,N_43137,N_44326);
nand U45164 (N_45164,N_44234,N_44966);
and U45165 (N_45165,N_43513,N_43210);
xnor U45166 (N_45166,N_43531,N_44909);
nand U45167 (N_45167,N_44461,N_43892);
nand U45168 (N_45168,N_42583,N_44150);
nand U45169 (N_45169,N_44114,N_42756);
nor U45170 (N_45170,N_44193,N_44457);
xor U45171 (N_45171,N_42874,N_44905);
or U45172 (N_45172,N_44247,N_43702);
nand U45173 (N_45173,N_43485,N_44760);
and U45174 (N_45174,N_43792,N_43332);
nor U45175 (N_45175,N_42514,N_43713);
and U45176 (N_45176,N_44256,N_43891);
nor U45177 (N_45177,N_44624,N_44802);
nor U45178 (N_45178,N_43666,N_43015);
nor U45179 (N_45179,N_42781,N_43779);
and U45180 (N_45180,N_43497,N_44587);
nor U45181 (N_45181,N_43715,N_42650);
and U45182 (N_45182,N_42683,N_43425);
nand U45183 (N_45183,N_44398,N_43529);
or U45184 (N_45184,N_44390,N_44701);
and U45185 (N_45185,N_44446,N_43008);
nand U45186 (N_45186,N_43186,N_44066);
xor U45187 (N_45187,N_43300,N_43000);
nand U45188 (N_45188,N_44817,N_42701);
and U45189 (N_45189,N_44283,N_43464);
xnor U45190 (N_45190,N_43928,N_44971);
and U45191 (N_45191,N_43041,N_43383);
or U45192 (N_45192,N_44964,N_43838);
nor U45193 (N_45193,N_44362,N_44261);
nor U45194 (N_45194,N_44711,N_44875);
nand U45195 (N_45195,N_44619,N_43649);
xnor U45196 (N_45196,N_44391,N_44202);
nor U45197 (N_45197,N_43446,N_44630);
xor U45198 (N_45198,N_43059,N_43108);
nand U45199 (N_45199,N_44704,N_43694);
nor U45200 (N_45200,N_43449,N_44908);
and U45201 (N_45201,N_42562,N_43154);
nor U45202 (N_45202,N_44545,N_44931);
or U45203 (N_45203,N_43975,N_43551);
or U45204 (N_45204,N_44593,N_44871);
nor U45205 (N_45205,N_43844,N_43350);
xnor U45206 (N_45206,N_44472,N_44020);
nor U45207 (N_45207,N_44260,N_43948);
nand U45208 (N_45208,N_43334,N_42892);
nor U45209 (N_45209,N_43143,N_43109);
and U45210 (N_45210,N_43794,N_44001);
xor U45211 (N_45211,N_42596,N_44395);
xnor U45212 (N_45212,N_42670,N_44665);
and U45213 (N_45213,N_44497,N_44938);
xnor U45214 (N_45214,N_42856,N_43128);
nor U45215 (N_45215,N_44085,N_43748);
and U45216 (N_45216,N_43155,N_42863);
xnor U45217 (N_45217,N_43553,N_42561);
or U45218 (N_45218,N_44181,N_44124);
and U45219 (N_45219,N_42712,N_43825);
or U45220 (N_45220,N_43095,N_44990);
or U45221 (N_45221,N_42928,N_44529);
or U45222 (N_45222,N_43981,N_44280);
or U45223 (N_45223,N_42765,N_43125);
xnor U45224 (N_45224,N_44911,N_43525);
xor U45225 (N_45225,N_43573,N_43759);
nor U45226 (N_45226,N_43633,N_42914);
xnor U45227 (N_45227,N_44946,N_43547);
nor U45228 (N_45228,N_42718,N_42913);
nand U45229 (N_45229,N_43458,N_44282);
or U45230 (N_45230,N_42981,N_42639);
and U45231 (N_45231,N_44749,N_44201);
and U45232 (N_45232,N_43459,N_44050);
xnor U45233 (N_45233,N_44319,N_42879);
or U45234 (N_45234,N_43919,N_42950);
or U45235 (N_45235,N_43631,N_44585);
xor U45236 (N_45236,N_44705,N_43208);
nand U45237 (N_45237,N_43004,N_43739);
and U45238 (N_45238,N_43111,N_42637);
nand U45239 (N_45239,N_42500,N_43368);
xor U45240 (N_45240,N_44761,N_44778);
xnor U45241 (N_45241,N_42677,N_44211);
or U45242 (N_45242,N_43068,N_44935);
or U45243 (N_45243,N_44574,N_44806);
nand U45244 (N_45244,N_43093,N_42621);
nor U45245 (N_45245,N_42899,N_43226);
xnor U45246 (N_45246,N_43903,N_43821);
nor U45247 (N_45247,N_42935,N_44933);
or U45248 (N_45248,N_44367,N_42541);
and U45249 (N_45249,N_43810,N_44330);
and U45250 (N_45250,N_44107,N_43196);
nand U45251 (N_45251,N_44987,N_42716);
nor U45252 (N_45252,N_43454,N_42896);
or U45253 (N_45253,N_44378,N_42832);
or U45254 (N_45254,N_43696,N_43594);
and U45255 (N_45255,N_42806,N_42711);
nand U45256 (N_45256,N_43624,N_44813);
nor U45257 (N_45257,N_44983,N_43249);
or U45258 (N_45258,N_44582,N_43415);
xor U45259 (N_45259,N_42848,N_43653);
nand U45260 (N_45260,N_44048,N_43869);
nand U45261 (N_45261,N_44648,N_43690);
and U45262 (N_45262,N_43050,N_42954);
nor U45263 (N_45263,N_44278,N_43407);
or U45264 (N_45264,N_44486,N_44292);
nor U45265 (N_45265,N_43071,N_44104);
xor U45266 (N_45266,N_43431,N_42545);
nor U45267 (N_45267,N_44616,N_44266);
and U45268 (N_45268,N_44456,N_43061);
nor U45269 (N_45269,N_44289,N_44008);
nand U45270 (N_45270,N_42884,N_43480);
nand U45271 (N_45271,N_44428,N_42590);
nand U45272 (N_45272,N_44044,N_43612);
nor U45273 (N_45273,N_44055,N_43889);
or U45274 (N_45274,N_42635,N_43269);
and U45275 (N_45275,N_43432,N_43391);
and U45276 (N_45276,N_44258,N_44943);
nor U45277 (N_45277,N_44508,N_44915);
nor U45278 (N_45278,N_43443,N_44236);
xor U45279 (N_45279,N_44757,N_44645);
or U45280 (N_45280,N_43721,N_43187);
nand U45281 (N_45281,N_43574,N_44100);
nor U45282 (N_45282,N_42904,N_43776);
and U45283 (N_45283,N_44838,N_44653);
nor U45284 (N_45284,N_42519,N_44361);
nand U45285 (N_45285,N_42658,N_43229);
and U45286 (N_45286,N_43149,N_43403);
nor U45287 (N_45287,N_44803,N_44808);
and U45288 (N_45288,N_42688,N_44206);
nand U45289 (N_45289,N_44141,N_44991);
nor U45290 (N_45290,N_44453,N_44411);
nor U45291 (N_45291,N_44062,N_44490);
xnor U45292 (N_45292,N_43418,N_42926);
nand U45293 (N_45293,N_42811,N_44858);
or U45294 (N_45294,N_44734,N_43915);
xor U45295 (N_45295,N_44631,N_43705);
or U45296 (N_45296,N_44392,N_44239);
xnor U45297 (N_45297,N_43227,N_44495);
nand U45298 (N_45298,N_44730,N_44632);
nand U45299 (N_45299,N_44090,N_44203);
nor U45300 (N_45300,N_44707,N_43114);
nand U45301 (N_45301,N_43254,N_43430);
or U45302 (N_45302,N_42671,N_44810);
nor U45303 (N_45303,N_43863,N_43421);
nor U45304 (N_45304,N_42709,N_43289);
or U45305 (N_45305,N_43133,N_44021);
nor U45306 (N_45306,N_43392,N_42860);
or U45307 (N_45307,N_42697,N_44249);
and U45308 (N_45308,N_43890,N_43586);
nand U45309 (N_45309,N_43835,N_43009);
xor U45310 (N_45310,N_43593,N_43369);
and U45311 (N_45311,N_44922,N_42733);
or U45312 (N_45312,N_43764,N_43053);
xnor U45313 (N_45313,N_43657,N_43395);
nor U45314 (N_45314,N_44768,N_42618);
xor U45315 (N_45315,N_42841,N_43255);
xnor U45316 (N_45316,N_43761,N_43830);
or U45317 (N_45317,N_43950,N_44856);
nor U45318 (N_45318,N_44474,N_43885);
or U45319 (N_45319,N_42537,N_43783);
xor U45320 (N_45320,N_43183,N_44385);
and U45321 (N_45321,N_44333,N_43433);
nand U45322 (N_45322,N_44345,N_43563);
xor U45323 (N_45323,N_44060,N_44144);
nor U45324 (N_45324,N_44136,N_44799);
nor U45325 (N_45325,N_44654,N_43601);
and U45326 (N_45326,N_44982,N_42789);
xnor U45327 (N_45327,N_44560,N_43828);
xnor U45328 (N_45328,N_42738,N_42611);
nor U45329 (N_45329,N_44079,N_43888);
xor U45330 (N_45330,N_44432,N_42962);
xnor U45331 (N_45331,N_43352,N_44609);
nand U45332 (N_45332,N_43957,N_44923);
xor U45333 (N_45333,N_43662,N_44690);
xnor U45334 (N_45334,N_43843,N_42773);
nand U45335 (N_45335,N_44466,N_44231);
xor U45336 (N_45336,N_44182,N_42744);
nand U45337 (N_45337,N_43752,N_44878);
nor U45338 (N_45338,N_42776,N_42760);
xnor U45339 (N_45339,N_44192,N_42869);
xor U45340 (N_45340,N_44303,N_43853);
nor U45341 (N_45341,N_42749,N_44015);
and U45342 (N_45342,N_44597,N_44823);
xor U45343 (N_45343,N_43509,N_43092);
xor U45344 (N_45344,N_42943,N_44007);
and U45345 (N_45345,N_44088,N_44454);
or U45346 (N_45346,N_43176,N_44314);
or U45347 (N_45347,N_44171,N_42571);
nor U45348 (N_45348,N_42814,N_43503);
nor U45349 (N_45349,N_43655,N_44095);
xor U45350 (N_45350,N_44888,N_44547);
nor U45351 (N_45351,N_44520,N_44714);
nor U45352 (N_45352,N_44769,N_42762);
xnor U45353 (N_45353,N_43451,N_42548);
or U45354 (N_45354,N_44037,N_43158);
nand U45355 (N_45355,N_44059,N_42589);
nand U45356 (N_45356,N_42694,N_44792);
or U45357 (N_45357,N_43782,N_43470);
or U45358 (N_45358,N_43656,N_44506);
xor U45359 (N_45359,N_44845,N_44153);
or U45360 (N_45360,N_43145,N_43939);
nor U45361 (N_45361,N_43506,N_43780);
and U45362 (N_45362,N_43019,N_44591);
nand U45363 (N_45363,N_42802,N_43800);
or U45364 (N_45364,N_43047,N_42952);
nand U45365 (N_45365,N_43734,N_43572);
or U45366 (N_45366,N_43270,N_44290);
xnor U45367 (N_45367,N_43051,N_44369);
xor U45368 (N_45368,N_42939,N_43166);
xor U45369 (N_45369,N_43893,N_44644);
or U45370 (N_45370,N_43945,N_42784);
nand U45371 (N_45371,N_43074,N_44900);
or U45372 (N_45372,N_43801,N_43684);
or U45373 (N_45373,N_43493,N_44318);
and U45374 (N_45374,N_42704,N_44628);
and U45375 (N_45375,N_44480,N_43217);
and U45376 (N_45376,N_42865,N_44642);
xor U45377 (N_45377,N_43606,N_43279);
xor U45378 (N_45378,N_43706,N_43735);
nor U45379 (N_45379,N_43566,N_44788);
xor U45380 (N_45380,N_43303,N_43946);
xnor U45381 (N_45381,N_42647,N_44967);
and U45382 (N_45382,N_42633,N_44944);
and U45383 (N_45383,N_42523,N_44219);
nand U45384 (N_45384,N_43209,N_43930);
nor U45385 (N_45385,N_43536,N_43283);
nor U45386 (N_45386,N_43688,N_44646);
nor U45387 (N_45387,N_43686,N_42564);
nor U45388 (N_45388,N_43294,N_44729);
nor U45389 (N_45389,N_43195,N_43521);
nand U45390 (N_45390,N_43355,N_44470);
nor U45391 (N_45391,N_44599,N_43918);
xnor U45392 (N_45392,N_42964,N_44825);
nand U45393 (N_45393,N_42728,N_44296);
and U45394 (N_45394,N_44637,N_42970);
nor U45395 (N_45395,N_44601,N_44353);
nor U45396 (N_45396,N_43923,N_43274);
and U45397 (N_45397,N_43032,N_42741);
xor U45398 (N_45398,N_43023,N_43512);
nand U45399 (N_45399,N_44424,N_44742);
nor U45400 (N_45400,N_43630,N_43550);
or U45401 (N_45401,N_43661,N_44140);
xor U45402 (N_45402,N_43580,N_44930);
and U45403 (N_45403,N_43100,N_44627);
or U45404 (N_45404,N_43170,N_43867);
nand U45405 (N_45405,N_44876,N_42859);
xor U45406 (N_45406,N_44307,N_43685);
or U45407 (N_45407,N_44094,N_43876);
and U45408 (N_45408,N_43152,N_43747);
xor U45409 (N_45409,N_44886,N_44526);
nand U45410 (N_45410,N_43766,N_43072);
and U45411 (N_45411,N_44573,N_43295);
or U45412 (N_45412,N_42967,N_43789);
or U45413 (N_45413,N_44833,N_42922);
xor U45414 (N_45414,N_43880,N_43216);
or U45415 (N_45415,N_44535,N_43124);
nor U45416 (N_45416,N_43589,N_44351);
and U45417 (N_45417,N_42539,N_43386);
nand U45418 (N_45418,N_42629,N_43084);
nor U45419 (N_45419,N_44862,N_43608);
and U45420 (N_45420,N_44414,N_43907);
xnor U45421 (N_45421,N_43839,N_42916);
and U45422 (N_45422,N_44158,N_44879);
xor U45423 (N_45423,N_44039,N_44014);
xor U45424 (N_45424,N_42948,N_44953);
xor U45425 (N_45425,N_44431,N_42565);
or U45426 (N_45426,N_43495,N_43738);
nand U45427 (N_45427,N_44612,N_43045);
xor U45428 (N_45428,N_43374,N_43060);
or U45429 (N_45429,N_42576,N_44302);
nor U45430 (N_45430,N_44178,N_44516);
and U45431 (N_45431,N_43017,N_42903);
nor U45432 (N_45432,N_42513,N_44370);
xnor U45433 (N_45433,N_44641,N_43771);
nand U45434 (N_45434,N_43401,N_44409);
nand U45435 (N_45435,N_43381,N_44379);
nand U45436 (N_45436,N_42508,N_44965);
or U45437 (N_45437,N_42992,N_44070);
nand U45438 (N_45438,N_43035,N_44084);
xnor U45439 (N_45439,N_43492,N_44503);
or U45440 (N_45440,N_43429,N_42820);
or U45441 (N_45441,N_43440,N_44415);
nor U45442 (N_45442,N_42923,N_43538);
xor U45443 (N_45443,N_44183,N_43922);
or U45444 (N_45444,N_43938,N_42616);
or U45445 (N_45445,N_43318,N_43539);
xnor U45446 (N_45446,N_44067,N_43862);
nor U45447 (N_45447,N_43916,N_44187);
and U45448 (N_45448,N_43746,N_44819);
nand U45449 (N_45449,N_44340,N_44677);
xnor U45450 (N_45450,N_43831,N_42730);
or U45451 (N_45451,N_43313,N_43206);
nor U45452 (N_45452,N_42581,N_43972);
nor U45453 (N_45453,N_43774,N_43762);
nor U45454 (N_45454,N_43201,N_43722);
nor U45455 (N_45455,N_43438,N_43474);
and U45456 (N_45456,N_44464,N_43190);
nand U45457 (N_45457,N_43253,N_43416);
nand U45458 (N_45458,N_42975,N_44606);
or U45459 (N_45459,N_44747,N_43214);
nor U45460 (N_45460,N_43319,N_44312);
or U45461 (N_45461,N_43377,N_44200);
and U45462 (N_45462,N_43665,N_44073);
nor U45463 (N_45463,N_44626,N_42812);
nor U45464 (N_45464,N_43895,N_44342);
nor U45465 (N_45465,N_42573,N_42657);
nand U45466 (N_45466,N_43131,N_44331);
nand U45467 (N_45467,N_44636,N_42608);
and U45468 (N_45468,N_43376,N_43564);
or U45469 (N_45469,N_44745,N_43769);
nand U45470 (N_45470,N_43742,N_44873);
nand U45471 (N_45471,N_44167,N_42921);
or U45472 (N_45472,N_42845,N_44012);
and U45473 (N_45473,N_42663,N_44689);
nand U45474 (N_45474,N_44270,N_44664);
nor U45475 (N_45475,N_43827,N_44155);
nor U45476 (N_45476,N_42870,N_44404);
xnor U45477 (N_45477,N_43317,N_42990);
nor U45478 (N_45478,N_42659,N_44267);
nand U45479 (N_45479,N_44986,N_44822);
or U45480 (N_45480,N_44295,N_44118);
or U45481 (N_45481,N_42752,N_42842);
and U45482 (N_45482,N_42721,N_44981);
xor U45483 (N_45483,N_43750,N_43400);
nand U45484 (N_45484,N_44359,N_42999);
nand U45485 (N_45485,N_44798,N_44984);
nand U45486 (N_45486,N_44865,N_44610);
nand U45487 (N_45487,N_43634,N_42724);
nor U45488 (N_45488,N_43191,N_42693);
or U45489 (N_45489,N_43030,N_43846);
nor U45490 (N_45490,N_44316,N_42909);
nor U45491 (N_45491,N_44117,N_42714);
or U45492 (N_45492,N_43924,N_43977);
and U45493 (N_45493,N_43266,N_44811);
nor U45494 (N_45494,N_44096,N_43510);
and U45495 (N_45495,N_44818,N_44793);
nand U45496 (N_45496,N_44402,N_44238);
or U45497 (N_45497,N_44985,N_44386);
or U45498 (N_45498,N_43337,N_44577);
nand U45499 (N_45499,N_42790,N_43663);
nor U45500 (N_45500,N_44568,N_42817);
or U45501 (N_45501,N_44651,N_43016);
nand U45502 (N_45502,N_43054,N_44356);
and U45503 (N_45503,N_44383,N_43615);
or U45504 (N_45504,N_43147,N_43628);
or U45505 (N_45505,N_43086,N_43618);
nand U45506 (N_45506,N_44578,N_42844);
xnor U45507 (N_45507,N_43526,N_44241);
xnor U45508 (N_45508,N_44496,N_43037);
nand U45509 (N_45509,N_43457,N_43463);
or U45510 (N_45510,N_43184,N_44210);
nand U45511 (N_45511,N_44892,N_43864);
and U45512 (N_45512,N_44363,N_43426);
nand U45513 (N_45513,N_43714,N_43452);
nand U45514 (N_45514,N_44859,N_43961);
or U45515 (N_45515,N_42805,N_44684);
or U45516 (N_45516,N_44667,N_44068);
xnor U45517 (N_45517,N_43408,N_44052);
and U45518 (N_45518,N_44598,N_44450);
nor U45519 (N_45519,N_44510,N_44724);
xnor U45520 (N_45520,N_43641,N_42558);
and U45521 (N_45521,N_43366,N_42567);
and U45522 (N_45522,N_43840,N_44406);
nand U45523 (N_45523,N_43478,N_43785);
or U45524 (N_45524,N_44121,N_43523);
nand U45525 (N_45525,N_43097,N_43850);
nand U45526 (N_45526,N_44174,N_44388);
and U45527 (N_45527,N_44826,N_42900);
nand U45528 (N_45528,N_43602,N_43894);
xnor U45529 (N_45529,N_43901,N_42654);
or U45530 (N_45530,N_44305,N_42778);
xnor U45531 (N_45531,N_42604,N_43384);
or U45532 (N_45532,N_42858,N_42739);
nor U45533 (N_45533,N_42592,N_43687);
nand U45534 (N_45534,N_44228,N_43784);
nand U45535 (N_45535,N_43284,N_43469);
or U45536 (N_45536,N_44146,N_43658);
and U45537 (N_45537,N_43132,N_42597);
or U45538 (N_45538,N_44056,N_43342);
nand U45539 (N_45539,N_43561,N_44349);
xnor U45540 (N_45540,N_42886,N_44961);
or U45541 (N_45541,N_43331,N_44384);
xnor U45542 (N_45542,N_43359,N_42649);
or U45543 (N_45543,N_42885,N_43942);
xor U45544 (N_45544,N_43882,N_43067);
xnor U45545 (N_45545,N_43707,N_43728);
nand U45546 (N_45546,N_42800,N_43276);
nor U45547 (N_45547,N_43077,N_44458);
nor U45548 (N_45548,N_43062,N_43476);
and U45549 (N_45549,N_42680,N_43848);
and U45550 (N_45550,N_43994,N_44166);
nor U45551 (N_45551,N_43836,N_43417);
or U45552 (N_45552,N_43066,N_43382);
xnor U45553 (N_45553,N_44805,N_43180);
nor U45554 (N_45554,N_44539,N_43816);
nor U45555 (N_45555,N_44467,N_44932);
xor U45556 (N_45556,N_44035,N_42665);
nor U45557 (N_45557,N_43410,N_43065);
nand U45558 (N_45558,N_43327,N_44198);
nand U45559 (N_45559,N_44442,N_43763);
xnor U45560 (N_45560,N_42609,N_44509);
xnor U45561 (N_45561,N_43178,N_43483);
or U45562 (N_45562,N_44942,N_43231);
xor U45563 (N_45563,N_44579,N_44416);
nand U45564 (N_45564,N_44026,N_42521);
nand U45565 (N_45565,N_44759,N_43263);
nand U45566 (N_45566,N_42905,N_44003);
or U45567 (N_45567,N_43955,N_42725);
or U45568 (N_45568,N_43194,N_44213);
and U45569 (N_45569,N_43031,N_43046);
xor U45570 (N_45570,N_43315,N_42750);
nor U45571 (N_45571,N_42772,N_44229);
nor U45572 (N_45572,N_43832,N_44168);
nand U45573 (N_45573,N_42620,N_44306);
nor U45574 (N_45574,N_44410,N_43179);
or U45575 (N_45575,N_44829,N_42840);
xor U45576 (N_45576,N_43291,N_43716);
and U45577 (N_45577,N_43456,N_44243);
and U45578 (N_45578,N_43034,N_44740);
nand U45579 (N_45579,N_42867,N_42557);
nand U45580 (N_45580,N_43242,N_44732);
nand U45581 (N_45581,N_43765,N_42612);
and U45582 (N_45582,N_44753,N_44691);
xor U45583 (N_45583,N_43585,N_44122);
nand U45584 (N_45584,N_44465,N_43013);
nand U45585 (N_45585,N_44024,N_44973);
and U45586 (N_45586,N_44899,N_44901);
and U45587 (N_45587,N_44253,N_43379);
and U45588 (N_45588,N_43091,N_44254);
and U45589 (N_45589,N_44400,N_44978);
nand U45590 (N_45590,N_43600,N_43645);
nand U45591 (N_45591,N_44925,N_44038);
nor U45592 (N_45592,N_44031,N_43936);
xor U45593 (N_45593,N_44584,N_42510);
xnor U45594 (N_45594,N_42661,N_43489);
nor U45595 (N_45595,N_44695,N_43394);
nor U45596 (N_45596,N_44780,N_44658);
xor U45597 (N_45597,N_43434,N_42580);
or U45598 (N_45598,N_44963,N_42757);
nand U45599 (N_45599,N_42763,N_43874);
nand U45600 (N_45600,N_43198,N_43360);
or U45601 (N_45601,N_43101,N_43258);
nor U45602 (N_45602,N_43135,N_44727);
and U45603 (N_45603,N_43157,N_44590);
nand U45604 (N_45604,N_43823,N_43937);
xnor U45605 (N_45605,N_43625,N_42626);
nor U45606 (N_45606,N_43638,N_43144);
or U45607 (N_45607,N_43259,N_44502);
nor U45608 (N_45608,N_42700,N_42852);
nand U45609 (N_45609,N_43396,N_44782);
xnor U45610 (N_45610,N_42632,N_44920);
xnor U45611 (N_45611,N_44857,N_44904);
xnor U45612 (N_45612,N_44710,N_44413);
and U45613 (N_45613,N_43837,N_43292);
xnor U45614 (N_45614,N_42644,N_44575);
nor U45615 (N_45615,N_43309,N_44517);
or U45616 (N_45616,N_44098,N_43301);
xor U45617 (N_45617,N_42664,N_44870);
xnor U45618 (N_45618,N_43680,N_42882);
nand U45619 (N_45619,N_43250,N_42824);
or U45620 (N_45620,N_43052,N_43277);
xnor U45621 (N_45621,N_43859,N_44103);
or U45622 (N_45622,N_43020,N_42717);
nor U45623 (N_45623,N_43999,N_44752);
xor U45624 (N_45624,N_42615,N_43507);
nor U45625 (N_45625,N_43751,N_44807);
and U45626 (N_45626,N_43163,N_43420);
nor U45627 (N_45627,N_44180,N_43727);
nand U45628 (N_45628,N_44188,N_44002);
xnor U45629 (N_45629,N_44726,N_42522);
or U45630 (N_45630,N_44230,N_43620);
nand U45631 (N_45631,N_43482,N_44719);
xor U45632 (N_45632,N_43515,N_42971);
nor U45633 (N_45633,N_44071,N_44844);
xnor U45634 (N_45634,N_42771,N_43679);
nand U45635 (N_45635,N_44891,N_43861);
xnor U45636 (N_45636,N_43501,N_43570);
or U45637 (N_45637,N_43675,N_43791);
nor U45638 (N_45638,N_44928,N_44321);
and U45639 (N_45639,N_43385,N_43271);
nor U45640 (N_45640,N_44374,N_43960);
nand U45641 (N_45641,N_43335,N_44693);
or U45642 (N_45642,N_42731,N_43243);
nand U45643 (N_45643,N_42946,N_43998);
or U45644 (N_45644,N_43632,N_43010);
and U45645 (N_45645,N_42794,N_42682);
and U45646 (N_45646,N_43508,N_43635);
and U45647 (N_45647,N_43151,N_44447);
xor U45648 (N_45648,N_42669,N_43648);
nor U45649 (N_45649,N_43683,N_43592);
nand U45650 (N_45650,N_43678,N_44864);
and U45651 (N_45651,N_44285,N_43005);
and U45652 (N_45652,N_42906,N_44116);
nor U45653 (N_45653,N_43790,N_44789);
nand U45654 (N_45654,N_43857,N_44968);
and U45655 (N_45655,N_44540,N_44861);
nand U45656 (N_45656,N_44308,N_44478);
xnor U45657 (N_45657,N_44723,N_44077);
xor U45658 (N_45658,N_44519,N_43344);
nand U45659 (N_45659,N_42504,N_44309);
xor U45660 (N_45660,N_43069,N_42755);
nand U45661 (N_45661,N_44421,N_43595);
or U45662 (N_45662,N_42656,N_44018);
xor U45663 (N_45663,N_44785,N_44248);
nand U45664 (N_45664,N_43803,N_43571);
nor U45665 (N_45665,N_44663,N_44222);
nand U45666 (N_45666,N_43753,N_42606);
and U45667 (N_45667,N_42568,N_44602);
and U45668 (N_45668,N_44119,N_43348);
xnor U45669 (N_45669,N_44754,N_42873);
or U45670 (N_45670,N_42614,N_44425);
nand U45671 (N_45671,N_42546,N_42910);
nand U45672 (N_45672,N_44998,N_44134);
and U45673 (N_45673,N_44783,N_43324);
xor U45674 (N_45674,N_44418,N_44551);
xor U45675 (N_45675,N_43349,N_44074);
nor U45676 (N_45676,N_43312,N_42808);
nand U45677 (N_45677,N_44232,N_42818);
xnor U45678 (N_45678,N_44449,N_43724);
nor U45679 (N_45679,N_44929,N_44699);
and U45680 (N_45680,N_44473,N_43558);
nor U45681 (N_45681,N_44294,N_44286);
nand U45682 (N_45682,N_43905,N_42779);
nand U45683 (N_45683,N_44934,N_43361);
nor U45684 (N_45684,N_42945,N_42681);
or U45685 (N_45685,N_44683,N_44767);
xor U45686 (N_45686,N_43177,N_44064);
nand U45687 (N_45687,N_42827,N_44498);
xor U45688 (N_45688,N_44380,N_43479);
nor U45689 (N_45689,N_43623,N_43346);
or U45690 (N_45690,N_44214,N_44160);
nand U45691 (N_45691,N_43940,N_43904);
and U45692 (N_45692,N_43056,N_43484);
and U45693 (N_45693,N_43555,N_43697);
nand U45694 (N_45694,N_42996,N_44608);
xnor U45695 (N_45695,N_42719,N_44974);
nor U45696 (N_45696,N_44401,N_44518);
and U45697 (N_45697,N_42524,N_44828);
xnor U45698 (N_45698,N_43787,N_44471);
xnor U45699 (N_45699,N_44816,N_44279);
or U45700 (N_45700,N_43590,N_43952);
xnor U45701 (N_45701,N_43218,N_42973);
nor U45702 (N_45702,N_42624,N_43806);
nand U45703 (N_45703,N_42610,N_44208);
xor U45704 (N_45704,N_43175,N_44194);
xnor U45705 (N_45705,N_43272,N_44957);
or U45706 (N_45706,N_44507,N_43181);
and U45707 (N_45707,N_42668,N_42816);
and U45708 (N_45708,N_44435,N_43496);
nand U45709 (N_45709,N_42983,N_44227);
nand U45710 (N_45710,N_44556,N_43841);
and U45711 (N_45711,N_44053,N_42854);
or U45712 (N_45712,N_44523,N_42619);
or U45713 (N_45713,N_43043,N_44919);
xor U45714 (N_45714,N_44427,N_42607);
or U45715 (N_45715,N_43098,N_42974);
nor U45716 (N_45716,N_44544,N_44281);
xnor U45717 (N_45717,N_43311,N_44777);
or U45718 (N_45718,N_43105,N_43228);
nand U45719 (N_45719,N_44940,N_44335);
nand U45720 (N_45720,N_43587,N_44448);
xor U45721 (N_45721,N_44849,N_42628);
nand U45722 (N_45722,N_44357,N_42894);
xnor U45723 (N_45723,N_44894,N_43213);
xor U45724 (N_45724,N_43304,N_44697);
xnor U45725 (N_45725,N_43537,N_42652);
nand U45726 (N_45726,N_44958,N_44299);
xor U45727 (N_45727,N_44310,N_44226);
xor U45728 (N_45728,N_44840,N_44956);
nor U45729 (N_45729,N_44440,N_44170);
nand U45730 (N_45730,N_42708,N_44311);
xnor U45731 (N_45731,N_43991,N_43519);
nor U45732 (N_45732,N_43472,N_44921);
or U45733 (N_45733,N_44162,N_44781);
nor U45734 (N_45734,N_43730,N_42501);
nand U45735 (N_45735,N_43729,N_43219);
nor U45736 (N_45736,N_44809,N_44439);
or U45737 (N_45737,N_43205,N_43756);
nand U45738 (N_45738,N_44851,N_42622);
nor U45739 (N_45739,N_42998,N_43811);
nor U45740 (N_45740,N_43511,N_44476);
xnor U45741 (N_45741,N_44504,N_44364);
nand U45742 (N_45742,N_44868,N_42807);
nor U45743 (N_45743,N_42907,N_44586);
xor U45744 (N_45744,N_43103,N_44625);
and U45745 (N_45745,N_42825,N_44513);
or U45746 (N_45746,N_43567,N_43112);
xor U45747 (N_45747,N_44703,N_42917);
or U45748 (N_45748,N_44669,N_43116);
xor U45749 (N_45749,N_42627,N_44438);
and U45750 (N_45750,N_44939,N_43712);
or U45751 (N_45751,N_43168,N_43740);
nand U45752 (N_45752,N_43073,N_43085);
nand U45753 (N_45753,N_42925,N_44534);
and U45754 (N_45754,N_44106,N_44197);
and U45755 (N_45755,N_42696,N_43490);
xor U45756 (N_45756,N_44784,N_43200);
nor U45757 (N_45757,N_44477,N_43424);
or U45758 (N_45758,N_44086,N_44884);
nand U45759 (N_45759,N_44772,N_44887);
nand U45760 (N_45760,N_43979,N_43122);
and U45761 (N_45761,N_44288,N_43995);
nor U45762 (N_45762,N_44051,N_42570);
xor U45763 (N_45763,N_44895,N_44854);
and U45764 (N_45764,N_44172,N_43252);
or U45765 (N_45765,N_44533,N_43978);
or U45766 (N_45766,N_44101,N_43399);
xnor U45767 (N_45767,N_42929,N_42857);
and U45768 (N_45768,N_44487,N_42809);
nor U45769 (N_45769,N_43708,N_44538);
and U45770 (N_45770,N_43793,N_43797);
nand U45771 (N_45771,N_42520,N_44615);
nor U45772 (N_45772,N_43667,N_44045);
xnor U45773 (N_45773,N_44685,N_43225);
or U45774 (N_45774,N_44137,N_43441);
and U45775 (N_45775,N_44135,N_44976);
and U45776 (N_45776,N_42986,N_44528);
or U45777 (N_45777,N_43887,N_44455);
xor U45778 (N_45778,N_44365,N_43287);
xnor U45779 (N_45779,N_44163,N_44820);
xor U45780 (N_45780,N_43011,N_42793);
or U45781 (N_45781,N_43881,N_43966);
nand U45782 (N_45782,N_43475,N_44043);
nand U45783 (N_45783,N_43954,N_43435);
nand U45784 (N_45784,N_42535,N_42579);
and U45785 (N_45785,N_43692,N_43090);
nand U45786 (N_45786,N_43965,N_43405);
or U45787 (N_45787,N_42798,N_43980);
xor U45788 (N_45788,N_44323,N_44399);
nor U45789 (N_45789,N_44366,N_43262);
xnor U45790 (N_45790,N_44237,N_42871);
or U45791 (N_45791,N_44755,N_44110);
and U45792 (N_45792,N_44488,N_42968);
and U45793 (N_45793,N_43514,N_44537);
nor U45794 (N_45794,N_44962,N_43189);
nand U45795 (N_45795,N_44735,N_43908);
nand U45796 (N_45796,N_42691,N_44758);
and U45797 (N_45797,N_43261,N_44327);
or U45798 (N_45798,N_44629,N_42891);
or U45799 (N_45799,N_44687,N_43603);
or U45800 (N_45800,N_42768,N_42927);
nor U45801 (N_45801,N_44246,N_43182);
or U45802 (N_45802,N_43126,N_42588);
nor U45803 (N_45803,N_44131,N_42835);
and U45804 (N_45804,N_43953,N_43909);
nand U45805 (N_45805,N_42930,N_44536);
and U45806 (N_45806,N_44570,N_44546);
nand U45807 (N_45807,N_42912,N_44511);
xnor U45808 (N_45808,N_44675,N_43445);
and U45809 (N_45809,N_44199,N_44164);
and U45810 (N_45810,N_43963,N_42743);
nor U45811 (N_45811,N_44341,N_44988);
nor U45812 (N_45812,N_44483,N_44874);
or U45813 (N_45813,N_43247,N_44678);
nand U45814 (N_45814,N_44893,N_44492);
or U45815 (N_45815,N_43057,N_44138);
nor U45816 (N_45816,N_43860,N_43676);
and U45817 (N_45817,N_42687,N_44563);
or U45818 (N_45818,N_44033,N_42897);
nor U45819 (N_45819,N_43286,N_42958);
or U45820 (N_45820,N_44959,N_44329);
or U45821 (N_45821,N_43798,N_42651);
xnor U45822 (N_45822,N_44751,N_43238);
nand U45823 (N_45823,N_43854,N_44047);
nor U45824 (N_45824,N_44834,N_43375);
or U45825 (N_45825,N_43591,N_44924);
nand U45826 (N_45826,N_42861,N_43530);
or U45827 (N_45827,N_44739,N_44611);
xor U45828 (N_45828,N_44259,N_43969);
or U45829 (N_45829,N_44006,N_43902);
or U45830 (N_45830,N_43499,N_44355);
and U45831 (N_45831,N_43351,N_43007);
xnor U45832 (N_45832,N_42689,N_44681);
xor U45833 (N_45833,N_44429,N_42705);
xnor U45834 (N_45834,N_44850,N_44224);
or U45835 (N_45835,N_44089,N_43328);
and U45836 (N_45836,N_44527,N_42502);
or U45837 (N_45837,N_42582,N_43674);
xor U45838 (N_45838,N_44949,N_44004);
or U45839 (N_45839,N_44656,N_43777);
nand U45840 (N_45840,N_43450,N_42613);
and U45841 (N_45841,N_42594,N_43870);
or U45842 (N_45842,N_44682,N_43036);
nand U45843 (N_45843,N_44408,N_43578);
xnor U45844 (N_45844,N_42710,N_43544);
xor U45845 (N_45845,N_44770,N_43164);
or U45846 (N_45846,N_43234,N_42572);
or U45847 (N_45847,N_44830,N_44566);
and U45848 (N_45848,N_44061,N_44522);
nor U45849 (N_45849,N_43212,N_43248);
nand U45850 (N_45850,N_44423,N_42720);
nand U45851 (N_45851,N_43542,N_43654);
and U45852 (N_45852,N_44469,N_44054);
or U45853 (N_45853,N_44860,N_43367);
and U45854 (N_45854,N_44148,N_43044);
nand U45855 (N_45855,N_43398,N_44087);
and U45856 (N_45856,N_43720,N_43925);
nand U45857 (N_45857,N_43079,N_44655);
xnor U45858 (N_45858,N_43669,N_42801);
nor U45859 (N_45859,N_43741,N_44994);
nor U45860 (N_45860,N_43868,N_43121);
nand U45861 (N_45861,N_42877,N_44161);
nor U45862 (N_45862,N_43532,N_44766);
and U45863 (N_45863,N_42828,N_43160);
xnor U45864 (N_45864,N_43280,N_42932);
xor U45865 (N_45865,N_42505,N_44273);
nor U45866 (N_45866,N_42679,N_43083);
nor U45867 (N_45867,N_42642,N_43754);
nand U45868 (N_45868,N_43604,N_42506);
or U45869 (N_45869,N_43817,N_42960);
nand U45870 (N_45870,N_43719,N_42706);
nand U45871 (N_45871,N_43146,N_44903);
xnor U45872 (N_45872,N_43677,N_44652);
nor U45873 (N_45873,N_43970,N_44926);
or U45874 (N_45874,N_43380,N_43643);
xor U45875 (N_45875,N_43723,N_44670);
xor U45876 (N_45876,N_43110,N_43080);
and U45877 (N_45877,N_43818,N_42553);
or U45878 (N_45878,N_43033,N_42949);
or U45879 (N_45879,N_42595,N_44207);
xor U45880 (N_45880,N_43388,N_44553);
nand U45881 (N_45881,N_42544,N_42646);
or U45882 (N_45882,N_43650,N_42920);
xor U45883 (N_45883,N_44620,N_44554);
nor U45884 (N_45884,N_42723,N_43106);
or U45885 (N_45885,N_44177,N_42770);
nor U45886 (N_45886,N_43964,N_44204);
xor U45887 (N_45887,N_43583,N_44970);
nor U45888 (N_45888,N_44257,N_42833);
nand U45889 (N_45889,N_43001,N_42530);
or U45890 (N_45890,N_42965,N_43082);
xor U45891 (N_45891,N_44128,N_44298);
nand U45892 (N_45892,N_44338,N_43237);
and U45893 (N_45893,N_44890,N_44265);
xnor U45894 (N_45894,N_42586,N_43668);
and U45895 (N_45895,N_43282,N_42585);
and U45896 (N_45896,N_44129,N_42944);
nor U45897 (N_45897,N_42978,N_44555);
or U45898 (N_45898,N_44130,N_43148);
and U45899 (N_45899,N_42774,N_42551);
and U45900 (N_45900,N_44422,N_43767);
or U45901 (N_45901,N_43293,N_42853);
or U45902 (N_45902,N_43875,N_43370);
nand U45903 (N_45903,N_43826,N_44948);
nand U45904 (N_45904,N_44036,N_43129);
xor U45905 (N_45905,N_43244,N_43598);
nor U45906 (N_45906,N_42766,N_43522);
nand U45907 (N_45907,N_43673,N_44017);
nand U45908 (N_45908,N_42525,N_44791);
or U45909 (N_45909,N_43813,N_42780);
nand U45910 (N_45910,N_43636,N_43468);
xor U45911 (N_45911,N_42837,N_44756);
nor U45912 (N_45912,N_44142,N_43281);
or U45913 (N_45913,N_44205,N_44019);
nand U45914 (N_45914,N_43340,N_44744);
or U45915 (N_45915,N_42796,N_42953);
nand U45916 (N_45916,N_44936,N_44328);
nand U45917 (N_45917,N_42695,N_44376);
and U45918 (N_45918,N_44350,N_44271);
or U45919 (N_45919,N_43897,N_44344);
or U45920 (N_45920,N_42660,N_43533);
nor U45921 (N_45921,N_44132,N_44115);
or U45922 (N_45922,N_42575,N_42692);
nand U45923 (N_45923,N_44127,N_42549);
nand U45924 (N_45924,N_42713,N_44877);
xnor U45925 (N_45925,N_43022,N_44063);
nand U45926 (N_45926,N_43851,N_42829);
or U45927 (N_45927,N_42881,N_43505);
and U45928 (N_45928,N_43799,N_44133);
or U45929 (N_45929,N_42555,N_44814);
or U45930 (N_45930,N_44541,N_44264);
and U45931 (N_45931,N_43302,N_43967);
or U45932 (N_45932,N_43310,N_43557);
nand U45933 (N_45933,N_42799,N_43140);
or U45934 (N_45934,N_42878,N_43524);
xnor U45935 (N_45935,N_44196,N_43442);
nand U45936 (N_45936,N_42847,N_42804);
nor U45937 (N_45937,N_44867,N_43173);
nor U45938 (N_45938,N_44221,N_44542);
nand U45939 (N_45939,N_43597,N_44889);
nor U45940 (N_45940,N_43617,N_44482);
nand U45941 (N_45941,N_43371,N_43596);
xor U45942 (N_45942,N_43899,N_43659);
or U45943 (N_45943,N_44332,N_44337);
nand U45944 (N_45944,N_44728,N_43699);
or U45945 (N_45945,N_42577,N_43865);
and U45946 (N_45946,N_44176,N_43781);
or U45947 (N_45947,N_43824,N_44287);
xnor U45948 (N_45948,N_43099,N_44698);
or U45949 (N_45949,N_43581,N_44339);
nor U45950 (N_45950,N_43387,N_43744);
nand U45951 (N_45951,N_44368,N_43517);
xnor U45952 (N_45952,N_43856,N_43932);
or U45953 (N_45953,N_43356,N_43232);
or U45954 (N_45954,N_44293,N_42898);
or U45955 (N_45955,N_44564,N_44277);
or U45956 (N_45956,N_44885,N_43343);
nand U45957 (N_45957,N_44185,N_43627);
nand U45958 (N_45958,N_44082,N_44898);
and U45959 (N_45959,N_44152,N_43439);
and U45960 (N_45960,N_44112,N_42819);
xor U45961 (N_45961,N_43477,N_42742);
xnor U45962 (N_45962,N_44459,N_44081);
and U45963 (N_45963,N_43884,N_44358);
nand U45964 (N_45964,N_44405,N_44773);
nand U45965 (N_45965,N_42821,N_43786);
nand U45966 (N_45966,N_44165,N_44846);
and U45967 (N_45967,N_43251,N_43185);
nor U45968 (N_45968,N_43136,N_43575);
or U45969 (N_45969,N_44634,N_44672);
xnor U45970 (N_45970,N_44561,N_42777);
xor U45971 (N_45971,N_43285,N_44979);
and U45972 (N_45972,N_43552,N_43913);
nor U45973 (N_45973,N_43906,N_43773);
xor U45974 (N_45974,N_43795,N_43599);
xnor U45975 (N_45975,N_44603,N_44567);
xor U45976 (N_45976,N_43926,N_43120);
xor U45977 (N_45977,N_43819,N_43345);
nor U45978 (N_45978,N_43220,N_44097);
or U45979 (N_45979,N_43737,N_44883);
or U45980 (N_45980,N_44475,N_44869);
xnor U45981 (N_45981,N_43088,N_42826);
nor U45982 (N_45982,N_43778,N_43012);
and U45983 (N_45983,N_42783,N_44235);
xnor U45984 (N_45984,N_44215,N_42638);
xor U45985 (N_45985,N_43444,N_44191);
and U45986 (N_45986,N_43404,N_44853);
nand U45987 (N_45987,N_44748,N_43569);
and U45988 (N_45988,N_43504,N_44525);
nor U45989 (N_45989,N_44113,N_44159);
xnor U45990 (N_45990,N_42566,N_44175);
nand U45991 (N_45991,N_43584,N_44494);
nand U45992 (N_45992,N_42767,N_43353);
nand U45993 (N_45993,N_44099,N_43174);
nor U45994 (N_45994,N_43075,N_44407);
and U45995 (N_45995,N_42956,N_44721);
nand U45996 (N_45996,N_43834,N_44659);
or U45997 (N_45997,N_44343,N_43471);
xnor U45998 (N_45998,N_42518,N_43670);
or U45999 (N_45999,N_44852,N_43138);
xor U46000 (N_46000,N_42662,N_44046);
nand U46001 (N_46001,N_44647,N_43855);
or U46002 (N_46002,N_43235,N_44532);
xnor U46003 (N_46003,N_43815,N_44969);
or U46004 (N_46004,N_43562,N_43297);
nand U46005 (N_46005,N_42655,N_43025);
or U46006 (N_46006,N_44635,N_43221);
or U46007 (N_46007,N_44600,N_43494);
nand U46008 (N_46008,N_43681,N_42674);
nor U46009 (N_46009,N_44916,N_42736);
nand U46010 (N_46010,N_44080,N_43804);
and U46011 (N_46011,N_42648,N_44149);
nand U46012 (N_46012,N_43162,N_44346);
nand U46013 (N_46013,N_44848,N_44382);
nor U46014 (N_46014,N_44543,N_42699);
xnor U46015 (N_46015,N_43024,N_44233);
and U46016 (N_46016,N_42791,N_43829);
or U46017 (N_46017,N_42690,N_43167);
xnor U46018 (N_46018,N_42883,N_44765);
and U46019 (N_46019,N_43265,N_43912);
nand U46020 (N_46020,N_42969,N_44034);
nand U46021 (N_46021,N_42751,N_44836);
nor U46022 (N_46022,N_43070,N_44481);
or U46023 (N_46023,N_44245,N_44831);
nand U46024 (N_46024,N_44897,N_42729);
nand U46025 (N_46025,N_42529,N_42889);
nand U46026 (N_46026,N_44123,N_43165);
xnor U46027 (N_46027,N_44242,N_42995);
nand U46028 (N_46028,N_43807,N_43448);
nand U46029 (N_46029,N_43113,N_43956);
and U46030 (N_46030,N_43703,N_42507);
or U46031 (N_46031,N_44855,N_43055);
or U46032 (N_46032,N_44022,N_43006);
nor U46033 (N_46033,N_43362,N_44479);
or U46034 (N_46034,N_43622,N_43871);
nor U46035 (N_46035,N_42788,N_43357);
or U46036 (N_46036,N_42887,N_44173);
and U46037 (N_46037,N_43760,N_44945);
xnor U46038 (N_46038,N_42512,N_43736);
and U46039 (N_46039,N_43014,N_43996);
and U46040 (N_46040,N_44420,N_43364);
nand U46041 (N_46041,N_42754,N_43320);
and U46042 (N_46042,N_44301,N_42947);
or U46043 (N_46043,N_44125,N_44881);
nand U46044 (N_46044,N_44102,N_42895);
nand U46045 (N_46045,N_42623,N_44065);
and U46046 (N_46046,N_42797,N_43406);
or U46047 (N_46047,N_44372,N_44169);
nor U46048 (N_46048,N_44741,N_42987);
and U46049 (N_46049,N_43487,N_43118);
xnor U46050 (N_46050,N_44225,N_44941);
and U46051 (N_46051,N_44317,N_42993);
or U46052 (N_46052,N_43749,N_43437);
or U46053 (N_46053,N_43959,N_42980);
or U46054 (N_46054,N_43171,N_43717);
xor U46055 (N_46055,N_43701,N_43027);
nor U46056 (N_46056,N_44688,N_43971);
nor U46057 (N_46057,N_43486,N_43534);
nand U46058 (N_46058,N_44223,N_44444);
or U46059 (N_46059,N_44394,N_44716);
nor U46060 (N_46060,N_43947,N_44980);
and U46061 (N_46061,N_43997,N_43172);
nor U46062 (N_46062,N_43516,N_43543);
xnor U46063 (N_46063,N_42547,N_42936);
nand U46064 (N_46064,N_44717,N_44975);
or U46065 (N_46065,N_44558,N_42722);
nor U46066 (N_46066,N_43192,N_42550);
and U46067 (N_46067,N_44120,N_44320);
xor U46068 (N_46068,N_42554,N_43693);
or U46069 (N_46069,N_44218,N_42503);
xnor U46070 (N_46070,N_44016,N_44075);
or U46071 (N_46071,N_42963,N_44154);
xnor U46072 (N_46072,N_42672,N_44300);
xor U46073 (N_46073,N_43491,N_43197);
nor U46074 (N_46074,N_44576,N_44795);
xor U46075 (N_46075,N_43973,N_43540);
and U46076 (N_46076,N_44377,N_43929);
or U46077 (N_46077,N_44692,N_44696);
nand U46078 (N_46078,N_43664,N_44764);
or U46079 (N_46079,N_42758,N_43239);
or U46080 (N_46080,N_44209,N_43560);
xor U46081 (N_46081,N_42782,N_44815);
nand U46082 (N_46082,N_43700,N_44032);
or U46083 (N_46083,N_44521,N_42737);
or U46084 (N_46084,N_42941,N_43390);
and U46085 (N_46085,N_44091,N_43159);
xor U46086 (N_46086,N_43461,N_42972);
xor U46087 (N_46087,N_44863,N_42830);
xor U46088 (N_46088,N_43616,N_44297);
xor U46089 (N_46089,N_44837,N_43161);
xnor U46090 (N_46090,N_43142,N_42630);
xor U46091 (N_46091,N_43063,N_43878);
and U46092 (N_46092,N_43267,N_43428);
nand U46093 (N_46093,N_42598,N_44706);
and U46094 (N_46094,N_44841,N_42533);
or U46095 (N_46095,N_42893,N_42748);
or U46096 (N_46096,N_44725,N_44313);
nor U46097 (N_46097,N_42625,N_43933);
xnor U46098 (N_46098,N_42584,N_43652);
nor U46099 (N_46099,N_43985,N_44436);
and U46100 (N_46100,N_42740,N_44720);
or U46101 (N_46101,N_43528,N_44468);
nor U46102 (N_46102,N_43436,N_43812);
nor U46103 (N_46103,N_44412,N_43064);
nor U46104 (N_46104,N_44671,N_43920);
nor U46105 (N_46105,N_43018,N_43556);
nand U46106 (N_46106,N_43646,N_44030);
nand U46107 (N_46107,N_42599,N_44272);
and U46108 (N_46108,N_44952,N_44605);
nor U46109 (N_46109,N_44661,N_43347);
nor U46110 (N_46110,N_42785,N_42715);
xor U46111 (N_46111,N_42560,N_43156);
and U46112 (N_46112,N_44571,N_43931);
xnor U46113 (N_46113,N_43814,N_44794);
nand U46114 (N_46114,N_44662,N_43040);
nor U46115 (N_46115,N_42676,N_43833);
xor U46116 (N_46116,N_44092,N_43378);
nor U46117 (N_46117,N_44437,N_42994);
and U46118 (N_46118,N_42686,N_44025);
or U46119 (N_46119,N_44737,N_43153);
xnor U46120 (N_46120,N_43873,N_43886);
or U46121 (N_46121,N_42634,N_43096);
nor U46122 (N_46122,N_44255,N_44592);
nand U46123 (N_46123,N_43268,N_43193);
nand U46124 (N_46124,N_42851,N_44484);
nand U46125 (N_46125,N_43866,N_42988);
or U46126 (N_46126,N_44955,N_43314);
xor U46127 (N_46127,N_44673,N_43230);
xor U46128 (N_46128,N_42938,N_44650);
or U46129 (N_46129,N_43306,N_43076);
or U46130 (N_46130,N_43927,N_44913);
and U46131 (N_46131,N_44776,N_44426);
and U46132 (N_46132,N_44790,N_44005);
or U46133 (N_46133,N_42666,N_43695);
and U46134 (N_46134,N_43241,N_44040);
nand U46135 (N_46135,N_44360,N_44269);
xor U46136 (N_46136,N_42775,N_43914);
nor U46137 (N_46137,N_43535,N_44010);
nor U46138 (N_46138,N_43104,N_44715);
nor U46139 (N_46139,N_43518,N_43548);
and U46140 (N_46140,N_44800,N_43048);
nor U46141 (N_46141,N_44639,N_44722);
nor U46142 (N_46142,N_44960,N_44334);
xnor U46143 (N_46143,N_43466,N_44896);
nand U46144 (N_46144,N_43898,N_44489);
nor U46145 (N_46145,N_43672,N_43246);
xor U46146 (N_46146,N_43488,N_44550);
nor U46147 (N_46147,N_43541,N_42563);
xor U46148 (N_46148,N_43021,N_43316);
nor U46149 (N_46149,N_44354,N_42531);
or U46150 (N_46150,N_42984,N_42538);
xor U46151 (N_46151,N_43130,N_44396);
nand U46152 (N_46152,N_44996,N_44093);
nand U46153 (N_46153,N_44596,N_43393);
or U46154 (N_46154,N_43002,N_44910);
nand U46155 (N_46155,N_44076,N_43921);
nand U46156 (N_46156,N_42703,N_44607);
xnor U46157 (N_46157,N_44572,N_43726);
or U46158 (N_46158,N_42872,N_44244);
xnor U46159 (N_46159,N_43757,N_44589);
and U46160 (N_46160,N_43768,N_42511);
and U46161 (N_46161,N_43460,N_42976);
nor U46162 (N_46162,N_43414,N_44195);
xor U46163 (N_46163,N_42961,N_43992);
nand U46164 (N_46164,N_43582,N_42849);
nor U46165 (N_46165,N_42746,N_44738);
nand U46166 (N_46166,N_44842,N_42792);
xor U46167 (N_46167,N_43900,N_44524);
xnor U46168 (N_46168,N_43660,N_44371);
and U46169 (N_46169,N_44145,N_42982);
or U46170 (N_46170,N_44872,N_44775);
or U46171 (N_46171,N_42745,N_43257);
and U46172 (N_46172,N_44666,N_44679);
or U46173 (N_46173,N_44618,N_44393);
nor U46174 (N_46174,N_42591,N_43990);
or U46175 (N_46175,N_43139,N_43278);
nor U46176 (N_46176,N_44562,N_44565);
nor U46177 (N_46177,N_43691,N_43453);
nor U46178 (N_46178,N_44762,N_43802);
xor U46179 (N_46179,N_42540,N_42600);
nor U46180 (N_46180,N_42890,N_44643);
xor U46181 (N_46181,N_44736,N_44835);
and U46182 (N_46182,N_42678,N_44434);
xnor U46183 (N_46183,N_42759,N_44514);
xnor U46184 (N_46184,N_42839,N_43842);
nor U46185 (N_46185,N_43413,N_42868);
nor U46186 (N_46186,N_42933,N_43204);
or U46187 (N_46187,N_42985,N_43150);
xor U46188 (N_46188,N_43689,N_44622);
nand U46189 (N_46189,N_42951,N_44763);
xor U46190 (N_46190,N_44731,N_42675);
nor U46191 (N_46191,N_42726,N_44375);
or U46192 (N_46192,N_43264,N_43520);
nand U46193 (N_46193,N_42934,N_44617);
xor U46194 (N_46194,N_44252,N_43465);
xnor U46195 (N_46195,N_43123,N_44451);
nor U46196 (N_46196,N_44569,N_43619);
xor U46197 (N_46197,N_44011,N_42641);
xnor U46198 (N_46198,N_44029,N_43788);
xnor U46199 (N_46199,N_44640,N_43772);
or U46200 (N_46200,N_44832,N_42836);
xnor U46201 (N_46201,N_44108,N_44604);
nand U46202 (N_46202,N_43808,N_42587);
xor U46203 (N_46203,N_44847,N_43500);
nand U46204 (N_46204,N_44284,N_44069);
xor U46205 (N_46205,N_43389,N_43288);
and U46206 (N_46206,N_44275,N_44668);
nor U46207 (N_46207,N_42734,N_43354);
nor U46208 (N_46208,N_43671,N_43644);
xnor U46209 (N_46209,N_44072,N_43637);
nand U46210 (N_46210,N_44460,N_44151);
or U46211 (N_46211,N_44325,N_43745);
nor U46212 (N_46212,N_42732,N_43858);
or U46213 (N_46213,N_44595,N_43078);
and U46214 (N_46214,N_44463,N_44462);
nor U46215 (N_46215,N_43879,N_43958);
nand U46216 (N_46216,N_44189,N_43710);
and U46217 (N_46217,N_42813,N_44276);
nor U46218 (N_46218,N_44179,N_42957);
nand U46219 (N_46219,N_44997,N_44548);
xor U46220 (N_46220,N_43365,N_44882);
and U46221 (N_46221,N_43847,N_44827);
nand U46222 (N_46222,N_43718,N_43260);
xnor U46223 (N_46223,N_43211,N_43029);
nand U46224 (N_46224,N_43363,N_44709);
nor U46225 (N_46225,N_44917,N_44250);
nand U46226 (N_46226,N_42795,N_44013);
and U46227 (N_46227,N_43809,N_43409);
xor U46228 (N_46228,N_43941,N_44373);
or U46229 (N_46229,N_44906,N_44797);
xor U46230 (N_46230,N_43554,N_42924);
xor U46231 (N_46231,N_43559,N_43568);
xnor U46232 (N_46232,N_43911,N_43775);
and U46233 (N_46233,N_44009,N_44485);
nand U46234 (N_46234,N_43579,N_44614);
nand U46235 (N_46235,N_42601,N_42532);
xnor U46236 (N_46236,N_42834,N_42761);
or U46237 (N_46237,N_44397,N_43731);
xnor U46238 (N_46238,N_43993,N_44217);
nand U46239 (N_46239,N_42846,N_42977);
nor U46240 (N_46240,N_44694,N_43910);
nand U46241 (N_46241,N_43042,N_43968);
or U46242 (N_46242,N_42815,N_43236);
and U46243 (N_46243,N_44927,N_43207);
xnor U46244 (N_46244,N_42605,N_43613);
nor U46245 (N_46245,N_43102,N_42864);
xor U46246 (N_46246,N_44156,N_44274);
and U46247 (N_46247,N_43003,N_42901);
nor U46248 (N_46248,N_44804,N_43422);
nand U46249 (N_46249,N_44581,N_44937);
or U46250 (N_46250,N_42791,N_43147);
or U46251 (N_46251,N_42948,N_42734);
nand U46252 (N_46252,N_43925,N_44913);
and U46253 (N_46253,N_42577,N_42688);
xor U46254 (N_46254,N_43080,N_43277);
or U46255 (N_46255,N_43020,N_43563);
xnor U46256 (N_46256,N_42946,N_42698);
and U46257 (N_46257,N_44357,N_43554);
and U46258 (N_46258,N_44312,N_42640);
and U46259 (N_46259,N_43626,N_44566);
or U46260 (N_46260,N_43907,N_44397);
or U46261 (N_46261,N_44866,N_43367);
nor U46262 (N_46262,N_44867,N_43167);
and U46263 (N_46263,N_43276,N_43196);
nand U46264 (N_46264,N_43462,N_43643);
xor U46265 (N_46265,N_44339,N_43746);
nor U46266 (N_46266,N_43043,N_44457);
or U46267 (N_46267,N_43581,N_42991);
xnor U46268 (N_46268,N_44595,N_43488);
nand U46269 (N_46269,N_44085,N_42567);
and U46270 (N_46270,N_42644,N_42978);
and U46271 (N_46271,N_44589,N_43514);
nor U46272 (N_46272,N_42663,N_43013);
nor U46273 (N_46273,N_44523,N_42627);
nand U46274 (N_46274,N_44752,N_43895);
and U46275 (N_46275,N_43197,N_42831);
nand U46276 (N_46276,N_44855,N_44070);
xor U46277 (N_46277,N_44846,N_44233);
nor U46278 (N_46278,N_42941,N_44799);
xor U46279 (N_46279,N_44520,N_44226);
xnor U46280 (N_46280,N_43632,N_42855);
or U46281 (N_46281,N_44042,N_44404);
xor U46282 (N_46282,N_42924,N_43075);
xor U46283 (N_46283,N_44381,N_43460);
or U46284 (N_46284,N_44139,N_42633);
nor U46285 (N_46285,N_43456,N_43999);
nor U46286 (N_46286,N_44573,N_44261);
and U46287 (N_46287,N_42503,N_43489);
xor U46288 (N_46288,N_44077,N_42929);
or U46289 (N_46289,N_43614,N_42765);
xor U46290 (N_46290,N_43598,N_44949);
or U46291 (N_46291,N_43809,N_43915);
or U46292 (N_46292,N_43957,N_42664);
nand U46293 (N_46293,N_43278,N_42936);
or U46294 (N_46294,N_44244,N_44544);
and U46295 (N_46295,N_44096,N_44451);
and U46296 (N_46296,N_43289,N_42757);
or U46297 (N_46297,N_44320,N_43215);
xor U46298 (N_46298,N_43650,N_44883);
and U46299 (N_46299,N_44278,N_44149);
nand U46300 (N_46300,N_43561,N_44280);
and U46301 (N_46301,N_44295,N_43410);
nand U46302 (N_46302,N_43183,N_43114);
or U46303 (N_46303,N_43873,N_42895);
and U46304 (N_46304,N_42593,N_44222);
xor U46305 (N_46305,N_44573,N_43721);
or U46306 (N_46306,N_44509,N_42722);
nor U46307 (N_46307,N_44177,N_43116);
and U46308 (N_46308,N_43091,N_42561);
xor U46309 (N_46309,N_44723,N_44696);
and U46310 (N_46310,N_44950,N_44289);
nor U46311 (N_46311,N_44845,N_42884);
nand U46312 (N_46312,N_44433,N_43820);
nor U46313 (N_46313,N_44948,N_44975);
and U46314 (N_46314,N_44675,N_44539);
xnor U46315 (N_46315,N_43494,N_43685);
and U46316 (N_46316,N_44272,N_42906);
xnor U46317 (N_46317,N_44123,N_43147);
or U46318 (N_46318,N_44533,N_42995);
nor U46319 (N_46319,N_44322,N_43241);
xnor U46320 (N_46320,N_43209,N_42688);
and U46321 (N_46321,N_43687,N_44051);
xor U46322 (N_46322,N_43960,N_43410);
nor U46323 (N_46323,N_44863,N_44541);
xor U46324 (N_46324,N_42537,N_44576);
nand U46325 (N_46325,N_43060,N_42591);
nand U46326 (N_46326,N_43225,N_43429);
and U46327 (N_46327,N_44678,N_43644);
and U46328 (N_46328,N_44195,N_44531);
nor U46329 (N_46329,N_44860,N_44460);
nor U46330 (N_46330,N_43059,N_43442);
xor U46331 (N_46331,N_43078,N_44043);
or U46332 (N_46332,N_44769,N_42794);
nand U46333 (N_46333,N_43050,N_43528);
and U46334 (N_46334,N_42606,N_43243);
and U46335 (N_46335,N_43865,N_43682);
and U46336 (N_46336,N_42522,N_44092);
nand U46337 (N_46337,N_44069,N_44306);
xnor U46338 (N_46338,N_44801,N_43156);
and U46339 (N_46339,N_43466,N_44176);
or U46340 (N_46340,N_43019,N_42944);
and U46341 (N_46341,N_43047,N_44453);
nand U46342 (N_46342,N_44183,N_43289);
nor U46343 (N_46343,N_43613,N_44787);
or U46344 (N_46344,N_43314,N_44397);
or U46345 (N_46345,N_44738,N_44589);
and U46346 (N_46346,N_42693,N_44483);
nand U46347 (N_46347,N_44521,N_42878);
and U46348 (N_46348,N_43357,N_42933);
or U46349 (N_46349,N_43122,N_43433);
nor U46350 (N_46350,N_43424,N_43784);
xor U46351 (N_46351,N_43276,N_43607);
nor U46352 (N_46352,N_42818,N_42613);
nand U46353 (N_46353,N_44481,N_44245);
nand U46354 (N_46354,N_42939,N_43670);
and U46355 (N_46355,N_43818,N_44531);
nand U46356 (N_46356,N_44657,N_43595);
nand U46357 (N_46357,N_42999,N_43652);
and U46358 (N_46358,N_43807,N_43994);
xnor U46359 (N_46359,N_43916,N_44047);
xor U46360 (N_46360,N_43415,N_44722);
or U46361 (N_46361,N_44884,N_42886);
or U46362 (N_46362,N_44676,N_44138);
xnor U46363 (N_46363,N_43665,N_42766);
xor U46364 (N_46364,N_43291,N_42625);
nor U46365 (N_46365,N_44946,N_44516);
and U46366 (N_46366,N_43439,N_42518);
xor U46367 (N_46367,N_42923,N_44620);
and U46368 (N_46368,N_43507,N_44430);
nor U46369 (N_46369,N_44583,N_43497);
or U46370 (N_46370,N_44229,N_43467);
and U46371 (N_46371,N_44471,N_43198);
or U46372 (N_46372,N_44539,N_44749);
xnor U46373 (N_46373,N_43647,N_42862);
xnor U46374 (N_46374,N_42867,N_42694);
nor U46375 (N_46375,N_42905,N_44105);
or U46376 (N_46376,N_44544,N_43458);
and U46377 (N_46377,N_44416,N_44884);
and U46378 (N_46378,N_44906,N_42834);
xnor U46379 (N_46379,N_43123,N_44485);
or U46380 (N_46380,N_42609,N_44427);
and U46381 (N_46381,N_43952,N_43644);
nand U46382 (N_46382,N_44451,N_44704);
nor U46383 (N_46383,N_43217,N_44392);
nand U46384 (N_46384,N_42531,N_44081);
or U46385 (N_46385,N_44375,N_42695);
nand U46386 (N_46386,N_44985,N_43125);
nor U46387 (N_46387,N_44601,N_44273);
or U46388 (N_46388,N_42838,N_43134);
and U46389 (N_46389,N_42932,N_44254);
or U46390 (N_46390,N_44278,N_44462);
nor U46391 (N_46391,N_44365,N_43735);
nor U46392 (N_46392,N_44538,N_44381);
nand U46393 (N_46393,N_43213,N_44313);
and U46394 (N_46394,N_44419,N_43720);
nand U46395 (N_46395,N_43452,N_43118);
xnor U46396 (N_46396,N_44290,N_42801);
xnor U46397 (N_46397,N_44063,N_43052);
nor U46398 (N_46398,N_43230,N_43191);
xnor U46399 (N_46399,N_43105,N_44120);
or U46400 (N_46400,N_43307,N_44585);
xnor U46401 (N_46401,N_43234,N_42985);
nor U46402 (N_46402,N_43103,N_43673);
or U46403 (N_46403,N_43870,N_43427);
nor U46404 (N_46404,N_44219,N_43768);
nor U46405 (N_46405,N_44969,N_43117);
nor U46406 (N_46406,N_44886,N_44091);
nor U46407 (N_46407,N_44177,N_43219);
xnor U46408 (N_46408,N_42882,N_44077);
nor U46409 (N_46409,N_42689,N_43246);
or U46410 (N_46410,N_43988,N_44543);
nor U46411 (N_46411,N_43647,N_44514);
and U46412 (N_46412,N_44789,N_43849);
nand U46413 (N_46413,N_42571,N_43203);
nor U46414 (N_46414,N_43417,N_42961);
or U46415 (N_46415,N_44230,N_44759);
and U46416 (N_46416,N_43924,N_43858);
nor U46417 (N_46417,N_44859,N_42817);
nand U46418 (N_46418,N_43698,N_44692);
xnor U46419 (N_46419,N_44367,N_44325);
nor U46420 (N_46420,N_43683,N_43340);
nor U46421 (N_46421,N_43962,N_42776);
nor U46422 (N_46422,N_44245,N_44214);
and U46423 (N_46423,N_44486,N_43055);
nor U46424 (N_46424,N_43174,N_44191);
and U46425 (N_46425,N_44092,N_43640);
nand U46426 (N_46426,N_43922,N_44827);
nand U46427 (N_46427,N_43482,N_43631);
and U46428 (N_46428,N_42630,N_42770);
xor U46429 (N_46429,N_43404,N_42909);
xnor U46430 (N_46430,N_44878,N_42815);
nor U46431 (N_46431,N_43188,N_43986);
or U46432 (N_46432,N_44230,N_43202);
nand U46433 (N_46433,N_43613,N_42681);
and U46434 (N_46434,N_44097,N_44988);
xor U46435 (N_46435,N_42996,N_44946);
or U46436 (N_46436,N_42710,N_43855);
nand U46437 (N_46437,N_43347,N_44275);
and U46438 (N_46438,N_43511,N_44427);
or U46439 (N_46439,N_43913,N_44294);
or U46440 (N_46440,N_42561,N_42697);
nor U46441 (N_46441,N_44271,N_43843);
nor U46442 (N_46442,N_44262,N_43765);
xnor U46443 (N_46443,N_44314,N_43683);
xnor U46444 (N_46444,N_42546,N_42659);
nor U46445 (N_46445,N_44329,N_43320);
nor U46446 (N_46446,N_42555,N_43927);
xnor U46447 (N_46447,N_44675,N_43206);
and U46448 (N_46448,N_44412,N_43094);
xor U46449 (N_46449,N_44395,N_43589);
or U46450 (N_46450,N_42604,N_44518);
and U46451 (N_46451,N_42580,N_44906);
and U46452 (N_46452,N_43731,N_43872);
nor U46453 (N_46453,N_43024,N_42847);
and U46454 (N_46454,N_43798,N_44571);
nand U46455 (N_46455,N_42699,N_44561);
and U46456 (N_46456,N_43777,N_44892);
xnor U46457 (N_46457,N_44067,N_42723);
nand U46458 (N_46458,N_44088,N_43994);
or U46459 (N_46459,N_44074,N_43073);
nand U46460 (N_46460,N_44427,N_44729);
or U46461 (N_46461,N_44242,N_43004);
or U46462 (N_46462,N_43496,N_43411);
or U46463 (N_46463,N_44828,N_42729);
xor U46464 (N_46464,N_42950,N_42686);
and U46465 (N_46465,N_43785,N_44008);
nor U46466 (N_46466,N_42953,N_44041);
or U46467 (N_46467,N_43542,N_42973);
nor U46468 (N_46468,N_43741,N_43439);
or U46469 (N_46469,N_42558,N_44494);
and U46470 (N_46470,N_43906,N_44426);
and U46471 (N_46471,N_44561,N_42851);
xor U46472 (N_46472,N_43460,N_44076);
nor U46473 (N_46473,N_43547,N_43595);
and U46474 (N_46474,N_42648,N_42905);
or U46475 (N_46475,N_43068,N_44969);
and U46476 (N_46476,N_43641,N_44648);
nor U46477 (N_46477,N_43237,N_42649);
and U46478 (N_46478,N_44995,N_42541);
nand U46479 (N_46479,N_44725,N_43714);
xnor U46480 (N_46480,N_44093,N_44438);
and U46481 (N_46481,N_42817,N_43939);
xnor U46482 (N_46482,N_43447,N_44356);
nand U46483 (N_46483,N_43665,N_43315);
nand U46484 (N_46484,N_44355,N_42910);
xor U46485 (N_46485,N_43175,N_44245);
or U46486 (N_46486,N_44179,N_43201);
xnor U46487 (N_46487,N_43094,N_42666);
nand U46488 (N_46488,N_44673,N_42743);
xor U46489 (N_46489,N_43028,N_43704);
nand U46490 (N_46490,N_43127,N_44502);
nand U46491 (N_46491,N_44588,N_43887);
or U46492 (N_46492,N_42597,N_44096);
nor U46493 (N_46493,N_44165,N_42993);
xnor U46494 (N_46494,N_44608,N_42861);
xnor U46495 (N_46495,N_43854,N_43439);
or U46496 (N_46496,N_42902,N_44460);
or U46497 (N_46497,N_44363,N_44348);
nand U46498 (N_46498,N_44868,N_42916);
nand U46499 (N_46499,N_43564,N_43834);
nor U46500 (N_46500,N_43634,N_44073);
or U46501 (N_46501,N_44267,N_44305);
nor U46502 (N_46502,N_43537,N_44097);
nor U46503 (N_46503,N_42660,N_44754);
or U46504 (N_46504,N_42512,N_42716);
nor U46505 (N_46505,N_42769,N_44721);
nor U46506 (N_46506,N_43352,N_43269);
xor U46507 (N_46507,N_44232,N_43048);
nand U46508 (N_46508,N_42668,N_42769);
nand U46509 (N_46509,N_43699,N_43848);
nor U46510 (N_46510,N_44682,N_43690);
and U46511 (N_46511,N_42702,N_42552);
nor U46512 (N_46512,N_43639,N_43685);
nor U46513 (N_46513,N_44177,N_44158);
and U46514 (N_46514,N_44877,N_43112);
nand U46515 (N_46515,N_43073,N_43414);
nand U46516 (N_46516,N_43104,N_44760);
nor U46517 (N_46517,N_43080,N_44562);
xnor U46518 (N_46518,N_43882,N_44760);
nor U46519 (N_46519,N_44604,N_43949);
and U46520 (N_46520,N_44217,N_43403);
and U46521 (N_46521,N_44115,N_43344);
nand U46522 (N_46522,N_44255,N_43188);
xnor U46523 (N_46523,N_42812,N_44445);
and U46524 (N_46524,N_44252,N_44861);
or U46525 (N_46525,N_43296,N_42826);
xnor U46526 (N_46526,N_42536,N_43168);
nand U46527 (N_46527,N_44576,N_43066);
xnor U46528 (N_46528,N_43987,N_44719);
nor U46529 (N_46529,N_43814,N_43730);
or U46530 (N_46530,N_42913,N_44045);
nand U46531 (N_46531,N_43947,N_43483);
or U46532 (N_46532,N_44545,N_42929);
nand U46533 (N_46533,N_44861,N_44402);
nor U46534 (N_46534,N_43842,N_43956);
nand U46535 (N_46535,N_42995,N_44722);
or U46536 (N_46536,N_43038,N_43084);
nand U46537 (N_46537,N_43705,N_42745);
nor U46538 (N_46538,N_43402,N_42864);
xor U46539 (N_46539,N_43316,N_43019);
or U46540 (N_46540,N_43907,N_43100);
and U46541 (N_46541,N_43534,N_44035);
and U46542 (N_46542,N_43289,N_42671);
nand U46543 (N_46543,N_43428,N_42987);
and U46544 (N_46544,N_44301,N_43603);
nor U46545 (N_46545,N_43920,N_44153);
nand U46546 (N_46546,N_44972,N_44367);
or U46547 (N_46547,N_44908,N_44559);
nand U46548 (N_46548,N_44434,N_44759);
and U46549 (N_46549,N_44283,N_42826);
and U46550 (N_46550,N_42906,N_42641);
or U46551 (N_46551,N_44440,N_43529);
xor U46552 (N_46552,N_43768,N_44478);
nand U46553 (N_46553,N_42585,N_44569);
nand U46554 (N_46554,N_43335,N_43898);
and U46555 (N_46555,N_44133,N_44989);
or U46556 (N_46556,N_42764,N_44188);
nor U46557 (N_46557,N_43283,N_44584);
and U46558 (N_46558,N_43801,N_42756);
xnor U46559 (N_46559,N_44415,N_43481);
nand U46560 (N_46560,N_44546,N_44571);
xnor U46561 (N_46561,N_43385,N_43147);
nor U46562 (N_46562,N_44002,N_42735);
nand U46563 (N_46563,N_44266,N_44554);
xor U46564 (N_46564,N_44326,N_43201);
nor U46565 (N_46565,N_42663,N_44621);
and U46566 (N_46566,N_42827,N_43122);
xor U46567 (N_46567,N_44264,N_44941);
or U46568 (N_46568,N_43115,N_43512);
and U46569 (N_46569,N_42512,N_44417);
nor U46570 (N_46570,N_44093,N_43103);
and U46571 (N_46571,N_42969,N_43919);
xnor U46572 (N_46572,N_44942,N_43888);
nand U46573 (N_46573,N_44106,N_43699);
xnor U46574 (N_46574,N_43348,N_42690);
or U46575 (N_46575,N_44251,N_43226);
xor U46576 (N_46576,N_44357,N_42758);
xnor U46577 (N_46577,N_44502,N_43762);
nor U46578 (N_46578,N_43193,N_42988);
and U46579 (N_46579,N_43885,N_44150);
nor U46580 (N_46580,N_43422,N_43741);
nand U46581 (N_46581,N_43250,N_44419);
or U46582 (N_46582,N_43254,N_42944);
nor U46583 (N_46583,N_42522,N_43549);
and U46584 (N_46584,N_43822,N_43703);
and U46585 (N_46585,N_43980,N_44563);
and U46586 (N_46586,N_42727,N_44235);
or U46587 (N_46587,N_43881,N_42924);
nor U46588 (N_46588,N_44893,N_43759);
nor U46589 (N_46589,N_44534,N_43881);
xnor U46590 (N_46590,N_43365,N_44599);
nand U46591 (N_46591,N_44163,N_44039);
nor U46592 (N_46592,N_43137,N_43682);
nand U46593 (N_46593,N_42581,N_44830);
nand U46594 (N_46594,N_44814,N_44686);
and U46595 (N_46595,N_44969,N_44254);
xnor U46596 (N_46596,N_44002,N_43761);
and U46597 (N_46597,N_43034,N_42698);
nor U46598 (N_46598,N_42829,N_43361);
nand U46599 (N_46599,N_44161,N_43316);
or U46600 (N_46600,N_42641,N_42502);
nand U46601 (N_46601,N_44321,N_44723);
nand U46602 (N_46602,N_43961,N_44505);
nand U46603 (N_46603,N_42539,N_43284);
nand U46604 (N_46604,N_44657,N_44695);
xor U46605 (N_46605,N_43676,N_42954);
xnor U46606 (N_46606,N_43939,N_43799);
and U46607 (N_46607,N_43126,N_42702);
and U46608 (N_46608,N_44029,N_43175);
or U46609 (N_46609,N_42664,N_44757);
or U46610 (N_46610,N_44492,N_44408);
or U46611 (N_46611,N_43516,N_43171);
and U46612 (N_46612,N_42751,N_44819);
and U46613 (N_46613,N_44065,N_43498);
xor U46614 (N_46614,N_44638,N_43842);
nand U46615 (N_46615,N_44045,N_44918);
nor U46616 (N_46616,N_44824,N_44563);
or U46617 (N_46617,N_42551,N_44057);
and U46618 (N_46618,N_44190,N_44996);
nor U46619 (N_46619,N_44380,N_44592);
nand U46620 (N_46620,N_43677,N_42831);
xnor U46621 (N_46621,N_42917,N_44635);
xor U46622 (N_46622,N_42842,N_44286);
xor U46623 (N_46623,N_42856,N_43950);
nor U46624 (N_46624,N_44230,N_44265);
xor U46625 (N_46625,N_44170,N_44930);
and U46626 (N_46626,N_43183,N_44571);
or U46627 (N_46627,N_43466,N_43342);
xor U46628 (N_46628,N_43077,N_42873);
xor U46629 (N_46629,N_44885,N_44956);
or U46630 (N_46630,N_44616,N_43464);
nand U46631 (N_46631,N_42841,N_43623);
xor U46632 (N_46632,N_42725,N_44639);
nand U46633 (N_46633,N_42993,N_44467);
nand U46634 (N_46634,N_44999,N_44350);
or U46635 (N_46635,N_42596,N_42508);
nor U46636 (N_46636,N_43180,N_44591);
nor U46637 (N_46637,N_44253,N_44504);
nand U46638 (N_46638,N_43016,N_44689);
xor U46639 (N_46639,N_43996,N_44957);
xnor U46640 (N_46640,N_42501,N_42775);
or U46641 (N_46641,N_44845,N_42527);
or U46642 (N_46642,N_44208,N_43913);
nor U46643 (N_46643,N_42766,N_44574);
and U46644 (N_46644,N_43240,N_44516);
and U46645 (N_46645,N_44706,N_43912);
or U46646 (N_46646,N_44367,N_43265);
xnor U46647 (N_46647,N_43371,N_42924);
and U46648 (N_46648,N_44311,N_43462);
and U46649 (N_46649,N_42697,N_43840);
nand U46650 (N_46650,N_44716,N_44756);
or U46651 (N_46651,N_43750,N_43729);
and U46652 (N_46652,N_44480,N_43401);
and U46653 (N_46653,N_44918,N_44708);
nand U46654 (N_46654,N_44405,N_43280);
nand U46655 (N_46655,N_42954,N_43254);
nor U46656 (N_46656,N_42630,N_44696);
nand U46657 (N_46657,N_43526,N_43201);
and U46658 (N_46658,N_44223,N_44787);
nor U46659 (N_46659,N_42958,N_42892);
xor U46660 (N_46660,N_44451,N_42874);
and U46661 (N_46661,N_44196,N_44577);
nor U46662 (N_46662,N_43905,N_44468);
nor U46663 (N_46663,N_44168,N_42675);
nor U46664 (N_46664,N_44019,N_44596);
nor U46665 (N_46665,N_44550,N_44793);
nor U46666 (N_46666,N_43075,N_44809);
xor U46667 (N_46667,N_42622,N_44037);
or U46668 (N_46668,N_44101,N_44045);
or U46669 (N_46669,N_43552,N_44119);
nand U46670 (N_46670,N_44785,N_42789);
and U46671 (N_46671,N_44819,N_43613);
nand U46672 (N_46672,N_43281,N_43696);
or U46673 (N_46673,N_42663,N_44940);
or U46674 (N_46674,N_43075,N_43045);
nand U46675 (N_46675,N_43995,N_43444);
nor U46676 (N_46676,N_43296,N_43201);
nor U46677 (N_46677,N_43632,N_43062);
or U46678 (N_46678,N_43394,N_43705);
nor U46679 (N_46679,N_44067,N_44336);
and U46680 (N_46680,N_43388,N_43611);
nor U46681 (N_46681,N_43046,N_44401);
or U46682 (N_46682,N_44565,N_42916);
and U46683 (N_46683,N_44059,N_42703);
and U46684 (N_46684,N_44304,N_44934);
and U46685 (N_46685,N_42970,N_42973);
and U46686 (N_46686,N_43550,N_43988);
nand U46687 (N_46687,N_42577,N_44746);
xor U46688 (N_46688,N_43200,N_42664);
xnor U46689 (N_46689,N_43274,N_44312);
nor U46690 (N_46690,N_43415,N_43879);
and U46691 (N_46691,N_42937,N_42626);
nor U46692 (N_46692,N_42673,N_43467);
or U46693 (N_46693,N_43019,N_42788);
nor U46694 (N_46694,N_42885,N_44381);
and U46695 (N_46695,N_43425,N_43076);
nor U46696 (N_46696,N_42713,N_43580);
nor U46697 (N_46697,N_42597,N_44161);
nor U46698 (N_46698,N_44683,N_43807);
nand U46699 (N_46699,N_43915,N_43806);
xor U46700 (N_46700,N_44785,N_42769);
xnor U46701 (N_46701,N_43398,N_44464);
nor U46702 (N_46702,N_43400,N_43551);
and U46703 (N_46703,N_44200,N_43363);
and U46704 (N_46704,N_42913,N_44824);
nor U46705 (N_46705,N_44987,N_44431);
xor U46706 (N_46706,N_44988,N_43717);
nor U46707 (N_46707,N_42953,N_43036);
nor U46708 (N_46708,N_42934,N_44600);
and U46709 (N_46709,N_44914,N_44892);
xnor U46710 (N_46710,N_42994,N_44393);
xnor U46711 (N_46711,N_43067,N_43818);
xnor U46712 (N_46712,N_44604,N_43002);
and U46713 (N_46713,N_42999,N_43389);
and U46714 (N_46714,N_42760,N_44889);
and U46715 (N_46715,N_42766,N_44247);
and U46716 (N_46716,N_44280,N_44500);
nor U46717 (N_46717,N_43518,N_44562);
nor U46718 (N_46718,N_43860,N_43351);
and U46719 (N_46719,N_42712,N_43712);
xor U46720 (N_46720,N_44252,N_44540);
and U46721 (N_46721,N_43229,N_44833);
and U46722 (N_46722,N_42637,N_44104);
and U46723 (N_46723,N_44063,N_44599);
and U46724 (N_46724,N_42584,N_44976);
nor U46725 (N_46725,N_44368,N_44040);
nor U46726 (N_46726,N_44483,N_42880);
and U46727 (N_46727,N_42645,N_42757);
nand U46728 (N_46728,N_43003,N_44172);
nor U46729 (N_46729,N_44908,N_43411);
and U46730 (N_46730,N_42942,N_44773);
nand U46731 (N_46731,N_42855,N_42978);
and U46732 (N_46732,N_42946,N_43122);
or U46733 (N_46733,N_43513,N_42979);
nand U46734 (N_46734,N_44938,N_42662);
nand U46735 (N_46735,N_44123,N_43359);
nor U46736 (N_46736,N_44914,N_43171);
xor U46737 (N_46737,N_44581,N_42895);
xnor U46738 (N_46738,N_42753,N_43224);
nor U46739 (N_46739,N_44412,N_44382);
nand U46740 (N_46740,N_44411,N_43636);
nand U46741 (N_46741,N_44033,N_43523);
nor U46742 (N_46742,N_43209,N_44427);
nand U46743 (N_46743,N_43869,N_42568);
nand U46744 (N_46744,N_43818,N_44855);
and U46745 (N_46745,N_43102,N_43296);
or U46746 (N_46746,N_43941,N_44962);
nand U46747 (N_46747,N_44647,N_44812);
or U46748 (N_46748,N_44628,N_44240);
and U46749 (N_46749,N_43662,N_44345);
xor U46750 (N_46750,N_43955,N_43548);
nand U46751 (N_46751,N_44633,N_44150);
xor U46752 (N_46752,N_44555,N_42739);
and U46753 (N_46753,N_42910,N_43741);
nand U46754 (N_46754,N_43020,N_42578);
nand U46755 (N_46755,N_44811,N_43326);
or U46756 (N_46756,N_43923,N_44917);
or U46757 (N_46757,N_42835,N_44732);
xnor U46758 (N_46758,N_43170,N_44104);
nand U46759 (N_46759,N_44210,N_43749);
nand U46760 (N_46760,N_42709,N_44469);
nor U46761 (N_46761,N_43465,N_43968);
nor U46762 (N_46762,N_43238,N_42518);
nand U46763 (N_46763,N_44884,N_42797);
and U46764 (N_46764,N_42675,N_43003);
and U46765 (N_46765,N_43361,N_43778);
or U46766 (N_46766,N_43274,N_44841);
or U46767 (N_46767,N_43807,N_44880);
nor U46768 (N_46768,N_43042,N_42684);
nor U46769 (N_46769,N_43235,N_44748);
xor U46770 (N_46770,N_43714,N_42713);
and U46771 (N_46771,N_44476,N_44436);
nand U46772 (N_46772,N_44959,N_44948);
nor U46773 (N_46773,N_44466,N_44909);
and U46774 (N_46774,N_44368,N_44405);
nor U46775 (N_46775,N_43862,N_44418);
nor U46776 (N_46776,N_43073,N_44660);
nor U46777 (N_46777,N_44357,N_42995);
nand U46778 (N_46778,N_42593,N_43822);
nand U46779 (N_46779,N_43820,N_43742);
and U46780 (N_46780,N_43504,N_44159);
nand U46781 (N_46781,N_43312,N_43273);
nor U46782 (N_46782,N_42980,N_42768);
nand U46783 (N_46783,N_43268,N_43495);
nor U46784 (N_46784,N_44188,N_44680);
or U46785 (N_46785,N_43462,N_42669);
or U46786 (N_46786,N_44479,N_42507);
nor U46787 (N_46787,N_43764,N_44985);
nor U46788 (N_46788,N_44478,N_44422);
nand U46789 (N_46789,N_42935,N_42597);
nor U46790 (N_46790,N_43724,N_44639);
and U46791 (N_46791,N_42575,N_44528);
nor U46792 (N_46792,N_42540,N_43445);
xor U46793 (N_46793,N_44737,N_43649);
and U46794 (N_46794,N_43237,N_43631);
xnor U46795 (N_46795,N_43717,N_44391);
or U46796 (N_46796,N_43725,N_43018);
nor U46797 (N_46797,N_43935,N_42800);
and U46798 (N_46798,N_43048,N_44720);
or U46799 (N_46799,N_44727,N_44075);
and U46800 (N_46800,N_43114,N_44081);
nor U46801 (N_46801,N_44458,N_44804);
and U46802 (N_46802,N_43275,N_43950);
nor U46803 (N_46803,N_44654,N_44561);
nor U46804 (N_46804,N_44166,N_43652);
and U46805 (N_46805,N_43055,N_44854);
and U46806 (N_46806,N_44600,N_44589);
xor U46807 (N_46807,N_44265,N_43046);
nand U46808 (N_46808,N_43950,N_43048);
nor U46809 (N_46809,N_42548,N_43525);
xor U46810 (N_46810,N_43590,N_44015);
xnor U46811 (N_46811,N_43191,N_43897);
xnor U46812 (N_46812,N_43870,N_43857);
xor U46813 (N_46813,N_44223,N_43534);
nor U46814 (N_46814,N_42801,N_44009);
nor U46815 (N_46815,N_44495,N_43555);
xor U46816 (N_46816,N_43538,N_43240);
nand U46817 (N_46817,N_44299,N_44509);
xor U46818 (N_46818,N_42654,N_44569);
xnor U46819 (N_46819,N_44530,N_44864);
nand U46820 (N_46820,N_44453,N_44935);
nand U46821 (N_46821,N_44214,N_44014);
and U46822 (N_46822,N_44334,N_43498);
or U46823 (N_46823,N_44332,N_43514);
or U46824 (N_46824,N_43892,N_44040);
nor U46825 (N_46825,N_44423,N_42931);
or U46826 (N_46826,N_44741,N_43369);
nor U46827 (N_46827,N_43706,N_44727);
or U46828 (N_46828,N_44329,N_43158);
nor U46829 (N_46829,N_42899,N_42637);
or U46830 (N_46830,N_43271,N_43950);
and U46831 (N_46831,N_44519,N_42652);
and U46832 (N_46832,N_44647,N_43643);
or U46833 (N_46833,N_43885,N_43738);
xnor U46834 (N_46834,N_42557,N_44885);
nand U46835 (N_46835,N_44062,N_44090);
and U46836 (N_46836,N_43245,N_44677);
or U46837 (N_46837,N_44036,N_42803);
xnor U46838 (N_46838,N_43171,N_43956);
nor U46839 (N_46839,N_44447,N_44151);
or U46840 (N_46840,N_44505,N_44546);
xor U46841 (N_46841,N_44937,N_44705);
nor U46842 (N_46842,N_44870,N_42792);
or U46843 (N_46843,N_43980,N_44687);
nand U46844 (N_46844,N_44399,N_43341);
or U46845 (N_46845,N_44426,N_42501);
or U46846 (N_46846,N_44999,N_44175);
or U46847 (N_46847,N_44827,N_43472);
or U46848 (N_46848,N_43717,N_42564);
xnor U46849 (N_46849,N_43260,N_44065);
nor U46850 (N_46850,N_43351,N_44535);
nand U46851 (N_46851,N_44218,N_44779);
nand U46852 (N_46852,N_43862,N_43577);
nor U46853 (N_46853,N_42701,N_44363);
and U46854 (N_46854,N_42668,N_44977);
or U46855 (N_46855,N_44306,N_44089);
xnor U46856 (N_46856,N_44931,N_43229);
and U46857 (N_46857,N_44946,N_42762);
and U46858 (N_46858,N_43908,N_43004);
nand U46859 (N_46859,N_44770,N_43860);
xnor U46860 (N_46860,N_43658,N_43332);
nor U46861 (N_46861,N_44891,N_43770);
nand U46862 (N_46862,N_44015,N_44217);
xor U46863 (N_46863,N_44421,N_43575);
nand U46864 (N_46864,N_42689,N_44925);
nand U46865 (N_46865,N_42596,N_43494);
and U46866 (N_46866,N_43759,N_44205);
xnor U46867 (N_46867,N_44403,N_44931);
xnor U46868 (N_46868,N_43670,N_44367);
nand U46869 (N_46869,N_44839,N_44938);
nand U46870 (N_46870,N_43044,N_43464);
nand U46871 (N_46871,N_43881,N_44997);
or U46872 (N_46872,N_43169,N_43043);
xor U46873 (N_46873,N_44217,N_43324);
nand U46874 (N_46874,N_44849,N_42778);
xnor U46875 (N_46875,N_44574,N_42833);
or U46876 (N_46876,N_44055,N_43542);
nand U46877 (N_46877,N_43467,N_43110);
xor U46878 (N_46878,N_44973,N_43906);
nor U46879 (N_46879,N_44286,N_42636);
nand U46880 (N_46880,N_44039,N_43652);
and U46881 (N_46881,N_44033,N_43099);
or U46882 (N_46882,N_42587,N_44201);
xnor U46883 (N_46883,N_44956,N_43825);
and U46884 (N_46884,N_44468,N_43903);
xor U46885 (N_46885,N_43773,N_42719);
xor U46886 (N_46886,N_42781,N_43168);
nor U46887 (N_46887,N_42828,N_43418);
nand U46888 (N_46888,N_44883,N_44844);
xor U46889 (N_46889,N_44424,N_44957);
or U46890 (N_46890,N_43069,N_42597);
or U46891 (N_46891,N_44833,N_44089);
nor U46892 (N_46892,N_43025,N_42782);
xor U46893 (N_46893,N_42763,N_43376);
or U46894 (N_46894,N_43443,N_44254);
nor U46895 (N_46895,N_42945,N_43144);
and U46896 (N_46896,N_43813,N_43964);
nor U46897 (N_46897,N_42936,N_43754);
and U46898 (N_46898,N_44143,N_44692);
nor U46899 (N_46899,N_44006,N_42933);
and U46900 (N_46900,N_42729,N_42630);
nor U46901 (N_46901,N_44454,N_43190);
and U46902 (N_46902,N_44831,N_43288);
xnor U46903 (N_46903,N_42516,N_44023);
xor U46904 (N_46904,N_44822,N_42649);
nand U46905 (N_46905,N_44850,N_43213);
xnor U46906 (N_46906,N_44951,N_44120);
xnor U46907 (N_46907,N_43993,N_44502);
nor U46908 (N_46908,N_44893,N_43469);
nor U46909 (N_46909,N_44764,N_44278);
nor U46910 (N_46910,N_43365,N_44244);
nor U46911 (N_46911,N_42638,N_43333);
xor U46912 (N_46912,N_43388,N_44089);
or U46913 (N_46913,N_42585,N_42992);
nand U46914 (N_46914,N_42687,N_42846);
xnor U46915 (N_46915,N_43380,N_44279);
xor U46916 (N_46916,N_43910,N_44672);
xnor U46917 (N_46917,N_44043,N_43002);
and U46918 (N_46918,N_43429,N_44360);
nand U46919 (N_46919,N_43648,N_43516);
and U46920 (N_46920,N_43827,N_43197);
nand U46921 (N_46921,N_44608,N_43289);
or U46922 (N_46922,N_44897,N_43296);
nand U46923 (N_46923,N_42564,N_44847);
nor U46924 (N_46924,N_44837,N_43569);
xor U46925 (N_46925,N_43199,N_44200);
and U46926 (N_46926,N_44690,N_44791);
nand U46927 (N_46927,N_43488,N_44527);
nand U46928 (N_46928,N_42963,N_44870);
nand U46929 (N_46929,N_44027,N_44920);
nor U46930 (N_46930,N_44630,N_42723);
nand U46931 (N_46931,N_42530,N_42694);
nor U46932 (N_46932,N_44782,N_42802);
nor U46933 (N_46933,N_42738,N_42505);
and U46934 (N_46934,N_43897,N_42664);
nand U46935 (N_46935,N_43893,N_44777);
and U46936 (N_46936,N_43960,N_43751);
nor U46937 (N_46937,N_43096,N_44506);
xor U46938 (N_46938,N_42762,N_42947);
and U46939 (N_46939,N_43652,N_44107);
nand U46940 (N_46940,N_42949,N_43075);
nor U46941 (N_46941,N_44256,N_44324);
nand U46942 (N_46942,N_42943,N_42685);
or U46943 (N_46943,N_44261,N_43389);
xnor U46944 (N_46944,N_44074,N_44141);
xor U46945 (N_46945,N_42835,N_43185);
and U46946 (N_46946,N_44589,N_43758);
or U46947 (N_46947,N_44363,N_43643);
xnor U46948 (N_46948,N_42525,N_43928);
xor U46949 (N_46949,N_44188,N_42726);
nor U46950 (N_46950,N_44532,N_43861);
and U46951 (N_46951,N_44830,N_44353);
or U46952 (N_46952,N_43885,N_44583);
nor U46953 (N_46953,N_43989,N_43485);
xor U46954 (N_46954,N_43113,N_42676);
xor U46955 (N_46955,N_44002,N_44951);
nor U46956 (N_46956,N_43006,N_43454);
nor U46957 (N_46957,N_43149,N_43370);
nand U46958 (N_46958,N_43596,N_43969);
nand U46959 (N_46959,N_44944,N_44374);
and U46960 (N_46960,N_44949,N_43963);
nor U46961 (N_46961,N_44535,N_42671);
and U46962 (N_46962,N_42859,N_44743);
and U46963 (N_46963,N_43040,N_42681);
nand U46964 (N_46964,N_42619,N_44620);
xor U46965 (N_46965,N_43947,N_42846);
nand U46966 (N_46966,N_43651,N_43215);
xnor U46967 (N_46967,N_42667,N_43375);
nand U46968 (N_46968,N_44456,N_43095);
nor U46969 (N_46969,N_42903,N_44945);
nor U46970 (N_46970,N_44234,N_44587);
nor U46971 (N_46971,N_44335,N_44530);
nor U46972 (N_46972,N_43200,N_42586);
nor U46973 (N_46973,N_43043,N_43917);
nor U46974 (N_46974,N_42983,N_43547);
xor U46975 (N_46975,N_43542,N_42613);
or U46976 (N_46976,N_44971,N_44357);
and U46977 (N_46977,N_44241,N_44860);
nor U46978 (N_46978,N_44892,N_43132);
and U46979 (N_46979,N_44466,N_43252);
or U46980 (N_46980,N_44194,N_44492);
xnor U46981 (N_46981,N_43052,N_43828);
nor U46982 (N_46982,N_44177,N_44265);
nor U46983 (N_46983,N_43265,N_43453);
or U46984 (N_46984,N_44746,N_43483);
xnor U46985 (N_46985,N_43242,N_43122);
nand U46986 (N_46986,N_44351,N_43401);
or U46987 (N_46987,N_44689,N_43761);
and U46988 (N_46988,N_44592,N_42706);
xnor U46989 (N_46989,N_43764,N_43933);
and U46990 (N_46990,N_43150,N_43671);
or U46991 (N_46991,N_43406,N_42669);
and U46992 (N_46992,N_43456,N_43638);
nor U46993 (N_46993,N_43090,N_43314);
xor U46994 (N_46994,N_43675,N_42975);
and U46995 (N_46995,N_43475,N_43310);
nor U46996 (N_46996,N_44721,N_43405);
or U46997 (N_46997,N_44911,N_44035);
xnor U46998 (N_46998,N_44791,N_44918);
or U46999 (N_46999,N_43299,N_43561);
xnor U47000 (N_47000,N_43028,N_44363);
xnor U47001 (N_47001,N_42788,N_44360);
xor U47002 (N_47002,N_44579,N_43647);
and U47003 (N_47003,N_42619,N_43805);
or U47004 (N_47004,N_43607,N_44995);
or U47005 (N_47005,N_43955,N_44505);
or U47006 (N_47006,N_43253,N_44192);
and U47007 (N_47007,N_44788,N_43679);
and U47008 (N_47008,N_43783,N_43862);
or U47009 (N_47009,N_43074,N_42691);
and U47010 (N_47010,N_42910,N_42725);
and U47011 (N_47011,N_43687,N_44082);
or U47012 (N_47012,N_44509,N_43362);
and U47013 (N_47013,N_42882,N_42837);
nand U47014 (N_47014,N_42814,N_43208);
xor U47015 (N_47015,N_43892,N_43233);
or U47016 (N_47016,N_43784,N_44743);
or U47017 (N_47017,N_44082,N_43192);
xor U47018 (N_47018,N_43352,N_44378);
nand U47019 (N_47019,N_43003,N_44039);
xor U47020 (N_47020,N_43391,N_44856);
nand U47021 (N_47021,N_43931,N_43411);
nor U47022 (N_47022,N_44400,N_43899);
xor U47023 (N_47023,N_44749,N_42685);
and U47024 (N_47024,N_44014,N_42634);
and U47025 (N_47025,N_44817,N_43926);
or U47026 (N_47026,N_42859,N_42957);
nor U47027 (N_47027,N_43245,N_43966);
nand U47028 (N_47028,N_44598,N_42753);
and U47029 (N_47029,N_44329,N_44912);
and U47030 (N_47030,N_44161,N_44501);
nand U47031 (N_47031,N_42844,N_42550);
xor U47032 (N_47032,N_43915,N_44419);
nor U47033 (N_47033,N_43934,N_43141);
xnor U47034 (N_47034,N_43902,N_43280);
xor U47035 (N_47035,N_44524,N_43695);
nor U47036 (N_47036,N_43556,N_43064);
nor U47037 (N_47037,N_44707,N_43738);
or U47038 (N_47038,N_42585,N_42949);
and U47039 (N_47039,N_43539,N_44814);
xnor U47040 (N_47040,N_42655,N_43343);
nor U47041 (N_47041,N_43776,N_44836);
xor U47042 (N_47042,N_42824,N_43476);
and U47043 (N_47043,N_43814,N_43259);
nor U47044 (N_47044,N_44721,N_43569);
nand U47045 (N_47045,N_44625,N_43544);
and U47046 (N_47046,N_44717,N_43782);
xor U47047 (N_47047,N_42841,N_43423);
nand U47048 (N_47048,N_43823,N_44118);
xor U47049 (N_47049,N_44489,N_44892);
xnor U47050 (N_47050,N_44526,N_43492);
xnor U47051 (N_47051,N_43809,N_44367);
or U47052 (N_47052,N_43558,N_42647);
nor U47053 (N_47053,N_44142,N_43466);
nand U47054 (N_47054,N_43459,N_44561);
nor U47055 (N_47055,N_44075,N_42720);
nand U47056 (N_47056,N_44426,N_44221);
or U47057 (N_47057,N_42830,N_42628);
and U47058 (N_47058,N_43856,N_43214);
nand U47059 (N_47059,N_44153,N_43488);
nor U47060 (N_47060,N_44626,N_44435);
nand U47061 (N_47061,N_43803,N_44954);
nor U47062 (N_47062,N_42758,N_42768);
or U47063 (N_47063,N_42578,N_44744);
xor U47064 (N_47064,N_44297,N_44113);
or U47065 (N_47065,N_43040,N_42687);
and U47066 (N_47066,N_43911,N_43046);
nor U47067 (N_47067,N_44451,N_43196);
and U47068 (N_47068,N_42807,N_43928);
nor U47069 (N_47069,N_44033,N_43218);
nand U47070 (N_47070,N_43951,N_44572);
nor U47071 (N_47071,N_43453,N_42687);
nand U47072 (N_47072,N_44187,N_44278);
and U47073 (N_47073,N_43634,N_43574);
or U47074 (N_47074,N_43802,N_43794);
or U47075 (N_47075,N_43576,N_42887);
xnor U47076 (N_47076,N_43413,N_44743);
and U47077 (N_47077,N_43474,N_44861);
nor U47078 (N_47078,N_44017,N_43232);
and U47079 (N_47079,N_43716,N_42600);
or U47080 (N_47080,N_44381,N_43910);
nor U47081 (N_47081,N_43731,N_44055);
nand U47082 (N_47082,N_44975,N_44579);
or U47083 (N_47083,N_43841,N_44959);
and U47084 (N_47084,N_44685,N_43756);
and U47085 (N_47085,N_44435,N_44674);
xor U47086 (N_47086,N_43895,N_42896);
and U47087 (N_47087,N_44554,N_44448);
and U47088 (N_47088,N_43962,N_42780);
nand U47089 (N_47089,N_42882,N_44746);
xor U47090 (N_47090,N_43630,N_43405);
xor U47091 (N_47091,N_44478,N_44891);
or U47092 (N_47092,N_42956,N_43446);
xor U47093 (N_47093,N_44901,N_44911);
or U47094 (N_47094,N_43752,N_43228);
nand U47095 (N_47095,N_44374,N_44953);
and U47096 (N_47096,N_42547,N_43989);
xnor U47097 (N_47097,N_43178,N_44505);
nor U47098 (N_47098,N_43061,N_42730);
or U47099 (N_47099,N_43382,N_44335);
nor U47100 (N_47100,N_44329,N_43886);
or U47101 (N_47101,N_42512,N_42780);
nand U47102 (N_47102,N_43255,N_42877);
nor U47103 (N_47103,N_43996,N_44452);
or U47104 (N_47104,N_42809,N_43336);
xor U47105 (N_47105,N_43353,N_43073);
nand U47106 (N_47106,N_42523,N_44213);
or U47107 (N_47107,N_43998,N_42604);
nand U47108 (N_47108,N_43622,N_44685);
or U47109 (N_47109,N_44714,N_44829);
xor U47110 (N_47110,N_44073,N_42643);
and U47111 (N_47111,N_43804,N_43806);
xnor U47112 (N_47112,N_42670,N_43005);
or U47113 (N_47113,N_44022,N_43618);
or U47114 (N_47114,N_42578,N_44336);
nand U47115 (N_47115,N_43388,N_42582);
and U47116 (N_47116,N_44205,N_42671);
and U47117 (N_47117,N_43483,N_43070);
or U47118 (N_47118,N_44054,N_43660);
or U47119 (N_47119,N_43187,N_43777);
nand U47120 (N_47120,N_43791,N_43574);
nor U47121 (N_47121,N_44275,N_43982);
or U47122 (N_47122,N_44280,N_43415);
and U47123 (N_47123,N_43000,N_44498);
and U47124 (N_47124,N_44850,N_44475);
and U47125 (N_47125,N_44871,N_43671);
or U47126 (N_47126,N_43758,N_43616);
nor U47127 (N_47127,N_43306,N_43299);
and U47128 (N_47128,N_42626,N_43473);
nor U47129 (N_47129,N_43776,N_42548);
or U47130 (N_47130,N_44782,N_44013);
or U47131 (N_47131,N_44366,N_42708);
or U47132 (N_47132,N_42740,N_44193);
and U47133 (N_47133,N_44603,N_44534);
nand U47134 (N_47134,N_42565,N_43892);
xor U47135 (N_47135,N_43596,N_44718);
or U47136 (N_47136,N_42607,N_43320);
or U47137 (N_47137,N_44420,N_43973);
and U47138 (N_47138,N_44962,N_43663);
and U47139 (N_47139,N_42522,N_44822);
nand U47140 (N_47140,N_44881,N_43783);
xnor U47141 (N_47141,N_43919,N_43884);
nor U47142 (N_47142,N_42508,N_44953);
nor U47143 (N_47143,N_42504,N_43759);
nand U47144 (N_47144,N_43407,N_44970);
nor U47145 (N_47145,N_44650,N_44241);
or U47146 (N_47146,N_42718,N_42730);
nor U47147 (N_47147,N_43421,N_43708);
xor U47148 (N_47148,N_44738,N_43684);
xor U47149 (N_47149,N_44697,N_44546);
and U47150 (N_47150,N_44685,N_43359);
nor U47151 (N_47151,N_43580,N_44821);
nor U47152 (N_47152,N_44293,N_43541);
or U47153 (N_47153,N_44529,N_44133);
and U47154 (N_47154,N_43869,N_43790);
xor U47155 (N_47155,N_44551,N_44368);
and U47156 (N_47156,N_44746,N_44800);
nor U47157 (N_47157,N_43329,N_42563);
and U47158 (N_47158,N_44085,N_44455);
xnor U47159 (N_47159,N_43778,N_43803);
nand U47160 (N_47160,N_43938,N_43187);
xnor U47161 (N_47161,N_43421,N_44078);
and U47162 (N_47162,N_44068,N_42982);
and U47163 (N_47163,N_43574,N_43987);
or U47164 (N_47164,N_43705,N_43747);
and U47165 (N_47165,N_43606,N_43420);
and U47166 (N_47166,N_43432,N_43705);
xnor U47167 (N_47167,N_42838,N_44473);
and U47168 (N_47168,N_43692,N_44309);
and U47169 (N_47169,N_43184,N_43938);
xnor U47170 (N_47170,N_42649,N_43271);
xnor U47171 (N_47171,N_44862,N_43760);
xor U47172 (N_47172,N_42861,N_43570);
xnor U47173 (N_47173,N_43430,N_43911);
xor U47174 (N_47174,N_42884,N_43383);
or U47175 (N_47175,N_44273,N_42824);
nand U47176 (N_47176,N_42934,N_44199);
and U47177 (N_47177,N_44221,N_44157);
nand U47178 (N_47178,N_44668,N_43735);
nor U47179 (N_47179,N_43397,N_44155);
xor U47180 (N_47180,N_42589,N_43382);
and U47181 (N_47181,N_44961,N_43957);
or U47182 (N_47182,N_43443,N_44295);
xnor U47183 (N_47183,N_42807,N_43367);
and U47184 (N_47184,N_44270,N_43374);
and U47185 (N_47185,N_42654,N_43021);
xor U47186 (N_47186,N_42987,N_44405);
nor U47187 (N_47187,N_42790,N_43260);
or U47188 (N_47188,N_42937,N_43988);
nor U47189 (N_47189,N_44885,N_43276);
nor U47190 (N_47190,N_44432,N_42542);
nand U47191 (N_47191,N_43119,N_43395);
xor U47192 (N_47192,N_44198,N_42526);
and U47193 (N_47193,N_44302,N_44239);
and U47194 (N_47194,N_42976,N_43713);
xor U47195 (N_47195,N_43674,N_43645);
xnor U47196 (N_47196,N_44440,N_42557);
or U47197 (N_47197,N_43136,N_43160);
nor U47198 (N_47198,N_43306,N_44212);
or U47199 (N_47199,N_43812,N_44202);
xnor U47200 (N_47200,N_43568,N_44483);
xor U47201 (N_47201,N_43748,N_44611);
nor U47202 (N_47202,N_43910,N_44873);
and U47203 (N_47203,N_43214,N_44095);
nor U47204 (N_47204,N_43101,N_43625);
and U47205 (N_47205,N_43650,N_43579);
and U47206 (N_47206,N_44888,N_44300);
nor U47207 (N_47207,N_42687,N_44565);
or U47208 (N_47208,N_43521,N_44637);
nand U47209 (N_47209,N_44181,N_42576);
xnor U47210 (N_47210,N_42518,N_42763);
and U47211 (N_47211,N_44840,N_44534);
and U47212 (N_47212,N_42601,N_44992);
nand U47213 (N_47213,N_44139,N_44445);
nand U47214 (N_47214,N_43423,N_44223);
and U47215 (N_47215,N_44666,N_44712);
xor U47216 (N_47216,N_42667,N_44116);
xnor U47217 (N_47217,N_42753,N_43051);
and U47218 (N_47218,N_43562,N_43306);
nand U47219 (N_47219,N_43839,N_44992);
or U47220 (N_47220,N_43131,N_44427);
and U47221 (N_47221,N_44964,N_44046);
nand U47222 (N_47222,N_42708,N_44853);
nor U47223 (N_47223,N_42997,N_44590);
nor U47224 (N_47224,N_43341,N_43096);
or U47225 (N_47225,N_44597,N_43822);
or U47226 (N_47226,N_44872,N_44351);
xnor U47227 (N_47227,N_42617,N_44030);
nand U47228 (N_47228,N_43196,N_43804);
nand U47229 (N_47229,N_44487,N_43683);
and U47230 (N_47230,N_43848,N_43705);
or U47231 (N_47231,N_44994,N_43958);
nor U47232 (N_47232,N_44141,N_42812);
or U47233 (N_47233,N_43548,N_43582);
nor U47234 (N_47234,N_43125,N_43243);
nand U47235 (N_47235,N_42868,N_44002);
or U47236 (N_47236,N_43502,N_44760);
xnor U47237 (N_47237,N_42602,N_43631);
or U47238 (N_47238,N_43054,N_43053);
xor U47239 (N_47239,N_44009,N_43774);
or U47240 (N_47240,N_43572,N_43107);
and U47241 (N_47241,N_43528,N_44317);
or U47242 (N_47242,N_44383,N_43045);
and U47243 (N_47243,N_43710,N_44702);
nor U47244 (N_47244,N_42543,N_42960);
xnor U47245 (N_47245,N_44816,N_44323);
or U47246 (N_47246,N_43049,N_43328);
nand U47247 (N_47247,N_42734,N_44698);
and U47248 (N_47248,N_42631,N_44203);
or U47249 (N_47249,N_43938,N_44220);
nand U47250 (N_47250,N_44072,N_44715);
nor U47251 (N_47251,N_43542,N_42718);
nor U47252 (N_47252,N_43289,N_44340);
xnor U47253 (N_47253,N_43705,N_43275);
nand U47254 (N_47254,N_44255,N_42948);
xor U47255 (N_47255,N_44710,N_43895);
or U47256 (N_47256,N_42938,N_42592);
nand U47257 (N_47257,N_44882,N_43419);
nand U47258 (N_47258,N_43459,N_44166);
and U47259 (N_47259,N_43512,N_44090);
xnor U47260 (N_47260,N_42804,N_43241);
xor U47261 (N_47261,N_43117,N_44402);
nor U47262 (N_47262,N_44526,N_42689);
nor U47263 (N_47263,N_44187,N_44582);
or U47264 (N_47264,N_44715,N_42945);
xor U47265 (N_47265,N_42702,N_43162);
or U47266 (N_47266,N_43863,N_43856);
and U47267 (N_47267,N_43228,N_44936);
nor U47268 (N_47268,N_44548,N_43908);
nand U47269 (N_47269,N_44862,N_44515);
nor U47270 (N_47270,N_43387,N_44959);
and U47271 (N_47271,N_44020,N_44740);
or U47272 (N_47272,N_42851,N_44555);
xor U47273 (N_47273,N_44135,N_44275);
or U47274 (N_47274,N_42730,N_44850);
or U47275 (N_47275,N_44144,N_43673);
and U47276 (N_47276,N_42908,N_44753);
xnor U47277 (N_47277,N_44438,N_44432);
or U47278 (N_47278,N_44409,N_44541);
nand U47279 (N_47279,N_43522,N_43179);
nor U47280 (N_47280,N_44016,N_42525);
xnor U47281 (N_47281,N_42973,N_44066);
nand U47282 (N_47282,N_43227,N_43027);
or U47283 (N_47283,N_43483,N_43653);
nand U47284 (N_47284,N_43051,N_44756);
and U47285 (N_47285,N_44352,N_44251);
xor U47286 (N_47286,N_42738,N_42916);
and U47287 (N_47287,N_43342,N_44317);
and U47288 (N_47288,N_43740,N_44726);
nor U47289 (N_47289,N_42732,N_42548);
xnor U47290 (N_47290,N_42936,N_44047);
nand U47291 (N_47291,N_44167,N_42693);
and U47292 (N_47292,N_43155,N_42591);
xnor U47293 (N_47293,N_43891,N_44926);
or U47294 (N_47294,N_44715,N_44992);
xor U47295 (N_47295,N_43797,N_43741);
xnor U47296 (N_47296,N_43762,N_42538);
nand U47297 (N_47297,N_43753,N_44633);
or U47298 (N_47298,N_44924,N_44127);
xor U47299 (N_47299,N_44146,N_44630);
or U47300 (N_47300,N_42763,N_43168);
and U47301 (N_47301,N_43353,N_44392);
nand U47302 (N_47302,N_44269,N_43969);
and U47303 (N_47303,N_43363,N_42648);
nand U47304 (N_47304,N_44094,N_43353);
and U47305 (N_47305,N_44768,N_43701);
nand U47306 (N_47306,N_42839,N_42727);
nand U47307 (N_47307,N_44616,N_43579);
nor U47308 (N_47308,N_44251,N_43661);
xor U47309 (N_47309,N_43085,N_44629);
and U47310 (N_47310,N_43084,N_44966);
or U47311 (N_47311,N_43202,N_43805);
and U47312 (N_47312,N_44492,N_42691);
and U47313 (N_47313,N_43311,N_43039);
and U47314 (N_47314,N_44147,N_43987);
and U47315 (N_47315,N_44489,N_42975);
nand U47316 (N_47316,N_44094,N_42747);
xnor U47317 (N_47317,N_42539,N_42800);
or U47318 (N_47318,N_44363,N_44547);
or U47319 (N_47319,N_42647,N_44936);
nor U47320 (N_47320,N_43790,N_42633);
nor U47321 (N_47321,N_44182,N_42998);
and U47322 (N_47322,N_44788,N_44493);
and U47323 (N_47323,N_43279,N_43094);
nand U47324 (N_47324,N_43447,N_43872);
and U47325 (N_47325,N_44717,N_42643);
nand U47326 (N_47326,N_42922,N_44801);
nand U47327 (N_47327,N_42735,N_43992);
or U47328 (N_47328,N_44765,N_43089);
and U47329 (N_47329,N_42685,N_43286);
and U47330 (N_47330,N_43340,N_44276);
or U47331 (N_47331,N_43565,N_44500);
or U47332 (N_47332,N_44560,N_44659);
xnor U47333 (N_47333,N_44548,N_43071);
and U47334 (N_47334,N_44060,N_42825);
xor U47335 (N_47335,N_43300,N_43322);
nand U47336 (N_47336,N_44742,N_42817);
nor U47337 (N_47337,N_43129,N_43900);
xor U47338 (N_47338,N_43297,N_44575);
nor U47339 (N_47339,N_44734,N_43396);
and U47340 (N_47340,N_43370,N_42545);
and U47341 (N_47341,N_42989,N_44907);
or U47342 (N_47342,N_43131,N_43055);
and U47343 (N_47343,N_42601,N_44153);
and U47344 (N_47344,N_44583,N_42633);
or U47345 (N_47345,N_43698,N_42742);
xor U47346 (N_47346,N_44922,N_43613);
nand U47347 (N_47347,N_43232,N_43283);
or U47348 (N_47348,N_44026,N_43003);
or U47349 (N_47349,N_43395,N_44772);
nor U47350 (N_47350,N_43629,N_43541);
and U47351 (N_47351,N_44016,N_42943);
nor U47352 (N_47352,N_44543,N_43879);
xnor U47353 (N_47353,N_42650,N_43305);
and U47354 (N_47354,N_44703,N_43018);
xor U47355 (N_47355,N_43868,N_44302);
nor U47356 (N_47356,N_43964,N_43383);
and U47357 (N_47357,N_42819,N_44677);
nand U47358 (N_47358,N_42723,N_44645);
nand U47359 (N_47359,N_44531,N_43030);
or U47360 (N_47360,N_43358,N_43198);
xnor U47361 (N_47361,N_44221,N_43733);
nor U47362 (N_47362,N_44752,N_43755);
nand U47363 (N_47363,N_42633,N_44625);
or U47364 (N_47364,N_43709,N_44158);
or U47365 (N_47365,N_44471,N_44490);
and U47366 (N_47366,N_44944,N_44298);
or U47367 (N_47367,N_43396,N_44795);
xnor U47368 (N_47368,N_42982,N_44811);
or U47369 (N_47369,N_43990,N_43005);
nand U47370 (N_47370,N_43143,N_42697);
nor U47371 (N_47371,N_43572,N_44873);
xnor U47372 (N_47372,N_43465,N_42593);
or U47373 (N_47373,N_43235,N_43103);
and U47374 (N_47374,N_43367,N_43019);
nand U47375 (N_47375,N_44239,N_44346);
nor U47376 (N_47376,N_43977,N_43212);
nor U47377 (N_47377,N_44838,N_42806);
or U47378 (N_47378,N_43747,N_44379);
nand U47379 (N_47379,N_43143,N_43129);
xnor U47380 (N_47380,N_43074,N_44180);
nor U47381 (N_47381,N_44920,N_43840);
and U47382 (N_47382,N_43065,N_42590);
xnor U47383 (N_47383,N_42560,N_44243);
nand U47384 (N_47384,N_42753,N_43776);
and U47385 (N_47385,N_44431,N_44198);
xor U47386 (N_47386,N_43762,N_44482);
and U47387 (N_47387,N_44626,N_44306);
nand U47388 (N_47388,N_43657,N_44120);
or U47389 (N_47389,N_43216,N_43556);
or U47390 (N_47390,N_42800,N_44309);
nand U47391 (N_47391,N_44107,N_42757);
nand U47392 (N_47392,N_43987,N_42831);
nor U47393 (N_47393,N_44979,N_44946);
or U47394 (N_47394,N_43239,N_43308);
or U47395 (N_47395,N_44810,N_43422);
or U47396 (N_47396,N_43071,N_42666);
nand U47397 (N_47397,N_44434,N_43724);
nand U47398 (N_47398,N_44992,N_42779);
xnor U47399 (N_47399,N_44119,N_42544);
nor U47400 (N_47400,N_43212,N_44077);
nand U47401 (N_47401,N_44446,N_43293);
nand U47402 (N_47402,N_43530,N_42909);
and U47403 (N_47403,N_44840,N_43689);
or U47404 (N_47404,N_42810,N_43572);
and U47405 (N_47405,N_43834,N_44364);
and U47406 (N_47406,N_43925,N_44291);
nor U47407 (N_47407,N_43304,N_43877);
and U47408 (N_47408,N_44827,N_43931);
and U47409 (N_47409,N_43108,N_43348);
nor U47410 (N_47410,N_43672,N_43977);
and U47411 (N_47411,N_44185,N_43875);
nand U47412 (N_47412,N_42913,N_43152);
nor U47413 (N_47413,N_43828,N_42587);
nand U47414 (N_47414,N_43903,N_44475);
nand U47415 (N_47415,N_44443,N_42619);
or U47416 (N_47416,N_43018,N_44673);
xor U47417 (N_47417,N_44986,N_44499);
xnor U47418 (N_47418,N_42999,N_44677);
nand U47419 (N_47419,N_42658,N_44227);
xnor U47420 (N_47420,N_44517,N_43574);
and U47421 (N_47421,N_43322,N_44275);
nor U47422 (N_47422,N_44604,N_43437);
or U47423 (N_47423,N_43624,N_44584);
or U47424 (N_47424,N_43583,N_44836);
nor U47425 (N_47425,N_44180,N_43094);
and U47426 (N_47426,N_43610,N_43915);
or U47427 (N_47427,N_44072,N_43801);
or U47428 (N_47428,N_42569,N_44674);
or U47429 (N_47429,N_44032,N_43879);
or U47430 (N_47430,N_44625,N_44136);
nor U47431 (N_47431,N_44375,N_43641);
nor U47432 (N_47432,N_43432,N_42814);
nand U47433 (N_47433,N_43160,N_44687);
nor U47434 (N_47434,N_43566,N_44123);
and U47435 (N_47435,N_42940,N_42903);
or U47436 (N_47436,N_44721,N_43917);
nor U47437 (N_47437,N_42968,N_43575);
or U47438 (N_47438,N_43970,N_43139);
nor U47439 (N_47439,N_43071,N_44977);
nand U47440 (N_47440,N_44406,N_43588);
nand U47441 (N_47441,N_44938,N_43604);
nand U47442 (N_47442,N_43474,N_44031);
nand U47443 (N_47443,N_44416,N_44736);
or U47444 (N_47444,N_43972,N_43271);
nand U47445 (N_47445,N_44859,N_42771);
nand U47446 (N_47446,N_42719,N_43114);
or U47447 (N_47447,N_44366,N_42702);
or U47448 (N_47448,N_43558,N_43623);
nor U47449 (N_47449,N_42826,N_44277);
nand U47450 (N_47450,N_44378,N_42509);
and U47451 (N_47451,N_44356,N_44987);
nand U47452 (N_47452,N_44014,N_44822);
nor U47453 (N_47453,N_43673,N_43772);
xor U47454 (N_47454,N_44566,N_43103);
nand U47455 (N_47455,N_43762,N_44669);
nand U47456 (N_47456,N_44692,N_43890);
and U47457 (N_47457,N_43264,N_43656);
xor U47458 (N_47458,N_43363,N_43020);
nand U47459 (N_47459,N_44790,N_44360);
or U47460 (N_47460,N_43857,N_44670);
nor U47461 (N_47461,N_44634,N_44664);
nor U47462 (N_47462,N_44329,N_42930);
and U47463 (N_47463,N_43405,N_43913);
and U47464 (N_47464,N_44597,N_43505);
nor U47465 (N_47465,N_44365,N_43957);
or U47466 (N_47466,N_44272,N_44980);
and U47467 (N_47467,N_44990,N_43822);
xnor U47468 (N_47468,N_44590,N_44897);
xor U47469 (N_47469,N_44413,N_42724);
or U47470 (N_47470,N_44227,N_43681);
nor U47471 (N_47471,N_44584,N_44044);
nor U47472 (N_47472,N_43101,N_42517);
or U47473 (N_47473,N_43553,N_43992);
nor U47474 (N_47474,N_44215,N_44223);
nand U47475 (N_47475,N_43845,N_42725);
or U47476 (N_47476,N_44594,N_44362);
xor U47477 (N_47477,N_43058,N_42761);
or U47478 (N_47478,N_44438,N_44731);
and U47479 (N_47479,N_43368,N_43745);
or U47480 (N_47480,N_42711,N_43040);
nor U47481 (N_47481,N_42695,N_44974);
nor U47482 (N_47482,N_44259,N_44027);
nor U47483 (N_47483,N_44820,N_44628);
and U47484 (N_47484,N_44777,N_43761);
nand U47485 (N_47485,N_44112,N_44094);
xor U47486 (N_47486,N_43704,N_44500);
or U47487 (N_47487,N_44627,N_43445);
and U47488 (N_47488,N_44953,N_44234);
and U47489 (N_47489,N_44219,N_43179);
nor U47490 (N_47490,N_43031,N_43682);
nand U47491 (N_47491,N_42860,N_44210);
and U47492 (N_47492,N_42620,N_42733);
or U47493 (N_47493,N_44522,N_43211);
xor U47494 (N_47494,N_43904,N_44369);
and U47495 (N_47495,N_42816,N_43957);
xor U47496 (N_47496,N_44530,N_42773);
nand U47497 (N_47497,N_44115,N_44119);
and U47498 (N_47498,N_42959,N_43728);
xnor U47499 (N_47499,N_44794,N_44709);
xnor U47500 (N_47500,N_45054,N_45510);
nor U47501 (N_47501,N_47197,N_45204);
and U47502 (N_47502,N_46743,N_46499);
xor U47503 (N_47503,N_46457,N_45970);
xor U47504 (N_47504,N_45177,N_45543);
xor U47505 (N_47505,N_46265,N_46857);
xor U47506 (N_47506,N_45211,N_45646);
nand U47507 (N_47507,N_47348,N_47010);
and U47508 (N_47508,N_47017,N_46945);
nand U47509 (N_47509,N_46599,N_46205);
nor U47510 (N_47510,N_46395,N_46113);
or U47511 (N_47511,N_47246,N_45459);
and U47512 (N_47512,N_46199,N_47373);
nand U47513 (N_47513,N_45294,N_46699);
nor U47514 (N_47514,N_47486,N_46950);
nor U47515 (N_47515,N_45585,N_45805);
and U47516 (N_47516,N_47125,N_47257);
nor U47517 (N_47517,N_46559,N_46569);
and U47518 (N_47518,N_47371,N_45963);
and U47519 (N_47519,N_45097,N_45765);
nor U47520 (N_47520,N_46180,N_46316);
nor U47521 (N_47521,N_45352,N_46157);
or U47522 (N_47522,N_47492,N_45514);
nor U47523 (N_47523,N_46823,N_45045);
or U47524 (N_47524,N_46261,N_45881);
and U47525 (N_47525,N_46749,N_47222);
and U47526 (N_47526,N_45600,N_45768);
or U47527 (N_47527,N_46879,N_45184);
or U47528 (N_47528,N_45152,N_46610);
nor U47529 (N_47529,N_45428,N_47377);
nand U47530 (N_47530,N_47354,N_47387);
and U47531 (N_47531,N_47198,N_47108);
nand U47532 (N_47532,N_45863,N_45739);
xor U47533 (N_47533,N_46688,N_46022);
nor U47534 (N_47534,N_45453,N_45784);
xor U47535 (N_47535,N_45532,N_47288);
nand U47536 (N_47536,N_45393,N_46542);
and U47537 (N_47537,N_45205,N_45363);
and U47538 (N_47538,N_46168,N_46509);
or U47539 (N_47539,N_45327,N_47165);
and U47540 (N_47540,N_47478,N_45912);
nand U47541 (N_47541,N_46755,N_47013);
nor U47542 (N_47542,N_45182,N_46474);
or U47543 (N_47543,N_47410,N_45122);
or U47544 (N_47544,N_46731,N_47335);
or U47545 (N_47545,N_45006,N_46463);
nand U47546 (N_47546,N_47475,N_46141);
nor U47547 (N_47547,N_45893,N_46767);
or U47548 (N_47548,N_45155,N_45228);
xor U47549 (N_47549,N_45396,N_45917);
or U47550 (N_47550,N_47375,N_47468);
nor U47551 (N_47551,N_45435,N_47226);
and U47552 (N_47552,N_46119,N_46937);
xnor U47553 (N_47553,N_47160,N_45340);
xnor U47554 (N_47554,N_46271,N_46270);
nor U47555 (N_47555,N_45521,N_45918);
xnor U47556 (N_47556,N_46618,N_45538);
or U47557 (N_47557,N_46919,N_47298);
and U47558 (N_47558,N_46829,N_46279);
xnor U47559 (N_47559,N_45458,N_45021);
nand U47560 (N_47560,N_45198,N_47183);
and U47561 (N_47561,N_45418,N_47404);
xnor U47562 (N_47562,N_46131,N_45989);
and U47563 (N_47563,N_46605,N_45564);
nor U47564 (N_47564,N_45406,N_46775);
and U47565 (N_47565,N_45984,N_46764);
or U47566 (N_47566,N_45381,N_45433);
nor U47567 (N_47567,N_46303,N_46813);
nor U47568 (N_47568,N_47359,N_46304);
xnor U47569 (N_47569,N_45391,N_46811);
and U47570 (N_47570,N_45120,N_45879);
nand U47571 (N_47571,N_45309,N_46295);
xor U47572 (N_47572,N_47086,N_47497);
nor U47573 (N_47573,N_45560,N_46149);
or U47574 (N_47574,N_47031,N_45566);
nand U47575 (N_47575,N_45050,N_45799);
xor U47576 (N_47576,N_46790,N_46447);
nor U47577 (N_47577,N_46747,N_46153);
or U47578 (N_47578,N_45596,N_46932);
nor U47579 (N_47579,N_46333,N_47083);
nor U47580 (N_47580,N_46514,N_46694);
and U47581 (N_47581,N_45154,N_45470);
nand U47582 (N_47582,N_45807,N_45827);
nand U47583 (N_47583,N_47364,N_45100);
nand U47584 (N_47584,N_45474,N_46120);
nor U47585 (N_47585,N_45246,N_45826);
nand U47586 (N_47586,N_47403,N_45713);
or U47587 (N_47587,N_45878,N_45606);
and U47588 (N_47588,N_46837,N_45562);
nand U47589 (N_47589,N_46982,N_46573);
and U47590 (N_47590,N_46492,N_45056);
or U47591 (N_47591,N_45550,N_46906);
and U47592 (N_47592,N_46976,N_46148);
nor U47593 (N_47593,N_46072,N_47337);
and U47594 (N_47594,N_45892,N_45462);
nand U47595 (N_47595,N_47191,N_47161);
and U47596 (N_47596,N_45592,N_46292);
and U47597 (N_47597,N_45476,N_45871);
xnor U47598 (N_47598,N_46810,N_47418);
and U47599 (N_47599,N_45192,N_45452);
nor U47600 (N_47600,N_46478,N_45854);
nand U47601 (N_47601,N_45516,N_46834);
nor U47602 (N_47602,N_47232,N_47319);
nand U47603 (N_47603,N_45783,N_45282);
nor U47604 (N_47604,N_46563,N_46912);
nand U47605 (N_47605,N_46000,N_46415);
or U47606 (N_47606,N_47392,N_45068);
xnor U47607 (N_47607,N_45414,N_46870);
nor U47608 (N_47608,N_45319,N_45426);
or U47609 (N_47609,N_46795,N_47442);
nor U47610 (N_47610,N_46904,N_45561);
and U47611 (N_47611,N_45176,N_45110);
nand U47612 (N_47612,N_47391,N_46323);
or U47613 (N_47613,N_47467,N_46515);
nor U47614 (N_47614,N_46601,N_45896);
nand U47615 (N_47615,N_45390,N_46355);
and U47616 (N_47616,N_46343,N_47098);
and U47617 (N_47617,N_47065,N_47106);
or U47618 (N_47618,N_45326,N_46472);
nor U47619 (N_47619,N_45049,N_46505);
nor U47620 (N_47620,N_47015,N_45785);
xnor U47621 (N_47621,N_45343,N_45051);
or U47622 (N_47622,N_45798,N_45541);
xnor U47623 (N_47623,N_45643,N_45368);
and U47624 (N_47624,N_46252,N_45345);
or U47625 (N_47625,N_46554,N_45446);
nor U47626 (N_47626,N_47368,N_46535);
nor U47627 (N_47627,N_45577,N_45866);
nand U47628 (N_47628,N_47394,N_47118);
xor U47629 (N_47629,N_46329,N_47050);
nand U47630 (N_47630,N_46911,N_46382);
nand U47631 (N_47631,N_47320,N_45681);
and U47632 (N_47632,N_47097,N_46284);
nand U47633 (N_47633,N_47437,N_46628);
nor U47634 (N_47634,N_45786,N_45818);
nor U47635 (N_47635,N_45266,N_46787);
xnor U47636 (N_47636,N_45316,N_46695);
or U47637 (N_47637,N_45598,N_47251);
nor U47638 (N_47638,N_47349,N_46549);
or U47639 (N_47639,N_45667,N_45138);
nor U47640 (N_47640,N_46645,N_45355);
xor U47641 (N_47641,N_46909,N_46154);
and U47642 (N_47642,N_45972,N_47292);
nand U47643 (N_47643,N_45948,N_46449);
and U47644 (N_47644,N_46405,N_46521);
xor U47645 (N_47645,N_45517,N_45243);
nand U47646 (N_47646,N_45447,N_45329);
or U47647 (N_47647,N_46267,N_46724);
and U47648 (N_47648,N_46972,N_45528);
xnor U47649 (N_47649,N_45167,N_47301);
nand U47650 (N_47650,N_46916,N_45145);
xor U47651 (N_47651,N_46793,N_46207);
nor U47652 (N_47652,N_45075,N_45481);
nand U47653 (N_47653,N_45280,N_46309);
nor U47654 (N_47654,N_46626,N_45523);
and U47655 (N_47655,N_47293,N_45947);
nand U47656 (N_47656,N_46864,N_46989);
nor U47657 (N_47657,N_45501,N_45583);
or U47658 (N_47658,N_45581,N_46105);
nand U47659 (N_47659,N_46954,N_46381);
and U47660 (N_47660,N_45720,N_46018);
nand U47661 (N_47661,N_47149,N_46680);
xnor U47662 (N_47662,N_46788,N_47011);
and U47663 (N_47663,N_47234,N_46312);
and U47664 (N_47664,N_46780,N_46967);
and U47665 (N_47665,N_45109,N_46566);
or U47666 (N_47666,N_46745,N_45370);
nor U47667 (N_47667,N_45618,N_45819);
xnor U47668 (N_47668,N_47248,N_47169);
xor U47669 (N_47669,N_47090,N_46838);
nand U47670 (N_47670,N_45662,N_46806);
nand U47671 (N_47671,N_47489,N_45968);
nor U47672 (N_47672,N_47019,N_45868);
or U47673 (N_47673,N_46371,N_47122);
nand U47674 (N_47674,N_45227,N_46112);
and U47675 (N_47675,N_45835,N_47300);
nand U47676 (N_47676,N_46190,N_45465);
or U47677 (N_47677,N_47473,N_46920);
nor U47678 (N_47678,N_46944,N_46773);
or U47679 (N_47679,N_46173,N_45808);
or U47680 (N_47680,N_46663,N_45718);
xor U47681 (N_47681,N_47179,N_46956);
xnor U47682 (N_47682,N_47444,N_46783);
or U47683 (N_47683,N_46987,N_46869);
and U47684 (N_47684,N_45650,N_46210);
or U47685 (N_47685,N_45519,N_46721);
and U47686 (N_47686,N_47295,N_46875);
or U47687 (N_47687,N_45487,N_46975);
or U47688 (N_47688,N_45450,N_47395);
nor U47689 (N_47689,N_46452,N_45952);
nor U47690 (N_47690,N_45616,N_45131);
and U47691 (N_47691,N_45873,N_45960);
xnor U47692 (N_47692,N_46936,N_46513);
nor U47693 (N_47693,N_45945,N_45530);
xor U47694 (N_47694,N_45694,N_45953);
xor U47695 (N_47695,N_45730,N_47376);
xnor U47696 (N_47696,N_45235,N_46299);
or U47697 (N_47697,N_46416,N_47303);
xnor U47698 (N_47698,N_47408,N_46727);
nand U47699 (N_47699,N_46871,N_46971);
nand U47700 (N_47700,N_46071,N_46289);
xor U47701 (N_47701,N_47210,N_47341);
and U47702 (N_47702,N_47070,N_45312);
xor U47703 (N_47703,N_45283,N_47220);
nor U47704 (N_47704,N_46523,N_45306);
xnor U47705 (N_47705,N_45734,N_46816);
nand U47706 (N_47706,N_45195,N_45727);
and U47707 (N_47707,N_45492,N_45877);
and U47708 (N_47708,N_45978,N_46953);
xor U47709 (N_47709,N_47150,N_46849);
nand U47710 (N_47710,N_46052,N_45471);
xnor U47711 (N_47711,N_46178,N_45810);
or U47712 (N_47712,N_46502,N_45437);
nand U47713 (N_47713,N_46019,N_46596);
nand U47714 (N_47714,N_46127,N_45388);
and U47715 (N_47715,N_47052,N_46692);
xor U47716 (N_47716,N_45086,N_47170);
xor U47717 (N_47717,N_46651,N_46058);
nand U47718 (N_47718,N_46774,N_45518);
nand U47719 (N_47719,N_45876,N_46209);
or U47720 (N_47720,N_46101,N_46527);
nand U47721 (N_47721,N_45889,N_46337);
nor U47722 (N_47722,N_45956,N_47036);
and U47723 (N_47723,N_45701,N_45148);
or U47724 (N_47724,N_45536,N_46438);
nor U47725 (N_47725,N_46188,N_46958);
xnor U47726 (N_47726,N_46044,N_47254);
or U47727 (N_47727,N_46929,N_46193);
xnor U47728 (N_47728,N_47075,N_45602);
or U47729 (N_47729,N_47272,N_45922);
nor U47730 (N_47730,N_47326,N_45104);
xor U47731 (N_47731,N_45130,N_46082);
or U47732 (N_47732,N_45369,N_46934);
nor U47733 (N_47733,N_47464,N_45020);
and U47734 (N_47734,N_46574,N_46589);
xnor U47735 (N_47735,N_45321,N_45842);
nor U47736 (N_47736,N_45942,N_45376);
or U47737 (N_47737,N_45715,N_46933);
nor U47738 (N_47738,N_46025,N_46256);
or U47739 (N_47739,N_46232,N_45062);
nand U47740 (N_47740,N_46595,N_46012);
xnor U47741 (N_47741,N_46181,N_47476);
or U47742 (N_47742,N_47455,N_45677);
nand U47743 (N_47743,N_45674,N_46225);
nor U47744 (N_47744,N_45128,N_46135);
or U47745 (N_47745,N_45609,N_45199);
and U47746 (N_47746,N_45242,N_45034);
xor U47747 (N_47747,N_46317,N_47422);
or U47748 (N_47748,N_47152,N_46147);
nor U47749 (N_47749,N_45706,N_46443);
nor U47750 (N_47750,N_46822,N_47067);
xor U47751 (N_47751,N_45931,N_47005);
nand U47752 (N_47752,N_45895,N_45307);
and U47753 (N_47753,N_46796,N_46288);
and U47754 (N_47754,N_46216,N_45024);
nor U47755 (N_47755,N_46177,N_46801);
nand U47756 (N_47756,N_46506,N_46576);
nand U47757 (N_47757,N_45157,N_46003);
or U47758 (N_47758,N_45082,N_45351);
nor U47759 (N_47759,N_46241,N_45454);
and U47760 (N_47760,N_46394,N_45838);
and U47761 (N_47761,N_46679,N_47109);
nand U47762 (N_47762,N_45615,N_46620);
nor U47763 (N_47763,N_47176,N_46732);
and U47764 (N_47764,N_47379,N_46196);
xor U47765 (N_47765,N_45737,N_47001);
or U47766 (N_47766,N_45332,N_45624);
nor U47767 (N_47767,N_46378,N_47463);
and U47768 (N_47768,N_45257,N_46377);
xor U47769 (N_47769,N_46862,N_47207);
nand U47770 (N_47770,N_45553,N_45248);
nor U47771 (N_47771,N_47402,N_46674);
or U47772 (N_47772,N_46826,N_45143);
or U47773 (N_47773,N_45744,N_45822);
and U47774 (N_47774,N_45439,N_46686);
and U47775 (N_47775,N_46089,N_46957);
nor U47776 (N_47776,N_46202,N_45241);
or U47777 (N_47777,N_45796,N_47482);
nand U47778 (N_47778,N_46244,N_47143);
nor U47779 (N_47779,N_46062,N_46517);
xor U47780 (N_47780,N_45318,N_46898);
or U47781 (N_47781,N_47003,N_46669);
nor U47782 (N_47782,N_47397,N_47038);
or U47783 (N_47783,N_47494,N_46363);
or U47784 (N_47784,N_45974,N_46078);
or U47785 (N_47785,N_46307,N_46100);
and U47786 (N_47786,N_45411,N_45404);
or U47787 (N_47787,N_46151,N_45627);
nand U47788 (N_47788,N_45855,N_45412);
nor U47789 (N_47789,N_47315,N_45179);
or U47790 (N_47790,N_45508,N_45716);
xor U47791 (N_47791,N_46219,N_46994);
or U47792 (N_47792,N_45007,N_45840);
xnor U47793 (N_47793,N_45567,N_47488);
xnor U47794 (N_47794,N_46621,N_46516);
nor U47795 (N_47795,N_46214,N_46922);
nor U47796 (N_47796,N_45679,N_45031);
nand U47797 (N_47797,N_46725,N_45621);
nor U47798 (N_47798,N_46541,N_45569);
xor U47799 (N_47799,N_45683,N_47092);
or U47800 (N_47800,N_46325,N_46518);
and U47801 (N_47801,N_47120,N_45019);
and U47802 (N_47802,N_47068,N_45353);
nor U47803 (N_47803,N_45524,N_45310);
and U47804 (N_47804,N_45346,N_46080);
xor U47805 (N_47805,N_45788,N_46035);
or U47806 (N_47806,N_47278,N_46006);
xnor U47807 (N_47807,N_47474,N_45688);
xor U47808 (N_47808,N_46186,N_47131);
or U47809 (N_47809,N_46239,N_45548);
and U47810 (N_47810,N_45026,N_46741);
xor U47811 (N_47811,N_45431,N_46771);
xnor U47812 (N_47812,N_45486,N_46411);
nand U47813 (N_47813,N_46708,N_46665);
and U47814 (N_47814,N_45502,N_47247);
nand U47815 (N_47815,N_45664,N_45975);
nor U47816 (N_47816,N_46029,N_46040);
and U47817 (N_47817,N_45407,N_47496);
and U47818 (N_47818,N_46092,N_46495);
and U47819 (N_47819,N_46166,N_47325);
nand U47820 (N_47820,N_46020,N_46122);
nand U47821 (N_47821,N_45913,N_46426);
nand U47822 (N_47822,N_46555,N_47267);
nor U47823 (N_47823,N_47260,N_46736);
xnor U47824 (N_47824,N_45311,N_47366);
xnor U47825 (N_47825,N_46497,N_45747);
and U47826 (N_47826,N_46852,N_46968);
or U47827 (N_47827,N_47470,N_46306);
nor U47828 (N_47828,N_46921,N_46602);
xor U47829 (N_47829,N_46700,N_47020);
or U47830 (N_47830,N_46756,N_46066);
nand U47831 (N_47831,N_46877,N_46844);
xnor U47832 (N_47832,N_46619,N_47499);
or U47833 (N_47833,N_46588,N_45595);
nand U47834 (N_47834,N_45721,N_47243);
nand U47835 (N_47835,N_46045,N_47256);
and U47836 (N_47836,N_46750,N_45885);
and U47837 (N_47837,N_45513,N_46013);
and U47838 (N_47838,N_47205,N_46797);
nor U47839 (N_47839,N_47330,N_47206);
nor U47840 (N_47840,N_47144,N_45187);
nor U47841 (N_47841,N_46630,N_45758);
xor U47842 (N_47842,N_46524,N_47009);
and U47843 (N_47843,N_45977,N_46161);
nor U47844 (N_47844,N_46866,N_45183);
nand U47845 (N_47845,N_46245,N_45253);
and U47846 (N_47846,N_46201,N_46489);
and U47847 (N_47847,N_45073,N_45633);
or U47848 (N_47848,N_47268,N_46341);
or U47849 (N_47849,N_45905,N_47438);
xor U47850 (N_47850,N_46636,N_45812);
and U47851 (N_47851,N_46735,N_45696);
xor U47852 (N_47852,N_45920,N_47324);
xnor U47853 (N_47853,N_45834,N_45180);
or U47854 (N_47854,N_46730,N_45262);
nor U47855 (N_47855,N_45373,N_45946);
and U47856 (N_47856,N_46768,N_46717);
nand U47857 (N_47857,N_45995,N_46712);
and U47858 (N_47858,N_46140,N_45599);
nor U47859 (N_47859,N_46675,N_46462);
nand U47860 (N_47860,N_46393,N_45274);
nor U47861 (N_47861,N_46691,N_45766);
xor U47862 (N_47862,N_47262,N_46427);
nand U47863 (N_47863,N_46404,N_45601);
xnor U47864 (N_47864,N_45137,N_45728);
xor U47865 (N_47865,N_45668,N_47269);
nand U47866 (N_47866,N_46136,N_45815);
and U47867 (N_47867,N_45959,N_47209);
xnor U47868 (N_47868,N_47155,N_45237);
nand U47869 (N_47869,N_45746,N_45413);
and U47870 (N_47870,N_46658,N_45982);
nand U47871 (N_47871,N_47338,N_46991);
and U47872 (N_47872,N_45557,N_45654);
nor U47873 (N_47873,N_45638,N_46234);
and U47874 (N_47874,N_47175,N_45273);
or U47875 (N_47875,N_45490,N_45379);
xor U47876 (N_47876,N_45079,N_46034);
and U47877 (N_47877,N_47177,N_47213);
nand U47878 (N_47878,N_47360,N_47157);
xor U47879 (N_47879,N_46272,N_46752);
nor U47880 (N_47880,N_46762,N_47225);
nor U47881 (N_47881,N_46264,N_45537);
xor U47882 (N_47882,N_46562,N_47327);
xnor U47883 (N_47883,N_46908,N_47104);
nor U47884 (N_47884,N_45193,N_46028);
xor U47885 (N_47885,N_46361,N_46017);
xor U47886 (N_47886,N_45580,N_46758);
or U47887 (N_47887,N_46580,N_46734);
nand U47888 (N_47888,N_47171,N_47045);
and U47889 (N_47889,N_45121,N_46726);
nor U47890 (N_47890,N_46941,N_47481);
nor U47891 (N_47891,N_47336,N_45238);
or U47892 (N_47892,N_47424,N_45202);
nand U47893 (N_47893,N_45289,N_45099);
nand U47894 (N_47894,N_46792,N_46423);
and U47895 (N_47895,N_45658,N_45707);
or U47896 (N_47896,N_46269,N_45083);
or U47897 (N_47897,N_47182,N_46597);
xor U47898 (N_47898,N_47353,N_47201);
and U47899 (N_47899,N_45231,N_45297);
or U47900 (N_47900,N_47283,N_45617);
nor U47901 (N_47901,N_45801,N_45443);
and U47902 (N_47902,N_47087,N_46410);
or U47903 (N_47903,N_47066,N_45880);
nand U47904 (N_47904,N_46999,N_45219);
or U47905 (N_47905,N_47261,N_46318);
nor U47906 (N_47906,N_46375,N_45702);
nor U47907 (N_47907,N_45623,N_45132);
nand U47908 (N_47908,N_45690,N_45259);
and U47909 (N_47909,N_45055,N_46339);
xnor U47910 (N_47910,N_45856,N_45276);
and U47911 (N_47911,N_46760,N_46093);
xor U47912 (N_47912,N_45457,N_45657);
nand U47913 (N_47913,N_45691,N_45698);
nor U47914 (N_47914,N_47224,N_46414);
nand U47915 (N_47915,N_47378,N_45763);
and U47916 (N_47916,N_46099,N_47334);
nor U47917 (N_47917,N_47483,N_45709);
nand U47918 (N_47918,N_46627,N_45572);
and U47919 (N_47919,N_46412,N_45999);
xor U47920 (N_47920,N_47119,N_45094);
xor U47921 (N_47921,N_47469,N_46440);
or U47922 (N_47922,N_45882,N_45542);
and U47923 (N_47923,N_47216,N_45405);
and U47924 (N_47924,N_46467,N_47372);
nor U47925 (N_47925,N_45330,N_45001);
or U47926 (N_47926,N_45908,N_45022);
and U47927 (N_47927,N_46334,N_46431);
nand U47928 (N_47928,N_46631,N_45813);
xnor U47929 (N_47929,N_46676,N_47048);
nand U47930 (N_47930,N_45047,N_45467);
nand U47931 (N_47931,N_47047,N_45787);
or U47932 (N_47932,N_46835,N_45849);
nor U47933 (N_47933,N_45214,N_45649);
xor U47934 (N_47934,N_45539,N_46081);
or U47935 (N_47935,N_45797,N_46682);
nand U47936 (N_47936,N_45399,N_45781);
or U47937 (N_47937,N_47282,N_46847);
and U47938 (N_47938,N_45013,N_47164);
nand U47939 (N_47939,N_45589,N_46860);
nand U47940 (N_47940,N_47082,N_46004);
and U47941 (N_47941,N_47495,N_46884);
xnor U47942 (N_47942,N_45949,N_45301);
xnor U47943 (N_47943,N_45299,N_47227);
nor U47944 (N_47944,N_46108,N_46946);
and U47945 (N_47945,N_46073,N_46508);
nand U47946 (N_47946,N_45194,N_45772);
and U47947 (N_47947,N_45582,N_45852);
xnor U47948 (N_47948,N_45093,N_46159);
or U47949 (N_47949,N_47071,N_45263);
or U47950 (N_47950,N_46503,N_47331);
nor U47951 (N_47951,N_46453,N_47145);
nand U47952 (N_47952,N_45255,N_46237);
or U47953 (N_47953,N_46470,N_47297);
and U47954 (N_47954,N_46890,N_47200);
nor U47955 (N_47955,N_45899,N_45637);
or U47956 (N_47956,N_46498,N_46907);
nand U47957 (N_47957,N_46403,N_45377);
xnor U47958 (N_47958,N_46077,N_46704);
and U47959 (N_47959,N_46054,N_45916);
nand U47960 (N_47960,N_46947,N_46327);
or U47961 (N_47961,N_45239,N_45841);
nor U47962 (N_47962,N_47398,N_45985);
or U47963 (N_47963,N_46742,N_45547);
nand U47964 (N_47964,N_45244,N_46273);
and U47965 (N_47965,N_47317,N_47113);
nor U47966 (N_47966,N_46711,N_45040);
or U47967 (N_47967,N_45017,N_46294);
nand U47968 (N_47968,N_45622,N_45046);
nor U47969 (N_47969,N_45287,N_45894);
nor U47970 (N_47970,N_45267,N_46642);
nand U47971 (N_47971,N_46370,N_45284);
or U47972 (N_47972,N_47252,N_45305);
nor U47973 (N_47973,N_46814,N_46685);
and U47974 (N_47974,N_45697,N_45349);
nor U47975 (N_47975,N_45794,N_46778);
or U47976 (N_47976,N_46887,N_46384);
nor U47977 (N_47977,N_45843,N_46718);
and U47978 (N_47978,N_46301,N_46995);
xor U47979 (N_47979,N_46939,N_46298);
and U47980 (N_47980,N_46226,N_45139);
nor U47981 (N_47981,N_45515,N_46182);
or U47982 (N_47982,N_45037,N_47188);
nand U47983 (N_47983,N_47195,N_45570);
and U47984 (N_47984,N_46359,N_45846);
and U47985 (N_47985,N_45230,N_45910);
xor U47986 (N_47986,N_45188,N_47416);
xor U47987 (N_47987,N_46859,N_46152);
xnor U47988 (N_47988,N_47352,N_46023);
nand U47989 (N_47989,N_46090,N_45969);
xnor U47990 (N_47990,N_47244,N_46753);
nor U47991 (N_47991,N_45671,N_45669);
xor U47992 (N_47992,N_45344,N_45904);
and U47993 (N_47993,N_46038,N_46354);
or U47994 (N_47994,N_46534,N_46970);
or U47995 (N_47995,N_45229,N_45200);
nor U47996 (N_47996,N_45990,N_46442);
nor U47997 (N_47997,N_45087,N_45764);
xnor U47998 (N_47998,N_46710,N_46399);
or U47999 (N_47999,N_46435,N_46615);
nand U48000 (N_48000,N_46046,N_47415);
and U48001 (N_48001,N_45575,N_46132);
nand U48002 (N_48002,N_46635,N_45171);
and U48003 (N_48003,N_46668,N_47032);
nand U48004 (N_48004,N_46121,N_47037);
and U48005 (N_48005,N_45261,N_47409);
xnor U48006 (N_48006,N_46656,N_46379);
nor U48007 (N_48007,N_45686,N_45400);
and U48008 (N_48008,N_46009,N_47008);
and U48009 (N_48009,N_45484,N_46229);
or U48010 (N_48010,N_45756,N_47187);
nand U48011 (N_48011,N_45504,N_46662);
nor U48012 (N_48012,N_47228,N_45277);
and U48013 (N_48013,N_47007,N_46344);
xor U48014 (N_48014,N_46433,N_45264);
and U48015 (N_48015,N_46043,N_45980);
or U48016 (N_48016,N_46349,N_47132);
and U48017 (N_48017,N_46728,N_47350);
and U48018 (N_48018,N_46102,N_47189);
nand U48019 (N_48019,N_45961,N_46218);
or U48020 (N_48020,N_47456,N_46943);
or U48021 (N_48021,N_45106,N_46723);
xnor U48022 (N_48022,N_46639,N_46213);
and U48023 (N_48023,N_45708,N_45417);
nand U48024 (N_48024,N_45178,N_46400);
and U48025 (N_48025,N_45030,N_45924);
nand U48026 (N_48026,N_45987,N_45060);
xor U48027 (N_48027,N_45939,N_46772);
nor U48028 (N_48028,N_45190,N_46007);
nand U48029 (N_48029,N_46417,N_46118);
nor U48030 (N_48030,N_45278,N_46465);
or U48031 (N_48031,N_46567,N_46150);
or U48032 (N_48032,N_45095,N_46206);
nor U48033 (N_48033,N_47363,N_45160);
nand U48034 (N_48034,N_45498,N_45210);
and U48035 (N_48035,N_45028,N_45742);
nor U48036 (N_48036,N_47328,N_46114);
nand U48037 (N_48037,N_46296,N_45755);
nor U48038 (N_48038,N_45422,N_47072);
and U48039 (N_48039,N_46927,N_46143);
and U48040 (N_48040,N_46179,N_47156);
xnor U48041 (N_48041,N_46784,N_46165);
nand U48042 (N_48042,N_45463,N_46484);
nor U48043 (N_48043,N_45113,N_45647);
or U48044 (N_48044,N_45844,N_45919);
nor U48045 (N_48045,N_45314,N_45303);
xor U48046 (N_48046,N_46998,N_45998);
nand U48047 (N_48047,N_46821,N_45048);
or U48048 (N_48048,N_47406,N_46374);
or U48049 (N_48049,N_47432,N_46458);
and U48050 (N_48050,N_45911,N_46231);
and U48051 (N_48051,N_45092,N_45361);
or U48052 (N_48052,N_46759,N_46538);
or U48053 (N_48053,N_46955,N_47280);
xnor U48054 (N_48054,N_47355,N_47436);
or U48055 (N_48055,N_45091,N_46137);
and U48056 (N_48056,N_47487,N_45757);
xnor U48057 (N_48057,N_46854,N_46798);
nor U48058 (N_48058,N_46133,N_45008);
and U48059 (N_48059,N_45884,N_47208);
xor U48060 (N_48060,N_45966,N_46262);
xnor U48061 (N_48061,N_46278,N_45976);
and U48062 (N_48062,N_45375,N_45556);
nand U48063 (N_48063,N_47142,N_46861);
and U48064 (N_48064,N_45850,N_46525);
nor U48065 (N_48065,N_45365,N_47351);
nand U48066 (N_48066,N_45153,N_46156);
nor U48067 (N_48067,N_45166,N_45067);
and U48068 (N_48068,N_47347,N_47333);
and U48069 (N_48069,N_47085,N_46079);
nand U48070 (N_48070,N_46347,N_47178);
and U48071 (N_48071,N_46926,N_46888);
xnor U48072 (N_48072,N_45372,N_45397);
nand U48073 (N_48073,N_45509,N_45061);
and U48074 (N_48074,N_46504,N_45545);
and U48075 (N_48075,N_46480,N_47382);
xnor U48076 (N_48076,N_46195,N_47389);
nor U48077 (N_48077,N_45057,N_47420);
nand U48078 (N_48078,N_45415,N_46128);
nor U48079 (N_48079,N_46894,N_46794);
nor U48080 (N_48080,N_47212,N_46938);
nand U48081 (N_48081,N_45635,N_45102);
xnor U48082 (N_48082,N_47014,N_47466);
xnor U48083 (N_48083,N_45342,N_45434);
xor U48084 (N_48084,N_45655,N_47253);
xnor U48085 (N_48085,N_47241,N_46986);
xor U48086 (N_48086,N_46702,N_45325);
xor U48087 (N_48087,N_46051,N_46348);
xor U48088 (N_48088,N_47345,N_45482);
or U48089 (N_48089,N_45169,N_45295);
nand U48090 (N_48090,N_47124,N_46625);
nor U48091 (N_48091,N_46536,N_45666);
or U48092 (N_48092,N_45731,N_46129);
or U48093 (N_48093,N_45802,N_47230);
nor U48094 (N_48094,N_46705,N_46510);
or U48095 (N_48095,N_45358,N_45029);
nor U48096 (N_48096,N_46047,N_46598);
nand U48097 (N_48097,N_46098,N_46291);
nand U48098 (N_48098,N_45724,N_46406);
xnor U48099 (N_48099,N_47238,N_46770);
and U48100 (N_48100,N_45288,N_45903);
xnor U48101 (N_48101,N_47114,N_46067);
nand U48102 (N_48102,N_46545,N_47029);
xnor U48103 (N_48103,N_45806,N_45098);
and U48104 (N_48104,N_45529,N_45108);
and U48105 (N_48105,N_47110,N_45425);
nor U48106 (N_48106,N_45663,N_45223);
or U48107 (N_48107,N_47126,N_46249);
and U48108 (N_48108,N_46990,N_47286);
nand U48109 (N_48109,N_47421,N_45773);
nand U48110 (N_48110,N_46024,N_45359);
and U48111 (N_48111,N_45639,N_46880);
nand U48112 (N_48112,N_45232,N_47308);
and U48113 (N_48113,N_45907,N_45018);
or U48114 (N_48114,N_45625,N_46130);
nand U48115 (N_48115,N_45254,N_45292);
nor U48116 (N_48116,N_46786,N_45170);
and U48117 (N_48117,N_46268,N_45304);
xnor U48118 (N_48118,N_45964,N_47281);
nand U48119 (N_48119,N_45902,N_45432);
xor U48120 (N_48120,N_47435,N_47034);
and U48121 (N_48121,N_45366,N_46979);
nor U48122 (N_48122,N_47459,N_46319);
and U48123 (N_48123,N_46543,N_46981);
nor U48124 (N_48124,N_46531,N_45607);
nand U48125 (N_48125,N_45071,N_45778);
nand U48126 (N_48126,N_46418,N_45955);
xor U48127 (N_48127,N_45930,N_45925);
nor U48128 (N_48128,N_45455,N_47100);
and U48129 (N_48129,N_46923,N_46050);
nor U48130 (N_48130,N_45700,N_47088);
or U48131 (N_48131,N_47356,N_47451);
or U48132 (N_48132,N_45298,N_45936);
or U48133 (N_48133,N_45371,N_47302);
xnor U48134 (N_48134,N_45038,N_46386);
nand U48135 (N_48135,N_45675,N_45684);
nor U48136 (N_48136,N_47103,N_47384);
or U48137 (N_48137,N_47215,N_45940);
and U48138 (N_48138,N_47316,N_47130);
xnor U48139 (N_48139,N_47388,N_45401);
or U48140 (N_48140,N_45563,N_46607);
and U48141 (N_48141,N_45997,N_45735);
or U48142 (N_48142,N_45468,N_46230);
and U48143 (N_48143,N_46473,N_46592);
nor U48144 (N_48144,N_46429,N_46039);
or U48145 (N_48145,N_45832,N_47417);
or U48146 (N_48146,N_47199,N_46530);
nor U48147 (N_48147,N_46706,N_47458);
xnor U48148 (N_48148,N_47343,N_46451);
xor U48149 (N_48149,N_46063,N_45578);
or U48150 (N_48150,N_46701,N_45631);
and U48151 (N_48151,N_47294,N_47039);
nor U48152 (N_48152,N_45090,N_46738);
and U48153 (N_48153,N_45234,N_45559);
nand U48154 (N_48154,N_47027,N_45507);
xor U48155 (N_48155,N_45612,N_46253);
nand U48156 (N_48156,N_45793,N_45676);
xor U48157 (N_48157,N_45551,N_45489);
nor U48158 (N_48158,N_45573,N_46690);
or U48159 (N_48159,N_46479,N_46434);
nand U48160 (N_48160,N_46959,N_46116);
nand U48161 (N_48161,N_45792,N_46096);
and U48162 (N_48162,N_46962,N_47358);
xnor U48163 (N_48163,N_46224,N_46617);
or U48164 (N_48164,N_45485,N_45419);
nor U48165 (N_48165,N_46459,N_46609);
xor U48166 (N_48166,N_46633,N_46867);
nand U48167 (N_48167,N_46647,N_47053);
xnor U48168 (N_48168,N_46330,N_46221);
nand U48169 (N_48169,N_47202,N_46897);
nor U48170 (N_48170,N_47290,N_45937);
nand U48171 (N_48171,N_45540,N_46117);
or U48172 (N_48172,N_47309,N_46840);
nand U48173 (N_48173,N_47344,N_46197);
or U48174 (N_48174,N_46600,N_45591);
or U48175 (N_48175,N_46653,N_46896);
and U48176 (N_48176,N_45641,N_47480);
nor U48177 (N_48177,N_46407,N_46948);
and U48178 (N_48178,N_45461,N_46565);
xor U48179 (N_48179,N_45587,N_46266);
or U48180 (N_48180,N_47049,N_47321);
nor U48181 (N_48181,N_47184,N_47060);
nand U48182 (N_48182,N_45535,N_47023);
nor U48183 (N_48183,N_46352,N_47265);
or U48184 (N_48184,N_47147,N_46520);
nor U48185 (N_48185,N_46553,N_46293);
nand U48186 (N_48186,N_47074,N_45080);
xor U48187 (N_48187,N_45313,N_45389);
or U48188 (N_48188,N_46215,N_47270);
or U48189 (N_48189,N_45865,N_45367);
and U48190 (N_48190,N_47386,N_45268);
or U48191 (N_48191,N_47166,N_45072);
or U48192 (N_48192,N_46254,N_46198);
nor U48193 (N_48193,N_45125,N_47434);
xnor U48194 (N_48194,N_45944,N_47370);
and U48195 (N_48195,N_46367,N_45042);
nor U48196 (N_48196,N_46983,N_46637);
xor U48197 (N_48197,N_45058,N_46913);
and U48198 (N_48198,N_46606,N_45270);
xor U48199 (N_48199,N_46751,N_47313);
and U48200 (N_48200,N_47185,N_47096);
xnor U48201 (N_48201,N_47233,N_45348);
or U48202 (N_48202,N_45493,N_46831);
nand U48203 (N_48203,N_45337,N_47465);
nor U48204 (N_48204,N_45480,N_46171);
xor U48205 (N_48205,N_45965,N_46049);
nand U48206 (N_48206,N_47221,N_46827);
nor U48207 (N_48207,N_45673,N_46891);
xnor U48208 (N_48208,N_45014,N_45135);
xor U48209 (N_48209,N_45009,N_46448);
nand U48210 (N_48210,N_45993,N_47425);
and U48211 (N_48211,N_47258,N_45584);
or U48212 (N_48212,N_45957,N_45743);
nand U48213 (N_48213,N_45499,N_46376);
nor U48214 (N_48214,N_47493,N_45041);
nor U48215 (N_48215,N_45909,N_47285);
nor U48216 (N_48216,N_45334,N_47407);
xor U48217 (N_48217,N_45790,N_46984);
nor U48218 (N_48218,N_46212,N_46342);
and U48219 (N_48219,N_46285,N_46546);
nor U48220 (N_48220,N_47449,N_45124);
and U48221 (N_48221,N_46372,N_47172);
or U48222 (N_48222,N_46302,N_45460);
or U48223 (N_48223,N_45848,N_47390);
xor U48224 (N_48224,N_45196,N_46123);
or U48225 (N_48225,N_46491,N_45478);
xnor U48226 (N_48226,N_46611,N_46997);
xnor U48227 (N_48227,N_45839,N_47077);
nand U48228 (N_48228,N_46086,N_47430);
or U48229 (N_48229,N_45302,N_45604);
or U48230 (N_48230,N_46698,N_46855);
xnor U48231 (N_48231,N_46088,N_47259);
nand U48232 (N_48232,N_47450,N_46203);
nor U48233 (N_48233,N_46666,N_46402);
or U48234 (N_48234,N_47173,N_47423);
or U48235 (N_48235,N_46126,N_46667);
and U48236 (N_48236,N_46977,N_46766);
and U48237 (N_48237,N_45845,N_46655);
and U48238 (N_48238,N_46564,N_45035);
nand U48239 (N_48239,N_47026,N_47412);
and U48240 (N_48240,N_47374,N_45981);
nor U48241 (N_48241,N_45165,N_46482);
nor U48242 (N_48242,N_47099,N_45215);
nand U48243 (N_48243,N_46036,N_45693);
xnor U48244 (N_48244,N_46583,N_45382);
xnor U48245 (N_48245,N_45864,N_45296);
nand U48246 (N_48246,N_47194,N_46324);
nand U48247 (N_48247,N_46924,N_47231);
or U48248 (N_48248,N_46008,N_47385);
xor U48249 (N_48249,N_45943,N_45992);
or U48250 (N_48250,N_46155,N_45336);
and U48251 (N_48251,N_45488,N_45991);
or U48252 (N_48252,N_46321,N_46882);
and U48253 (N_48253,N_46624,N_47304);
nor U48254 (N_48254,N_47310,N_45438);
and U48255 (N_48255,N_46290,N_46961);
and U48256 (N_48256,N_46581,N_47139);
or U48257 (N_48257,N_47057,N_47380);
and U48258 (N_48258,N_45293,N_47472);
xor U48259 (N_48259,N_45811,N_46808);
or U48260 (N_48260,N_46250,N_47112);
nor U48261 (N_48261,N_46843,N_45077);
nand U48262 (N_48262,N_47095,N_46189);
nor U48263 (N_48263,N_45149,N_45123);
xnor U48264 (N_48264,N_45874,N_46560);
nor U48265 (N_48265,N_46872,N_45275);
or U48266 (N_48266,N_46208,N_45660);
nand U48267 (N_48267,N_47146,N_47312);
and U48268 (N_48268,N_45201,N_46903);
nand U48269 (N_48269,N_46992,N_45033);
and U48270 (N_48270,N_45290,N_46041);
nor U48271 (N_48271,N_46659,N_47393);
and U48272 (N_48272,N_46027,N_45661);
nand U48273 (N_48273,N_47078,N_45497);
and U48274 (N_48274,N_46436,N_46069);
nor U48275 (N_48275,N_46754,N_46901);
nor U48276 (N_48276,N_45129,N_47426);
xnor U48277 (N_48277,N_45341,N_45632);
or U48278 (N_48278,N_46969,N_46577);
nor U48279 (N_48279,N_45436,N_45526);
or U48280 (N_48280,N_46661,N_45420);
nand U48281 (N_48281,N_45249,N_45774);
xnor U48282 (N_48282,N_47477,N_46585);
nand U48283 (N_48283,N_46488,N_45096);
nand U48284 (N_48284,N_46106,N_45883);
or U48285 (N_48285,N_47148,N_46850);
nand U48286 (N_48286,N_45105,N_45780);
or U48287 (N_48287,N_46238,N_46748);
or U48288 (N_48288,N_46275,N_46248);
xnor U48289 (N_48289,N_46640,N_45552);
and U48290 (N_48290,N_45350,N_46952);
nor U48291 (N_48291,N_46886,N_47102);
and U48292 (N_48292,N_46644,N_45546);
xnor U48293 (N_48293,N_46900,N_45207);
nand U48294 (N_48294,N_47291,N_46973);
xor U48295 (N_48295,N_46996,N_46091);
and U48296 (N_48296,N_46255,N_45112);
or U48297 (N_48297,N_46413,N_46362);
or U48298 (N_48298,N_47318,N_47080);
nor U48299 (N_48299,N_46582,N_46703);
nor U48300 (N_48300,N_45076,N_45767);
xor U48301 (N_48301,N_45645,N_45829);
and U48302 (N_48302,N_45216,N_46828);
and U48303 (N_48303,N_45935,N_45648);
xor U48304 (N_48304,N_46087,N_47223);
or U48305 (N_48305,N_46111,N_46134);
nor U48306 (N_48306,N_46053,N_46236);
xor U48307 (N_48307,N_46322,N_45914);
nand U48308 (N_48308,N_46030,N_46070);
or U48309 (N_48309,N_45144,N_46863);
xnor U48310 (N_48310,N_46807,N_47457);
nand U48311 (N_48311,N_46401,N_47128);
and U48312 (N_48312,N_46720,N_46949);
nand U48313 (N_48313,N_46115,N_45220);
nor U48314 (N_48314,N_47107,N_46528);
and U48315 (N_48315,N_45383,N_47135);
nor U48316 (N_48316,N_46328,N_45386);
and U48317 (N_48317,N_47168,N_45286);
xnor U48318 (N_48318,N_46819,N_45568);
or U48319 (N_48319,N_46222,N_47162);
nor U48320 (N_48320,N_45217,N_47445);
or U48321 (N_48321,N_46345,N_45579);
and U48322 (N_48322,N_47242,N_46746);
or U48323 (N_48323,N_46175,N_47399);
nor U48324 (N_48324,N_45862,N_46162);
nor U48325 (N_48325,N_46353,N_45172);
and U48326 (N_48326,N_45652,N_46163);
or U48327 (N_48327,N_45464,N_45360);
or U48328 (N_48328,N_47279,N_46409);
and U48329 (N_48329,N_46833,N_45928);
and U48330 (N_48330,N_46260,N_45320);
nand U48331 (N_48331,N_45967,N_46441);
nand U48332 (N_48332,N_46660,N_45081);
nor U48333 (N_48333,N_45771,N_46461);
xor U48334 (N_48334,N_46713,N_45809);
and U48335 (N_48335,N_46389,N_46868);
nand U48336 (N_48336,N_45782,N_46885);
and U48337 (N_48337,N_45870,N_45549);
nor U48338 (N_48338,N_46332,N_47245);
and U48339 (N_48339,N_46714,N_45753);
xnor U48340 (N_48340,N_45979,N_46876);
nor U48341 (N_48341,N_45525,N_45115);
xor U48342 (N_48342,N_46277,N_46928);
or U48343 (N_48343,N_47340,N_45483);
xor U48344 (N_48344,N_45206,N_45380);
or U48345 (N_48345,N_47263,N_45147);
nor U48346 (N_48346,N_45712,N_46512);
and U48347 (N_48347,N_45636,N_46902);
and U48348 (N_48348,N_45711,N_45175);
and U48349 (N_48349,N_46002,N_46103);
nor U48350 (N_48350,N_45830,N_46641);
or U48351 (N_48351,N_47255,N_46925);
nand U48352 (N_48352,N_45656,N_46464);
nand U48353 (N_48353,N_46297,N_47365);
xnor U48354 (N_48354,N_45356,N_47174);
nor U48355 (N_48355,N_45659,N_45710);
or U48356 (N_48356,N_45136,N_46235);
nand U48357 (N_48357,N_45134,N_45779);
and U48358 (N_48358,N_45374,N_46258);
xor U48359 (N_48359,N_47167,N_46185);
or U48360 (N_48360,N_46777,N_46501);
nor U48361 (N_48361,N_47448,N_45186);
or U48362 (N_48362,N_46037,N_45906);
nor U48363 (N_48363,N_46846,N_45836);
xnor U48364 (N_48364,N_45173,N_45398);
xor U48365 (N_48365,N_45837,N_46763);
and U48366 (N_48366,N_46507,N_47453);
or U48367 (N_48367,N_45565,N_46358);
or U48368 (N_48368,N_46883,N_46300);
or U48369 (N_48369,N_46733,N_45544);
or U48370 (N_48370,N_47093,N_46430);
nor U48371 (N_48371,N_45628,N_47446);
xor U48372 (N_48372,N_45005,N_47004);
and U48373 (N_48373,N_46980,N_45597);
xor U48374 (N_48374,N_46697,N_45754);
or U48375 (N_48375,N_47190,N_46719);
xor U48376 (N_48376,N_45150,N_46313);
nor U48377 (N_48377,N_46074,N_45168);
nand U48378 (N_48378,N_47237,N_46556);
or U48379 (N_48379,N_46789,N_46848);
nor U48380 (N_48380,N_46160,N_45151);
or U48381 (N_48381,N_47186,N_46124);
nand U48382 (N_48382,N_47021,N_46026);
and U48383 (N_48383,N_47273,N_45324);
xor U48384 (N_48384,N_45174,N_47266);
nor U48385 (N_48385,N_45472,N_46836);
nand U48386 (N_48386,N_47033,N_45736);
nand U48387 (N_48387,N_45614,N_46865);
nand U48388 (N_48388,N_46557,N_45875);
or U48389 (N_48389,N_47117,N_47236);
xor U48390 (N_48390,N_45158,N_45250);
nor U48391 (N_48391,N_45983,N_45692);
and U48392 (N_48392,N_45495,N_45680);
xnor U48393 (N_48393,N_46097,N_46455);
nand U48394 (N_48394,N_47405,N_45500);
nand U48395 (N_48395,N_45859,N_47006);
and U48396 (N_48396,N_45473,N_46233);
xor U48397 (N_48397,N_46014,N_46550);
and U48398 (N_48398,N_47214,N_47138);
nand U48399 (N_48399,N_45036,N_46357);
or U48400 (N_48400,N_45886,N_45611);
xor U48401 (N_48401,N_45872,N_47137);
nand U48402 (N_48402,N_45951,N_47381);
or U48403 (N_48403,N_46832,N_45685);
and U48404 (N_48404,N_47123,N_45423);
nand U48405 (N_48405,N_45338,N_47044);
or U48406 (N_48406,N_45469,N_46064);
nor U48407 (N_48407,N_46539,N_47461);
or U48408 (N_48408,N_46326,N_46351);
xnor U48409 (N_48409,N_46526,N_46757);
or U48410 (N_48410,N_47229,N_45226);
and U48411 (N_48411,N_45240,N_45496);
or U48412 (N_48412,N_45308,N_46856);
or U48413 (N_48413,N_47030,N_46396);
and U48414 (N_48414,N_46579,N_45089);
or U48415 (N_48415,N_47040,N_45440);
nand U48416 (N_48416,N_46192,N_45759);
and U48417 (N_48417,N_45392,N_46940);
nor U48418 (N_48418,N_46511,N_45315);
xnor U48419 (N_48419,N_46125,N_46346);
nand U48420 (N_48420,N_45078,N_47129);
nor U48421 (N_48421,N_45533,N_46586);
or U48422 (N_48422,N_46446,N_45084);
and U48423 (N_48423,N_45479,N_46494);
or U48424 (N_48424,N_46424,N_47025);
nor U48425 (N_48425,N_45717,N_46533);
or U48426 (N_48426,N_46673,N_45847);
nand U48427 (N_48427,N_47151,N_46740);
nand U48428 (N_48428,N_47158,N_45410);
nor U48429 (N_48429,N_46042,N_47427);
nor U48430 (N_48430,N_46873,N_46247);
or U48431 (N_48431,N_46005,N_46496);
nand U48432 (N_48432,N_46469,N_46001);
nor U48433 (N_48433,N_45938,N_47357);
nand U48434 (N_48434,N_46761,N_45448);
and U48435 (N_48435,N_46519,N_47367);
and U48436 (N_48436,N_47235,N_45828);
or U48437 (N_48437,N_45554,N_46568);
or U48438 (N_48438,N_45300,N_47043);
or U48439 (N_48439,N_45522,N_45923);
or U48440 (N_48440,N_46677,N_45451);
xnor U48441 (N_48441,N_45449,N_46356);
xnor U48442 (N_48442,N_47218,N_46765);
nand U48443 (N_48443,N_47396,N_46010);
nand U48444 (N_48444,N_46696,N_46481);
nand U48445 (N_48445,N_45527,N_45745);
xor U48446 (N_48446,N_45729,N_47277);
and U48447 (N_48447,N_47101,N_45678);
nor U48448 (N_48448,N_47305,N_45354);
xnor U48449 (N_48449,N_45901,N_46729);
or U48450 (N_48450,N_46364,N_45221);
and U48451 (N_48451,N_45751,N_45775);
nand U48452 (N_48452,N_47063,N_45114);
or U48453 (N_48453,N_45233,N_46373);
nand U48454 (N_48454,N_46360,N_47274);
xnor U48455 (N_48455,N_46881,N_46283);
and U48456 (N_48456,N_46804,N_45594);
xor U48457 (N_48457,N_46387,N_45161);
and U48458 (N_48458,N_46652,N_46428);
or U48459 (N_48459,N_47163,N_45762);
nand U48460 (N_48460,N_46791,N_45869);
and U48461 (N_48461,N_47217,N_45218);
nand U48462 (N_48462,N_45689,N_46841);
nor U48463 (N_48463,N_45824,N_47342);
xnor U48464 (N_48464,N_46144,N_45408);
nand U48465 (N_48465,N_46032,N_45789);
nand U48466 (N_48466,N_45427,N_47141);
nand U48467 (N_48467,N_47192,N_46439);
nor U48468 (N_48468,N_46572,N_45630);
or U48469 (N_48469,N_45603,N_45586);
xor U48470 (N_48470,N_45421,N_45191);
xnor U48471 (N_48471,N_46820,N_46522);
xor U48472 (N_48472,N_46654,N_46964);
nor U48473 (N_48473,N_47433,N_45456);
or U48474 (N_48474,N_45212,N_46281);
and U48475 (N_48475,N_45733,N_45117);
nor U48476 (N_48476,N_45142,N_45861);
or U48477 (N_48477,N_45384,N_45831);
nand U48478 (N_48478,N_46408,N_46930);
and U48479 (N_48479,N_46471,N_46942);
nor U48480 (N_48480,N_45052,N_46110);
and U48481 (N_48481,N_46657,N_45491);
nand U48482 (N_48482,N_47002,N_46935);
xor U48483 (N_48483,N_46892,N_45395);
nor U48484 (N_48484,N_46368,N_46183);
or U48485 (N_48485,N_45088,N_46243);
nor U48486 (N_48486,N_45291,N_46227);
and U48487 (N_48487,N_46335,N_46187);
nand U48488 (N_48488,N_46689,N_45347);
nor U48489 (N_48489,N_47180,N_46487);
xnor U48490 (N_48490,N_45285,N_46779);
and U48491 (N_48491,N_46276,N_45004);
or U48492 (N_48492,N_45732,N_45159);
and U48493 (N_48493,N_46910,N_46061);
and U48494 (N_48494,N_46397,N_45888);
or U48495 (N_48495,N_45044,N_47127);
xor U48496 (N_48496,N_47275,N_47452);
nand U48497 (N_48497,N_47056,N_45245);
and U48498 (N_48498,N_46311,N_47413);
and U48499 (N_48499,N_46905,N_46812);
xnor U48500 (N_48500,N_47490,N_45726);
or U48501 (N_48501,N_46616,N_46537);
and U48502 (N_48502,N_46614,N_45803);
nand U48503 (N_48503,N_46385,N_45203);
nor U48504 (N_48504,N_46830,N_45695);
or U48505 (N_48505,N_45185,N_45279);
or U48506 (N_48506,N_46172,N_46366);
nand U48507 (N_48507,N_45323,N_45777);
xor U48508 (N_48508,N_47249,N_47051);
and U48509 (N_48509,N_46059,N_47239);
nor U48510 (N_48510,N_47076,N_45222);
or U48511 (N_48511,N_46246,N_45003);
nand U48512 (N_48512,N_45503,N_45898);
nand U48513 (N_48513,N_47094,N_45642);
nor U48514 (N_48514,N_45063,N_46593);
and U48515 (N_48515,N_47089,N_45915);
or U48516 (N_48516,N_45511,N_47024);
xor U48517 (N_48517,N_46011,N_47485);
xor U48518 (N_48518,N_46460,N_46167);
xor U48519 (N_48519,N_45927,N_45085);
or U48520 (N_48520,N_47111,N_46383);
nor U48521 (N_48521,N_46604,N_45069);
or U48522 (N_48522,N_45629,N_45506);
or U48523 (N_48523,N_47204,N_45357);
nand U48524 (N_48524,N_45613,N_46802);
xor U48525 (N_48525,N_46951,N_45653);
nor U48526 (N_48526,N_45385,N_47276);
and U48527 (N_48527,N_45534,N_47401);
xor U48528 (N_48528,N_45505,N_46174);
or U48529 (N_48529,N_45394,N_47462);
and U48530 (N_48530,N_46874,N_46815);
and U48531 (N_48531,N_45335,N_46191);
and U48532 (N_48532,N_46365,N_45258);
or U48533 (N_48533,N_45023,N_45973);
nor U48534 (N_48534,N_46450,N_46432);
or U48535 (N_48535,N_46263,N_47250);
nor U48536 (N_48536,N_46575,N_45900);
and U48537 (N_48537,N_47284,N_46839);
xnor U48538 (N_48538,N_46398,N_46388);
and U48539 (N_48539,N_47105,N_45634);
nor U48540 (N_48540,N_45163,N_45833);
nand U48541 (N_48541,N_45053,N_45402);
or U48542 (N_48542,N_47323,N_47134);
and U48543 (N_48543,N_45651,N_45926);
nand U48544 (N_48544,N_46075,N_45015);
xnor U48545 (N_48545,N_46454,N_45760);
nand U48546 (N_48546,N_46242,N_46456);
nand U48547 (N_48547,N_45820,N_46960);
and U48548 (N_48548,N_46547,N_45699);
nor U48549 (N_48549,N_45929,N_47271);
nand U48550 (N_48550,N_45986,N_46315);
nand U48551 (N_48551,N_46314,N_45851);
xnor U48552 (N_48552,N_46419,N_47332);
or U48553 (N_48553,N_45590,N_45890);
or U48554 (N_48554,N_47140,N_46632);
or U48555 (N_48555,N_45574,N_46138);
xnor U48556 (N_48556,N_46817,N_46421);
nand U48557 (N_48557,N_46638,N_45588);
or U48558 (N_48558,N_45800,N_45761);
xnor U48559 (N_48559,N_45466,N_47443);
and U48560 (N_48560,N_45010,N_46490);
nor U48561 (N_48561,N_46781,N_47133);
nor U48562 (N_48562,N_46340,N_45281);
nor U48563 (N_48563,N_46094,N_46282);
nand U48564 (N_48564,N_45260,N_46809);
nand U48565 (N_48565,N_46629,N_45860);
and U48566 (N_48566,N_45722,N_47041);
or U48567 (N_48567,N_45994,N_45672);
or U48568 (N_48568,N_46622,N_46842);
nand U48569 (N_48569,N_45531,N_46286);
nor U48570 (N_48570,N_45682,N_46744);
or U48571 (N_48571,N_47454,N_45741);
nand U48572 (N_48572,N_45719,N_47059);
xnor U48573 (N_48573,N_46978,N_45738);
nor U48574 (N_48574,N_45064,N_47362);
and U48575 (N_48575,N_45988,N_45605);
or U48576 (N_48576,N_45853,N_45610);
nand U48577 (N_48577,N_45111,N_45941);
nand U48578 (N_48578,N_45817,N_46914);
nand U48579 (N_48579,N_46672,N_46145);
nand U48580 (N_48580,N_46493,N_46425);
xor U48581 (N_48581,N_47084,N_46931);
nand U48582 (N_48582,N_45687,N_47058);
nor U48583 (N_48583,N_45225,N_46965);
nand U48584 (N_48584,N_46084,N_45429);
or U48585 (N_48585,N_46917,N_46320);
and U48586 (N_48586,N_46057,N_45016);
xor U48587 (N_48587,N_45236,N_46805);
xor U48588 (N_48588,N_47339,N_45403);
nand U48589 (N_48589,N_46858,N_45059);
and U48590 (N_48590,N_45477,N_46548);
or U48591 (N_48591,N_46558,N_46176);
or U48592 (N_48592,N_46613,N_46257);
or U48593 (N_48593,N_46015,N_46076);
nor U48594 (N_48594,N_45644,N_45932);
xnor U48595 (N_48595,N_47153,N_46065);
or U48596 (N_48596,N_46693,N_46095);
or U48597 (N_48597,N_45958,N_46678);
or U48598 (N_48598,N_46825,N_46737);
xnor U48599 (N_48599,N_45208,N_47079);
nand U48600 (N_48600,N_45619,N_45750);
nand U48601 (N_48601,N_46709,N_46722);
or U48602 (N_48602,N_46670,N_45027);
xor U48603 (N_48603,N_46085,N_45043);
xor U48604 (N_48604,N_46200,N_46477);
nand U48605 (N_48605,N_47042,N_46060);
xor U48606 (N_48606,N_46707,N_46475);
xor U48607 (N_48607,N_45271,N_45025);
nor U48608 (N_48608,N_45795,N_45441);
or U48609 (N_48609,N_46305,N_47016);
nor U48610 (N_48610,N_45740,N_45164);
nand U48611 (N_48611,N_45933,N_45133);
nor U48612 (N_48612,N_46338,N_46142);
or U48613 (N_48613,N_46608,N_45252);
or U48614 (N_48614,N_46083,N_45247);
and U48615 (N_48615,N_47447,N_45065);
and U48616 (N_48616,N_46184,N_46785);
xnor U48617 (N_48617,N_46420,N_46587);
and U48618 (N_48618,N_45858,N_45816);
and U48619 (N_48619,N_46974,N_47479);
and U48620 (N_48620,N_46664,N_46164);
nand U48621 (N_48621,N_45197,N_45665);
and U48622 (N_48622,N_46552,N_47369);
nand U48623 (N_48623,N_46048,N_46650);
or U48624 (N_48624,N_45442,N_47240);
xor U48625 (N_48625,N_47028,N_45770);
and U48626 (N_48626,N_47193,N_45705);
nor U48627 (N_48627,N_45074,N_47203);
nand U48628 (N_48628,N_46468,N_46228);
and U48629 (N_48629,N_45364,N_45140);
nor U48630 (N_48630,N_46800,N_46769);
xor U48631 (N_48631,N_45520,N_46803);
nor U48632 (N_48632,N_45494,N_46818);
nand U48633 (N_48633,N_46612,N_47287);
or U48634 (N_48634,N_47296,N_46988);
or U48635 (N_48635,N_45409,N_46169);
or U48636 (N_48636,N_47411,N_47073);
and U48637 (N_48637,N_45213,N_45825);
nand U48638 (N_48638,N_45328,N_47439);
nor U48639 (N_48639,N_45670,N_46895);
nor U48640 (N_48640,N_47361,N_46963);
or U48641 (N_48641,N_45703,N_45269);
nand U48642 (N_48642,N_45857,N_46590);
nor U48643 (N_48643,N_45339,N_46422);
or U48644 (N_48644,N_47121,N_46915);
xor U48645 (N_48645,N_46331,N_47414);
or U48646 (N_48646,N_46390,N_47219);
nand U48647 (N_48647,N_45118,N_46623);
nor U48648 (N_48648,N_46476,N_45814);
or U48649 (N_48649,N_45887,N_45954);
and U48650 (N_48650,N_45256,N_45430);
nand U48651 (N_48651,N_45748,N_46107);
and U48652 (N_48652,N_45039,N_46845);
or U48653 (N_48653,N_45224,N_45119);
xor U48654 (N_48654,N_46310,N_46466);
or U48655 (N_48655,N_47062,N_45571);
or U48656 (N_48656,N_46170,N_46918);
and U48657 (N_48657,N_46561,N_46739);
nand U48658 (N_48658,N_45608,N_46500);
nand U48659 (N_48659,N_47484,N_47012);
nand U48660 (N_48660,N_45002,N_46648);
nor U48661 (N_48661,N_46139,N_45416);
and U48662 (N_48662,N_45317,N_45769);
and U48663 (N_48663,N_45804,N_45127);
xor U48664 (N_48664,N_45576,N_46716);
and U48665 (N_48665,N_47035,N_46223);
and U48666 (N_48666,N_47314,N_46681);
or U48667 (N_48667,N_46274,N_45934);
and U48668 (N_48668,N_46993,N_47307);
nand U48669 (N_48669,N_47211,N_45101);
nand U48670 (N_48670,N_46280,N_46715);
nand U48671 (N_48671,N_47428,N_45897);
or U48672 (N_48672,N_46899,N_45012);
and U48673 (N_48673,N_45424,N_45714);
nor U48674 (N_48674,N_46445,N_45116);
or U48675 (N_48675,N_45971,N_47400);
or U48676 (N_48676,N_46532,N_46824);
xnor U48677 (N_48677,N_45823,N_47136);
nor U48678 (N_48678,N_47000,N_45265);
or U48679 (N_48679,N_45103,N_46486);
nand U48680 (N_48680,N_47441,N_47061);
and U48681 (N_48681,N_46570,N_46671);
xor U48682 (N_48682,N_46158,N_47431);
or U48683 (N_48683,N_45146,N_45011);
nand U48684 (N_48684,N_46485,N_46649);
and U48685 (N_48685,N_46591,N_47419);
or U48686 (N_48686,N_45387,N_45821);
nor U48687 (N_48687,N_45066,N_45475);
nor U48688 (N_48688,N_46392,N_46109);
nand U48689 (N_48689,N_46350,N_47264);
nand U48690 (N_48690,N_47306,N_46851);
and U48691 (N_48691,N_45000,N_46251);
nor U48692 (N_48692,N_46194,N_46021);
nor U48693 (N_48693,N_47289,N_46483);
nand U48694 (N_48694,N_46146,N_45445);
and U48695 (N_48695,N_45362,N_46055);
and U48696 (N_48696,N_46578,N_45867);
and U48697 (N_48697,N_45209,N_47383);
nor U48698 (N_48698,N_45156,N_46893);
nand U48699 (N_48699,N_46985,N_46799);
xor U48700 (N_48700,N_45996,N_46529);
or U48701 (N_48701,N_45331,N_47159);
or U48702 (N_48702,N_46369,N_47091);
or U48703 (N_48703,N_45891,N_46551);
or U48704 (N_48704,N_47018,N_45723);
nand U48705 (N_48705,N_46056,N_46544);
or U48706 (N_48706,N_45181,N_46776);
and U48707 (N_48707,N_45640,N_47460);
nand U48708 (N_48708,N_45921,N_45251);
or U48709 (N_48709,N_46603,N_45107);
nand U48710 (N_48710,N_47181,N_46217);
nand U48711 (N_48711,N_47311,N_46444);
xnor U48712 (N_48712,N_45032,N_45704);
or U48713 (N_48713,N_47081,N_46308);
xor U48714 (N_48714,N_46684,N_46683);
and U48715 (N_48715,N_45749,N_47055);
and U48716 (N_48716,N_46068,N_45593);
xor U48717 (N_48717,N_46031,N_47329);
xnor U48718 (N_48718,N_47022,N_47471);
nand U48719 (N_48719,N_46584,N_45444);
nor U48720 (N_48720,N_46259,N_46966);
nor U48721 (N_48721,N_45791,N_46540);
and U48722 (N_48722,N_45141,N_46220);
xor U48723 (N_48723,N_46104,N_45070);
and U48724 (N_48724,N_45950,N_47491);
nand U48725 (N_48725,N_46016,N_46336);
nand U48726 (N_48726,N_46287,N_45962);
nand U48727 (N_48727,N_47322,N_47064);
and U48728 (N_48728,N_45162,N_46634);
and U48729 (N_48729,N_46646,N_46391);
xnor U48730 (N_48730,N_45620,N_47498);
nor U48731 (N_48731,N_47046,N_45322);
and U48732 (N_48732,N_47116,N_46571);
or U48733 (N_48733,N_47299,N_45626);
nor U48734 (N_48734,N_46782,N_47196);
xnor U48735 (N_48735,N_46211,N_47115);
nor U48736 (N_48736,N_46889,N_45558);
and U48737 (N_48737,N_46594,N_46853);
and U48738 (N_48738,N_45725,N_45752);
or U48739 (N_48739,N_45126,N_46437);
nor U48740 (N_48740,N_47154,N_46687);
nand U48741 (N_48741,N_45272,N_46204);
nand U48742 (N_48742,N_45333,N_46643);
nor U48743 (N_48743,N_45776,N_46380);
and U48744 (N_48744,N_45378,N_47069);
and U48745 (N_48745,N_47440,N_45512);
nand U48746 (N_48746,N_47429,N_47054);
xor U48747 (N_48747,N_45189,N_46033);
or U48748 (N_48748,N_45555,N_46878);
or U48749 (N_48749,N_47346,N_46240);
and U48750 (N_48750,N_47271,N_46383);
and U48751 (N_48751,N_47416,N_46698);
or U48752 (N_48752,N_45712,N_46683);
nor U48753 (N_48753,N_47261,N_47188);
nand U48754 (N_48754,N_45964,N_47280);
xnor U48755 (N_48755,N_45609,N_46215);
nor U48756 (N_48756,N_47082,N_45666);
nand U48757 (N_48757,N_47063,N_47417);
xor U48758 (N_48758,N_47128,N_46562);
or U48759 (N_48759,N_45658,N_46864);
or U48760 (N_48760,N_45820,N_45582);
or U48761 (N_48761,N_45337,N_46641);
or U48762 (N_48762,N_46314,N_46656);
nor U48763 (N_48763,N_46141,N_46867);
nand U48764 (N_48764,N_45942,N_46703);
nor U48765 (N_48765,N_47366,N_46084);
and U48766 (N_48766,N_46197,N_47369);
nand U48767 (N_48767,N_47392,N_45867);
and U48768 (N_48768,N_46232,N_45548);
or U48769 (N_48769,N_45592,N_46782);
or U48770 (N_48770,N_45191,N_46756);
xnor U48771 (N_48771,N_46781,N_47490);
and U48772 (N_48772,N_46774,N_46813);
nand U48773 (N_48773,N_46447,N_45934);
xor U48774 (N_48774,N_45552,N_47368);
nor U48775 (N_48775,N_45072,N_45196);
nand U48776 (N_48776,N_45222,N_46714);
nor U48777 (N_48777,N_46670,N_45178);
or U48778 (N_48778,N_46006,N_47005);
nor U48779 (N_48779,N_47245,N_46424);
or U48780 (N_48780,N_46271,N_45296);
and U48781 (N_48781,N_45630,N_46274);
and U48782 (N_48782,N_45530,N_45543);
and U48783 (N_48783,N_45198,N_45913);
nor U48784 (N_48784,N_46439,N_45208);
nand U48785 (N_48785,N_45064,N_46491);
xnor U48786 (N_48786,N_45380,N_46812);
nand U48787 (N_48787,N_45934,N_45272);
nand U48788 (N_48788,N_47024,N_45001);
nor U48789 (N_48789,N_45490,N_45730);
xor U48790 (N_48790,N_45810,N_46096);
xnor U48791 (N_48791,N_46573,N_46799);
and U48792 (N_48792,N_46612,N_45941);
xor U48793 (N_48793,N_45493,N_47422);
and U48794 (N_48794,N_47121,N_45424);
or U48795 (N_48795,N_45728,N_45145);
nand U48796 (N_48796,N_46640,N_46348);
and U48797 (N_48797,N_45429,N_45953);
xnor U48798 (N_48798,N_46770,N_45329);
and U48799 (N_48799,N_45977,N_45322);
and U48800 (N_48800,N_45108,N_45102);
and U48801 (N_48801,N_45198,N_46246);
nand U48802 (N_48802,N_45975,N_46588);
nor U48803 (N_48803,N_46219,N_45656);
xnor U48804 (N_48804,N_45495,N_45655);
or U48805 (N_48805,N_47373,N_46194);
nor U48806 (N_48806,N_47170,N_47065);
or U48807 (N_48807,N_47468,N_46522);
nor U48808 (N_48808,N_45928,N_45379);
or U48809 (N_48809,N_46552,N_45967);
nor U48810 (N_48810,N_46750,N_46991);
and U48811 (N_48811,N_45451,N_45858);
nor U48812 (N_48812,N_45892,N_45404);
nor U48813 (N_48813,N_45158,N_46710);
nand U48814 (N_48814,N_46943,N_46936);
xnor U48815 (N_48815,N_45591,N_46444);
xor U48816 (N_48816,N_46875,N_46014);
nand U48817 (N_48817,N_46560,N_46268);
xor U48818 (N_48818,N_46022,N_46627);
nand U48819 (N_48819,N_45750,N_47317);
nor U48820 (N_48820,N_47182,N_47391);
nand U48821 (N_48821,N_46444,N_46997);
and U48822 (N_48822,N_46525,N_46042);
or U48823 (N_48823,N_47004,N_45526);
xor U48824 (N_48824,N_46326,N_46821);
xnor U48825 (N_48825,N_47315,N_45864);
xor U48826 (N_48826,N_46972,N_45794);
and U48827 (N_48827,N_46968,N_45008);
xnor U48828 (N_48828,N_45311,N_45061);
xor U48829 (N_48829,N_45074,N_46158);
or U48830 (N_48830,N_46219,N_45189);
nand U48831 (N_48831,N_45717,N_47151);
xor U48832 (N_48832,N_46568,N_45229);
xnor U48833 (N_48833,N_47310,N_47264);
nand U48834 (N_48834,N_46212,N_45995);
nor U48835 (N_48835,N_45754,N_46680);
xnor U48836 (N_48836,N_47474,N_47455);
nand U48837 (N_48837,N_46981,N_46108);
nand U48838 (N_48838,N_45991,N_45449);
or U48839 (N_48839,N_45390,N_46342);
nand U48840 (N_48840,N_46031,N_47348);
or U48841 (N_48841,N_45963,N_47125);
or U48842 (N_48842,N_46192,N_46627);
xnor U48843 (N_48843,N_47176,N_46025);
or U48844 (N_48844,N_46153,N_47015);
and U48845 (N_48845,N_46714,N_45921);
or U48846 (N_48846,N_45334,N_45703);
nor U48847 (N_48847,N_45089,N_46386);
nor U48848 (N_48848,N_47454,N_46008);
xnor U48849 (N_48849,N_45981,N_46975);
nor U48850 (N_48850,N_46434,N_47394);
xor U48851 (N_48851,N_46514,N_46276);
nor U48852 (N_48852,N_45747,N_45157);
nand U48853 (N_48853,N_46698,N_46128);
and U48854 (N_48854,N_46417,N_46437);
and U48855 (N_48855,N_45843,N_47107);
nor U48856 (N_48856,N_45976,N_46605);
or U48857 (N_48857,N_47402,N_47030);
nand U48858 (N_48858,N_45063,N_45921);
nand U48859 (N_48859,N_47305,N_45992);
xor U48860 (N_48860,N_46332,N_46165);
and U48861 (N_48861,N_46676,N_46283);
or U48862 (N_48862,N_46944,N_47298);
xnor U48863 (N_48863,N_46070,N_46658);
and U48864 (N_48864,N_47256,N_46663);
and U48865 (N_48865,N_46032,N_45371);
nor U48866 (N_48866,N_47442,N_46395);
nor U48867 (N_48867,N_45303,N_46255);
or U48868 (N_48868,N_46978,N_47115);
and U48869 (N_48869,N_46180,N_46987);
nor U48870 (N_48870,N_46469,N_45187);
nor U48871 (N_48871,N_46856,N_47277);
or U48872 (N_48872,N_45836,N_45206);
nor U48873 (N_48873,N_46183,N_46182);
and U48874 (N_48874,N_47294,N_47109);
and U48875 (N_48875,N_46460,N_46674);
xnor U48876 (N_48876,N_47452,N_46031);
nor U48877 (N_48877,N_47448,N_45718);
nor U48878 (N_48878,N_45423,N_45071);
nand U48879 (N_48879,N_45132,N_47445);
nand U48880 (N_48880,N_46189,N_46025);
and U48881 (N_48881,N_46198,N_47257);
nand U48882 (N_48882,N_46160,N_45326);
or U48883 (N_48883,N_46869,N_45027);
and U48884 (N_48884,N_45915,N_47333);
nand U48885 (N_48885,N_46413,N_45981);
nand U48886 (N_48886,N_46808,N_45425);
nor U48887 (N_48887,N_45050,N_45213);
and U48888 (N_48888,N_47129,N_45711);
xnor U48889 (N_48889,N_46053,N_45524);
or U48890 (N_48890,N_46164,N_46408);
or U48891 (N_48891,N_45550,N_46621);
xor U48892 (N_48892,N_46145,N_45052);
or U48893 (N_48893,N_46780,N_46025);
xnor U48894 (N_48894,N_47253,N_46478);
and U48895 (N_48895,N_45154,N_45646);
xnor U48896 (N_48896,N_47046,N_45552);
nor U48897 (N_48897,N_45527,N_47171);
and U48898 (N_48898,N_46774,N_46288);
and U48899 (N_48899,N_45939,N_46990);
nand U48900 (N_48900,N_46337,N_45868);
or U48901 (N_48901,N_45288,N_45961);
nor U48902 (N_48902,N_47155,N_46004);
or U48903 (N_48903,N_46898,N_45718);
nor U48904 (N_48904,N_46093,N_45543);
and U48905 (N_48905,N_45728,N_45028);
or U48906 (N_48906,N_47286,N_46412);
nor U48907 (N_48907,N_46240,N_45551);
nand U48908 (N_48908,N_47230,N_45538);
nand U48909 (N_48909,N_46252,N_47111);
xnor U48910 (N_48910,N_45144,N_45781);
nor U48911 (N_48911,N_45610,N_46480);
and U48912 (N_48912,N_46387,N_45003);
and U48913 (N_48913,N_46995,N_46963);
xor U48914 (N_48914,N_46296,N_45400);
xor U48915 (N_48915,N_46481,N_47308);
xor U48916 (N_48916,N_47028,N_45475);
and U48917 (N_48917,N_45490,N_46889);
or U48918 (N_48918,N_45797,N_45454);
nor U48919 (N_48919,N_45112,N_45755);
or U48920 (N_48920,N_47258,N_45670);
xor U48921 (N_48921,N_45889,N_46738);
xor U48922 (N_48922,N_47212,N_45642);
nand U48923 (N_48923,N_46017,N_46450);
xnor U48924 (N_48924,N_45846,N_45143);
and U48925 (N_48925,N_47041,N_45686);
nor U48926 (N_48926,N_45580,N_46895);
nor U48927 (N_48927,N_46431,N_45205);
and U48928 (N_48928,N_45806,N_45124);
or U48929 (N_48929,N_46300,N_45831);
nor U48930 (N_48930,N_45872,N_46635);
nor U48931 (N_48931,N_45218,N_46449);
nand U48932 (N_48932,N_47334,N_47217);
and U48933 (N_48933,N_45422,N_45353);
xor U48934 (N_48934,N_46981,N_45192);
or U48935 (N_48935,N_45196,N_46410);
nand U48936 (N_48936,N_45892,N_47150);
nor U48937 (N_48937,N_45805,N_46243);
or U48938 (N_48938,N_47006,N_45914);
and U48939 (N_48939,N_47167,N_46145);
nand U48940 (N_48940,N_45186,N_45291);
or U48941 (N_48941,N_46625,N_47370);
and U48942 (N_48942,N_46264,N_45425);
and U48943 (N_48943,N_45649,N_45103);
nand U48944 (N_48944,N_47092,N_45886);
or U48945 (N_48945,N_45665,N_46583);
nor U48946 (N_48946,N_46073,N_45345);
xnor U48947 (N_48947,N_46089,N_47110);
nor U48948 (N_48948,N_45961,N_45647);
or U48949 (N_48949,N_45465,N_46021);
nor U48950 (N_48950,N_46616,N_45478);
or U48951 (N_48951,N_45758,N_46054);
nor U48952 (N_48952,N_45882,N_45393);
nand U48953 (N_48953,N_46905,N_47446);
nor U48954 (N_48954,N_47342,N_45288);
or U48955 (N_48955,N_46789,N_47172);
xor U48956 (N_48956,N_46927,N_46066);
nand U48957 (N_48957,N_47182,N_46398);
and U48958 (N_48958,N_47117,N_47119);
nor U48959 (N_48959,N_47074,N_46004);
nor U48960 (N_48960,N_46224,N_45375);
xnor U48961 (N_48961,N_45714,N_45677);
and U48962 (N_48962,N_47165,N_45976);
nand U48963 (N_48963,N_45429,N_45394);
or U48964 (N_48964,N_46327,N_45957);
xnor U48965 (N_48965,N_46192,N_45926);
nand U48966 (N_48966,N_45537,N_46718);
nor U48967 (N_48967,N_45259,N_45227);
nor U48968 (N_48968,N_45239,N_47482);
and U48969 (N_48969,N_45936,N_45666);
nor U48970 (N_48970,N_45500,N_45956);
nand U48971 (N_48971,N_46990,N_45059);
xnor U48972 (N_48972,N_45830,N_46218);
xor U48973 (N_48973,N_47309,N_46617);
xnor U48974 (N_48974,N_46107,N_46974);
and U48975 (N_48975,N_45063,N_46671);
xnor U48976 (N_48976,N_46280,N_46974);
and U48977 (N_48977,N_47326,N_46189);
xnor U48978 (N_48978,N_45063,N_45947);
or U48979 (N_48979,N_46850,N_45121);
nand U48980 (N_48980,N_45371,N_46734);
nand U48981 (N_48981,N_47296,N_46922);
or U48982 (N_48982,N_45101,N_46780);
or U48983 (N_48983,N_45039,N_47295);
nand U48984 (N_48984,N_47193,N_45164);
and U48985 (N_48985,N_46164,N_47355);
nand U48986 (N_48986,N_46847,N_46904);
and U48987 (N_48987,N_45214,N_45312);
or U48988 (N_48988,N_46725,N_46866);
nand U48989 (N_48989,N_45011,N_45445);
or U48990 (N_48990,N_47272,N_46953);
nand U48991 (N_48991,N_45830,N_46911);
nor U48992 (N_48992,N_47319,N_46140);
nor U48993 (N_48993,N_45996,N_46354);
nand U48994 (N_48994,N_45674,N_46249);
nand U48995 (N_48995,N_46021,N_46467);
or U48996 (N_48996,N_46330,N_45065);
nor U48997 (N_48997,N_45279,N_47191);
or U48998 (N_48998,N_47481,N_46629);
nand U48999 (N_48999,N_45378,N_46762);
xnor U49000 (N_49000,N_45391,N_46462);
or U49001 (N_49001,N_46490,N_46421);
and U49002 (N_49002,N_45935,N_47261);
or U49003 (N_49003,N_46002,N_47495);
nand U49004 (N_49004,N_45657,N_45237);
xor U49005 (N_49005,N_46665,N_45060);
or U49006 (N_49006,N_46864,N_46761);
nand U49007 (N_49007,N_45948,N_45907);
nor U49008 (N_49008,N_45550,N_46517);
or U49009 (N_49009,N_45677,N_47316);
and U49010 (N_49010,N_46440,N_45794);
xnor U49011 (N_49011,N_45853,N_47407);
nor U49012 (N_49012,N_46912,N_47058);
nand U49013 (N_49013,N_47031,N_45094);
nand U49014 (N_49014,N_45249,N_45247);
xnor U49015 (N_49015,N_47449,N_47271);
or U49016 (N_49016,N_45724,N_46099);
nand U49017 (N_49017,N_47411,N_46239);
and U49018 (N_49018,N_46781,N_45719);
nand U49019 (N_49019,N_46270,N_45849);
nor U49020 (N_49020,N_46800,N_47434);
nor U49021 (N_49021,N_45931,N_45615);
xor U49022 (N_49022,N_45169,N_45212);
nand U49023 (N_49023,N_47000,N_46703);
or U49024 (N_49024,N_45077,N_46316);
nand U49025 (N_49025,N_47206,N_46501);
or U49026 (N_49026,N_46144,N_46146);
xnor U49027 (N_49027,N_46910,N_45056);
and U49028 (N_49028,N_46085,N_47017);
and U49029 (N_49029,N_47446,N_45345);
nor U49030 (N_49030,N_47162,N_45652);
nand U49031 (N_49031,N_45606,N_47027);
xor U49032 (N_49032,N_45118,N_47032);
xor U49033 (N_49033,N_45824,N_47372);
nor U49034 (N_49034,N_46503,N_47011);
xnor U49035 (N_49035,N_46243,N_47042);
xor U49036 (N_49036,N_47247,N_45653);
xnor U49037 (N_49037,N_47263,N_47060);
nor U49038 (N_49038,N_46786,N_46421);
and U49039 (N_49039,N_46139,N_46235);
nand U49040 (N_49040,N_45095,N_47381);
or U49041 (N_49041,N_46334,N_45439);
and U49042 (N_49042,N_45122,N_46534);
nand U49043 (N_49043,N_45314,N_46028);
nor U49044 (N_49044,N_45119,N_46497);
or U49045 (N_49045,N_45950,N_45690);
or U49046 (N_49046,N_47474,N_46753);
or U49047 (N_49047,N_45464,N_47489);
and U49048 (N_49048,N_46583,N_46610);
xor U49049 (N_49049,N_45356,N_47295);
and U49050 (N_49050,N_45828,N_45955);
xnor U49051 (N_49051,N_45627,N_45394);
nor U49052 (N_49052,N_45651,N_47278);
nor U49053 (N_49053,N_46833,N_47045);
nor U49054 (N_49054,N_45446,N_45021);
and U49055 (N_49055,N_45507,N_45033);
nand U49056 (N_49056,N_45740,N_46469);
xor U49057 (N_49057,N_46099,N_47482);
or U49058 (N_49058,N_45286,N_46995);
nor U49059 (N_49059,N_46534,N_46854);
nand U49060 (N_49060,N_46863,N_45142);
and U49061 (N_49061,N_45190,N_45327);
nor U49062 (N_49062,N_45030,N_46572);
or U49063 (N_49063,N_46782,N_47212);
nand U49064 (N_49064,N_47262,N_46751);
nor U49065 (N_49065,N_47420,N_45113);
or U49066 (N_49066,N_45547,N_47491);
xor U49067 (N_49067,N_47160,N_46417);
and U49068 (N_49068,N_46090,N_45705);
nor U49069 (N_49069,N_46417,N_47116);
and U49070 (N_49070,N_46085,N_45150);
or U49071 (N_49071,N_46340,N_46617);
or U49072 (N_49072,N_46391,N_46529);
and U49073 (N_49073,N_46201,N_46312);
and U49074 (N_49074,N_47403,N_45405);
and U49075 (N_49075,N_45741,N_45921);
nand U49076 (N_49076,N_47377,N_45390);
xor U49077 (N_49077,N_45183,N_46255);
or U49078 (N_49078,N_45964,N_46066);
or U49079 (N_49079,N_45187,N_46414);
nor U49080 (N_49080,N_45708,N_45562);
nor U49081 (N_49081,N_47051,N_45074);
nor U49082 (N_49082,N_45398,N_45915);
or U49083 (N_49083,N_45418,N_45622);
nand U49084 (N_49084,N_47455,N_46338);
and U49085 (N_49085,N_47175,N_47114);
nand U49086 (N_49086,N_45873,N_47408);
or U49087 (N_49087,N_46110,N_46324);
and U49088 (N_49088,N_46891,N_45388);
nor U49089 (N_49089,N_46402,N_45412);
and U49090 (N_49090,N_47463,N_47449);
xnor U49091 (N_49091,N_46350,N_45534);
nor U49092 (N_49092,N_45277,N_47380);
or U49093 (N_49093,N_45380,N_46292);
or U49094 (N_49094,N_45523,N_45833);
nand U49095 (N_49095,N_46403,N_45667);
xnor U49096 (N_49096,N_45994,N_45509);
nand U49097 (N_49097,N_45039,N_45066);
xnor U49098 (N_49098,N_47285,N_47099);
nand U49099 (N_49099,N_46893,N_47475);
or U49100 (N_49100,N_47078,N_47134);
xor U49101 (N_49101,N_46473,N_46338);
nor U49102 (N_49102,N_47209,N_45740);
nand U49103 (N_49103,N_47450,N_46794);
nand U49104 (N_49104,N_46067,N_45651);
nor U49105 (N_49105,N_47338,N_46867);
nor U49106 (N_49106,N_45198,N_45045);
nor U49107 (N_49107,N_45516,N_46680);
nor U49108 (N_49108,N_45870,N_45365);
nor U49109 (N_49109,N_46254,N_47312);
or U49110 (N_49110,N_45569,N_46054);
xnor U49111 (N_49111,N_45816,N_45328);
and U49112 (N_49112,N_47288,N_45808);
or U49113 (N_49113,N_45687,N_47216);
xor U49114 (N_49114,N_45086,N_45198);
nor U49115 (N_49115,N_45528,N_45996);
and U49116 (N_49116,N_45115,N_45665);
nor U49117 (N_49117,N_47082,N_46037);
nand U49118 (N_49118,N_47023,N_45845);
nor U49119 (N_49119,N_45297,N_46876);
nand U49120 (N_49120,N_46297,N_45789);
nand U49121 (N_49121,N_46462,N_45059);
xnor U49122 (N_49122,N_45839,N_45655);
and U49123 (N_49123,N_45371,N_46995);
xnor U49124 (N_49124,N_47198,N_45212);
xor U49125 (N_49125,N_47111,N_47253);
and U49126 (N_49126,N_47116,N_45300);
nand U49127 (N_49127,N_46018,N_45616);
xor U49128 (N_49128,N_46760,N_47342);
or U49129 (N_49129,N_45904,N_46697);
and U49130 (N_49130,N_45521,N_45994);
and U49131 (N_49131,N_45821,N_45794);
nand U49132 (N_49132,N_46615,N_45726);
xnor U49133 (N_49133,N_46873,N_45820);
or U49134 (N_49134,N_46950,N_45589);
xor U49135 (N_49135,N_45889,N_46003);
or U49136 (N_49136,N_45573,N_46783);
nand U49137 (N_49137,N_45572,N_46888);
xnor U49138 (N_49138,N_46778,N_46415);
nor U49139 (N_49139,N_45170,N_46776);
or U49140 (N_49140,N_46639,N_45087);
or U49141 (N_49141,N_46121,N_46239);
or U49142 (N_49142,N_45391,N_47149);
nand U49143 (N_49143,N_47311,N_45282);
xor U49144 (N_49144,N_45156,N_46652);
or U49145 (N_49145,N_46290,N_46835);
or U49146 (N_49146,N_45752,N_46462);
or U49147 (N_49147,N_46002,N_45267);
nor U49148 (N_49148,N_45219,N_47106);
nor U49149 (N_49149,N_45862,N_45244);
nand U49150 (N_49150,N_45340,N_47134);
or U49151 (N_49151,N_45472,N_45183);
or U49152 (N_49152,N_47138,N_46466);
xor U49153 (N_49153,N_45769,N_45228);
or U49154 (N_49154,N_46810,N_46325);
nand U49155 (N_49155,N_47396,N_47014);
and U49156 (N_49156,N_45027,N_46279);
nor U49157 (N_49157,N_45586,N_45693);
and U49158 (N_49158,N_45387,N_46745);
xnor U49159 (N_49159,N_46283,N_45391);
nor U49160 (N_49160,N_45756,N_45096);
xor U49161 (N_49161,N_47239,N_45172);
nor U49162 (N_49162,N_46717,N_45145);
and U49163 (N_49163,N_46862,N_47339);
xnor U49164 (N_49164,N_45524,N_45324);
nor U49165 (N_49165,N_45707,N_47226);
nor U49166 (N_49166,N_45657,N_46010);
xnor U49167 (N_49167,N_47342,N_46321);
xor U49168 (N_49168,N_46236,N_45187);
xnor U49169 (N_49169,N_45074,N_46783);
nand U49170 (N_49170,N_46547,N_45920);
or U49171 (N_49171,N_46152,N_45316);
and U49172 (N_49172,N_45784,N_46286);
nor U49173 (N_49173,N_46727,N_46981);
and U49174 (N_49174,N_47351,N_45020);
and U49175 (N_49175,N_46191,N_46478);
and U49176 (N_49176,N_45938,N_46340);
nand U49177 (N_49177,N_45780,N_46396);
nand U49178 (N_49178,N_45929,N_46797);
nor U49179 (N_49179,N_45174,N_46659);
nand U49180 (N_49180,N_47458,N_45893);
xnor U49181 (N_49181,N_46443,N_45517);
and U49182 (N_49182,N_46576,N_45333);
and U49183 (N_49183,N_46068,N_45462);
or U49184 (N_49184,N_46850,N_46331);
or U49185 (N_49185,N_46454,N_47426);
nand U49186 (N_49186,N_45783,N_45290);
or U49187 (N_49187,N_46855,N_45638);
or U49188 (N_49188,N_46821,N_45285);
nand U49189 (N_49189,N_47376,N_47046);
and U49190 (N_49190,N_47182,N_45953);
xnor U49191 (N_49191,N_45631,N_46525);
xor U49192 (N_49192,N_45737,N_45618);
and U49193 (N_49193,N_45714,N_46256);
xor U49194 (N_49194,N_46337,N_46628);
xor U49195 (N_49195,N_45521,N_47468);
or U49196 (N_49196,N_45447,N_46079);
nor U49197 (N_49197,N_46022,N_46421);
nor U49198 (N_49198,N_45769,N_46959);
nand U49199 (N_49199,N_47196,N_46436);
and U49200 (N_49200,N_47181,N_46509);
and U49201 (N_49201,N_47163,N_45478);
nor U49202 (N_49202,N_46083,N_45459);
nor U49203 (N_49203,N_46464,N_46496);
nor U49204 (N_49204,N_45697,N_47443);
and U49205 (N_49205,N_47113,N_45395);
or U49206 (N_49206,N_45523,N_47103);
nor U49207 (N_49207,N_45869,N_46169);
or U49208 (N_49208,N_46049,N_47042);
and U49209 (N_49209,N_46397,N_46314);
nor U49210 (N_49210,N_45250,N_45778);
nor U49211 (N_49211,N_47351,N_47250);
xor U49212 (N_49212,N_45175,N_45923);
nor U49213 (N_49213,N_45420,N_46522);
nor U49214 (N_49214,N_46467,N_46250);
or U49215 (N_49215,N_45905,N_45365);
nor U49216 (N_49216,N_47049,N_45132);
nor U49217 (N_49217,N_46180,N_45972);
xor U49218 (N_49218,N_46842,N_45727);
nor U49219 (N_49219,N_46934,N_47496);
xor U49220 (N_49220,N_45990,N_45322);
and U49221 (N_49221,N_45600,N_45252);
or U49222 (N_49222,N_45445,N_47242);
or U49223 (N_49223,N_46534,N_46334);
nor U49224 (N_49224,N_45744,N_45043);
nand U49225 (N_49225,N_45557,N_47259);
and U49226 (N_49226,N_45307,N_46313);
nand U49227 (N_49227,N_45388,N_47124);
or U49228 (N_49228,N_45002,N_45215);
or U49229 (N_49229,N_46048,N_45574);
xor U49230 (N_49230,N_46169,N_47027);
and U49231 (N_49231,N_45729,N_45596);
nor U49232 (N_49232,N_47451,N_45793);
or U49233 (N_49233,N_46619,N_45734);
or U49234 (N_49234,N_46203,N_45367);
nor U49235 (N_49235,N_45812,N_47459);
nand U49236 (N_49236,N_46553,N_47082);
xnor U49237 (N_49237,N_45950,N_45961);
xnor U49238 (N_49238,N_46014,N_46171);
xnor U49239 (N_49239,N_45152,N_46453);
or U49240 (N_49240,N_47306,N_46005);
and U49241 (N_49241,N_45041,N_45865);
nand U49242 (N_49242,N_47456,N_46983);
and U49243 (N_49243,N_46947,N_46005);
nand U49244 (N_49244,N_47481,N_45895);
xor U49245 (N_49245,N_46890,N_46565);
and U49246 (N_49246,N_47429,N_45878);
nor U49247 (N_49247,N_46195,N_46301);
nor U49248 (N_49248,N_46068,N_45772);
and U49249 (N_49249,N_47159,N_47419);
or U49250 (N_49250,N_46963,N_47176);
or U49251 (N_49251,N_47303,N_46681);
xor U49252 (N_49252,N_45052,N_46358);
nand U49253 (N_49253,N_46053,N_45630);
nor U49254 (N_49254,N_45124,N_46658);
and U49255 (N_49255,N_45597,N_46303);
or U49256 (N_49256,N_45794,N_46557);
nor U49257 (N_49257,N_45517,N_47412);
and U49258 (N_49258,N_45565,N_45443);
xor U49259 (N_49259,N_46662,N_46054);
and U49260 (N_49260,N_45312,N_46255);
nor U49261 (N_49261,N_46427,N_46863);
and U49262 (N_49262,N_45847,N_45392);
nand U49263 (N_49263,N_45086,N_46606);
nor U49264 (N_49264,N_45325,N_47329);
nand U49265 (N_49265,N_47441,N_45155);
xor U49266 (N_49266,N_46905,N_46581);
nand U49267 (N_49267,N_46186,N_46045);
or U49268 (N_49268,N_47457,N_47229);
or U49269 (N_49269,N_45805,N_46446);
and U49270 (N_49270,N_46778,N_45163);
or U49271 (N_49271,N_47188,N_45664);
and U49272 (N_49272,N_45693,N_46762);
or U49273 (N_49273,N_46656,N_45241);
nor U49274 (N_49274,N_45094,N_46702);
xnor U49275 (N_49275,N_46967,N_46209);
nor U49276 (N_49276,N_46751,N_46834);
nand U49277 (N_49277,N_45670,N_47332);
nor U49278 (N_49278,N_47386,N_45337);
or U49279 (N_49279,N_46983,N_46487);
nand U49280 (N_49280,N_46509,N_45444);
or U49281 (N_49281,N_46121,N_47174);
or U49282 (N_49282,N_47173,N_46625);
xor U49283 (N_49283,N_45613,N_46177);
and U49284 (N_49284,N_46351,N_45572);
nand U49285 (N_49285,N_46063,N_46868);
nand U49286 (N_49286,N_45914,N_45150);
xnor U49287 (N_49287,N_46243,N_45057);
xnor U49288 (N_49288,N_46097,N_45751);
nor U49289 (N_49289,N_47338,N_45170);
nand U49290 (N_49290,N_45969,N_46449);
nor U49291 (N_49291,N_45995,N_46629);
and U49292 (N_49292,N_47160,N_45149);
xor U49293 (N_49293,N_46435,N_45622);
nand U49294 (N_49294,N_45258,N_46651);
or U49295 (N_49295,N_47276,N_46063);
xor U49296 (N_49296,N_46966,N_47082);
xnor U49297 (N_49297,N_45694,N_46760);
nand U49298 (N_49298,N_46979,N_46031);
xor U49299 (N_49299,N_45293,N_45368);
or U49300 (N_49300,N_46892,N_46346);
nand U49301 (N_49301,N_45331,N_46652);
nor U49302 (N_49302,N_45153,N_47380);
nand U49303 (N_49303,N_46878,N_45671);
or U49304 (N_49304,N_47283,N_45810);
xnor U49305 (N_49305,N_45456,N_47116);
nand U49306 (N_49306,N_46866,N_47133);
nand U49307 (N_49307,N_46087,N_45221);
xor U49308 (N_49308,N_46657,N_45277);
nand U49309 (N_49309,N_45538,N_46076);
nand U49310 (N_49310,N_47252,N_46364);
nand U49311 (N_49311,N_46636,N_45055);
xor U49312 (N_49312,N_45732,N_45399);
nand U49313 (N_49313,N_47426,N_45432);
or U49314 (N_49314,N_46791,N_46565);
nand U49315 (N_49315,N_46358,N_46204);
nand U49316 (N_49316,N_47041,N_46725);
nand U49317 (N_49317,N_46081,N_46077);
or U49318 (N_49318,N_46759,N_45920);
xnor U49319 (N_49319,N_45700,N_45669);
and U49320 (N_49320,N_45512,N_45391);
xor U49321 (N_49321,N_47173,N_46415);
and U49322 (N_49322,N_45632,N_46947);
xor U49323 (N_49323,N_47226,N_45668);
and U49324 (N_49324,N_46849,N_47194);
nor U49325 (N_49325,N_45571,N_45240);
and U49326 (N_49326,N_45717,N_46857);
nor U49327 (N_49327,N_46328,N_47096);
nor U49328 (N_49328,N_45561,N_46359);
nand U49329 (N_49329,N_45254,N_47004);
xor U49330 (N_49330,N_46286,N_47082);
and U49331 (N_49331,N_47028,N_46503);
and U49332 (N_49332,N_45059,N_47316);
nor U49333 (N_49333,N_45164,N_45543);
or U49334 (N_49334,N_46172,N_45585);
or U49335 (N_49335,N_47342,N_46392);
and U49336 (N_49336,N_46515,N_47430);
and U49337 (N_49337,N_46540,N_46042);
nand U49338 (N_49338,N_46330,N_45217);
and U49339 (N_49339,N_45542,N_46386);
and U49340 (N_49340,N_45332,N_45513);
and U49341 (N_49341,N_47107,N_46587);
nor U49342 (N_49342,N_46322,N_46376);
xnor U49343 (N_49343,N_47285,N_47058);
and U49344 (N_49344,N_45392,N_45084);
nor U49345 (N_49345,N_45020,N_46183);
and U49346 (N_49346,N_45100,N_45668);
xor U49347 (N_49347,N_45075,N_47140);
nor U49348 (N_49348,N_46386,N_47058);
and U49349 (N_49349,N_45327,N_46993);
nand U49350 (N_49350,N_46789,N_45787);
xnor U49351 (N_49351,N_45144,N_47402);
nor U49352 (N_49352,N_45173,N_47393);
nand U49353 (N_49353,N_47373,N_45465);
xor U49354 (N_49354,N_45238,N_46267);
and U49355 (N_49355,N_47450,N_45211);
or U49356 (N_49356,N_47346,N_46767);
nor U49357 (N_49357,N_45605,N_45108);
and U49358 (N_49358,N_46128,N_45414);
and U49359 (N_49359,N_46266,N_45631);
and U49360 (N_49360,N_45314,N_45277);
or U49361 (N_49361,N_46566,N_46202);
or U49362 (N_49362,N_45563,N_46046);
xnor U49363 (N_49363,N_47398,N_46139);
nor U49364 (N_49364,N_46356,N_47189);
or U49365 (N_49365,N_46399,N_46125);
nand U49366 (N_49366,N_47024,N_45382);
xor U49367 (N_49367,N_46183,N_46013);
or U49368 (N_49368,N_45729,N_45733);
nor U49369 (N_49369,N_46894,N_46957);
xnor U49370 (N_49370,N_46645,N_46623);
nand U49371 (N_49371,N_47324,N_45758);
xor U49372 (N_49372,N_46890,N_46356);
nand U49373 (N_49373,N_45288,N_46100);
xnor U49374 (N_49374,N_45670,N_47041);
and U49375 (N_49375,N_45304,N_45337);
or U49376 (N_49376,N_45349,N_47069);
nor U49377 (N_49377,N_46147,N_46157);
and U49378 (N_49378,N_45906,N_46172);
xnor U49379 (N_49379,N_46316,N_46500);
xnor U49380 (N_49380,N_46501,N_45876);
nand U49381 (N_49381,N_47307,N_47465);
nor U49382 (N_49382,N_45070,N_46264);
nand U49383 (N_49383,N_46057,N_46712);
xor U49384 (N_49384,N_46432,N_45782);
and U49385 (N_49385,N_45179,N_46500);
xnor U49386 (N_49386,N_45223,N_45317);
nand U49387 (N_49387,N_47020,N_46889);
nand U49388 (N_49388,N_46270,N_46945);
and U49389 (N_49389,N_46039,N_45831);
or U49390 (N_49390,N_46679,N_46825);
or U49391 (N_49391,N_45853,N_47355);
and U49392 (N_49392,N_46905,N_46862);
and U49393 (N_49393,N_45700,N_45987);
nor U49394 (N_49394,N_45011,N_46320);
nor U49395 (N_49395,N_46186,N_47035);
xnor U49396 (N_49396,N_46479,N_45908);
nor U49397 (N_49397,N_45269,N_45655);
or U49398 (N_49398,N_47454,N_46364);
or U49399 (N_49399,N_47374,N_45969);
and U49400 (N_49400,N_45267,N_46488);
xor U49401 (N_49401,N_46122,N_45591);
nand U49402 (N_49402,N_45618,N_47130);
or U49403 (N_49403,N_47422,N_46480);
or U49404 (N_49404,N_45680,N_45259);
or U49405 (N_49405,N_46177,N_46563);
and U49406 (N_49406,N_45636,N_47187);
xnor U49407 (N_49407,N_45005,N_46808);
or U49408 (N_49408,N_46721,N_46834);
nor U49409 (N_49409,N_45559,N_45456);
xnor U49410 (N_49410,N_45242,N_46852);
nor U49411 (N_49411,N_47226,N_47357);
xnor U49412 (N_49412,N_45472,N_47195);
or U49413 (N_49413,N_45618,N_45511);
nand U49414 (N_49414,N_45329,N_47126);
xor U49415 (N_49415,N_47155,N_45858);
or U49416 (N_49416,N_45097,N_45388);
or U49417 (N_49417,N_45408,N_45644);
nor U49418 (N_49418,N_45091,N_47244);
xnor U49419 (N_49419,N_47418,N_47090);
xor U49420 (N_49420,N_45315,N_45373);
or U49421 (N_49421,N_46365,N_47052);
xnor U49422 (N_49422,N_45559,N_47482);
or U49423 (N_49423,N_45681,N_46815);
nor U49424 (N_49424,N_45702,N_47244);
nand U49425 (N_49425,N_46299,N_45352);
nand U49426 (N_49426,N_45978,N_47240);
nor U49427 (N_49427,N_45766,N_45189);
or U49428 (N_49428,N_46735,N_46430);
or U49429 (N_49429,N_46847,N_46723);
nor U49430 (N_49430,N_45382,N_45561);
nor U49431 (N_49431,N_45933,N_45627);
or U49432 (N_49432,N_46163,N_46959);
nand U49433 (N_49433,N_47328,N_47033);
or U49434 (N_49434,N_46636,N_45640);
or U49435 (N_49435,N_45051,N_47477);
or U49436 (N_49436,N_45480,N_47357);
nor U49437 (N_49437,N_46897,N_45677);
nand U49438 (N_49438,N_45401,N_46075);
nor U49439 (N_49439,N_46531,N_45580);
and U49440 (N_49440,N_45136,N_46489);
nor U49441 (N_49441,N_46221,N_47105);
nor U49442 (N_49442,N_45847,N_45741);
and U49443 (N_49443,N_45459,N_47128);
xnor U49444 (N_49444,N_45958,N_46817);
or U49445 (N_49445,N_47383,N_46472);
nand U49446 (N_49446,N_46945,N_45630);
nor U49447 (N_49447,N_45305,N_46406);
nand U49448 (N_49448,N_47390,N_46328);
or U49449 (N_49449,N_46255,N_47122);
and U49450 (N_49450,N_45130,N_45747);
nor U49451 (N_49451,N_46246,N_47333);
nor U49452 (N_49452,N_45207,N_46447);
nand U49453 (N_49453,N_45084,N_46935);
xnor U49454 (N_49454,N_45502,N_45292);
and U49455 (N_49455,N_46816,N_46610);
or U49456 (N_49456,N_46043,N_45372);
nor U49457 (N_49457,N_46944,N_46065);
and U49458 (N_49458,N_45486,N_46668);
nor U49459 (N_49459,N_46138,N_45518);
and U49460 (N_49460,N_45340,N_45170);
nor U49461 (N_49461,N_46296,N_45670);
nor U49462 (N_49462,N_46494,N_46665);
and U49463 (N_49463,N_45822,N_46937);
and U49464 (N_49464,N_46532,N_46886);
nor U49465 (N_49465,N_45686,N_46971);
and U49466 (N_49466,N_45545,N_47175);
and U49467 (N_49467,N_45421,N_46757);
and U49468 (N_49468,N_45377,N_47006);
nand U49469 (N_49469,N_45003,N_46700);
nor U49470 (N_49470,N_46619,N_45336);
xnor U49471 (N_49471,N_46633,N_45163);
or U49472 (N_49472,N_47086,N_46313);
or U49473 (N_49473,N_45392,N_45137);
nor U49474 (N_49474,N_45799,N_45226);
and U49475 (N_49475,N_45774,N_46769);
xnor U49476 (N_49476,N_45410,N_47168);
xnor U49477 (N_49477,N_45606,N_45513);
or U49478 (N_49478,N_45260,N_46191);
and U49479 (N_49479,N_47441,N_46792);
or U49480 (N_49480,N_46736,N_45189);
nand U49481 (N_49481,N_45743,N_46846);
nand U49482 (N_49482,N_47038,N_46045);
nor U49483 (N_49483,N_46314,N_46937);
nand U49484 (N_49484,N_45331,N_46976);
xnor U49485 (N_49485,N_46214,N_45328);
xnor U49486 (N_49486,N_46823,N_45156);
nor U49487 (N_49487,N_46170,N_46458);
xor U49488 (N_49488,N_46289,N_47284);
nor U49489 (N_49489,N_46988,N_46684);
xnor U49490 (N_49490,N_46103,N_46243);
nor U49491 (N_49491,N_45873,N_46176);
xor U49492 (N_49492,N_46895,N_45913);
xnor U49493 (N_49493,N_46474,N_47145);
xor U49494 (N_49494,N_46541,N_47004);
nor U49495 (N_49495,N_46310,N_47385);
xor U49496 (N_49496,N_46820,N_47241);
xnor U49497 (N_49497,N_45628,N_46970);
and U49498 (N_49498,N_47418,N_45092);
and U49499 (N_49499,N_46647,N_46043);
and U49500 (N_49500,N_46628,N_47124);
nand U49501 (N_49501,N_45357,N_45061);
or U49502 (N_49502,N_47064,N_47093);
nor U49503 (N_49503,N_45392,N_45329);
xor U49504 (N_49504,N_47496,N_47164);
nand U49505 (N_49505,N_45263,N_46698);
or U49506 (N_49506,N_45541,N_46789);
nand U49507 (N_49507,N_47446,N_45320);
xor U49508 (N_49508,N_45535,N_47079);
or U49509 (N_49509,N_46083,N_46261);
xnor U49510 (N_49510,N_47201,N_46778);
nor U49511 (N_49511,N_47474,N_46704);
nor U49512 (N_49512,N_46065,N_45506);
or U49513 (N_49513,N_45319,N_45239);
nor U49514 (N_49514,N_47459,N_47491);
or U49515 (N_49515,N_46204,N_46379);
xor U49516 (N_49516,N_47152,N_46404);
xnor U49517 (N_49517,N_46421,N_46980);
xor U49518 (N_49518,N_46001,N_45398);
xor U49519 (N_49519,N_47426,N_45845);
nand U49520 (N_49520,N_46553,N_47312);
nand U49521 (N_49521,N_45084,N_46774);
or U49522 (N_49522,N_46883,N_46718);
and U49523 (N_49523,N_45380,N_46280);
or U49524 (N_49524,N_46497,N_46568);
and U49525 (N_49525,N_46619,N_47133);
xor U49526 (N_49526,N_45522,N_45986);
nor U49527 (N_49527,N_45679,N_46134);
or U49528 (N_49528,N_45265,N_45982);
or U49529 (N_49529,N_46746,N_45681);
nor U49530 (N_49530,N_45196,N_46598);
and U49531 (N_49531,N_47481,N_45460);
nor U49532 (N_49532,N_45867,N_46934);
nor U49533 (N_49533,N_45504,N_47013);
nand U49534 (N_49534,N_47338,N_45777);
nor U49535 (N_49535,N_46815,N_45294);
or U49536 (N_49536,N_46252,N_46901);
xnor U49537 (N_49537,N_45032,N_46124);
nor U49538 (N_49538,N_45038,N_46275);
xor U49539 (N_49539,N_46939,N_46395);
nor U49540 (N_49540,N_45105,N_46240);
xor U49541 (N_49541,N_46674,N_47294);
or U49542 (N_49542,N_47162,N_45163);
and U49543 (N_49543,N_47487,N_46352);
or U49544 (N_49544,N_45599,N_47302);
xor U49545 (N_49545,N_45516,N_45431);
and U49546 (N_49546,N_46910,N_46912);
nor U49547 (N_49547,N_45919,N_47339);
nor U49548 (N_49548,N_46146,N_45534);
nand U49549 (N_49549,N_45056,N_45675);
and U49550 (N_49550,N_46602,N_45133);
nor U49551 (N_49551,N_45012,N_46613);
nand U49552 (N_49552,N_45765,N_46714);
and U49553 (N_49553,N_45337,N_47262);
and U49554 (N_49554,N_45538,N_45461);
and U49555 (N_49555,N_45236,N_46710);
nand U49556 (N_49556,N_45339,N_46536);
nor U49557 (N_49557,N_46629,N_46566);
nand U49558 (N_49558,N_45451,N_45266);
xnor U49559 (N_49559,N_45391,N_46019);
or U49560 (N_49560,N_45172,N_46656);
nand U49561 (N_49561,N_45606,N_47288);
xor U49562 (N_49562,N_45842,N_45380);
nor U49563 (N_49563,N_45424,N_46258);
nand U49564 (N_49564,N_47091,N_46627);
and U49565 (N_49565,N_47385,N_45509);
and U49566 (N_49566,N_45200,N_45173);
or U49567 (N_49567,N_46311,N_45293);
nand U49568 (N_49568,N_45596,N_47407);
nand U49569 (N_49569,N_46133,N_45154);
or U49570 (N_49570,N_46761,N_46144);
nand U49571 (N_49571,N_45239,N_45010);
xor U49572 (N_49572,N_46904,N_45051);
xor U49573 (N_49573,N_47209,N_45441);
or U49574 (N_49574,N_47004,N_46385);
xnor U49575 (N_49575,N_46691,N_46670);
nand U49576 (N_49576,N_45598,N_45173);
or U49577 (N_49577,N_46581,N_47273);
nand U49578 (N_49578,N_46479,N_45460);
and U49579 (N_49579,N_47072,N_45479);
nor U49580 (N_49580,N_46723,N_46341);
and U49581 (N_49581,N_45636,N_46416);
or U49582 (N_49582,N_47326,N_46222);
and U49583 (N_49583,N_45759,N_47466);
nor U49584 (N_49584,N_45618,N_47167);
nor U49585 (N_49585,N_47202,N_46508);
or U49586 (N_49586,N_47132,N_46792);
xor U49587 (N_49587,N_45853,N_46406);
or U49588 (N_49588,N_45641,N_45639);
or U49589 (N_49589,N_47389,N_45009);
nor U49590 (N_49590,N_46058,N_45132);
nand U49591 (N_49591,N_46982,N_46659);
and U49592 (N_49592,N_47040,N_45078);
xnor U49593 (N_49593,N_46172,N_45100);
xnor U49594 (N_49594,N_46523,N_45404);
xor U49595 (N_49595,N_45779,N_45019);
xor U49596 (N_49596,N_46565,N_47022);
and U49597 (N_49597,N_46084,N_45483);
xor U49598 (N_49598,N_47020,N_46604);
and U49599 (N_49599,N_46541,N_46672);
nor U49600 (N_49600,N_47450,N_47072);
nand U49601 (N_49601,N_47227,N_45802);
nand U49602 (N_49602,N_45851,N_46533);
or U49603 (N_49603,N_45566,N_46675);
or U49604 (N_49604,N_46730,N_46182);
nand U49605 (N_49605,N_46880,N_47346);
and U49606 (N_49606,N_46424,N_45994);
xor U49607 (N_49607,N_46139,N_47430);
nor U49608 (N_49608,N_45800,N_47422);
nor U49609 (N_49609,N_45925,N_46903);
and U49610 (N_49610,N_47352,N_45461);
nand U49611 (N_49611,N_46547,N_45309);
nand U49612 (N_49612,N_45314,N_46293);
or U49613 (N_49613,N_45445,N_45821);
xnor U49614 (N_49614,N_45608,N_46279);
nor U49615 (N_49615,N_47373,N_47324);
nor U49616 (N_49616,N_45012,N_45899);
nand U49617 (N_49617,N_46025,N_46080);
nor U49618 (N_49618,N_46938,N_45408);
or U49619 (N_49619,N_46414,N_46801);
nor U49620 (N_49620,N_45089,N_45680);
and U49621 (N_49621,N_45595,N_46976);
or U49622 (N_49622,N_46182,N_46610);
and U49623 (N_49623,N_46736,N_47155);
or U49624 (N_49624,N_46726,N_46238);
and U49625 (N_49625,N_46428,N_45572);
xor U49626 (N_49626,N_47376,N_46654);
nor U49627 (N_49627,N_47177,N_46035);
nor U49628 (N_49628,N_45852,N_46704);
xor U49629 (N_49629,N_46046,N_45687);
nand U49630 (N_49630,N_46017,N_46498);
and U49631 (N_49631,N_46989,N_46427);
and U49632 (N_49632,N_47058,N_45432);
xnor U49633 (N_49633,N_46010,N_47336);
xnor U49634 (N_49634,N_46730,N_46376);
or U49635 (N_49635,N_46831,N_46015);
or U49636 (N_49636,N_45449,N_45508);
nand U49637 (N_49637,N_45971,N_47174);
and U49638 (N_49638,N_46008,N_46734);
nor U49639 (N_49639,N_45197,N_46035);
and U49640 (N_49640,N_46608,N_46530);
nor U49641 (N_49641,N_45424,N_45747);
nand U49642 (N_49642,N_45759,N_46466);
nand U49643 (N_49643,N_46069,N_46182);
xnor U49644 (N_49644,N_46238,N_45734);
and U49645 (N_49645,N_47285,N_46025);
and U49646 (N_49646,N_45565,N_46476);
or U49647 (N_49647,N_45563,N_45030);
nand U49648 (N_49648,N_45110,N_47492);
nand U49649 (N_49649,N_45998,N_45132);
or U49650 (N_49650,N_46815,N_46863);
nor U49651 (N_49651,N_45861,N_46564);
nand U49652 (N_49652,N_47126,N_45742);
nand U49653 (N_49653,N_45917,N_47077);
xor U49654 (N_49654,N_45875,N_45869);
and U49655 (N_49655,N_47206,N_46125);
nand U49656 (N_49656,N_47062,N_46172);
xnor U49657 (N_49657,N_45819,N_45692);
nor U49658 (N_49658,N_47394,N_46491);
and U49659 (N_49659,N_46789,N_47115);
nor U49660 (N_49660,N_46946,N_47277);
nor U49661 (N_49661,N_45587,N_45307);
nand U49662 (N_49662,N_45140,N_45210);
or U49663 (N_49663,N_46245,N_46770);
and U49664 (N_49664,N_45221,N_46968);
nor U49665 (N_49665,N_47069,N_46740);
xnor U49666 (N_49666,N_45866,N_45766);
and U49667 (N_49667,N_45231,N_47449);
nor U49668 (N_49668,N_46034,N_46697);
nand U49669 (N_49669,N_46868,N_46869);
and U49670 (N_49670,N_46144,N_46603);
or U49671 (N_49671,N_45886,N_45161);
xor U49672 (N_49672,N_45925,N_46926);
xnor U49673 (N_49673,N_47377,N_45914);
and U49674 (N_49674,N_45506,N_46334);
xor U49675 (N_49675,N_47426,N_47128);
or U49676 (N_49676,N_45387,N_45731);
xnor U49677 (N_49677,N_46371,N_46877);
nand U49678 (N_49678,N_47203,N_45727);
nand U49679 (N_49679,N_46023,N_47430);
or U49680 (N_49680,N_45878,N_45024);
or U49681 (N_49681,N_46314,N_46725);
nor U49682 (N_49682,N_46875,N_46091);
xor U49683 (N_49683,N_45717,N_47244);
nand U49684 (N_49684,N_45482,N_46767);
nor U49685 (N_49685,N_46736,N_47386);
xnor U49686 (N_49686,N_47024,N_45246);
and U49687 (N_49687,N_45124,N_46628);
xor U49688 (N_49688,N_46927,N_46017);
or U49689 (N_49689,N_45800,N_45702);
nand U49690 (N_49690,N_45065,N_46423);
and U49691 (N_49691,N_45505,N_47478);
and U49692 (N_49692,N_46607,N_46532);
xor U49693 (N_49693,N_45014,N_47008);
and U49694 (N_49694,N_47294,N_45868);
nand U49695 (N_49695,N_46558,N_45973);
nor U49696 (N_49696,N_47104,N_45825);
nand U49697 (N_49697,N_45546,N_45544);
and U49698 (N_49698,N_45579,N_46913);
nand U49699 (N_49699,N_45447,N_46086);
nor U49700 (N_49700,N_45131,N_45179);
xor U49701 (N_49701,N_47334,N_47152);
and U49702 (N_49702,N_46748,N_45278);
and U49703 (N_49703,N_45406,N_45798);
nor U49704 (N_49704,N_47424,N_47129);
nor U49705 (N_49705,N_46753,N_46022);
nand U49706 (N_49706,N_46751,N_46780);
nand U49707 (N_49707,N_45220,N_46551);
or U49708 (N_49708,N_45658,N_45987);
and U49709 (N_49709,N_47208,N_47111);
or U49710 (N_49710,N_45383,N_46314);
nand U49711 (N_49711,N_45858,N_45801);
nand U49712 (N_49712,N_45905,N_46250);
and U49713 (N_49713,N_46952,N_45525);
nor U49714 (N_49714,N_46502,N_46429);
nor U49715 (N_49715,N_46387,N_46054);
nor U49716 (N_49716,N_45359,N_45658);
and U49717 (N_49717,N_45033,N_46951);
or U49718 (N_49718,N_45707,N_47439);
xnor U49719 (N_49719,N_47020,N_45563);
or U49720 (N_49720,N_46252,N_47060);
or U49721 (N_49721,N_45629,N_47452);
nand U49722 (N_49722,N_46228,N_46655);
nand U49723 (N_49723,N_46891,N_46246);
or U49724 (N_49724,N_46838,N_46577);
nor U49725 (N_49725,N_47118,N_46819);
and U49726 (N_49726,N_46126,N_46528);
or U49727 (N_49727,N_45127,N_46284);
xor U49728 (N_49728,N_47073,N_45709);
xor U49729 (N_49729,N_47114,N_47019);
nand U49730 (N_49730,N_47269,N_45176);
xor U49731 (N_49731,N_45231,N_46103);
xor U49732 (N_49732,N_46288,N_45158);
nor U49733 (N_49733,N_47170,N_47205);
and U49734 (N_49734,N_45718,N_45136);
or U49735 (N_49735,N_47167,N_46234);
nand U49736 (N_49736,N_46854,N_47356);
and U49737 (N_49737,N_46286,N_45824);
nand U49738 (N_49738,N_46846,N_47385);
or U49739 (N_49739,N_46321,N_46541);
and U49740 (N_49740,N_47367,N_46855);
nor U49741 (N_49741,N_46266,N_45424);
nor U49742 (N_49742,N_45620,N_46761);
and U49743 (N_49743,N_45885,N_45495);
nor U49744 (N_49744,N_45593,N_46339);
and U49745 (N_49745,N_47358,N_45147);
nand U49746 (N_49746,N_46175,N_45042);
nor U49747 (N_49747,N_47265,N_46247);
nor U49748 (N_49748,N_47458,N_45358);
nand U49749 (N_49749,N_46155,N_46753);
xnor U49750 (N_49750,N_46650,N_45478);
nor U49751 (N_49751,N_47028,N_46285);
nor U49752 (N_49752,N_45729,N_45747);
nand U49753 (N_49753,N_45489,N_46207);
nor U49754 (N_49754,N_46517,N_47234);
nor U49755 (N_49755,N_46308,N_45266);
or U49756 (N_49756,N_47468,N_46437);
and U49757 (N_49757,N_45579,N_46257);
or U49758 (N_49758,N_45481,N_46690);
or U49759 (N_49759,N_45103,N_47485);
nor U49760 (N_49760,N_46664,N_46180);
xor U49761 (N_49761,N_45031,N_46759);
or U49762 (N_49762,N_45693,N_45675);
xnor U49763 (N_49763,N_45340,N_45477);
or U49764 (N_49764,N_47399,N_46744);
nor U49765 (N_49765,N_46591,N_47201);
nor U49766 (N_49766,N_45479,N_45892);
nor U49767 (N_49767,N_46608,N_45983);
xor U49768 (N_49768,N_47087,N_47486);
nor U49769 (N_49769,N_46134,N_45740);
xnor U49770 (N_49770,N_46698,N_46254);
nand U49771 (N_49771,N_46243,N_45848);
nor U49772 (N_49772,N_45528,N_45050);
nor U49773 (N_49773,N_46197,N_46081);
xnor U49774 (N_49774,N_45567,N_45998);
or U49775 (N_49775,N_45514,N_46276);
xor U49776 (N_49776,N_45286,N_45255);
xor U49777 (N_49777,N_45510,N_46313);
nor U49778 (N_49778,N_46306,N_46336);
or U49779 (N_49779,N_45587,N_47420);
nand U49780 (N_49780,N_47041,N_45550);
nor U49781 (N_49781,N_47223,N_45782);
and U49782 (N_49782,N_46739,N_46707);
nor U49783 (N_49783,N_46768,N_45127);
nand U49784 (N_49784,N_46253,N_45000);
and U49785 (N_49785,N_45262,N_45333);
or U49786 (N_49786,N_46540,N_46810);
nand U49787 (N_49787,N_45403,N_46807);
xnor U49788 (N_49788,N_46546,N_45969);
or U49789 (N_49789,N_45797,N_46981);
or U49790 (N_49790,N_45174,N_45525);
nor U49791 (N_49791,N_45726,N_45589);
and U49792 (N_49792,N_46721,N_46070);
xor U49793 (N_49793,N_46122,N_47460);
or U49794 (N_49794,N_46856,N_45136);
and U49795 (N_49795,N_46766,N_45631);
xnor U49796 (N_49796,N_45815,N_46666);
and U49797 (N_49797,N_45743,N_46661);
xor U49798 (N_49798,N_47398,N_46949);
and U49799 (N_49799,N_46214,N_45842);
or U49800 (N_49800,N_47380,N_45422);
xnor U49801 (N_49801,N_46779,N_45976);
xor U49802 (N_49802,N_45731,N_46048);
nand U49803 (N_49803,N_46807,N_46086);
nor U49804 (N_49804,N_45018,N_45825);
nand U49805 (N_49805,N_46804,N_46286);
and U49806 (N_49806,N_45894,N_46050);
and U49807 (N_49807,N_45187,N_45470);
nor U49808 (N_49808,N_47001,N_46927);
xor U49809 (N_49809,N_45555,N_45557);
and U49810 (N_49810,N_47066,N_47464);
xor U49811 (N_49811,N_46633,N_45783);
nor U49812 (N_49812,N_47099,N_46837);
nor U49813 (N_49813,N_45393,N_47316);
and U49814 (N_49814,N_45005,N_45974);
xor U49815 (N_49815,N_46330,N_45290);
nor U49816 (N_49816,N_45361,N_45238);
nor U49817 (N_49817,N_46551,N_45952);
nor U49818 (N_49818,N_45230,N_46908);
xor U49819 (N_49819,N_46453,N_45084);
xnor U49820 (N_49820,N_45142,N_47000);
nand U49821 (N_49821,N_46329,N_46075);
or U49822 (N_49822,N_47123,N_46795);
xnor U49823 (N_49823,N_46506,N_45954);
nor U49824 (N_49824,N_46951,N_46856);
or U49825 (N_49825,N_46430,N_46181);
nor U49826 (N_49826,N_45999,N_46882);
xnor U49827 (N_49827,N_46405,N_45517);
xor U49828 (N_49828,N_47118,N_46125);
xnor U49829 (N_49829,N_45237,N_46427);
nand U49830 (N_49830,N_46754,N_47310);
nand U49831 (N_49831,N_45011,N_47138);
or U49832 (N_49832,N_46706,N_46848);
and U49833 (N_49833,N_45694,N_45709);
nor U49834 (N_49834,N_46768,N_45973);
nor U49835 (N_49835,N_45718,N_46492);
and U49836 (N_49836,N_46875,N_45182);
nand U49837 (N_49837,N_47416,N_45402);
or U49838 (N_49838,N_46702,N_45754);
and U49839 (N_49839,N_46135,N_47184);
or U49840 (N_49840,N_45918,N_45146);
nor U49841 (N_49841,N_45040,N_45679);
nand U49842 (N_49842,N_46054,N_45156);
xnor U49843 (N_49843,N_45474,N_46503);
or U49844 (N_49844,N_45411,N_47021);
nand U49845 (N_49845,N_47007,N_45554);
xnor U49846 (N_49846,N_46873,N_47059);
nand U49847 (N_49847,N_46630,N_46534);
or U49848 (N_49848,N_46165,N_45915);
and U49849 (N_49849,N_46837,N_45853);
xor U49850 (N_49850,N_45265,N_45878);
xor U49851 (N_49851,N_47248,N_46230);
nand U49852 (N_49852,N_46628,N_45016);
and U49853 (N_49853,N_46741,N_46772);
xnor U49854 (N_49854,N_46560,N_45104);
and U49855 (N_49855,N_45474,N_45512);
xor U49856 (N_49856,N_46502,N_45144);
nand U49857 (N_49857,N_47180,N_46084);
nor U49858 (N_49858,N_46388,N_46293);
and U49859 (N_49859,N_47268,N_46183);
or U49860 (N_49860,N_46429,N_46484);
nand U49861 (N_49861,N_46105,N_45245);
nand U49862 (N_49862,N_47443,N_46313);
and U49863 (N_49863,N_45937,N_47013);
nor U49864 (N_49864,N_45979,N_46955);
nor U49865 (N_49865,N_47476,N_45913);
and U49866 (N_49866,N_46115,N_45994);
or U49867 (N_49867,N_46050,N_45304);
nor U49868 (N_49868,N_45453,N_46988);
nor U49869 (N_49869,N_47011,N_47149);
and U49870 (N_49870,N_45058,N_45220);
xor U49871 (N_49871,N_46696,N_46584);
xor U49872 (N_49872,N_45144,N_47236);
and U49873 (N_49873,N_45608,N_46903);
or U49874 (N_49874,N_45568,N_46799);
and U49875 (N_49875,N_45615,N_45417);
nand U49876 (N_49876,N_46248,N_46234);
nand U49877 (N_49877,N_46636,N_46742);
nor U49878 (N_49878,N_45906,N_45865);
and U49879 (N_49879,N_46243,N_46156);
and U49880 (N_49880,N_46077,N_46477);
nor U49881 (N_49881,N_46964,N_45372);
or U49882 (N_49882,N_46174,N_47313);
nor U49883 (N_49883,N_46251,N_46310);
nand U49884 (N_49884,N_46217,N_46361);
xor U49885 (N_49885,N_45180,N_46177);
nor U49886 (N_49886,N_47489,N_46957);
and U49887 (N_49887,N_46903,N_45596);
nor U49888 (N_49888,N_45484,N_47375);
nand U49889 (N_49889,N_45788,N_46796);
nand U49890 (N_49890,N_46083,N_45859);
or U49891 (N_49891,N_46321,N_45085);
or U49892 (N_49892,N_46278,N_47361);
or U49893 (N_49893,N_45329,N_46977);
nor U49894 (N_49894,N_46079,N_47431);
nor U49895 (N_49895,N_46114,N_46594);
or U49896 (N_49896,N_45907,N_46838);
or U49897 (N_49897,N_46253,N_47409);
nand U49898 (N_49898,N_46843,N_46928);
or U49899 (N_49899,N_45830,N_46270);
nand U49900 (N_49900,N_46790,N_45220);
xnor U49901 (N_49901,N_46496,N_45589);
nor U49902 (N_49902,N_46968,N_47310);
nand U49903 (N_49903,N_45151,N_45661);
and U49904 (N_49904,N_45402,N_46593);
xor U49905 (N_49905,N_47056,N_45284);
nor U49906 (N_49906,N_46088,N_45858);
xor U49907 (N_49907,N_47019,N_46671);
and U49908 (N_49908,N_46470,N_46185);
nand U49909 (N_49909,N_46237,N_46908);
or U49910 (N_49910,N_46785,N_47341);
nor U49911 (N_49911,N_47234,N_47198);
or U49912 (N_49912,N_46046,N_45655);
xnor U49913 (N_49913,N_45901,N_46523);
and U49914 (N_49914,N_46644,N_46339);
and U49915 (N_49915,N_45933,N_46049);
and U49916 (N_49916,N_47254,N_45783);
nor U49917 (N_49917,N_46327,N_45725);
or U49918 (N_49918,N_46094,N_47319);
nor U49919 (N_49919,N_45409,N_46770);
nand U49920 (N_49920,N_45245,N_46652);
nand U49921 (N_49921,N_45572,N_47023);
xnor U49922 (N_49922,N_45779,N_45677);
and U49923 (N_49923,N_45290,N_45210);
and U49924 (N_49924,N_45841,N_45101);
nor U49925 (N_49925,N_45006,N_45827);
xnor U49926 (N_49926,N_45949,N_45668);
or U49927 (N_49927,N_45397,N_47010);
nor U49928 (N_49928,N_46656,N_47220);
or U49929 (N_49929,N_46963,N_45358);
nor U49930 (N_49930,N_46138,N_45746);
nand U49931 (N_49931,N_46229,N_46813);
and U49932 (N_49932,N_45238,N_46894);
nor U49933 (N_49933,N_45501,N_46643);
nand U49934 (N_49934,N_46688,N_45553);
xnor U49935 (N_49935,N_45945,N_45879);
or U49936 (N_49936,N_45475,N_45665);
xnor U49937 (N_49937,N_46752,N_45885);
nand U49938 (N_49938,N_45384,N_45451);
nor U49939 (N_49939,N_45355,N_45256);
xnor U49940 (N_49940,N_46988,N_46839);
or U49941 (N_49941,N_45966,N_46991);
or U49942 (N_49942,N_47212,N_45267);
xor U49943 (N_49943,N_45893,N_47403);
nor U49944 (N_49944,N_45577,N_46143);
nor U49945 (N_49945,N_46505,N_45249);
nor U49946 (N_49946,N_47035,N_45165);
xor U49947 (N_49947,N_46740,N_45197);
or U49948 (N_49948,N_45842,N_46723);
or U49949 (N_49949,N_45995,N_45759);
and U49950 (N_49950,N_45027,N_46284);
xnor U49951 (N_49951,N_46858,N_46941);
nor U49952 (N_49952,N_46078,N_45350);
and U49953 (N_49953,N_45351,N_45559);
nand U49954 (N_49954,N_47436,N_46813);
nor U49955 (N_49955,N_45779,N_47097);
nand U49956 (N_49956,N_45261,N_46405);
nor U49957 (N_49957,N_47332,N_47495);
nor U49958 (N_49958,N_46010,N_45723);
or U49959 (N_49959,N_45160,N_46706);
or U49960 (N_49960,N_45126,N_46618);
xor U49961 (N_49961,N_47055,N_45370);
or U49962 (N_49962,N_45716,N_46200);
nand U49963 (N_49963,N_46167,N_47027);
xnor U49964 (N_49964,N_47214,N_46025);
or U49965 (N_49965,N_46094,N_45876);
and U49966 (N_49966,N_46155,N_46355);
and U49967 (N_49967,N_46409,N_45212);
xnor U49968 (N_49968,N_46606,N_45616);
and U49969 (N_49969,N_46527,N_47211);
nor U49970 (N_49970,N_45127,N_46660);
xor U49971 (N_49971,N_47150,N_46716);
nor U49972 (N_49972,N_45962,N_45202);
and U49973 (N_49973,N_47474,N_46933);
and U49974 (N_49974,N_46372,N_45856);
nand U49975 (N_49975,N_46369,N_46198);
nor U49976 (N_49976,N_46477,N_45707);
and U49977 (N_49977,N_45050,N_46589);
nand U49978 (N_49978,N_45675,N_46248);
and U49979 (N_49979,N_45159,N_45702);
and U49980 (N_49980,N_46793,N_46262);
nor U49981 (N_49981,N_45231,N_45036);
xor U49982 (N_49982,N_47142,N_45541);
or U49983 (N_49983,N_46264,N_46151);
nand U49984 (N_49984,N_46617,N_47476);
nand U49985 (N_49985,N_45077,N_45116);
nand U49986 (N_49986,N_45200,N_45198);
nor U49987 (N_49987,N_45228,N_46570);
nand U49988 (N_49988,N_46799,N_46639);
nor U49989 (N_49989,N_47200,N_45239);
xor U49990 (N_49990,N_45915,N_45187);
or U49991 (N_49991,N_46114,N_45338);
nand U49992 (N_49992,N_46360,N_46029);
and U49993 (N_49993,N_46810,N_46524);
nor U49994 (N_49994,N_47494,N_47344);
or U49995 (N_49995,N_46376,N_45876);
and U49996 (N_49996,N_45109,N_47145);
nand U49997 (N_49997,N_45648,N_45929);
or U49998 (N_49998,N_46583,N_45054);
nand U49999 (N_49999,N_45021,N_47259);
or UO_0 (O_0,N_47580,N_49371);
nand UO_1 (O_1,N_49880,N_49320);
nor UO_2 (O_2,N_47854,N_49216);
or UO_3 (O_3,N_49489,N_49501);
or UO_4 (O_4,N_48805,N_49256);
and UO_5 (O_5,N_49364,N_49615);
nand UO_6 (O_6,N_48110,N_48327);
nor UO_7 (O_7,N_49473,N_47723);
nor UO_8 (O_8,N_48982,N_48939);
or UO_9 (O_9,N_48920,N_49813);
nor UO_10 (O_10,N_49893,N_49062);
nand UO_11 (O_11,N_49982,N_49550);
nor UO_12 (O_12,N_48838,N_49449);
or UO_13 (O_13,N_48663,N_47559);
nor UO_14 (O_14,N_48355,N_48202);
and UO_15 (O_15,N_48343,N_47655);
or UO_16 (O_16,N_48551,N_48117);
nand UO_17 (O_17,N_49163,N_48038);
and UO_18 (O_18,N_48547,N_48857);
nor UO_19 (O_19,N_48568,N_48774);
or UO_20 (O_20,N_49013,N_48477);
xnor UO_21 (O_21,N_49992,N_47540);
and UO_22 (O_22,N_47567,N_48375);
or UO_23 (O_23,N_49093,N_48740);
nand UO_24 (O_24,N_48712,N_47735);
or UO_25 (O_25,N_47566,N_48742);
and UO_26 (O_26,N_48772,N_48086);
or UO_27 (O_27,N_48445,N_47676);
xnor UO_28 (O_28,N_47983,N_48408);
or UO_29 (O_29,N_47576,N_48042);
nor UO_30 (O_30,N_48680,N_49418);
and UO_31 (O_31,N_47949,N_48539);
xor UO_32 (O_32,N_47713,N_48161);
or UO_33 (O_33,N_48192,N_47890);
nor UO_34 (O_34,N_47515,N_49560);
or UO_35 (O_35,N_49767,N_47654);
nand UO_36 (O_36,N_48111,N_49978);
or UO_37 (O_37,N_47702,N_49235);
nor UO_38 (O_38,N_48501,N_48827);
and UO_39 (O_39,N_48321,N_49580);
or UO_40 (O_40,N_49243,N_48357);
or UO_41 (O_41,N_47948,N_48993);
xor UO_42 (O_42,N_48065,N_49931);
xnor UO_43 (O_43,N_49472,N_49361);
nand UO_44 (O_44,N_48144,N_49174);
nor UO_45 (O_45,N_48279,N_48107);
or UO_46 (O_46,N_48531,N_47920);
nor UO_47 (O_47,N_48840,N_48260);
xnor UO_48 (O_48,N_49374,N_47614);
xnor UO_49 (O_49,N_49040,N_48284);
or UO_50 (O_50,N_49369,N_49884);
xor UO_51 (O_51,N_48536,N_48781);
and UO_52 (O_52,N_48308,N_47751);
xnor UO_53 (O_53,N_49810,N_48130);
nor UO_54 (O_54,N_48808,N_49469);
nand UO_55 (O_55,N_48055,N_48009);
or UO_56 (O_56,N_48549,N_48913);
xnor UO_57 (O_57,N_47767,N_49249);
xnor UO_58 (O_58,N_48618,N_48407);
nor UO_59 (O_59,N_49822,N_48550);
xnor UO_60 (O_60,N_48719,N_49898);
nor UO_61 (O_61,N_49100,N_48344);
nand UO_62 (O_62,N_48912,N_48608);
nand UO_63 (O_63,N_48815,N_49347);
nor UO_64 (O_64,N_48325,N_48701);
nor UO_65 (O_65,N_49005,N_47901);
nand UO_66 (O_66,N_49983,N_48019);
nand UO_67 (O_67,N_49530,N_48219);
xor UO_68 (O_68,N_49520,N_47869);
and UO_69 (O_69,N_48820,N_49303);
or UO_70 (O_70,N_48890,N_47985);
or UO_71 (O_71,N_48090,N_49824);
nor UO_72 (O_72,N_49494,N_48892);
and UO_73 (O_73,N_49994,N_47938);
and UO_74 (O_74,N_49466,N_48413);
and UO_75 (O_75,N_49358,N_48900);
xnor UO_76 (O_76,N_49948,N_48709);
nand UO_77 (O_77,N_49833,N_49873);
or UO_78 (O_78,N_49535,N_48611);
or UO_79 (O_79,N_49655,N_49363);
xnor UO_80 (O_80,N_49806,N_47777);
or UO_81 (O_81,N_48995,N_48236);
nor UO_82 (O_82,N_48366,N_49099);
and UO_83 (O_83,N_48856,N_49230);
nand UO_84 (O_84,N_48552,N_49792);
nand UO_85 (O_85,N_49667,N_47677);
and UO_86 (O_86,N_48185,N_47894);
and UO_87 (O_87,N_48271,N_47916);
and UO_88 (O_88,N_47990,N_49507);
and UO_89 (O_89,N_49206,N_48410);
nand UO_90 (O_90,N_47957,N_47733);
xnor UO_91 (O_91,N_48240,N_49599);
nor UO_92 (O_92,N_49526,N_49248);
xor UO_93 (O_93,N_49962,N_49740);
nand UO_94 (O_94,N_49323,N_49537);
or UO_95 (O_95,N_47906,N_49447);
nand UO_96 (O_96,N_49777,N_49729);
and UO_97 (O_97,N_47881,N_49279);
xnor UO_98 (O_98,N_48962,N_48356);
or UO_99 (O_99,N_48613,N_49857);
and UO_100 (O_100,N_49272,N_47675);
nand UO_101 (O_101,N_49171,N_48937);
nand UO_102 (O_102,N_49139,N_48761);
xnor UO_103 (O_103,N_47952,N_48254);
and UO_104 (O_104,N_49794,N_49190);
xor UO_105 (O_105,N_48797,N_48959);
and UO_106 (O_106,N_48670,N_47650);
or UO_107 (O_107,N_49016,N_49342);
or UO_108 (O_108,N_47831,N_48770);
xor UO_109 (O_109,N_47725,N_48052);
and UO_110 (O_110,N_48186,N_49886);
and UO_111 (O_111,N_47910,N_48545);
nor UO_112 (O_112,N_48275,N_49207);
nand UO_113 (O_113,N_47928,N_49313);
nor UO_114 (O_114,N_49020,N_48591);
nand UO_115 (O_115,N_47662,N_49928);
nand UO_116 (O_116,N_48004,N_48380);
xnor UO_117 (O_117,N_48403,N_49670);
and UO_118 (O_118,N_47592,N_48690);
nor UO_119 (O_119,N_48949,N_49879);
or UO_120 (O_120,N_47571,N_49198);
nand UO_121 (O_121,N_49021,N_48878);
nor UO_122 (O_122,N_48699,N_48302);
or UO_123 (O_123,N_49628,N_47716);
and UO_124 (O_124,N_47871,N_48832);
nor UO_125 (O_125,N_48510,N_47583);
or UO_126 (O_126,N_48746,N_48923);
nand UO_127 (O_127,N_48030,N_49470);
nand UO_128 (O_128,N_48929,N_49155);
or UO_129 (O_129,N_47714,N_47989);
and UO_130 (O_130,N_47841,N_49122);
and UO_131 (O_131,N_49865,N_49043);
nand UO_132 (O_132,N_47754,N_49722);
nand UO_133 (O_133,N_48533,N_47904);
or UO_134 (O_134,N_48062,N_49430);
nor UO_135 (O_135,N_48603,N_49999);
and UO_136 (O_136,N_49294,N_47726);
nand UO_137 (O_137,N_48232,N_49312);
and UO_138 (O_138,N_49421,N_48886);
nor UO_139 (O_139,N_47613,N_48902);
nor UO_140 (O_140,N_49901,N_47855);
and UO_141 (O_141,N_48685,N_48830);
nand UO_142 (O_142,N_48852,N_48596);
and UO_143 (O_143,N_47525,N_48732);
nor UO_144 (O_144,N_49586,N_48012);
or UO_145 (O_145,N_49710,N_48765);
xor UO_146 (O_146,N_49338,N_48535);
xor UO_147 (O_147,N_48693,N_48530);
or UO_148 (O_148,N_48368,N_49738);
xnor UO_149 (O_149,N_48792,N_48661);
nor UO_150 (O_150,N_48191,N_49402);
or UO_151 (O_151,N_48930,N_47742);
and UO_152 (O_152,N_49675,N_48493);
xor UO_153 (O_153,N_49072,N_48096);
and UO_154 (O_154,N_48140,N_47744);
or UO_155 (O_155,N_48882,N_47924);
nand UO_156 (O_156,N_49913,N_48919);
xor UO_157 (O_157,N_49169,N_47674);
and UO_158 (O_158,N_48983,N_49149);
or UO_159 (O_159,N_49483,N_48903);
and UO_160 (O_160,N_47545,N_48835);
nor UO_161 (O_161,N_48138,N_47641);
and UO_162 (O_162,N_48296,N_47623);
xnor UO_163 (O_163,N_48441,N_48068);
and UO_164 (O_164,N_48958,N_49681);
nor UO_165 (O_165,N_49297,N_48925);
or UO_166 (O_166,N_48187,N_47709);
or UO_167 (O_167,N_48394,N_48115);
and UO_168 (O_168,N_49227,N_48149);
nand UO_169 (O_169,N_49377,N_49378);
nor UO_170 (O_170,N_48581,N_49337);
xor UO_171 (O_171,N_49245,N_49391);
nand UO_172 (O_172,N_49394,N_49219);
or UO_173 (O_173,N_48504,N_49173);
or UO_174 (O_174,N_48378,N_47642);
nand UO_175 (O_175,N_49268,N_49673);
xor UO_176 (O_176,N_48524,N_49410);
xor UO_177 (O_177,N_47937,N_49701);
and UO_178 (O_178,N_49776,N_49785);
nand UO_179 (O_179,N_47762,N_49588);
nand UO_180 (O_180,N_48584,N_48035);
nor UO_181 (O_181,N_49633,N_49465);
nand UO_182 (O_182,N_49053,N_48965);
and UO_183 (O_183,N_48854,N_49622);
or UO_184 (O_184,N_49420,N_49028);
or UO_185 (O_185,N_48287,N_48927);
nand UO_186 (O_186,N_49741,N_49253);
or UO_187 (O_187,N_47973,N_48973);
xor UO_188 (O_188,N_49298,N_48577);
and UO_189 (O_189,N_49422,N_48570);
or UO_190 (O_190,N_49559,N_49208);
xnor UO_191 (O_191,N_48862,N_49168);
nor UO_192 (O_192,N_48682,N_48312);
nor UO_193 (O_193,N_48330,N_48217);
xnor UO_194 (O_194,N_49456,N_49282);
or UO_195 (O_195,N_48258,N_49566);
nor UO_196 (O_196,N_47847,N_48726);
nor UO_197 (O_197,N_49247,N_49136);
xnor UO_198 (O_198,N_48871,N_49400);
or UO_199 (O_199,N_49764,N_47679);
nand UO_200 (O_200,N_47737,N_49582);
nor UO_201 (O_201,N_48988,N_47579);
or UO_202 (O_202,N_47564,N_49625);
or UO_203 (O_203,N_48266,N_48869);
nor UO_204 (O_204,N_49784,N_49499);
nand UO_205 (O_205,N_49343,N_47543);
or UO_206 (O_206,N_48969,N_48724);
nand UO_207 (O_207,N_48294,N_48331);
or UO_208 (O_208,N_48448,N_49787);
and UO_209 (O_209,N_49316,N_48909);
or UO_210 (O_210,N_48388,N_49842);
nor UO_211 (O_211,N_48780,N_47886);
nand UO_212 (O_212,N_47604,N_49441);
or UO_213 (O_213,N_47731,N_49089);
xor UO_214 (O_214,N_49646,N_48645);
nor UO_215 (O_215,N_49195,N_49172);
xor UO_216 (O_216,N_49284,N_48692);
and UO_217 (O_217,N_47562,N_47892);
nor UO_218 (O_218,N_47982,N_49736);
xor UO_219 (O_219,N_49295,N_49632);
xnor UO_220 (O_220,N_49866,N_48938);
xor UO_221 (O_221,N_49647,N_48595);
or UO_222 (O_222,N_49370,N_49527);
and UO_223 (O_223,N_48710,N_48752);
xnor UO_224 (O_224,N_48195,N_48006);
or UO_225 (O_225,N_47774,N_48422);
nand UO_226 (O_226,N_49360,N_48861);
or UO_227 (O_227,N_48048,N_47805);
xnor UO_228 (O_228,N_49024,N_49367);
or UO_229 (O_229,N_47599,N_48679);
nand UO_230 (O_230,N_47658,N_49797);
or UO_231 (O_231,N_48114,N_47801);
nand UO_232 (O_232,N_48200,N_49678);
xnor UO_233 (O_233,N_49627,N_47556);
nand UO_234 (O_234,N_48961,N_49322);
nand UO_235 (O_235,N_48429,N_49604);
and UO_236 (O_236,N_48750,N_49837);
xnor UO_237 (O_237,N_48390,N_49061);
or UO_238 (O_238,N_48437,N_47585);
and UO_239 (O_239,N_49228,N_49471);
nor UO_240 (O_240,N_49073,N_47836);
or UO_241 (O_241,N_49652,N_49751);
nand UO_242 (O_242,N_48371,N_49576);
or UO_243 (O_243,N_49821,N_48346);
nand UO_244 (O_244,N_49657,N_48461);
xor UO_245 (O_245,N_48879,N_49540);
nand UO_246 (O_246,N_47999,N_49944);
nor UO_247 (O_247,N_47551,N_48257);
nor UO_248 (O_248,N_48348,N_49334);
or UO_249 (O_249,N_48332,N_47776);
or UO_250 (O_250,N_48087,N_47612);
xnor UO_251 (O_251,N_49350,N_48480);
xnor UO_252 (O_252,N_48858,N_48451);
nand UO_253 (O_253,N_49607,N_47729);
nand UO_254 (O_254,N_48771,N_48132);
nor UO_255 (O_255,N_48521,N_47902);
or UO_256 (O_256,N_47979,N_49444);
nor UO_257 (O_257,N_48458,N_49146);
nand UO_258 (O_258,N_49427,N_48809);
and UO_259 (O_259,N_49927,N_48142);
nand UO_260 (O_260,N_47561,N_48867);
nor UO_261 (O_261,N_48075,N_49862);
or UO_262 (O_262,N_49570,N_48311);
nor UO_263 (O_263,N_48415,N_49068);
and UO_264 (O_264,N_48665,N_49092);
and UO_265 (O_265,N_48083,N_49086);
nand UO_266 (O_266,N_48970,N_48310);
nor UO_267 (O_267,N_49330,N_48617);
nor UO_268 (O_268,N_48743,N_48070);
nand UO_269 (O_269,N_49424,N_48383);
or UO_270 (O_270,N_49423,N_49845);
xor UO_271 (O_271,N_47514,N_47833);
or UO_272 (O_272,N_48876,N_48245);
or UO_273 (O_273,N_49548,N_49727);
and UO_274 (O_274,N_49179,N_49803);
and UO_275 (O_275,N_47644,N_48518);
nand UO_276 (O_276,N_48498,N_49936);
xor UO_277 (O_277,N_49734,N_49809);
nand UO_278 (O_278,N_48756,N_49695);
nand UO_279 (O_279,N_48528,N_48206);
and UO_280 (O_280,N_47789,N_49014);
or UO_281 (O_281,N_49079,N_48024);
nand UO_282 (O_282,N_48031,N_49194);
or UO_283 (O_283,N_49603,N_48382);
and UO_284 (O_284,N_49754,N_47548);
xnor UO_285 (O_285,N_47997,N_48241);
or UO_286 (O_286,N_48265,N_49869);
and UO_287 (O_287,N_47670,N_47897);
xor UO_288 (O_288,N_49595,N_47877);
xor UO_289 (O_289,N_48606,N_47505);
xnor UO_290 (O_290,N_48704,N_47967);
nor UO_291 (O_291,N_49409,N_49831);
and UO_292 (O_292,N_48264,N_49849);
nand UO_293 (O_293,N_49443,N_47965);
and UO_294 (O_294,N_49800,N_48252);
xnor UO_295 (O_295,N_49356,N_47528);
or UO_296 (O_296,N_49906,N_48060);
or UO_297 (O_297,N_48324,N_48678);
nand UO_298 (O_298,N_49166,N_49060);
xnor UO_299 (O_299,N_49706,N_49065);
xor UO_300 (O_300,N_48507,N_49140);
nand UO_301 (O_301,N_47539,N_48872);
and UO_302 (O_302,N_48837,N_49629);
and UO_303 (O_303,N_47602,N_49623);
or UO_304 (O_304,N_49197,N_49708);
xor UO_305 (O_305,N_48339,N_48691);
xnor UO_306 (O_306,N_49047,N_48529);
or UO_307 (O_307,N_48826,N_48667);
and UO_308 (O_308,N_49055,N_48370);
and UO_309 (O_309,N_49445,N_48351);
or UO_310 (O_310,N_49131,N_49574);
xor UO_311 (O_311,N_48464,N_48306);
and UO_312 (O_312,N_48141,N_47740);
nand UO_313 (O_313,N_48505,N_48406);
and UO_314 (O_314,N_49691,N_48102);
or UO_315 (O_315,N_49916,N_48384);
nor UO_316 (O_316,N_48492,N_49329);
xnor UO_317 (O_317,N_47589,N_48885);
nor UO_318 (O_318,N_49010,N_47511);
nand UO_319 (O_319,N_49150,N_47582);
or UO_320 (O_320,N_48011,N_48419);
or UO_321 (O_321,N_48788,N_48555);
nand UO_322 (O_322,N_48513,N_49032);
xnor UO_323 (O_323,N_48466,N_49658);
and UO_324 (O_324,N_48433,N_48478);
nand UO_325 (O_325,N_49383,N_48653);
nand UO_326 (O_326,N_49119,N_49209);
nor UO_327 (O_327,N_47680,N_47653);
nand UO_328 (O_328,N_48696,N_48801);
xor UO_329 (O_329,N_49861,N_48850);
nand UO_330 (O_330,N_48082,N_47667);
nand UO_331 (O_331,N_49460,N_47581);
nand UO_332 (O_332,N_48672,N_48899);
and UO_333 (O_333,N_49379,N_49500);
xor UO_334 (O_334,N_49293,N_49154);
xor UO_335 (O_335,N_48677,N_47747);
nor UO_336 (O_336,N_47666,N_49731);
and UO_337 (O_337,N_49232,N_47531);
nand UO_338 (O_338,N_49083,N_48798);
or UO_339 (O_339,N_49897,N_48588);
xor UO_340 (O_340,N_49307,N_48320);
nand UO_341 (O_341,N_48669,N_48424);
or UO_342 (O_342,N_49276,N_47668);
and UO_343 (O_343,N_48123,N_49735);
xnor UO_344 (O_344,N_47624,N_48301);
xor UO_345 (O_345,N_48565,N_48490);
or UO_346 (O_346,N_48508,N_49143);
and UO_347 (O_347,N_49805,N_47988);
xnor UO_348 (O_348,N_49022,N_49640);
or UO_349 (O_349,N_49593,N_49656);
and UO_350 (O_350,N_49674,N_48046);
xor UO_351 (O_351,N_48485,N_48379);
or UO_352 (O_352,N_49502,N_49528);
or UO_353 (O_353,N_49853,N_49000);
nand UO_354 (O_354,N_49683,N_48463);
nor UO_355 (O_355,N_49795,N_48722);
nand UO_356 (O_356,N_49988,N_49608);
or UO_357 (O_357,N_48034,N_47934);
xnor UO_358 (O_358,N_49668,N_48465);
or UO_359 (O_359,N_49462,N_49644);
nand UO_360 (O_360,N_48675,N_49493);
nor UO_361 (O_361,N_49707,N_49711);
nand UO_362 (O_362,N_49807,N_49920);
nor UO_363 (O_363,N_49152,N_47784);
xor UO_364 (O_364,N_49917,N_47885);
xor UO_365 (O_365,N_49868,N_48566);
xnor UO_366 (O_366,N_48713,N_49182);
nand UO_367 (O_367,N_48762,N_48579);
and UO_368 (O_368,N_47739,N_49375);
nand UO_369 (O_369,N_49568,N_48749);
xnor UO_370 (O_370,N_47537,N_47665);
or UO_371 (O_371,N_47526,N_49684);
or UO_372 (O_372,N_49895,N_49258);
and UO_373 (O_373,N_48334,N_48715);
nand UO_374 (O_374,N_48362,N_48328);
nor UO_375 (O_375,N_47970,N_49859);
or UO_376 (O_376,N_48975,N_47608);
and UO_377 (O_377,N_49968,N_48818);
xnor UO_378 (O_378,N_49121,N_48127);
and UO_379 (O_379,N_48790,N_48883);
and UO_380 (O_380,N_47943,N_47752);
xnor UO_381 (O_381,N_48196,N_49035);
and UO_382 (O_382,N_49511,N_48483);
xnor UO_383 (O_383,N_48889,N_47698);
xor UO_384 (O_384,N_49737,N_48457);
or UO_385 (O_385,N_47683,N_49932);
and UO_386 (O_386,N_48354,N_48439);
nor UO_387 (O_387,N_48853,N_48474);
or UO_388 (O_388,N_48720,N_49091);
xor UO_389 (O_389,N_47763,N_48204);
and UO_390 (O_390,N_49941,N_49934);
xor UO_391 (O_391,N_49720,N_48554);
or UO_392 (O_392,N_48649,N_48643);
nor UO_393 (O_393,N_48033,N_48246);
or UO_394 (O_394,N_49301,N_49645);
or UO_395 (O_395,N_47617,N_48174);
and UO_396 (O_396,N_49244,N_49698);
nor UO_397 (O_397,N_47693,N_49225);
or UO_398 (O_398,N_48242,N_47980);
nand UO_399 (O_399,N_49183,N_48015);
nor UO_400 (O_400,N_49218,N_47977);
and UO_401 (O_401,N_48844,N_49894);
xnor UO_402 (O_402,N_49521,N_49848);
or UO_403 (O_403,N_47756,N_48162);
nand UO_404 (O_404,N_48077,N_49964);
nor UO_405 (O_405,N_47874,N_49362);
nor UO_406 (O_406,N_47945,N_47637);
and UO_407 (O_407,N_49651,N_49408);
nor UO_408 (O_408,N_49503,N_48706);
xnor UO_409 (O_409,N_47656,N_49027);
xnor UO_410 (O_410,N_47931,N_49191);
nand UO_411 (O_411,N_49946,N_47758);
xor UO_412 (O_412,N_48164,N_47879);
and UO_413 (O_413,N_48952,N_48108);
nor UO_414 (O_414,N_47984,N_49867);
and UO_415 (O_415,N_48751,N_49662);
nand UO_416 (O_416,N_49546,N_49610);
nor UO_417 (O_417,N_49478,N_47663);
and UO_418 (O_418,N_49257,N_47711);
or UO_419 (O_419,N_48175,N_48432);
xnor UO_420 (O_420,N_47597,N_47659);
and UO_421 (O_421,N_49271,N_49984);
and UO_422 (O_422,N_48340,N_48233);
and UO_423 (O_423,N_49193,N_49440);
and UO_424 (O_424,N_48342,N_49529);
and UO_425 (O_425,N_47810,N_48847);
or UO_426 (O_426,N_48932,N_49125);
and UO_427 (O_427,N_49349,N_48874);
or UO_428 (O_428,N_48776,N_49545);
and UO_429 (O_429,N_48273,N_48986);
nor UO_430 (O_430,N_49355,N_47816);
or UO_431 (O_431,N_49957,N_48253);
nand UO_432 (O_432,N_49732,N_49929);
xnor UO_433 (O_433,N_48951,N_48182);
xnor UO_434 (O_434,N_49649,N_47821);
and UO_435 (O_435,N_48974,N_47768);
or UO_436 (O_436,N_47813,N_47701);
and UO_437 (O_437,N_48003,N_49843);
nor UO_438 (O_438,N_49600,N_48314);
nand UO_439 (O_439,N_47760,N_47799);
or UO_440 (O_440,N_47862,N_49816);
and UO_441 (O_441,N_48147,N_49716);
xnor UO_442 (O_442,N_49543,N_47504);
nor UO_443 (O_443,N_48814,N_48361);
nor UO_444 (O_444,N_47958,N_48101);
and UO_445 (O_445,N_49554,N_47827);
and UO_446 (O_446,N_49517,N_47893);
nor UO_447 (O_447,N_47909,N_49054);
xor UO_448 (O_448,N_48036,N_48526);
and UO_449 (O_449,N_49796,N_49963);
nand UO_450 (O_450,N_48179,N_49057);
xor UO_451 (O_451,N_47502,N_49660);
xor UO_452 (O_452,N_49260,N_49592);
nor UO_453 (O_453,N_48274,N_49203);
and UO_454 (O_454,N_48664,N_47689);
and UO_455 (O_455,N_48702,N_47941);
and UO_456 (O_456,N_49752,N_49385);
and UO_457 (O_457,N_48532,N_48599);
xnor UO_458 (O_458,N_48673,N_49763);
or UO_459 (O_459,N_48911,N_49281);
nand UO_460 (O_460,N_47640,N_48683);
nand UO_461 (O_461,N_47630,N_48151);
xor UO_462 (O_462,N_48040,N_48404);
and UO_463 (O_463,N_48578,N_47880);
xor UO_464 (O_464,N_47746,N_49778);
nand UO_465 (O_465,N_49856,N_48631);
and UO_466 (O_466,N_47552,N_48402);
xnor UO_467 (O_467,N_47765,N_48178);
nand UO_468 (O_468,N_49419,N_49538);
and UO_469 (O_469,N_48697,N_48481);
nor UO_470 (O_470,N_47738,N_49542);
xnor UO_471 (O_471,N_49184,N_47569);
nand UO_472 (O_472,N_47621,N_49614);
nor UO_473 (O_473,N_48904,N_48262);
nand UO_474 (O_474,N_49650,N_48405);
and UO_475 (O_475,N_48707,N_48527);
or UO_476 (O_476,N_48159,N_48557);
and UO_477 (O_477,N_48304,N_48897);
nor UO_478 (O_478,N_49261,N_49951);
nor UO_479 (O_479,N_48373,N_48560);
and UO_480 (O_480,N_49002,N_47783);
or UO_481 (O_481,N_49240,N_48793);
and UO_482 (O_482,N_47809,N_49976);
and UO_483 (O_483,N_49264,N_48764);
nand UO_484 (O_484,N_47598,N_48278);
or UO_485 (O_485,N_49464,N_49045);
and UO_486 (O_486,N_49819,N_47806);
nor UO_487 (O_487,N_49346,N_49986);
xnor UO_488 (O_488,N_48625,N_47594);
xor UO_489 (O_489,N_48450,N_48243);
or UO_490 (O_490,N_48968,N_47769);
xnor UO_491 (O_491,N_48455,N_48352);
or UO_492 (O_492,N_49860,N_47523);
and UO_493 (O_493,N_49685,N_49486);
nor UO_494 (O_494,N_48305,N_49158);
nand UO_495 (O_495,N_49433,N_49101);
xnor UO_496 (O_496,N_48081,N_49405);
or UO_497 (O_497,N_47724,N_49270);
nand UO_498 (O_498,N_48285,N_47927);
nor UO_499 (O_499,N_49274,N_47820);
nor UO_500 (O_500,N_47529,N_48594);
nor UO_501 (O_501,N_49863,N_48280);
nand UO_502 (O_502,N_48639,N_48747);
and UO_503 (O_503,N_49786,N_47944);
nand UO_504 (O_504,N_48979,N_48126);
or UO_505 (O_505,N_49145,N_49739);
xor UO_506 (O_506,N_49196,N_48165);
xnor UO_507 (O_507,N_49359,N_47578);
nand UO_508 (O_508,N_49048,N_48128);
and UO_509 (O_509,N_49575,N_48586);
nor UO_510 (O_510,N_48152,N_48244);
or UO_511 (O_511,N_48157,N_49745);
nand UO_512 (O_512,N_49354,N_47753);
nand UO_513 (O_513,N_48261,N_48870);
and UO_514 (O_514,N_49215,N_49001);
or UO_515 (O_515,N_48777,N_49531);
nand UO_516 (O_516,N_49098,N_48222);
or UO_517 (O_517,N_49509,N_48263);
nand UO_518 (O_518,N_48020,N_49998);
nand UO_519 (O_519,N_47745,N_47922);
nand UO_520 (O_520,N_47596,N_48976);
nand UO_521 (O_521,N_48652,N_49373);
nand UO_522 (O_522,N_48802,N_49105);
xnor UO_523 (O_523,N_49156,N_49746);
nor UO_524 (O_524,N_49573,N_48456);
nor UO_525 (O_525,N_48488,N_49760);
xnor UO_526 (O_526,N_48967,N_49563);
nor UO_527 (O_527,N_47895,N_48435);
nor UO_528 (O_528,N_49890,N_49990);
nand UO_529 (O_529,N_49508,N_48650);
xor UO_530 (O_530,N_47625,N_49417);
nand UO_531 (O_531,N_47870,N_48748);
nand UO_532 (O_532,N_48829,N_49266);
and UO_533 (O_533,N_47509,N_49761);
nor UO_534 (O_534,N_49023,N_47542);
nor UO_535 (O_535,N_48372,N_49669);
nand UO_536 (O_536,N_47757,N_47518);
or UO_537 (O_537,N_49613,N_49468);
or UO_538 (O_538,N_47778,N_49426);
nand UO_539 (O_539,N_47527,N_49631);
xor UO_540 (O_540,N_49715,N_47946);
nand UO_541 (O_541,N_49581,N_48616);
xor UO_542 (O_542,N_48199,N_48646);
nand UO_543 (O_543,N_48917,N_49463);
nor UO_544 (O_544,N_48896,N_48092);
nand UO_545 (O_545,N_49938,N_49770);
and UO_546 (O_546,N_49768,N_49971);
nand UO_547 (O_547,N_49799,N_49498);
nor UO_548 (O_548,N_49340,N_49484);
xor UO_549 (O_549,N_48471,N_47969);
nor UO_550 (O_550,N_47876,N_48898);
xnor UO_551 (O_551,N_47773,N_47811);
or UO_552 (O_552,N_47521,N_49609);
xnor UO_553 (O_553,N_49973,N_47684);
nor UO_554 (O_554,N_49980,N_48010);
and UO_555 (O_555,N_49159,N_49157);
and UO_556 (O_556,N_49481,N_49029);
xnor UO_557 (O_557,N_48239,N_47878);
or UO_558 (O_558,N_48633,N_47708);
xnor UO_559 (O_559,N_47796,N_49115);
and UO_560 (O_560,N_48991,N_49479);
nor UO_561 (O_561,N_47883,N_47535);
and UO_562 (O_562,N_48905,N_48946);
or UO_563 (O_563,N_47699,N_48880);
or UO_564 (O_564,N_49721,N_48166);
nand UO_565 (O_565,N_47823,N_49459);
nor UO_566 (O_566,N_47717,N_48908);
or UO_567 (O_567,N_49438,N_49031);
nand UO_568 (O_568,N_48884,N_48943);
or UO_569 (O_569,N_49714,N_49128);
nor UO_570 (O_570,N_49606,N_49648);
xnor UO_571 (O_571,N_49454,N_49620);
nand UO_572 (O_572,N_49801,N_48572);
nor UO_573 (O_573,N_48635,N_47759);
or UO_574 (O_574,N_49003,N_49214);
or UO_575 (O_575,N_49789,N_49049);
nor UO_576 (O_576,N_49730,N_47794);
nor UO_577 (O_577,N_48597,N_48738);
nor UO_578 (O_578,N_49914,N_49137);
xnor UO_579 (O_579,N_47971,N_49827);
xor UO_580 (O_580,N_49304,N_48453);
or UO_581 (O_581,N_48224,N_49557);
xor UO_582 (O_582,N_49536,N_49510);
nand UO_583 (O_583,N_47903,N_48449);
nor UO_584 (O_584,N_48948,N_47950);
or UO_585 (O_585,N_48516,N_48695);
nor UO_586 (O_586,N_49432,N_48816);
and UO_587 (O_587,N_47712,N_49496);
nand UO_588 (O_588,N_49275,N_48177);
and UO_589 (O_589,N_49050,N_49344);
nand UO_590 (O_590,N_48769,N_48421);
and UO_591 (O_591,N_47695,N_48796);
nand UO_592 (O_592,N_49017,N_49317);
or UO_593 (O_593,N_47936,N_48323);
xor UO_594 (O_594,N_48438,N_48783);
or UO_595 (O_595,N_47730,N_49129);
and UO_596 (O_596,N_48014,N_48299);
or UO_597 (O_597,N_49826,N_49170);
nand UO_598 (O_598,N_48071,N_49779);
or UO_599 (O_599,N_48745,N_49309);
nand UO_600 (O_600,N_47646,N_48767);
xnor UO_601 (O_601,N_47618,N_47771);
nor UO_602 (O_602,N_49012,N_49598);
and UO_603 (O_603,N_49448,N_48576);
or UO_604 (O_604,N_49758,N_49713);
or UO_605 (O_605,N_48700,N_47887);
nor UO_606 (O_606,N_48487,N_47547);
and UO_607 (O_607,N_49889,N_49724);
nor UO_608 (O_608,N_49933,N_48607);
or UO_609 (O_609,N_47975,N_47852);
or UO_610 (O_610,N_49522,N_48721);
or UO_611 (O_611,N_49775,N_48017);
nand UO_612 (O_612,N_49584,N_49058);
and UO_613 (O_613,N_47800,N_48733);
nor UO_614 (O_614,N_47803,N_49686);
nor UO_615 (O_615,N_49905,N_48160);
nand UO_616 (O_616,N_48105,N_48215);
nand UO_617 (O_617,N_49549,N_49900);
xnor UO_618 (O_618,N_49106,N_49967);
or UO_619 (O_619,N_48520,N_48290);
nor UO_620 (O_620,N_49221,N_48918);
and UO_621 (O_621,N_48176,N_48725);
nand UO_622 (O_622,N_47616,N_49943);
and UO_623 (O_623,N_48039,N_49280);
and UO_624 (O_624,N_48051,N_48063);
or UO_625 (O_625,N_48605,N_49975);
and UO_626 (O_626,N_49491,N_49783);
nand UO_627 (O_627,N_49991,N_49039);
and UO_628 (O_628,N_49116,N_47575);
nor UO_629 (O_629,N_48148,N_48313);
or UO_630 (O_630,N_49401,N_48634);
or UO_631 (O_631,N_47645,N_49591);
or UO_632 (O_632,N_49742,N_49429);
and UO_633 (O_633,N_49995,N_49911);
xor UO_634 (O_634,N_48289,N_48183);
nor UO_635 (O_635,N_49782,N_49368);
nand UO_636 (O_636,N_49780,N_48915);
nor UO_637 (O_637,N_49103,N_48440);
and UO_638 (O_638,N_49876,N_48868);
nor UO_639 (O_639,N_48118,N_48763);
xor UO_640 (O_640,N_47636,N_48249);
or UO_641 (O_641,N_49504,N_47914);
nand UO_642 (O_642,N_49555,N_48966);
nor UO_643 (O_643,N_48694,N_47824);
and UO_644 (O_644,N_49829,N_48999);
nand UO_645 (O_645,N_48172,N_48377);
or UO_646 (O_646,N_47933,N_49619);
nor UO_647 (O_647,N_47998,N_48078);
nor UO_648 (O_648,N_49970,N_47550);
xnor UO_649 (O_649,N_47839,N_49063);
nand UO_650 (O_650,N_49416,N_47891);
nand UO_651 (O_651,N_48153,N_49328);
nor UO_652 (O_652,N_49888,N_49387);
and UO_653 (O_653,N_49160,N_48981);
and UO_654 (O_654,N_49425,N_49286);
xnor UO_655 (O_655,N_48604,N_48475);
and UO_656 (O_656,N_48234,N_48662);
nor UO_657 (O_657,N_48256,N_49518);
nor UO_658 (O_658,N_49132,N_49224);
or UO_659 (O_659,N_49825,N_48674);
or UO_660 (O_660,N_48562,N_48811);
xnor UO_661 (O_661,N_47588,N_48298);
nor UO_662 (O_662,N_49386,N_48523);
and UO_663 (O_663,N_47587,N_48602);
and UO_664 (O_664,N_49388,N_49544);
nor UO_665 (O_665,N_47995,N_47593);
xnor UO_666 (O_666,N_48624,N_49220);
xor UO_667 (O_667,N_49326,N_48129);
nand UO_668 (O_668,N_48411,N_49009);
nand UO_669 (O_669,N_47918,N_49692);
or UO_670 (O_670,N_48391,N_48259);
and UO_671 (O_671,N_49743,N_47986);
or UO_672 (O_672,N_48454,N_48489);
nor UO_673 (O_673,N_49955,N_48583);
nand UO_674 (O_674,N_48519,N_49398);
xnor UO_675 (O_675,N_49952,N_47568);
xnor UO_676 (O_676,N_48369,N_47691);
nor UO_677 (O_677,N_48960,N_47673);
and UO_678 (O_678,N_48590,N_47775);
nand UO_679 (O_679,N_48546,N_48647);
or UO_680 (O_680,N_47687,N_48573);
or UO_681 (O_681,N_49870,N_47710);
nand UO_682 (O_682,N_49492,N_49283);
nor UO_683 (O_683,N_49457,N_49700);
or UO_684 (O_684,N_49041,N_48648);
nand UO_685 (O_685,N_48297,N_48427);
or UO_686 (O_686,N_48718,N_48089);
xor UO_687 (O_687,N_48281,N_48760);
and UO_688 (O_688,N_47959,N_47956);
xnor UO_689 (O_689,N_48657,N_49590);
xnor UO_690 (O_690,N_48171,N_48980);
and UO_691 (O_691,N_48345,N_47842);
xnor UO_692 (O_692,N_48877,N_47857);
xor UO_693 (O_693,N_48541,N_48389);
xnor UO_694 (O_694,N_48623,N_47610);
nand UO_695 (O_695,N_48103,N_47797);
xnor UO_696 (O_696,N_49396,N_48553);
nor UO_697 (O_697,N_48642,N_49665);
xor UO_698 (O_698,N_49664,N_49109);
and UO_699 (O_699,N_48385,N_49175);
xor UO_700 (O_700,N_48119,N_49406);
xnor UO_701 (O_701,N_48116,N_47672);
xnor UO_702 (O_702,N_49878,N_49165);
xor UO_703 (O_703,N_49514,N_49719);
and UO_704 (O_704,N_48775,N_48235);
nand UO_705 (O_705,N_48836,N_49516);
or UO_706 (O_706,N_49395,N_49376);
xor UO_707 (O_707,N_49151,N_48091);
nand UO_708 (O_708,N_48218,N_49331);
nand UO_709 (O_709,N_48131,N_49310);
xor UO_710 (O_710,N_47634,N_47908);
nor UO_711 (O_711,N_49663,N_49059);
and UO_712 (O_712,N_48088,N_48431);
and UO_713 (O_713,N_49909,N_49318);
and UO_714 (O_714,N_48423,N_49308);
and UO_715 (O_715,N_48381,N_49688);
nand UO_716 (O_716,N_49138,N_48587);
nor UO_717 (O_717,N_49475,N_48758);
and UO_718 (O_718,N_48580,N_48399);
and UO_719 (O_719,N_48223,N_47619);
nor UO_720 (O_720,N_47817,N_49987);
xnor UO_721 (O_721,N_49565,N_48998);
or UO_722 (O_722,N_48316,N_49036);
nor UO_723 (O_723,N_49693,N_49412);
and UO_724 (O_724,N_49153,N_48768);
nor UO_725 (O_725,N_49512,N_49497);
or UO_726 (O_726,N_49082,N_49748);
nor UO_727 (O_727,N_48766,N_49108);
nand UO_728 (O_728,N_49823,N_48825);
nor UO_729 (O_729,N_49924,N_49102);
xnor UO_730 (O_730,N_49630,N_47755);
and UO_731 (O_731,N_49912,N_48135);
nand UO_732 (O_732,N_47963,N_47506);
nand UO_733 (O_733,N_48250,N_49181);
or UO_734 (O_734,N_49025,N_49246);
and UO_735 (O_735,N_47832,N_48412);
or UO_736 (O_736,N_48924,N_48338);
xnor UO_737 (O_737,N_48716,N_47872);
xor UO_738 (O_738,N_49945,N_47899);
and UO_739 (O_739,N_49450,N_49832);
and UO_740 (O_740,N_48396,N_49793);
and UO_741 (O_741,N_47843,N_48730);
nand UO_742 (O_742,N_48538,N_49222);
and UO_743 (O_743,N_47818,N_47516);
nand UO_744 (O_744,N_49993,N_49682);
xnor UO_745 (O_745,N_48326,N_48841);
or UO_746 (O_746,N_47930,N_47743);
nor UO_747 (O_747,N_49696,N_48703);
or UO_748 (O_748,N_47981,N_47907);
or UO_749 (O_749,N_48632,N_47786);
or UO_750 (O_750,N_48134,N_49704);
nand UO_751 (O_751,N_48828,N_48336);
or UO_752 (O_752,N_49892,N_47912);
nand UO_753 (O_753,N_48708,N_48600);
nand UO_754 (O_754,N_48016,N_48397);
xnor UO_755 (O_755,N_48181,N_49858);
or UO_756 (O_756,N_49596,N_47722);
nand UO_757 (O_757,N_49488,N_47802);
nand UO_758 (O_758,N_49534,N_49874);
or UO_759 (O_759,N_48001,N_48689);
and UO_760 (O_760,N_49044,N_47560);
xnor UO_761 (O_761,N_49774,N_48942);
or UO_762 (O_762,N_48335,N_49269);
xor UO_763 (O_763,N_48085,N_48786);
nand UO_764 (O_764,N_48659,N_48782);
and UO_765 (O_765,N_49127,N_49381);
xnor UO_766 (O_766,N_48851,N_48277);
xor UO_767 (O_767,N_48916,N_49712);
nand UO_768 (O_768,N_48270,N_49142);
xor UO_769 (O_769,N_49004,N_49515);
and UO_770 (O_770,N_48150,N_47923);
or UO_771 (O_771,N_48211,N_48363);
nand UO_772 (O_772,N_47830,N_48154);
nor UO_773 (O_773,N_48137,N_48064);
nor UO_774 (O_774,N_47538,N_49855);
or UO_775 (O_775,N_48957,N_47639);
and UO_776 (O_776,N_48163,N_48864);
or UO_777 (O_777,N_47546,N_48887);
xor UO_778 (O_778,N_48337,N_49838);
nand UO_779 (O_779,N_49533,N_49567);
and UO_780 (O_780,N_49130,N_48027);
xor UO_781 (O_781,N_47868,N_47508);
xor UO_782 (O_782,N_47856,N_49558);
xnor UO_783 (O_783,N_47900,N_48935);
or UO_784 (O_784,N_47741,N_49506);
nand UO_785 (O_785,N_49141,N_49757);
nor UO_786 (O_786,N_48789,N_48374);
and UO_787 (O_787,N_47845,N_48099);
or UO_788 (O_788,N_48209,N_49111);
nand UO_789 (O_789,N_48734,N_48687);
or UO_790 (O_790,N_49327,N_49026);
xor UO_791 (O_791,N_48460,N_47960);
and UO_792 (O_792,N_49587,N_48574);
and UO_793 (O_793,N_48146,N_48963);
and UO_794 (O_794,N_49126,N_47524);
nor UO_795 (O_795,N_48512,N_48100);
and UO_796 (O_796,N_49033,N_47860);
xor UO_797 (O_797,N_49697,N_49285);
nand UO_798 (O_798,N_48994,N_47700);
or UO_799 (O_799,N_49234,N_49335);
or UO_800 (O_800,N_47812,N_48468);
xor UO_801 (O_801,N_49178,N_49201);
xor UO_802 (O_802,N_49452,N_48367);
nand UO_803 (O_803,N_49818,N_49840);
or UO_804 (O_804,N_47867,N_48443);
nand UO_805 (O_805,N_48655,N_49960);
and UO_806 (O_806,N_48585,N_49380);
nor UO_807 (O_807,N_49766,N_49135);
or UO_808 (O_808,N_49847,N_48660);
xnor UO_809 (O_809,N_49850,N_49887);
xnor UO_810 (O_810,N_48341,N_47622);
nor UO_811 (O_811,N_48681,N_49299);
nand UO_812 (O_812,N_48630,N_48891);
nand UO_813 (O_813,N_47520,N_47788);
nor UO_814 (O_814,N_48548,N_47607);
or UO_815 (O_815,N_47849,N_49547);
and UO_816 (O_816,N_48881,N_49015);
xnor UO_817 (O_817,N_49180,N_47911);
xnor UO_818 (O_818,N_49921,N_47595);
and UO_819 (O_819,N_49882,N_47727);
nand UO_820 (O_820,N_49985,N_49718);
xor UO_821 (O_821,N_48926,N_48522);
xor UO_822 (O_822,N_47522,N_48084);
nor UO_823 (O_823,N_47972,N_48400);
and UO_824 (O_824,N_48728,N_49439);
nor UO_825 (O_825,N_49654,N_48401);
nand UO_826 (O_826,N_49167,N_48947);
nor UO_827 (O_827,N_48452,N_48267);
and UO_828 (O_828,N_48459,N_47947);
xnor UO_829 (O_829,N_47819,N_48420);
nor UO_830 (O_830,N_48276,N_48426);
and UO_831 (O_831,N_49689,N_49872);
nor UO_832 (O_832,N_48189,N_49407);
nand UO_833 (O_833,N_47690,N_49428);
xor UO_834 (O_834,N_49597,N_49357);
nor UO_835 (O_835,N_48614,N_48741);
nor UO_836 (O_836,N_47734,N_49051);
or UO_837 (O_837,N_49877,N_48013);
xor UO_838 (O_838,N_49090,N_48817);
nor UO_839 (O_839,N_47541,N_48364);
or UO_840 (O_840,N_48469,N_49262);
xor UO_841 (O_841,N_47835,N_49844);
or UO_842 (O_842,N_49353,N_47861);
and UO_843 (O_843,N_48755,N_48711);
or UO_844 (O_844,N_48225,N_48727);
and UO_845 (O_845,N_49699,N_48418);
nand UO_846 (O_846,N_49291,N_49578);
or UO_847 (O_847,N_49110,N_48514);
or UO_848 (O_848,N_49213,N_48145);
nor UO_849 (O_849,N_49616,N_47859);
and UO_850 (O_850,N_49431,N_48839);
or UO_851 (O_851,N_48282,N_48293);
xor UO_852 (O_852,N_47761,N_47992);
and UO_853 (O_853,N_48803,N_47785);
nor UO_854 (O_854,N_49830,N_49384);
nand UO_855 (O_855,N_49052,N_49680);
or UO_856 (O_856,N_49661,N_48509);
and UO_857 (O_857,N_48053,N_48169);
or UO_858 (O_858,N_48292,N_48737);
nor UO_859 (O_859,N_48525,N_47682);
and UO_860 (O_860,N_47815,N_47565);
xnor UO_861 (O_861,N_49321,N_47889);
and UO_862 (O_862,N_48008,N_49852);
and UO_863 (O_863,N_47605,N_48247);
xor UO_864 (O_864,N_49278,N_49458);
and UO_865 (O_865,N_48120,N_49839);
and UO_866 (O_866,N_49828,N_49277);
xnor UO_867 (O_867,N_47932,N_49332);
nor UO_868 (O_868,N_49114,N_49919);
or UO_869 (O_869,N_48170,N_48944);
nor UO_870 (O_870,N_48644,N_49034);
nor UO_871 (O_871,N_48953,N_49097);
xor UO_872 (O_872,N_49075,N_48188);
nor UO_873 (O_873,N_49601,N_49659);
xor UO_874 (O_874,N_49080,N_48446);
and UO_875 (O_875,N_48619,N_48495);
or UO_876 (O_876,N_49676,N_49042);
nor UO_877 (O_877,N_48018,N_49148);
nand UO_878 (O_878,N_49679,N_49773);
nand UO_879 (O_879,N_48824,N_48987);
nand UO_880 (O_880,N_48609,N_48859);
xor UO_881 (O_881,N_48823,N_48705);
xor UO_882 (O_882,N_49896,N_49750);
and UO_883 (O_883,N_49164,N_49733);
xnor UO_884 (O_884,N_48821,N_48698);
xor UO_885 (O_885,N_48941,N_47657);
nor UO_886 (O_886,N_48910,N_49638);
nand UO_887 (O_887,N_48112,N_48268);
or UO_888 (O_888,N_48804,N_48497);
nor UO_889 (O_889,N_48156,N_47858);
nand UO_890 (O_890,N_49290,N_49302);
nor UO_891 (O_891,N_49480,N_48515);
xor UO_892 (O_892,N_48540,N_47828);
and UO_893 (O_893,N_48436,N_47875);
nand UO_894 (O_894,N_49096,N_48049);
xnor UO_895 (O_895,N_47865,N_49617);
nor UO_896 (O_896,N_48238,N_47584);
nand UO_897 (O_897,N_48041,N_47748);
nand UO_898 (O_898,N_48476,N_47558);
nor UO_899 (O_899,N_48922,N_49802);
nand UO_900 (O_900,N_48658,N_48977);
nand UO_901 (O_901,N_48104,N_49989);
or UO_902 (O_902,N_49399,N_48744);
nand UO_903 (O_903,N_47962,N_48472);
nand UO_904 (O_904,N_48228,N_47779);
or UO_905 (O_905,N_48023,N_48785);
nand UO_906 (O_906,N_48914,N_49255);
or UO_907 (O_907,N_49212,N_49056);
nand UO_908 (O_908,N_49446,N_48739);
and UO_909 (O_909,N_47840,N_48637);
and UO_910 (O_910,N_48575,N_49404);
and UO_911 (O_911,N_48251,N_49273);
nand UO_912 (O_912,N_49238,N_49037);
nand UO_913 (O_913,N_48799,N_49577);
nand UO_914 (O_914,N_49564,N_49569);
and UO_915 (O_915,N_48888,N_47838);
or UO_916 (O_916,N_48865,N_49624);
and UO_917 (O_917,N_49413,N_49885);
nand UO_918 (O_918,N_47728,N_48022);
nand UO_919 (O_919,N_48318,N_48444);
or UO_920 (O_920,N_48307,N_47649);
nand UO_921 (O_921,N_49038,N_48109);
xor UO_922 (O_922,N_49594,N_47896);
nand UO_923 (O_923,N_49390,N_48193);
or UO_924 (O_924,N_49926,N_47706);
nor UO_925 (O_925,N_49192,N_47804);
nor UO_926 (O_926,N_47925,N_47532);
nor UO_927 (O_927,N_48893,N_48688);
nand UO_928 (O_928,N_48353,N_48184);
or UO_929 (O_929,N_49891,N_48365);
nor UO_930 (O_930,N_48155,N_48972);
and UO_931 (O_931,N_48231,N_49634);
nor UO_932 (O_932,N_48955,N_48628);
xor UO_933 (O_933,N_49442,N_48286);
or UO_934 (O_934,N_49296,N_48059);
nand UO_935 (O_935,N_49846,N_48800);
or UO_936 (O_936,N_49922,N_49250);
nand UO_937 (O_937,N_48167,N_48723);
or UO_938 (O_938,N_49602,N_48230);
nor UO_939 (O_939,N_49541,N_48080);
or UO_940 (O_940,N_49947,N_47732);
nand UO_941 (O_941,N_48360,N_49694);
and UO_942 (O_942,N_49341,N_49107);
or UO_943 (O_943,N_47720,N_49556);
and UO_944 (O_944,N_47940,N_49372);
xor UO_945 (O_945,N_48794,N_48213);
or UO_946 (O_946,N_49339,N_48731);
and UO_947 (O_947,N_48168,N_47798);
nor UO_948 (O_948,N_49202,N_48350);
nor UO_949 (O_949,N_49605,N_49910);
or UO_950 (O_950,N_49324,N_48125);
xnor UO_951 (O_951,N_48676,N_48620);
and UO_952 (O_952,N_49467,N_49239);
and UO_953 (O_953,N_48567,N_47609);
nand UO_954 (O_954,N_48007,N_48194);
or UO_955 (O_955,N_47766,N_49969);
or UO_956 (O_956,N_49611,N_47628);
xnor UO_957 (O_957,N_47633,N_49519);
xor UO_958 (O_958,N_47848,N_49123);
and UO_959 (O_959,N_49871,N_48205);
nand UO_960 (O_960,N_49325,N_49671);
or UO_961 (O_961,N_49007,N_48210);
and UO_962 (O_962,N_47629,N_47671);
nand UO_963 (O_963,N_48303,N_49300);
and UO_964 (O_964,N_47549,N_48442);
nand UO_965 (O_965,N_49069,N_48598);
nand UO_966 (O_966,N_48534,N_49804);
nor UO_967 (O_967,N_48753,N_48054);
or UO_968 (O_968,N_48283,N_48569);
or UO_969 (O_969,N_49185,N_49455);
or UO_970 (O_970,N_47707,N_48359);
nand UO_971 (O_971,N_48028,N_48349);
nand UO_972 (O_972,N_49231,N_49018);
or UO_973 (O_973,N_47793,N_48139);
nor UO_974 (O_974,N_47976,N_49788);
and UO_975 (O_975,N_47704,N_49918);
nor UO_976 (O_976,N_48807,N_49287);
and UO_977 (O_977,N_48848,N_49094);
nor UO_978 (O_978,N_49074,N_49030);
nand UO_979 (O_979,N_48425,N_47780);
nand UO_980 (O_980,N_49333,N_49875);
xnor UO_981 (O_981,N_48317,N_49241);
or UO_982 (O_982,N_49254,N_47638);
or UO_983 (O_983,N_49189,N_49067);
xor UO_984 (O_984,N_49981,N_47782);
nor UO_985 (O_985,N_49233,N_49979);
xor UO_986 (O_986,N_49147,N_48395);
nand UO_987 (O_987,N_48073,N_48029);
nor UO_988 (O_988,N_49930,N_47718);
nor UO_989 (O_989,N_49461,N_48032);
nor UO_990 (O_990,N_48906,N_49345);
or UO_991 (O_991,N_49414,N_47661);
or UO_992 (O_992,N_47781,N_47517);
nor UO_993 (O_993,N_48484,N_47513);
xnor UO_994 (O_994,N_47563,N_47825);
or UO_995 (O_995,N_48496,N_47787);
nand UO_996 (O_996,N_49702,N_48050);
nand UO_997 (O_997,N_48500,N_48779);
xnor UO_998 (O_998,N_49070,N_48656);
nor UO_999 (O_999,N_49186,N_49046);
nand UO_1000 (O_1000,N_48467,N_48855);
nor UO_1001 (O_1001,N_49834,N_47615);
xor UO_1002 (O_1002,N_48729,N_48482);
nor UO_1003 (O_1003,N_48005,N_49643);
nor UO_1004 (O_1004,N_47500,N_47822);
and UO_1005 (O_1005,N_47954,N_49841);
xor UO_1006 (O_1006,N_48901,N_49725);
nand UO_1007 (O_1007,N_48846,N_49562);
and UO_1008 (O_1008,N_48309,N_49087);
nor UO_1009 (O_1009,N_49956,N_49267);
xor UO_1010 (O_1010,N_48589,N_49904);
nand UO_1011 (O_1011,N_48047,N_48447);
or UO_1012 (O_1012,N_48058,N_47555);
nand UO_1013 (O_1013,N_47632,N_48543);
xor UO_1014 (O_1014,N_47929,N_49505);
or UO_1015 (O_1015,N_48025,N_49723);
and UO_1016 (O_1016,N_49161,N_48971);
nand UO_1017 (O_1017,N_48061,N_47996);
or UO_1018 (O_1018,N_48076,N_49289);
and UO_1019 (O_1019,N_47572,N_47510);
xor UO_1020 (O_1020,N_49965,N_48074);
or UO_1021 (O_1021,N_48736,N_49755);
xor UO_1022 (O_1022,N_49621,N_47898);
xnor UO_1023 (O_1023,N_48666,N_47577);
nand UO_1024 (O_1024,N_48622,N_49977);
xnor UO_1025 (O_1025,N_49008,N_48097);
xor UO_1026 (O_1026,N_49653,N_48831);
and UO_1027 (O_1027,N_47987,N_49618);
and UO_1028 (O_1028,N_47519,N_48473);
and UO_1029 (O_1029,N_49200,N_47669);
xor UO_1030 (O_1030,N_48601,N_48686);
xnor UO_1031 (O_1031,N_48787,N_48221);
or UO_1032 (O_1032,N_49583,N_49881);
xor UO_1033 (O_1033,N_48502,N_49477);
or UO_1034 (O_1034,N_49996,N_48754);
and UO_1035 (O_1035,N_48641,N_47501);
or UO_1036 (O_1036,N_49958,N_48173);
nand UO_1037 (O_1037,N_48810,N_49078);
nand UO_1038 (O_1038,N_48759,N_48158);
or UO_1039 (O_1039,N_47620,N_47586);
nand UO_1040 (O_1040,N_49539,N_49251);
xnor UO_1041 (O_1041,N_49064,N_47888);
xor UO_1042 (O_1042,N_49162,N_48226);
and UO_1043 (O_1043,N_47574,N_47951);
nor UO_1044 (O_1044,N_47536,N_47749);
and UO_1045 (O_1045,N_49854,N_49790);
and UO_1046 (O_1046,N_48940,N_49923);
nor UO_1047 (O_1047,N_48636,N_49081);
xor UO_1048 (O_1048,N_49690,N_49709);
nand UO_1049 (O_1049,N_49836,N_47678);
nor UO_1050 (O_1050,N_47792,N_48057);
or UO_1051 (O_1051,N_47905,N_49561);
nand UO_1052 (O_1052,N_48564,N_48220);
nor UO_1053 (O_1053,N_48079,N_48295);
nor UO_1054 (O_1054,N_48561,N_47533);
nor UO_1055 (O_1055,N_47770,N_47590);
xnor UO_1056 (O_1056,N_48795,N_48248);
nand UO_1057 (O_1057,N_49382,N_49236);
xnor UO_1058 (O_1058,N_48430,N_49814);
nand UO_1059 (O_1059,N_49728,N_48791);
xor UO_1060 (O_1060,N_49188,N_48997);
or UO_1061 (O_1061,N_47850,N_47626);
nand UO_1062 (O_1062,N_49113,N_48629);
or UO_1063 (O_1063,N_47882,N_48198);
and UO_1064 (O_1064,N_49532,N_49937);
or UO_1065 (O_1065,N_48043,N_48098);
nor UO_1066 (O_1066,N_48558,N_48907);
nor UO_1067 (O_1067,N_47697,N_48491);
or UO_1068 (O_1068,N_49259,N_49393);
nor UO_1069 (O_1069,N_48978,N_49639);
nand UO_1070 (O_1070,N_48434,N_47692);
nand UO_1071 (O_1071,N_47966,N_48773);
nor UO_1072 (O_1072,N_47681,N_49348);
and UO_1073 (O_1073,N_47829,N_49579);
xor UO_1074 (O_1074,N_47853,N_48416);
xnor UO_1075 (O_1075,N_48984,N_49940);
nor UO_1076 (O_1076,N_48486,N_48610);
nand UO_1077 (O_1077,N_49798,N_47696);
nor UO_1078 (O_1078,N_49263,N_49950);
and UO_1079 (O_1079,N_49959,N_49336);
xor UO_1080 (O_1080,N_47750,N_49292);
xor UO_1081 (O_1081,N_47993,N_49134);
or UO_1082 (O_1082,N_48928,N_48992);
nand UO_1083 (O_1083,N_49315,N_49705);
xnor UO_1084 (O_1084,N_48612,N_47651);
nor UO_1085 (O_1085,N_47611,N_48990);
and UO_1086 (O_1086,N_48866,N_47915);
nor UO_1087 (O_1087,N_49808,N_49411);
nor UO_1088 (O_1088,N_49436,N_47648);
or UO_1089 (O_1089,N_48517,N_49482);
xnor UO_1090 (O_1090,N_49753,N_49762);
and UO_1091 (O_1091,N_47791,N_48833);
nand UO_1092 (O_1092,N_48229,N_49571);
or UO_1093 (O_1093,N_48121,N_49311);
and UO_1094 (O_1094,N_49772,N_48037);
nor UO_1095 (O_1095,N_49223,N_49552);
and UO_1096 (O_1096,N_48849,N_48954);
and UO_1097 (O_1097,N_48592,N_47736);
and UO_1098 (O_1098,N_49513,N_47643);
nand UO_1099 (O_1099,N_49759,N_47664);
xor UO_1100 (O_1100,N_48376,N_47652);
nor UO_1101 (O_1101,N_49949,N_47660);
and UO_1102 (O_1102,N_48834,N_49403);
and UO_1103 (O_1103,N_48333,N_49902);
xor UO_1104 (O_1104,N_48996,N_48428);
and UO_1105 (O_1105,N_48934,N_48621);
xnor UO_1106 (O_1106,N_49392,N_48000);
nand UO_1107 (O_1107,N_49306,N_48122);
nand UO_1108 (O_1108,N_49351,N_48985);
and UO_1109 (O_1109,N_48822,N_47764);
and UO_1110 (O_1110,N_48207,N_48668);
or UO_1111 (O_1111,N_49899,N_48544);
nand UO_1112 (O_1112,N_47942,N_47939);
nand UO_1113 (O_1113,N_49811,N_49352);
nand UO_1114 (O_1114,N_48227,N_48542);
nor UO_1115 (O_1115,N_48387,N_49771);
xnor UO_1116 (O_1116,N_47686,N_49434);
and UO_1117 (O_1117,N_47631,N_48315);
and UO_1118 (O_1118,N_49817,N_49226);
or UO_1119 (O_1119,N_48571,N_48735);
nand UO_1120 (O_1120,N_49997,N_48002);
and UO_1121 (O_1121,N_48095,N_48045);
and UO_1122 (O_1122,N_49435,N_49204);
xnor UO_1123 (O_1123,N_49124,N_49851);
nand UO_1124 (O_1124,N_49820,N_48143);
nand UO_1125 (O_1125,N_47715,N_48778);
nor UO_1126 (O_1126,N_48875,N_48640);
and UO_1127 (O_1127,N_49726,N_49769);
nor UO_1128 (O_1128,N_48845,N_49972);
or UO_1129 (O_1129,N_48272,N_47603);
xor UO_1130 (O_1130,N_48094,N_48069);
and UO_1131 (O_1131,N_48503,N_49071);
nand UO_1132 (O_1132,N_48819,N_49485);
or UO_1133 (O_1133,N_49437,N_48964);
and UO_1134 (O_1134,N_47917,N_48654);
or UO_1135 (O_1135,N_49397,N_48470);
nor UO_1136 (O_1136,N_47553,N_48255);
or UO_1137 (O_1137,N_48717,N_47961);
nand UO_1138 (O_1138,N_48180,N_47955);
nor UO_1139 (O_1139,N_49495,N_49077);
xnor UO_1140 (O_1140,N_48895,N_49237);
nor UO_1141 (O_1141,N_47772,N_49765);
nor UO_1142 (O_1142,N_48398,N_49553);
nand UO_1143 (O_1143,N_49229,N_49703);
and UO_1144 (O_1144,N_47919,N_49961);
nor UO_1145 (O_1145,N_49211,N_48462);
nand UO_1146 (O_1146,N_48393,N_49915);
xor UO_1147 (O_1147,N_49749,N_49199);
or UO_1148 (O_1148,N_49626,N_47685);
xor UO_1149 (O_1149,N_49641,N_48417);
nor UO_1150 (O_1150,N_48392,N_49095);
and UO_1151 (O_1151,N_49939,N_49112);
and UO_1152 (O_1152,N_49205,N_49265);
nor UO_1153 (O_1153,N_47953,N_47935);
nand UO_1154 (O_1154,N_48936,N_49791);
and UO_1155 (O_1155,N_48300,N_49319);
or UO_1156 (O_1156,N_49451,N_48873);
xor UO_1157 (O_1157,N_48208,N_49252);
or UO_1158 (O_1158,N_47694,N_48863);
or UO_1159 (O_1159,N_48237,N_49966);
or UO_1160 (O_1160,N_48067,N_48945);
nor UO_1161 (O_1161,N_49076,N_48021);
or UO_1162 (O_1162,N_48812,N_49642);
and UO_1163 (O_1163,N_49117,N_47557);
or UO_1164 (O_1164,N_48757,N_49019);
and UO_1165 (O_1165,N_47573,N_48056);
nand UO_1166 (O_1166,N_49490,N_48197);
nor UO_1167 (O_1167,N_48593,N_47851);
nand UO_1168 (O_1168,N_48556,N_48627);
or UO_1169 (O_1169,N_49903,N_49476);
nor UO_1170 (O_1170,N_48813,N_47703);
xor UO_1171 (O_1171,N_49672,N_47994);
nand UO_1172 (O_1172,N_48989,N_48494);
nand UO_1173 (O_1173,N_49717,N_48124);
or UO_1174 (O_1174,N_47534,N_48269);
xnor UO_1175 (O_1175,N_49104,N_49666);
nand UO_1176 (O_1176,N_48956,N_48214);
nand UO_1177 (O_1177,N_48026,N_48950);
xnor UO_1178 (O_1178,N_49088,N_47884);
or UO_1179 (O_1179,N_49120,N_49487);
xor UO_1180 (O_1180,N_49365,N_49133);
or UO_1181 (O_1181,N_49572,N_48684);
nor UO_1182 (O_1182,N_48671,N_49744);
xnor UO_1183 (O_1183,N_48931,N_48479);
xnor UO_1184 (O_1184,N_49953,N_47601);
nand UO_1185 (O_1185,N_49415,N_48638);
and UO_1186 (O_1186,N_49474,N_49366);
or UO_1187 (O_1187,N_49084,N_48113);
xor UO_1188 (O_1188,N_48106,N_47814);
nand UO_1189 (O_1189,N_48347,N_48066);
xor UO_1190 (O_1190,N_47507,N_49305);
xor UO_1191 (O_1191,N_47968,N_47530);
xor UO_1192 (O_1192,N_49812,N_47873);
or UO_1193 (O_1193,N_49974,N_48288);
and UO_1194 (O_1194,N_48506,N_49525);
nor UO_1195 (O_1195,N_49288,N_47846);
and UO_1196 (O_1196,N_49524,N_48582);
and UO_1197 (O_1197,N_47991,N_48414);
nand UO_1198 (O_1198,N_48537,N_48860);
nand UO_1199 (O_1199,N_49176,N_48933);
xor UO_1200 (O_1200,N_49453,N_49815);
or UO_1201 (O_1201,N_49585,N_47795);
or UO_1202 (O_1202,N_49242,N_48626);
xnor UO_1203 (O_1203,N_47591,N_48921);
and UO_1204 (O_1204,N_48072,N_47863);
or UO_1205 (O_1205,N_47807,N_49935);
nand UO_1206 (O_1206,N_49954,N_49066);
or UO_1207 (O_1207,N_48190,N_48044);
or UO_1208 (O_1208,N_49925,N_49210);
nand UO_1209 (O_1209,N_48409,N_49217);
and UO_1210 (O_1210,N_49144,N_49006);
and UO_1211 (O_1211,N_49118,N_49551);
nand UO_1212 (O_1212,N_48216,N_48615);
nand UO_1213 (O_1213,N_47544,N_49085);
or UO_1214 (O_1214,N_48212,N_49187);
and UO_1215 (O_1215,N_47688,N_48319);
or UO_1216 (O_1216,N_48714,N_47866);
nor UO_1217 (O_1217,N_49589,N_47826);
nor UO_1218 (O_1218,N_47790,N_48511);
nand UO_1219 (O_1219,N_48133,N_47606);
nand UO_1220 (O_1220,N_47974,N_48386);
and UO_1221 (O_1221,N_48499,N_47834);
xnor UO_1222 (O_1222,N_47913,N_47808);
xor UO_1223 (O_1223,N_48322,N_49942);
nand UO_1224 (O_1224,N_48563,N_49756);
xnor UO_1225 (O_1225,N_47554,N_47964);
xor UO_1226 (O_1226,N_47721,N_47647);
and UO_1227 (O_1227,N_49523,N_48358);
and UO_1228 (O_1228,N_49636,N_48203);
and UO_1229 (O_1229,N_47837,N_49687);
nand UO_1230 (O_1230,N_49314,N_47705);
xnor UO_1231 (O_1231,N_49612,N_47512);
nand UO_1232 (O_1232,N_47570,N_47503);
xor UO_1233 (O_1233,N_49389,N_49177);
nor UO_1234 (O_1234,N_49864,N_47926);
nand UO_1235 (O_1235,N_48329,N_48842);
nor UO_1236 (O_1236,N_48559,N_49635);
or UO_1237 (O_1237,N_48136,N_48291);
and UO_1238 (O_1238,N_47864,N_49747);
and UO_1239 (O_1239,N_48784,N_47600);
nand UO_1240 (O_1240,N_48894,N_48651);
nor UO_1241 (O_1241,N_47844,N_48843);
and UO_1242 (O_1242,N_47978,N_47921);
nand UO_1243 (O_1243,N_49011,N_49637);
or UO_1244 (O_1244,N_49677,N_48201);
or UO_1245 (O_1245,N_48806,N_49883);
or UO_1246 (O_1246,N_49835,N_47627);
nand UO_1247 (O_1247,N_48093,N_49781);
or UO_1248 (O_1248,N_47719,N_49908);
nor UO_1249 (O_1249,N_47635,N_49907);
xor UO_1250 (O_1250,N_49150,N_49005);
nor UO_1251 (O_1251,N_47955,N_47532);
nor UO_1252 (O_1252,N_48558,N_48125);
xnor UO_1253 (O_1253,N_49047,N_48232);
or UO_1254 (O_1254,N_47580,N_47782);
xor UO_1255 (O_1255,N_47959,N_48248);
nor UO_1256 (O_1256,N_49617,N_48540);
or UO_1257 (O_1257,N_48213,N_47685);
xnor UO_1258 (O_1258,N_49547,N_49417);
nand UO_1259 (O_1259,N_47603,N_48488);
or UO_1260 (O_1260,N_47846,N_49424);
and UO_1261 (O_1261,N_47992,N_47827);
nor UO_1262 (O_1262,N_49741,N_49032);
xor UO_1263 (O_1263,N_47530,N_47652);
or UO_1264 (O_1264,N_48715,N_49308);
or UO_1265 (O_1265,N_48137,N_47895);
and UO_1266 (O_1266,N_48461,N_49659);
xor UO_1267 (O_1267,N_49421,N_49846);
and UO_1268 (O_1268,N_47912,N_49905);
nand UO_1269 (O_1269,N_49690,N_49940);
or UO_1270 (O_1270,N_49980,N_48988);
or UO_1271 (O_1271,N_48387,N_49531);
and UO_1272 (O_1272,N_47551,N_48125);
and UO_1273 (O_1273,N_49971,N_49911);
nor UO_1274 (O_1274,N_47826,N_49619);
or UO_1275 (O_1275,N_49224,N_48077);
nor UO_1276 (O_1276,N_49955,N_47972);
nor UO_1277 (O_1277,N_48577,N_49702);
and UO_1278 (O_1278,N_47532,N_47787);
nor UO_1279 (O_1279,N_48413,N_49930);
or UO_1280 (O_1280,N_49478,N_48563);
nand UO_1281 (O_1281,N_48725,N_48903);
and UO_1282 (O_1282,N_48370,N_49210);
or UO_1283 (O_1283,N_47700,N_48515);
and UO_1284 (O_1284,N_49697,N_48509);
xnor UO_1285 (O_1285,N_47818,N_49156);
nor UO_1286 (O_1286,N_48906,N_49382);
or UO_1287 (O_1287,N_48969,N_48826);
xnor UO_1288 (O_1288,N_48257,N_48761);
and UO_1289 (O_1289,N_47529,N_47719);
and UO_1290 (O_1290,N_48855,N_48546);
xor UO_1291 (O_1291,N_48852,N_47902);
nor UO_1292 (O_1292,N_48677,N_49806);
nand UO_1293 (O_1293,N_49297,N_49098);
or UO_1294 (O_1294,N_47658,N_49071);
or UO_1295 (O_1295,N_48995,N_49057);
xnor UO_1296 (O_1296,N_49655,N_48265);
nor UO_1297 (O_1297,N_49423,N_49246);
or UO_1298 (O_1298,N_49798,N_47857);
xor UO_1299 (O_1299,N_47870,N_48239);
nor UO_1300 (O_1300,N_48372,N_48645);
and UO_1301 (O_1301,N_49782,N_47568);
or UO_1302 (O_1302,N_49963,N_49962);
xor UO_1303 (O_1303,N_49589,N_47864);
nand UO_1304 (O_1304,N_48946,N_48257);
nor UO_1305 (O_1305,N_48102,N_47782);
nand UO_1306 (O_1306,N_49786,N_48714);
or UO_1307 (O_1307,N_49339,N_48126);
or UO_1308 (O_1308,N_49895,N_49468);
nand UO_1309 (O_1309,N_49228,N_49576);
nor UO_1310 (O_1310,N_47653,N_49558);
or UO_1311 (O_1311,N_48876,N_47607);
nand UO_1312 (O_1312,N_49335,N_48960);
nand UO_1313 (O_1313,N_48470,N_49327);
nand UO_1314 (O_1314,N_49747,N_48976);
or UO_1315 (O_1315,N_49374,N_47505);
or UO_1316 (O_1316,N_49037,N_49213);
and UO_1317 (O_1317,N_48203,N_49743);
or UO_1318 (O_1318,N_49665,N_49195);
xor UO_1319 (O_1319,N_48730,N_48217);
xor UO_1320 (O_1320,N_49092,N_49568);
xnor UO_1321 (O_1321,N_49343,N_47994);
and UO_1322 (O_1322,N_48503,N_49179);
xnor UO_1323 (O_1323,N_48080,N_49477);
or UO_1324 (O_1324,N_49670,N_49761);
nor UO_1325 (O_1325,N_48197,N_48347);
nor UO_1326 (O_1326,N_49106,N_49447);
xnor UO_1327 (O_1327,N_47535,N_48233);
or UO_1328 (O_1328,N_48075,N_48847);
nand UO_1329 (O_1329,N_49784,N_48856);
nand UO_1330 (O_1330,N_49792,N_49225);
xnor UO_1331 (O_1331,N_48639,N_48048);
nand UO_1332 (O_1332,N_47733,N_49727);
xor UO_1333 (O_1333,N_48120,N_48977);
or UO_1334 (O_1334,N_48676,N_47934);
nand UO_1335 (O_1335,N_48786,N_49621);
or UO_1336 (O_1336,N_48002,N_47801);
xnor UO_1337 (O_1337,N_49419,N_47973);
nor UO_1338 (O_1338,N_48608,N_48941);
xor UO_1339 (O_1339,N_49346,N_48741);
xnor UO_1340 (O_1340,N_49566,N_47707);
and UO_1341 (O_1341,N_48053,N_48103);
xnor UO_1342 (O_1342,N_48522,N_49911);
or UO_1343 (O_1343,N_49150,N_48480);
and UO_1344 (O_1344,N_48230,N_48136);
nor UO_1345 (O_1345,N_47604,N_49588);
or UO_1346 (O_1346,N_49499,N_48619);
and UO_1347 (O_1347,N_49496,N_49527);
xor UO_1348 (O_1348,N_49527,N_49729);
xnor UO_1349 (O_1349,N_48278,N_49216);
or UO_1350 (O_1350,N_48139,N_49153);
nor UO_1351 (O_1351,N_48972,N_47811);
nand UO_1352 (O_1352,N_47533,N_49745);
or UO_1353 (O_1353,N_48660,N_48534);
or UO_1354 (O_1354,N_49076,N_48515);
nand UO_1355 (O_1355,N_48797,N_49302);
xnor UO_1356 (O_1356,N_47989,N_49593);
or UO_1357 (O_1357,N_48780,N_49559);
and UO_1358 (O_1358,N_48479,N_48035);
or UO_1359 (O_1359,N_48808,N_49195);
xor UO_1360 (O_1360,N_48795,N_49372);
and UO_1361 (O_1361,N_49573,N_48984);
and UO_1362 (O_1362,N_48592,N_48439);
and UO_1363 (O_1363,N_48369,N_48941);
nor UO_1364 (O_1364,N_49862,N_47748);
nand UO_1365 (O_1365,N_49352,N_49570);
nor UO_1366 (O_1366,N_49846,N_47955);
or UO_1367 (O_1367,N_49356,N_49123);
nand UO_1368 (O_1368,N_47978,N_48648);
xnor UO_1369 (O_1369,N_48985,N_48380);
xnor UO_1370 (O_1370,N_49185,N_48117);
nand UO_1371 (O_1371,N_48293,N_48376);
and UO_1372 (O_1372,N_49271,N_49979);
xnor UO_1373 (O_1373,N_49589,N_49107);
nand UO_1374 (O_1374,N_48201,N_47655);
nor UO_1375 (O_1375,N_48752,N_49497);
and UO_1376 (O_1376,N_48780,N_48770);
nand UO_1377 (O_1377,N_49290,N_49939);
nand UO_1378 (O_1378,N_48186,N_49956);
and UO_1379 (O_1379,N_48937,N_49396);
nand UO_1380 (O_1380,N_49867,N_49527);
xor UO_1381 (O_1381,N_48059,N_47567);
or UO_1382 (O_1382,N_49177,N_48607);
xnor UO_1383 (O_1383,N_48391,N_48191);
or UO_1384 (O_1384,N_48920,N_48056);
or UO_1385 (O_1385,N_48596,N_49327);
xnor UO_1386 (O_1386,N_49187,N_49823);
and UO_1387 (O_1387,N_48005,N_48490);
nor UO_1388 (O_1388,N_49184,N_48877);
or UO_1389 (O_1389,N_48103,N_49132);
or UO_1390 (O_1390,N_49920,N_49714);
xnor UO_1391 (O_1391,N_48327,N_47866);
xor UO_1392 (O_1392,N_47979,N_49281);
nor UO_1393 (O_1393,N_49979,N_48042);
xnor UO_1394 (O_1394,N_49595,N_48413);
or UO_1395 (O_1395,N_49209,N_49705);
and UO_1396 (O_1396,N_49057,N_48045);
xor UO_1397 (O_1397,N_48900,N_48955);
nor UO_1398 (O_1398,N_48575,N_48493);
nand UO_1399 (O_1399,N_48624,N_47582);
or UO_1400 (O_1400,N_49443,N_48187);
xor UO_1401 (O_1401,N_49452,N_49922);
nand UO_1402 (O_1402,N_49763,N_49977);
nand UO_1403 (O_1403,N_48187,N_49831);
or UO_1404 (O_1404,N_48302,N_48740);
nand UO_1405 (O_1405,N_49387,N_49866);
or UO_1406 (O_1406,N_49162,N_48737);
nor UO_1407 (O_1407,N_48396,N_48891);
and UO_1408 (O_1408,N_47678,N_49489);
or UO_1409 (O_1409,N_49542,N_48317);
nor UO_1410 (O_1410,N_48343,N_49839);
xnor UO_1411 (O_1411,N_49943,N_47572);
nand UO_1412 (O_1412,N_48710,N_48016);
or UO_1413 (O_1413,N_49081,N_49918);
or UO_1414 (O_1414,N_47955,N_48679);
or UO_1415 (O_1415,N_48508,N_47999);
nand UO_1416 (O_1416,N_49151,N_47788);
or UO_1417 (O_1417,N_48833,N_47581);
nand UO_1418 (O_1418,N_49229,N_48192);
and UO_1419 (O_1419,N_49300,N_48240);
and UO_1420 (O_1420,N_49130,N_48905);
nand UO_1421 (O_1421,N_47697,N_49143);
and UO_1422 (O_1422,N_49058,N_49485);
and UO_1423 (O_1423,N_49682,N_49283);
nand UO_1424 (O_1424,N_49923,N_49036);
xor UO_1425 (O_1425,N_49781,N_48205);
nand UO_1426 (O_1426,N_49499,N_48267);
xor UO_1427 (O_1427,N_47903,N_49252);
nor UO_1428 (O_1428,N_47584,N_48698);
nand UO_1429 (O_1429,N_47522,N_47923);
or UO_1430 (O_1430,N_47964,N_48155);
and UO_1431 (O_1431,N_48002,N_47570);
nand UO_1432 (O_1432,N_49067,N_48015);
and UO_1433 (O_1433,N_49611,N_49830);
or UO_1434 (O_1434,N_48048,N_48587);
nand UO_1435 (O_1435,N_48676,N_48456);
or UO_1436 (O_1436,N_49490,N_47575);
nor UO_1437 (O_1437,N_47661,N_49862);
and UO_1438 (O_1438,N_48470,N_49515);
nand UO_1439 (O_1439,N_48604,N_47628);
nor UO_1440 (O_1440,N_48437,N_48296);
nand UO_1441 (O_1441,N_49187,N_48161);
nor UO_1442 (O_1442,N_48672,N_47912);
xnor UO_1443 (O_1443,N_49135,N_49894);
nand UO_1444 (O_1444,N_48281,N_48123);
or UO_1445 (O_1445,N_49320,N_47960);
nor UO_1446 (O_1446,N_48269,N_48762);
and UO_1447 (O_1447,N_48521,N_49772);
xor UO_1448 (O_1448,N_48911,N_49885);
and UO_1449 (O_1449,N_47917,N_49752);
xor UO_1450 (O_1450,N_49131,N_48955);
xor UO_1451 (O_1451,N_48243,N_49094);
nor UO_1452 (O_1452,N_48692,N_48107);
or UO_1453 (O_1453,N_49051,N_49029);
nor UO_1454 (O_1454,N_47613,N_48484);
xnor UO_1455 (O_1455,N_48171,N_47746);
xnor UO_1456 (O_1456,N_49281,N_47821);
and UO_1457 (O_1457,N_48440,N_48208);
nor UO_1458 (O_1458,N_47616,N_48266);
or UO_1459 (O_1459,N_49629,N_47602);
nand UO_1460 (O_1460,N_49791,N_48783);
or UO_1461 (O_1461,N_49709,N_49457);
nor UO_1462 (O_1462,N_48898,N_49473);
xnor UO_1463 (O_1463,N_49286,N_48234);
xor UO_1464 (O_1464,N_49251,N_48565);
and UO_1465 (O_1465,N_49792,N_48404);
nand UO_1466 (O_1466,N_48370,N_47871);
and UO_1467 (O_1467,N_48525,N_49773);
xor UO_1468 (O_1468,N_49192,N_49274);
or UO_1469 (O_1469,N_48170,N_49611);
or UO_1470 (O_1470,N_49580,N_49134);
or UO_1471 (O_1471,N_49121,N_49947);
xnor UO_1472 (O_1472,N_49251,N_49200);
and UO_1473 (O_1473,N_47764,N_48528);
or UO_1474 (O_1474,N_47692,N_47618);
or UO_1475 (O_1475,N_49264,N_48652);
or UO_1476 (O_1476,N_49014,N_48441);
nor UO_1477 (O_1477,N_48526,N_47577);
nand UO_1478 (O_1478,N_47887,N_47892);
xnor UO_1479 (O_1479,N_47514,N_48427);
nand UO_1480 (O_1480,N_48038,N_47864);
nand UO_1481 (O_1481,N_48122,N_47724);
and UO_1482 (O_1482,N_49947,N_48828);
xnor UO_1483 (O_1483,N_47736,N_48022);
nand UO_1484 (O_1484,N_49561,N_49833);
or UO_1485 (O_1485,N_49289,N_49060);
nor UO_1486 (O_1486,N_49007,N_49293);
nor UO_1487 (O_1487,N_49406,N_49179);
and UO_1488 (O_1488,N_47506,N_48315);
nor UO_1489 (O_1489,N_49179,N_48777);
and UO_1490 (O_1490,N_49537,N_49651);
or UO_1491 (O_1491,N_48771,N_49093);
nor UO_1492 (O_1492,N_49966,N_49427);
xor UO_1493 (O_1493,N_48053,N_49984);
or UO_1494 (O_1494,N_48121,N_49178);
xor UO_1495 (O_1495,N_47671,N_47815);
xor UO_1496 (O_1496,N_49111,N_48796);
or UO_1497 (O_1497,N_49857,N_48926);
xor UO_1498 (O_1498,N_48673,N_49896);
nor UO_1499 (O_1499,N_49829,N_47546);
and UO_1500 (O_1500,N_49138,N_48750);
xor UO_1501 (O_1501,N_47921,N_47938);
nor UO_1502 (O_1502,N_49189,N_49738);
xnor UO_1503 (O_1503,N_48286,N_48054);
nand UO_1504 (O_1504,N_49057,N_48117);
or UO_1505 (O_1505,N_48234,N_48070);
or UO_1506 (O_1506,N_48918,N_47687);
nand UO_1507 (O_1507,N_49279,N_48033);
xnor UO_1508 (O_1508,N_48931,N_48504);
and UO_1509 (O_1509,N_49721,N_49537);
and UO_1510 (O_1510,N_49764,N_49478);
xnor UO_1511 (O_1511,N_48031,N_48105);
or UO_1512 (O_1512,N_48968,N_49398);
nand UO_1513 (O_1513,N_48113,N_49597);
nor UO_1514 (O_1514,N_48415,N_48416);
and UO_1515 (O_1515,N_47913,N_49164);
nand UO_1516 (O_1516,N_48944,N_47741);
nand UO_1517 (O_1517,N_48578,N_48470);
xor UO_1518 (O_1518,N_48878,N_49747);
xor UO_1519 (O_1519,N_48267,N_47714);
nor UO_1520 (O_1520,N_47954,N_49830);
and UO_1521 (O_1521,N_48365,N_49231);
nand UO_1522 (O_1522,N_48581,N_47963);
or UO_1523 (O_1523,N_48482,N_48117);
nor UO_1524 (O_1524,N_48194,N_48144);
xnor UO_1525 (O_1525,N_48562,N_49657);
xnor UO_1526 (O_1526,N_47500,N_49404);
and UO_1527 (O_1527,N_49239,N_47838);
or UO_1528 (O_1528,N_49588,N_49272);
nand UO_1529 (O_1529,N_48801,N_49689);
nand UO_1530 (O_1530,N_47875,N_48298);
or UO_1531 (O_1531,N_48911,N_47978);
nor UO_1532 (O_1532,N_49533,N_47665);
nor UO_1533 (O_1533,N_49711,N_47672);
or UO_1534 (O_1534,N_48741,N_49646);
xor UO_1535 (O_1535,N_48215,N_47881);
nor UO_1536 (O_1536,N_47713,N_47693);
or UO_1537 (O_1537,N_48390,N_48956);
nand UO_1538 (O_1538,N_49553,N_48861);
nor UO_1539 (O_1539,N_48920,N_47596);
and UO_1540 (O_1540,N_49119,N_49893);
nor UO_1541 (O_1541,N_47894,N_47966);
xnor UO_1542 (O_1542,N_48017,N_48927);
nor UO_1543 (O_1543,N_49111,N_49431);
or UO_1544 (O_1544,N_49675,N_48196);
nand UO_1545 (O_1545,N_49757,N_49779);
or UO_1546 (O_1546,N_48483,N_47772);
nand UO_1547 (O_1547,N_47712,N_48069);
nor UO_1548 (O_1548,N_49544,N_49137);
nand UO_1549 (O_1549,N_47882,N_47616);
or UO_1550 (O_1550,N_47874,N_49236);
and UO_1551 (O_1551,N_47944,N_49479);
xor UO_1552 (O_1552,N_47760,N_49617);
nor UO_1553 (O_1553,N_47882,N_49257);
xor UO_1554 (O_1554,N_49470,N_49938);
nor UO_1555 (O_1555,N_48442,N_47612);
xor UO_1556 (O_1556,N_49097,N_48359);
or UO_1557 (O_1557,N_49677,N_47967);
xor UO_1558 (O_1558,N_49453,N_49440);
nand UO_1559 (O_1559,N_49586,N_47601);
nor UO_1560 (O_1560,N_49565,N_49268);
or UO_1561 (O_1561,N_49255,N_49458);
and UO_1562 (O_1562,N_49344,N_47512);
nor UO_1563 (O_1563,N_47690,N_49711);
and UO_1564 (O_1564,N_48507,N_47906);
and UO_1565 (O_1565,N_49647,N_49139);
and UO_1566 (O_1566,N_49451,N_48438);
xnor UO_1567 (O_1567,N_48441,N_49989);
nor UO_1568 (O_1568,N_48614,N_48149);
or UO_1569 (O_1569,N_48717,N_49970);
xor UO_1570 (O_1570,N_48317,N_48365);
nand UO_1571 (O_1571,N_47913,N_47856);
and UO_1572 (O_1572,N_48128,N_47956);
and UO_1573 (O_1573,N_49266,N_49394);
xnor UO_1574 (O_1574,N_48039,N_48710);
nor UO_1575 (O_1575,N_47880,N_48388);
xor UO_1576 (O_1576,N_49804,N_48891);
nand UO_1577 (O_1577,N_47796,N_48214);
and UO_1578 (O_1578,N_48060,N_47751);
or UO_1579 (O_1579,N_48059,N_49432);
nor UO_1580 (O_1580,N_47709,N_49582);
xnor UO_1581 (O_1581,N_49621,N_48870);
nand UO_1582 (O_1582,N_47700,N_49237);
and UO_1583 (O_1583,N_48441,N_47955);
nor UO_1584 (O_1584,N_48725,N_49025);
nor UO_1585 (O_1585,N_48403,N_47684);
or UO_1586 (O_1586,N_49607,N_47508);
or UO_1587 (O_1587,N_49506,N_48584);
nand UO_1588 (O_1588,N_47830,N_49624);
nand UO_1589 (O_1589,N_48217,N_49734);
and UO_1590 (O_1590,N_47554,N_48902);
and UO_1591 (O_1591,N_47523,N_48942);
nand UO_1592 (O_1592,N_49940,N_47786);
xor UO_1593 (O_1593,N_48187,N_49772);
xnor UO_1594 (O_1594,N_49603,N_48401);
xnor UO_1595 (O_1595,N_49375,N_49384);
nand UO_1596 (O_1596,N_49093,N_47888);
xor UO_1597 (O_1597,N_48511,N_49072);
nand UO_1598 (O_1598,N_47636,N_49249);
and UO_1599 (O_1599,N_47788,N_47602);
nor UO_1600 (O_1600,N_48420,N_49283);
xnor UO_1601 (O_1601,N_47847,N_48262);
or UO_1602 (O_1602,N_49044,N_49592);
xnor UO_1603 (O_1603,N_48605,N_49251);
and UO_1604 (O_1604,N_47791,N_47790);
or UO_1605 (O_1605,N_49713,N_48936);
or UO_1606 (O_1606,N_48644,N_49233);
or UO_1607 (O_1607,N_49608,N_49389);
nor UO_1608 (O_1608,N_48785,N_48611);
xor UO_1609 (O_1609,N_48983,N_48234);
nor UO_1610 (O_1610,N_49519,N_47787);
or UO_1611 (O_1611,N_48993,N_47825);
xor UO_1612 (O_1612,N_49350,N_48145);
nand UO_1613 (O_1613,N_48405,N_49127);
nor UO_1614 (O_1614,N_48499,N_49002);
and UO_1615 (O_1615,N_49540,N_49108);
nand UO_1616 (O_1616,N_47775,N_49524);
nor UO_1617 (O_1617,N_48140,N_49297);
xor UO_1618 (O_1618,N_49206,N_49453);
nor UO_1619 (O_1619,N_48247,N_48355);
nand UO_1620 (O_1620,N_48440,N_49210);
and UO_1621 (O_1621,N_49494,N_49222);
nor UO_1622 (O_1622,N_48150,N_49930);
and UO_1623 (O_1623,N_47715,N_48446);
or UO_1624 (O_1624,N_49004,N_48592);
and UO_1625 (O_1625,N_49151,N_47909);
nand UO_1626 (O_1626,N_49917,N_47825);
nor UO_1627 (O_1627,N_48497,N_49616);
xnor UO_1628 (O_1628,N_47636,N_47656);
xor UO_1629 (O_1629,N_49738,N_48618);
nand UO_1630 (O_1630,N_49355,N_48975);
and UO_1631 (O_1631,N_47534,N_49699);
nand UO_1632 (O_1632,N_48354,N_49606);
xor UO_1633 (O_1633,N_48485,N_49018);
nor UO_1634 (O_1634,N_49339,N_47538);
xor UO_1635 (O_1635,N_47783,N_48977);
and UO_1636 (O_1636,N_48896,N_48266);
nand UO_1637 (O_1637,N_49289,N_49032);
nor UO_1638 (O_1638,N_49792,N_48438);
and UO_1639 (O_1639,N_47720,N_48796);
and UO_1640 (O_1640,N_49612,N_49565);
xor UO_1641 (O_1641,N_49806,N_49308);
xnor UO_1642 (O_1642,N_48027,N_49196);
nor UO_1643 (O_1643,N_48325,N_48729);
nand UO_1644 (O_1644,N_47628,N_49696);
xnor UO_1645 (O_1645,N_49455,N_47568);
nor UO_1646 (O_1646,N_49455,N_49784);
or UO_1647 (O_1647,N_49190,N_47761);
or UO_1648 (O_1648,N_48786,N_49372);
and UO_1649 (O_1649,N_47565,N_49401);
or UO_1650 (O_1650,N_48347,N_49503);
or UO_1651 (O_1651,N_48932,N_47620);
xnor UO_1652 (O_1652,N_48518,N_49146);
or UO_1653 (O_1653,N_49429,N_49959);
or UO_1654 (O_1654,N_49572,N_48672);
xnor UO_1655 (O_1655,N_48643,N_49336);
xor UO_1656 (O_1656,N_47855,N_48675);
nor UO_1657 (O_1657,N_49725,N_49932);
nor UO_1658 (O_1658,N_49042,N_48886);
or UO_1659 (O_1659,N_48631,N_48265);
xnor UO_1660 (O_1660,N_47714,N_49919);
nor UO_1661 (O_1661,N_48508,N_47776);
and UO_1662 (O_1662,N_49852,N_47688);
nor UO_1663 (O_1663,N_47910,N_48619);
nor UO_1664 (O_1664,N_49417,N_48417);
xnor UO_1665 (O_1665,N_48451,N_49572);
nor UO_1666 (O_1666,N_49542,N_48723);
nor UO_1667 (O_1667,N_47666,N_47663);
or UO_1668 (O_1668,N_48176,N_49071);
nor UO_1669 (O_1669,N_48798,N_49270);
nand UO_1670 (O_1670,N_49822,N_47904);
nand UO_1671 (O_1671,N_48863,N_49204);
xor UO_1672 (O_1672,N_49116,N_49254);
and UO_1673 (O_1673,N_48061,N_47867);
and UO_1674 (O_1674,N_48281,N_48826);
and UO_1675 (O_1675,N_48729,N_49641);
or UO_1676 (O_1676,N_47780,N_49063);
nand UO_1677 (O_1677,N_47687,N_48578);
or UO_1678 (O_1678,N_47970,N_48361);
or UO_1679 (O_1679,N_49220,N_49336);
xnor UO_1680 (O_1680,N_47601,N_49396);
nor UO_1681 (O_1681,N_48979,N_47906);
nand UO_1682 (O_1682,N_47690,N_47540);
and UO_1683 (O_1683,N_48388,N_48344);
and UO_1684 (O_1684,N_48943,N_47578);
nand UO_1685 (O_1685,N_48847,N_47990);
nor UO_1686 (O_1686,N_47688,N_47746);
or UO_1687 (O_1687,N_49303,N_49802);
nor UO_1688 (O_1688,N_49314,N_48878);
nand UO_1689 (O_1689,N_47857,N_49290);
and UO_1690 (O_1690,N_49197,N_49416);
xnor UO_1691 (O_1691,N_48917,N_48379);
xnor UO_1692 (O_1692,N_49828,N_48871);
or UO_1693 (O_1693,N_48720,N_48173);
xnor UO_1694 (O_1694,N_49340,N_48126);
or UO_1695 (O_1695,N_47778,N_48797);
nor UO_1696 (O_1696,N_48862,N_48920);
or UO_1697 (O_1697,N_48294,N_49498);
and UO_1698 (O_1698,N_48240,N_49269);
and UO_1699 (O_1699,N_49772,N_47875);
or UO_1700 (O_1700,N_49159,N_49104);
or UO_1701 (O_1701,N_47997,N_49661);
and UO_1702 (O_1702,N_49957,N_47744);
and UO_1703 (O_1703,N_49523,N_48156);
or UO_1704 (O_1704,N_47864,N_48367);
nand UO_1705 (O_1705,N_47713,N_48982);
and UO_1706 (O_1706,N_49409,N_48269);
nand UO_1707 (O_1707,N_49608,N_49490);
nor UO_1708 (O_1708,N_48979,N_49159);
nor UO_1709 (O_1709,N_49009,N_47534);
nor UO_1710 (O_1710,N_49887,N_48452);
and UO_1711 (O_1711,N_48239,N_47505);
xnor UO_1712 (O_1712,N_48974,N_47564);
nand UO_1713 (O_1713,N_48343,N_48000);
xor UO_1714 (O_1714,N_49546,N_48774);
and UO_1715 (O_1715,N_48444,N_49174);
and UO_1716 (O_1716,N_47935,N_48371);
nand UO_1717 (O_1717,N_47869,N_48255);
xor UO_1718 (O_1718,N_47868,N_47599);
nand UO_1719 (O_1719,N_47506,N_48314);
and UO_1720 (O_1720,N_47774,N_48466);
xor UO_1721 (O_1721,N_49441,N_48020);
nor UO_1722 (O_1722,N_48786,N_48413);
nand UO_1723 (O_1723,N_48419,N_49694);
or UO_1724 (O_1724,N_48256,N_48077);
nand UO_1725 (O_1725,N_48254,N_48753);
and UO_1726 (O_1726,N_49709,N_49517);
xnor UO_1727 (O_1727,N_48738,N_48163);
xnor UO_1728 (O_1728,N_48465,N_49241);
xnor UO_1729 (O_1729,N_49205,N_49315);
nor UO_1730 (O_1730,N_47629,N_49105);
or UO_1731 (O_1731,N_49958,N_48571);
and UO_1732 (O_1732,N_47728,N_48636);
or UO_1733 (O_1733,N_48108,N_49800);
nand UO_1734 (O_1734,N_49685,N_49340);
and UO_1735 (O_1735,N_47926,N_47937);
and UO_1736 (O_1736,N_49413,N_49263);
or UO_1737 (O_1737,N_49571,N_49093);
or UO_1738 (O_1738,N_48893,N_48722);
nand UO_1739 (O_1739,N_48014,N_49689);
and UO_1740 (O_1740,N_48959,N_49770);
xor UO_1741 (O_1741,N_49488,N_47655);
or UO_1742 (O_1742,N_47657,N_49458);
nor UO_1743 (O_1743,N_48318,N_49993);
nor UO_1744 (O_1744,N_48564,N_48725);
and UO_1745 (O_1745,N_48123,N_47985);
nor UO_1746 (O_1746,N_49554,N_49736);
and UO_1747 (O_1747,N_49138,N_48970);
and UO_1748 (O_1748,N_47946,N_48072);
or UO_1749 (O_1749,N_48985,N_48134);
xnor UO_1750 (O_1750,N_48989,N_48025);
and UO_1751 (O_1751,N_49536,N_49124);
nand UO_1752 (O_1752,N_49472,N_47886);
nand UO_1753 (O_1753,N_49366,N_48652);
nor UO_1754 (O_1754,N_49454,N_49373);
nor UO_1755 (O_1755,N_49405,N_48340);
nor UO_1756 (O_1756,N_48084,N_48500);
xnor UO_1757 (O_1757,N_48081,N_49366);
and UO_1758 (O_1758,N_48793,N_49918);
or UO_1759 (O_1759,N_49609,N_48254);
and UO_1760 (O_1760,N_48167,N_47874);
xnor UO_1761 (O_1761,N_47525,N_47529);
or UO_1762 (O_1762,N_48047,N_48860);
or UO_1763 (O_1763,N_47786,N_47635);
nand UO_1764 (O_1764,N_49419,N_49990);
xor UO_1765 (O_1765,N_49033,N_48917);
nand UO_1766 (O_1766,N_48268,N_48003);
and UO_1767 (O_1767,N_47571,N_48798);
xnor UO_1768 (O_1768,N_48700,N_48633);
nand UO_1769 (O_1769,N_48018,N_48729);
and UO_1770 (O_1770,N_48490,N_48726);
xnor UO_1771 (O_1771,N_48110,N_48558);
xor UO_1772 (O_1772,N_47581,N_47828);
nor UO_1773 (O_1773,N_49370,N_49157);
xor UO_1774 (O_1774,N_49438,N_48902);
xor UO_1775 (O_1775,N_48426,N_49394);
and UO_1776 (O_1776,N_48785,N_49351);
nand UO_1777 (O_1777,N_49589,N_48877);
xnor UO_1778 (O_1778,N_48501,N_47678);
nor UO_1779 (O_1779,N_48018,N_49118);
nor UO_1780 (O_1780,N_49000,N_47745);
nor UO_1781 (O_1781,N_49051,N_48719);
nor UO_1782 (O_1782,N_49206,N_49824);
and UO_1783 (O_1783,N_48200,N_47589);
nand UO_1784 (O_1784,N_48208,N_49384);
and UO_1785 (O_1785,N_47849,N_49985);
xor UO_1786 (O_1786,N_47973,N_49001);
nand UO_1787 (O_1787,N_49911,N_49906);
xnor UO_1788 (O_1788,N_47718,N_48273);
nor UO_1789 (O_1789,N_48574,N_49938);
xor UO_1790 (O_1790,N_49919,N_49972);
xnor UO_1791 (O_1791,N_49602,N_49556);
or UO_1792 (O_1792,N_47502,N_47922);
or UO_1793 (O_1793,N_49688,N_49010);
or UO_1794 (O_1794,N_48896,N_49115);
nand UO_1795 (O_1795,N_47997,N_47976);
or UO_1796 (O_1796,N_49948,N_47978);
nor UO_1797 (O_1797,N_47585,N_47911);
nand UO_1798 (O_1798,N_48969,N_48393);
xor UO_1799 (O_1799,N_48078,N_49919);
and UO_1800 (O_1800,N_48658,N_49014);
or UO_1801 (O_1801,N_48601,N_48524);
or UO_1802 (O_1802,N_48129,N_47815);
nor UO_1803 (O_1803,N_48189,N_48131);
and UO_1804 (O_1804,N_48234,N_49856);
nor UO_1805 (O_1805,N_49786,N_49928);
nor UO_1806 (O_1806,N_49089,N_48992);
xor UO_1807 (O_1807,N_48981,N_49013);
nor UO_1808 (O_1808,N_48058,N_49480);
xor UO_1809 (O_1809,N_48309,N_47847);
nor UO_1810 (O_1810,N_48867,N_48245);
nor UO_1811 (O_1811,N_48707,N_48163);
nor UO_1812 (O_1812,N_48581,N_48922);
or UO_1813 (O_1813,N_49780,N_47577);
xnor UO_1814 (O_1814,N_49585,N_49901);
or UO_1815 (O_1815,N_49400,N_49633);
xor UO_1816 (O_1816,N_49579,N_47776);
and UO_1817 (O_1817,N_48267,N_48765);
nor UO_1818 (O_1818,N_49613,N_49845);
and UO_1819 (O_1819,N_48513,N_49106);
nand UO_1820 (O_1820,N_48479,N_48895);
and UO_1821 (O_1821,N_49356,N_48220);
nor UO_1822 (O_1822,N_47945,N_49703);
xor UO_1823 (O_1823,N_49289,N_49393);
nand UO_1824 (O_1824,N_47737,N_47750);
nand UO_1825 (O_1825,N_49023,N_47533);
and UO_1826 (O_1826,N_49507,N_48388);
nand UO_1827 (O_1827,N_48672,N_48739);
xor UO_1828 (O_1828,N_49986,N_49572);
and UO_1829 (O_1829,N_48965,N_49041);
nand UO_1830 (O_1830,N_48642,N_49676);
nor UO_1831 (O_1831,N_48738,N_49753);
nand UO_1832 (O_1832,N_49196,N_49671);
nor UO_1833 (O_1833,N_48177,N_49801);
nand UO_1834 (O_1834,N_49218,N_48964);
or UO_1835 (O_1835,N_48054,N_47794);
nor UO_1836 (O_1836,N_48139,N_49647);
xor UO_1837 (O_1837,N_49312,N_47535);
xnor UO_1838 (O_1838,N_49155,N_48191);
xnor UO_1839 (O_1839,N_48635,N_48853);
nor UO_1840 (O_1840,N_49127,N_47591);
and UO_1841 (O_1841,N_49614,N_47736);
and UO_1842 (O_1842,N_48786,N_47766);
or UO_1843 (O_1843,N_49019,N_49792);
nor UO_1844 (O_1844,N_48014,N_48198);
nand UO_1845 (O_1845,N_47648,N_48620);
and UO_1846 (O_1846,N_48415,N_48201);
xnor UO_1847 (O_1847,N_48085,N_49622);
and UO_1848 (O_1848,N_49656,N_48901);
or UO_1849 (O_1849,N_48565,N_48678);
nand UO_1850 (O_1850,N_47777,N_48610);
or UO_1851 (O_1851,N_48179,N_49765);
nor UO_1852 (O_1852,N_49007,N_48598);
nor UO_1853 (O_1853,N_48996,N_49707);
and UO_1854 (O_1854,N_49557,N_48460);
nor UO_1855 (O_1855,N_48363,N_47958);
or UO_1856 (O_1856,N_47956,N_49330);
nand UO_1857 (O_1857,N_48232,N_49351);
or UO_1858 (O_1858,N_49276,N_49965);
and UO_1859 (O_1859,N_48223,N_48496);
nand UO_1860 (O_1860,N_47588,N_47514);
xor UO_1861 (O_1861,N_49844,N_48324);
nor UO_1862 (O_1862,N_47899,N_47838);
nand UO_1863 (O_1863,N_48823,N_48832);
xor UO_1864 (O_1864,N_49862,N_48412);
xnor UO_1865 (O_1865,N_48693,N_47715);
and UO_1866 (O_1866,N_49301,N_49551);
xnor UO_1867 (O_1867,N_49571,N_48107);
nand UO_1868 (O_1868,N_48474,N_48176);
nor UO_1869 (O_1869,N_49164,N_49076);
and UO_1870 (O_1870,N_48681,N_47769);
nand UO_1871 (O_1871,N_49386,N_47945);
and UO_1872 (O_1872,N_48807,N_48017);
nor UO_1873 (O_1873,N_48346,N_48459);
or UO_1874 (O_1874,N_49356,N_48676);
xor UO_1875 (O_1875,N_49868,N_47621);
or UO_1876 (O_1876,N_47807,N_48379);
nor UO_1877 (O_1877,N_48827,N_48247);
and UO_1878 (O_1878,N_47500,N_48396);
nand UO_1879 (O_1879,N_47878,N_48781);
nand UO_1880 (O_1880,N_48550,N_47675);
and UO_1881 (O_1881,N_48017,N_48453);
nor UO_1882 (O_1882,N_47510,N_49463);
xnor UO_1883 (O_1883,N_48527,N_48146);
or UO_1884 (O_1884,N_47789,N_48963);
xnor UO_1885 (O_1885,N_47830,N_48114);
or UO_1886 (O_1886,N_49147,N_48819);
nand UO_1887 (O_1887,N_48220,N_49117);
and UO_1888 (O_1888,N_48486,N_49456);
or UO_1889 (O_1889,N_49982,N_49268);
nor UO_1890 (O_1890,N_49467,N_49123);
xnor UO_1891 (O_1891,N_47782,N_47747);
or UO_1892 (O_1892,N_49106,N_49243);
and UO_1893 (O_1893,N_49110,N_49123);
and UO_1894 (O_1894,N_47585,N_48787);
or UO_1895 (O_1895,N_48899,N_49467);
xnor UO_1896 (O_1896,N_49624,N_49382);
nand UO_1897 (O_1897,N_47510,N_47989);
or UO_1898 (O_1898,N_49884,N_48010);
or UO_1899 (O_1899,N_48696,N_47557);
or UO_1900 (O_1900,N_49368,N_48842);
xor UO_1901 (O_1901,N_48543,N_48463);
and UO_1902 (O_1902,N_49996,N_49957);
or UO_1903 (O_1903,N_47793,N_47903);
nand UO_1904 (O_1904,N_47530,N_48126);
nand UO_1905 (O_1905,N_48407,N_47658);
nor UO_1906 (O_1906,N_49610,N_49551);
nor UO_1907 (O_1907,N_48403,N_49239);
and UO_1908 (O_1908,N_49430,N_49421);
nor UO_1909 (O_1909,N_47558,N_48623);
and UO_1910 (O_1910,N_47742,N_49341);
nand UO_1911 (O_1911,N_49020,N_49151);
or UO_1912 (O_1912,N_48269,N_49068);
nor UO_1913 (O_1913,N_48591,N_49834);
and UO_1914 (O_1914,N_48104,N_48012);
and UO_1915 (O_1915,N_48186,N_48147);
nand UO_1916 (O_1916,N_48140,N_49516);
nor UO_1917 (O_1917,N_49684,N_49882);
or UO_1918 (O_1918,N_48084,N_48688);
nor UO_1919 (O_1919,N_47644,N_49311);
xnor UO_1920 (O_1920,N_47786,N_47550);
xor UO_1921 (O_1921,N_48836,N_49584);
and UO_1922 (O_1922,N_47628,N_49562);
and UO_1923 (O_1923,N_49832,N_48893);
xnor UO_1924 (O_1924,N_49212,N_48862);
xnor UO_1925 (O_1925,N_48902,N_49046);
and UO_1926 (O_1926,N_49111,N_48189);
or UO_1927 (O_1927,N_47963,N_48671);
nand UO_1928 (O_1928,N_49993,N_49929);
nand UO_1929 (O_1929,N_49618,N_49549);
and UO_1930 (O_1930,N_47620,N_48641);
nor UO_1931 (O_1931,N_49807,N_49801);
nand UO_1932 (O_1932,N_48627,N_47905);
or UO_1933 (O_1933,N_47501,N_49431);
nand UO_1934 (O_1934,N_47938,N_48112);
nand UO_1935 (O_1935,N_48983,N_48379);
xor UO_1936 (O_1936,N_48584,N_48887);
nor UO_1937 (O_1937,N_49916,N_48182);
or UO_1938 (O_1938,N_48709,N_47899);
nand UO_1939 (O_1939,N_49323,N_47667);
and UO_1940 (O_1940,N_49951,N_49566);
or UO_1941 (O_1941,N_49099,N_49756);
xnor UO_1942 (O_1942,N_48378,N_49952);
nor UO_1943 (O_1943,N_47975,N_47933);
or UO_1944 (O_1944,N_47587,N_49191);
nor UO_1945 (O_1945,N_49262,N_49376);
nor UO_1946 (O_1946,N_47990,N_49129);
nor UO_1947 (O_1947,N_47946,N_49628);
xor UO_1948 (O_1948,N_47596,N_48187);
or UO_1949 (O_1949,N_48609,N_49018);
nor UO_1950 (O_1950,N_48667,N_48697);
or UO_1951 (O_1951,N_47553,N_49936);
nor UO_1952 (O_1952,N_48239,N_48311);
xor UO_1953 (O_1953,N_49480,N_48476);
nor UO_1954 (O_1954,N_49979,N_49991);
nand UO_1955 (O_1955,N_47594,N_49299);
nor UO_1956 (O_1956,N_47776,N_48669);
nor UO_1957 (O_1957,N_48699,N_49636);
xnor UO_1958 (O_1958,N_49925,N_49578);
xor UO_1959 (O_1959,N_47879,N_49675);
and UO_1960 (O_1960,N_48185,N_48458);
and UO_1961 (O_1961,N_49912,N_47823);
nor UO_1962 (O_1962,N_48317,N_49373);
and UO_1963 (O_1963,N_47555,N_49789);
or UO_1964 (O_1964,N_49976,N_48260);
nand UO_1965 (O_1965,N_49891,N_49264);
xnor UO_1966 (O_1966,N_49277,N_47606);
and UO_1967 (O_1967,N_49961,N_48506);
nand UO_1968 (O_1968,N_47734,N_49623);
nand UO_1969 (O_1969,N_48380,N_48798);
or UO_1970 (O_1970,N_49496,N_49070);
xor UO_1971 (O_1971,N_48009,N_48651);
or UO_1972 (O_1972,N_49797,N_48410);
xnor UO_1973 (O_1973,N_47914,N_48001);
nand UO_1974 (O_1974,N_47950,N_49197);
or UO_1975 (O_1975,N_49013,N_48038);
nor UO_1976 (O_1976,N_48207,N_49839);
nor UO_1977 (O_1977,N_47555,N_47756);
xnor UO_1978 (O_1978,N_48629,N_49835);
xnor UO_1979 (O_1979,N_49938,N_49025);
xnor UO_1980 (O_1980,N_49681,N_49870);
xnor UO_1981 (O_1981,N_47782,N_48262);
or UO_1982 (O_1982,N_49735,N_47622);
nor UO_1983 (O_1983,N_48389,N_48443);
nor UO_1984 (O_1984,N_47851,N_49536);
nor UO_1985 (O_1985,N_48964,N_48959);
and UO_1986 (O_1986,N_48824,N_48091);
or UO_1987 (O_1987,N_49772,N_49611);
or UO_1988 (O_1988,N_49586,N_48097);
and UO_1989 (O_1989,N_49011,N_49328);
and UO_1990 (O_1990,N_49092,N_48333);
or UO_1991 (O_1991,N_49151,N_47768);
nor UO_1992 (O_1992,N_49054,N_49240);
and UO_1993 (O_1993,N_49803,N_48916);
nor UO_1994 (O_1994,N_49524,N_49370);
and UO_1995 (O_1995,N_48454,N_49161);
xor UO_1996 (O_1996,N_49966,N_48190);
or UO_1997 (O_1997,N_48552,N_49942);
xnor UO_1998 (O_1998,N_47705,N_48008);
nand UO_1999 (O_1999,N_49394,N_49052);
nand UO_2000 (O_2000,N_49414,N_47615);
and UO_2001 (O_2001,N_48856,N_49044);
or UO_2002 (O_2002,N_47586,N_47921);
nor UO_2003 (O_2003,N_49629,N_49252);
nor UO_2004 (O_2004,N_49517,N_49092);
and UO_2005 (O_2005,N_49957,N_47619);
nand UO_2006 (O_2006,N_48577,N_47597);
xnor UO_2007 (O_2007,N_49724,N_49111);
xor UO_2008 (O_2008,N_48709,N_49496);
or UO_2009 (O_2009,N_49103,N_47743);
nand UO_2010 (O_2010,N_48391,N_48084);
nor UO_2011 (O_2011,N_49240,N_48696);
xor UO_2012 (O_2012,N_47649,N_47650);
and UO_2013 (O_2013,N_49821,N_47913);
or UO_2014 (O_2014,N_49386,N_49593);
or UO_2015 (O_2015,N_47754,N_49069);
or UO_2016 (O_2016,N_47746,N_47987);
nand UO_2017 (O_2017,N_48886,N_48304);
nand UO_2018 (O_2018,N_49886,N_48543);
and UO_2019 (O_2019,N_48115,N_49130);
nor UO_2020 (O_2020,N_47988,N_48573);
nand UO_2021 (O_2021,N_48007,N_48707);
or UO_2022 (O_2022,N_48632,N_48605);
and UO_2023 (O_2023,N_47821,N_49187);
or UO_2024 (O_2024,N_49630,N_48145);
or UO_2025 (O_2025,N_48919,N_49365);
nand UO_2026 (O_2026,N_49831,N_47513);
nor UO_2027 (O_2027,N_49822,N_48903);
or UO_2028 (O_2028,N_48674,N_47817);
and UO_2029 (O_2029,N_48918,N_47516);
or UO_2030 (O_2030,N_48218,N_49970);
nand UO_2031 (O_2031,N_48909,N_47820);
nor UO_2032 (O_2032,N_48210,N_47861);
nand UO_2033 (O_2033,N_48489,N_49252);
xnor UO_2034 (O_2034,N_49780,N_49403);
nand UO_2035 (O_2035,N_47976,N_48463);
xor UO_2036 (O_2036,N_47693,N_47789);
and UO_2037 (O_2037,N_47912,N_47825);
nor UO_2038 (O_2038,N_49204,N_49582);
or UO_2039 (O_2039,N_47987,N_49875);
or UO_2040 (O_2040,N_47817,N_48601);
nor UO_2041 (O_2041,N_48596,N_47732);
or UO_2042 (O_2042,N_48407,N_49293);
or UO_2043 (O_2043,N_48728,N_49836);
nor UO_2044 (O_2044,N_49325,N_47843);
and UO_2045 (O_2045,N_49399,N_49255);
or UO_2046 (O_2046,N_47716,N_47634);
nand UO_2047 (O_2047,N_49609,N_49326);
or UO_2048 (O_2048,N_48483,N_48560);
and UO_2049 (O_2049,N_49159,N_47999);
or UO_2050 (O_2050,N_49695,N_49576);
nor UO_2051 (O_2051,N_48707,N_49941);
nor UO_2052 (O_2052,N_49041,N_49791);
and UO_2053 (O_2053,N_48945,N_49763);
xor UO_2054 (O_2054,N_49437,N_49596);
and UO_2055 (O_2055,N_48839,N_48903);
xor UO_2056 (O_2056,N_48582,N_47725);
nor UO_2057 (O_2057,N_47574,N_49827);
and UO_2058 (O_2058,N_48139,N_48590);
nand UO_2059 (O_2059,N_48395,N_49730);
and UO_2060 (O_2060,N_49381,N_48217);
xnor UO_2061 (O_2061,N_47549,N_49957);
nor UO_2062 (O_2062,N_47971,N_48450);
nand UO_2063 (O_2063,N_49596,N_49169);
nand UO_2064 (O_2064,N_48451,N_47687);
xnor UO_2065 (O_2065,N_48050,N_47830);
or UO_2066 (O_2066,N_48052,N_48964);
nand UO_2067 (O_2067,N_47606,N_49740);
nor UO_2068 (O_2068,N_49006,N_48234);
and UO_2069 (O_2069,N_48503,N_49808);
or UO_2070 (O_2070,N_48026,N_47648);
xnor UO_2071 (O_2071,N_48174,N_48669);
or UO_2072 (O_2072,N_48016,N_49859);
or UO_2073 (O_2073,N_48146,N_48652);
xor UO_2074 (O_2074,N_49317,N_49645);
or UO_2075 (O_2075,N_47606,N_48376);
nand UO_2076 (O_2076,N_49121,N_49460);
xnor UO_2077 (O_2077,N_48464,N_48546);
xor UO_2078 (O_2078,N_48515,N_48128);
nand UO_2079 (O_2079,N_49504,N_47760);
nand UO_2080 (O_2080,N_47521,N_48071);
and UO_2081 (O_2081,N_48930,N_47989);
and UO_2082 (O_2082,N_48175,N_48628);
nor UO_2083 (O_2083,N_47962,N_49477);
nor UO_2084 (O_2084,N_49172,N_49800);
and UO_2085 (O_2085,N_49666,N_48647);
xor UO_2086 (O_2086,N_49015,N_48156);
xnor UO_2087 (O_2087,N_48366,N_49174);
nand UO_2088 (O_2088,N_49030,N_49368);
nor UO_2089 (O_2089,N_47658,N_48947);
nor UO_2090 (O_2090,N_48411,N_48187);
nor UO_2091 (O_2091,N_49321,N_47635);
xnor UO_2092 (O_2092,N_48362,N_47967);
xnor UO_2093 (O_2093,N_48420,N_49194);
and UO_2094 (O_2094,N_47879,N_48488);
or UO_2095 (O_2095,N_49494,N_47701);
or UO_2096 (O_2096,N_49952,N_48084);
nor UO_2097 (O_2097,N_47887,N_49992);
or UO_2098 (O_2098,N_48454,N_49063);
or UO_2099 (O_2099,N_47814,N_49817);
and UO_2100 (O_2100,N_49493,N_48783);
or UO_2101 (O_2101,N_49445,N_49906);
and UO_2102 (O_2102,N_49382,N_48649);
or UO_2103 (O_2103,N_47864,N_48246);
nand UO_2104 (O_2104,N_48917,N_48546);
and UO_2105 (O_2105,N_47562,N_48157);
xor UO_2106 (O_2106,N_47647,N_48790);
or UO_2107 (O_2107,N_49967,N_49801);
or UO_2108 (O_2108,N_48870,N_49886);
or UO_2109 (O_2109,N_48798,N_49013);
xor UO_2110 (O_2110,N_49754,N_48289);
and UO_2111 (O_2111,N_48449,N_48995);
nand UO_2112 (O_2112,N_48703,N_47744);
xnor UO_2113 (O_2113,N_47970,N_47560);
nor UO_2114 (O_2114,N_49959,N_48788);
or UO_2115 (O_2115,N_48489,N_47726);
nand UO_2116 (O_2116,N_48242,N_48227);
and UO_2117 (O_2117,N_48287,N_49601);
and UO_2118 (O_2118,N_47500,N_49081);
and UO_2119 (O_2119,N_49197,N_48532);
xor UO_2120 (O_2120,N_49364,N_47582);
nand UO_2121 (O_2121,N_48639,N_48770);
nand UO_2122 (O_2122,N_48699,N_48711);
or UO_2123 (O_2123,N_49330,N_48611);
or UO_2124 (O_2124,N_48965,N_48659);
nor UO_2125 (O_2125,N_48905,N_49803);
nand UO_2126 (O_2126,N_47898,N_48901);
xnor UO_2127 (O_2127,N_49746,N_49166);
and UO_2128 (O_2128,N_49785,N_48756);
xnor UO_2129 (O_2129,N_49750,N_47971);
or UO_2130 (O_2130,N_48736,N_47688);
nand UO_2131 (O_2131,N_49344,N_48028);
nand UO_2132 (O_2132,N_47737,N_47508);
nor UO_2133 (O_2133,N_47897,N_48660);
nor UO_2134 (O_2134,N_49083,N_49763);
nand UO_2135 (O_2135,N_49481,N_48712);
nand UO_2136 (O_2136,N_48330,N_49094);
nand UO_2137 (O_2137,N_49803,N_48626);
xnor UO_2138 (O_2138,N_49646,N_48622);
nand UO_2139 (O_2139,N_49057,N_47775);
or UO_2140 (O_2140,N_47859,N_49798);
or UO_2141 (O_2141,N_47548,N_47522);
and UO_2142 (O_2142,N_49374,N_47844);
nor UO_2143 (O_2143,N_48282,N_49426);
nand UO_2144 (O_2144,N_49228,N_49590);
and UO_2145 (O_2145,N_49144,N_49436);
nor UO_2146 (O_2146,N_48742,N_49505);
or UO_2147 (O_2147,N_48387,N_48023);
nor UO_2148 (O_2148,N_47993,N_48970);
xnor UO_2149 (O_2149,N_49028,N_49151);
xor UO_2150 (O_2150,N_48641,N_49119);
xor UO_2151 (O_2151,N_49714,N_49996);
and UO_2152 (O_2152,N_47735,N_47963);
or UO_2153 (O_2153,N_49942,N_47949);
nand UO_2154 (O_2154,N_49731,N_48405);
and UO_2155 (O_2155,N_48361,N_49020);
nand UO_2156 (O_2156,N_49975,N_49107);
nand UO_2157 (O_2157,N_48283,N_49489);
nand UO_2158 (O_2158,N_48892,N_49396);
nor UO_2159 (O_2159,N_48086,N_47898);
or UO_2160 (O_2160,N_49040,N_48817);
xnor UO_2161 (O_2161,N_49654,N_48414);
xor UO_2162 (O_2162,N_48365,N_49875);
xnor UO_2163 (O_2163,N_48011,N_49824);
and UO_2164 (O_2164,N_49696,N_48084);
or UO_2165 (O_2165,N_49941,N_48070);
xnor UO_2166 (O_2166,N_49344,N_49684);
or UO_2167 (O_2167,N_48804,N_47525);
xor UO_2168 (O_2168,N_48356,N_48871);
nand UO_2169 (O_2169,N_49310,N_47966);
nor UO_2170 (O_2170,N_49153,N_48821);
and UO_2171 (O_2171,N_49993,N_49647);
and UO_2172 (O_2172,N_47777,N_48330);
or UO_2173 (O_2173,N_48492,N_48540);
or UO_2174 (O_2174,N_48079,N_47929);
and UO_2175 (O_2175,N_47833,N_49393);
nand UO_2176 (O_2176,N_48099,N_47739);
nor UO_2177 (O_2177,N_49817,N_48584);
and UO_2178 (O_2178,N_48273,N_48260);
xnor UO_2179 (O_2179,N_49610,N_49298);
nor UO_2180 (O_2180,N_49050,N_49670);
and UO_2181 (O_2181,N_49785,N_48413);
nor UO_2182 (O_2182,N_49843,N_47518);
and UO_2183 (O_2183,N_49461,N_48681);
or UO_2184 (O_2184,N_49430,N_48893);
or UO_2185 (O_2185,N_47527,N_48581);
nor UO_2186 (O_2186,N_49443,N_48897);
nand UO_2187 (O_2187,N_48539,N_49583);
nor UO_2188 (O_2188,N_49789,N_48815);
nor UO_2189 (O_2189,N_48993,N_47981);
nand UO_2190 (O_2190,N_48307,N_48721);
nand UO_2191 (O_2191,N_48610,N_48113);
xnor UO_2192 (O_2192,N_48313,N_48382);
and UO_2193 (O_2193,N_49718,N_49773);
nor UO_2194 (O_2194,N_49905,N_48171);
xor UO_2195 (O_2195,N_47907,N_48269);
or UO_2196 (O_2196,N_47845,N_49178);
and UO_2197 (O_2197,N_48050,N_48600);
nor UO_2198 (O_2198,N_48876,N_49543);
or UO_2199 (O_2199,N_49775,N_49662);
or UO_2200 (O_2200,N_49405,N_49321);
or UO_2201 (O_2201,N_49162,N_49834);
and UO_2202 (O_2202,N_47890,N_48364);
nor UO_2203 (O_2203,N_48050,N_47974);
and UO_2204 (O_2204,N_48616,N_48545);
nand UO_2205 (O_2205,N_48232,N_47748);
xnor UO_2206 (O_2206,N_47884,N_47741);
xnor UO_2207 (O_2207,N_48605,N_49027);
or UO_2208 (O_2208,N_49457,N_48737);
or UO_2209 (O_2209,N_48943,N_48123);
and UO_2210 (O_2210,N_48119,N_47827);
and UO_2211 (O_2211,N_47576,N_48076);
nor UO_2212 (O_2212,N_49148,N_47644);
nor UO_2213 (O_2213,N_47789,N_49169);
xnor UO_2214 (O_2214,N_48780,N_49565);
nand UO_2215 (O_2215,N_48092,N_48900);
nand UO_2216 (O_2216,N_48998,N_49889);
and UO_2217 (O_2217,N_49548,N_49223);
nand UO_2218 (O_2218,N_48809,N_48683);
nand UO_2219 (O_2219,N_48424,N_47671);
or UO_2220 (O_2220,N_47535,N_49527);
or UO_2221 (O_2221,N_49979,N_47557);
or UO_2222 (O_2222,N_48220,N_49429);
nor UO_2223 (O_2223,N_47727,N_47745);
xor UO_2224 (O_2224,N_49647,N_49042);
xnor UO_2225 (O_2225,N_48678,N_48642);
nor UO_2226 (O_2226,N_47626,N_48110);
and UO_2227 (O_2227,N_48958,N_48080);
nand UO_2228 (O_2228,N_49235,N_49255);
and UO_2229 (O_2229,N_48848,N_49674);
and UO_2230 (O_2230,N_48743,N_48818);
or UO_2231 (O_2231,N_48797,N_48897);
and UO_2232 (O_2232,N_49570,N_49797);
and UO_2233 (O_2233,N_49038,N_47929);
xor UO_2234 (O_2234,N_47738,N_47677);
xor UO_2235 (O_2235,N_47735,N_48164);
and UO_2236 (O_2236,N_48703,N_48274);
nand UO_2237 (O_2237,N_49655,N_49337);
and UO_2238 (O_2238,N_47876,N_48960);
nand UO_2239 (O_2239,N_49062,N_49048);
nand UO_2240 (O_2240,N_49982,N_47621);
and UO_2241 (O_2241,N_49238,N_49411);
or UO_2242 (O_2242,N_49542,N_49362);
and UO_2243 (O_2243,N_49533,N_49834);
nor UO_2244 (O_2244,N_48646,N_48712);
and UO_2245 (O_2245,N_48332,N_49687);
xor UO_2246 (O_2246,N_48155,N_47532);
xnor UO_2247 (O_2247,N_48257,N_47995);
xor UO_2248 (O_2248,N_47741,N_49749);
or UO_2249 (O_2249,N_49116,N_48034);
nor UO_2250 (O_2250,N_48146,N_49005);
nor UO_2251 (O_2251,N_47924,N_49895);
nand UO_2252 (O_2252,N_49479,N_49553);
nor UO_2253 (O_2253,N_48945,N_48052);
xnor UO_2254 (O_2254,N_48175,N_48778);
or UO_2255 (O_2255,N_49805,N_49987);
or UO_2256 (O_2256,N_48145,N_47772);
nor UO_2257 (O_2257,N_48113,N_47703);
xor UO_2258 (O_2258,N_47988,N_48642);
nor UO_2259 (O_2259,N_49146,N_47592);
xnor UO_2260 (O_2260,N_49075,N_48078);
and UO_2261 (O_2261,N_47663,N_48456);
and UO_2262 (O_2262,N_49090,N_48695);
nand UO_2263 (O_2263,N_48752,N_48337);
or UO_2264 (O_2264,N_48419,N_47628);
nor UO_2265 (O_2265,N_49656,N_49729);
nand UO_2266 (O_2266,N_47501,N_49514);
or UO_2267 (O_2267,N_49160,N_48831);
or UO_2268 (O_2268,N_48766,N_48853);
nor UO_2269 (O_2269,N_48575,N_49399);
xnor UO_2270 (O_2270,N_48233,N_48544);
nand UO_2271 (O_2271,N_48814,N_49740);
or UO_2272 (O_2272,N_48715,N_48268);
nand UO_2273 (O_2273,N_48180,N_48243);
nor UO_2274 (O_2274,N_49004,N_49512);
and UO_2275 (O_2275,N_48655,N_49641);
and UO_2276 (O_2276,N_49016,N_49123);
or UO_2277 (O_2277,N_49718,N_48585);
nor UO_2278 (O_2278,N_49032,N_47683);
and UO_2279 (O_2279,N_48734,N_49314);
nand UO_2280 (O_2280,N_49017,N_47979);
and UO_2281 (O_2281,N_49946,N_48516);
or UO_2282 (O_2282,N_48220,N_49524);
and UO_2283 (O_2283,N_49653,N_49480);
nor UO_2284 (O_2284,N_49745,N_48410);
and UO_2285 (O_2285,N_49292,N_49359);
nor UO_2286 (O_2286,N_49965,N_49996);
nor UO_2287 (O_2287,N_48983,N_48741);
nand UO_2288 (O_2288,N_48974,N_47731);
or UO_2289 (O_2289,N_49803,N_49815);
or UO_2290 (O_2290,N_49697,N_49249);
xor UO_2291 (O_2291,N_49931,N_48671);
and UO_2292 (O_2292,N_49127,N_47702);
and UO_2293 (O_2293,N_49551,N_49915);
nor UO_2294 (O_2294,N_47810,N_48771);
and UO_2295 (O_2295,N_47560,N_47525);
nand UO_2296 (O_2296,N_49344,N_49601);
xor UO_2297 (O_2297,N_49340,N_49235);
nand UO_2298 (O_2298,N_48128,N_48786);
and UO_2299 (O_2299,N_49022,N_49926);
and UO_2300 (O_2300,N_48198,N_48127);
nor UO_2301 (O_2301,N_47810,N_47617);
nor UO_2302 (O_2302,N_48963,N_48185);
nand UO_2303 (O_2303,N_49088,N_48715);
nor UO_2304 (O_2304,N_47851,N_49098);
or UO_2305 (O_2305,N_48486,N_49569);
xnor UO_2306 (O_2306,N_48938,N_48302);
nor UO_2307 (O_2307,N_47920,N_47950);
nand UO_2308 (O_2308,N_48181,N_47782);
nand UO_2309 (O_2309,N_49725,N_49864);
nand UO_2310 (O_2310,N_48153,N_47738);
xor UO_2311 (O_2311,N_49759,N_47614);
xor UO_2312 (O_2312,N_49613,N_48603);
and UO_2313 (O_2313,N_49562,N_47914);
nand UO_2314 (O_2314,N_49700,N_48849);
xor UO_2315 (O_2315,N_48201,N_49077);
nand UO_2316 (O_2316,N_49571,N_47645);
or UO_2317 (O_2317,N_47535,N_47575);
nand UO_2318 (O_2318,N_49511,N_49814);
or UO_2319 (O_2319,N_48448,N_49713);
and UO_2320 (O_2320,N_48492,N_49321);
and UO_2321 (O_2321,N_49489,N_47661);
nor UO_2322 (O_2322,N_47531,N_48528);
nand UO_2323 (O_2323,N_49017,N_49256);
and UO_2324 (O_2324,N_47766,N_47925);
or UO_2325 (O_2325,N_49872,N_48987);
nor UO_2326 (O_2326,N_48385,N_47576);
xor UO_2327 (O_2327,N_49904,N_47892);
nand UO_2328 (O_2328,N_48261,N_48158);
and UO_2329 (O_2329,N_49931,N_48361);
xor UO_2330 (O_2330,N_49451,N_49741);
xor UO_2331 (O_2331,N_48760,N_49508);
and UO_2332 (O_2332,N_49465,N_48619);
and UO_2333 (O_2333,N_48867,N_47984);
xnor UO_2334 (O_2334,N_48982,N_49083);
xnor UO_2335 (O_2335,N_47752,N_47557);
nor UO_2336 (O_2336,N_48770,N_49200);
nor UO_2337 (O_2337,N_49154,N_47524);
and UO_2338 (O_2338,N_48549,N_49946);
nand UO_2339 (O_2339,N_49097,N_48480);
or UO_2340 (O_2340,N_49391,N_47517);
nor UO_2341 (O_2341,N_48297,N_47845);
and UO_2342 (O_2342,N_48146,N_48508);
and UO_2343 (O_2343,N_47917,N_48396);
nor UO_2344 (O_2344,N_49673,N_47802);
and UO_2345 (O_2345,N_47646,N_49177);
xor UO_2346 (O_2346,N_48357,N_48531);
and UO_2347 (O_2347,N_49522,N_47994);
xnor UO_2348 (O_2348,N_48286,N_49609);
or UO_2349 (O_2349,N_48121,N_47642);
xor UO_2350 (O_2350,N_49479,N_48011);
nand UO_2351 (O_2351,N_47919,N_47900);
and UO_2352 (O_2352,N_49275,N_49816);
xor UO_2353 (O_2353,N_48325,N_48261);
nand UO_2354 (O_2354,N_48557,N_49787);
or UO_2355 (O_2355,N_48578,N_47879);
and UO_2356 (O_2356,N_47775,N_47886);
xnor UO_2357 (O_2357,N_48812,N_48582);
nor UO_2358 (O_2358,N_47581,N_49116);
nor UO_2359 (O_2359,N_48809,N_49438);
nor UO_2360 (O_2360,N_49175,N_47910);
or UO_2361 (O_2361,N_49802,N_49847);
or UO_2362 (O_2362,N_49511,N_49304);
and UO_2363 (O_2363,N_49471,N_47685);
and UO_2364 (O_2364,N_49307,N_49842);
xnor UO_2365 (O_2365,N_49450,N_48767);
or UO_2366 (O_2366,N_49445,N_47820);
nand UO_2367 (O_2367,N_48770,N_48194);
nand UO_2368 (O_2368,N_49201,N_48981);
nor UO_2369 (O_2369,N_47897,N_47790);
nor UO_2370 (O_2370,N_49882,N_48046);
xnor UO_2371 (O_2371,N_47763,N_47907);
nand UO_2372 (O_2372,N_48514,N_49690);
nor UO_2373 (O_2373,N_49754,N_47787);
and UO_2374 (O_2374,N_49303,N_49158);
nor UO_2375 (O_2375,N_49123,N_49854);
nand UO_2376 (O_2376,N_47862,N_49091);
or UO_2377 (O_2377,N_49547,N_48179);
xor UO_2378 (O_2378,N_48305,N_48652);
nor UO_2379 (O_2379,N_47658,N_48051);
xor UO_2380 (O_2380,N_48381,N_49367);
or UO_2381 (O_2381,N_49069,N_48952);
nand UO_2382 (O_2382,N_48683,N_49880);
nor UO_2383 (O_2383,N_47512,N_49219);
and UO_2384 (O_2384,N_48329,N_49488);
nor UO_2385 (O_2385,N_49818,N_49882);
or UO_2386 (O_2386,N_49907,N_49024);
and UO_2387 (O_2387,N_49572,N_47614);
nand UO_2388 (O_2388,N_48176,N_48260);
or UO_2389 (O_2389,N_47982,N_48862);
nand UO_2390 (O_2390,N_49155,N_47627);
nor UO_2391 (O_2391,N_48478,N_48721);
and UO_2392 (O_2392,N_47854,N_49081);
xnor UO_2393 (O_2393,N_49667,N_48857);
or UO_2394 (O_2394,N_48420,N_48893);
or UO_2395 (O_2395,N_49780,N_49846);
and UO_2396 (O_2396,N_47537,N_48587);
or UO_2397 (O_2397,N_49685,N_49591);
xor UO_2398 (O_2398,N_48099,N_48661);
and UO_2399 (O_2399,N_48962,N_49310);
or UO_2400 (O_2400,N_48206,N_49449);
or UO_2401 (O_2401,N_49645,N_48960);
or UO_2402 (O_2402,N_48741,N_48605);
or UO_2403 (O_2403,N_48043,N_47958);
and UO_2404 (O_2404,N_48158,N_47567);
nor UO_2405 (O_2405,N_49807,N_49661);
xnor UO_2406 (O_2406,N_49270,N_47549);
and UO_2407 (O_2407,N_48965,N_49706);
nand UO_2408 (O_2408,N_48847,N_49144);
or UO_2409 (O_2409,N_49282,N_49094);
and UO_2410 (O_2410,N_49502,N_49410);
nor UO_2411 (O_2411,N_49095,N_48965);
nand UO_2412 (O_2412,N_49249,N_49778);
and UO_2413 (O_2413,N_48974,N_49599);
and UO_2414 (O_2414,N_48210,N_49031);
xnor UO_2415 (O_2415,N_49891,N_49921);
nand UO_2416 (O_2416,N_49241,N_48125);
xor UO_2417 (O_2417,N_48070,N_47539);
nand UO_2418 (O_2418,N_48613,N_48931);
xnor UO_2419 (O_2419,N_47958,N_48431);
xor UO_2420 (O_2420,N_47517,N_49020);
nor UO_2421 (O_2421,N_49177,N_49690);
nand UO_2422 (O_2422,N_49272,N_48833);
and UO_2423 (O_2423,N_48126,N_47942);
and UO_2424 (O_2424,N_49606,N_47947);
nand UO_2425 (O_2425,N_49078,N_48100);
and UO_2426 (O_2426,N_48972,N_48865);
or UO_2427 (O_2427,N_49935,N_47638);
xnor UO_2428 (O_2428,N_47858,N_49398);
or UO_2429 (O_2429,N_48883,N_49525);
nor UO_2430 (O_2430,N_48781,N_47534);
xor UO_2431 (O_2431,N_49791,N_48914);
and UO_2432 (O_2432,N_48227,N_47561);
or UO_2433 (O_2433,N_49484,N_49936);
xnor UO_2434 (O_2434,N_48469,N_49913);
nor UO_2435 (O_2435,N_48077,N_47854);
nor UO_2436 (O_2436,N_49158,N_47950);
nand UO_2437 (O_2437,N_48967,N_48923);
nor UO_2438 (O_2438,N_49047,N_48156);
or UO_2439 (O_2439,N_48027,N_48814);
xnor UO_2440 (O_2440,N_49038,N_48267);
or UO_2441 (O_2441,N_48123,N_49539);
and UO_2442 (O_2442,N_48166,N_49432);
and UO_2443 (O_2443,N_49988,N_49496);
and UO_2444 (O_2444,N_48452,N_48045);
xnor UO_2445 (O_2445,N_48254,N_48932);
and UO_2446 (O_2446,N_49965,N_48866);
nand UO_2447 (O_2447,N_47545,N_49618);
and UO_2448 (O_2448,N_48830,N_49595);
nor UO_2449 (O_2449,N_49040,N_49797);
or UO_2450 (O_2450,N_48362,N_47535);
nand UO_2451 (O_2451,N_49753,N_49399);
nand UO_2452 (O_2452,N_48055,N_47736);
nor UO_2453 (O_2453,N_47570,N_47751);
and UO_2454 (O_2454,N_47824,N_48318);
xnor UO_2455 (O_2455,N_49746,N_47557);
and UO_2456 (O_2456,N_49112,N_48621);
nor UO_2457 (O_2457,N_48719,N_47897);
xnor UO_2458 (O_2458,N_48075,N_49316);
nor UO_2459 (O_2459,N_47575,N_47611);
nand UO_2460 (O_2460,N_48159,N_47789);
nand UO_2461 (O_2461,N_48679,N_49071);
and UO_2462 (O_2462,N_48010,N_48502);
or UO_2463 (O_2463,N_48311,N_49946);
and UO_2464 (O_2464,N_48505,N_48115);
nor UO_2465 (O_2465,N_49191,N_48002);
or UO_2466 (O_2466,N_49695,N_49489);
and UO_2467 (O_2467,N_48581,N_48185);
xnor UO_2468 (O_2468,N_49772,N_48362);
or UO_2469 (O_2469,N_49292,N_48483);
nand UO_2470 (O_2470,N_49640,N_48073);
or UO_2471 (O_2471,N_49656,N_47961);
or UO_2472 (O_2472,N_47797,N_49647);
or UO_2473 (O_2473,N_47854,N_48284);
and UO_2474 (O_2474,N_49323,N_49114);
xor UO_2475 (O_2475,N_47514,N_47675);
and UO_2476 (O_2476,N_49029,N_49449);
nor UO_2477 (O_2477,N_49093,N_49444);
nor UO_2478 (O_2478,N_47892,N_47910);
nand UO_2479 (O_2479,N_48489,N_47760);
or UO_2480 (O_2480,N_48707,N_47831);
and UO_2481 (O_2481,N_49780,N_49423);
or UO_2482 (O_2482,N_48005,N_47710);
and UO_2483 (O_2483,N_48765,N_49290);
nor UO_2484 (O_2484,N_49396,N_49229);
xnor UO_2485 (O_2485,N_48250,N_47837);
nor UO_2486 (O_2486,N_49630,N_47857);
xor UO_2487 (O_2487,N_49342,N_48601);
xnor UO_2488 (O_2488,N_49091,N_48071);
and UO_2489 (O_2489,N_49707,N_49448);
and UO_2490 (O_2490,N_49832,N_48112);
and UO_2491 (O_2491,N_49364,N_49286);
and UO_2492 (O_2492,N_49843,N_48137);
and UO_2493 (O_2493,N_47881,N_49321);
xor UO_2494 (O_2494,N_49247,N_49352);
nor UO_2495 (O_2495,N_47911,N_47881);
and UO_2496 (O_2496,N_47822,N_49914);
nor UO_2497 (O_2497,N_47757,N_48622);
nand UO_2498 (O_2498,N_49969,N_49210);
and UO_2499 (O_2499,N_47500,N_48867);
and UO_2500 (O_2500,N_49642,N_48904);
xnor UO_2501 (O_2501,N_49769,N_49810);
nor UO_2502 (O_2502,N_47845,N_48855);
nor UO_2503 (O_2503,N_48815,N_48765);
nand UO_2504 (O_2504,N_49994,N_48218);
nor UO_2505 (O_2505,N_49920,N_48374);
nor UO_2506 (O_2506,N_47630,N_48801);
nor UO_2507 (O_2507,N_49995,N_48868);
xnor UO_2508 (O_2508,N_48786,N_47843);
or UO_2509 (O_2509,N_49917,N_48760);
nand UO_2510 (O_2510,N_47738,N_48950);
or UO_2511 (O_2511,N_48299,N_48707);
or UO_2512 (O_2512,N_48012,N_49176);
or UO_2513 (O_2513,N_49438,N_49575);
or UO_2514 (O_2514,N_49388,N_49734);
xnor UO_2515 (O_2515,N_48171,N_49368);
xnor UO_2516 (O_2516,N_47582,N_47623);
nand UO_2517 (O_2517,N_48611,N_48362);
or UO_2518 (O_2518,N_48033,N_48038);
or UO_2519 (O_2519,N_48461,N_49627);
and UO_2520 (O_2520,N_48594,N_48948);
and UO_2521 (O_2521,N_48607,N_49442);
nor UO_2522 (O_2522,N_48039,N_49741);
xor UO_2523 (O_2523,N_48281,N_49544);
nor UO_2524 (O_2524,N_48803,N_49897);
and UO_2525 (O_2525,N_47714,N_49804);
nor UO_2526 (O_2526,N_49383,N_47627);
or UO_2527 (O_2527,N_49846,N_48517);
and UO_2528 (O_2528,N_48206,N_48529);
or UO_2529 (O_2529,N_47869,N_49224);
nand UO_2530 (O_2530,N_49940,N_49972);
xor UO_2531 (O_2531,N_48198,N_49939);
or UO_2532 (O_2532,N_49108,N_49177);
and UO_2533 (O_2533,N_49226,N_49867);
xnor UO_2534 (O_2534,N_49823,N_49210);
or UO_2535 (O_2535,N_48651,N_48557);
nand UO_2536 (O_2536,N_48730,N_47655);
xor UO_2537 (O_2537,N_49368,N_49823);
or UO_2538 (O_2538,N_49068,N_49191);
or UO_2539 (O_2539,N_49594,N_48749);
nor UO_2540 (O_2540,N_49493,N_48110);
nor UO_2541 (O_2541,N_48352,N_48694);
nand UO_2542 (O_2542,N_49552,N_48439);
xor UO_2543 (O_2543,N_48250,N_48186);
nor UO_2544 (O_2544,N_48318,N_48734);
and UO_2545 (O_2545,N_48238,N_48792);
nor UO_2546 (O_2546,N_49931,N_48568);
nand UO_2547 (O_2547,N_48418,N_48191);
xor UO_2548 (O_2548,N_47955,N_49039);
nand UO_2549 (O_2549,N_49911,N_49212);
and UO_2550 (O_2550,N_49761,N_48653);
or UO_2551 (O_2551,N_48720,N_49752);
and UO_2552 (O_2552,N_47699,N_49948);
and UO_2553 (O_2553,N_49114,N_49285);
xor UO_2554 (O_2554,N_48802,N_49415);
xor UO_2555 (O_2555,N_47842,N_49438);
nand UO_2556 (O_2556,N_49484,N_48605);
or UO_2557 (O_2557,N_49323,N_49041);
or UO_2558 (O_2558,N_49335,N_47651);
nor UO_2559 (O_2559,N_49620,N_47968);
or UO_2560 (O_2560,N_48197,N_49028);
nand UO_2561 (O_2561,N_47778,N_47680);
and UO_2562 (O_2562,N_49188,N_49996);
xnor UO_2563 (O_2563,N_49925,N_49385);
nor UO_2564 (O_2564,N_47941,N_48487);
xnor UO_2565 (O_2565,N_48528,N_47821);
and UO_2566 (O_2566,N_48481,N_49219);
nor UO_2567 (O_2567,N_48708,N_48839);
nor UO_2568 (O_2568,N_48191,N_48654);
and UO_2569 (O_2569,N_48101,N_48884);
xor UO_2570 (O_2570,N_49157,N_47871);
nor UO_2571 (O_2571,N_47769,N_48756);
nor UO_2572 (O_2572,N_49691,N_48879);
nand UO_2573 (O_2573,N_47698,N_49166);
xor UO_2574 (O_2574,N_49887,N_48387);
and UO_2575 (O_2575,N_48800,N_48829);
nand UO_2576 (O_2576,N_48915,N_48640);
or UO_2577 (O_2577,N_48841,N_48574);
and UO_2578 (O_2578,N_47911,N_49645);
xnor UO_2579 (O_2579,N_48293,N_49114);
nor UO_2580 (O_2580,N_49356,N_48341);
or UO_2581 (O_2581,N_49280,N_49876);
nor UO_2582 (O_2582,N_47927,N_49151);
or UO_2583 (O_2583,N_47822,N_48793);
xor UO_2584 (O_2584,N_49007,N_47998);
or UO_2585 (O_2585,N_49811,N_48886);
xnor UO_2586 (O_2586,N_49587,N_49249);
or UO_2587 (O_2587,N_49838,N_49111);
or UO_2588 (O_2588,N_48177,N_49612);
and UO_2589 (O_2589,N_47552,N_48568);
nand UO_2590 (O_2590,N_48546,N_48919);
or UO_2591 (O_2591,N_49834,N_47766);
or UO_2592 (O_2592,N_49831,N_48333);
nand UO_2593 (O_2593,N_47563,N_48702);
or UO_2594 (O_2594,N_48580,N_49723);
xnor UO_2595 (O_2595,N_48565,N_49346);
or UO_2596 (O_2596,N_48007,N_48613);
nand UO_2597 (O_2597,N_47671,N_48068);
xnor UO_2598 (O_2598,N_49794,N_48912);
nor UO_2599 (O_2599,N_47652,N_49733);
nand UO_2600 (O_2600,N_49807,N_48524);
xnor UO_2601 (O_2601,N_49639,N_48998);
xnor UO_2602 (O_2602,N_47578,N_49881);
nor UO_2603 (O_2603,N_47854,N_49168);
and UO_2604 (O_2604,N_49118,N_49941);
nand UO_2605 (O_2605,N_47948,N_48917);
and UO_2606 (O_2606,N_48416,N_47978);
xnor UO_2607 (O_2607,N_49469,N_47529);
nor UO_2608 (O_2608,N_47535,N_48074);
nor UO_2609 (O_2609,N_49033,N_47676);
or UO_2610 (O_2610,N_49443,N_49835);
xnor UO_2611 (O_2611,N_48183,N_49827);
and UO_2612 (O_2612,N_49110,N_49609);
xnor UO_2613 (O_2613,N_48353,N_47594);
xnor UO_2614 (O_2614,N_48162,N_48110);
or UO_2615 (O_2615,N_48188,N_49964);
and UO_2616 (O_2616,N_49508,N_48955);
or UO_2617 (O_2617,N_47702,N_49464);
nand UO_2618 (O_2618,N_48149,N_47840);
nor UO_2619 (O_2619,N_49116,N_49151);
nor UO_2620 (O_2620,N_48112,N_47833);
and UO_2621 (O_2621,N_49574,N_49580);
nand UO_2622 (O_2622,N_49189,N_48395);
xnor UO_2623 (O_2623,N_49916,N_47943);
xor UO_2624 (O_2624,N_49261,N_49714);
xnor UO_2625 (O_2625,N_49872,N_49532);
or UO_2626 (O_2626,N_49775,N_49874);
nand UO_2627 (O_2627,N_48443,N_48162);
xnor UO_2628 (O_2628,N_49780,N_49895);
xnor UO_2629 (O_2629,N_48520,N_49060);
nand UO_2630 (O_2630,N_49139,N_48530);
or UO_2631 (O_2631,N_49352,N_49104);
xor UO_2632 (O_2632,N_48924,N_49867);
nand UO_2633 (O_2633,N_49883,N_47684);
or UO_2634 (O_2634,N_49265,N_48468);
nor UO_2635 (O_2635,N_49111,N_48104);
and UO_2636 (O_2636,N_49042,N_49618);
xor UO_2637 (O_2637,N_49784,N_48912);
nor UO_2638 (O_2638,N_49309,N_48410);
xnor UO_2639 (O_2639,N_48355,N_47834);
or UO_2640 (O_2640,N_49340,N_49273);
nor UO_2641 (O_2641,N_48107,N_49556);
xor UO_2642 (O_2642,N_49284,N_47997);
nor UO_2643 (O_2643,N_49507,N_49302);
nand UO_2644 (O_2644,N_47642,N_49187);
and UO_2645 (O_2645,N_49650,N_49923);
and UO_2646 (O_2646,N_49603,N_48066);
xor UO_2647 (O_2647,N_47807,N_48843);
or UO_2648 (O_2648,N_49863,N_47880);
or UO_2649 (O_2649,N_49522,N_49822);
xnor UO_2650 (O_2650,N_47759,N_49298);
or UO_2651 (O_2651,N_48688,N_49066);
nand UO_2652 (O_2652,N_49920,N_49967);
xnor UO_2653 (O_2653,N_48091,N_48297);
xnor UO_2654 (O_2654,N_48205,N_49432);
nor UO_2655 (O_2655,N_49093,N_49851);
nand UO_2656 (O_2656,N_49704,N_48290);
and UO_2657 (O_2657,N_49101,N_49860);
or UO_2658 (O_2658,N_47745,N_48998);
nor UO_2659 (O_2659,N_47544,N_49682);
or UO_2660 (O_2660,N_49744,N_49641);
and UO_2661 (O_2661,N_48471,N_48973);
nand UO_2662 (O_2662,N_49122,N_49017);
nor UO_2663 (O_2663,N_49614,N_49254);
and UO_2664 (O_2664,N_47797,N_47847);
or UO_2665 (O_2665,N_48508,N_47514);
or UO_2666 (O_2666,N_48005,N_48406);
nand UO_2667 (O_2667,N_47619,N_48148);
nand UO_2668 (O_2668,N_49319,N_49459);
xnor UO_2669 (O_2669,N_47609,N_48141);
or UO_2670 (O_2670,N_49731,N_49634);
nor UO_2671 (O_2671,N_49517,N_49674);
nand UO_2672 (O_2672,N_47950,N_49461);
nand UO_2673 (O_2673,N_49123,N_49104);
or UO_2674 (O_2674,N_49840,N_48688);
or UO_2675 (O_2675,N_47957,N_49271);
nand UO_2676 (O_2676,N_48178,N_48169);
xnor UO_2677 (O_2677,N_48133,N_49134);
nand UO_2678 (O_2678,N_49862,N_47626);
xnor UO_2679 (O_2679,N_47770,N_49413);
or UO_2680 (O_2680,N_48994,N_49434);
and UO_2681 (O_2681,N_49594,N_49444);
and UO_2682 (O_2682,N_47578,N_47819);
nor UO_2683 (O_2683,N_48800,N_49759);
or UO_2684 (O_2684,N_49276,N_47794);
nor UO_2685 (O_2685,N_49775,N_48008);
xor UO_2686 (O_2686,N_48996,N_48562);
and UO_2687 (O_2687,N_48943,N_49480);
xnor UO_2688 (O_2688,N_48476,N_48321);
xnor UO_2689 (O_2689,N_48123,N_49770);
nor UO_2690 (O_2690,N_47928,N_49246);
nor UO_2691 (O_2691,N_48696,N_49226);
xnor UO_2692 (O_2692,N_48863,N_48183);
and UO_2693 (O_2693,N_47735,N_48987);
xor UO_2694 (O_2694,N_47891,N_48021);
xor UO_2695 (O_2695,N_47978,N_49312);
and UO_2696 (O_2696,N_48144,N_48227);
or UO_2697 (O_2697,N_49066,N_48952);
and UO_2698 (O_2698,N_48697,N_49219);
xor UO_2699 (O_2699,N_49187,N_49732);
xnor UO_2700 (O_2700,N_47781,N_49128);
nand UO_2701 (O_2701,N_49606,N_47583);
xnor UO_2702 (O_2702,N_48392,N_47971);
and UO_2703 (O_2703,N_48247,N_48188);
or UO_2704 (O_2704,N_48831,N_49831);
and UO_2705 (O_2705,N_47885,N_47954);
nand UO_2706 (O_2706,N_48413,N_49263);
xnor UO_2707 (O_2707,N_47729,N_48915);
and UO_2708 (O_2708,N_48897,N_47725);
or UO_2709 (O_2709,N_48113,N_48459);
or UO_2710 (O_2710,N_48061,N_47884);
and UO_2711 (O_2711,N_48981,N_49726);
and UO_2712 (O_2712,N_49530,N_47915);
nand UO_2713 (O_2713,N_49126,N_47684);
nand UO_2714 (O_2714,N_47526,N_49771);
nand UO_2715 (O_2715,N_48810,N_49349);
xnor UO_2716 (O_2716,N_49732,N_49719);
nor UO_2717 (O_2717,N_49702,N_49332);
nor UO_2718 (O_2718,N_49158,N_48077);
xnor UO_2719 (O_2719,N_47780,N_48371);
xor UO_2720 (O_2720,N_49353,N_48164);
nand UO_2721 (O_2721,N_47688,N_49229);
nand UO_2722 (O_2722,N_48556,N_48317);
or UO_2723 (O_2723,N_48541,N_49623);
or UO_2724 (O_2724,N_48200,N_49935);
nand UO_2725 (O_2725,N_49545,N_48697);
xor UO_2726 (O_2726,N_49580,N_48845);
and UO_2727 (O_2727,N_48909,N_48531);
nand UO_2728 (O_2728,N_47751,N_48290);
nor UO_2729 (O_2729,N_49056,N_47603);
xor UO_2730 (O_2730,N_47669,N_49048);
and UO_2731 (O_2731,N_49707,N_49756);
nor UO_2732 (O_2732,N_48725,N_49834);
or UO_2733 (O_2733,N_48223,N_49499);
xor UO_2734 (O_2734,N_47712,N_49699);
and UO_2735 (O_2735,N_49385,N_47648);
or UO_2736 (O_2736,N_48920,N_49076);
nand UO_2737 (O_2737,N_49033,N_48070);
nand UO_2738 (O_2738,N_48750,N_49868);
or UO_2739 (O_2739,N_48344,N_49461);
nor UO_2740 (O_2740,N_49237,N_48426);
or UO_2741 (O_2741,N_48321,N_49301);
nand UO_2742 (O_2742,N_48285,N_48643);
xor UO_2743 (O_2743,N_49401,N_48136);
nand UO_2744 (O_2744,N_49311,N_48449);
nand UO_2745 (O_2745,N_49078,N_47868);
or UO_2746 (O_2746,N_47933,N_47525);
or UO_2747 (O_2747,N_49292,N_49377);
and UO_2748 (O_2748,N_48969,N_47766);
nor UO_2749 (O_2749,N_48462,N_49766);
xnor UO_2750 (O_2750,N_49870,N_48319);
nand UO_2751 (O_2751,N_49842,N_49522);
xor UO_2752 (O_2752,N_49517,N_47779);
nor UO_2753 (O_2753,N_47785,N_48947);
and UO_2754 (O_2754,N_48449,N_49153);
or UO_2755 (O_2755,N_47619,N_48461);
or UO_2756 (O_2756,N_49864,N_47929);
nand UO_2757 (O_2757,N_48460,N_48075);
nand UO_2758 (O_2758,N_48910,N_49978);
nor UO_2759 (O_2759,N_48495,N_49602);
xor UO_2760 (O_2760,N_49000,N_49116);
nor UO_2761 (O_2761,N_48165,N_47862);
xnor UO_2762 (O_2762,N_49612,N_49900);
nand UO_2763 (O_2763,N_49594,N_48502);
or UO_2764 (O_2764,N_48639,N_47872);
or UO_2765 (O_2765,N_48225,N_48841);
nor UO_2766 (O_2766,N_48078,N_48723);
and UO_2767 (O_2767,N_47528,N_49816);
nand UO_2768 (O_2768,N_49668,N_49712);
or UO_2769 (O_2769,N_49831,N_48526);
nor UO_2770 (O_2770,N_48229,N_47939);
nor UO_2771 (O_2771,N_47571,N_48005);
nor UO_2772 (O_2772,N_49446,N_47703);
or UO_2773 (O_2773,N_48350,N_48674);
nand UO_2774 (O_2774,N_47982,N_47810);
xnor UO_2775 (O_2775,N_48486,N_47918);
nor UO_2776 (O_2776,N_49844,N_47579);
nor UO_2777 (O_2777,N_48641,N_49587);
xor UO_2778 (O_2778,N_49598,N_48435);
or UO_2779 (O_2779,N_48554,N_49753);
or UO_2780 (O_2780,N_48840,N_47745);
nor UO_2781 (O_2781,N_49991,N_48503);
nand UO_2782 (O_2782,N_48516,N_49732);
or UO_2783 (O_2783,N_48751,N_49295);
nand UO_2784 (O_2784,N_49106,N_47784);
nand UO_2785 (O_2785,N_47659,N_48282);
xor UO_2786 (O_2786,N_49570,N_48009);
or UO_2787 (O_2787,N_49904,N_48930);
and UO_2788 (O_2788,N_49896,N_48272);
and UO_2789 (O_2789,N_48295,N_47732);
nor UO_2790 (O_2790,N_48200,N_48336);
xor UO_2791 (O_2791,N_49156,N_48371);
nor UO_2792 (O_2792,N_48553,N_48589);
and UO_2793 (O_2793,N_47899,N_48299);
nor UO_2794 (O_2794,N_49583,N_49311);
nand UO_2795 (O_2795,N_47692,N_48153);
or UO_2796 (O_2796,N_48873,N_48836);
nand UO_2797 (O_2797,N_48706,N_48404);
xnor UO_2798 (O_2798,N_47904,N_48046);
nand UO_2799 (O_2799,N_48880,N_49597);
nand UO_2800 (O_2800,N_48748,N_49396);
and UO_2801 (O_2801,N_48056,N_48566);
and UO_2802 (O_2802,N_48775,N_49679);
xnor UO_2803 (O_2803,N_48211,N_48673);
and UO_2804 (O_2804,N_48076,N_47872);
nor UO_2805 (O_2805,N_48840,N_49509);
nor UO_2806 (O_2806,N_48169,N_48026);
or UO_2807 (O_2807,N_48045,N_49777);
nand UO_2808 (O_2808,N_48266,N_49113);
nand UO_2809 (O_2809,N_48292,N_49232);
nor UO_2810 (O_2810,N_49666,N_48498);
and UO_2811 (O_2811,N_48191,N_47588);
xnor UO_2812 (O_2812,N_48816,N_49983);
or UO_2813 (O_2813,N_49102,N_49690);
nor UO_2814 (O_2814,N_49032,N_49434);
nor UO_2815 (O_2815,N_48570,N_49554);
or UO_2816 (O_2816,N_48560,N_49191);
nand UO_2817 (O_2817,N_49967,N_47682);
nand UO_2818 (O_2818,N_48868,N_49390);
or UO_2819 (O_2819,N_48883,N_48386);
xnor UO_2820 (O_2820,N_48496,N_47956);
and UO_2821 (O_2821,N_48144,N_47581);
and UO_2822 (O_2822,N_47752,N_48205);
nor UO_2823 (O_2823,N_47765,N_47549);
nor UO_2824 (O_2824,N_49897,N_47620);
xnor UO_2825 (O_2825,N_49367,N_48297);
xnor UO_2826 (O_2826,N_48963,N_48156);
and UO_2827 (O_2827,N_48738,N_48067);
or UO_2828 (O_2828,N_47850,N_47621);
xor UO_2829 (O_2829,N_49992,N_49561);
nor UO_2830 (O_2830,N_48657,N_49317);
nor UO_2831 (O_2831,N_49207,N_49571);
or UO_2832 (O_2832,N_47517,N_48938);
nand UO_2833 (O_2833,N_48987,N_48670);
or UO_2834 (O_2834,N_49899,N_49662);
nor UO_2835 (O_2835,N_48779,N_49281);
xor UO_2836 (O_2836,N_48578,N_49093);
xor UO_2837 (O_2837,N_48870,N_48365);
or UO_2838 (O_2838,N_49320,N_49832);
xor UO_2839 (O_2839,N_48186,N_49481);
nand UO_2840 (O_2840,N_48159,N_48099);
nand UO_2841 (O_2841,N_47767,N_47544);
and UO_2842 (O_2842,N_49336,N_49267);
or UO_2843 (O_2843,N_47720,N_49322);
nor UO_2844 (O_2844,N_49650,N_48469);
xnor UO_2845 (O_2845,N_47692,N_48910);
xnor UO_2846 (O_2846,N_47608,N_47578);
xor UO_2847 (O_2847,N_48349,N_48557);
nand UO_2848 (O_2848,N_49831,N_48613);
and UO_2849 (O_2849,N_48173,N_47847);
nor UO_2850 (O_2850,N_48130,N_48355);
xnor UO_2851 (O_2851,N_49172,N_48423);
and UO_2852 (O_2852,N_47886,N_48847);
nand UO_2853 (O_2853,N_48828,N_47637);
or UO_2854 (O_2854,N_49787,N_48522);
and UO_2855 (O_2855,N_49310,N_49334);
xor UO_2856 (O_2856,N_48704,N_49660);
nand UO_2857 (O_2857,N_49506,N_49777);
nor UO_2858 (O_2858,N_49540,N_47678);
nand UO_2859 (O_2859,N_49920,N_49433);
and UO_2860 (O_2860,N_49392,N_49524);
nor UO_2861 (O_2861,N_49376,N_48495);
xor UO_2862 (O_2862,N_49890,N_47939);
xnor UO_2863 (O_2863,N_49853,N_48808);
nor UO_2864 (O_2864,N_47755,N_49188);
nand UO_2865 (O_2865,N_49611,N_49100);
or UO_2866 (O_2866,N_48169,N_48190);
and UO_2867 (O_2867,N_48551,N_48548);
nand UO_2868 (O_2868,N_49259,N_49327);
xor UO_2869 (O_2869,N_48465,N_48474);
xnor UO_2870 (O_2870,N_48265,N_49315);
xor UO_2871 (O_2871,N_49516,N_48993);
nand UO_2872 (O_2872,N_49707,N_49373);
nand UO_2873 (O_2873,N_49996,N_47620);
xor UO_2874 (O_2874,N_48998,N_48579);
or UO_2875 (O_2875,N_48572,N_47937);
and UO_2876 (O_2876,N_49918,N_48452);
nand UO_2877 (O_2877,N_49413,N_49979);
nand UO_2878 (O_2878,N_49741,N_47806);
nor UO_2879 (O_2879,N_47575,N_48174);
nand UO_2880 (O_2880,N_49162,N_47585);
or UO_2881 (O_2881,N_49189,N_47659);
and UO_2882 (O_2882,N_49238,N_48236);
and UO_2883 (O_2883,N_47810,N_49862);
or UO_2884 (O_2884,N_47904,N_48624);
nand UO_2885 (O_2885,N_47700,N_49821);
xnor UO_2886 (O_2886,N_49175,N_48631);
nor UO_2887 (O_2887,N_49683,N_48884);
nor UO_2888 (O_2888,N_48016,N_47602);
or UO_2889 (O_2889,N_47955,N_48882);
xor UO_2890 (O_2890,N_48444,N_49916);
or UO_2891 (O_2891,N_48857,N_49688);
xnor UO_2892 (O_2892,N_48908,N_49366);
xnor UO_2893 (O_2893,N_49612,N_48280);
nor UO_2894 (O_2894,N_49121,N_49630);
or UO_2895 (O_2895,N_49211,N_49384);
and UO_2896 (O_2896,N_48790,N_48553);
or UO_2897 (O_2897,N_48107,N_48624);
or UO_2898 (O_2898,N_49243,N_49296);
and UO_2899 (O_2899,N_48788,N_49573);
nand UO_2900 (O_2900,N_48819,N_47661);
nand UO_2901 (O_2901,N_49793,N_48983);
xnor UO_2902 (O_2902,N_48083,N_48189);
xnor UO_2903 (O_2903,N_47996,N_49675);
nor UO_2904 (O_2904,N_48124,N_47514);
xor UO_2905 (O_2905,N_48169,N_47985);
nor UO_2906 (O_2906,N_49391,N_48058);
or UO_2907 (O_2907,N_48051,N_47580);
nor UO_2908 (O_2908,N_48837,N_48915);
or UO_2909 (O_2909,N_49221,N_48625);
or UO_2910 (O_2910,N_48748,N_48015);
and UO_2911 (O_2911,N_47641,N_48566);
xnor UO_2912 (O_2912,N_48350,N_49681);
and UO_2913 (O_2913,N_49252,N_48256);
xor UO_2914 (O_2914,N_48578,N_49143);
nor UO_2915 (O_2915,N_48982,N_48563);
nor UO_2916 (O_2916,N_49882,N_48400);
nor UO_2917 (O_2917,N_48182,N_49239);
nand UO_2918 (O_2918,N_48383,N_48760);
or UO_2919 (O_2919,N_48926,N_48148);
xor UO_2920 (O_2920,N_49080,N_49940);
xor UO_2921 (O_2921,N_48872,N_49901);
and UO_2922 (O_2922,N_47504,N_48712);
nand UO_2923 (O_2923,N_48061,N_48485);
or UO_2924 (O_2924,N_49166,N_48912);
xor UO_2925 (O_2925,N_47782,N_49211);
or UO_2926 (O_2926,N_49337,N_48606);
and UO_2927 (O_2927,N_48814,N_48170);
or UO_2928 (O_2928,N_47930,N_49541);
nand UO_2929 (O_2929,N_49764,N_49392);
nor UO_2930 (O_2930,N_48106,N_47610);
nand UO_2931 (O_2931,N_48184,N_48571);
or UO_2932 (O_2932,N_49754,N_48409);
nand UO_2933 (O_2933,N_48022,N_49561);
nor UO_2934 (O_2934,N_48633,N_47741);
nor UO_2935 (O_2935,N_49869,N_49348);
nand UO_2936 (O_2936,N_49342,N_48945);
nand UO_2937 (O_2937,N_49261,N_49323);
nor UO_2938 (O_2938,N_48750,N_49495);
nor UO_2939 (O_2939,N_49409,N_47586);
or UO_2940 (O_2940,N_49395,N_49229);
and UO_2941 (O_2941,N_49338,N_47618);
nand UO_2942 (O_2942,N_49418,N_49571);
nand UO_2943 (O_2943,N_48304,N_48623);
or UO_2944 (O_2944,N_48026,N_47665);
xnor UO_2945 (O_2945,N_48613,N_48325);
nand UO_2946 (O_2946,N_48506,N_47662);
or UO_2947 (O_2947,N_48477,N_47879);
and UO_2948 (O_2948,N_49901,N_49547);
xor UO_2949 (O_2949,N_49270,N_49501);
nor UO_2950 (O_2950,N_47840,N_48758);
and UO_2951 (O_2951,N_49910,N_49852);
nand UO_2952 (O_2952,N_47509,N_48604);
and UO_2953 (O_2953,N_49811,N_49827);
or UO_2954 (O_2954,N_49547,N_49019);
nand UO_2955 (O_2955,N_48683,N_49161);
nand UO_2956 (O_2956,N_49692,N_49943);
nand UO_2957 (O_2957,N_48111,N_48735);
nand UO_2958 (O_2958,N_49463,N_49664);
nand UO_2959 (O_2959,N_48406,N_49004);
nor UO_2960 (O_2960,N_48759,N_49391);
nor UO_2961 (O_2961,N_48883,N_48292);
nor UO_2962 (O_2962,N_48610,N_48393);
xnor UO_2963 (O_2963,N_49843,N_47856);
or UO_2964 (O_2964,N_47737,N_48539);
or UO_2965 (O_2965,N_49484,N_47972);
nor UO_2966 (O_2966,N_48452,N_48943);
and UO_2967 (O_2967,N_49248,N_49271);
and UO_2968 (O_2968,N_49674,N_48401);
nor UO_2969 (O_2969,N_48875,N_49177);
nor UO_2970 (O_2970,N_48777,N_48652);
nand UO_2971 (O_2971,N_48846,N_48774);
xor UO_2972 (O_2972,N_47892,N_49250);
or UO_2973 (O_2973,N_47760,N_47749);
nor UO_2974 (O_2974,N_47843,N_48016);
nand UO_2975 (O_2975,N_47884,N_48718);
nor UO_2976 (O_2976,N_47858,N_49314);
nor UO_2977 (O_2977,N_48306,N_47573);
nor UO_2978 (O_2978,N_48966,N_49849);
and UO_2979 (O_2979,N_49274,N_49017);
and UO_2980 (O_2980,N_48213,N_49581);
nor UO_2981 (O_2981,N_49212,N_47527);
xnor UO_2982 (O_2982,N_49298,N_49636);
or UO_2983 (O_2983,N_49102,N_47554);
nand UO_2984 (O_2984,N_48460,N_49464);
or UO_2985 (O_2985,N_47581,N_48555);
nand UO_2986 (O_2986,N_47891,N_49137);
or UO_2987 (O_2987,N_47813,N_49591);
xnor UO_2988 (O_2988,N_49654,N_48108);
or UO_2989 (O_2989,N_48792,N_48286);
and UO_2990 (O_2990,N_49995,N_47858);
nor UO_2991 (O_2991,N_48082,N_49356);
nand UO_2992 (O_2992,N_48562,N_48578);
or UO_2993 (O_2993,N_47909,N_48085);
or UO_2994 (O_2994,N_47685,N_48971);
or UO_2995 (O_2995,N_47882,N_48247);
nor UO_2996 (O_2996,N_49835,N_47815);
xor UO_2997 (O_2997,N_48121,N_48240);
nor UO_2998 (O_2998,N_49679,N_47646);
nor UO_2999 (O_2999,N_49101,N_49537);
nor UO_3000 (O_3000,N_49628,N_47519);
xnor UO_3001 (O_3001,N_49861,N_48944);
nand UO_3002 (O_3002,N_47865,N_47916);
and UO_3003 (O_3003,N_47517,N_48865);
or UO_3004 (O_3004,N_49054,N_48367);
nor UO_3005 (O_3005,N_49279,N_47642);
xor UO_3006 (O_3006,N_48889,N_49578);
nand UO_3007 (O_3007,N_48065,N_48973);
or UO_3008 (O_3008,N_49411,N_48140);
or UO_3009 (O_3009,N_48932,N_48408);
or UO_3010 (O_3010,N_49978,N_48883);
xor UO_3011 (O_3011,N_48209,N_47718);
or UO_3012 (O_3012,N_49431,N_48662);
nor UO_3013 (O_3013,N_48307,N_48259);
nor UO_3014 (O_3014,N_48577,N_48237);
xnor UO_3015 (O_3015,N_48563,N_47723);
nor UO_3016 (O_3016,N_49243,N_48906);
nand UO_3017 (O_3017,N_47855,N_48762);
xnor UO_3018 (O_3018,N_48106,N_49771);
nor UO_3019 (O_3019,N_48913,N_48843);
nor UO_3020 (O_3020,N_48479,N_47848);
or UO_3021 (O_3021,N_47932,N_48494);
or UO_3022 (O_3022,N_49154,N_48187);
nand UO_3023 (O_3023,N_49320,N_47549);
nand UO_3024 (O_3024,N_49084,N_49865);
or UO_3025 (O_3025,N_49596,N_49514);
nand UO_3026 (O_3026,N_47926,N_49381);
and UO_3027 (O_3027,N_49115,N_49482);
nand UO_3028 (O_3028,N_47785,N_49974);
and UO_3029 (O_3029,N_48461,N_48574);
xor UO_3030 (O_3030,N_49393,N_47828);
or UO_3031 (O_3031,N_47990,N_48064);
nand UO_3032 (O_3032,N_49914,N_48837);
and UO_3033 (O_3033,N_49278,N_48083);
nor UO_3034 (O_3034,N_49668,N_48638);
or UO_3035 (O_3035,N_47723,N_48878);
nor UO_3036 (O_3036,N_49791,N_48424);
nor UO_3037 (O_3037,N_48667,N_48946);
and UO_3038 (O_3038,N_48794,N_49979);
or UO_3039 (O_3039,N_48077,N_49768);
xnor UO_3040 (O_3040,N_48269,N_49471);
xnor UO_3041 (O_3041,N_48671,N_48020);
nand UO_3042 (O_3042,N_48246,N_47674);
nor UO_3043 (O_3043,N_47780,N_49502);
xnor UO_3044 (O_3044,N_48540,N_48184);
xor UO_3045 (O_3045,N_48981,N_48768);
xor UO_3046 (O_3046,N_47917,N_49013);
nand UO_3047 (O_3047,N_49431,N_49539);
nor UO_3048 (O_3048,N_48110,N_49815);
and UO_3049 (O_3049,N_48711,N_49647);
xor UO_3050 (O_3050,N_49337,N_48404);
xnor UO_3051 (O_3051,N_48436,N_48387);
xnor UO_3052 (O_3052,N_48938,N_49321);
and UO_3053 (O_3053,N_48566,N_48317);
nand UO_3054 (O_3054,N_48563,N_48649);
and UO_3055 (O_3055,N_48579,N_49985);
nor UO_3056 (O_3056,N_48410,N_47897);
or UO_3057 (O_3057,N_48218,N_48718);
nand UO_3058 (O_3058,N_48490,N_49995);
nand UO_3059 (O_3059,N_49426,N_48011);
xor UO_3060 (O_3060,N_49851,N_49070);
nor UO_3061 (O_3061,N_49549,N_48211);
and UO_3062 (O_3062,N_48456,N_49278);
nand UO_3063 (O_3063,N_49600,N_48210);
or UO_3064 (O_3064,N_49787,N_47883);
and UO_3065 (O_3065,N_47753,N_48790);
nor UO_3066 (O_3066,N_47627,N_49552);
xor UO_3067 (O_3067,N_47790,N_48456);
or UO_3068 (O_3068,N_48384,N_49190);
nand UO_3069 (O_3069,N_49044,N_49888);
and UO_3070 (O_3070,N_48581,N_48575);
or UO_3071 (O_3071,N_48771,N_49889);
xnor UO_3072 (O_3072,N_47604,N_48538);
nand UO_3073 (O_3073,N_49193,N_49143);
and UO_3074 (O_3074,N_49204,N_49877);
nor UO_3075 (O_3075,N_48348,N_49882);
or UO_3076 (O_3076,N_47506,N_49266);
and UO_3077 (O_3077,N_49616,N_47582);
nor UO_3078 (O_3078,N_48083,N_48902);
nor UO_3079 (O_3079,N_48566,N_48348);
or UO_3080 (O_3080,N_48283,N_49453);
xnor UO_3081 (O_3081,N_48299,N_48811);
or UO_3082 (O_3082,N_49586,N_47517);
nand UO_3083 (O_3083,N_49835,N_48944);
or UO_3084 (O_3084,N_49395,N_48114);
or UO_3085 (O_3085,N_48434,N_48384);
xnor UO_3086 (O_3086,N_48665,N_49624);
and UO_3087 (O_3087,N_49971,N_48756);
xor UO_3088 (O_3088,N_49032,N_47978);
nand UO_3089 (O_3089,N_48433,N_49780);
xnor UO_3090 (O_3090,N_49723,N_47646);
nand UO_3091 (O_3091,N_48322,N_49110);
nor UO_3092 (O_3092,N_47976,N_47924);
and UO_3093 (O_3093,N_49282,N_47838);
nor UO_3094 (O_3094,N_48614,N_47665);
and UO_3095 (O_3095,N_49205,N_48633);
nor UO_3096 (O_3096,N_48921,N_49389);
nor UO_3097 (O_3097,N_48790,N_49046);
nand UO_3098 (O_3098,N_48635,N_48615);
and UO_3099 (O_3099,N_48136,N_48428);
nor UO_3100 (O_3100,N_49770,N_48063);
xor UO_3101 (O_3101,N_49174,N_49582);
nand UO_3102 (O_3102,N_48621,N_49024);
and UO_3103 (O_3103,N_47541,N_49758);
xnor UO_3104 (O_3104,N_47894,N_48307);
nor UO_3105 (O_3105,N_48789,N_48783);
nand UO_3106 (O_3106,N_48405,N_49951);
or UO_3107 (O_3107,N_49747,N_48713);
nor UO_3108 (O_3108,N_47504,N_48954);
xnor UO_3109 (O_3109,N_47975,N_49513);
xor UO_3110 (O_3110,N_49530,N_48181);
nand UO_3111 (O_3111,N_47678,N_47818);
xor UO_3112 (O_3112,N_48591,N_49015);
nand UO_3113 (O_3113,N_48922,N_49679);
or UO_3114 (O_3114,N_48479,N_49409);
nand UO_3115 (O_3115,N_48486,N_49950);
nor UO_3116 (O_3116,N_49100,N_48864);
and UO_3117 (O_3117,N_47868,N_48807);
nor UO_3118 (O_3118,N_48849,N_48537);
nand UO_3119 (O_3119,N_47525,N_48308);
nor UO_3120 (O_3120,N_48314,N_49088);
nand UO_3121 (O_3121,N_49515,N_48809);
nand UO_3122 (O_3122,N_48380,N_48196);
or UO_3123 (O_3123,N_47843,N_47839);
nor UO_3124 (O_3124,N_49889,N_48352);
nand UO_3125 (O_3125,N_49783,N_47744);
and UO_3126 (O_3126,N_49280,N_49833);
nand UO_3127 (O_3127,N_48237,N_47543);
nor UO_3128 (O_3128,N_47624,N_49255);
and UO_3129 (O_3129,N_47863,N_47579);
nor UO_3130 (O_3130,N_47571,N_47636);
nor UO_3131 (O_3131,N_48015,N_48998);
and UO_3132 (O_3132,N_49490,N_49054);
or UO_3133 (O_3133,N_48793,N_48453);
or UO_3134 (O_3134,N_49228,N_49749);
and UO_3135 (O_3135,N_47956,N_48974);
and UO_3136 (O_3136,N_49352,N_48398);
xnor UO_3137 (O_3137,N_48896,N_49459);
or UO_3138 (O_3138,N_49954,N_49598);
nor UO_3139 (O_3139,N_49762,N_49031);
or UO_3140 (O_3140,N_47654,N_47622);
and UO_3141 (O_3141,N_49593,N_48477);
nand UO_3142 (O_3142,N_48664,N_47532);
and UO_3143 (O_3143,N_49479,N_48474);
xnor UO_3144 (O_3144,N_49615,N_48786);
and UO_3145 (O_3145,N_48386,N_48302);
or UO_3146 (O_3146,N_48829,N_49828);
nor UO_3147 (O_3147,N_49586,N_48830);
nand UO_3148 (O_3148,N_48158,N_48831);
nor UO_3149 (O_3149,N_48944,N_47833);
or UO_3150 (O_3150,N_48404,N_49281);
nor UO_3151 (O_3151,N_49871,N_48569);
nand UO_3152 (O_3152,N_48653,N_49354);
nand UO_3153 (O_3153,N_47892,N_48343);
nand UO_3154 (O_3154,N_49309,N_49313);
nand UO_3155 (O_3155,N_47934,N_49679);
nand UO_3156 (O_3156,N_47796,N_49335);
xnor UO_3157 (O_3157,N_47657,N_49128);
or UO_3158 (O_3158,N_47564,N_48770);
or UO_3159 (O_3159,N_48571,N_49934);
nand UO_3160 (O_3160,N_49850,N_47931);
nor UO_3161 (O_3161,N_48143,N_49002);
and UO_3162 (O_3162,N_47668,N_47915);
or UO_3163 (O_3163,N_48804,N_49561);
nor UO_3164 (O_3164,N_48787,N_49704);
xor UO_3165 (O_3165,N_47590,N_47609);
xnor UO_3166 (O_3166,N_48054,N_48635);
or UO_3167 (O_3167,N_48060,N_49921);
and UO_3168 (O_3168,N_49652,N_49658);
and UO_3169 (O_3169,N_48660,N_48481);
nor UO_3170 (O_3170,N_48712,N_48574);
or UO_3171 (O_3171,N_49738,N_47987);
nor UO_3172 (O_3172,N_47769,N_48557);
nand UO_3173 (O_3173,N_48282,N_48509);
and UO_3174 (O_3174,N_47827,N_47940);
xor UO_3175 (O_3175,N_48525,N_48405);
nor UO_3176 (O_3176,N_48214,N_49991);
nor UO_3177 (O_3177,N_48297,N_48945);
and UO_3178 (O_3178,N_49350,N_49089);
nand UO_3179 (O_3179,N_47549,N_48879);
nor UO_3180 (O_3180,N_49141,N_47961);
nand UO_3181 (O_3181,N_48381,N_47614);
xor UO_3182 (O_3182,N_49908,N_48911);
xor UO_3183 (O_3183,N_48143,N_48465);
and UO_3184 (O_3184,N_48103,N_48927);
and UO_3185 (O_3185,N_48785,N_47758);
xor UO_3186 (O_3186,N_48585,N_49363);
xor UO_3187 (O_3187,N_49712,N_49655);
nor UO_3188 (O_3188,N_48321,N_47837);
and UO_3189 (O_3189,N_49415,N_49138);
nand UO_3190 (O_3190,N_47594,N_48978);
and UO_3191 (O_3191,N_48244,N_49126);
nand UO_3192 (O_3192,N_49222,N_48222);
nand UO_3193 (O_3193,N_48635,N_49880);
xor UO_3194 (O_3194,N_47766,N_48539);
or UO_3195 (O_3195,N_47641,N_48255);
nor UO_3196 (O_3196,N_49214,N_48150);
nor UO_3197 (O_3197,N_49151,N_48208);
or UO_3198 (O_3198,N_48203,N_49758);
or UO_3199 (O_3199,N_48866,N_48337);
and UO_3200 (O_3200,N_48275,N_48880);
and UO_3201 (O_3201,N_47788,N_47610);
nor UO_3202 (O_3202,N_49223,N_48962);
xor UO_3203 (O_3203,N_48530,N_49772);
or UO_3204 (O_3204,N_49452,N_49081);
xnor UO_3205 (O_3205,N_47694,N_49990);
xnor UO_3206 (O_3206,N_48454,N_49742);
nor UO_3207 (O_3207,N_48730,N_47634);
nand UO_3208 (O_3208,N_48206,N_49791);
or UO_3209 (O_3209,N_48923,N_48611);
nor UO_3210 (O_3210,N_49361,N_48954);
nand UO_3211 (O_3211,N_48744,N_49348);
xnor UO_3212 (O_3212,N_49738,N_47841);
nor UO_3213 (O_3213,N_49932,N_47774);
nor UO_3214 (O_3214,N_48329,N_47826);
nor UO_3215 (O_3215,N_48153,N_48926);
nor UO_3216 (O_3216,N_48120,N_49587);
xnor UO_3217 (O_3217,N_49097,N_48521);
and UO_3218 (O_3218,N_48562,N_47980);
nor UO_3219 (O_3219,N_48827,N_48802);
or UO_3220 (O_3220,N_49570,N_49279);
and UO_3221 (O_3221,N_49886,N_47953);
xor UO_3222 (O_3222,N_48801,N_47602);
nor UO_3223 (O_3223,N_49075,N_49721);
xor UO_3224 (O_3224,N_48678,N_48824);
and UO_3225 (O_3225,N_48169,N_49477);
nand UO_3226 (O_3226,N_47730,N_48748);
nor UO_3227 (O_3227,N_49139,N_48880);
nand UO_3228 (O_3228,N_48960,N_47563);
xnor UO_3229 (O_3229,N_48146,N_49208);
nor UO_3230 (O_3230,N_49585,N_49519);
and UO_3231 (O_3231,N_49506,N_48173);
nor UO_3232 (O_3232,N_49965,N_47605);
xnor UO_3233 (O_3233,N_48431,N_48705);
xor UO_3234 (O_3234,N_49651,N_49453);
nand UO_3235 (O_3235,N_48092,N_48234);
and UO_3236 (O_3236,N_49802,N_49299);
xor UO_3237 (O_3237,N_49121,N_49492);
or UO_3238 (O_3238,N_47722,N_47979);
xnor UO_3239 (O_3239,N_48704,N_48591);
or UO_3240 (O_3240,N_47667,N_49205);
or UO_3241 (O_3241,N_49534,N_49276);
nor UO_3242 (O_3242,N_49362,N_48835);
nor UO_3243 (O_3243,N_49569,N_49494);
or UO_3244 (O_3244,N_48577,N_48223);
nand UO_3245 (O_3245,N_49463,N_47639);
nor UO_3246 (O_3246,N_49501,N_47624);
nand UO_3247 (O_3247,N_47796,N_48865);
nor UO_3248 (O_3248,N_49611,N_47839);
nand UO_3249 (O_3249,N_48474,N_49209);
nor UO_3250 (O_3250,N_49610,N_48643);
and UO_3251 (O_3251,N_47968,N_48314);
nand UO_3252 (O_3252,N_49811,N_47892);
nor UO_3253 (O_3253,N_48615,N_49719);
nand UO_3254 (O_3254,N_47868,N_47645);
xnor UO_3255 (O_3255,N_48566,N_48478);
or UO_3256 (O_3256,N_49998,N_47501);
and UO_3257 (O_3257,N_49658,N_48815);
xor UO_3258 (O_3258,N_47530,N_48747);
or UO_3259 (O_3259,N_49988,N_48044);
nand UO_3260 (O_3260,N_48077,N_47526);
or UO_3261 (O_3261,N_48823,N_48668);
or UO_3262 (O_3262,N_49724,N_48296);
and UO_3263 (O_3263,N_48919,N_48370);
or UO_3264 (O_3264,N_48711,N_47622);
or UO_3265 (O_3265,N_48107,N_47936);
or UO_3266 (O_3266,N_47998,N_48827);
nor UO_3267 (O_3267,N_49265,N_48428);
nor UO_3268 (O_3268,N_48834,N_48121);
xnor UO_3269 (O_3269,N_48867,N_47830);
nor UO_3270 (O_3270,N_48565,N_49774);
xnor UO_3271 (O_3271,N_48991,N_49002);
nand UO_3272 (O_3272,N_49571,N_49074);
and UO_3273 (O_3273,N_49993,N_49257);
xnor UO_3274 (O_3274,N_48404,N_47817);
xor UO_3275 (O_3275,N_48116,N_48819);
or UO_3276 (O_3276,N_49867,N_47981);
and UO_3277 (O_3277,N_48968,N_49299);
xor UO_3278 (O_3278,N_49726,N_47882);
nor UO_3279 (O_3279,N_47796,N_49040);
and UO_3280 (O_3280,N_47629,N_49265);
or UO_3281 (O_3281,N_47639,N_49251);
and UO_3282 (O_3282,N_48586,N_48971);
or UO_3283 (O_3283,N_49368,N_47647);
xor UO_3284 (O_3284,N_47791,N_48607);
xor UO_3285 (O_3285,N_49465,N_49511);
nand UO_3286 (O_3286,N_47847,N_48860);
xor UO_3287 (O_3287,N_47661,N_49203);
and UO_3288 (O_3288,N_48759,N_49469);
nor UO_3289 (O_3289,N_49377,N_49566);
nand UO_3290 (O_3290,N_49648,N_49379);
xor UO_3291 (O_3291,N_48002,N_49236);
xor UO_3292 (O_3292,N_49409,N_49351);
and UO_3293 (O_3293,N_48770,N_47558);
or UO_3294 (O_3294,N_48513,N_49437);
and UO_3295 (O_3295,N_49579,N_48762);
nand UO_3296 (O_3296,N_49814,N_49827);
xnor UO_3297 (O_3297,N_47986,N_49562);
nor UO_3298 (O_3298,N_49822,N_48766);
nor UO_3299 (O_3299,N_49042,N_47783);
xnor UO_3300 (O_3300,N_49689,N_48831);
and UO_3301 (O_3301,N_47578,N_49608);
xor UO_3302 (O_3302,N_47968,N_49346);
or UO_3303 (O_3303,N_49599,N_48625);
and UO_3304 (O_3304,N_49831,N_48856);
nor UO_3305 (O_3305,N_49001,N_49861);
xor UO_3306 (O_3306,N_48096,N_47805);
and UO_3307 (O_3307,N_48746,N_47502);
and UO_3308 (O_3308,N_48032,N_47572);
xor UO_3309 (O_3309,N_49817,N_48419);
xnor UO_3310 (O_3310,N_48430,N_48003);
nand UO_3311 (O_3311,N_49154,N_47960);
or UO_3312 (O_3312,N_49173,N_48124);
nor UO_3313 (O_3313,N_48066,N_48653);
nor UO_3314 (O_3314,N_48210,N_48566);
and UO_3315 (O_3315,N_47598,N_49558);
nor UO_3316 (O_3316,N_49559,N_48932);
nor UO_3317 (O_3317,N_49511,N_48374);
nand UO_3318 (O_3318,N_47726,N_49395);
xnor UO_3319 (O_3319,N_48878,N_49934);
or UO_3320 (O_3320,N_48428,N_48490);
nand UO_3321 (O_3321,N_48857,N_48685);
and UO_3322 (O_3322,N_47789,N_48261);
xor UO_3323 (O_3323,N_49204,N_49221);
nor UO_3324 (O_3324,N_47530,N_47778);
and UO_3325 (O_3325,N_49483,N_48041);
and UO_3326 (O_3326,N_48031,N_48024);
nor UO_3327 (O_3327,N_48857,N_48879);
and UO_3328 (O_3328,N_48803,N_48858);
xnor UO_3329 (O_3329,N_48675,N_49336);
nand UO_3330 (O_3330,N_49693,N_48701);
and UO_3331 (O_3331,N_48902,N_49540);
and UO_3332 (O_3332,N_48997,N_48703);
nor UO_3333 (O_3333,N_47598,N_49210);
or UO_3334 (O_3334,N_48486,N_49369);
and UO_3335 (O_3335,N_49294,N_49522);
and UO_3336 (O_3336,N_49047,N_49338);
nand UO_3337 (O_3337,N_47781,N_47971);
xnor UO_3338 (O_3338,N_47597,N_48714);
and UO_3339 (O_3339,N_49401,N_47953);
nand UO_3340 (O_3340,N_48791,N_48025);
nor UO_3341 (O_3341,N_48543,N_48612);
xnor UO_3342 (O_3342,N_48211,N_49063);
nor UO_3343 (O_3343,N_49949,N_48871);
and UO_3344 (O_3344,N_47940,N_48677);
and UO_3345 (O_3345,N_48475,N_47928);
or UO_3346 (O_3346,N_49584,N_49019);
or UO_3347 (O_3347,N_49703,N_49758);
and UO_3348 (O_3348,N_48999,N_48549);
or UO_3349 (O_3349,N_49473,N_48882);
xor UO_3350 (O_3350,N_48843,N_47685);
nor UO_3351 (O_3351,N_48314,N_48930);
or UO_3352 (O_3352,N_47574,N_48237);
xnor UO_3353 (O_3353,N_48723,N_49167);
xor UO_3354 (O_3354,N_49382,N_49379);
nand UO_3355 (O_3355,N_47779,N_49111);
nor UO_3356 (O_3356,N_49119,N_48740);
or UO_3357 (O_3357,N_48118,N_49358);
nand UO_3358 (O_3358,N_48792,N_47954);
and UO_3359 (O_3359,N_48281,N_49563);
nor UO_3360 (O_3360,N_49026,N_48082);
or UO_3361 (O_3361,N_49177,N_49577);
or UO_3362 (O_3362,N_49803,N_48829);
nand UO_3363 (O_3363,N_48147,N_49122);
or UO_3364 (O_3364,N_49930,N_48860);
nand UO_3365 (O_3365,N_49618,N_48745);
and UO_3366 (O_3366,N_48734,N_48178);
or UO_3367 (O_3367,N_47592,N_48452);
xnor UO_3368 (O_3368,N_48927,N_48515);
and UO_3369 (O_3369,N_48201,N_49845);
nor UO_3370 (O_3370,N_48148,N_47711);
xor UO_3371 (O_3371,N_47811,N_48265);
nor UO_3372 (O_3372,N_48533,N_49678);
nand UO_3373 (O_3373,N_49396,N_47530);
nor UO_3374 (O_3374,N_49707,N_49784);
xnor UO_3375 (O_3375,N_48825,N_49848);
nor UO_3376 (O_3376,N_48809,N_49865);
and UO_3377 (O_3377,N_48768,N_49217);
xor UO_3378 (O_3378,N_48103,N_49503);
nand UO_3379 (O_3379,N_48837,N_49483);
nand UO_3380 (O_3380,N_47769,N_49822);
nor UO_3381 (O_3381,N_48255,N_47539);
nor UO_3382 (O_3382,N_47762,N_49441);
nand UO_3383 (O_3383,N_49099,N_49320);
nand UO_3384 (O_3384,N_48502,N_47884);
nor UO_3385 (O_3385,N_48702,N_49426);
and UO_3386 (O_3386,N_48365,N_49201);
nor UO_3387 (O_3387,N_47900,N_48647);
nand UO_3388 (O_3388,N_47893,N_48932);
nand UO_3389 (O_3389,N_49266,N_48773);
nand UO_3390 (O_3390,N_49342,N_49507);
or UO_3391 (O_3391,N_48849,N_47832);
or UO_3392 (O_3392,N_48553,N_49218);
nand UO_3393 (O_3393,N_49888,N_48455);
xor UO_3394 (O_3394,N_48766,N_49741);
or UO_3395 (O_3395,N_47607,N_48403);
and UO_3396 (O_3396,N_49045,N_48150);
nor UO_3397 (O_3397,N_48038,N_48763);
xnor UO_3398 (O_3398,N_49185,N_47803);
nand UO_3399 (O_3399,N_49956,N_48998);
xnor UO_3400 (O_3400,N_47571,N_49455);
xor UO_3401 (O_3401,N_47765,N_49741);
and UO_3402 (O_3402,N_48293,N_48032);
and UO_3403 (O_3403,N_48650,N_48815);
xnor UO_3404 (O_3404,N_49389,N_48359);
nor UO_3405 (O_3405,N_49537,N_49645);
nand UO_3406 (O_3406,N_49090,N_49468);
or UO_3407 (O_3407,N_49613,N_47766);
nand UO_3408 (O_3408,N_48102,N_49422);
nand UO_3409 (O_3409,N_49036,N_49691);
and UO_3410 (O_3410,N_47768,N_48023);
xor UO_3411 (O_3411,N_49683,N_49182);
or UO_3412 (O_3412,N_48874,N_47817);
nor UO_3413 (O_3413,N_49615,N_49419);
and UO_3414 (O_3414,N_48343,N_49855);
nand UO_3415 (O_3415,N_48939,N_48849);
xnor UO_3416 (O_3416,N_49607,N_49325);
or UO_3417 (O_3417,N_48497,N_49509);
nand UO_3418 (O_3418,N_47649,N_48602);
or UO_3419 (O_3419,N_48031,N_48943);
or UO_3420 (O_3420,N_49548,N_49322);
or UO_3421 (O_3421,N_47827,N_47917);
and UO_3422 (O_3422,N_49274,N_48816);
nand UO_3423 (O_3423,N_49238,N_48244);
xor UO_3424 (O_3424,N_48827,N_48144);
and UO_3425 (O_3425,N_48969,N_48691);
xor UO_3426 (O_3426,N_49189,N_48457);
nand UO_3427 (O_3427,N_47763,N_49670);
and UO_3428 (O_3428,N_48823,N_49652);
and UO_3429 (O_3429,N_47693,N_47731);
nand UO_3430 (O_3430,N_49382,N_47678);
nor UO_3431 (O_3431,N_49839,N_48942);
nand UO_3432 (O_3432,N_47997,N_47514);
and UO_3433 (O_3433,N_49501,N_49059);
xnor UO_3434 (O_3434,N_49320,N_47527);
nand UO_3435 (O_3435,N_47759,N_49354);
and UO_3436 (O_3436,N_49362,N_48860);
nand UO_3437 (O_3437,N_48951,N_49265);
and UO_3438 (O_3438,N_47646,N_49709);
nor UO_3439 (O_3439,N_47721,N_48970);
or UO_3440 (O_3440,N_49218,N_47513);
nor UO_3441 (O_3441,N_49099,N_49120);
and UO_3442 (O_3442,N_47752,N_49844);
nor UO_3443 (O_3443,N_48463,N_49616);
xor UO_3444 (O_3444,N_48575,N_48674);
xnor UO_3445 (O_3445,N_48702,N_49915);
or UO_3446 (O_3446,N_49652,N_48728);
nand UO_3447 (O_3447,N_48830,N_49277);
nor UO_3448 (O_3448,N_48343,N_49171);
nor UO_3449 (O_3449,N_49869,N_47901);
nand UO_3450 (O_3450,N_49738,N_48150);
or UO_3451 (O_3451,N_47570,N_48545);
nand UO_3452 (O_3452,N_48395,N_49100);
or UO_3453 (O_3453,N_49437,N_49007);
xnor UO_3454 (O_3454,N_48291,N_48272);
and UO_3455 (O_3455,N_49513,N_47595);
or UO_3456 (O_3456,N_48733,N_49662);
or UO_3457 (O_3457,N_48607,N_49228);
nand UO_3458 (O_3458,N_48511,N_49464);
nor UO_3459 (O_3459,N_49151,N_48779);
or UO_3460 (O_3460,N_49945,N_49210);
nand UO_3461 (O_3461,N_49724,N_48989);
nand UO_3462 (O_3462,N_48746,N_48444);
xnor UO_3463 (O_3463,N_49559,N_48442);
and UO_3464 (O_3464,N_47732,N_48335);
xor UO_3465 (O_3465,N_49103,N_47668);
nor UO_3466 (O_3466,N_48204,N_48487);
xnor UO_3467 (O_3467,N_49836,N_48635);
nand UO_3468 (O_3468,N_49103,N_48818);
and UO_3469 (O_3469,N_48379,N_48776);
and UO_3470 (O_3470,N_48594,N_49497);
or UO_3471 (O_3471,N_49819,N_47962);
nand UO_3472 (O_3472,N_48304,N_48811);
or UO_3473 (O_3473,N_47641,N_49560);
or UO_3474 (O_3474,N_47833,N_48908);
and UO_3475 (O_3475,N_48247,N_48002);
xor UO_3476 (O_3476,N_49169,N_48851);
nor UO_3477 (O_3477,N_48272,N_49225);
xnor UO_3478 (O_3478,N_47976,N_49376);
nor UO_3479 (O_3479,N_48165,N_49990);
xor UO_3480 (O_3480,N_49582,N_49108);
nor UO_3481 (O_3481,N_48962,N_49353);
and UO_3482 (O_3482,N_48331,N_48543);
and UO_3483 (O_3483,N_48614,N_48469);
xor UO_3484 (O_3484,N_48356,N_47950);
nand UO_3485 (O_3485,N_49192,N_48657);
nand UO_3486 (O_3486,N_49215,N_47584);
nand UO_3487 (O_3487,N_49175,N_47778);
and UO_3488 (O_3488,N_48738,N_49487);
nand UO_3489 (O_3489,N_48132,N_47535);
and UO_3490 (O_3490,N_48683,N_49829);
nor UO_3491 (O_3491,N_49721,N_48197);
and UO_3492 (O_3492,N_49787,N_47924);
nand UO_3493 (O_3493,N_49080,N_48728);
xor UO_3494 (O_3494,N_49768,N_48758);
and UO_3495 (O_3495,N_48673,N_49460);
and UO_3496 (O_3496,N_49622,N_49751);
and UO_3497 (O_3497,N_48339,N_47898);
nand UO_3498 (O_3498,N_48927,N_49673);
and UO_3499 (O_3499,N_48413,N_49594);
nand UO_3500 (O_3500,N_47707,N_49018);
nand UO_3501 (O_3501,N_49016,N_48013);
xor UO_3502 (O_3502,N_49836,N_48845);
or UO_3503 (O_3503,N_48924,N_48614);
nand UO_3504 (O_3504,N_47553,N_49525);
or UO_3505 (O_3505,N_48339,N_49364);
or UO_3506 (O_3506,N_49800,N_48054);
xor UO_3507 (O_3507,N_48564,N_49966);
and UO_3508 (O_3508,N_48092,N_49075);
xnor UO_3509 (O_3509,N_49833,N_48738);
xnor UO_3510 (O_3510,N_49738,N_48153);
nand UO_3511 (O_3511,N_49137,N_48373);
nor UO_3512 (O_3512,N_49465,N_48499);
nor UO_3513 (O_3513,N_48202,N_49673);
nor UO_3514 (O_3514,N_48569,N_48230);
xor UO_3515 (O_3515,N_49791,N_48067);
and UO_3516 (O_3516,N_48907,N_49401);
or UO_3517 (O_3517,N_48315,N_48941);
nand UO_3518 (O_3518,N_47906,N_48484);
nand UO_3519 (O_3519,N_48189,N_49425);
nor UO_3520 (O_3520,N_48283,N_49866);
xnor UO_3521 (O_3521,N_48229,N_49140);
and UO_3522 (O_3522,N_49609,N_49896);
nand UO_3523 (O_3523,N_49605,N_49140);
nand UO_3524 (O_3524,N_47962,N_47718);
nand UO_3525 (O_3525,N_49237,N_48286);
or UO_3526 (O_3526,N_49583,N_47622);
and UO_3527 (O_3527,N_48128,N_48088);
nor UO_3528 (O_3528,N_49370,N_49899);
xor UO_3529 (O_3529,N_47628,N_48459);
nand UO_3530 (O_3530,N_49235,N_49756);
nor UO_3531 (O_3531,N_47675,N_49456);
and UO_3532 (O_3532,N_48668,N_49124);
and UO_3533 (O_3533,N_49705,N_49031);
nor UO_3534 (O_3534,N_49366,N_49245);
or UO_3535 (O_3535,N_49153,N_49186);
nor UO_3536 (O_3536,N_49618,N_48168);
nand UO_3537 (O_3537,N_48526,N_48046);
or UO_3538 (O_3538,N_49044,N_49846);
and UO_3539 (O_3539,N_49459,N_48152);
nor UO_3540 (O_3540,N_48942,N_47655);
or UO_3541 (O_3541,N_49047,N_49919);
xor UO_3542 (O_3542,N_48853,N_49367);
and UO_3543 (O_3543,N_47601,N_48532);
nand UO_3544 (O_3544,N_49424,N_48878);
and UO_3545 (O_3545,N_48691,N_48513);
nand UO_3546 (O_3546,N_49844,N_49108);
or UO_3547 (O_3547,N_47855,N_48837);
nor UO_3548 (O_3548,N_49573,N_48542);
nand UO_3549 (O_3549,N_49038,N_49830);
nor UO_3550 (O_3550,N_48512,N_49087);
xnor UO_3551 (O_3551,N_48203,N_47599);
nand UO_3552 (O_3552,N_48933,N_47958);
nor UO_3553 (O_3553,N_48450,N_48884);
xnor UO_3554 (O_3554,N_49146,N_47788);
nand UO_3555 (O_3555,N_48409,N_48534);
or UO_3556 (O_3556,N_48838,N_49562);
xor UO_3557 (O_3557,N_47512,N_47596);
xor UO_3558 (O_3558,N_49023,N_49475);
nand UO_3559 (O_3559,N_48516,N_49559);
nor UO_3560 (O_3560,N_48804,N_49809);
xor UO_3561 (O_3561,N_48893,N_48529);
xnor UO_3562 (O_3562,N_49653,N_48543);
xor UO_3563 (O_3563,N_49077,N_49345);
nand UO_3564 (O_3564,N_49372,N_49330);
or UO_3565 (O_3565,N_48061,N_49373);
and UO_3566 (O_3566,N_49304,N_49877);
or UO_3567 (O_3567,N_47603,N_47664);
xnor UO_3568 (O_3568,N_47723,N_47984);
or UO_3569 (O_3569,N_47633,N_49306);
nor UO_3570 (O_3570,N_47949,N_49116);
or UO_3571 (O_3571,N_48212,N_49806);
xnor UO_3572 (O_3572,N_49011,N_49129);
or UO_3573 (O_3573,N_47823,N_49950);
and UO_3574 (O_3574,N_48912,N_49229);
nand UO_3575 (O_3575,N_48402,N_48384);
xor UO_3576 (O_3576,N_49638,N_48230);
nand UO_3577 (O_3577,N_48121,N_48576);
nand UO_3578 (O_3578,N_48944,N_49950);
and UO_3579 (O_3579,N_48977,N_47887);
and UO_3580 (O_3580,N_48783,N_49101);
or UO_3581 (O_3581,N_48024,N_49116);
xnor UO_3582 (O_3582,N_47557,N_48253);
and UO_3583 (O_3583,N_49835,N_47643);
xor UO_3584 (O_3584,N_48542,N_48359);
or UO_3585 (O_3585,N_48227,N_47545);
nand UO_3586 (O_3586,N_47736,N_49840);
xor UO_3587 (O_3587,N_49285,N_49465);
xnor UO_3588 (O_3588,N_49553,N_47741);
xor UO_3589 (O_3589,N_48101,N_49715);
nor UO_3590 (O_3590,N_49890,N_47968);
nor UO_3591 (O_3591,N_48799,N_48184);
and UO_3592 (O_3592,N_48081,N_48149);
or UO_3593 (O_3593,N_49364,N_48223);
or UO_3594 (O_3594,N_48005,N_48761);
nand UO_3595 (O_3595,N_47765,N_48966);
and UO_3596 (O_3596,N_49321,N_48530);
and UO_3597 (O_3597,N_48684,N_49508);
nand UO_3598 (O_3598,N_49785,N_49048);
or UO_3599 (O_3599,N_49797,N_49912);
nand UO_3600 (O_3600,N_49435,N_47529);
and UO_3601 (O_3601,N_48208,N_49477);
or UO_3602 (O_3602,N_48915,N_49590);
or UO_3603 (O_3603,N_48976,N_49549);
xor UO_3604 (O_3604,N_47764,N_47747);
and UO_3605 (O_3605,N_47779,N_49976);
nand UO_3606 (O_3606,N_49812,N_49690);
xor UO_3607 (O_3607,N_48127,N_49088);
or UO_3608 (O_3608,N_49374,N_48290);
nand UO_3609 (O_3609,N_48635,N_48661);
nand UO_3610 (O_3610,N_47589,N_48663);
nor UO_3611 (O_3611,N_48752,N_48787);
nand UO_3612 (O_3612,N_48853,N_49129);
nand UO_3613 (O_3613,N_48624,N_48748);
nand UO_3614 (O_3614,N_49123,N_47869);
and UO_3615 (O_3615,N_49478,N_47830);
xnor UO_3616 (O_3616,N_47568,N_47926);
nor UO_3617 (O_3617,N_49174,N_48705);
or UO_3618 (O_3618,N_49993,N_49085);
or UO_3619 (O_3619,N_47817,N_49050);
and UO_3620 (O_3620,N_48393,N_49438);
xor UO_3621 (O_3621,N_48351,N_48384);
xor UO_3622 (O_3622,N_49759,N_49536);
or UO_3623 (O_3623,N_48180,N_47500);
nand UO_3624 (O_3624,N_48964,N_49925);
xor UO_3625 (O_3625,N_48689,N_48400);
nand UO_3626 (O_3626,N_47938,N_47987);
nand UO_3627 (O_3627,N_49043,N_48337);
nor UO_3628 (O_3628,N_48762,N_49572);
xnor UO_3629 (O_3629,N_47751,N_49258);
nand UO_3630 (O_3630,N_47700,N_48052);
nor UO_3631 (O_3631,N_48236,N_47663);
nor UO_3632 (O_3632,N_49379,N_48127);
or UO_3633 (O_3633,N_47893,N_48468);
and UO_3634 (O_3634,N_48227,N_49610);
and UO_3635 (O_3635,N_48067,N_48289);
nand UO_3636 (O_3636,N_49458,N_48065);
xnor UO_3637 (O_3637,N_49136,N_48976);
nand UO_3638 (O_3638,N_47612,N_47732);
xnor UO_3639 (O_3639,N_49229,N_49026);
and UO_3640 (O_3640,N_47591,N_47798);
or UO_3641 (O_3641,N_49769,N_47798);
or UO_3642 (O_3642,N_49407,N_48033);
and UO_3643 (O_3643,N_48846,N_47519);
and UO_3644 (O_3644,N_48377,N_49326);
nand UO_3645 (O_3645,N_47723,N_49148);
or UO_3646 (O_3646,N_49167,N_47935);
and UO_3647 (O_3647,N_48329,N_49425);
and UO_3648 (O_3648,N_48660,N_48650);
nand UO_3649 (O_3649,N_49473,N_48494);
xnor UO_3650 (O_3650,N_48330,N_48434);
and UO_3651 (O_3651,N_48612,N_48762);
nor UO_3652 (O_3652,N_49808,N_49042);
xnor UO_3653 (O_3653,N_47847,N_49999);
and UO_3654 (O_3654,N_49246,N_48324);
nand UO_3655 (O_3655,N_49360,N_48653);
nor UO_3656 (O_3656,N_48691,N_48525);
nor UO_3657 (O_3657,N_48700,N_49069);
nand UO_3658 (O_3658,N_47565,N_49391);
and UO_3659 (O_3659,N_47900,N_48752);
or UO_3660 (O_3660,N_48726,N_48920);
or UO_3661 (O_3661,N_48217,N_47943);
xnor UO_3662 (O_3662,N_48194,N_48594);
or UO_3663 (O_3663,N_47984,N_49075);
or UO_3664 (O_3664,N_48704,N_49051);
nand UO_3665 (O_3665,N_48185,N_48350);
nand UO_3666 (O_3666,N_48328,N_48725);
and UO_3667 (O_3667,N_48060,N_48215);
and UO_3668 (O_3668,N_48215,N_49064);
xnor UO_3669 (O_3669,N_49902,N_47835);
or UO_3670 (O_3670,N_48821,N_49774);
or UO_3671 (O_3671,N_49282,N_47966);
xnor UO_3672 (O_3672,N_47629,N_48691);
xnor UO_3673 (O_3673,N_49569,N_47797);
xor UO_3674 (O_3674,N_49018,N_49173);
nand UO_3675 (O_3675,N_49928,N_48744);
and UO_3676 (O_3676,N_48960,N_48794);
nand UO_3677 (O_3677,N_47771,N_47661);
and UO_3678 (O_3678,N_49505,N_48773);
and UO_3679 (O_3679,N_47917,N_49788);
or UO_3680 (O_3680,N_48624,N_48824);
nand UO_3681 (O_3681,N_48162,N_49175);
xnor UO_3682 (O_3682,N_48386,N_48475);
and UO_3683 (O_3683,N_47900,N_47734);
and UO_3684 (O_3684,N_48611,N_49371);
or UO_3685 (O_3685,N_48561,N_48895);
or UO_3686 (O_3686,N_47817,N_47583);
nand UO_3687 (O_3687,N_48261,N_48713);
and UO_3688 (O_3688,N_47827,N_48185);
xnor UO_3689 (O_3689,N_48246,N_49733);
and UO_3690 (O_3690,N_49551,N_49861);
xnor UO_3691 (O_3691,N_49551,N_48771);
and UO_3692 (O_3692,N_49298,N_49952);
xnor UO_3693 (O_3693,N_48116,N_48616);
and UO_3694 (O_3694,N_49844,N_47641);
nand UO_3695 (O_3695,N_48861,N_49311);
and UO_3696 (O_3696,N_48001,N_49365);
or UO_3697 (O_3697,N_49493,N_47592);
xnor UO_3698 (O_3698,N_49678,N_49950);
and UO_3699 (O_3699,N_47569,N_47722);
and UO_3700 (O_3700,N_48193,N_47605);
or UO_3701 (O_3701,N_47969,N_48447);
or UO_3702 (O_3702,N_48325,N_49069);
and UO_3703 (O_3703,N_49475,N_49127);
and UO_3704 (O_3704,N_47868,N_48778);
nor UO_3705 (O_3705,N_48811,N_48866);
or UO_3706 (O_3706,N_48533,N_47826);
nand UO_3707 (O_3707,N_48039,N_49148);
or UO_3708 (O_3708,N_49753,N_48774);
or UO_3709 (O_3709,N_48137,N_49275);
nor UO_3710 (O_3710,N_49913,N_48847);
or UO_3711 (O_3711,N_47843,N_47542);
and UO_3712 (O_3712,N_48055,N_47594);
and UO_3713 (O_3713,N_47699,N_47792);
nand UO_3714 (O_3714,N_49777,N_48862);
or UO_3715 (O_3715,N_48162,N_48047);
nand UO_3716 (O_3716,N_48384,N_49220);
nand UO_3717 (O_3717,N_49104,N_49303);
and UO_3718 (O_3718,N_49524,N_49908);
xor UO_3719 (O_3719,N_49087,N_48793);
and UO_3720 (O_3720,N_48627,N_47621);
and UO_3721 (O_3721,N_49679,N_49473);
or UO_3722 (O_3722,N_47691,N_49015);
nor UO_3723 (O_3723,N_49277,N_49518);
nand UO_3724 (O_3724,N_49486,N_47905);
nor UO_3725 (O_3725,N_48120,N_49692);
xnor UO_3726 (O_3726,N_48222,N_49017);
nor UO_3727 (O_3727,N_49738,N_49477);
or UO_3728 (O_3728,N_48478,N_47875);
or UO_3729 (O_3729,N_48828,N_48638);
nand UO_3730 (O_3730,N_48748,N_47535);
nor UO_3731 (O_3731,N_49702,N_47844);
or UO_3732 (O_3732,N_47587,N_48362);
or UO_3733 (O_3733,N_49503,N_47948);
nor UO_3734 (O_3734,N_47943,N_48895);
xor UO_3735 (O_3735,N_48313,N_47562);
and UO_3736 (O_3736,N_49669,N_47645);
nand UO_3737 (O_3737,N_49947,N_49763);
nand UO_3738 (O_3738,N_49587,N_48543);
and UO_3739 (O_3739,N_47544,N_48494);
xnor UO_3740 (O_3740,N_47644,N_48806);
and UO_3741 (O_3741,N_48028,N_47611);
xor UO_3742 (O_3742,N_49522,N_48260);
nand UO_3743 (O_3743,N_47502,N_49360);
and UO_3744 (O_3744,N_48456,N_49545);
and UO_3745 (O_3745,N_48511,N_47888);
or UO_3746 (O_3746,N_48530,N_48016);
nand UO_3747 (O_3747,N_49728,N_49805);
or UO_3748 (O_3748,N_48449,N_49579);
xnor UO_3749 (O_3749,N_48776,N_49871);
and UO_3750 (O_3750,N_49175,N_49869);
nor UO_3751 (O_3751,N_49244,N_47761);
xor UO_3752 (O_3752,N_48107,N_49312);
and UO_3753 (O_3753,N_47965,N_47973);
xor UO_3754 (O_3754,N_49764,N_48467);
nand UO_3755 (O_3755,N_48567,N_47731);
nand UO_3756 (O_3756,N_48038,N_48934);
and UO_3757 (O_3757,N_49750,N_47580);
and UO_3758 (O_3758,N_47558,N_47661);
nor UO_3759 (O_3759,N_49298,N_48702);
xor UO_3760 (O_3760,N_49073,N_47840);
or UO_3761 (O_3761,N_48790,N_49600);
nand UO_3762 (O_3762,N_49885,N_47896);
nand UO_3763 (O_3763,N_49011,N_49922);
and UO_3764 (O_3764,N_49279,N_48662);
and UO_3765 (O_3765,N_47859,N_49533);
or UO_3766 (O_3766,N_49783,N_48569);
nand UO_3767 (O_3767,N_48287,N_48153);
xor UO_3768 (O_3768,N_48185,N_49687);
and UO_3769 (O_3769,N_48357,N_49104);
xor UO_3770 (O_3770,N_49031,N_48692);
and UO_3771 (O_3771,N_49280,N_48592);
xor UO_3772 (O_3772,N_49483,N_48323);
and UO_3773 (O_3773,N_48385,N_47909);
and UO_3774 (O_3774,N_48088,N_48178);
xnor UO_3775 (O_3775,N_49321,N_49052);
xnor UO_3776 (O_3776,N_47970,N_48162);
or UO_3777 (O_3777,N_48024,N_49964);
xnor UO_3778 (O_3778,N_47786,N_49741);
or UO_3779 (O_3779,N_48734,N_49003);
or UO_3780 (O_3780,N_49123,N_49927);
and UO_3781 (O_3781,N_48031,N_48674);
or UO_3782 (O_3782,N_49087,N_48098);
xor UO_3783 (O_3783,N_48621,N_49521);
or UO_3784 (O_3784,N_49964,N_49594);
nand UO_3785 (O_3785,N_49488,N_48499);
xor UO_3786 (O_3786,N_47980,N_48268);
xor UO_3787 (O_3787,N_49936,N_49600);
or UO_3788 (O_3788,N_48108,N_48435);
nor UO_3789 (O_3789,N_49420,N_48306);
xnor UO_3790 (O_3790,N_48156,N_49128);
xor UO_3791 (O_3791,N_48367,N_48431);
nor UO_3792 (O_3792,N_48883,N_48880);
or UO_3793 (O_3793,N_49390,N_49834);
or UO_3794 (O_3794,N_47709,N_49412);
or UO_3795 (O_3795,N_48165,N_47549);
and UO_3796 (O_3796,N_49998,N_49935);
or UO_3797 (O_3797,N_47832,N_48941);
nand UO_3798 (O_3798,N_47529,N_49669);
and UO_3799 (O_3799,N_49198,N_48634);
or UO_3800 (O_3800,N_49947,N_49253);
nand UO_3801 (O_3801,N_49077,N_48480);
or UO_3802 (O_3802,N_47659,N_49389);
and UO_3803 (O_3803,N_49571,N_47904);
or UO_3804 (O_3804,N_48974,N_49100);
or UO_3805 (O_3805,N_49533,N_48393);
xnor UO_3806 (O_3806,N_47633,N_49406);
xor UO_3807 (O_3807,N_48901,N_48453);
or UO_3808 (O_3808,N_49116,N_49921);
nand UO_3809 (O_3809,N_49583,N_49477);
nor UO_3810 (O_3810,N_49415,N_47882);
xor UO_3811 (O_3811,N_48433,N_49993);
nor UO_3812 (O_3812,N_48228,N_48929);
xnor UO_3813 (O_3813,N_48231,N_49693);
and UO_3814 (O_3814,N_48093,N_48289);
nor UO_3815 (O_3815,N_49541,N_47567);
or UO_3816 (O_3816,N_48059,N_49180);
xor UO_3817 (O_3817,N_49187,N_48035);
nor UO_3818 (O_3818,N_47791,N_48494);
nor UO_3819 (O_3819,N_49072,N_49610);
nand UO_3820 (O_3820,N_48753,N_48227);
nand UO_3821 (O_3821,N_49867,N_48685);
xor UO_3822 (O_3822,N_49464,N_47572);
nor UO_3823 (O_3823,N_47935,N_49458);
xor UO_3824 (O_3824,N_49177,N_48906);
nor UO_3825 (O_3825,N_48543,N_49661);
or UO_3826 (O_3826,N_49434,N_48735);
and UO_3827 (O_3827,N_48515,N_48908);
or UO_3828 (O_3828,N_48012,N_49913);
xor UO_3829 (O_3829,N_47835,N_49360);
nor UO_3830 (O_3830,N_49732,N_49399);
xor UO_3831 (O_3831,N_49924,N_47917);
nor UO_3832 (O_3832,N_48537,N_48800);
or UO_3833 (O_3833,N_47927,N_48476);
nor UO_3834 (O_3834,N_49744,N_49931);
and UO_3835 (O_3835,N_49563,N_49500);
xnor UO_3836 (O_3836,N_47789,N_49460);
nand UO_3837 (O_3837,N_47553,N_48001);
xor UO_3838 (O_3838,N_47534,N_49023);
xor UO_3839 (O_3839,N_48941,N_47791);
or UO_3840 (O_3840,N_49559,N_49346);
or UO_3841 (O_3841,N_48032,N_48422);
nand UO_3842 (O_3842,N_47656,N_49639);
nor UO_3843 (O_3843,N_48234,N_48525);
and UO_3844 (O_3844,N_49418,N_49239);
nor UO_3845 (O_3845,N_48482,N_48283);
and UO_3846 (O_3846,N_47899,N_49966);
nand UO_3847 (O_3847,N_47853,N_48726);
and UO_3848 (O_3848,N_49912,N_49413);
nand UO_3849 (O_3849,N_49660,N_47820);
nand UO_3850 (O_3850,N_49046,N_49690);
and UO_3851 (O_3851,N_48200,N_49759);
or UO_3852 (O_3852,N_48109,N_49689);
nand UO_3853 (O_3853,N_48681,N_49310);
or UO_3854 (O_3854,N_49930,N_48864);
nand UO_3855 (O_3855,N_49156,N_49800);
or UO_3856 (O_3856,N_48975,N_48808);
xor UO_3857 (O_3857,N_47701,N_49862);
nand UO_3858 (O_3858,N_48101,N_49172);
nor UO_3859 (O_3859,N_49915,N_48421);
xnor UO_3860 (O_3860,N_49318,N_47856);
or UO_3861 (O_3861,N_48245,N_48815);
xor UO_3862 (O_3862,N_47982,N_49024);
nand UO_3863 (O_3863,N_49313,N_49168);
xor UO_3864 (O_3864,N_48440,N_49303);
nand UO_3865 (O_3865,N_49676,N_48148);
and UO_3866 (O_3866,N_47975,N_48475);
nor UO_3867 (O_3867,N_49988,N_48603);
nand UO_3868 (O_3868,N_48765,N_48717);
or UO_3869 (O_3869,N_48405,N_49198);
nand UO_3870 (O_3870,N_49185,N_48709);
and UO_3871 (O_3871,N_49451,N_49432);
and UO_3872 (O_3872,N_48018,N_47568);
nor UO_3873 (O_3873,N_47578,N_47764);
or UO_3874 (O_3874,N_48090,N_49683);
nor UO_3875 (O_3875,N_47731,N_47894);
nand UO_3876 (O_3876,N_48774,N_49051);
or UO_3877 (O_3877,N_49720,N_48481);
or UO_3878 (O_3878,N_49087,N_47589);
nor UO_3879 (O_3879,N_48543,N_49936);
or UO_3880 (O_3880,N_48148,N_47909);
and UO_3881 (O_3881,N_47536,N_49046);
nor UO_3882 (O_3882,N_49991,N_48050);
nor UO_3883 (O_3883,N_48506,N_49292);
nor UO_3884 (O_3884,N_49884,N_48077);
xnor UO_3885 (O_3885,N_49390,N_49018);
and UO_3886 (O_3886,N_47793,N_49892);
nand UO_3887 (O_3887,N_47916,N_47903);
nand UO_3888 (O_3888,N_48724,N_47707);
xnor UO_3889 (O_3889,N_47906,N_49319);
nand UO_3890 (O_3890,N_49695,N_48422);
or UO_3891 (O_3891,N_48219,N_49961);
xnor UO_3892 (O_3892,N_48560,N_48970);
and UO_3893 (O_3893,N_49054,N_48772);
xor UO_3894 (O_3894,N_47589,N_48379);
nand UO_3895 (O_3895,N_48379,N_48030);
xnor UO_3896 (O_3896,N_49422,N_49859);
and UO_3897 (O_3897,N_48854,N_47646);
nand UO_3898 (O_3898,N_47589,N_49500);
nor UO_3899 (O_3899,N_49077,N_49015);
or UO_3900 (O_3900,N_48106,N_49299);
nand UO_3901 (O_3901,N_47846,N_48944);
nor UO_3902 (O_3902,N_49770,N_48967);
or UO_3903 (O_3903,N_47832,N_47811);
nand UO_3904 (O_3904,N_49260,N_48286);
nand UO_3905 (O_3905,N_47859,N_47965);
and UO_3906 (O_3906,N_48887,N_47653);
or UO_3907 (O_3907,N_48214,N_49823);
and UO_3908 (O_3908,N_48605,N_48240);
xor UO_3909 (O_3909,N_47764,N_48301);
and UO_3910 (O_3910,N_49496,N_49519);
or UO_3911 (O_3911,N_47929,N_47640);
or UO_3912 (O_3912,N_47632,N_47694);
or UO_3913 (O_3913,N_49737,N_48850);
xnor UO_3914 (O_3914,N_48911,N_49406);
and UO_3915 (O_3915,N_49143,N_49140);
or UO_3916 (O_3916,N_49783,N_49194);
xnor UO_3917 (O_3917,N_49147,N_49519);
xnor UO_3918 (O_3918,N_48230,N_48270);
nand UO_3919 (O_3919,N_49592,N_47673);
and UO_3920 (O_3920,N_48251,N_48126);
xor UO_3921 (O_3921,N_48991,N_49027);
and UO_3922 (O_3922,N_49823,N_49537);
and UO_3923 (O_3923,N_48325,N_49717);
or UO_3924 (O_3924,N_49162,N_48908);
xnor UO_3925 (O_3925,N_49088,N_49630);
xor UO_3926 (O_3926,N_48260,N_48810);
or UO_3927 (O_3927,N_48833,N_47982);
xor UO_3928 (O_3928,N_49873,N_49338);
and UO_3929 (O_3929,N_47581,N_49228);
or UO_3930 (O_3930,N_48878,N_48428);
or UO_3931 (O_3931,N_47574,N_48694);
nor UO_3932 (O_3932,N_49718,N_49252);
nor UO_3933 (O_3933,N_48272,N_48554);
nand UO_3934 (O_3934,N_48636,N_48196);
nor UO_3935 (O_3935,N_47704,N_48726);
and UO_3936 (O_3936,N_49778,N_47603);
nor UO_3937 (O_3937,N_48753,N_49781);
and UO_3938 (O_3938,N_49745,N_48945);
nor UO_3939 (O_3939,N_48451,N_49320);
or UO_3940 (O_3940,N_47579,N_49650);
or UO_3941 (O_3941,N_49189,N_48612);
xor UO_3942 (O_3942,N_49665,N_49342);
and UO_3943 (O_3943,N_48350,N_48982);
nor UO_3944 (O_3944,N_48273,N_48714);
nand UO_3945 (O_3945,N_48900,N_48399);
nand UO_3946 (O_3946,N_48190,N_49920);
xnor UO_3947 (O_3947,N_49324,N_49538);
nor UO_3948 (O_3948,N_49420,N_47615);
or UO_3949 (O_3949,N_49630,N_49727);
nand UO_3950 (O_3950,N_48128,N_47733);
nor UO_3951 (O_3951,N_48444,N_49392);
nor UO_3952 (O_3952,N_48407,N_48325);
nor UO_3953 (O_3953,N_48380,N_49385);
nand UO_3954 (O_3954,N_48497,N_48453);
nand UO_3955 (O_3955,N_47890,N_47966);
xor UO_3956 (O_3956,N_47519,N_47940);
or UO_3957 (O_3957,N_47708,N_49806);
or UO_3958 (O_3958,N_49834,N_49210);
xnor UO_3959 (O_3959,N_49995,N_49954);
or UO_3960 (O_3960,N_49220,N_48170);
nor UO_3961 (O_3961,N_49594,N_48264);
nor UO_3962 (O_3962,N_48836,N_48831);
nor UO_3963 (O_3963,N_49693,N_49181);
and UO_3964 (O_3964,N_48653,N_49607);
xor UO_3965 (O_3965,N_48007,N_47952);
xnor UO_3966 (O_3966,N_48691,N_49421);
or UO_3967 (O_3967,N_48237,N_47971);
nand UO_3968 (O_3968,N_47676,N_49597);
xnor UO_3969 (O_3969,N_48656,N_48582);
or UO_3970 (O_3970,N_49297,N_49415);
and UO_3971 (O_3971,N_49219,N_48050);
xnor UO_3972 (O_3972,N_48873,N_48355);
xnor UO_3973 (O_3973,N_48808,N_49593);
nand UO_3974 (O_3974,N_48407,N_47517);
xor UO_3975 (O_3975,N_48183,N_49982);
xor UO_3976 (O_3976,N_49279,N_47534);
or UO_3977 (O_3977,N_47755,N_47948);
nand UO_3978 (O_3978,N_49627,N_49725);
nor UO_3979 (O_3979,N_48054,N_49260);
or UO_3980 (O_3980,N_49116,N_48237);
or UO_3981 (O_3981,N_48076,N_48416);
or UO_3982 (O_3982,N_49412,N_48692);
xnor UO_3983 (O_3983,N_48786,N_48502);
nand UO_3984 (O_3984,N_49726,N_48297);
or UO_3985 (O_3985,N_49177,N_48099);
xor UO_3986 (O_3986,N_47620,N_48631);
and UO_3987 (O_3987,N_49038,N_49199);
and UO_3988 (O_3988,N_48887,N_48864);
or UO_3989 (O_3989,N_49556,N_49754);
xor UO_3990 (O_3990,N_49649,N_48310);
or UO_3991 (O_3991,N_48590,N_49895);
nand UO_3992 (O_3992,N_49213,N_49287);
and UO_3993 (O_3993,N_49549,N_49568);
nor UO_3994 (O_3994,N_47640,N_49989);
or UO_3995 (O_3995,N_47576,N_48416);
and UO_3996 (O_3996,N_47739,N_49244);
nand UO_3997 (O_3997,N_49576,N_49355);
xnor UO_3998 (O_3998,N_48313,N_48758);
or UO_3999 (O_3999,N_48643,N_48337);
nor UO_4000 (O_4000,N_48883,N_48581);
xnor UO_4001 (O_4001,N_47518,N_49715);
or UO_4002 (O_4002,N_49970,N_47866);
xor UO_4003 (O_4003,N_49675,N_49157);
xnor UO_4004 (O_4004,N_48972,N_48697);
or UO_4005 (O_4005,N_49796,N_47778);
xnor UO_4006 (O_4006,N_49136,N_47549);
nand UO_4007 (O_4007,N_48000,N_49711);
xnor UO_4008 (O_4008,N_48438,N_49438);
and UO_4009 (O_4009,N_48342,N_47534);
nand UO_4010 (O_4010,N_48682,N_48539);
xor UO_4011 (O_4011,N_49865,N_48752);
nand UO_4012 (O_4012,N_48122,N_49982);
nor UO_4013 (O_4013,N_47638,N_49528);
and UO_4014 (O_4014,N_49682,N_47649);
nor UO_4015 (O_4015,N_48937,N_49112);
nand UO_4016 (O_4016,N_48323,N_48386);
xor UO_4017 (O_4017,N_47542,N_49452);
and UO_4018 (O_4018,N_49371,N_49226);
or UO_4019 (O_4019,N_48066,N_47898);
nor UO_4020 (O_4020,N_49680,N_49017);
nor UO_4021 (O_4021,N_48634,N_48259);
xnor UO_4022 (O_4022,N_48557,N_48593);
xor UO_4023 (O_4023,N_49096,N_48960);
and UO_4024 (O_4024,N_48815,N_48785);
xnor UO_4025 (O_4025,N_48889,N_49259);
nor UO_4026 (O_4026,N_48459,N_49631);
and UO_4027 (O_4027,N_47612,N_49952);
and UO_4028 (O_4028,N_47836,N_49081);
nor UO_4029 (O_4029,N_47888,N_48025);
and UO_4030 (O_4030,N_49961,N_47719);
nor UO_4031 (O_4031,N_49863,N_47649);
nand UO_4032 (O_4032,N_49783,N_49631);
xnor UO_4033 (O_4033,N_48121,N_48186);
nor UO_4034 (O_4034,N_47778,N_47914);
xor UO_4035 (O_4035,N_48102,N_49836);
nor UO_4036 (O_4036,N_48406,N_49584);
or UO_4037 (O_4037,N_49359,N_49935);
or UO_4038 (O_4038,N_48757,N_49669);
or UO_4039 (O_4039,N_48001,N_48278);
and UO_4040 (O_4040,N_47907,N_49148);
nand UO_4041 (O_4041,N_47541,N_49637);
nor UO_4042 (O_4042,N_49184,N_49739);
xor UO_4043 (O_4043,N_48521,N_49888);
xor UO_4044 (O_4044,N_48808,N_47898);
xnor UO_4045 (O_4045,N_48767,N_48465);
and UO_4046 (O_4046,N_47553,N_48994);
xnor UO_4047 (O_4047,N_48444,N_49842);
xor UO_4048 (O_4048,N_49109,N_49946);
nor UO_4049 (O_4049,N_49908,N_49721);
nor UO_4050 (O_4050,N_48766,N_48208);
and UO_4051 (O_4051,N_48626,N_48465);
and UO_4052 (O_4052,N_49659,N_49998);
xor UO_4053 (O_4053,N_49510,N_48875);
nor UO_4054 (O_4054,N_48764,N_48022);
nor UO_4055 (O_4055,N_47652,N_48155);
and UO_4056 (O_4056,N_49604,N_48006);
and UO_4057 (O_4057,N_49013,N_49273);
xnor UO_4058 (O_4058,N_49643,N_49571);
xnor UO_4059 (O_4059,N_48821,N_47920);
xnor UO_4060 (O_4060,N_49675,N_47623);
nand UO_4061 (O_4061,N_48205,N_48065);
nor UO_4062 (O_4062,N_49843,N_48383);
nor UO_4063 (O_4063,N_47891,N_49684);
or UO_4064 (O_4064,N_48722,N_47829);
nand UO_4065 (O_4065,N_48671,N_48806);
nor UO_4066 (O_4066,N_48072,N_47862);
or UO_4067 (O_4067,N_48535,N_47853);
and UO_4068 (O_4068,N_48260,N_49792);
xnor UO_4069 (O_4069,N_49023,N_48404);
and UO_4070 (O_4070,N_48353,N_49338);
nor UO_4071 (O_4071,N_49629,N_49965);
xnor UO_4072 (O_4072,N_47593,N_48189);
nand UO_4073 (O_4073,N_48844,N_48420);
nor UO_4074 (O_4074,N_49225,N_48983);
or UO_4075 (O_4075,N_48391,N_48376);
nor UO_4076 (O_4076,N_48150,N_47524);
xor UO_4077 (O_4077,N_49821,N_47670);
and UO_4078 (O_4078,N_49143,N_47517);
nand UO_4079 (O_4079,N_47913,N_49459);
nand UO_4080 (O_4080,N_49543,N_47590);
nor UO_4081 (O_4081,N_48434,N_49149);
xnor UO_4082 (O_4082,N_48284,N_49344);
or UO_4083 (O_4083,N_48494,N_48059);
xor UO_4084 (O_4084,N_48727,N_47799);
nor UO_4085 (O_4085,N_49076,N_49162);
or UO_4086 (O_4086,N_48469,N_49242);
or UO_4087 (O_4087,N_48449,N_49712);
xnor UO_4088 (O_4088,N_49351,N_47507);
xor UO_4089 (O_4089,N_47686,N_48062);
nor UO_4090 (O_4090,N_49847,N_49361);
xnor UO_4091 (O_4091,N_48447,N_47747);
nor UO_4092 (O_4092,N_49745,N_47956);
or UO_4093 (O_4093,N_47543,N_47723);
or UO_4094 (O_4094,N_49582,N_49366);
nor UO_4095 (O_4095,N_49126,N_49568);
xor UO_4096 (O_4096,N_49642,N_47544);
nand UO_4097 (O_4097,N_47867,N_49456);
xnor UO_4098 (O_4098,N_49039,N_48877);
or UO_4099 (O_4099,N_48702,N_48081);
nand UO_4100 (O_4100,N_49159,N_49619);
xnor UO_4101 (O_4101,N_47845,N_48395);
nor UO_4102 (O_4102,N_47665,N_47673);
nor UO_4103 (O_4103,N_49118,N_49812);
or UO_4104 (O_4104,N_47585,N_47523);
and UO_4105 (O_4105,N_48301,N_48705);
nor UO_4106 (O_4106,N_48541,N_48191);
and UO_4107 (O_4107,N_48809,N_47924);
or UO_4108 (O_4108,N_47539,N_48463);
or UO_4109 (O_4109,N_49073,N_49030);
or UO_4110 (O_4110,N_49378,N_48826);
and UO_4111 (O_4111,N_49281,N_47619);
nor UO_4112 (O_4112,N_47549,N_48172);
nor UO_4113 (O_4113,N_49851,N_48311);
nand UO_4114 (O_4114,N_47967,N_49207);
nand UO_4115 (O_4115,N_49408,N_48863);
and UO_4116 (O_4116,N_48365,N_48519);
or UO_4117 (O_4117,N_48256,N_49732);
nand UO_4118 (O_4118,N_49309,N_48484);
and UO_4119 (O_4119,N_48625,N_48343);
and UO_4120 (O_4120,N_48228,N_49779);
xnor UO_4121 (O_4121,N_48733,N_49481);
xnor UO_4122 (O_4122,N_48529,N_47822);
nand UO_4123 (O_4123,N_49782,N_49121);
xnor UO_4124 (O_4124,N_48679,N_49018);
and UO_4125 (O_4125,N_48244,N_47707);
or UO_4126 (O_4126,N_48531,N_49126);
nand UO_4127 (O_4127,N_48171,N_49939);
and UO_4128 (O_4128,N_49235,N_49205);
xor UO_4129 (O_4129,N_49350,N_48053);
nor UO_4130 (O_4130,N_49513,N_47534);
nand UO_4131 (O_4131,N_47810,N_47546);
xor UO_4132 (O_4132,N_49309,N_49438);
nor UO_4133 (O_4133,N_48727,N_49178);
or UO_4134 (O_4134,N_49658,N_48644);
nor UO_4135 (O_4135,N_48330,N_49247);
xor UO_4136 (O_4136,N_49012,N_49679);
nand UO_4137 (O_4137,N_48975,N_49717);
nor UO_4138 (O_4138,N_49330,N_48600);
or UO_4139 (O_4139,N_49666,N_47906);
nor UO_4140 (O_4140,N_49080,N_48905);
or UO_4141 (O_4141,N_48131,N_48641);
and UO_4142 (O_4142,N_48940,N_49028);
and UO_4143 (O_4143,N_48702,N_47759);
nor UO_4144 (O_4144,N_48872,N_47916);
xnor UO_4145 (O_4145,N_48261,N_47622);
and UO_4146 (O_4146,N_49417,N_48751);
or UO_4147 (O_4147,N_47846,N_48533);
nor UO_4148 (O_4148,N_49723,N_47552);
and UO_4149 (O_4149,N_48256,N_49608);
nor UO_4150 (O_4150,N_49441,N_48044);
xor UO_4151 (O_4151,N_49416,N_48821);
nor UO_4152 (O_4152,N_48050,N_47704);
and UO_4153 (O_4153,N_49189,N_48565);
and UO_4154 (O_4154,N_48484,N_49166);
or UO_4155 (O_4155,N_48336,N_49064);
or UO_4156 (O_4156,N_48835,N_49774);
and UO_4157 (O_4157,N_47814,N_49211);
nand UO_4158 (O_4158,N_49562,N_48780);
and UO_4159 (O_4159,N_49298,N_47678);
nor UO_4160 (O_4160,N_47900,N_49055);
nand UO_4161 (O_4161,N_49298,N_48178);
xnor UO_4162 (O_4162,N_48568,N_49674);
nor UO_4163 (O_4163,N_49994,N_49648);
or UO_4164 (O_4164,N_49263,N_49699);
xnor UO_4165 (O_4165,N_48514,N_49776);
nand UO_4166 (O_4166,N_48558,N_48444);
xnor UO_4167 (O_4167,N_48872,N_47721);
nor UO_4168 (O_4168,N_48209,N_49283);
xor UO_4169 (O_4169,N_47571,N_47547);
nor UO_4170 (O_4170,N_47524,N_49232);
nor UO_4171 (O_4171,N_48366,N_48433);
or UO_4172 (O_4172,N_49700,N_48996);
nand UO_4173 (O_4173,N_48125,N_48228);
and UO_4174 (O_4174,N_49559,N_47595);
or UO_4175 (O_4175,N_49395,N_48725);
and UO_4176 (O_4176,N_49911,N_48589);
nor UO_4177 (O_4177,N_49241,N_49427);
xnor UO_4178 (O_4178,N_49699,N_48753);
and UO_4179 (O_4179,N_49835,N_48382);
xnor UO_4180 (O_4180,N_49324,N_48986);
and UO_4181 (O_4181,N_49398,N_49489);
or UO_4182 (O_4182,N_49913,N_49433);
nand UO_4183 (O_4183,N_47976,N_49801);
and UO_4184 (O_4184,N_49985,N_47934);
or UO_4185 (O_4185,N_47776,N_47930);
xnor UO_4186 (O_4186,N_48182,N_49177);
or UO_4187 (O_4187,N_49831,N_49583);
or UO_4188 (O_4188,N_48490,N_48663);
nor UO_4189 (O_4189,N_47822,N_47794);
nand UO_4190 (O_4190,N_49764,N_48976);
nand UO_4191 (O_4191,N_49588,N_49363);
nand UO_4192 (O_4192,N_48384,N_49037);
or UO_4193 (O_4193,N_48919,N_48193);
xnor UO_4194 (O_4194,N_47754,N_48866);
xnor UO_4195 (O_4195,N_47834,N_48203);
or UO_4196 (O_4196,N_48035,N_48876);
and UO_4197 (O_4197,N_49930,N_48163);
and UO_4198 (O_4198,N_49082,N_47704);
or UO_4199 (O_4199,N_47685,N_48264);
xnor UO_4200 (O_4200,N_49249,N_49268);
xnor UO_4201 (O_4201,N_48205,N_48469);
nor UO_4202 (O_4202,N_48875,N_49692);
xnor UO_4203 (O_4203,N_48334,N_49599);
nor UO_4204 (O_4204,N_47510,N_48984);
nor UO_4205 (O_4205,N_49853,N_48946);
nand UO_4206 (O_4206,N_49332,N_48795);
and UO_4207 (O_4207,N_49524,N_49685);
or UO_4208 (O_4208,N_49343,N_48082);
or UO_4209 (O_4209,N_48373,N_49737);
nand UO_4210 (O_4210,N_47548,N_49362);
nand UO_4211 (O_4211,N_49201,N_48798);
or UO_4212 (O_4212,N_49808,N_49397);
nor UO_4213 (O_4213,N_49443,N_48397);
nor UO_4214 (O_4214,N_49433,N_49915);
nand UO_4215 (O_4215,N_48083,N_48710);
xnor UO_4216 (O_4216,N_48513,N_48422);
nand UO_4217 (O_4217,N_49921,N_48664);
nand UO_4218 (O_4218,N_49328,N_48933);
and UO_4219 (O_4219,N_49983,N_48697);
and UO_4220 (O_4220,N_48771,N_48483);
xor UO_4221 (O_4221,N_49769,N_49590);
and UO_4222 (O_4222,N_47761,N_47505);
and UO_4223 (O_4223,N_49140,N_48332);
and UO_4224 (O_4224,N_47620,N_47864);
xnor UO_4225 (O_4225,N_48818,N_49175);
or UO_4226 (O_4226,N_49845,N_48594);
and UO_4227 (O_4227,N_47730,N_48226);
nor UO_4228 (O_4228,N_48878,N_49618);
xor UO_4229 (O_4229,N_48313,N_49381);
xnor UO_4230 (O_4230,N_49997,N_48494);
and UO_4231 (O_4231,N_47639,N_48076);
xor UO_4232 (O_4232,N_49597,N_47956);
and UO_4233 (O_4233,N_48517,N_49570);
or UO_4234 (O_4234,N_48341,N_48676);
nand UO_4235 (O_4235,N_49745,N_49753);
xnor UO_4236 (O_4236,N_47511,N_47779);
xnor UO_4237 (O_4237,N_48284,N_48893);
xor UO_4238 (O_4238,N_48906,N_48148);
or UO_4239 (O_4239,N_47573,N_48246);
or UO_4240 (O_4240,N_49299,N_49744);
nand UO_4241 (O_4241,N_48471,N_47826);
xnor UO_4242 (O_4242,N_49439,N_49935);
nor UO_4243 (O_4243,N_49953,N_49421);
nor UO_4244 (O_4244,N_49920,N_48155);
xnor UO_4245 (O_4245,N_48815,N_48544);
or UO_4246 (O_4246,N_48080,N_47761);
nand UO_4247 (O_4247,N_49025,N_49184);
and UO_4248 (O_4248,N_49391,N_49075);
and UO_4249 (O_4249,N_48471,N_48893);
nor UO_4250 (O_4250,N_48281,N_48027);
xnor UO_4251 (O_4251,N_49907,N_48603);
or UO_4252 (O_4252,N_48641,N_48202);
and UO_4253 (O_4253,N_48280,N_48985);
xnor UO_4254 (O_4254,N_49964,N_48642);
nand UO_4255 (O_4255,N_48012,N_48026);
nand UO_4256 (O_4256,N_47809,N_48310);
xnor UO_4257 (O_4257,N_49640,N_48274);
nor UO_4258 (O_4258,N_49272,N_48177);
and UO_4259 (O_4259,N_47526,N_49826);
nor UO_4260 (O_4260,N_48686,N_47501);
xnor UO_4261 (O_4261,N_48903,N_49324);
nor UO_4262 (O_4262,N_48493,N_49163);
or UO_4263 (O_4263,N_48527,N_49631);
xnor UO_4264 (O_4264,N_48053,N_48016);
nor UO_4265 (O_4265,N_47640,N_48330);
and UO_4266 (O_4266,N_49599,N_49008);
nor UO_4267 (O_4267,N_48816,N_49398);
and UO_4268 (O_4268,N_48635,N_48947);
or UO_4269 (O_4269,N_49713,N_48300);
or UO_4270 (O_4270,N_49313,N_47668);
xnor UO_4271 (O_4271,N_49009,N_48564);
nand UO_4272 (O_4272,N_48377,N_47559);
nor UO_4273 (O_4273,N_48464,N_47971);
or UO_4274 (O_4274,N_48019,N_49894);
nand UO_4275 (O_4275,N_48779,N_48813);
nor UO_4276 (O_4276,N_49751,N_48698);
nor UO_4277 (O_4277,N_49942,N_48938);
nand UO_4278 (O_4278,N_49990,N_47854);
or UO_4279 (O_4279,N_47528,N_48770);
nand UO_4280 (O_4280,N_48862,N_47592);
and UO_4281 (O_4281,N_49895,N_49926);
or UO_4282 (O_4282,N_48877,N_49252);
nand UO_4283 (O_4283,N_47930,N_48378);
nand UO_4284 (O_4284,N_47632,N_48231);
nor UO_4285 (O_4285,N_49941,N_48104);
nand UO_4286 (O_4286,N_48734,N_48875);
and UO_4287 (O_4287,N_49601,N_48365);
or UO_4288 (O_4288,N_48689,N_48521);
or UO_4289 (O_4289,N_47728,N_49344);
xor UO_4290 (O_4290,N_48966,N_48446);
nand UO_4291 (O_4291,N_47572,N_47629);
nand UO_4292 (O_4292,N_48928,N_49905);
and UO_4293 (O_4293,N_47672,N_47575);
and UO_4294 (O_4294,N_48460,N_49290);
or UO_4295 (O_4295,N_49243,N_47956);
nor UO_4296 (O_4296,N_49937,N_48906);
nor UO_4297 (O_4297,N_49481,N_49904);
nand UO_4298 (O_4298,N_48447,N_49714);
nor UO_4299 (O_4299,N_47758,N_49247);
nand UO_4300 (O_4300,N_48442,N_47705);
nand UO_4301 (O_4301,N_49509,N_47737);
nand UO_4302 (O_4302,N_48496,N_48506);
and UO_4303 (O_4303,N_49755,N_47610);
xnor UO_4304 (O_4304,N_47869,N_48591);
nand UO_4305 (O_4305,N_49047,N_47623);
and UO_4306 (O_4306,N_48797,N_48939);
or UO_4307 (O_4307,N_49040,N_48136);
xor UO_4308 (O_4308,N_48024,N_49076);
and UO_4309 (O_4309,N_49455,N_48447);
nand UO_4310 (O_4310,N_48442,N_48260);
nor UO_4311 (O_4311,N_48259,N_48745);
nand UO_4312 (O_4312,N_49740,N_48376);
or UO_4313 (O_4313,N_48004,N_48884);
nand UO_4314 (O_4314,N_48831,N_49498);
xnor UO_4315 (O_4315,N_47867,N_49262);
and UO_4316 (O_4316,N_48376,N_49758);
or UO_4317 (O_4317,N_47795,N_48030);
nor UO_4318 (O_4318,N_49064,N_47851);
and UO_4319 (O_4319,N_47721,N_48004);
or UO_4320 (O_4320,N_48546,N_47708);
or UO_4321 (O_4321,N_48526,N_48177);
xor UO_4322 (O_4322,N_49083,N_49019);
xnor UO_4323 (O_4323,N_49504,N_49004);
xnor UO_4324 (O_4324,N_49112,N_48817);
xnor UO_4325 (O_4325,N_48187,N_47940);
or UO_4326 (O_4326,N_49948,N_48083);
and UO_4327 (O_4327,N_47901,N_49108);
xnor UO_4328 (O_4328,N_49131,N_49068);
nor UO_4329 (O_4329,N_48695,N_47583);
xor UO_4330 (O_4330,N_48911,N_49720);
and UO_4331 (O_4331,N_49947,N_49972);
nand UO_4332 (O_4332,N_48658,N_49838);
xor UO_4333 (O_4333,N_49330,N_48266);
or UO_4334 (O_4334,N_47720,N_49604);
nor UO_4335 (O_4335,N_48191,N_47730);
nor UO_4336 (O_4336,N_48114,N_48532);
nand UO_4337 (O_4337,N_49356,N_49830);
xnor UO_4338 (O_4338,N_49878,N_49370);
or UO_4339 (O_4339,N_48504,N_48015);
nand UO_4340 (O_4340,N_47663,N_47640);
and UO_4341 (O_4341,N_49315,N_49480);
nor UO_4342 (O_4342,N_49915,N_49721);
nor UO_4343 (O_4343,N_48612,N_47899);
and UO_4344 (O_4344,N_48012,N_48784);
xor UO_4345 (O_4345,N_48510,N_49068);
xnor UO_4346 (O_4346,N_47962,N_47808);
nor UO_4347 (O_4347,N_47879,N_48754);
xor UO_4348 (O_4348,N_49063,N_47531);
nand UO_4349 (O_4349,N_48307,N_49877);
nand UO_4350 (O_4350,N_47760,N_47791);
nor UO_4351 (O_4351,N_49925,N_48369);
nor UO_4352 (O_4352,N_49981,N_47681);
and UO_4353 (O_4353,N_47529,N_49180);
nand UO_4354 (O_4354,N_48497,N_49784);
or UO_4355 (O_4355,N_47879,N_48084);
nand UO_4356 (O_4356,N_49070,N_48189);
xnor UO_4357 (O_4357,N_48692,N_48317);
and UO_4358 (O_4358,N_49702,N_48266);
or UO_4359 (O_4359,N_47748,N_47698);
nor UO_4360 (O_4360,N_48519,N_47508);
or UO_4361 (O_4361,N_48602,N_48364);
or UO_4362 (O_4362,N_48574,N_47548);
or UO_4363 (O_4363,N_48757,N_49695);
xnor UO_4364 (O_4364,N_49746,N_48069);
and UO_4365 (O_4365,N_48807,N_49099);
and UO_4366 (O_4366,N_48265,N_47796);
nor UO_4367 (O_4367,N_47650,N_49108);
nor UO_4368 (O_4368,N_48380,N_49793);
or UO_4369 (O_4369,N_48158,N_49782);
nor UO_4370 (O_4370,N_48609,N_49037);
nor UO_4371 (O_4371,N_49545,N_47597);
or UO_4372 (O_4372,N_47854,N_49789);
nand UO_4373 (O_4373,N_49635,N_48183);
nor UO_4374 (O_4374,N_49709,N_48820);
nor UO_4375 (O_4375,N_48097,N_48269);
nand UO_4376 (O_4376,N_47628,N_49634);
nand UO_4377 (O_4377,N_49957,N_48524);
and UO_4378 (O_4378,N_48662,N_47824);
nand UO_4379 (O_4379,N_49316,N_48649);
nand UO_4380 (O_4380,N_47800,N_48144);
xor UO_4381 (O_4381,N_48951,N_49136);
and UO_4382 (O_4382,N_47731,N_48837);
or UO_4383 (O_4383,N_47503,N_48844);
nand UO_4384 (O_4384,N_47591,N_49766);
and UO_4385 (O_4385,N_48981,N_48626);
xor UO_4386 (O_4386,N_48290,N_47786);
nor UO_4387 (O_4387,N_48491,N_49063);
nor UO_4388 (O_4388,N_48653,N_47631);
or UO_4389 (O_4389,N_49862,N_49050);
or UO_4390 (O_4390,N_47774,N_48661);
xor UO_4391 (O_4391,N_48350,N_48041);
xnor UO_4392 (O_4392,N_49818,N_48258);
and UO_4393 (O_4393,N_48763,N_48153);
xnor UO_4394 (O_4394,N_49392,N_48491);
and UO_4395 (O_4395,N_49020,N_48027);
xor UO_4396 (O_4396,N_47520,N_48491);
or UO_4397 (O_4397,N_49049,N_49802);
xnor UO_4398 (O_4398,N_47735,N_49049);
or UO_4399 (O_4399,N_48379,N_48466);
xor UO_4400 (O_4400,N_48603,N_49578);
xnor UO_4401 (O_4401,N_49384,N_48417);
xor UO_4402 (O_4402,N_49669,N_49674);
or UO_4403 (O_4403,N_47825,N_47789);
xnor UO_4404 (O_4404,N_47838,N_49200);
xnor UO_4405 (O_4405,N_47528,N_48318);
nand UO_4406 (O_4406,N_49973,N_49711);
nor UO_4407 (O_4407,N_48110,N_47807);
nor UO_4408 (O_4408,N_49430,N_48727);
nor UO_4409 (O_4409,N_48307,N_49993);
nand UO_4410 (O_4410,N_49058,N_49987);
and UO_4411 (O_4411,N_48592,N_48897);
or UO_4412 (O_4412,N_48847,N_48979);
and UO_4413 (O_4413,N_47760,N_49395);
nand UO_4414 (O_4414,N_49731,N_47661);
nand UO_4415 (O_4415,N_48865,N_48143);
xnor UO_4416 (O_4416,N_48201,N_47602);
or UO_4417 (O_4417,N_48352,N_49692);
and UO_4418 (O_4418,N_48767,N_49681);
nor UO_4419 (O_4419,N_49974,N_49774);
xnor UO_4420 (O_4420,N_48000,N_49456);
xor UO_4421 (O_4421,N_49565,N_49443);
and UO_4422 (O_4422,N_49178,N_49379);
nor UO_4423 (O_4423,N_49037,N_48890);
or UO_4424 (O_4424,N_49507,N_49157);
nand UO_4425 (O_4425,N_48912,N_49393);
xor UO_4426 (O_4426,N_49668,N_49830);
nand UO_4427 (O_4427,N_49626,N_47689);
nor UO_4428 (O_4428,N_49475,N_47563);
xor UO_4429 (O_4429,N_47993,N_47836);
nor UO_4430 (O_4430,N_49942,N_49762);
or UO_4431 (O_4431,N_48874,N_48898);
nand UO_4432 (O_4432,N_48816,N_47899);
xor UO_4433 (O_4433,N_48877,N_47968);
nor UO_4434 (O_4434,N_49997,N_48224);
nor UO_4435 (O_4435,N_49695,N_48327);
nor UO_4436 (O_4436,N_47891,N_48709);
nand UO_4437 (O_4437,N_48739,N_47838);
nand UO_4438 (O_4438,N_48599,N_49006);
and UO_4439 (O_4439,N_49761,N_48240);
nand UO_4440 (O_4440,N_49680,N_48798);
or UO_4441 (O_4441,N_47847,N_49944);
xnor UO_4442 (O_4442,N_49981,N_48639);
or UO_4443 (O_4443,N_47881,N_49116);
nand UO_4444 (O_4444,N_49147,N_49504);
xor UO_4445 (O_4445,N_48924,N_47560);
and UO_4446 (O_4446,N_47784,N_48582);
and UO_4447 (O_4447,N_49660,N_47817);
xnor UO_4448 (O_4448,N_47806,N_47978);
and UO_4449 (O_4449,N_48239,N_48840);
nand UO_4450 (O_4450,N_48525,N_47508);
nor UO_4451 (O_4451,N_49493,N_49627);
and UO_4452 (O_4452,N_49987,N_49243);
nor UO_4453 (O_4453,N_48881,N_48021);
nand UO_4454 (O_4454,N_49598,N_48532);
nor UO_4455 (O_4455,N_48998,N_48401);
nand UO_4456 (O_4456,N_48422,N_49645);
or UO_4457 (O_4457,N_49250,N_47936);
xnor UO_4458 (O_4458,N_47556,N_48732);
and UO_4459 (O_4459,N_49308,N_49948);
and UO_4460 (O_4460,N_48309,N_48809);
or UO_4461 (O_4461,N_49013,N_49794);
nor UO_4462 (O_4462,N_47662,N_49124);
and UO_4463 (O_4463,N_47547,N_49049);
or UO_4464 (O_4464,N_49306,N_49159);
or UO_4465 (O_4465,N_48825,N_49271);
nor UO_4466 (O_4466,N_48253,N_48814);
xnor UO_4467 (O_4467,N_47833,N_48227);
nor UO_4468 (O_4468,N_48798,N_48050);
xnor UO_4469 (O_4469,N_48509,N_49131);
and UO_4470 (O_4470,N_48587,N_49769);
xnor UO_4471 (O_4471,N_48943,N_47999);
and UO_4472 (O_4472,N_49947,N_47536);
and UO_4473 (O_4473,N_48132,N_49714);
nand UO_4474 (O_4474,N_49611,N_49376);
and UO_4475 (O_4475,N_49176,N_47920);
xnor UO_4476 (O_4476,N_49253,N_48034);
nand UO_4477 (O_4477,N_49476,N_48882);
and UO_4478 (O_4478,N_48660,N_49677);
and UO_4479 (O_4479,N_49308,N_48923);
or UO_4480 (O_4480,N_49387,N_48708);
and UO_4481 (O_4481,N_47821,N_48833);
or UO_4482 (O_4482,N_48247,N_47735);
nand UO_4483 (O_4483,N_49462,N_47844);
nor UO_4484 (O_4484,N_47670,N_48675);
xnor UO_4485 (O_4485,N_49872,N_47628);
nand UO_4486 (O_4486,N_47523,N_48538);
and UO_4487 (O_4487,N_49968,N_49514);
xnor UO_4488 (O_4488,N_48889,N_47553);
nor UO_4489 (O_4489,N_48809,N_48235);
and UO_4490 (O_4490,N_49547,N_49178);
nand UO_4491 (O_4491,N_49494,N_47938);
nor UO_4492 (O_4492,N_48389,N_48383);
or UO_4493 (O_4493,N_49375,N_49359);
and UO_4494 (O_4494,N_48344,N_49908);
or UO_4495 (O_4495,N_47668,N_48930);
nor UO_4496 (O_4496,N_49372,N_48753);
nor UO_4497 (O_4497,N_49610,N_47803);
and UO_4498 (O_4498,N_48188,N_49332);
nor UO_4499 (O_4499,N_48327,N_49583);
xnor UO_4500 (O_4500,N_49409,N_48964);
nand UO_4501 (O_4501,N_49453,N_47629);
nand UO_4502 (O_4502,N_49176,N_49992);
xor UO_4503 (O_4503,N_47698,N_49739);
nand UO_4504 (O_4504,N_48636,N_48294);
or UO_4505 (O_4505,N_48937,N_49459);
or UO_4506 (O_4506,N_49223,N_49759);
and UO_4507 (O_4507,N_48949,N_47741);
or UO_4508 (O_4508,N_49410,N_49217);
xnor UO_4509 (O_4509,N_47766,N_47614);
nor UO_4510 (O_4510,N_49347,N_49714);
and UO_4511 (O_4511,N_48287,N_49488);
and UO_4512 (O_4512,N_49732,N_47902);
xnor UO_4513 (O_4513,N_48542,N_48307);
nor UO_4514 (O_4514,N_47864,N_49309);
and UO_4515 (O_4515,N_47599,N_47783);
and UO_4516 (O_4516,N_49307,N_47538);
nand UO_4517 (O_4517,N_49737,N_49825);
nor UO_4518 (O_4518,N_48678,N_48210);
nand UO_4519 (O_4519,N_49290,N_48196);
xnor UO_4520 (O_4520,N_49977,N_48604);
xor UO_4521 (O_4521,N_48241,N_48421);
or UO_4522 (O_4522,N_49220,N_47931);
xor UO_4523 (O_4523,N_49869,N_47786);
nor UO_4524 (O_4524,N_47996,N_47869);
xor UO_4525 (O_4525,N_49561,N_48506);
or UO_4526 (O_4526,N_49861,N_49761);
nor UO_4527 (O_4527,N_48490,N_48166);
xor UO_4528 (O_4528,N_49203,N_49218);
xor UO_4529 (O_4529,N_49799,N_49351);
xor UO_4530 (O_4530,N_49611,N_49508);
and UO_4531 (O_4531,N_49906,N_48904);
and UO_4532 (O_4532,N_49925,N_49613);
and UO_4533 (O_4533,N_49042,N_49365);
nor UO_4534 (O_4534,N_49366,N_47795);
xnor UO_4535 (O_4535,N_48129,N_49598);
or UO_4536 (O_4536,N_49544,N_49214);
nor UO_4537 (O_4537,N_48880,N_48429);
or UO_4538 (O_4538,N_47773,N_48597);
nand UO_4539 (O_4539,N_49016,N_49385);
nand UO_4540 (O_4540,N_48611,N_48346);
and UO_4541 (O_4541,N_48372,N_49127);
nor UO_4542 (O_4542,N_49224,N_49055);
or UO_4543 (O_4543,N_48708,N_48618);
xor UO_4544 (O_4544,N_47939,N_49638);
nand UO_4545 (O_4545,N_47635,N_48345);
and UO_4546 (O_4546,N_49467,N_49277);
nor UO_4547 (O_4547,N_47787,N_49405);
nor UO_4548 (O_4548,N_49764,N_49673);
xor UO_4549 (O_4549,N_49794,N_48681);
or UO_4550 (O_4550,N_49871,N_49738);
nand UO_4551 (O_4551,N_48259,N_48591);
and UO_4552 (O_4552,N_47859,N_48804);
nor UO_4553 (O_4553,N_48451,N_49938);
and UO_4554 (O_4554,N_48373,N_49859);
nor UO_4555 (O_4555,N_48722,N_49965);
and UO_4556 (O_4556,N_49771,N_49104);
nor UO_4557 (O_4557,N_49512,N_49222);
nor UO_4558 (O_4558,N_48592,N_47714);
nand UO_4559 (O_4559,N_48055,N_49195);
or UO_4560 (O_4560,N_47713,N_48562);
and UO_4561 (O_4561,N_49790,N_48358);
and UO_4562 (O_4562,N_48577,N_48010);
and UO_4563 (O_4563,N_49810,N_49323);
and UO_4564 (O_4564,N_48703,N_47796);
xor UO_4565 (O_4565,N_49607,N_47880);
nor UO_4566 (O_4566,N_47575,N_49907);
nor UO_4567 (O_4567,N_48342,N_49011);
nor UO_4568 (O_4568,N_47824,N_49486);
xnor UO_4569 (O_4569,N_47709,N_49451);
or UO_4570 (O_4570,N_47795,N_47675);
nor UO_4571 (O_4571,N_47697,N_47606);
and UO_4572 (O_4572,N_49793,N_48035);
and UO_4573 (O_4573,N_48802,N_47942);
or UO_4574 (O_4574,N_48713,N_49297);
and UO_4575 (O_4575,N_48793,N_49344);
or UO_4576 (O_4576,N_48308,N_49618);
or UO_4577 (O_4577,N_48779,N_49966);
xor UO_4578 (O_4578,N_49890,N_49880);
or UO_4579 (O_4579,N_49811,N_49884);
xnor UO_4580 (O_4580,N_49866,N_48485);
and UO_4581 (O_4581,N_48974,N_47927);
nor UO_4582 (O_4582,N_48832,N_48783);
or UO_4583 (O_4583,N_48366,N_48877);
xor UO_4584 (O_4584,N_48342,N_47870);
xnor UO_4585 (O_4585,N_49043,N_47651);
nand UO_4586 (O_4586,N_47565,N_48328);
and UO_4587 (O_4587,N_49455,N_48997);
and UO_4588 (O_4588,N_47610,N_48481);
and UO_4589 (O_4589,N_49395,N_48494);
nand UO_4590 (O_4590,N_47965,N_49758);
and UO_4591 (O_4591,N_49913,N_48688);
nor UO_4592 (O_4592,N_49224,N_48635);
nand UO_4593 (O_4593,N_49422,N_47643);
nand UO_4594 (O_4594,N_48529,N_48272);
xnor UO_4595 (O_4595,N_47542,N_49424);
and UO_4596 (O_4596,N_47592,N_49578);
xnor UO_4597 (O_4597,N_47686,N_47857);
or UO_4598 (O_4598,N_47529,N_49433);
and UO_4599 (O_4599,N_48591,N_49361);
nand UO_4600 (O_4600,N_49196,N_48442);
and UO_4601 (O_4601,N_49247,N_48801);
xnor UO_4602 (O_4602,N_49341,N_48875);
nand UO_4603 (O_4603,N_49165,N_47918);
or UO_4604 (O_4604,N_47931,N_47633);
or UO_4605 (O_4605,N_49401,N_49071);
and UO_4606 (O_4606,N_48327,N_48853);
xor UO_4607 (O_4607,N_47867,N_48865);
or UO_4608 (O_4608,N_49301,N_47536);
or UO_4609 (O_4609,N_49674,N_49315);
xor UO_4610 (O_4610,N_49847,N_49244);
xor UO_4611 (O_4611,N_47532,N_48127);
xnor UO_4612 (O_4612,N_49333,N_49432);
or UO_4613 (O_4613,N_49352,N_49550);
and UO_4614 (O_4614,N_49746,N_48091);
xor UO_4615 (O_4615,N_48099,N_48617);
nor UO_4616 (O_4616,N_48660,N_49980);
xnor UO_4617 (O_4617,N_48152,N_49996);
xor UO_4618 (O_4618,N_49241,N_49669);
xnor UO_4619 (O_4619,N_48952,N_48067);
nor UO_4620 (O_4620,N_48782,N_49881);
nor UO_4621 (O_4621,N_49846,N_48697);
and UO_4622 (O_4622,N_48009,N_49828);
nor UO_4623 (O_4623,N_47736,N_49731);
xor UO_4624 (O_4624,N_48290,N_48444);
nor UO_4625 (O_4625,N_48811,N_48459);
xnor UO_4626 (O_4626,N_49658,N_48767);
and UO_4627 (O_4627,N_49106,N_49198);
nand UO_4628 (O_4628,N_49175,N_48565);
and UO_4629 (O_4629,N_49605,N_49712);
nand UO_4630 (O_4630,N_49855,N_47716);
nor UO_4631 (O_4631,N_49873,N_48422);
xnor UO_4632 (O_4632,N_48450,N_48879);
nand UO_4633 (O_4633,N_49071,N_48536);
nor UO_4634 (O_4634,N_48575,N_47911);
or UO_4635 (O_4635,N_49326,N_48258);
nor UO_4636 (O_4636,N_49577,N_48614);
nor UO_4637 (O_4637,N_49777,N_47783);
and UO_4638 (O_4638,N_49243,N_49314);
nor UO_4639 (O_4639,N_48154,N_47502);
and UO_4640 (O_4640,N_48365,N_47816);
nand UO_4641 (O_4641,N_47993,N_49431);
xor UO_4642 (O_4642,N_49321,N_49291);
nand UO_4643 (O_4643,N_48138,N_48114);
nor UO_4644 (O_4644,N_47664,N_48918);
nand UO_4645 (O_4645,N_47966,N_47914);
xnor UO_4646 (O_4646,N_47884,N_48528);
or UO_4647 (O_4647,N_48405,N_49576);
and UO_4648 (O_4648,N_47856,N_49821);
xor UO_4649 (O_4649,N_48480,N_49962);
or UO_4650 (O_4650,N_49383,N_48379);
nor UO_4651 (O_4651,N_48880,N_47906);
and UO_4652 (O_4652,N_47986,N_49728);
nand UO_4653 (O_4653,N_48699,N_49167);
nand UO_4654 (O_4654,N_48956,N_49264);
xor UO_4655 (O_4655,N_49871,N_48147);
or UO_4656 (O_4656,N_49239,N_47791);
and UO_4657 (O_4657,N_49977,N_48437);
or UO_4658 (O_4658,N_49356,N_49476);
xnor UO_4659 (O_4659,N_49366,N_48988);
xnor UO_4660 (O_4660,N_49498,N_48034);
xor UO_4661 (O_4661,N_47945,N_48810);
or UO_4662 (O_4662,N_49167,N_49678);
xor UO_4663 (O_4663,N_48368,N_49724);
and UO_4664 (O_4664,N_49257,N_48955);
xor UO_4665 (O_4665,N_48770,N_49267);
nand UO_4666 (O_4666,N_47509,N_49923);
and UO_4667 (O_4667,N_47582,N_47638);
or UO_4668 (O_4668,N_49420,N_48677);
or UO_4669 (O_4669,N_48214,N_48475);
and UO_4670 (O_4670,N_49967,N_49123);
xnor UO_4671 (O_4671,N_49172,N_49506);
nor UO_4672 (O_4672,N_48279,N_47516);
or UO_4673 (O_4673,N_49951,N_48863);
xor UO_4674 (O_4674,N_48541,N_49053);
and UO_4675 (O_4675,N_47695,N_49033);
nand UO_4676 (O_4676,N_49077,N_48993);
nand UO_4677 (O_4677,N_49053,N_49844);
xor UO_4678 (O_4678,N_49315,N_49524);
xor UO_4679 (O_4679,N_49580,N_48669);
xnor UO_4680 (O_4680,N_47554,N_49261);
or UO_4681 (O_4681,N_47800,N_49474);
nor UO_4682 (O_4682,N_49990,N_48867);
and UO_4683 (O_4683,N_49708,N_48563);
nand UO_4684 (O_4684,N_48409,N_48429);
or UO_4685 (O_4685,N_49929,N_48988);
or UO_4686 (O_4686,N_49914,N_47814);
and UO_4687 (O_4687,N_49521,N_48133);
or UO_4688 (O_4688,N_48899,N_49599);
or UO_4689 (O_4689,N_49905,N_49880);
xnor UO_4690 (O_4690,N_48015,N_49214);
or UO_4691 (O_4691,N_47761,N_47546);
and UO_4692 (O_4692,N_49815,N_48094);
or UO_4693 (O_4693,N_48599,N_48281);
or UO_4694 (O_4694,N_49247,N_48810);
or UO_4695 (O_4695,N_49748,N_48337);
xor UO_4696 (O_4696,N_48194,N_49320);
nor UO_4697 (O_4697,N_47565,N_48521);
nand UO_4698 (O_4698,N_47725,N_49104);
nor UO_4699 (O_4699,N_48743,N_49047);
nand UO_4700 (O_4700,N_48199,N_48956);
or UO_4701 (O_4701,N_49380,N_47660);
or UO_4702 (O_4702,N_49484,N_48448);
nand UO_4703 (O_4703,N_48608,N_49507);
and UO_4704 (O_4704,N_49250,N_49505);
xor UO_4705 (O_4705,N_49186,N_47712);
xor UO_4706 (O_4706,N_49700,N_49491);
nand UO_4707 (O_4707,N_48902,N_49406);
nor UO_4708 (O_4708,N_48374,N_48135);
nand UO_4709 (O_4709,N_48961,N_49131);
nand UO_4710 (O_4710,N_49102,N_48817);
nand UO_4711 (O_4711,N_49765,N_49503);
and UO_4712 (O_4712,N_48616,N_47836);
nand UO_4713 (O_4713,N_48509,N_49163);
nor UO_4714 (O_4714,N_47583,N_49218);
and UO_4715 (O_4715,N_49181,N_49709);
and UO_4716 (O_4716,N_49022,N_48092);
and UO_4717 (O_4717,N_48159,N_48058);
and UO_4718 (O_4718,N_48795,N_49955);
and UO_4719 (O_4719,N_48391,N_47855);
nor UO_4720 (O_4720,N_48586,N_49829);
and UO_4721 (O_4721,N_48189,N_47946);
nand UO_4722 (O_4722,N_49083,N_48410);
nand UO_4723 (O_4723,N_49828,N_49420);
nand UO_4724 (O_4724,N_48963,N_49389);
or UO_4725 (O_4725,N_48366,N_47595);
xor UO_4726 (O_4726,N_49984,N_49951);
nand UO_4727 (O_4727,N_49041,N_47950);
or UO_4728 (O_4728,N_47996,N_49350);
or UO_4729 (O_4729,N_49614,N_49572);
and UO_4730 (O_4730,N_48203,N_47807);
and UO_4731 (O_4731,N_49228,N_48344);
and UO_4732 (O_4732,N_48146,N_49400);
and UO_4733 (O_4733,N_49494,N_48235);
or UO_4734 (O_4734,N_49973,N_49319);
nand UO_4735 (O_4735,N_48662,N_47563);
xor UO_4736 (O_4736,N_48049,N_48358);
xor UO_4737 (O_4737,N_47525,N_49748);
or UO_4738 (O_4738,N_48431,N_49995);
nor UO_4739 (O_4739,N_47811,N_48468);
xnor UO_4740 (O_4740,N_49583,N_48658);
and UO_4741 (O_4741,N_47986,N_49150);
nand UO_4742 (O_4742,N_48189,N_47533);
xnor UO_4743 (O_4743,N_49738,N_49111);
or UO_4744 (O_4744,N_49828,N_49209);
and UO_4745 (O_4745,N_49843,N_47885);
and UO_4746 (O_4746,N_48479,N_48706);
and UO_4747 (O_4747,N_48752,N_48014);
and UO_4748 (O_4748,N_49802,N_49565);
or UO_4749 (O_4749,N_48517,N_48741);
nor UO_4750 (O_4750,N_48151,N_49657);
xor UO_4751 (O_4751,N_47630,N_49366);
or UO_4752 (O_4752,N_49220,N_49805);
nand UO_4753 (O_4753,N_49555,N_48794);
nand UO_4754 (O_4754,N_48670,N_47825);
nor UO_4755 (O_4755,N_49163,N_49707);
nand UO_4756 (O_4756,N_47608,N_47540);
or UO_4757 (O_4757,N_49877,N_49097);
xnor UO_4758 (O_4758,N_48917,N_48270);
nor UO_4759 (O_4759,N_47546,N_48547);
nor UO_4760 (O_4760,N_48905,N_48607);
nor UO_4761 (O_4761,N_49674,N_47521);
or UO_4762 (O_4762,N_48165,N_48836);
xnor UO_4763 (O_4763,N_47789,N_49849);
and UO_4764 (O_4764,N_47554,N_47834);
and UO_4765 (O_4765,N_49723,N_47645);
or UO_4766 (O_4766,N_47561,N_47596);
or UO_4767 (O_4767,N_48419,N_49982);
or UO_4768 (O_4768,N_47852,N_49925);
and UO_4769 (O_4769,N_48945,N_48855);
nor UO_4770 (O_4770,N_48772,N_49620);
xor UO_4771 (O_4771,N_48410,N_49267);
and UO_4772 (O_4772,N_49663,N_48682);
or UO_4773 (O_4773,N_48738,N_47844);
xor UO_4774 (O_4774,N_49576,N_49007);
or UO_4775 (O_4775,N_47666,N_48216);
nor UO_4776 (O_4776,N_49417,N_49307);
xnor UO_4777 (O_4777,N_48846,N_49432);
nand UO_4778 (O_4778,N_49256,N_47971);
xor UO_4779 (O_4779,N_49125,N_47725);
nor UO_4780 (O_4780,N_48314,N_48962);
nand UO_4781 (O_4781,N_49486,N_49937);
or UO_4782 (O_4782,N_49752,N_48219);
and UO_4783 (O_4783,N_49035,N_47675);
or UO_4784 (O_4784,N_49565,N_48305);
nor UO_4785 (O_4785,N_48012,N_47663);
xnor UO_4786 (O_4786,N_47516,N_47630);
or UO_4787 (O_4787,N_49933,N_48807);
nand UO_4788 (O_4788,N_49094,N_47751);
nand UO_4789 (O_4789,N_48314,N_49277);
or UO_4790 (O_4790,N_48075,N_48659);
nor UO_4791 (O_4791,N_47562,N_49709);
xor UO_4792 (O_4792,N_48458,N_49151);
or UO_4793 (O_4793,N_47798,N_47947);
or UO_4794 (O_4794,N_48383,N_48997);
nand UO_4795 (O_4795,N_49610,N_47808);
nor UO_4796 (O_4796,N_49441,N_47767);
nor UO_4797 (O_4797,N_48629,N_48737);
or UO_4798 (O_4798,N_47665,N_49392);
nor UO_4799 (O_4799,N_49703,N_48016);
nor UO_4800 (O_4800,N_48926,N_47556);
nor UO_4801 (O_4801,N_49896,N_48403);
nand UO_4802 (O_4802,N_49803,N_49541);
xnor UO_4803 (O_4803,N_48978,N_49670);
nor UO_4804 (O_4804,N_48828,N_49881);
nor UO_4805 (O_4805,N_48342,N_47543);
nor UO_4806 (O_4806,N_48404,N_49395);
nor UO_4807 (O_4807,N_48795,N_48291);
nor UO_4808 (O_4808,N_48746,N_49298);
nand UO_4809 (O_4809,N_49697,N_48207);
nor UO_4810 (O_4810,N_49383,N_49600);
nand UO_4811 (O_4811,N_48610,N_48216);
and UO_4812 (O_4812,N_48711,N_49070);
and UO_4813 (O_4813,N_49652,N_47834);
or UO_4814 (O_4814,N_48592,N_48041);
nand UO_4815 (O_4815,N_49138,N_48324);
or UO_4816 (O_4816,N_48157,N_48140);
or UO_4817 (O_4817,N_49480,N_48647);
xor UO_4818 (O_4818,N_49829,N_49077);
xor UO_4819 (O_4819,N_49438,N_48337);
and UO_4820 (O_4820,N_48464,N_47699);
nand UO_4821 (O_4821,N_48593,N_47502);
or UO_4822 (O_4822,N_49100,N_48572);
and UO_4823 (O_4823,N_48217,N_48808);
and UO_4824 (O_4824,N_48147,N_47512);
nor UO_4825 (O_4825,N_47752,N_48417);
and UO_4826 (O_4826,N_49209,N_47908);
nand UO_4827 (O_4827,N_49153,N_48751);
or UO_4828 (O_4828,N_48863,N_49818);
nor UO_4829 (O_4829,N_48628,N_47675);
nand UO_4830 (O_4830,N_49490,N_48549);
nand UO_4831 (O_4831,N_48421,N_48032);
or UO_4832 (O_4832,N_49688,N_49968);
xnor UO_4833 (O_4833,N_47616,N_48321);
or UO_4834 (O_4834,N_48017,N_49231);
nand UO_4835 (O_4835,N_49838,N_49272);
or UO_4836 (O_4836,N_49055,N_48985);
or UO_4837 (O_4837,N_49958,N_47822);
and UO_4838 (O_4838,N_48660,N_49230);
nor UO_4839 (O_4839,N_47770,N_48417);
and UO_4840 (O_4840,N_47646,N_47569);
and UO_4841 (O_4841,N_48443,N_48822);
and UO_4842 (O_4842,N_49050,N_49422);
and UO_4843 (O_4843,N_49551,N_49078);
xnor UO_4844 (O_4844,N_47646,N_49350);
nor UO_4845 (O_4845,N_47847,N_47993);
xor UO_4846 (O_4846,N_48649,N_48730);
nor UO_4847 (O_4847,N_48551,N_48270);
nor UO_4848 (O_4848,N_47912,N_49479);
or UO_4849 (O_4849,N_49877,N_47956);
or UO_4850 (O_4850,N_49554,N_48092);
or UO_4851 (O_4851,N_47567,N_48390);
and UO_4852 (O_4852,N_49785,N_48364);
nand UO_4853 (O_4853,N_49405,N_47508);
nor UO_4854 (O_4854,N_48594,N_47681);
nor UO_4855 (O_4855,N_48178,N_47754);
nor UO_4856 (O_4856,N_48122,N_49063);
nor UO_4857 (O_4857,N_47503,N_48171);
or UO_4858 (O_4858,N_48065,N_49789);
and UO_4859 (O_4859,N_48377,N_47863);
nand UO_4860 (O_4860,N_48766,N_49347);
and UO_4861 (O_4861,N_49305,N_48740);
xor UO_4862 (O_4862,N_48315,N_47653);
nand UO_4863 (O_4863,N_48469,N_47772);
or UO_4864 (O_4864,N_47557,N_48207);
nand UO_4865 (O_4865,N_47974,N_47844);
or UO_4866 (O_4866,N_48284,N_49035);
nand UO_4867 (O_4867,N_48067,N_47684);
nor UO_4868 (O_4868,N_48507,N_48367);
nor UO_4869 (O_4869,N_48406,N_49395);
or UO_4870 (O_4870,N_49665,N_47501);
nor UO_4871 (O_4871,N_49878,N_48434);
or UO_4872 (O_4872,N_49799,N_47616);
nand UO_4873 (O_4873,N_49514,N_49675);
or UO_4874 (O_4874,N_47763,N_48161);
and UO_4875 (O_4875,N_49814,N_48879);
or UO_4876 (O_4876,N_48870,N_47648);
or UO_4877 (O_4877,N_48928,N_48981);
or UO_4878 (O_4878,N_49458,N_49731);
or UO_4879 (O_4879,N_49492,N_49158);
nand UO_4880 (O_4880,N_49293,N_47991);
and UO_4881 (O_4881,N_48602,N_48469);
nand UO_4882 (O_4882,N_49946,N_47914);
nand UO_4883 (O_4883,N_48292,N_48223);
and UO_4884 (O_4884,N_49048,N_47643);
nor UO_4885 (O_4885,N_49685,N_47560);
xnor UO_4886 (O_4886,N_48373,N_49703);
or UO_4887 (O_4887,N_48347,N_48608);
nand UO_4888 (O_4888,N_48482,N_48233);
nand UO_4889 (O_4889,N_49653,N_49763);
nand UO_4890 (O_4890,N_48113,N_48591);
nand UO_4891 (O_4891,N_48335,N_49140);
or UO_4892 (O_4892,N_47577,N_48447);
and UO_4893 (O_4893,N_47641,N_48940);
and UO_4894 (O_4894,N_49808,N_48940);
or UO_4895 (O_4895,N_47917,N_48218);
or UO_4896 (O_4896,N_49603,N_49937);
xor UO_4897 (O_4897,N_48298,N_49893);
and UO_4898 (O_4898,N_49422,N_49775);
and UO_4899 (O_4899,N_48413,N_49601);
xnor UO_4900 (O_4900,N_49558,N_49190);
or UO_4901 (O_4901,N_49358,N_49278);
xnor UO_4902 (O_4902,N_47695,N_49512);
nand UO_4903 (O_4903,N_49369,N_48014);
nor UO_4904 (O_4904,N_48491,N_49759);
nand UO_4905 (O_4905,N_47955,N_47790);
or UO_4906 (O_4906,N_48074,N_47513);
nand UO_4907 (O_4907,N_48020,N_49519);
and UO_4908 (O_4908,N_48791,N_49164);
or UO_4909 (O_4909,N_47883,N_48653);
and UO_4910 (O_4910,N_48116,N_48612);
nor UO_4911 (O_4911,N_49926,N_49873);
nand UO_4912 (O_4912,N_49725,N_48938);
or UO_4913 (O_4913,N_48420,N_48211);
xor UO_4914 (O_4914,N_48882,N_49560);
or UO_4915 (O_4915,N_48437,N_47906);
or UO_4916 (O_4916,N_48270,N_47855);
or UO_4917 (O_4917,N_49826,N_48512);
nor UO_4918 (O_4918,N_49235,N_48351);
xnor UO_4919 (O_4919,N_47530,N_49380);
nor UO_4920 (O_4920,N_47877,N_47967);
and UO_4921 (O_4921,N_48928,N_49876);
xnor UO_4922 (O_4922,N_47549,N_49629);
xnor UO_4923 (O_4923,N_49316,N_49397);
nor UO_4924 (O_4924,N_47953,N_49338);
nand UO_4925 (O_4925,N_48597,N_47814);
and UO_4926 (O_4926,N_47951,N_49954);
and UO_4927 (O_4927,N_49125,N_49734);
and UO_4928 (O_4928,N_49679,N_49532);
and UO_4929 (O_4929,N_47501,N_49641);
nor UO_4930 (O_4930,N_49596,N_47965);
xnor UO_4931 (O_4931,N_48869,N_47711);
xor UO_4932 (O_4932,N_48420,N_48707);
nand UO_4933 (O_4933,N_49465,N_48901);
or UO_4934 (O_4934,N_49312,N_49145);
nand UO_4935 (O_4935,N_47828,N_48491);
nand UO_4936 (O_4936,N_48070,N_48472);
xnor UO_4937 (O_4937,N_48886,N_48603);
nand UO_4938 (O_4938,N_48226,N_49627);
and UO_4939 (O_4939,N_49941,N_48920);
or UO_4940 (O_4940,N_48890,N_48623);
nor UO_4941 (O_4941,N_49505,N_48305);
nand UO_4942 (O_4942,N_47772,N_49005);
xor UO_4943 (O_4943,N_48935,N_49780);
nand UO_4944 (O_4944,N_49306,N_48200);
nor UO_4945 (O_4945,N_49079,N_48882);
or UO_4946 (O_4946,N_49860,N_48477);
nand UO_4947 (O_4947,N_47973,N_48435);
xnor UO_4948 (O_4948,N_48613,N_49109);
xor UO_4949 (O_4949,N_48476,N_48154);
or UO_4950 (O_4950,N_49922,N_47810);
nor UO_4951 (O_4951,N_48042,N_48074);
nand UO_4952 (O_4952,N_48924,N_49025);
nor UO_4953 (O_4953,N_49374,N_47919);
xnor UO_4954 (O_4954,N_49531,N_48739);
or UO_4955 (O_4955,N_49656,N_47815);
or UO_4956 (O_4956,N_47722,N_48661);
nor UO_4957 (O_4957,N_48571,N_49990);
and UO_4958 (O_4958,N_47749,N_47544);
nand UO_4959 (O_4959,N_49931,N_48513);
nor UO_4960 (O_4960,N_47599,N_47692);
and UO_4961 (O_4961,N_49973,N_48586);
xor UO_4962 (O_4962,N_48784,N_47893);
nor UO_4963 (O_4963,N_49359,N_48948);
or UO_4964 (O_4964,N_49668,N_48516);
or UO_4965 (O_4965,N_49613,N_49795);
and UO_4966 (O_4966,N_47759,N_48872);
nand UO_4967 (O_4967,N_48420,N_49479);
xnor UO_4968 (O_4968,N_49702,N_49223);
nand UO_4969 (O_4969,N_49915,N_48654);
nor UO_4970 (O_4970,N_49938,N_49576);
and UO_4971 (O_4971,N_49667,N_47787);
or UO_4972 (O_4972,N_47946,N_48506);
nor UO_4973 (O_4973,N_48544,N_48465);
xnor UO_4974 (O_4974,N_48449,N_48418);
xor UO_4975 (O_4975,N_48143,N_48173);
nor UO_4976 (O_4976,N_48251,N_49646);
nand UO_4977 (O_4977,N_49898,N_49316);
nor UO_4978 (O_4978,N_47971,N_49261);
nand UO_4979 (O_4979,N_48346,N_48735);
xor UO_4980 (O_4980,N_47558,N_48545);
xor UO_4981 (O_4981,N_48028,N_48702);
nor UO_4982 (O_4982,N_47582,N_47773);
or UO_4983 (O_4983,N_47699,N_48064);
nand UO_4984 (O_4984,N_48757,N_48957);
and UO_4985 (O_4985,N_49957,N_48036);
xnor UO_4986 (O_4986,N_47780,N_49528);
or UO_4987 (O_4987,N_49497,N_47758);
or UO_4988 (O_4988,N_47771,N_49053);
nand UO_4989 (O_4989,N_48636,N_47752);
xnor UO_4990 (O_4990,N_47541,N_48368);
nand UO_4991 (O_4991,N_47985,N_49991);
xnor UO_4992 (O_4992,N_48358,N_48809);
or UO_4993 (O_4993,N_48978,N_47874);
xor UO_4994 (O_4994,N_48088,N_49802);
nor UO_4995 (O_4995,N_48084,N_49372);
nor UO_4996 (O_4996,N_48885,N_48343);
or UO_4997 (O_4997,N_49766,N_48163);
or UO_4998 (O_4998,N_47795,N_49599);
nor UO_4999 (O_4999,N_47719,N_47919);
endmodule