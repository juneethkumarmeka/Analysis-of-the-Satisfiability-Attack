module basic_2500_25000_3000_20_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_500,In_1795);
or U1 (N_1,In_2485,In_1519);
nand U2 (N_2,In_1417,In_390);
or U3 (N_3,In_511,In_251);
nor U4 (N_4,In_881,In_862);
or U5 (N_5,In_2258,In_1830);
nor U6 (N_6,In_2094,In_766);
or U7 (N_7,In_425,In_1171);
nand U8 (N_8,In_1527,In_2474);
xnor U9 (N_9,In_1266,In_1054);
and U10 (N_10,In_295,In_768);
and U11 (N_11,In_314,In_1977);
nor U12 (N_12,In_1227,In_1345);
nand U13 (N_13,In_2452,In_683);
and U14 (N_14,In_381,In_1604);
nor U15 (N_15,In_1620,In_2174);
xnor U16 (N_16,In_1837,In_1908);
nor U17 (N_17,In_576,In_859);
or U18 (N_18,In_1759,In_45);
and U19 (N_19,In_1636,In_1191);
or U20 (N_20,In_445,In_1913);
or U21 (N_21,In_312,In_586);
nand U22 (N_22,In_955,In_814);
and U23 (N_23,In_206,In_2017);
or U24 (N_24,In_578,In_2206);
nand U25 (N_25,In_1673,In_2427);
or U26 (N_26,In_1244,In_2337);
xor U27 (N_27,In_1972,In_49);
or U28 (N_28,In_374,In_310);
nor U29 (N_29,In_866,In_948);
or U30 (N_30,In_156,In_1066);
nor U31 (N_31,In_1863,In_1755);
or U32 (N_32,In_2104,In_2053);
nor U33 (N_33,In_1089,In_907);
nor U34 (N_34,In_272,In_2481);
nand U35 (N_35,In_2019,In_2272);
nor U36 (N_36,In_1707,In_1524);
xnor U37 (N_37,In_404,In_644);
and U38 (N_38,In_228,In_723);
or U39 (N_39,In_2252,In_595);
or U40 (N_40,In_707,In_599);
or U41 (N_41,In_136,In_983);
or U42 (N_42,In_2298,In_1333);
nand U43 (N_43,In_639,In_1176);
nor U44 (N_44,In_1082,In_491);
nor U45 (N_45,In_1923,In_575);
nand U46 (N_46,In_372,In_638);
nand U47 (N_47,In_2290,In_171);
and U48 (N_48,In_29,In_1009);
and U49 (N_49,In_188,In_232);
or U50 (N_50,In_761,In_973);
or U51 (N_51,In_564,In_2410);
nor U52 (N_52,In_1985,In_1563);
or U53 (N_53,In_2181,In_2393);
or U54 (N_54,In_468,In_2407);
nor U55 (N_55,In_2242,In_773);
and U56 (N_56,In_841,In_1570);
or U57 (N_57,In_914,In_622);
or U58 (N_58,In_598,In_2059);
nand U59 (N_59,In_223,In_79);
and U60 (N_60,In_642,In_2120);
nand U61 (N_61,In_2421,In_1632);
and U62 (N_62,In_1271,In_1617);
or U63 (N_63,In_884,In_158);
nor U64 (N_64,In_1722,In_2036);
nand U65 (N_65,In_1316,In_516);
nor U66 (N_66,In_1767,In_1646);
and U67 (N_67,In_2433,In_1926);
nand U68 (N_68,In_257,In_2003);
xnor U69 (N_69,In_498,In_679);
and U70 (N_70,In_967,In_918);
nand U71 (N_71,In_1145,In_2256);
or U72 (N_72,In_180,In_711);
or U73 (N_73,In_261,In_2346);
and U74 (N_74,In_1373,In_2005);
xor U75 (N_75,In_1700,In_1609);
xnor U76 (N_76,In_1403,In_406);
xor U77 (N_77,In_2445,In_1576);
xnor U78 (N_78,In_1947,In_2032);
or U79 (N_79,In_1588,In_1971);
or U80 (N_80,In_1282,In_2418);
nor U81 (N_81,In_1812,In_1553);
and U82 (N_82,In_1813,In_615);
nand U83 (N_83,In_2226,In_1615);
xnor U84 (N_84,In_1583,In_1849);
and U85 (N_85,In_702,In_538);
xnor U86 (N_86,In_1446,In_2330);
or U87 (N_87,In_1018,In_551);
nand U88 (N_88,In_1859,In_2498);
xor U89 (N_89,In_1442,In_926);
and U90 (N_90,In_1199,In_1855);
nor U91 (N_91,In_1091,In_1735);
and U92 (N_92,In_966,In_1818);
xor U93 (N_93,In_2012,In_360);
and U94 (N_94,In_1535,In_1703);
or U95 (N_95,In_1478,In_1106);
nand U96 (N_96,In_2083,In_376);
nor U97 (N_97,In_1851,In_2268);
nand U98 (N_98,In_623,In_910);
nand U99 (N_99,In_1844,In_2113);
nor U100 (N_100,In_661,In_852);
nor U101 (N_101,In_1674,In_1090);
nor U102 (N_102,In_1892,In_799);
and U103 (N_103,In_2428,In_1876);
and U104 (N_104,In_1183,In_2297);
xor U105 (N_105,In_2227,In_1189);
and U106 (N_106,In_958,In_552);
xor U107 (N_107,In_2231,In_1860);
nor U108 (N_108,In_1410,In_262);
and U109 (N_109,In_2187,In_2143);
or U110 (N_110,In_115,In_1888);
nor U111 (N_111,In_1815,In_978);
xnor U112 (N_112,In_1838,In_659);
nand U113 (N_113,In_1575,In_450);
and U114 (N_114,In_1224,In_2473);
nand U115 (N_115,In_2098,In_1081);
or U116 (N_116,In_1668,In_113);
or U117 (N_117,In_1079,In_2063);
or U118 (N_118,In_1612,In_747);
nand U119 (N_119,In_1414,In_1243);
and U120 (N_120,In_484,In_2049);
or U121 (N_121,In_1980,In_1672);
nand U122 (N_122,In_1026,In_1044);
nor U123 (N_123,In_1267,In_1301);
nand U124 (N_124,In_2347,In_1623);
xnor U125 (N_125,In_1512,In_2236);
or U126 (N_126,In_1823,In_413);
xnor U127 (N_127,In_1115,In_656);
xor U128 (N_128,In_351,In_2207);
and U129 (N_129,In_986,In_1577);
nor U130 (N_130,In_2399,In_2369);
or U131 (N_131,In_2025,In_2487);
xor U132 (N_132,In_1829,In_1470);
or U133 (N_133,In_1149,In_1146);
and U134 (N_134,In_1175,In_142);
nor U135 (N_135,In_2095,In_811);
nor U136 (N_136,In_728,In_31);
and U137 (N_137,In_2026,In_2101);
and U138 (N_138,In_1297,In_1537);
nand U139 (N_139,In_1702,In_2156);
or U140 (N_140,In_1928,In_1393);
nand U141 (N_141,In_1756,In_867);
nand U142 (N_142,In_1877,In_807);
xnor U143 (N_143,In_545,In_1704);
nor U144 (N_144,In_132,In_808);
and U145 (N_145,In_209,In_2130);
nand U146 (N_146,In_1174,In_2129);
nor U147 (N_147,In_1371,In_782);
and U148 (N_148,In_2315,In_1508);
and U149 (N_149,In_2189,In_1135);
and U150 (N_150,In_729,In_774);
or U151 (N_151,In_2389,In_621);
nand U152 (N_152,In_1606,In_2117);
nand U153 (N_153,In_1313,In_488);
xnor U154 (N_154,In_1254,In_449);
nor U155 (N_155,In_663,In_1596);
and U156 (N_156,In_410,In_1430);
nor U157 (N_157,In_1987,In_2230);
nor U158 (N_158,In_624,In_2416);
or U159 (N_159,In_467,In_1480);
nand U160 (N_160,In_178,In_522);
xor U161 (N_161,In_1386,In_1994);
nand U162 (N_162,In_2169,In_1320);
or U163 (N_163,In_2397,In_444);
and U164 (N_164,In_1083,In_509);
nor U165 (N_165,In_1151,In_9);
nor U166 (N_166,In_1685,In_1486);
nand U167 (N_167,In_980,In_1852);
or U168 (N_168,In_1825,In_1328);
and U169 (N_169,In_2106,In_1275);
or U170 (N_170,In_1692,In_474);
nor U171 (N_171,In_1073,In_377);
nor U172 (N_172,In_1317,In_704);
xnor U173 (N_173,In_668,In_632);
or U174 (N_174,In_739,In_101);
or U175 (N_175,In_2470,In_230);
and U176 (N_176,In_1148,In_1188);
nor U177 (N_177,In_181,In_2341);
nor U178 (N_178,In_529,In_327);
or U179 (N_179,In_1920,In_340);
xor U180 (N_180,In_1758,In_781);
xnor U181 (N_181,In_585,In_2304);
and U182 (N_182,In_3,In_60);
xor U183 (N_183,In_1228,In_890);
nor U184 (N_184,In_588,In_2343);
xnor U185 (N_185,In_2205,In_85);
or U186 (N_186,In_959,In_836);
xnor U187 (N_187,In_416,In_18);
nor U188 (N_188,In_458,In_665);
nor U189 (N_189,In_1868,In_1826);
nor U190 (N_190,In_87,In_2327);
nor U191 (N_191,In_2072,In_682);
and U192 (N_192,In_1551,In_2411);
nand U193 (N_193,In_893,In_160);
xor U194 (N_194,In_1638,In_2050);
nand U195 (N_195,In_1719,In_804);
xor U196 (N_196,In_2224,In_482);
and U197 (N_197,In_721,In_1717);
or U198 (N_198,In_645,In_1727);
xor U199 (N_199,In_2334,In_851);
nor U200 (N_200,In_350,In_2111);
nand U201 (N_201,In_647,In_74);
xor U202 (N_202,In_250,In_1491);
xor U203 (N_203,In_985,In_186);
and U204 (N_204,In_1233,In_2387);
or U205 (N_205,In_1593,In_428);
nand U206 (N_206,In_1982,In_987);
nand U207 (N_207,In_1421,In_903);
xnor U208 (N_208,In_1862,In_119);
xnor U209 (N_209,In_547,In_1520);
or U210 (N_210,In_1235,In_438);
nand U211 (N_211,In_1732,In_846);
and U212 (N_212,In_818,In_2405);
or U213 (N_213,In_1314,In_2430);
nand U214 (N_214,In_1016,In_935);
xnor U215 (N_215,In_50,In_1900);
xnor U216 (N_216,In_1602,In_195);
and U217 (N_217,In_238,In_790);
nand U218 (N_218,In_76,In_1751);
nand U219 (N_219,In_1781,In_199);
and U220 (N_220,In_1626,In_941);
nand U221 (N_221,In_651,In_1634);
xor U222 (N_222,In_464,In_2089);
or U223 (N_223,In_1348,In_969);
or U224 (N_224,In_453,In_1680);
nand U225 (N_225,In_1821,In_1912);
xnor U226 (N_226,In_2042,In_1848);
or U227 (N_227,In_752,In_686);
nand U228 (N_228,In_362,In_1810);
and U229 (N_229,In_972,In_57);
nor U230 (N_230,In_722,In_288);
nand U231 (N_231,In_1598,In_145);
xnor U232 (N_232,In_524,In_950);
nand U233 (N_233,In_1045,In_2168);
nand U234 (N_234,In_892,In_2426);
nand U235 (N_235,In_2008,In_2028);
nor U236 (N_236,In_2177,In_1773);
and U237 (N_237,In_777,In_213);
and U238 (N_238,In_845,In_2340);
and U239 (N_239,In_1204,In_2463);
nand U240 (N_240,In_394,In_1058);
xor U241 (N_241,In_681,In_714);
nor U242 (N_242,In_324,In_1032);
or U243 (N_243,In_1212,In_363);
or U244 (N_244,In_1681,In_2489);
or U245 (N_245,In_5,In_1565);
xor U246 (N_246,In_1622,In_889);
and U247 (N_247,In_258,In_2192);
or U248 (N_248,In_337,In_2217);
nand U249 (N_249,In_205,In_1041);
and U250 (N_250,In_717,In_2375);
xor U251 (N_251,In_2161,In_1178);
or U252 (N_252,In_22,In_326);
or U253 (N_253,In_1714,In_1768);
xor U254 (N_254,In_554,In_1276);
xor U255 (N_255,In_2066,In_202);
and U256 (N_256,In_2404,In_2110);
xor U257 (N_257,In_1656,In_2237);
xnor U258 (N_258,In_741,In_1578);
or U259 (N_259,In_103,In_2408);
or U260 (N_260,In_1745,In_179);
xnor U261 (N_261,In_2382,In_2204);
xor U262 (N_262,In_55,In_124);
and U263 (N_263,In_1422,In_2173);
nor U264 (N_264,In_123,In_2287);
and U265 (N_265,In_42,In_1841);
xor U266 (N_266,In_2317,In_541);
or U267 (N_267,In_1407,In_1186);
nor U268 (N_268,In_1309,In_2491);
nor U269 (N_269,In_1654,In_2086);
or U270 (N_270,In_1062,In_203);
or U271 (N_271,In_2071,In_749);
or U272 (N_272,In_1299,In_131);
or U273 (N_273,In_877,In_1479);
nand U274 (N_274,In_71,In_2260);
nor U275 (N_275,In_442,In_150);
and U276 (N_276,In_830,In_1419);
xnor U277 (N_277,In_190,In_1644);
nand U278 (N_278,In_2048,In_356);
and U279 (N_279,In_117,In_2141);
and U280 (N_280,In_1213,In_1500);
or U281 (N_281,In_2372,In_1774);
xor U282 (N_282,In_2447,In_1805);
nand U283 (N_283,In_1101,In_1302);
and U284 (N_284,In_2475,In_1440);
xor U285 (N_285,In_701,In_791);
nor U286 (N_286,In_1963,In_1725);
nor U287 (N_287,In_2085,In_2184);
nand U288 (N_288,In_330,In_307);
nand U289 (N_289,In_405,In_2185);
and U290 (N_290,In_1950,In_225);
xor U291 (N_291,In_151,In_1064);
and U292 (N_292,In_1540,In_838);
or U293 (N_293,In_2151,In_1181);
xor U294 (N_294,In_2370,In_2444);
or U295 (N_295,In_796,In_2203);
nor U296 (N_296,In_1984,In_993);
and U297 (N_297,In_2229,In_1449);
or U298 (N_298,In_1765,In_279);
nand U299 (N_299,In_1516,In_125);
and U300 (N_300,In_1902,In_408);
xnor U301 (N_301,In_162,In_154);
and U302 (N_302,In_2412,In_1701);
and U303 (N_303,In_1318,In_1836);
nor U304 (N_304,In_418,In_1285);
or U305 (N_305,In_2209,In_2016);
nor U306 (N_306,In_1010,In_1840);
and U307 (N_307,In_2270,In_557);
nor U308 (N_308,In_1803,In_100);
nor U309 (N_309,In_107,In_1200);
and U310 (N_310,In_1358,In_118);
and U311 (N_311,In_2241,In_1433);
nand U312 (N_312,In_17,In_2326);
xor U313 (N_313,In_1651,In_1791);
and U314 (N_314,In_420,In_692);
or U315 (N_315,In_610,In_1720);
xnor U316 (N_316,In_1214,In_1988);
nor U317 (N_317,In_765,In_1435);
and U318 (N_318,In_1772,In_2265);
nand U319 (N_319,In_1391,In_515);
nor U320 (N_320,In_2179,In_1931);
and U321 (N_321,In_1990,In_865);
nand U322 (N_322,In_2090,In_2157);
and U323 (N_323,In_2220,In_135);
nor U324 (N_324,In_1890,In_2312);
nor U325 (N_325,In_1517,In_1069);
nor U326 (N_326,In_1601,In_508);
nor U327 (N_327,In_2022,In_1635);
or U328 (N_328,In_1409,In_887);
or U329 (N_329,In_380,In_1322);
xor U330 (N_330,In_748,In_2001);
nor U331 (N_331,In_1019,In_1589);
or U332 (N_332,In_15,In_1143);
or U333 (N_333,In_1341,In_591);
or U334 (N_334,In_842,In_2009);
nand U335 (N_335,In_1363,In_1682);
or U336 (N_336,In_1154,In_253);
or U337 (N_337,In_684,In_2323);
and U338 (N_338,In_2103,In_367);
nand U339 (N_339,In_2118,In_412);
xnor U340 (N_340,In_1724,In_1441);
nand U341 (N_341,In_1690,In_580);
and U342 (N_342,In_1997,In_1142);
nand U343 (N_343,In_1108,In_1071);
or U344 (N_344,In_1377,In_664);
and U345 (N_345,In_2394,In_1780);
nor U346 (N_346,In_2422,In_1802);
or U347 (N_347,In_1922,In_1037);
and U348 (N_348,In_2044,In_2194);
xnor U349 (N_349,In_1933,In_587);
nand U350 (N_350,In_1878,In_1014);
nor U351 (N_351,In_2222,In_2338);
nor U352 (N_352,In_1484,In_1956);
and U353 (N_353,In_1132,In_1240);
xnor U354 (N_354,In_1853,In_168);
nor U355 (N_355,In_2450,In_1050);
nand U356 (N_356,In_1757,In_519);
nor U357 (N_357,In_823,In_30);
and U358 (N_358,In_1986,In_2378);
nand U359 (N_359,In_218,In_2216);
or U360 (N_360,In_759,In_934);
xnor U361 (N_361,In_690,In_1179);
nand U362 (N_362,In_1159,In_81);
nor U363 (N_363,In_1194,In_329);
nor U364 (N_364,In_2134,In_1574);
nand U365 (N_365,In_1505,In_108);
nand U366 (N_366,In_147,In_2497);
nor U367 (N_367,In_1924,In_1843);
nor U368 (N_368,In_1754,In_873);
and U369 (N_369,In_900,In_2305);
nand U370 (N_370,In_1828,In_2070);
nand U371 (N_371,In_553,In_2424);
nand U372 (N_372,In_1716,In_398);
or U373 (N_373,In_19,In_1499);
and U374 (N_374,In_732,In_1569);
nor U375 (N_375,In_1237,In_581);
and U376 (N_376,In_854,In_2243);
nor U377 (N_377,In_1097,In_988);
or U378 (N_378,In_2245,In_2176);
nor U379 (N_379,In_764,In_928);
nand U380 (N_380,In_385,In_409);
and U381 (N_381,In_1124,In_2225);
and U382 (N_382,In_1688,In_2438);
or U383 (N_383,In_528,In_455);
and U384 (N_384,In_775,In_16);
and U385 (N_385,In_2013,In_1279);
nor U386 (N_386,In_2136,In_2442);
nand U387 (N_387,In_56,In_938);
and U388 (N_388,In_1978,In_590);
nor U389 (N_389,In_1804,In_2054);
or U390 (N_390,In_1624,In_801);
xnor U391 (N_391,In_1518,In_1238);
xnor U392 (N_392,In_2339,In_283);
and U393 (N_393,In_2124,In_157);
nor U394 (N_394,In_1379,In_1437);
or U395 (N_395,In_384,In_84);
nor U396 (N_396,In_2011,In_1896);
nor U397 (N_397,In_1936,In_1662);
nor U398 (N_398,In_513,In_1221);
nor U399 (N_399,In_727,In_244);
xor U400 (N_400,In_1940,In_743);
nor U401 (N_401,In_1808,In_109);
and U402 (N_402,In_1362,In_2432);
nor U403 (N_403,In_1141,In_2076);
or U404 (N_404,In_2303,In_720);
nand U405 (N_405,In_567,In_738);
and U406 (N_406,In_1162,In_1263);
and U407 (N_407,In_1337,In_153);
nor U408 (N_408,In_1123,In_1585);
nand U409 (N_409,In_66,In_1550);
xnor U410 (N_410,In_104,In_165);
and U411 (N_411,In_2271,In_2152);
xor U412 (N_412,In_2302,In_964);
and U413 (N_413,In_122,In_2440);
xnor U414 (N_414,In_148,In_824);
nor U415 (N_415,In_129,In_63);
and U416 (N_416,In_2038,In_1942);
nor U417 (N_417,In_401,In_1432);
nor U418 (N_418,In_1954,In_2040);
and U419 (N_419,In_2449,In_451);
and U420 (N_420,In_2273,In_320);
and U421 (N_421,In_296,In_97);
or U422 (N_422,In_924,In_769);
and U423 (N_423,In_1528,In_1272);
nor U424 (N_424,In_137,In_28);
xor U425 (N_425,In_1586,In_1786);
xor U426 (N_426,In_1981,In_2259);
xnor U427 (N_427,In_2283,In_2029);
or U428 (N_428,In_1268,In_318);
and U429 (N_429,In_1995,In_1383);
xnor U430 (N_430,In_751,In_929);
nand U431 (N_431,In_2014,In_1944);
xor U432 (N_432,In_1152,In_1395);
or U433 (N_433,In_243,In_630);
nand U434 (N_434,In_2377,In_2280);
nor U435 (N_435,In_1937,In_1131);
or U436 (N_436,In_1898,In_1627);
nor U437 (N_437,In_589,In_1534);
nor U438 (N_438,In_895,In_1359);
nor U439 (N_439,In_1513,In_492);
nand U440 (N_440,In_423,In_1614);
nand U441 (N_441,In_1660,In_1822);
or U442 (N_442,In_878,In_396);
nor U443 (N_443,In_2281,In_370);
xnor U444 (N_444,In_883,In_1389);
xnor U445 (N_445,In_1870,In_436);
and U446 (N_446,In_73,In_2116);
and U447 (N_447,In_1356,In_735);
nand U448 (N_448,In_784,In_1364);
and U449 (N_449,In_315,In_677);
and U450 (N_450,In_2472,In_2039);
nor U451 (N_451,In_1114,In_2331);
and U452 (N_452,In_1501,In_1382);
nand U453 (N_453,In_1210,In_1412);
xnor U454 (N_454,In_2431,In_1678);
nor U455 (N_455,In_1733,In_321);
nand U456 (N_456,In_1798,In_229);
nand U457 (N_457,In_1230,In_2175);
nor U458 (N_458,In_694,In_1173);
nand U459 (N_459,In_2228,In_989);
xnor U460 (N_460,In_1424,In_968);
and U461 (N_461,In_1388,In_1052);
and U462 (N_462,In_1801,In_876);
nor U463 (N_463,In_979,In_1167);
and U464 (N_464,In_241,In_974);
xnor U465 (N_465,In_1229,In_1790);
or U466 (N_466,In_539,In_1974);
or U467 (N_467,In_1126,In_1879);
nor U468 (N_468,In_88,In_2379);
xor U469 (N_469,In_1728,In_604);
or U470 (N_470,In_1169,In_2464);
or U471 (N_471,In_2435,In_789);
and U472 (N_472,In_834,In_2494);
nor U473 (N_473,In_1854,In_2055);
nand U474 (N_474,In_2052,In_183);
or U475 (N_475,In_594,In_901);
nor U476 (N_476,In_1351,In_837);
or U477 (N_477,In_1915,In_952);
or U478 (N_478,In_1935,In_2434);
xor U479 (N_479,In_359,In_1335);
nand U480 (N_480,In_577,In_523);
nor U481 (N_481,In_2436,In_1443);
and U482 (N_482,In_670,In_2081);
or U483 (N_483,In_86,In_2329);
nand U484 (N_484,In_1679,In_2269);
xnor U485 (N_485,In_1579,In_2193);
nand U486 (N_486,In_1306,In_2277);
nand U487 (N_487,In_2420,In_164);
or U488 (N_488,In_1993,In_607);
xor U489 (N_489,In_816,In_335);
nand U490 (N_490,In_2202,In_143);
nand U491 (N_491,In_419,In_2368);
nor U492 (N_492,In_800,In_309);
and U493 (N_493,In_715,In_606);
and U494 (N_494,In_1789,In_712);
nand U495 (N_495,In_2353,In_1649);
nor U496 (N_496,In_1764,In_485);
or U497 (N_497,In_286,In_193);
and U498 (N_498,In_77,In_349);
or U499 (N_499,In_2469,In_317);
and U500 (N_500,In_1557,In_69);
nor U501 (N_501,In_637,In_1845);
nand U502 (N_502,In_249,In_696);
nand U503 (N_503,In_2301,In_1948);
xor U504 (N_504,In_1185,In_1436);
nor U505 (N_505,In_48,In_1526);
nand U506 (N_506,In_114,In_1451);
nand U507 (N_507,In_470,In_1642);
nand U508 (N_508,In_1560,In_259);
nor U509 (N_509,In_1655,In_754);
nor U510 (N_510,In_1008,In_1552);
and U511 (N_511,In_1705,In_688);
and U512 (N_512,In_2356,In_176);
nand U513 (N_513,In_2135,In_1340);
or U514 (N_514,In_2490,In_2092);
or U515 (N_515,In_112,In_303);
and U516 (N_516,In_407,In_1369);
or U517 (N_517,In_1426,In_583);
xnor U518 (N_518,In_1400,In_1487);
nor U519 (N_519,In_1399,In_2147);
or U520 (N_520,In_1895,In_1347);
and U521 (N_521,In_1469,In_2115);
xnor U522 (N_522,In_67,In_559);
and U523 (N_523,In_1998,In_2100);
or U524 (N_524,In_1633,In_1640);
nand U525 (N_525,In_1905,In_1203);
xnor U526 (N_526,In_1164,In_38);
nor U527 (N_527,In_1015,In_2201);
nor U528 (N_528,In_1160,In_271);
nand U529 (N_529,In_771,In_561);
nand U530 (N_530,In_2218,In_574);
and U531 (N_531,In_2276,In_1323);
nand U532 (N_532,In_2355,In_227);
xnor U533 (N_533,In_1797,In_2477);
and U534 (N_534,In_864,In_1127);
xor U535 (N_535,In_613,In_36);
and U536 (N_536,In_1125,In_1013);
nor U537 (N_537,In_221,In_783);
nand U538 (N_538,In_341,In_2159);
nor U539 (N_539,In_196,In_650);
and U540 (N_540,In_872,In_270);
nand U541 (N_541,In_273,In_563);
xnor U542 (N_542,In_182,In_1666);
nand U543 (N_543,In_2132,In_1689);
and U544 (N_544,In_1338,In_2171);
xnor U545 (N_545,In_2213,In_1111);
nor U546 (N_546,In_2250,In_1817);
xnor U547 (N_547,In_744,In_443);
xor U548 (N_548,In_786,In_2466);
nor U549 (N_549,In_92,In_456);
and U550 (N_550,In_1824,In_1357);
nor U551 (N_551,In_1249,In_459);
xnor U552 (N_552,In_2064,In_1402);
xor U553 (N_553,In_2233,In_1597);
or U554 (N_554,In_2371,In_2190);
or U555 (N_555,In_832,In_785);
nor U556 (N_556,In_1952,In_61);
nand U557 (N_557,In_471,In_2232);
and U558 (N_558,In_687,In_742);
nor U559 (N_559,In_2309,In_1161);
and U560 (N_560,In_863,In_1694);
or U561 (N_561,In_1246,In_1257);
nor U562 (N_562,In_1561,In_829);
and U563 (N_563,In_1833,In_1729);
or U564 (N_564,In_2126,In_2097);
or U565 (N_565,In_1819,In_2158);
and U566 (N_566,In_1507,In_1904);
and U567 (N_567,In_2131,In_1086);
and U568 (N_568,In_2021,In_700);
xnor U569 (N_569,In_24,In_1294);
nand U570 (N_570,In_1792,In_1771);
xor U571 (N_571,In_13,In_2319);
or U572 (N_572,In_1325,In_1321);
xor U573 (N_573,In_91,In_698);
or U574 (N_574,In_1088,In_608);
nor U575 (N_575,In_746,In_2395);
and U576 (N_576,In_276,In_568);
or U577 (N_577,In_1392,In_1497);
or U578 (N_578,In_226,In_247);
nor U579 (N_579,In_285,In_1510);
xor U580 (N_580,In_1939,In_861);
nand U581 (N_581,In_236,In_2150);
xor U582 (N_582,In_263,In_740);
and U583 (N_583,In_537,In_2164);
nor U584 (N_584,In_2170,In_301);
nor U585 (N_585,In_417,In_1630);
or U586 (N_586,In_212,In_2087);
or U587 (N_587,In_1628,In_1028);
nor U588 (N_588,In_58,In_507);
and U589 (N_589,In_344,In_2468);
or U590 (N_590,In_452,In_1133);
and U591 (N_591,In_502,In_2453);
xor U592 (N_592,In_797,In_1245);
nor U593 (N_593,In_936,In_770);
and U594 (N_594,In_953,In_2247);
or U595 (N_595,In_1003,In_219);
nor U596 (N_596,In_1531,In_1504);
nand U597 (N_597,In_434,In_693);
nand U598 (N_598,In_264,In_1450);
or U599 (N_599,In_1057,In_2460);
or U600 (N_600,In_220,In_1699);
and U601 (N_601,In_997,In_1949);
and U602 (N_602,In_933,In_1581);
or U603 (N_603,In_994,In_1590);
and U604 (N_604,In_51,In_347);
xnor U605 (N_605,In_441,In_885);
or U606 (N_606,In_1025,In_2084);
nand U607 (N_607,In_2386,In_1675);
and U608 (N_608,In_2360,In_1867);
xor U609 (N_609,In_1975,In_643);
and U610 (N_610,In_1372,In_1017);
nand U611 (N_611,In_1156,In_382);
and U612 (N_612,In_2383,In_497);
and U613 (N_613,In_1001,In_961);
nand U614 (N_614,In_1157,In_116);
and U615 (N_615,In_2023,In_501);
or U616 (N_616,In_2324,In_2244);
and U617 (N_617,In_121,In_1917);
nand U618 (N_618,In_1568,In_26);
or U619 (N_619,In_1599,In_1850);
nor U620 (N_620,In_1405,In_1763);
and U621 (N_621,In_1816,In_1903);
or U622 (N_622,In_1760,In_660);
xor U623 (N_623,In_1051,In_1349);
or U624 (N_624,In_1639,In_1138);
and U625 (N_625,In_336,In_1592);
nand U626 (N_626,In_1957,In_141);
and U627 (N_627,In_1921,In_805);
nand U628 (N_628,In_1308,In_1712);
nor U629 (N_629,In_1459,In_1049);
nor U630 (N_630,In_2080,In_981);
and U631 (N_631,In_965,In_1130);
and U632 (N_632,In_674,In_1884);
nor U633 (N_633,In_191,In_159);
or U634 (N_634,In_2145,In_1023);
or U635 (N_635,In_198,In_1669);
nor U636 (N_636,In_1063,In_1869);
xor U637 (N_637,In_1394,In_2183);
nand U638 (N_638,In_1255,In_1785);
xnor U639 (N_639,In_2180,In_339);
or U640 (N_640,In_627,In_1076);
and U641 (N_641,In_240,In_1094);
and U642 (N_642,In_282,In_1769);
xnor U643 (N_643,In_7,In_614);
nand U644 (N_644,In_1621,In_2367);
and U645 (N_645,In_1799,In_1814);
xor U646 (N_646,In_2349,In_655);
xnor U647 (N_647,In_2496,In_1070);
and U648 (N_648,In_2144,In_246);
nor U649 (N_649,In_937,In_821);
and U650 (N_650,In_358,In_2165);
or U651 (N_651,In_1384,In_1914);
xnor U652 (N_652,In_290,In_1342);
nor U653 (N_653,In_1536,In_1953);
and U654 (N_654,In_1036,In_281);
nor U655 (N_655,In_1288,In_487);
nor U656 (N_656,In_2391,In_1406);
and U657 (N_657,In_2114,In_2380);
or U658 (N_658,In_1242,In_1613);
xor U659 (N_659,In_1887,In_1858);
xor U660 (N_660,In_1571,In_2335);
nor U661 (N_661,In_2293,In_1150);
and U662 (N_662,In_1992,In_503);
xor U663 (N_663,In_776,In_634);
nand U664 (N_664,In_1021,In_59);
nor U665 (N_665,In_996,In_120);
and U666 (N_666,In_2061,In_1906);
xor U667 (N_667,In_1573,In_52);
or U668 (N_668,In_2140,In_128);
xnor U669 (N_669,In_266,In_1885);
or U670 (N_670,In_1300,In_427);
nor U671 (N_671,In_328,In_2031);
nor U672 (N_672,In_237,In_1205);
or U673 (N_673,In_631,In_27);
nor U674 (N_674,In_1461,In_667);
and U675 (N_675,In_2082,In_1368);
or U676 (N_676,In_2163,In_2037);
and U677 (N_677,In_2208,In_855);
or U678 (N_678,In_962,In_1269);
and U679 (N_679,In_2314,In_1172);
or U680 (N_680,In_139,In_1136);
xor U681 (N_681,In_2034,In_1502);
nand U682 (N_682,In_648,In_736);
nand U683 (N_683,In_919,In_1653);
or U684 (N_684,In_334,In_429);
nor U685 (N_685,In_2060,In_1206);
or U686 (N_686,In_1775,In_709);
nand U687 (N_687,In_2458,In_1147);
nor U688 (N_688,In_2010,In_820);
nor U689 (N_689,In_1396,In_1187);
and U690 (N_690,In_1696,In_304);
nand U691 (N_691,In_757,In_1880);
nor U692 (N_692,In_12,In_300);
nand U693 (N_693,In_1192,In_1207);
and U694 (N_694,In_1324,In_2196);
nand U695 (N_695,In_189,In_871);
nor U696 (N_696,In_14,In_1472);
nand U697 (N_697,In_1163,In_848);
xor U698 (N_698,In_931,In_2212);
nor U699 (N_699,In_2361,In_976);
and U700 (N_700,In_2499,In_1096);
nor U701 (N_701,In_472,In_2121);
nand U702 (N_702,In_1455,In_473);
nor U703 (N_703,In_2257,In_214);
and U704 (N_704,In_2020,In_1109);
xnor U705 (N_705,In_2308,In_1343);
nand U706 (N_706,In_795,In_1958);
and U707 (N_707,In_2316,In_486);
and U708 (N_708,In_1332,In_378);
xnor U709 (N_709,In_1493,In_810);
nor U710 (N_710,In_494,In_1964);
xnor U711 (N_711,In_43,In_975);
nor U712 (N_712,In_1556,In_1471);
nor U713 (N_713,In_1374,In_465);
or U714 (N_714,In_1498,In_806);
or U715 (N_715,In_756,In_1059);
or U716 (N_716,In_402,In_1281);
nor U717 (N_717,In_2105,In_83);
and U718 (N_718,In_548,In_1752);
and U719 (N_719,In_1739,In_905);
xnor U720 (N_720,In_1521,In_21);
and U721 (N_721,In_2300,In_2000);
nand U722 (N_722,In_2198,In_706);
and U723 (N_723,In_1695,In_2239);
xnor U724 (N_724,In_1591,In_1648);
or U725 (N_725,In_530,In_1731);
and U726 (N_726,In_779,In_2123);
nor U727 (N_727,In_1946,In_2311);
nand U728 (N_728,In_652,In_1208);
xor U729 (N_729,In_1899,In_493);
and U730 (N_730,In_1408,In_2024);
or U731 (N_731,In_1683,In_32);
and U732 (N_732,In_514,In_499);
or U733 (N_733,In_1734,In_1113);
nand U734 (N_734,In_1068,In_1468);
xnor U735 (N_735,In_163,In_1065);
nand U736 (N_736,In_430,In_254);
xor U737 (N_737,In_788,In_1962);
nand U738 (N_738,In_479,In_435);
xnor U739 (N_739,In_1259,In_490);
and U740 (N_740,In_260,In_825);
nor U741 (N_741,In_758,In_772);
xor U742 (N_742,In_2033,In_2492);
or U743 (N_743,In_2035,In_365);
or U744 (N_744,In_2088,In_1310);
xnor U745 (N_745,In_618,In_2437);
and U746 (N_746,In_1305,In_475);
nand U747 (N_747,In_217,In_1533);
xor U748 (N_748,In_175,In_1582);
nand U749 (N_749,In_1744,In_666);
or U750 (N_750,In_1239,In_827);
xnor U751 (N_751,In_831,In_1927);
xnor U752 (N_752,In_2321,In_2288);
and U753 (N_753,In_1693,In_1346);
nand U754 (N_754,In_1929,In_2069);
and U755 (N_755,In_2,In_277);
nand U756 (N_756,In_331,In_184);
nand U757 (N_757,In_945,In_2248);
nor U758 (N_758,In_1232,In_1303);
and U759 (N_759,In_1085,In_322);
xor U760 (N_760,In_658,In_1580);
nor U761 (N_761,In_544,In_956);
nand U762 (N_762,In_2483,In_1319);
xor U763 (N_763,In_146,In_2096);
xor U764 (N_764,In_1800,In_268);
or U765 (N_765,In_284,In_2099);
and U766 (N_766,In_1280,In_1100);
nor U767 (N_767,In_815,In_819);
nand U768 (N_768,In_1584,In_1448);
xor U769 (N_769,In_1522,In_2166);
nor U770 (N_770,In_731,In_1738);
and U771 (N_771,In_1216,In_1966);
xor U772 (N_772,In_512,In_1000);
xnor U773 (N_773,In_1494,In_1030);
xor U774 (N_774,In_1248,In_1298);
nand U775 (N_775,In_1664,In_1698);
or U776 (N_776,In_397,In_1930);
and U777 (N_777,In_1439,In_140);
nand U778 (N_778,In_65,In_2186);
or U779 (N_779,In_1119,In_555);
nor U780 (N_780,In_1857,In_1941);
and U781 (N_781,In_2133,In_1864);
nand U782 (N_782,In_603,In_1918);
nor U783 (N_783,In_1144,In_932);
nor U784 (N_784,In_1429,In_628);
or U785 (N_785,In_565,In_399);
and U786 (N_786,In_640,In_1261);
nor U787 (N_787,In_2068,In_1564);
xnor U788 (N_788,In_1661,In_2441);
or U789 (N_789,In_2146,In_817);
and U790 (N_790,In_1423,In_1572);
and U791 (N_791,In_616,In_1219);
xor U792 (N_792,In_1029,In_915);
and U793 (N_793,In_177,In_2047);
nor U794 (N_794,In_1353,In_1350);
or U795 (N_795,In_280,In_167);
or U796 (N_796,In_2462,In_943);
nand U797 (N_797,In_2401,In_1866);
or U798 (N_798,In_2396,In_605);
nor U799 (N_799,In_1077,In_636);
nor U800 (N_800,In_1020,In_1481);
xor U801 (N_801,In_760,In_138);
or U802 (N_802,In_462,In_224);
or U803 (N_803,In_289,In_2138);
nand U804 (N_804,In_856,In_1390);
or U805 (N_805,In_930,In_1002);
nand U806 (N_806,In_1007,In_323);
or U807 (N_807,In_478,In_1616);
and U808 (N_808,In_2350,In_870);
and U809 (N_809,In_1697,In_1641);
or U810 (N_810,In_906,In_1195);
nand U811 (N_811,In_1503,In_72);
nand U812 (N_812,In_1380,In_1901);
and U813 (N_813,In_1637,In_1139);
or U814 (N_814,In_1721,In_319);
and U815 (N_815,In_1525,In_2385);
xnor U816 (N_816,In_1787,In_2476);
xnor U817 (N_817,In_911,In_1741);
nor U818 (N_818,In_2234,In_626);
nand U819 (N_819,In_1355,In_673);
nor U820 (N_820,In_1663,In_35);
xor U821 (N_821,In_535,In_400);
and U822 (N_822,In_593,In_469);
nor U823 (N_823,In_946,In_235);
nand U824 (N_824,In_2374,In_1747);
nand U825 (N_825,In_1625,In_671);
xnor U826 (N_826,In_2357,In_354);
and U827 (N_827,In_1611,In_2295);
or U828 (N_828,In_1365,In_1490);
nand U829 (N_829,In_597,In_2348);
nand U830 (N_830,In_2398,In_6);
and U831 (N_831,In_753,In_2451);
or U832 (N_832,In_2249,In_844);
nor U833 (N_833,In_1033,In_0);
nor U834 (N_834,In_1289,In_2381);
nor U835 (N_835,In_719,In_1809);
nand U836 (N_836,In_1856,In_1907);
and U837 (N_837,In_853,In_1969);
nor U838 (N_838,In_2262,In_265);
xor U839 (N_839,In_2155,In_898);
or U840 (N_840,In_689,In_1976);
nand U841 (N_841,In_2409,In_1806);
and U842 (N_842,In_110,In_2235);
nor U843 (N_843,In_1006,In_239);
nor U844 (N_844,In_1562,In_2322);
nor U845 (N_845,In_2495,In_750);
and U846 (N_846,In_2320,In_395);
or U847 (N_847,In_542,In_1256);
or U848 (N_848,In_457,In_1897);
nand U849 (N_849,In_1004,In_278);
nor U850 (N_850,In_1375,In_1460);
or U851 (N_851,In_1881,In_2045);
or U852 (N_852,In_653,In_840);
or U853 (N_853,In_558,In_415);
and U854 (N_854,In_2128,In_1012);
and U855 (N_855,In_1530,In_1919);
nor U856 (N_856,In_792,In_98);
or U857 (N_857,In_1201,In_1378);
xnor U858 (N_858,In_204,In_1770);
xor U859 (N_859,In_504,In_1102);
nand U860 (N_860,In_1098,In_1506);
and U861 (N_861,In_2154,In_1473);
and U862 (N_862,In_149,In_992);
and U863 (N_863,In_1718,In_1691);
nand U864 (N_864,In_53,In_2160);
or U865 (N_865,In_1329,In_1554);
xnor U866 (N_866,In_1121,In_896);
and U867 (N_867,In_940,In_461);
and U868 (N_868,In_345,In_1783);
nor U869 (N_869,In_75,In_2006);
xor U870 (N_870,In_2199,In_835);
nor U871 (N_871,In_1107,In_2392);
or U872 (N_872,In_2167,In_2478);
xnor U873 (N_873,In_1827,In_886);
nand U874 (N_874,In_654,In_2465);
nor U875 (N_875,In_1056,In_984);
xor U876 (N_876,In_1260,In_1532);
xor U877 (N_877,In_1835,In_1165);
nand U878 (N_878,In_446,In_348);
and U879 (N_879,In_724,In_10);
or U880 (N_880,In_1456,In_526);
nand U881 (N_881,In_699,In_1043);
and U882 (N_882,In_89,In_1103);
nand U883 (N_883,In_570,In_922);
and U884 (N_884,In_1979,In_869);
and U885 (N_885,In_1709,In_371);
or U886 (N_886,In_1116,In_868);
xor U887 (N_887,In_1209,In_169);
nor U888 (N_888,In_252,In_245);
and U889 (N_889,In_1737,In_1462);
nand U890 (N_890,In_192,In_691);
nand U891 (N_891,In_1861,In_1222);
or U892 (N_892,In_1925,In_1659);
xnor U893 (N_893,In_560,In_133);
nor U894 (N_894,In_1587,In_1128);
nand U895 (N_895,In_1959,In_2195);
xnor U896 (N_896,In_248,In_2284);
and U897 (N_897,In_2285,In_388);
xnor U898 (N_898,In_1060,In_2275);
and U899 (N_899,In_550,In_1514);
and U900 (N_900,In_1748,In_2278);
xor U901 (N_901,In_2108,In_612);
or U902 (N_902,In_1762,In_1511);
nand U903 (N_903,In_102,In_2191);
and U904 (N_904,In_828,In_70);
and U905 (N_905,In_2291,In_601);
xnor U906 (N_906,In_437,In_1027);
nand U907 (N_907,In_46,In_1074);
xnor U908 (N_908,In_1284,In_2251);
or U909 (N_909,In_1477,In_1595);
or U910 (N_910,In_813,In_798);
and U911 (N_911,In_172,In_2413);
nand U912 (N_912,In_96,In_2366);
and U913 (N_913,In_2266,In_1197);
and U914 (N_914,In_1155,In_2263);
and U915 (N_915,In_2149,In_44);
nand U916 (N_916,In_161,In_2148);
xnor U917 (N_917,In_1295,In_1447);
nor U918 (N_918,In_957,In_897);
and U919 (N_919,In_460,In_1991);
nand U920 (N_920,In_1715,In_1753);
xor U921 (N_921,In_990,In_311);
nand U922 (N_922,In_1776,In_2051);
or U923 (N_923,In_1196,In_2122);
nor U924 (N_924,In_2403,In_2443);
nor U925 (N_925,In_860,In_33);
or U926 (N_926,In_2200,In_2459);
xor U927 (N_927,In_669,In_685);
and U928 (N_928,In_1352,In_1932);
nor U929 (N_929,In_448,In_1453);
xnor U930 (N_930,In_1961,In_2461);
and U931 (N_931,In_342,In_572);
and U932 (N_932,In_1547,In_879);
and U933 (N_933,In_2057,In_1676);
nor U934 (N_934,In_1431,In_411);
and U935 (N_935,In_1973,In_2390);
and U936 (N_936,In_439,In_600);
nor U937 (N_937,In_2267,In_1652);
nor U938 (N_938,In_333,In_316);
or U939 (N_939,In_1710,In_908);
xnor U940 (N_940,In_2292,In_1566);
and U941 (N_941,In_847,In_2294);
nor U942 (N_942,In_343,In_2041);
nor U943 (N_943,In_1782,In_477);
nor U944 (N_944,In_849,In_2102);
nand U945 (N_945,In_880,In_369);
nor U946 (N_946,In_2342,In_1686);
nor U947 (N_947,In_1140,In_1427);
nor U948 (N_948,In_216,In_294);
nand U949 (N_949,In_737,In_466);
or U950 (N_950,In_2091,In_2344);
or U951 (N_951,In_1067,In_1250);
or U952 (N_952,In_633,In_2210);
or U953 (N_953,In_2307,In_1454);
and U954 (N_954,In_1428,In_2373);
or U955 (N_955,In_2414,In_255);
nand U956 (N_956,In_1687,In_1270);
and U957 (N_957,In_426,In_1610);
and U958 (N_958,In_533,In_1726);
nand U959 (N_959,In_1761,In_352);
and U960 (N_960,In_1293,In_1796);
nor U961 (N_961,In_454,In_850);
xnor U962 (N_962,In_960,In_999);
nand U963 (N_963,In_1667,In_23);
xnor U964 (N_964,In_2153,In_1112);
or U965 (N_965,In_1344,In_1170);
xnor U966 (N_966,In_211,In_111);
nor U967 (N_967,In_134,In_695);
nor U968 (N_968,In_1366,In_2388);
xnor U969 (N_969,In_403,In_47);
nor U970 (N_970,In_39,In_1055);
nor U971 (N_971,In_291,In_368);
and U972 (N_972,In_308,In_2246);
nor U973 (N_973,In_571,In_646);
and U974 (N_974,In_1657,In_1080);
xnor U975 (N_975,In_34,In_1951);
nand U976 (N_976,In_1608,In_1118);
or U977 (N_977,In_1523,In_424);
xor U978 (N_978,In_267,In_1011);
xnor U979 (N_979,In_1645,In_1820);
nand U980 (N_980,In_2056,In_733);
and U981 (N_981,In_207,In_1723);
nand U982 (N_982,In_2127,In_364);
nor U983 (N_983,In_713,In_2067);
or U984 (N_984,In_2109,In_1292);
or U985 (N_985,In_2264,In_2454);
xor U986 (N_986,In_366,In_1618);
xor U987 (N_987,In_391,In_1647);
nor U988 (N_988,In_1463,In_130);
nor U989 (N_989,In_1488,In_812);
xnor U990 (N_990,In_1489,In_617);
xnor U991 (N_991,In_68,In_1252);
nor U992 (N_992,In_2078,In_1483);
nand U993 (N_993,In_1677,In_2027);
or U994 (N_994,In_126,In_2255);
xnor U995 (N_995,In_1258,In_705);
and U996 (N_996,In_1989,In_2402);
or U997 (N_997,In_1492,In_2423);
nand U998 (N_998,In_1234,In_1215);
or U999 (N_999,In_1053,In_2328);
nand U1000 (N_1000,In_947,In_780);
nor U1001 (N_1001,In_2215,In_353);
nor U1002 (N_1002,In_1330,In_2493);
and U1003 (N_1003,In_1104,In_904);
nor U1004 (N_1004,In_1381,In_2417);
nand U1005 (N_1005,In_767,In_2286);
xnor U1006 (N_1006,In_755,In_778);
and U1007 (N_1007,In_675,In_1539);
nor U1008 (N_1008,In_1241,In_2107);
and U1009 (N_1009,In_1778,In_496);
and U1010 (N_1010,In_1307,In_1545);
nor U1011 (N_1011,In_1122,In_2261);
xnor U1012 (N_1012,In_1743,In_1223);
or U1013 (N_1013,In_1889,In_313);
and U1014 (N_1014,In_1713,In_1283);
or U1015 (N_1015,In_386,In_1793);
nand U1016 (N_1016,In_152,In_166);
nand U1017 (N_1017,In_1311,In_1415);
and U1018 (N_1018,In_1046,In_1658);
nand U1019 (N_1019,In_194,In_355);
and U1020 (N_1020,In_1485,In_1397);
nand U1021 (N_1021,In_2299,In_649);
nand U1022 (N_1022,In_734,In_2079);
xor U1023 (N_1023,In_2351,In_37);
and U1024 (N_1024,In_393,In_1265);
nand U1025 (N_1025,In_913,In_745);
xor U1026 (N_1026,In_1603,In_680);
or U1027 (N_1027,In_1034,In_2456);
and U1028 (N_1028,In_510,In_1999);
or U1029 (N_1029,In_41,In_1134);
nor U1030 (N_1030,In_1274,In_222);
nor U1031 (N_1031,In_566,In_489);
nor U1032 (N_1032,In_1476,In_1464);
nor U1033 (N_1033,In_1166,In_495);
xor U1034 (N_1034,In_1943,In_1546);
nand U1035 (N_1035,In_793,In_1226);
or U1036 (N_1036,In_215,In_1549);
nor U1037 (N_1037,In_2073,In_506);
and U1038 (N_1038,In_520,In_2429);
xnor U1039 (N_1039,In_1048,In_562);
and U1040 (N_1040,In_1401,In_256);
or U1041 (N_1041,In_1452,In_1022);
xor U1042 (N_1042,In_298,In_90);
and U1043 (N_1043,In_641,In_2363);
or U1044 (N_1044,In_944,In_569);
xnor U1045 (N_1045,In_447,In_1934);
nand U1046 (N_1046,In_1370,In_708);
nor U1047 (N_1047,In_875,In_2046);
or U1048 (N_1048,In_338,In_4);
xnor U1049 (N_1049,In_579,In_609);
nand U1050 (N_1050,In_1193,In_1894);
nor U1051 (N_1051,In_1331,In_1794);
nand U1052 (N_1052,In_1273,In_2289);
nand U1053 (N_1053,In_1047,In_916);
nor U1054 (N_1054,In_1875,In_1965);
xor U1055 (N_1055,In_763,In_1871);
nor U1056 (N_1056,In_11,In_833);
or U1057 (N_1057,In_440,In_2211);
or U1058 (N_1058,In_1882,In_2484);
nand U1059 (N_1059,In_1559,In_1411);
nand U1060 (N_1060,In_1290,In_977);
nand U1061 (N_1061,In_1955,In_40);
nand U1062 (N_1062,In_676,In_970);
or U1063 (N_1063,In_389,In_1766);
or U1064 (N_1064,In_2352,In_1072);
nand U1065 (N_1065,In_1084,In_1198);
nand U1066 (N_1066,In_64,In_1278);
nand U1067 (N_1067,In_1445,In_234);
and U1068 (N_1068,In_2058,In_1418);
and U1069 (N_1069,In_1398,In_2062);
or U1070 (N_1070,In_1039,In_1842);
xor U1071 (N_1071,In_1184,In_197);
nor U1072 (N_1072,In_1360,In_822);
xor U1073 (N_1073,In_726,In_1262);
nor U1074 (N_1074,In_725,In_275);
or U1075 (N_1075,In_2137,In_662);
nand U1076 (N_1076,In_2279,In_1117);
nand U1077 (N_1077,In_620,In_1087);
and U1078 (N_1078,In_2139,In_794);
nand U1079 (N_1079,In_299,In_2482);
nor U1080 (N_1080,In_602,In_127);
xnor U1081 (N_1081,In_200,In_357);
or U1082 (N_1082,In_2075,In_730);
and U1083 (N_1083,In_187,In_2359);
nand U1084 (N_1084,In_954,In_518);
xnor U1085 (N_1085,In_1607,In_2015);
xnor U1086 (N_1086,In_899,In_82);
nand U1087 (N_1087,In_1457,In_995);
xnor U1088 (N_1088,In_170,In_826);
nand U1089 (N_1089,In_809,In_1708);
xor U1090 (N_1090,In_20,In_2471);
and U1091 (N_1091,In_2182,In_611);
and U1092 (N_1092,In_1831,In_2400);
or U1093 (N_1093,In_25,In_1075);
or U1094 (N_1094,In_1893,In_2448);
xor U1095 (N_1095,In_1031,In_1543);
nand U1096 (N_1096,In_1529,In_242);
nand U1097 (N_1097,In_2358,In_1750);
nand U1098 (N_1098,In_99,In_433);
and U1099 (N_1099,In_1779,In_1367);
nand U1100 (N_1100,In_762,In_1983);
nand U1101 (N_1101,In_703,In_1467);
nor U1102 (N_1102,In_2065,In_78);
or U1103 (N_1103,In_678,In_2112);
or U1104 (N_1104,In_1444,In_173);
or U1105 (N_1105,In_2384,In_93);
or U1106 (N_1106,In_332,In_2455);
nor U1107 (N_1107,In_2002,In_463);
and U1108 (N_1108,In_2415,In_540);
xnor U1109 (N_1109,In_1495,In_1541);
and U1110 (N_1110,In_1832,In_1416);
nand U1111 (N_1111,In_297,In_305);
nor U1112 (N_1112,In_1631,In_1264);
or U1113 (N_1113,In_373,In_1650);
nor U1114 (N_1114,In_1061,In_1129);
and U1115 (N_1115,In_949,In_1643);
and U1116 (N_1116,In_942,In_2254);
nor U1117 (N_1117,In_2354,In_1742);
xnor U1118 (N_1118,In_2188,In_1182);
xor U1119 (N_1119,In_1247,In_2376);
and U1120 (N_1120,In_1839,In_1099);
xnor U1121 (N_1121,In_2467,In_325);
and U1122 (N_1122,In_1558,In_549);
xnor U1123 (N_1123,In_1376,In_2446);
and U1124 (N_1124,In_527,In_2296);
xor U1125 (N_1125,In_1354,In_155);
or U1126 (N_1126,In_1251,In_1153);
or U1127 (N_1127,In_920,In_2043);
nor U1128 (N_1128,In_2238,In_2197);
or U1129 (N_1129,In_839,In_1385);
xnor U1130 (N_1130,In_2214,In_1220);
xnor U1131 (N_1131,In_2425,In_1865);
nor U1132 (N_1132,In_287,In_573);
nand U1133 (N_1133,In_210,In_1996);
xnor U1134 (N_1134,In_657,In_2074);
and U1135 (N_1135,In_787,In_2406);
and U1136 (N_1136,In_1291,In_1474);
or U1137 (N_1137,In_619,In_293);
nand U1138 (N_1138,In_1217,In_2004);
xor U1139 (N_1139,In_1158,In_421);
or U1140 (N_1140,In_2419,In_1567);
nand U1141 (N_1141,In_2325,In_1190);
nand U1142 (N_1142,In_80,In_874);
nand U1143 (N_1143,In_1711,In_1093);
xor U1144 (N_1144,In_2030,In_387);
nor U1145 (N_1145,In_1095,In_2219);
xnor U1146 (N_1146,In_1706,In_1847);
nand U1147 (N_1147,In_2345,In_2486);
nand U1148 (N_1148,In_1042,In_1807);
nand U1149 (N_1149,In_1600,In_476);
or U1150 (N_1150,In_1740,In_1434);
xnor U1151 (N_1151,In_106,In_1304);
and U1152 (N_1152,In_843,In_925);
xor U1153 (N_1153,In_2488,In_1296);
xor U1154 (N_1154,In_1035,In_998);
xor U1155 (N_1155,In_2223,In_185);
and U1156 (N_1156,In_346,In_543);
xor U1157 (N_1157,In_1040,In_963);
nor U1158 (N_1158,In_2119,In_1886);
xnor U1159 (N_1159,In_392,In_909);
xnor U1160 (N_1160,In_1404,In_1670);
and U1161 (N_1161,In_432,In_894);
nand U1162 (N_1162,In_1202,In_95);
xnor U1163 (N_1163,In_2365,In_2125);
nor U1164 (N_1164,In_1883,In_1811);
and U1165 (N_1165,In_1334,In_1960);
or U1166 (N_1166,In_1542,In_94);
nand U1167 (N_1167,In_1736,In_233);
and U1168 (N_1168,In_1548,In_2318);
nor U1169 (N_1169,In_1277,In_635);
xnor U1170 (N_1170,In_1253,In_1482);
and U1171 (N_1171,In_596,In_1105);
or U1172 (N_1172,In_1218,In_375);
and U1173 (N_1173,In_274,In_521);
and U1174 (N_1174,In_1730,In_546);
or U1175 (N_1175,In_1180,In_672);
nand U1176 (N_1176,In_1538,In_1092);
nand U1177 (N_1177,In_1629,In_2336);
or U1178 (N_1178,In_1420,In_2142);
nand U1179 (N_1179,In_2480,In_2439);
or U1180 (N_1180,In_1873,In_2162);
or U1181 (N_1181,In_505,In_1777);
nand U1182 (N_1182,In_536,In_1315);
and U1183 (N_1183,In_2178,In_697);
xnor U1184 (N_1184,In_1231,In_1872);
nor U1185 (N_1185,In_951,In_1788);
and U1186 (N_1186,In_1286,In_1749);
xnor U1187 (N_1187,In_144,In_1509);
xnor U1188 (N_1188,In_1834,In_592);
nand U1189 (N_1189,In_481,In_1024);
xnor U1190 (N_1190,In_1120,In_1970);
or U1191 (N_1191,In_1,In_269);
and U1192 (N_1192,In_1413,In_716);
xor U1193 (N_1193,In_1910,In_54);
xnor U1194 (N_1194,In_584,In_858);
or U1195 (N_1195,In_105,In_2240);
xnor U1196 (N_1196,In_991,In_2172);
xnor U1197 (N_1197,In_1938,In_857);
and U1198 (N_1198,In_1784,In_1911);
nor U1199 (N_1199,In_1605,In_802);
and U1200 (N_1200,In_1211,In_532);
xnor U1201 (N_1201,In_2362,In_1891);
nor U1202 (N_1202,In_912,In_379);
nand U1203 (N_1203,In_306,In_1326);
nand U1204 (N_1204,In_2364,In_1361);
or U1205 (N_1205,In_2221,In_1005);
nor U1206 (N_1206,In_201,In_1458);
and U1207 (N_1207,In_625,In_302);
nand U1208 (N_1208,In_921,In_1619);
and U1209 (N_1209,In_422,In_2333);
xor U1210 (N_1210,In_803,In_882);
nor U1211 (N_1211,In_888,In_1312);
nor U1212 (N_1212,In_2007,In_480);
nor U1213 (N_1213,In_1110,In_1515);
nand U1214 (N_1214,In_1671,In_8);
nand U1215 (N_1215,In_1336,In_1909);
nand U1216 (N_1216,In_1945,In_923);
xor U1217 (N_1217,In_1684,In_556);
nand U1218 (N_1218,In_1496,In_414);
nor U1219 (N_1219,In_1916,In_1968);
and U1220 (N_1220,In_62,In_582);
xor U1221 (N_1221,In_1594,In_1967);
or U1222 (N_1222,In_2274,In_1425);
nand U1223 (N_1223,In_383,In_2310);
and U1224 (N_1224,In_534,In_2018);
nor U1225 (N_1225,In_525,In_1327);
xor U1226 (N_1226,In_971,In_1387);
and U1227 (N_1227,In_2332,In_2457);
nor U1228 (N_1228,In_531,In_2093);
nand U1229 (N_1229,In_517,In_629);
nand U1230 (N_1230,In_902,In_710);
or U1231 (N_1231,In_483,In_1846);
nand U1232 (N_1232,In_1544,In_1874);
nor U1233 (N_1233,In_1465,In_927);
and U1234 (N_1234,In_1137,In_1746);
xor U1235 (N_1235,In_891,In_292);
nor U1236 (N_1236,In_2479,In_2313);
nand U1237 (N_1237,In_1168,In_2306);
and U1238 (N_1238,In_2077,In_1177);
or U1239 (N_1239,In_208,In_174);
nand U1240 (N_1240,In_1038,In_1225);
nor U1241 (N_1241,In_939,In_1339);
or U1242 (N_1242,In_1236,In_917);
xor U1243 (N_1243,In_1475,In_361);
or U1244 (N_1244,In_2282,In_431);
nand U1245 (N_1245,In_231,In_2253);
nor U1246 (N_1246,In_1287,In_1555);
xor U1247 (N_1247,In_1466,In_1665);
and U1248 (N_1248,In_982,In_1078);
nor U1249 (N_1249,In_718,In_1438);
or U1250 (N_1250,N_852,N_1063);
and U1251 (N_1251,N_347,N_1178);
xnor U1252 (N_1252,N_568,N_906);
and U1253 (N_1253,N_813,N_773);
nor U1254 (N_1254,N_241,N_677);
nor U1255 (N_1255,N_1187,N_1098);
nand U1256 (N_1256,N_889,N_166);
or U1257 (N_1257,N_960,N_595);
xor U1258 (N_1258,N_1044,N_474);
nand U1259 (N_1259,N_1239,N_571);
nor U1260 (N_1260,N_698,N_788);
and U1261 (N_1261,N_145,N_214);
or U1262 (N_1262,N_1212,N_395);
or U1263 (N_1263,N_130,N_134);
and U1264 (N_1264,N_397,N_566);
or U1265 (N_1265,N_486,N_503);
nand U1266 (N_1266,N_579,N_932);
nand U1267 (N_1267,N_1154,N_10);
or U1268 (N_1268,N_538,N_246);
or U1269 (N_1269,N_228,N_509);
xnor U1270 (N_1270,N_1195,N_602);
nand U1271 (N_1271,N_201,N_820);
and U1272 (N_1272,N_1113,N_294);
nor U1273 (N_1273,N_296,N_449);
and U1274 (N_1274,N_531,N_167);
xnor U1275 (N_1275,N_54,N_812);
nand U1276 (N_1276,N_922,N_1086);
or U1277 (N_1277,N_1043,N_890);
nand U1278 (N_1278,N_415,N_32);
or U1279 (N_1279,N_55,N_625);
or U1280 (N_1280,N_489,N_340);
nor U1281 (N_1281,N_876,N_101);
nand U1282 (N_1282,N_950,N_945);
or U1283 (N_1283,N_394,N_760);
nor U1284 (N_1284,N_716,N_1220);
xnor U1285 (N_1285,N_1146,N_758);
xnor U1286 (N_1286,N_836,N_409);
nand U1287 (N_1287,N_517,N_493);
and U1288 (N_1288,N_541,N_671);
nor U1289 (N_1289,N_1228,N_837);
nand U1290 (N_1290,N_1186,N_182);
and U1291 (N_1291,N_1218,N_557);
and U1292 (N_1292,N_258,N_968);
nor U1293 (N_1293,N_679,N_887);
xor U1294 (N_1294,N_412,N_631);
and U1295 (N_1295,N_648,N_361);
nor U1296 (N_1296,N_882,N_614);
nand U1297 (N_1297,N_877,N_6);
nor U1298 (N_1298,N_610,N_389);
and U1299 (N_1299,N_63,N_642);
nand U1300 (N_1300,N_424,N_643);
and U1301 (N_1301,N_382,N_172);
or U1302 (N_1302,N_985,N_535);
or U1303 (N_1303,N_243,N_159);
nand U1304 (N_1304,N_947,N_104);
and U1305 (N_1305,N_661,N_405);
nor U1306 (N_1306,N_1104,N_457);
and U1307 (N_1307,N_280,N_478);
nand U1308 (N_1308,N_810,N_963);
nand U1309 (N_1309,N_658,N_384);
nand U1310 (N_1310,N_881,N_1151);
xor U1311 (N_1311,N_750,N_608);
nand U1312 (N_1312,N_358,N_128);
xor U1313 (N_1313,N_1047,N_1100);
nor U1314 (N_1314,N_419,N_1059);
nand U1315 (N_1315,N_1153,N_1079);
or U1316 (N_1316,N_630,N_1164);
xnor U1317 (N_1317,N_849,N_589);
and U1318 (N_1318,N_133,N_597);
xnor U1319 (N_1319,N_999,N_833);
nor U1320 (N_1320,N_1062,N_834);
and U1321 (N_1321,N_867,N_547);
nand U1322 (N_1322,N_187,N_312);
nor U1323 (N_1323,N_1070,N_365);
nor U1324 (N_1324,N_34,N_1089);
xor U1325 (N_1325,N_640,N_649);
and U1326 (N_1326,N_757,N_324);
or U1327 (N_1327,N_224,N_1201);
and U1328 (N_1328,N_878,N_22);
nand U1329 (N_1329,N_49,N_184);
xnor U1330 (N_1330,N_697,N_426);
nor U1331 (N_1331,N_728,N_1046);
nand U1332 (N_1332,N_992,N_800);
nor U1333 (N_1333,N_238,N_617);
or U1334 (N_1334,N_1168,N_983);
and U1335 (N_1335,N_994,N_103);
and U1336 (N_1336,N_868,N_1072);
and U1337 (N_1337,N_357,N_297);
or U1338 (N_1338,N_809,N_718);
or U1339 (N_1339,N_1191,N_1221);
nand U1340 (N_1340,N_600,N_1129);
xor U1341 (N_1341,N_270,N_711);
nand U1342 (N_1342,N_441,N_1045);
nand U1343 (N_1343,N_633,N_399);
nor U1344 (N_1344,N_157,N_1161);
or U1345 (N_1345,N_117,N_298);
nor U1346 (N_1346,N_1031,N_148);
or U1347 (N_1347,N_1011,N_693);
nor U1348 (N_1348,N_91,N_739);
and U1349 (N_1349,N_993,N_545);
or U1350 (N_1350,N_220,N_713);
or U1351 (N_1351,N_856,N_843);
xnor U1352 (N_1352,N_1145,N_1193);
xor U1353 (N_1353,N_916,N_68);
xnor U1354 (N_1354,N_37,N_1049);
or U1355 (N_1355,N_522,N_937);
and U1356 (N_1356,N_460,N_721);
or U1357 (N_1357,N_929,N_607);
nand U1358 (N_1358,N_252,N_1209);
xor U1359 (N_1359,N_82,N_338);
and U1360 (N_1360,N_376,N_17);
nand U1361 (N_1361,N_569,N_348);
xnor U1362 (N_1362,N_1057,N_90);
and U1363 (N_1363,N_266,N_300);
xor U1364 (N_1364,N_984,N_612);
and U1365 (N_1365,N_761,N_110);
nand U1366 (N_1366,N_178,N_121);
nor U1367 (N_1367,N_248,N_436);
nand U1368 (N_1368,N_275,N_664);
nor U1369 (N_1369,N_722,N_1242);
nor U1370 (N_1370,N_359,N_1019);
and U1371 (N_1371,N_1035,N_907);
nand U1372 (N_1372,N_111,N_830);
and U1373 (N_1373,N_400,N_210);
and U1374 (N_1374,N_554,N_255);
and U1375 (N_1375,N_705,N_1233);
and U1376 (N_1376,N_520,N_1182);
nand U1377 (N_1377,N_969,N_583);
nand U1378 (N_1378,N_289,N_663);
nand U1379 (N_1379,N_1159,N_373);
or U1380 (N_1380,N_565,N_826);
or U1381 (N_1381,N_1094,N_885);
nand U1382 (N_1382,N_1054,N_479);
xor U1383 (N_1383,N_1244,N_841);
nand U1384 (N_1384,N_1010,N_870);
xor U1385 (N_1385,N_1222,N_370);
xnor U1386 (N_1386,N_539,N_949);
or U1387 (N_1387,N_644,N_551);
xor U1388 (N_1388,N_212,N_896);
xor U1389 (N_1389,N_206,N_952);
nor U1390 (N_1390,N_72,N_817);
nor U1391 (N_1391,N_585,N_979);
xor U1392 (N_1392,N_913,N_463);
nor U1393 (N_1393,N_18,N_793);
nand U1394 (N_1394,N_112,N_927);
and U1395 (N_1395,N_601,N_763);
or U1396 (N_1396,N_1002,N_292);
and U1397 (N_1397,N_28,N_410);
or U1398 (N_1398,N_550,N_1150);
nand U1399 (N_1399,N_578,N_323);
nand U1400 (N_1400,N_732,N_407);
nand U1401 (N_1401,N_895,N_518);
nand U1402 (N_1402,N_47,N_1246);
and U1403 (N_1403,N_288,N_1160);
nand U1404 (N_1404,N_1188,N_253);
nor U1405 (N_1405,N_1083,N_1119);
nor U1406 (N_1406,N_1249,N_835);
xnor U1407 (N_1407,N_781,N_329);
nand U1408 (N_1408,N_366,N_1040);
nand U1409 (N_1409,N_1141,N_417);
or U1410 (N_1410,N_94,N_1005);
and U1411 (N_1411,N_745,N_1200);
nor U1412 (N_1412,N_590,N_102);
or U1413 (N_1413,N_847,N_445);
or U1414 (N_1414,N_1015,N_832);
nor U1415 (N_1415,N_943,N_219);
and U1416 (N_1416,N_84,N_873);
nor U1417 (N_1417,N_1226,N_230);
or U1418 (N_1418,N_942,N_654);
and U1419 (N_1419,N_767,N_851);
nor U1420 (N_1420,N_466,N_706);
xnor U1421 (N_1421,N_914,N_899);
xnor U1422 (N_1422,N_66,N_435);
or U1423 (N_1423,N_337,N_468);
xor U1424 (N_1424,N_582,N_797);
and U1425 (N_1425,N_165,N_1241);
nor U1426 (N_1426,N_635,N_1058);
or U1427 (N_1427,N_310,N_456);
nand U1428 (N_1428,N_222,N_1197);
nor U1429 (N_1429,N_609,N_796);
xnor U1430 (N_1430,N_1078,N_421);
or U1431 (N_1431,N_137,N_501);
nor U1432 (N_1432,N_363,N_158);
nand U1433 (N_1433,N_0,N_923);
nand U1434 (N_1434,N_660,N_355);
and U1435 (N_1435,N_986,N_772);
nor U1436 (N_1436,N_532,N_284);
nand U1437 (N_1437,N_953,N_24);
nand U1438 (N_1438,N_598,N_154);
and U1439 (N_1439,N_342,N_221);
and U1440 (N_1440,N_933,N_1074);
or U1441 (N_1441,N_577,N_1225);
or U1442 (N_1442,N_736,N_552);
and U1443 (N_1443,N_36,N_406);
nor U1444 (N_1444,N_669,N_863);
or U1445 (N_1445,N_192,N_491);
or U1446 (N_1446,N_304,N_700);
xor U1447 (N_1447,N_276,N_688);
nor U1448 (N_1448,N_961,N_1003);
xor U1449 (N_1449,N_1184,N_317);
nand U1450 (N_1450,N_431,N_48);
xnor U1451 (N_1451,N_74,N_122);
nor U1452 (N_1452,N_524,N_143);
and U1453 (N_1453,N_1165,N_651);
nor U1454 (N_1454,N_808,N_622);
nand U1455 (N_1455,N_641,N_784);
and U1456 (N_1456,N_126,N_823);
xnor U1457 (N_1457,N_277,N_536);
or U1458 (N_1458,N_1190,N_1169);
or U1459 (N_1459,N_51,N_696);
nor U1460 (N_1460,N_469,N_401);
nor U1461 (N_1461,N_534,N_804);
nor U1462 (N_1462,N_754,N_756);
xnor U1463 (N_1463,N_782,N_429);
and U1464 (N_1464,N_1198,N_556);
and U1465 (N_1465,N_1215,N_958);
or U1466 (N_1466,N_328,N_869);
and U1467 (N_1467,N_519,N_416);
and U1468 (N_1468,N_1181,N_268);
xor U1469 (N_1469,N_1248,N_1042);
xnor U1470 (N_1470,N_254,N_1050);
xnor U1471 (N_1471,N_866,N_1167);
and U1472 (N_1472,N_325,N_1052);
xor U1473 (N_1473,N_864,N_404);
xor U1474 (N_1474,N_1053,N_1183);
nor U1475 (N_1475,N_26,N_777);
or U1476 (N_1476,N_141,N_1208);
or U1477 (N_1477,N_67,N_790);
and U1478 (N_1478,N_840,N_1223);
nand U1479 (N_1479,N_762,N_1111);
nor U1480 (N_1480,N_811,N_279);
and U1481 (N_1481,N_447,N_940);
and U1482 (N_1482,N_1158,N_910);
nor U1483 (N_1483,N_972,N_42);
nor U1484 (N_1484,N_657,N_801);
xor U1485 (N_1485,N_4,N_13);
or U1486 (N_1486,N_432,N_1224);
or U1487 (N_1487,N_1144,N_1173);
and U1488 (N_1488,N_89,N_88);
and U1489 (N_1489,N_588,N_803);
or U1490 (N_1490,N_549,N_99);
nand U1491 (N_1491,N_115,N_140);
or U1492 (N_1492,N_1134,N_1090);
xnor U1493 (N_1493,N_218,N_848);
nor U1494 (N_1494,N_171,N_461);
nand U1495 (N_1495,N_239,N_1084);
and U1496 (N_1496,N_307,N_638);
nor U1497 (N_1497,N_139,N_766);
nor U1498 (N_1498,N_393,N_560);
nor U1499 (N_1499,N_64,N_626);
or U1500 (N_1500,N_912,N_901);
or U1501 (N_1501,N_12,N_249);
and U1502 (N_1502,N_572,N_1009);
nor U1503 (N_1503,N_645,N_956);
nand U1504 (N_1504,N_473,N_967);
nor U1505 (N_1505,N_330,N_364);
nand U1506 (N_1506,N_161,N_1122);
xor U1507 (N_1507,N_458,N_995);
nor U1508 (N_1508,N_97,N_1147);
xnor U1509 (N_1509,N_1199,N_308);
nor U1510 (N_1510,N_1138,N_861);
and U1511 (N_1511,N_25,N_1117);
xnor U1512 (N_1512,N_240,N_681);
xor U1513 (N_1513,N_892,N_1120);
xor U1514 (N_1514,N_508,N_647);
or U1515 (N_1515,N_164,N_505);
xnor U1516 (N_1516,N_301,N_637);
nor U1517 (N_1517,N_792,N_236);
and U1518 (N_1518,N_379,N_1103);
nor U1519 (N_1519,N_1152,N_639);
xor U1520 (N_1520,N_707,N_225);
nor U1521 (N_1521,N_755,N_480);
nand U1522 (N_1522,N_720,N_1125);
nand U1523 (N_1523,N_198,N_694);
nor U1524 (N_1524,N_1234,N_770);
or U1525 (N_1525,N_938,N_886);
and U1526 (N_1526,N_386,N_894);
and U1527 (N_1527,N_1004,N_935);
xor U1528 (N_1528,N_839,N_387);
or U1529 (N_1529,N_41,N_1107);
or U1530 (N_1530,N_646,N_465);
nand U1531 (N_1531,N_1112,N_1000);
and U1532 (N_1532,N_987,N_290);
or U1533 (N_1533,N_1065,N_740);
xor U1534 (N_1534,N_525,N_699);
xor U1535 (N_1535,N_1109,N_936);
xor U1536 (N_1536,N_512,N_575);
nor U1537 (N_1537,N_799,N_81);
or U1538 (N_1538,N_341,N_996);
or U1539 (N_1539,N_229,N_771);
nor U1540 (N_1540,N_780,N_561);
or U1541 (N_1541,N_43,N_684);
xnor U1542 (N_1542,N_77,N_372);
nor U1543 (N_1543,N_682,N_1115);
nand U1544 (N_1544,N_1056,N_769);
and U1545 (N_1545,N_434,N_149);
xnor U1546 (N_1546,N_1230,N_305);
and U1547 (N_1547,N_1060,N_791);
or U1548 (N_1548,N_50,N_381);
xnor U1549 (N_1549,N_692,N_33);
nor U1550 (N_1550,N_69,N_917);
or U1551 (N_1551,N_976,N_377);
nor U1552 (N_1552,N_29,N_1028);
xnor U1553 (N_1553,N_888,N_391);
nand U1554 (N_1554,N_513,N_344);
or U1555 (N_1555,N_511,N_499);
and U1556 (N_1556,N_174,N_715);
nand U1557 (N_1557,N_1038,N_282);
or U1558 (N_1558,N_181,N_492);
nor U1559 (N_1559,N_127,N_319);
xnor U1560 (N_1560,N_1132,N_163);
xor U1561 (N_1561,N_540,N_1143);
and U1562 (N_1562,N_926,N_430);
xnor U1563 (N_1563,N_789,N_495);
xor U1564 (N_1564,N_388,N_118);
and U1565 (N_1565,N_1205,N_1022);
and U1566 (N_1566,N_1064,N_30);
or U1567 (N_1567,N_744,N_738);
or U1568 (N_1568,N_865,N_908);
or U1569 (N_1569,N_2,N_1024);
nor U1570 (N_1570,N_95,N_1245);
nor U1571 (N_1571,N_695,N_690);
or U1572 (N_1572,N_1092,N_1238);
nand U1573 (N_1573,N_235,N_712);
xor U1574 (N_1574,N_786,N_227);
nand U1575 (N_1575,N_189,N_1101);
and U1576 (N_1576,N_604,N_905);
xor U1577 (N_1577,N_58,N_911);
and U1578 (N_1578,N_313,N_1128);
and U1579 (N_1579,N_40,N_915);
nor U1580 (N_1580,N_234,N_859);
xnor U1581 (N_1581,N_1067,N_516);
and U1582 (N_1582,N_980,N_795);
xor U1583 (N_1583,N_733,N_403);
nor U1584 (N_1584,N_1162,N_874);
nand U1585 (N_1585,N_1105,N_476);
and U1586 (N_1586,N_9,N_398);
and U1587 (N_1587,N_665,N_119);
nor U1588 (N_1588,N_418,N_862);
xor U1589 (N_1589,N_815,N_76);
nand U1590 (N_1590,N_624,N_977);
nor U1591 (N_1591,N_202,N_131);
xor U1592 (N_1592,N_1127,N_632);
and U1593 (N_1593,N_683,N_1185);
nor U1594 (N_1594,N_217,N_701);
nor U1595 (N_1595,N_621,N_1088);
nor U1596 (N_1596,N_71,N_1247);
and U1597 (N_1597,N_959,N_880);
nor U1598 (N_1598,N_162,N_957);
nand U1599 (N_1599,N_558,N_749);
nor U1600 (N_1600,N_93,N_86);
and U1601 (N_1601,N_526,N_1126);
or U1602 (N_1602,N_1214,N_169);
nand U1603 (N_1603,N_484,N_180);
xnor U1604 (N_1604,N_717,N_332);
xnor U1605 (N_1605,N_15,N_822);
or U1606 (N_1606,N_352,N_596);
nor U1607 (N_1607,N_891,N_1227);
nand U1608 (N_1608,N_1135,N_629);
and U1609 (N_1609,N_351,N_785);
or U1610 (N_1610,N_921,N_623);
and U1611 (N_1611,N_396,N_455);
nor U1612 (N_1612,N_593,N_414);
nor U1613 (N_1613,N_1029,N_1108);
nor U1614 (N_1614,N_287,N_850);
and U1615 (N_1615,N_529,N_599);
xor U1616 (N_1616,N_844,N_1192);
or U1617 (N_1617,N_1068,N_260);
or U1618 (N_1618,N_521,N_1133);
xnor U1619 (N_1619,N_1155,N_667);
or U1620 (N_1620,N_1061,N_263);
nor U1621 (N_1621,N_685,N_783);
xor U1622 (N_1622,N_155,N_295);
nand U1623 (N_1623,N_1071,N_1020);
or U1624 (N_1624,N_966,N_204);
nor U1625 (N_1625,N_477,N_515);
xor U1626 (N_1626,N_1025,N_975);
or U1627 (N_1627,N_454,N_748);
and U1628 (N_1628,N_576,N_1194);
or U1629 (N_1629,N_132,N_636);
xor U1630 (N_1630,N_106,N_383);
nand U1631 (N_1631,N_444,N_439);
nor U1632 (N_1632,N_845,N_1124);
nand U1633 (N_1633,N_1177,N_346);
xnor U1634 (N_1634,N_497,N_490);
xor U1635 (N_1635,N_1077,N_618);
or U1636 (N_1636,N_1007,N_107);
or U1637 (N_1637,N_450,N_787);
nor U1638 (N_1638,N_52,N_35);
nor U1639 (N_1639,N_19,N_725);
and U1640 (N_1640,N_676,N_1166);
or U1641 (N_1641,N_83,N_213);
nand U1642 (N_1642,N_286,N_20);
xor U1643 (N_1643,N_356,N_842);
and U1644 (N_1644,N_303,N_537);
nor U1645 (N_1645,N_38,N_326);
or U1646 (N_1646,N_274,N_256);
nand U1647 (N_1647,N_142,N_354);
and U1648 (N_1648,N_498,N_928);
and U1649 (N_1649,N_186,N_299);
nor U1650 (N_1650,N_741,N_605);
nand U1651 (N_1651,N_205,N_655);
or U1652 (N_1652,N_116,N_269);
nand U1653 (N_1653,N_504,N_1017);
or U1654 (N_1654,N_440,N_483);
xor U1655 (N_1655,N_65,N_727);
nand U1656 (N_1656,N_23,N_487);
nor U1657 (N_1657,N_462,N_496);
and U1658 (N_1658,N_530,N_1116);
or U1659 (N_1659,N_514,N_990);
and U1660 (N_1660,N_233,N_232);
and U1661 (N_1661,N_973,N_125);
and U1662 (N_1662,N_1012,N_634);
nand U1663 (N_1663,N_724,N_1216);
and U1664 (N_1664,N_378,N_1231);
and U1665 (N_1665,N_413,N_1235);
or U1666 (N_1666,N_374,N_964);
or U1667 (N_1667,N_59,N_768);
and U1668 (N_1668,N_98,N_353);
nor U1669 (N_1669,N_675,N_778);
nor U1670 (N_1670,N_1032,N_574);
nor U1671 (N_1671,N_100,N_231);
nand U1672 (N_1672,N_802,N_931);
nor U1673 (N_1673,N_709,N_464);
or U1674 (N_1674,N_311,N_152);
nor U1675 (N_1675,N_652,N_500);
xor U1676 (N_1676,N_53,N_1172);
and U1677 (N_1677,N_672,N_242);
nor U1678 (N_1678,N_265,N_680);
or U1679 (N_1679,N_563,N_442);
xnor U1680 (N_1680,N_96,N_829);
xor U1681 (N_1681,N_616,N_1095);
xor U1682 (N_1682,N_302,N_743);
nand U1683 (N_1683,N_1097,N_362);
or U1684 (N_1684,N_613,N_257);
nor U1685 (N_1685,N_197,N_1157);
and U1686 (N_1686,N_11,N_314);
xor U1687 (N_1687,N_459,N_742);
nand U1688 (N_1688,N_185,N_726);
and U1689 (N_1689,N_1066,N_546);
xnor U1690 (N_1690,N_805,N_991);
and U1691 (N_1691,N_57,N_1023);
xor U1692 (N_1692,N_591,N_250);
nor U1693 (N_1693,N_860,N_1118);
and U1694 (N_1694,N_105,N_3);
and U1695 (N_1695,N_909,N_1174);
nand U1696 (N_1696,N_871,N_136);
nand U1697 (N_1697,N_428,N_587);
and U1698 (N_1698,N_1232,N_971);
nand U1699 (N_1699,N_1189,N_79);
and U1700 (N_1700,N_267,N_151);
nand U1701 (N_1701,N_448,N_44);
xor U1702 (N_1702,N_764,N_190);
or U1703 (N_1703,N_735,N_687);
xnor U1704 (N_1704,N_689,N_408);
nor U1705 (N_1705,N_1013,N_502);
nand U1706 (N_1706,N_668,N_271);
and U1707 (N_1707,N_349,N_1041);
or U1708 (N_1708,N_331,N_1087);
xnor U1709 (N_1709,N_855,N_427);
or U1710 (N_1710,N_262,N_392);
nand U1711 (N_1711,N_1027,N_606);
nand U1712 (N_1712,N_170,N_875);
and U1713 (N_1713,N_244,N_453);
or U1714 (N_1714,N_1106,N_203);
nand U1715 (N_1715,N_1139,N_320);
xor U1716 (N_1716,N_507,N_350);
nor U1717 (N_1717,N_437,N_974);
nor U1718 (N_1718,N_423,N_1210);
nor U1719 (N_1719,N_339,N_120);
xnor U1720 (N_1720,N_567,N_930);
nand U1721 (N_1721,N_1055,N_653);
or U1722 (N_1722,N_1081,N_542);
nor U1723 (N_1723,N_336,N_1148);
and U1724 (N_1724,N_109,N_918);
xor U1725 (N_1725,N_46,N_879);
or U1726 (N_1726,N_528,N_825);
or U1727 (N_1727,N_208,N_559);
or U1728 (N_1728,N_293,N_195);
nor U1729 (N_1729,N_1196,N_150);
nand U1730 (N_1730,N_108,N_85);
xnor U1731 (N_1731,N_135,N_1213);
or U1732 (N_1732,N_828,N_898);
or U1733 (N_1733,N_659,N_965);
or U1734 (N_1734,N_603,N_402);
nand U1735 (N_1735,N_61,N_798);
nor U1736 (N_1736,N_207,N_485);
or U1737 (N_1737,N_385,N_433);
xnor U1738 (N_1738,N_553,N_251);
nand U1739 (N_1739,N_704,N_734);
and U1740 (N_1740,N_138,N_708);
and U1741 (N_1741,N_806,N_1140);
or U1742 (N_1742,N_747,N_113);
xnor U1743 (N_1743,N_183,N_1123);
and U1744 (N_1744,N_584,N_1026);
xor U1745 (N_1745,N_494,N_1202);
nand U1746 (N_1746,N_375,N_273);
and U1747 (N_1747,N_129,N_818);
nor U1748 (N_1748,N_173,N_1080);
nor U1749 (N_1749,N_746,N_838);
and U1750 (N_1750,N_1211,N_1036);
and U1751 (N_1751,N_594,N_774);
xor U1752 (N_1752,N_1001,N_1243);
nor U1753 (N_1753,N_175,N_261);
and U1754 (N_1754,N_543,N_1240);
nand U1755 (N_1755,N_422,N_438);
or U1756 (N_1756,N_615,N_920);
xnor U1757 (N_1757,N_369,N_831);
and U1758 (N_1758,N_573,N_75);
and U1759 (N_1759,N_281,N_1037);
nor U1760 (N_1760,N_941,N_674);
xor U1761 (N_1761,N_794,N_730);
xnor U1762 (N_1762,N_1039,N_7);
nor U1763 (N_1763,N_819,N_345);
nor U1764 (N_1764,N_1229,N_592);
nor U1765 (N_1765,N_475,N_285);
nand U1766 (N_1766,N_1156,N_586);
or U1767 (N_1767,N_775,N_1180);
xnor U1768 (N_1768,N_1091,N_824);
nand U1769 (N_1769,N_998,N_555);
nor U1770 (N_1770,N_278,N_368);
and U1771 (N_1771,N_779,N_1021);
or U1772 (N_1772,N_425,N_343);
nor U1773 (N_1773,N_527,N_753);
and U1774 (N_1774,N_380,N_45);
or U1775 (N_1775,N_988,N_114);
and U1776 (N_1776,N_188,N_510);
nand U1777 (N_1777,N_723,N_223);
xor U1778 (N_1778,N_620,N_562);
xor U1779 (N_1779,N_1142,N_1006);
xnor U1780 (N_1780,N_731,N_283);
and U1781 (N_1781,N_946,N_884);
nand U1782 (N_1782,N_226,N_1099);
xor U1783 (N_1783,N_31,N_611);
nor U1784 (N_1784,N_306,N_264);
nor U1785 (N_1785,N_92,N_411);
xnor U1786 (N_1786,N_853,N_291);
or U1787 (N_1787,N_1179,N_944);
xnor U1788 (N_1788,N_56,N_1);
or U1789 (N_1789,N_367,N_327);
and U1790 (N_1790,N_934,N_160);
nor U1791 (N_1791,N_1014,N_955);
nor U1792 (N_1792,N_73,N_62);
xnor U1793 (N_1793,N_564,N_21);
nand U1794 (N_1794,N_872,N_752);
or U1795 (N_1795,N_467,N_673);
nor U1796 (N_1796,N_948,N_919);
nor U1797 (N_1797,N_1163,N_1076);
nor U1798 (N_1798,N_1217,N_177);
or U1799 (N_1799,N_821,N_334);
xnor U1800 (N_1800,N_1136,N_662);
or U1801 (N_1801,N_893,N_883);
xnor U1802 (N_1802,N_691,N_193);
or U1803 (N_1803,N_472,N_1203);
nor U1804 (N_1804,N_360,N_176);
nor U1805 (N_1805,N_335,N_978);
xor U1806 (N_1806,N_737,N_147);
and U1807 (N_1807,N_714,N_939);
nor U1808 (N_1808,N_1175,N_627);
and U1809 (N_1809,N_1170,N_776);
nand U1810 (N_1810,N_903,N_951);
and U1811 (N_1811,N_443,N_1093);
and U1812 (N_1812,N_702,N_1018);
nor U1813 (N_1813,N_1033,N_650);
or U1814 (N_1814,N_1237,N_1137);
nand U1815 (N_1815,N_548,N_807);
nor U1816 (N_1816,N_902,N_1030);
nand U1817 (N_1817,N_997,N_318);
or U1818 (N_1818,N_272,N_1069);
and U1819 (N_1819,N_765,N_156);
or U1820 (N_1820,N_1236,N_858);
or U1821 (N_1821,N_581,N_678);
nand U1822 (N_1822,N_1131,N_245);
or U1823 (N_1823,N_666,N_60);
nor U1824 (N_1824,N_322,N_989);
or U1825 (N_1825,N_482,N_1073);
or U1826 (N_1826,N_452,N_1008);
xnor U1827 (N_1827,N_390,N_315);
xor U1828 (N_1828,N_179,N_209);
and U1829 (N_1829,N_814,N_216);
xor U1830 (N_1830,N_686,N_619);
and U1831 (N_1831,N_1204,N_200);
xnor U1832 (N_1832,N_321,N_670);
nand U1833 (N_1833,N_70,N_962);
xor U1834 (N_1834,N_900,N_628);
or U1835 (N_1835,N_451,N_719);
nor U1836 (N_1836,N_196,N_1110);
and U1837 (N_1837,N_481,N_16);
nor U1838 (N_1838,N_420,N_827);
or U1839 (N_1839,N_710,N_8);
xnor U1840 (N_1840,N_124,N_925);
nand U1841 (N_1841,N_333,N_488);
or U1842 (N_1842,N_144,N_470);
nand U1843 (N_1843,N_194,N_199);
or U1844 (N_1844,N_87,N_924);
nor U1845 (N_1845,N_371,N_78);
xor U1846 (N_1846,N_80,N_1102);
or U1847 (N_1847,N_506,N_191);
nor U1848 (N_1848,N_1149,N_5);
xnor U1849 (N_1849,N_123,N_1207);
or U1850 (N_1850,N_247,N_1051);
nor U1851 (N_1851,N_857,N_846);
or U1852 (N_1852,N_1048,N_14);
or U1853 (N_1853,N_446,N_1130);
or U1854 (N_1854,N_954,N_759);
nor U1855 (N_1855,N_1075,N_904);
nor U1856 (N_1856,N_1085,N_471);
and U1857 (N_1857,N_168,N_39);
or U1858 (N_1858,N_544,N_1114);
and U1859 (N_1859,N_259,N_580);
nor U1860 (N_1860,N_703,N_215);
or U1861 (N_1861,N_316,N_1171);
or U1862 (N_1862,N_1096,N_1034);
xnor U1863 (N_1863,N_523,N_27);
nor U1864 (N_1864,N_729,N_309);
nand U1865 (N_1865,N_211,N_237);
nor U1866 (N_1866,N_533,N_1176);
xnor U1867 (N_1867,N_1016,N_1219);
nor U1868 (N_1868,N_982,N_981);
or U1869 (N_1869,N_153,N_816);
nor U1870 (N_1870,N_146,N_656);
and U1871 (N_1871,N_1206,N_1082);
or U1872 (N_1872,N_897,N_854);
nand U1873 (N_1873,N_570,N_751);
xor U1874 (N_1874,N_970,N_1121);
nand U1875 (N_1875,N_1097,N_1122);
nand U1876 (N_1876,N_348,N_327);
xnor U1877 (N_1877,N_102,N_562);
nor U1878 (N_1878,N_379,N_1131);
nand U1879 (N_1879,N_922,N_884);
and U1880 (N_1880,N_788,N_364);
and U1881 (N_1881,N_909,N_499);
nor U1882 (N_1882,N_12,N_911);
or U1883 (N_1883,N_298,N_99);
xor U1884 (N_1884,N_1195,N_813);
nand U1885 (N_1885,N_1108,N_881);
xor U1886 (N_1886,N_594,N_726);
xor U1887 (N_1887,N_446,N_742);
nand U1888 (N_1888,N_298,N_158);
and U1889 (N_1889,N_1104,N_911);
or U1890 (N_1890,N_517,N_60);
or U1891 (N_1891,N_775,N_1200);
xnor U1892 (N_1892,N_488,N_469);
nand U1893 (N_1893,N_960,N_504);
nor U1894 (N_1894,N_1010,N_199);
or U1895 (N_1895,N_114,N_224);
nor U1896 (N_1896,N_1092,N_1021);
nand U1897 (N_1897,N_977,N_1015);
nor U1898 (N_1898,N_240,N_210);
nor U1899 (N_1899,N_511,N_196);
nand U1900 (N_1900,N_1161,N_651);
xnor U1901 (N_1901,N_1004,N_866);
or U1902 (N_1902,N_157,N_559);
nor U1903 (N_1903,N_558,N_532);
and U1904 (N_1904,N_120,N_50);
nand U1905 (N_1905,N_169,N_630);
nor U1906 (N_1906,N_248,N_101);
or U1907 (N_1907,N_276,N_341);
or U1908 (N_1908,N_207,N_84);
or U1909 (N_1909,N_1001,N_338);
nor U1910 (N_1910,N_1232,N_612);
nand U1911 (N_1911,N_305,N_307);
nor U1912 (N_1912,N_1015,N_1169);
or U1913 (N_1913,N_777,N_473);
or U1914 (N_1914,N_1071,N_818);
nor U1915 (N_1915,N_322,N_562);
nand U1916 (N_1916,N_1217,N_683);
nand U1917 (N_1917,N_460,N_498);
nand U1918 (N_1918,N_916,N_945);
and U1919 (N_1919,N_55,N_1107);
nand U1920 (N_1920,N_1211,N_837);
xor U1921 (N_1921,N_113,N_978);
and U1922 (N_1922,N_111,N_289);
xnor U1923 (N_1923,N_466,N_1105);
nand U1924 (N_1924,N_236,N_73);
nor U1925 (N_1925,N_123,N_1055);
xnor U1926 (N_1926,N_1185,N_968);
xnor U1927 (N_1927,N_805,N_619);
or U1928 (N_1928,N_996,N_472);
xnor U1929 (N_1929,N_817,N_591);
and U1930 (N_1930,N_213,N_1221);
nand U1931 (N_1931,N_1060,N_216);
or U1932 (N_1932,N_258,N_57);
nand U1933 (N_1933,N_1219,N_239);
or U1934 (N_1934,N_1004,N_818);
nand U1935 (N_1935,N_563,N_292);
xor U1936 (N_1936,N_659,N_277);
nor U1937 (N_1937,N_1122,N_528);
and U1938 (N_1938,N_526,N_283);
nand U1939 (N_1939,N_618,N_244);
nand U1940 (N_1940,N_294,N_1211);
nor U1941 (N_1941,N_254,N_344);
nor U1942 (N_1942,N_925,N_112);
nor U1943 (N_1943,N_516,N_792);
and U1944 (N_1944,N_458,N_829);
nand U1945 (N_1945,N_981,N_853);
nand U1946 (N_1946,N_594,N_268);
or U1947 (N_1947,N_1209,N_14);
and U1948 (N_1948,N_972,N_503);
nor U1949 (N_1949,N_67,N_861);
xnor U1950 (N_1950,N_280,N_76);
or U1951 (N_1951,N_1041,N_471);
nor U1952 (N_1952,N_870,N_118);
nand U1953 (N_1953,N_128,N_697);
nand U1954 (N_1954,N_232,N_325);
xnor U1955 (N_1955,N_230,N_446);
and U1956 (N_1956,N_200,N_739);
xor U1957 (N_1957,N_712,N_432);
nor U1958 (N_1958,N_664,N_354);
nand U1959 (N_1959,N_996,N_305);
and U1960 (N_1960,N_857,N_419);
nor U1961 (N_1961,N_54,N_79);
xnor U1962 (N_1962,N_788,N_422);
or U1963 (N_1963,N_7,N_829);
xnor U1964 (N_1964,N_132,N_544);
xor U1965 (N_1965,N_979,N_785);
nand U1966 (N_1966,N_297,N_901);
or U1967 (N_1967,N_744,N_340);
or U1968 (N_1968,N_860,N_796);
and U1969 (N_1969,N_742,N_1227);
xnor U1970 (N_1970,N_1219,N_179);
xnor U1971 (N_1971,N_945,N_415);
or U1972 (N_1972,N_618,N_1175);
and U1973 (N_1973,N_85,N_1102);
or U1974 (N_1974,N_687,N_896);
and U1975 (N_1975,N_1215,N_836);
nand U1976 (N_1976,N_655,N_443);
or U1977 (N_1977,N_923,N_490);
nand U1978 (N_1978,N_813,N_260);
xnor U1979 (N_1979,N_916,N_62);
and U1980 (N_1980,N_147,N_978);
nand U1981 (N_1981,N_756,N_1054);
xor U1982 (N_1982,N_204,N_1189);
nor U1983 (N_1983,N_191,N_239);
nand U1984 (N_1984,N_430,N_170);
or U1985 (N_1985,N_563,N_807);
and U1986 (N_1986,N_649,N_1201);
nand U1987 (N_1987,N_10,N_987);
or U1988 (N_1988,N_329,N_839);
nand U1989 (N_1989,N_9,N_947);
nand U1990 (N_1990,N_1112,N_332);
and U1991 (N_1991,N_667,N_592);
nand U1992 (N_1992,N_590,N_831);
or U1993 (N_1993,N_433,N_145);
and U1994 (N_1994,N_472,N_521);
xor U1995 (N_1995,N_1208,N_1229);
nand U1996 (N_1996,N_1189,N_681);
or U1997 (N_1997,N_637,N_573);
or U1998 (N_1998,N_234,N_270);
or U1999 (N_1999,N_1123,N_512);
nor U2000 (N_2000,N_1049,N_1114);
or U2001 (N_2001,N_748,N_356);
or U2002 (N_2002,N_592,N_539);
or U2003 (N_2003,N_836,N_708);
and U2004 (N_2004,N_2,N_604);
nor U2005 (N_2005,N_387,N_755);
or U2006 (N_2006,N_47,N_805);
nor U2007 (N_2007,N_346,N_345);
and U2008 (N_2008,N_991,N_574);
or U2009 (N_2009,N_404,N_518);
or U2010 (N_2010,N_147,N_249);
nor U2011 (N_2011,N_327,N_225);
or U2012 (N_2012,N_951,N_422);
xnor U2013 (N_2013,N_837,N_696);
or U2014 (N_2014,N_288,N_761);
and U2015 (N_2015,N_1154,N_829);
nand U2016 (N_2016,N_375,N_27);
and U2017 (N_2017,N_1073,N_291);
nor U2018 (N_2018,N_684,N_554);
or U2019 (N_2019,N_353,N_101);
or U2020 (N_2020,N_919,N_718);
nor U2021 (N_2021,N_514,N_726);
nand U2022 (N_2022,N_72,N_471);
and U2023 (N_2023,N_314,N_111);
and U2024 (N_2024,N_1081,N_218);
and U2025 (N_2025,N_736,N_757);
xor U2026 (N_2026,N_715,N_1208);
nand U2027 (N_2027,N_197,N_854);
or U2028 (N_2028,N_1009,N_787);
nand U2029 (N_2029,N_1211,N_125);
or U2030 (N_2030,N_1183,N_387);
nor U2031 (N_2031,N_680,N_205);
and U2032 (N_2032,N_1233,N_512);
nor U2033 (N_2033,N_979,N_133);
xor U2034 (N_2034,N_887,N_790);
nand U2035 (N_2035,N_648,N_1);
xor U2036 (N_2036,N_722,N_748);
and U2037 (N_2037,N_256,N_138);
and U2038 (N_2038,N_500,N_37);
nand U2039 (N_2039,N_229,N_488);
nor U2040 (N_2040,N_1164,N_450);
and U2041 (N_2041,N_721,N_1017);
and U2042 (N_2042,N_259,N_1061);
xnor U2043 (N_2043,N_935,N_799);
nor U2044 (N_2044,N_971,N_1079);
nand U2045 (N_2045,N_733,N_594);
xnor U2046 (N_2046,N_1007,N_142);
and U2047 (N_2047,N_715,N_150);
xnor U2048 (N_2048,N_205,N_626);
xor U2049 (N_2049,N_800,N_1200);
and U2050 (N_2050,N_1030,N_425);
nand U2051 (N_2051,N_1038,N_891);
and U2052 (N_2052,N_974,N_240);
or U2053 (N_2053,N_18,N_441);
xor U2054 (N_2054,N_976,N_1160);
or U2055 (N_2055,N_677,N_1047);
nor U2056 (N_2056,N_268,N_781);
nand U2057 (N_2057,N_68,N_211);
nor U2058 (N_2058,N_926,N_1006);
and U2059 (N_2059,N_937,N_706);
nor U2060 (N_2060,N_43,N_149);
xor U2061 (N_2061,N_916,N_357);
and U2062 (N_2062,N_1170,N_665);
xor U2063 (N_2063,N_932,N_513);
xnor U2064 (N_2064,N_130,N_500);
or U2065 (N_2065,N_1040,N_711);
nor U2066 (N_2066,N_949,N_1190);
nand U2067 (N_2067,N_327,N_293);
nand U2068 (N_2068,N_1137,N_772);
nor U2069 (N_2069,N_1067,N_543);
xnor U2070 (N_2070,N_1008,N_219);
and U2071 (N_2071,N_657,N_426);
nor U2072 (N_2072,N_79,N_608);
and U2073 (N_2073,N_4,N_1151);
or U2074 (N_2074,N_710,N_467);
nor U2075 (N_2075,N_1059,N_677);
nand U2076 (N_2076,N_181,N_290);
xnor U2077 (N_2077,N_60,N_1125);
and U2078 (N_2078,N_66,N_616);
nor U2079 (N_2079,N_355,N_1152);
and U2080 (N_2080,N_650,N_361);
xor U2081 (N_2081,N_1066,N_1246);
xor U2082 (N_2082,N_716,N_778);
or U2083 (N_2083,N_64,N_615);
xnor U2084 (N_2084,N_1078,N_48);
nand U2085 (N_2085,N_385,N_848);
and U2086 (N_2086,N_361,N_515);
xnor U2087 (N_2087,N_463,N_788);
and U2088 (N_2088,N_696,N_200);
nand U2089 (N_2089,N_1163,N_1044);
or U2090 (N_2090,N_820,N_1080);
nand U2091 (N_2091,N_87,N_82);
and U2092 (N_2092,N_695,N_1103);
and U2093 (N_2093,N_33,N_1095);
and U2094 (N_2094,N_115,N_854);
and U2095 (N_2095,N_751,N_55);
and U2096 (N_2096,N_219,N_647);
xor U2097 (N_2097,N_210,N_721);
or U2098 (N_2098,N_1205,N_419);
nor U2099 (N_2099,N_165,N_890);
nand U2100 (N_2100,N_205,N_1180);
xor U2101 (N_2101,N_595,N_1126);
nand U2102 (N_2102,N_809,N_236);
nand U2103 (N_2103,N_611,N_616);
or U2104 (N_2104,N_903,N_1016);
nand U2105 (N_2105,N_384,N_640);
and U2106 (N_2106,N_535,N_702);
or U2107 (N_2107,N_985,N_297);
nor U2108 (N_2108,N_795,N_757);
or U2109 (N_2109,N_833,N_51);
and U2110 (N_2110,N_752,N_258);
nor U2111 (N_2111,N_1050,N_290);
and U2112 (N_2112,N_218,N_881);
and U2113 (N_2113,N_316,N_767);
or U2114 (N_2114,N_1249,N_358);
and U2115 (N_2115,N_71,N_534);
or U2116 (N_2116,N_696,N_663);
xnor U2117 (N_2117,N_84,N_431);
nand U2118 (N_2118,N_813,N_679);
and U2119 (N_2119,N_17,N_299);
nand U2120 (N_2120,N_620,N_475);
or U2121 (N_2121,N_1022,N_753);
nand U2122 (N_2122,N_672,N_1248);
nand U2123 (N_2123,N_1210,N_567);
or U2124 (N_2124,N_464,N_341);
or U2125 (N_2125,N_182,N_852);
nand U2126 (N_2126,N_626,N_536);
nor U2127 (N_2127,N_1071,N_364);
nor U2128 (N_2128,N_1233,N_903);
xor U2129 (N_2129,N_613,N_652);
and U2130 (N_2130,N_662,N_1137);
xnor U2131 (N_2131,N_999,N_246);
xor U2132 (N_2132,N_18,N_882);
nand U2133 (N_2133,N_320,N_1128);
nor U2134 (N_2134,N_833,N_542);
nand U2135 (N_2135,N_669,N_281);
xor U2136 (N_2136,N_114,N_919);
or U2137 (N_2137,N_599,N_1109);
xnor U2138 (N_2138,N_121,N_917);
and U2139 (N_2139,N_1157,N_299);
or U2140 (N_2140,N_1077,N_272);
or U2141 (N_2141,N_801,N_994);
nor U2142 (N_2142,N_1130,N_976);
or U2143 (N_2143,N_459,N_193);
xnor U2144 (N_2144,N_425,N_931);
nor U2145 (N_2145,N_61,N_172);
nor U2146 (N_2146,N_922,N_852);
or U2147 (N_2147,N_148,N_589);
nor U2148 (N_2148,N_1178,N_25);
nor U2149 (N_2149,N_175,N_876);
nand U2150 (N_2150,N_537,N_803);
and U2151 (N_2151,N_339,N_958);
or U2152 (N_2152,N_587,N_328);
or U2153 (N_2153,N_1003,N_173);
xor U2154 (N_2154,N_790,N_1033);
nand U2155 (N_2155,N_680,N_444);
xor U2156 (N_2156,N_801,N_52);
and U2157 (N_2157,N_659,N_720);
or U2158 (N_2158,N_51,N_107);
or U2159 (N_2159,N_795,N_402);
xnor U2160 (N_2160,N_933,N_916);
and U2161 (N_2161,N_441,N_684);
and U2162 (N_2162,N_447,N_113);
or U2163 (N_2163,N_354,N_289);
and U2164 (N_2164,N_514,N_276);
and U2165 (N_2165,N_1073,N_1006);
and U2166 (N_2166,N_806,N_777);
or U2167 (N_2167,N_1127,N_1091);
or U2168 (N_2168,N_288,N_1097);
xor U2169 (N_2169,N_215,N_598);
xor U2170 (N_2170,N_865,N_1196);
or U2171 (N_2171,N_109,N_1088);
and U2172 (N_2172,N_628,N_748);
nor U2173 (N_2173,N_226,N_14);
nor U2174 (N_2174,N_960,N_235);
and U2175 (N_2175,N_793,N_673);
xor U2176 (N_2176,N_697,N_1223);
or U2177 (N_2177,N_782,N_714);
nand U2178 (N_2178,N_946,N_262);
or U2179 (N_2179,N_813,N_238);
nand U2180 (N_2180,N_409,N_436);
nand U2181 (N_2181,N_505,N_957);
nand U2182 (N_2182,N_898,N_923);
nand U2183 (N_2183,N_1164,N_1071);
and U2184 (N_2184,N_432,N_524);
xor U2185 (N_2185,N_100,N_486);
nand U2186 (N_2186,N_140,N_94);
and U2187 (N_2187,N_1068,N_951);
or U2188 (N_2188,N_719,N_805);
nand U2189 (N_2189,N_852,N_357);
and U2190 (N_2190,N_1018,N_910);
or U2191 (N_2191,N_717,N_1243);
nor U2192 (N_2192,N_285,N_157);
or U2193 (N_2193,N_238,N_326);
nor U2194 (N_2194,N_680,N_591);
or U2195 (N_2195,N_491,N_1043);
xnor U2196 (N_2196,N_857,N_683);
xor U2197 (N_2197,N_783,N_991);
xnor U2198 (N_2198,N_542,N_608);
or U2199 (N_2199,N_1203,N_199);
or U2200 (N_2200,N_51,N_61);
nand U2201 (N_2201,N_196,N_449);
or U2202 (N_2202,N_410,N_471);
nand U2203 (N_2203,N_827,N_326);
nand U2204 (N_2204,N_982,N_1064);
and U2205 (N_2205,N_839,N_981);
nand U2206 (N_2206,N_316,N_434);
and U2207 (N_2207,N_707,N_400);
nor U2208 (N_2208,N_678,N_75);
and U2209 (N_2209,N_118,N_301);
and U2210 (N_2210,N_685,N_1125);
and U2211 (N_2211,N_176,N_932);
and U2212 (N_2212,N_462,N_1215);
nand U2213 (N_2213,N_241,N_31);
nand U2214 (N_2214,N_282,N_241);
or U2215 (N_2215,N_767,N_453);
xor U2216 (N_2216,N_815,N_106);
xor U2217 (N_2217,N_1017,N_781);
nand U2218 (N_2218,N_1084,N_132);
and U2219 (N_2219,N_515,N_97);
and U2220 (N_2220,N_552,N_674);
nand U2221 (N_2221,N_221,N_1112);
nor U2222 (N_2222,N_633,N_770);
nand U2223 (N_2223,N_647,N_369);
or U2224 (N_2224,N_965,N_350);
nor U2225 (N_2225,N_1000,N_437);
and U2226 (N_2226,N_408,N_1146);
and U2227 (N_2227,N_333,N_1004);
xnor U2228 (N_2228,N_871,N_1063);
or U2229 (N_2229,N_1027,N_17);
nand U2230 (N_2230,N_667,N_252);
nor U2231 (N_2231,N_411,N_1129);
xor U2232 (N_2232,N_159,N_41);
or U2233 (N_2233,N_728,N_513);
xnor U2234 (N_2234,N_1203,N_1092);
nand U2235 (N_2235,N_360,N_997);
xor U2236 (N_2236,N_232,N_54);
nand U2237 (N_2237,N_919,N_750);
nor U2238 (N_2238,N_398,N_208);
nand U2239 (N_2239,N_841,N_746);
nand U2240 (N_2240,N_243,N_787);
nand U2241 (N_2241,N_669,N_1239);
and U2242 (N_2242,N_923,N_675);
nand U2243 (N_2243,N_49,N_264);
and U2244 (N_2244,N_355,N_393);
xnor U2245 (N_2245,N_940,N_397);
nand U2246 (N_2246,N_352,N_397);
and U2247 (N_2247,N_317,N_1237);
and U2248 (N_2248,N_1198,N_392);
and U2249 (N_2249,N_1009,N_40);
xor U2250 (N_2250,N_453,N_411);
xnor U2251 (N_2251,N_132,N_1073);
nand U2252 (N_2252,N_330,N_1131);
or U2253 (N_2253,N_316,N_242);
or U2254 (N_2254,N_112,N_396);
and U2255 (N_2255,N_964,N_813);
or U2256 (N_2256,N_247,N_1006);
nand U2257 (N_2257,N_1046,N_227);
nand U2258 (N_2258,N_604,N_364);
xor U2259 (N_2259,N_1087,N_1226);
nand U2260 (N_2260,N_730,N_79);
or U2261 (N_2261,N_181,N_564);
xor U2262 (N_2262,N_32,N_808);
nor U2263 (N_2263,N_487,N_250);
or U2264 (N_2264,N_1085,N_703);
nand U2265 (N_2265,N_1203,N_1010);
nand U2266 (N_2266,N_229,N_895);
nor U2267 (N_2267,N_1019,N_242);
xor U2268 (N_2268,N_915,N_736);
or U2269 (N_2269,N_546,N_936);
and U2270 (N_2270,N_808,N_305);
nand U2271 (N_2271,N_448,N_184);
or U2272 (N_2272,N_592,N_409);
xor U2273 (N_2273,N_818,N_755);
and U2274 (N_2274,N_414,N_254);
nor U2275 (N_2275,N_861,N_821);
or U2276 (N_2276,N_722,N_1241);
or U2277 (N_2277,N_345,N_1148);
nor U2278 (N_2278,N_260,N_144);
or U2279 (N_2279,N_570,N_368);
and U2280 (N_2280,N_913,N_572);
nand U2281 (N_2281,N_1170,N_536);
or U2282 (N_2282,N_839,N_218);
nand U2283 (N_2283,N_620,N_950);
nand U2284 (N_2284,N_103,N_55);
and U2285 (N_2285,N_58,N_720);
and U2286 (N_2286,N_77,N_1045);
or U2287 (N_2287,N_1241,N_188);
or U2288 (N_2288,N_515,N_1079);
and U2289 (N_2289,N_543,N_970);
and U2290 (N_2290,N_874,N_246);
nand U2291 (N_2291,N_79,N_444);
or U2292 (N_2292,N_105,N_936);
xor U2293 (N_2293,N_604,N_1065);
xor U2294 (N_2294,N_926,N_670);
and U2295 (N_2295,N_840,N_598);
and U2296 (N_2296,N_80,N_645);
nand U2297 (N_2297,N_1140,N_518);
and U2298 (N_2298,N_976,N_23);
xnor U2299 (N_2299,N_1119,N_1017);
or U2300 (N_2300,N_69,N_238);
nand U2301 (N_2301,N_823,N_585);
nand U2302 (N_2302,N_302,N_122);
or U2303 (N_2303,N_971,N_525);
or U2304 (N_2304,N_228,N_525);
xnor U2305 (N_2305,N_792,N_1092);
nor U2306 (N_2306,N_1134,N_954);
or U2307 (N_2307,N_188,N_818);
or U2308 (N_2308,N_932,N_215);
nand U2309 (N_2309,N_514,N_718);
nor U2310 (N_2310,N_134,N_454);
or U2311 (N_2311,N_563,N_199);
xor U2312 (N_2312,N_674,N_252);
and U2313 (N_2313,N_1177,N_528);
nand U2314 (N_2314,N_996,N_1244);
xor U2315 (N_2315,N_215,N_202);
xor U2316 (N_2316,N_525,N_745);
or U2317 (N_2317,N_1203,N_129);
nand U2318 (N_2318,N_398,N_423);
nor U2319 (N_2319,N_458,N_490);
nand U2320 (N_2320,N_725,N_370);
nor U2321 (N_2321,N_393,N_258);
and U2322 (N_2322,N_961,N_891);
xor U2323 (N_2323,N_620,N_285);
or U2324 (N_2324,N_338,N_567);
nor U2325 (N_2325,N_727,N_1154);
xnor U2326 (N_2326,N_917,N_193);
xnor U2327 (N_2327,N_285,N_508);
and U2328 (N_2328,N_1225,N_1215);
or U2329 (N_2329,N_165,N_987);
and U2330 (N_2330,N_404,N_547);
nor U2331 (N_2331,N_410,N_869);
xnor U2332 (N_2332,N_1193,N_849);
and U2333 (N_2333,N_1240,N_1148);
nor U2334 (N_2334,N_977,N_191);
and U2335 (N_2335,N_1235,N_111);
and U2336 (N_2336,N_1057,N_423);
nor U2337 (N_2337,N_1223,N_890);
and U2338 (N_2338,N_428,N_737);
xnor U2339 (N_2339,N_1207,N_1105);
xnor U2340 (N_2340,N_634,N_883);
or U2341 (N_2341,N_819,N_28);
nand U2342 (N_2342,N_944,N_724);
or U2343 (N_2343,N_878,N_84);
nor U2344 (N_2344,N_795,N_785);
and U2345 (N_2345,N_1195,N_936);
or U2346 (N_2346,N_863,N_1000);
xor U2347 (N_2347,N_697,N_43);
and U2348 (N_2348,N_794,N_192);
or U2349 (N_2349,N_581,N_52);
xor U2350 (N_2350,N_1046,N_937);
nand U2351 (N_2351,N_50,N_457);
and U2352 (N_2352,N_397,N_442);
nand U2353 (N_2353,N_583,N_767);
and U2354 (N_2354,N_828,N_517);
nor U2355 (N_2355,N_98,N_1208);
nor U2356 (N_2356,N_348,N_555);
nand U2357 (N_2357,N_714,N_167);
or U2358 (N_2358,N_1147,N_924);
nand U2359 (N_2359,N_867,N_106);
or U2360 (N_2360,N_684,N_555);
nand U2361 (N_2361,N_410,N_1088);
and U2362 (N_2362,N_398,N_895);
nand U2363 (N_2363,N_1189,N_786);
or U2364 (N_2364,N_286,N_19);
and U2365 (N_2365,N_965,N_35);
and U2366 (N_2366,N_1068,N_1185);
nor U2367 (N_2367,N_15,N_1219);
nand U2368 (N_2368,N_513,N_234);
or U2369 (N_2369,N_1040,N_318);
nand U2370 (N_2370,N_1133,N_706);
and U2371 (N_2371,N_1151,N_923);
nor U2372 (N_2372,N_590,N_1214);
nand U2373 (N_2373,N_544,N_531);
or U2374 (N_2374,N_424,N_313);
and U2375 (N_2375,N_145,N_134);
and U2376 (N_2376,N_1183,N_426);
and U2377 (N_2377,N_676,N_586);
and U2378 (N_2378,N_648,N_469);
and U2379 (N_2379,N_233,N_628);
and U2380 (N_2380,N_1141,N_1161);
nand U2381 (N_2381,N_838,N_20);
xor U2382 (N_2382,N_1215,N_779);
nor U2383 (N_2383,N_351,N_1051);
xnor U2384 (N_2384,N_1040,N_1246);
nor U2385 (N_2385,N_1174,N_62);
and U2386 (N_2386,N_127,N_284);
nor U2387 (N_2387,N_73,N_289);
and U2388 (N_2388,N_129,N_470);
or U2389 (N_2389,N_1062,N_784);
and U2390 (N_2390,N_868,N_659);
nor U2391 (N_2391,N_933,N_912);
or U2392 (N_2392,N_220,N_420);
xnor U2393 (N_2393,N_87,N_973);
nand U2394 (N_2394,N_422,N_1128);
and U2395 (N_2395,N_599,N_630);
or U2396 (N_2396,N_572,N_375);
nor U2397 (N_2397,N_846,N_1002);
and U2398 (N_2398,N_161,N_1099);
and U2399 (N_2399,N_1145,N_547);
or U2400 (N_2400,N_563,N_313);
or U2401 (N_2401,N_301,N_1224);
nand U2402 (N_2402,N_407,N_493);
or U2403 (N_2403,N_767,N_986);
nor U2404 (N_2404,N_1094,N_1168);
xnor U2405 (N_2405,N_217,N_762);
and U2406 (N_2406,N_1206,N_219);
nand U2407 (N_2407,N_1072,N_42);
nor U2408 (N_2408,N_984,N_404);
or U2409 (N_2409,N_281,N_983);
nor U2410 (N_2410,N_214,N_1055);
nand U2411 (N_2411,N_525,N_229);
and U2412 (N_2412,N_396,N_597);
or U2413 (N_2413,N_90,N_601);
or U2414 (N_2414,N_180,N_1006);
and U2415 (N_2415,N_1007,N_22);
nand U2416 (N_2416,N_210,N_79);
nand U2417 (N_2417,N_537,N_504);
nand U2418 (N_2418,N_820,N_355);
xnor U2419 (N_2419,N_187,N_658);
nand U2420 (N_2420,N_236,N_623);
or U2421 (N_2421,N_1099,N_589);
nor U2422 (N_2422,N_725,N_225);
and U2423 (N_2423,N_208,N_607);
nor U2424 (N_2424,N_230,N_329);
nor U2425 (N_2425,N_884,N_299);
or U2426 (N_2426,N_640,N_901);
or U2427 (N_2427,N_732,N_255);
nand U2428 (N_2428,N_58,N_199);
and U2429 (N_2429,N_999,N_340);
and U2430 (N_2430,N_117,N_127);
nand U2431 (N_2431,N_326,N_948);
and U2432 (N_2432,N_442,N_404);
xor U2433 (N_2433,N_232,N_975);
or U2434 (N_2434,N_383,N_1141);
and U2435 (N_2435,N_210,N_1058);
nor U2436 (N_2436,N_289,N_213);
and U2437 (N_2437,N_457,N_816);
and U2438 (N_2438,N_383,N_221);
and U2439 (N_2439,N_466,N_367);
and U2440 (N_2440,N_1067,N_641);
and U2441 (N_2441,N_420,N_522);
or U2442 (N_2442,N_340,N_178);
xnor U2443 (N_2443,N_210,N_554);
nor U2444 (N_2444,N_507,N_1108);
xnor U2445 (N_2445,N_294,N_15);
nand U2446 (N_2446,N_924,N_425);
nand U2447 (N_2447,N_35,N_281);
nand U2448 (N_2448,N_1035,N_111);
or U2449 (N_2449,N_1105,N_1012);
nor U2450 (N_2450,N_376,N_953);
or U2451 (N_2451,N_38,N_143);
xor U2452 (N_2452,N_267,N_1031);
nand U2453 (N_2453,N_386,N_546);
xnor U2454 (N_2454,N_242,N_199);
or U2455 (N_2455,N_406,N_995);
nor U2456 (N_2456,N_1083,N_441);
and U2457 (N_2457,N_799,N_8);
or U2458 (N_2458,N_521,N_1214);
xnor U2459 (N_2459,N_1127,N_2);
and U2460 (N_2460,N_800,N_1160);
xor U2461 (N_2461,N_399,N_157);
or U2462 (N_2462,N_284,N_725);
nor U2463 (N_2463,N_815,N_635);
and U2464 (N_2464,N_136,N_611);
nand U2465 (N_2465,N_502,N_678);
xnor U2466 (N_2466,N_994,N_905);
or U2467 (N_2467,N_253,N_355);
xnor U2468 (N_2468,N_604,N_321);
xor U2469 (N_2469,N_406,N_824);
nor U2470 (N_2470,N_292,N_680);
or U2471 (N_2471,N_1102,N_247);
or U2472 (N_2472,N_925,N_1166);
or U2473 (N_2473,N_262,N_1140);
nor U2474 (N_2474,N_187,N_813);
or U2475 (N_2475,N_848,N_349);
or U2476 (N_2476,N_1128,N_59);
or U2477 (N_2477,N_852,N_786);
and U2478 (N_2478,N_865,N_66);
xor U2479 (N_2479,N_207,N_966);
and U2480 (N_2480,N_1078,N_19);
nand U2481 (N_2481,N_799,N_591);
nor U2482 (N_2482,N_958,N_562);
and U2483 (N_2483,N_874,N_28);
and U2484 (N_2484,N_1076,N_968);
nor U2485 (N_2485,N_234,N_505);
or U2486 (N_2486,N_1021,N_670);
xor U2487 (N_2487,N_196,N_1056);
nand U2488 (N_2488,N_97,N_982);
xor U2489 (N_2489,N_506,N_333);
nand U2490 (N_2490,N_649,N_711);
and U2491 (N_2491,N_473,N_724);
nand U2492 (N_2492,N_366,N_1075);
nor U2493 (N_2493,N_249,N_114);
nand U2494 (N_2494,N_56,N_944);
nand U2495 (N_2495,N_1182,N_357);
xnor U2496 (N_2496,N_522,N_491);
nor U2497 (N_2497,N_78,N_2);
nand U2498 (N_2498,N_1125,N_760);
xor U2499 (N_2499,N_81,N_1247);
and U2500 (N_2500,N_1540,N_1414);
and U2501 (N_2501,N_1738,N_1301);
xor U2502 (N_2502,N_2208,N_1591);
xnor U2503 (N_2503,N_2147,N_2296);
nor U2504 (N_2504,N_1658,N_1914);
and U2505 (N_2505,N_1880,N_2131);
nor U2506 (N_2506,N_1382,N_1327);
and U2507 (N_2507,N_1742,N_1948);
nand U2508 (N_2508,N_1273,N_2070);
and U2509 (N_2509,N_2285,N_2057);
or U2510 (N_2510,N_1443,N_2157);
nand U2511 (N_2511,N_1719,N_1830);
and U2512 (N_2512,N_1457,N_1625);
nand U2513 (N_2513,N_1252,N_1816);
nand U2514 (N_2514,N_2238,N_1602);
nor U2515 (N_2515,N_2470,N_2217);
and U2516 (N_2516,N_1458,N_1665);
or U2517 (N_2517,N_2306,N_1812);
nand U2518 (N_2518,N_1551,N_1779);
or U2519 (N_2519,N_1419,N_1297);
nor U2520 (N_2520,N_1901,N_1935);
nor U2521 (N_2521,N_2165,N_1426);
and U2522 (N_2522,N_2192,N_1789);
and U2523 (N_2523,N_2483,N_1579);
xnor U2524 (N_2524,N_2485,N_2198);
or U2525 (N_2525,N_2413,N_1436);
nor U2526 (N_2526,N_2126,N_1933);
nand U2527 (N_2527,N_2447,N_1520);
or U2528 (N_2528,N_2293,N_1349);
and U2529 (N_2529,N_2499,N_1384);
nand U2530 (N_2530,N_1438,N_2088);
and U2531 (N_2531,N_2325,N_1596);
and U2532 (N_2532,N_2497,N_1287);
nor U2533 (N_2533,N_2249,N_2024);
and U2534 (N_2534,N_2009,N_1844);
nor U2535 (N_2535,N_1839,N_2402);
nand U2536 (N_2536,N_2049,N_1931);
xnor U2537 (N_2537,N_2031,N_2185);
or U2538 (N_2538,N_1451,N_2167);
nor U2539 (N_2539,N_2168,N_1755);
nor U2540 (N_2540,N_1546,N_1364);
xnor U2541 (N_2541,N_1942,N_2032);
nand U2542 (N_2542,N_2055,N_2001);
xnor U2543 (N_2543,N_1547,N_1855);
or U2544 (N_2544,N_2098,N_1759);
xor U2545 (N_2545,N_1999,N_2458);
nand U2546 (N_2546,N_1652,N_2297);
xor U2547 (N_2547,N_1886,N_2415);
nor U2548 (N_2548,N_2466,N_1424);
or U2549 (N_2549,N_2344,N_2125);
nand U2550 (N_2550,N_1572,N_1396);
or U2551 (N_2551,N_1597,N_1638);
or U2552 (N_2552,N_1308,N_1867);
nand U2553 (N_2553,N_1295,N_2028);
xnor U2554 (N_2554,N_2003,N_2498);
and U2555 (N_2555,N_1427,N_2488);
nand U2556 (N_2556,N_1963,N_1869);
or U2557 (N_2557,N_2002,N_1410);
nand U2558 (N_2558,N_1666,N_2355);
nor U2559 (N_2559,N_1758,N_1422);
and U2560 (N_2560,N_1370,N_1537);
nand U2561 (N_2561,N_1473,N_1641);
and U2562 (N_2562,N_2013,N_1912);
xor U2563 (N_2563,N_1313,N_2120);
nand U2564 (N_2564,N_1987,N_1951);
and U2565 (N_2565,N_1745,N_1334);
or U2566 (N_2566,N_2023,N_2116);
nor U2567 (N_2567,N_1885,N_1762);
and U2568 (N_2568,N_2330,N_2036);
xnor U2569 (N_2569,N_1828,N_1944);
or U2570 (N_2570,N_2103,N_2428);
or U2571 (N_2571,N_2477,N_1896);
and U2572 (N_2572,N_1776,N_1329);
or U2573 (N_2573,N_1765,N_1791);
nand U2574 (N_2574,N_1592,N_2259);
and U2575 (N_2575,N_2121,N_1463);
nor U2576 (N_2576,N_1628,N_2457);
and U2577 (N_2577,N_2242,N_1324);
nor U2578 (N_2578,N_1395,N_1616);
or U2579 (N_2579,N_2341,N_1630);
nor U2580 (N_2580,N_2043,N_1411);
nand U2581 (N_2581,N_1345,N_2460);
or U2582 (N_2582,N_2310,N_2375);
nand U2583 (N_2583,N_2274,N_2058);
xor U2584 (N_2584,N_1864,N_2084);
nor U2585 (N_2585,N_2371,N_2317);
xor U2586 (N_2586,N_1826,N_2467);
and U2587 (N_2587,N_1900,N_1930);
xnor U2588 (N_2588,N_1744,N_1409);
nand U2589 (N_2589,N_1467,N_1711);
nand U2590 (N_2590,N_1518,N_2395);
and U2591 (N_2591,N_1918,N_2394);
or U2592 (N_2592,N_1437,N_2418);
xnor U2593 (N_2593,N_1967,N_1371);
or U2594 (N_2594,N_1674,N_1512);
and U2595 (N_2595,N_1965,N_1664);
or U2596 (N_2596,N_2450,N_2328);
xnor U2597 (N_2597,N_2454,N_2429);
and U2598 (N_2598,N_1388,N_2300);
nand U2599 (N_2599,N_2234,N_2456);
nor U2600 (N_2600,N_1307,N_2373);
or U2601 (N_2601,N_2484,N_1603);
xnor U2602 (N_2602,N_1815,N_2337);
and U2603 (N_2603,N_2236,N_1526);
nand U2604 (N_2604,N_1351,N_1701);
and U2605 (N_2605,N_1790,N_1848);
or U2606 (N_2606,N_1294,N_1585);
nor U2607 (N_2607,N_1906,N_1849);
and U2608 (N_2608,N_1763,N_1306);
nand U2609 (N_2609,N_1377,N_1574);
and U2610 (N_2610,N_2164,N_1890);
nand U2611 (N_2611,N_1584,N_1532);
nand U2612 (N_2612,N_2495,N_1651);
nor U2613 (N_2613,N_2348,N_2280);
or U2614 (N_2614,N_2246,N_1691);
or U2615 (N_2615,N_2307,N_2008);
nor U2616 (N_2616,N_2260,N_1996);
xor U2617 (N_2617,N_2427,N_2149);
nand U2618 (N_2618,N_1868,N_1398);
and U2619 (N_2619,N_2384,N_1983);
xnor U2620 (N_2620,N_2320,N_2374);
nand U2621 (N_2621,N_1977,N_2441);
nor U2622 (N_2622,N_1699,N_2091);
xnor U2623 (N_2623,N_1320,N_1391);
nand U2624 (N_2624,N_1562,N_1737);
or U2625 (N_2625,N_2151,N_1367);
nor U2626 (N_2626,N_1505,N_2482);
nand U2627 (N_2627,N_1400,N_1453);
xnor U2628 (N_2628,N_1749,N_1975);
nand U2629 (N_2629,N_1837,N_1279);
or U2630 (N_2630,N_1934,N_1966);
nor U2631 (N_2631,N_1843,N_1618);
nand U2632 (N_2632,N_1257,N_1973);
or U2633 (N_2633,N_2421,N_2301);
xnor U2634 (N_2634,N_1729,N_2468);
and U2635 (N_2635,N_2071,N_1293);
nand U2636 (N_2636,N_1978,N_1688);
nor U2637 (N_2637,N_2350,N_1800);
nand U2638 (N_2638,N_2132,N_1970);
nor U2639 (N_2639,N_1916,N_2107);
nor U2640 (N_2640,N_1560,N_2442);
nand U2641 (N_2641,N_2455,N_2490);
and U2642 (N_2642,N_1722,N_1379);
or U2643 (N_2643,N_2051,N_1797);
xor U2644 (N_2644,N_1622,N_2017);
nor U2645 (N_2645,N_2224,N_1363);
nor U2646 (N_2646,N_2291,N_1846);
and U2647 (N_2647,N_2085,N_2475);
nor U2648 (N_2648,N_1897,N_1700);
nor U2649 (N_2649,N_2273,N_2170);
and U2650 (N_2650,N_1444,N_1647);
and U2651 (N_2651,N_1835,N_1267);
or U2652 (N_2652,N_1642,N_2136);
or U2653 (N_2653,N_1459,N_2469);
and U2654 (N_2654,N_1998,N_1870);
nand U2655 (N_2655,N_1785,N_2389);
or U2656 (N_2656,N_1769,N_2119);
nor U2657 (N_2657,N_1863,N_2117);
or U2658 (N_2658,N_2445,N_1428);
and U2659 (N_2659,N_2409,N_2215);
or U2660 (N_2660,N_2486,N_1757);
nor U2661 (N_2661,N_1402,N_1736);
and U2662 (N_2662,N_1523,N_2183);
or U2663 (N_2663,N_1854,N_1552);
and U2664 (N_2664,N_1686,N_1620);
nor U2665 (N_2665,N_1281,N_2377);
and U2666 (N_2666,N_1872,N_2252);
nor U2667 (N_2667,N_2191,N_1381);
and U2668 (N_2668,N_1639,N_1475);
xor U2669 (N_2669,N_2053,N_1670);
or U2670 (N_2670,N_2451,N_2021);
nand U2671 (N_2671,N_2081,N_1932);
xnor U2672 (N_2672,N_2278,N_2175);
nand U2673 (N_2673,N_1360,N_1772);
nand U2674 (N_2674,N_1519,N_1393);
and U2675 (N_2675,N_1979,N_2263);
nand U2676 (N_2676,N_1764,N_1418);
xor U2677 (N_2677,N_2207,N_2265);
nor U2678 (N_2678,N_1578,N_1253);
nor U2679 (N_2679,N_1626,N_1332);
or U2680 (N_2680,N_1416,N_2063);
nor U2681 (N_2681,N_2166,N_1621);
or U2682 (N_2682,N_2290,N_2471);
and U2683 (N_2683,N_1817,N_2361);
nand U2684 (N_2684,N_1913,N_1530);
nand U2685 (N_2685,N_2171,N_1649);
or U2686 (N_2686,N_1866,N_2064);
nand U2687 (N_2687,N_2141,N_2476);
or U2688 (N_2688,N_2480,N_1731);
or U2689 (N_2689,N_1277,N_1365);
and U2690 (N_2690,N_1369,N_1623);
xor U2691 (N_2691,N_1950,N_1922);
nor U2692 (N_2692,N_1521,N_1671);
and U2693 (N_2693,N_2423,N_1629);
nand U2694 (N_2694,N_2050,N_2094);
xor U2695 (N_2695,N_2193,N_1412);
nor U2696 (N_2696,N_2379,N_2250);
or U2697 (N_2697,N_1811,N_2391);
nand U2698 (N_2698,N_1710,N_2133);
nand U2699 (N_2699,N_2177,N_2343);
nor U2700 (N_2700,N_1971,N_2027);
nand U2701 (N_2701,N_1268,N_2255);
or U2702 (N_2702,N_2010,N_2230);
nand U2703 (N_2703,N_1882,N_1305);
xnor U2704 (N_2704,N_2073,N_1448);
or U2705 (N_2705,N_1741,N_1425);
nor U2706 (N_2706,N_2083,N_2087);
and U2707 (N_2707,N_1838,N_1877);
xor U2708 (N_2708,N_1732,N_1894);
or U2709 (N_2709,N_2018,N_1392);
nand U2710 (N_2710,N_2179,N_1771);
nand U2711 (N_2711,N_1511,N_2294);
nand U2712 (N_2712,N_2172,N_1343);
and U2713 (N_2713,N_1794,N_1624);
nor U2714 (N_2714,N_1299,N_1468);
nand U2715 (N_2715,N_1946,N_1832);
or U2716 (N_2716,N_1804,N_2162);
nand U2717 (N_2717,N_1806,N_1290);
or U2718 (N_2718,N_1915,N_1827);
nand U2719 (N_2719,N_1285,N_1570);
xnor U2720 (N_2720,N_1743,N_1783);
or U2721 (N_2721,N_2268,N_1506);
xor U2722 (N_2722,N_1516,N_2438);
and U2723 (N_2723,N_1461,N_2491);
and U2724 (N_2724,N_1472,N_1819);
xnor U2725 (N_2725,N_1354,N_1452);
nand U2726 (N_2726,N_1366,N_2323);
nand U2727 (N_2727,N_2140,N_1420);
xnor U2728 (N_2728,N_2176,N_1362);
xor U2729 (N_2729,N_1545,N_1997);
nor U2730 (N_2730,N_1746,N_1407);
or U2731 (N_2731,N_2218,N_2440);
xnor U2732 (N_2732,N_1561,N_1397);
and U2733 (N_2733,N_1534,N_2315);
xnor U2734 (N_2734,N_1689,N_1445);
xor U2735 (N_2735,N_1300,N_2228);
xor U2736 (N_2736,N_2363,N_1254);
or U2737 (N_2737,N_1487,N_1539);
or U2738 (N_2738,N_1470,N_1627);
nand U2739 (N_2739,N_1928,N_2299);
or U2740 (N_2740,N_2349,N_1712);
nand U2741 (N_2741,N_2047,N_2453);
and U2742 (N_2742,N_1693,N_2335);
nor U2743 (N_2743,N_2181,N_2210);
or U2744 (N_2744,N_2241,N_2261);
xor U2745 (N_2745,N_1587,N_2331);
and U2746 (N_2746,N_2393,N_1605);
xor U2747 (N_2747,N_1822,N_1682);
nand U2748 (N_2748,N_2052,N_2005);
nand U2749 (N_2749,N_1964,N_1640);
nor U2750 (N_2750,N_2115,N_1271);
nand U2751 (N_2751,N_1613,N_2305);
and U2752 (N_2752,N_2340,N_1490);
xnor U2753 (N_2753,N_1735,N_1538);
or U2754 (N_2754,N_1535,N_2286);
or U2755 (N_2755,N_1713,N_1927);
and U2756 (N_2756,N_1333,N_2159);
nor U2757 (N_2757,N_1637,N_2396);
and U2758 (N_2758,N_1482,N_2308);
or U2759 (N_2759,N_2270,N_1566);
nand U2760 (N_2760,N_2101,N_1358);
nand U2761 (N_2761,N_1718,N_2096);
xor U2762 (N_2762,N_1588,N_1383);
and U2763 (N_2763,N_1992,N_1348);
nor U2764 (N_2764,N_1836,N_1795);
xnor U2765 (N_2765,N_1586,N_2046);
or U2766 (N_2766,N_2033,N_2435);
nand U2767 (N_2767,N_2358,N_1604);
nor U2768 (N_2768,N_2038,N_2045);
xnor U2769 (N_2769,N_1825,N_2245);
or U2770 (N_2770,N_2102,N_1251);
nand U2771 (N_2771,N_2411,N_2105);
or U2772 (N_2772,N_1694,N_1325);
or U2773 (N_2773,N_2016,N_2202);
xnor U2774 (N_2774,N_1801,N_2420);
nand U2775 (N_2775,N_2104,N_1903);
xnor U2776 (N_2776,N_1891,N_2206);
nand U2777 (N_2777,N_2266,N_1669);
or U2778 (N_2778,N_1346,N_1661);
xnor U2779 (N_2779,N_1960,N_1611);
nor U2780 (N_2780,N_2093,N_1884);
nor U2781 (N_2781,N_1947,N_2303);
or U2782 (N_2782,N_2431,N_2329);
xnor U2783 (N_2783,N_2370,N_1269);
xor U2784 (N_2784,N_2272,N_1646);
nand U2785 (N_2785,N_1980,N_2289);
xnor U2786 (N_2786,N_1726,N_1856);
xor U2787 (N_2787,N_1399,N_1595);
and U2788 (N_2788,N_2321,N_1949);
nor U2789 (N_2789,N_2231,N_1824);
nor U2790 (N_2790,N_1995,N_1565);
nand U2791 (N_2791,N_1401,N_2383);
and U2792 (N_2792,N_2425,N_2118);
nand U2793 (N_2793,N_2399,N_1808);
and U2794 (N_2794,N_1507,N_1953);
nand U2795 (N_2795,N_1703,N_1476);
or U2796 (N_2796,N_1421,N_2059);
nand U2797 (N_2797,N_2240,N_1697);
nor U2798 (N_2798,N_2302,N_1704);
and U2799 (N_2799,N_1974,N_2199);
nand U2800 (N_2800,N_1288,N_1527);
or U2801 (N_2801,N_1533,N_1727);
nor U2802 (N_2802,N_1413,N_1860);
or U2803 (N_2803,N_1865,N_1542);
nand U2804 (N_2804,N_1321,N_1357);
and U2805 (N_2805,N_1707,N_1728);
nor U2806 (N_2806,N_1986,N_2054);
or U2807 (N_2807,N_1594,N_1655);
and U2808 (N_2808,N_2180,N_1748);
xor U2809 (N_2809,N_1283,N_2424);
nand U2810 (N_2810,N_1972,N_1631);
nor U2811 (N_2811,N_2314,N_2353);
nor U2812 (N_2812,N_2067,N_1617);
nor U2813 (N_2813,N_1633,N_1676);
or U2814 (N_2814,N_1657,N_2026);
xor U2815 (N_2815,N_1715,N_2152);
nand U2816 (N_2816,N_1289,N_2042);
nand U2817 (N_2817,N_2444,N_1577);
and U2818 (N_2818,N_2360,N_1814);
xnor U2819 (N_2819,N_1368,N_1489);
or U2820 (N_2820,N_2127,N_2276);
and U2821 (N_2821,N_2022,N_2039);
xor U2822 (N_2822,N_2128,N_1553);
nor U2823 (N_2823,N_2462,N_2324);
nor U2824 (N_2824,N_1714,N_1644);
nor U2825 (N_2825,N_1575,N_1454);
xor U2826 (N_2826,N_2221,N_2367);
and U2827 (N_2827,N_2347,N_2474);
xnor U2828 (N_2828,N_2041,N_1667);
nand U2829 (N_2829,N_1840,N_1524);
xnor U2830 (N_2830,N_2075,N_1761);
and U2831 (N_2831,N_1705,N_2186);
nand U2832 (N_2832,N_1528,N_2015);
xnor U2833 (N_2833,N_1338,N_1834);
nor U2834 (N_2834,N_1990,N_1432);
and U2835 (N_2835,N_1494,N_2401);
or U2836 (N_2836,N_2122,N_1888);
xnor U2837 (N_2837,N_1310,N_1770);
and U2838 (N_2838,N_1282,N_1768);
and U2839 (N_2839,N_1925,N_1315);
nand U2840 (N_2840,N_1961,N_2311);
nand U2841 (N_2841,N_1612,N_1328);
and U2842 (N_2842,N_2214,N_1962);
nor U2843 (N_2843,N_1632,N_2376);
and U2844 (N_2844,N_2189,N_2106);
xnor U2845 (N_2845,N_2090,N_1635);
nand U2846 (N_2846,N_1350,N_2123);
or U2847 (N_2847,N_1514,N_1780);
or U2848 (N_2848,N_1417,N_1548);
xor U2849 (N_2849,N_1462,N_1439);
and U2850 (N_2850,N_1851,N_1721);
nand U2851 (N_2851,N_2086,N_2184);
xnor U2852 (N_2852,N_1389,N_2112);
or U2853 (N_2853,N_2196,N_1788);
nor U2854 (N_2854,N_2019,N_1309);
and U2855 (N_2855,N_1423,N_1430);
xor U2856 (N_2856,N_1879,N_1515);
nor U2857 (N_2857,N_1924,N_2212);
xnor U2858 (N_2858,N_2405,N_1390);
xnor U2859 (N_2859,N_1988,N_2173);
and U2860 (N_2860,N_1431,N_1576);
nand U2861 (N_2861,N_2351,N_2281);
nor U2862 (N_2862,N_1372,N_2235);
or U2863 (N_2863,N_1956,N_1564);
and U2864 (N_2864,N_1720,N_2044);
nor U2865 (N_2865,N_2333,N_1447);
and U2866 (N_2866,N_1280,N_1480);
nand U2867 (N_2867,N_1943,N_2388);
and U2868 (N_2868,N_1853,N_1276);
and U2869 (N_2869,N_1675,N_1292);
xor U2870 (N_2870,N_1660,N_2244);
and U2871 (N_2871,N_1650,N_2219);
or U2872 (N_2872,N_1483,N_2182);
or U2873 (N_2873,N_1919,N_2304);
and U2874 (N_2874,N_1460,N_1484);
or U2875 (N_2875,N_1902,N_2190);
nor U2876 (N_2876,N_2461,N_2188);
nand U2877 (N_2877,N_1581,N_2113);
or U2878 (N_2878,N_2146,N_2493);
nor U2879 (N_2879,N_1258,N_2412);
nor U2880 (N_2880,N_2381,N_1895);
nand U2881 (N_2881,N_1250,N_1857);
xnor U2882 (N_2882,N_2430,N_1598);
and U2883 (N_2883,N_1415,N_2326);
or U2884 (N_2884,N_1340,N_2327);
nand U2885 (N_2885,N_2264,N_1375);
and U2886 (N_2886,N_1861,N_2378);
and U2887 (N_2887,N_2439,N_2357);
nand U2888 (N_2888,N_1529,N_1493);
and U2889 (N_2889,N_1740,N_1643);
nor U2890 (N_2890,N_2034,N_2275);
nand U2891 (N_2891,N_2316,N_2161);
xnor U2892 (N_2892,N_2222,N_2097);
nand U2893 (N_2893,N_2257,N_1376);
xor U2894 (N_2894,N_1841,N_1708);
or U2895 (N_2895,N_1698,N_1898);
xnor U2896 (N_2896,N_2082,N_2332);
nor U2897 (N_2897,N_1993,N_1687);
nand U2898 (N_2898,N_1905,N_1497);
and U2899 (N_2899,N_2163,N_2248);
nand U2900 (N_2900,N_1751,N_2068);
nand U2901 (N_2901,N_1314,N_2233);
and U2902 (N_2902,N_2342,N_1272);
and U2903 (N_2903,N_1256,N_1823);
nand U2904 (N_2904,N_2200,N_2334);
or U2905 (N_2905,N_2220,N_2201);
nand U2906 (N_2906,N_1760,N_1766);
or U2907 (N_2907,N_1394,N_2322);
xnor U2908 (N_2908,N_1656,N_1829);
and U2909 (N_2909,N_2256,N_1873);
or U2910 (N_2910,N_1373,N_2400);
xor U2911 (N_2911,N_1673,N_1263);
nor U2912 (N_2912,N_1663,N_1734);
and U2913 (N_2913,N_2243,N_2473);
and U2914 (N_2914,N_1569,N_1648);
or U2915 (N_2915,N_1984,N_2029);
xor U2916 (N_2916,N_1502,N_2487);
or U2917 (N_2917,N_1668,N_2397);
and U2918 (N_2918,N_2143,N_2436);
and U2919 (N_2919,N_1752,N_1255);
nand U2920 (N_2920,N_2449,N_1481);
and U2921 (N_2921,N_1936,N_2359);
nand U2922 (N_2922,N_1404,N_1952);
nor U2923 (N_2923,N_1455,N_1387);
or U2924 (N_2924,N_1793,N_2492);
xnor U2925 (N_2925,N_2403,N_1347);
xor U2926 (N_2926,N_2432,N_1323);
xor U2927 (N_2927,N_1491,N_1336);
nand U2928 (N_2928,N_2336,N_2040);
and U2929 (N_2929,N_2066,N_1677);
xnor U2930 (N_2930,N_2223,N_1917);
or U2931 (N_2931,N_1270,N_1923);
xor U2932 (N_2932,N_2129,N_1680);
nor U2933 (N_2933,N_1355,N_1994);
and U2934 (N_2934,N_1469,N_1568);
or U2935 (N_2935,N_1920,N_2061);
nor U2936 (N_2936,N_2142,N_1503);
nor U2937 (N_2937,N_1260,N_2108);
and U2938 (N_2938,N_1774,N_1478);
nor U2939 (N_2939,N_1874,N_1938);
nand U2940 (N_2940,N_1796,N_1778);
xor U2941 (N_2941,N_2037,N_1842);
and U2942 (N_2942,N_2339,N_2446);
nand U2943 (N_2943,N_2416,N_1904);
and U2944 (N_2944,N_1887,N_2072);
xor U2945 (N_2945,N_1496,N_2144);
xor U2946 (N_2946,N_2417,N_2459);
and U2947 (N_2947,N_1702,N_2137);
or U2948 (N_2948,N_1831,N_2481);
or U2949 (N_2949,N_1802,N_1555);
or U2950 (N_2950,N_1302,N_1750);
and U2951 (N_2951,N_1821,N_1908);
and U2952 (N_2952,N_1549,N_1479);
and U2953 (N_2953,N_1787,N_2092);
nand U2954 (N_2954,N_2069,N_1352);
xor U2955 (N_2955,N_1264,N_2025);
xor U2956 (N_2956,N_1331,N_2392);
nor U2957 (N_2957,N_1809,N_2156);
or U2958 (N_2958,N_1777,N_2062);
and U2959 (N_2959,N_2489,N_1408);
and U2960 (N_2960,N_1775,N_2448);
or U2961 (N_2961,N_1807,N_1477);
or U2962 (N_2962,N_2150,N_1434);
or U2963 (N_2963,N_1982,N_1531);
xor U2964 (N_2964,N_1322,N_2312);
and U2965 (N_2965,N_2407,N_2213);
xor U2966 (N_2966,N_2443,N_2229);
xnor U2967 (N_2967,N_1653,N_2283);
xnor U2968 (N_2968,N_2203,N_2287);
xnor U2969 (N_2969,N_1724,N_1311);
nor U2970 (N_2970,N_2386,N_2267);
nor U2971 (N_2971,N_1405,N_1356);
xor U2972 (N_2972,N_1692,N_1261);
xor U2973 (N_2973,N_2362,N_1544);
and U2974 (N_2974,N_1850,N_1847);
or U2975 (N_2975,N_1683,N_1833);
xnor U2976 (N_2976,N_2089,N_1580);
nor U2977 (N_2977,N_1339,N_2295);
xor U2978 (N_2978,N_2030,N_1730);
nor U2979 (N_2979,N_1465,N_1403);
or U2980 (N_2980,N_2077,N_2111);
nor U2981 (N_2981,N_1563,N_2205);
or U2982 (N_2982,N_1558,N_1910);
nor U2983 (N_2983,N_1386,N_1509);
nand U2984 (N_2984,N_2318,N_2158);
or U2985 (N_2985,N_2465,N_2366);
xor U2986 (N_2986,N_1939,N_1504);
or U2987 (N_2987,N_1259,N_2434);
nor U2988 (N_2988,N_1679,N_1717);
or U2989 (N_2989,N_1862,N_1753);
nor U2990 (N_2990,N_1716,N_1706);
or U2991 (N_2991,N_1499,N_1298);
nor U2992 (N_2992,N_1940,N_1858);
xnor U2993 (N_2993,N_1685,N_1590);
nand U2994 (N_2994,N_1449,N_1926);
or U2995 (N_2995,N_2124,N_1291);
nand U2996 (N_2996,N_1275,N_1485);
nand U2997 (N_2997,N_2404,N_2364);
nand U2998 (N_2998,N_1456,N_1709);
and U2999 (N_2999,N_1344,N_2135);
or U3000 (N_3000,N_2309,N_1471);
nor U3001 (N_3001,N_2226,N_2284);
or U3002 (N_3002,N_1634,N_1601);
or U3003 (N_3003,N_1353,N_1303);
nor U3004 (N_3004,N_2109,N_1907);
xor U3005 (N_3005,N_1909,N_1464);
nand U3006 (N_3006,N_2437,N_1374);
nand U3007 (N_3007,N_2065,N_1792);
and U3008 (N_3008,N_1969,N_2368);
and U3009 (N_3009,N_2195,N_1337);
and U3010 (N_3010,N_1911,N_1747);
and U3011 (N_3011,N_1820,N_1296);
nand U3012 (N_3012,N_1892,N_1899);
xor U3013 (N_3013,N_2345,N_1341);
nor U3014 (N_3014,N_1889,N_2253);
and U3015 (N_3015,N_2433,N_2012);
xor U3016 (N_3016,N_2354,N_1610);
xor U3017 (N_3017,N_2074,N_2356);
xnor U3018 (N_3018,N_2398,N_1583);
nand U3019 (N_3019,N_1435,N_2076);
xor U3020 (N_3020,N_2372,N_1517);
xnor U3021 (N_3021,N_1662,N_2004);
nand U3022 (N_3022,N_1550,N_2365);
nor U3023 (N_3023,N_1522,N_2000);
or U3024 (N_3024,N_1607,N_2382);
nand U3025 (N_3025,N_2134,N_1262);
nor U3026 (N_3026,N_1818,N_2247);
or U3027 (N_3027,N_1782,N_1342);
or U3028 (N_3028,N_1845,N_1659);
or U3029 (N_3029,N_1989,N_1606);
nand U3030 (N_3030,N_1754,N_1695);
nand U3031 (N_3031,N_2478,N_1921);
xnor U3032 (N_3032,N_1361,N_2258);
xnor U3033 (N_3033,N_2239,N_2225);
and U3034 (N_3034,N_1474,N_1286);
nand U3035 (N_3035,N_1654,N_1559);
nor U3036 (N_3036,N_2035,N_1875);
nand U3037 (N_3037,N_1876,N_1543);
nand U3038 (N_3038,N_2204,N_1619);
xor U3039 (N_3039,N_2313,N_1739);
or U3040 (N_3040,N_1991,N_2078);
nor U3041 (N_3041,N_1798,N_2048);
or U3042 (N_3042,N_2155,N_2464);
xor U3043 (N_3043,N_1871,N_1859);
xnor U3044 (N_3044,N_1488,N_1466);
xnor U3045 (N_3045,N_2463,N_1330);
and U3046 (N_3046,N_2262,N_1881);
or U3047 (N_3047,N_2153,N_2352);
nor U3048 (N_3048,N_1805,N_1541);
and U3049 (N_3049,N_2232,N_2100);
and U3050 (N_3050,N_1557,N_1672);
xor U3051 (N_3051,N_1609,N_2479);
or U3052 (N_3052,N_1968,N_1599);
and U3053 (N_3053,N_2169,N_2410);
nor U3054 (N_3054,N_1945,N_2178);
xnor U3055 (N_3055,N_2406,N_1554);
and U3056 (N_3056,N_1513,N_1981);
nor U3057 (N_3057,N_1893,N_1786);
xor U3058 (N_3058,N_1385,N_2452);
and U3059 (N_3059,N_2279,N_1690);
and U3060 (N_3060,N_2227,N_2080);
nor U3061 (N_3061,N_1265,N_1536);
nand U3062 (N_3062,N_2319,N_2292);
xor U3063 (N_3063,N_2414,N_1510);
and U3064 (N_3064,N_1450,N_1937);
or U3065 (N_3065,N_2298,N_1852);
nor U3066 (N_3066,N_1976,N_1985);
nor U3067 (N_3067,N_2079,N_1941);
or U3068 (N_3068,N_2390,N_2197);
and U3069 (N_3069,N_1446,N_2237);
and U3070 (N_3070,N_2194,N_2422);
nor U3071 (N_3071,N_1442,N_1784);
nand U3072 (N_3072,N_2139,N_1615);
xnor U3073 (N_3073,N_2154,N_1756);
or U3074 (N_3074,N_1803,N_1957);
nor U3075 (N_3075,N_2472,N_1573);
or U3076 (N_3076,N_2254,N_2095);
nor U3077 (N_3077,N_2114,N_1378);
nor U3078 (N_3078,N_1318,N_1556);
nand U3079 (N_3079,N_1608,N_2014);
nand U3080 (N_3080,N_1878,N_1495);
nor U3081 (N_3081,N_1593,N_2174);
xor U3082 (N_3082,N_2007,N_1312);
nand U3083 (N_3083,N_1723,N_1684);
nor U3084 (N_3084,N_2211,N_2011);
xor U3085 (N_3085,N_1958,N_1929);
or U3086 (N_3086,N_1284,N_1955);
or U3087 (N_3087,N_1440,N_1406);
nand U3088 (N_3088,N_2346,N_2209);
xnor U3089 (N_3089,N_1600,N_2060);
nand U3090 (N_3090,N_2419,N_1429);
nor U3091 (N_3091,N_2148,N_2385);
nand U3092 (N_3092,N_2056,N_1498);
or U3093 (N_3093,N_2160,N_2187);
xor U3094 (N_3094,N_2251,N_2006);
xnor U3095 (N_3095,N_1767,N_1316);
nor U3096 (N_3096,N_2288,N_1678);
or U3097 (N_3097,N_1636,N_1589);
nor U3098 (N_3098,N_1266,N_1571);
and U3099 (N_3099,N_1380,N_1492);
xor U3100 (N_3100,N_2145,N_1508);
xor U3101 (N_3101,N_2496,N_1500);
or U3102 (N_3102,N_1696,N_1733);
or U3103 (N_3103,N_1326,N_1781);
or U3104 (N_3104,N_2282,N_2216);
and U3105 (N_3105,N_1725,N_1773);
and U3106 (N_3106,N_1799,N_2269);
and U3107 (N_3107,N_2387,N_2380);
and U3108 (N_3108,N_1501,N_1433);
and U3109 (N_3109,N_2130,N_1319);
nand U3110 (N_3110,N_1582,N_1359);
xor U3111 (N_3111,N_1810,N_1304);
nand U3112 (N_3112,N_2271,N_1813);
nor U3113 (N_3113,N_1278,N_2099);
nand U3114 (N_3114,N_2369,N_1525);
nor U3115 (N_3115,N_1954,N_1959);
and U3116 (N_3116,N_2494,N_2426);
nand U3117 (N_3117,N_1883,N_1567);
xor U3118 (N_3118,N_2110,N_1645);
nand U3119 (N_3119,N_2138,N_1317);
nand U3120 (N_3120,N_1681,N_1274);
and U3121 (N_3121,N_2408,N_2338);
nand U3122 (N_3122,N_1441,N_2020);
and U3123 (N_3123,N_1614,N_1335);
nor U3124 (N_3124,N_2277,N_1486);
or U3125 (N_3125,N_2330,N_1963);
and U3126 (N_3126,N_1337,N_2476);
xor U3127 (N_3127,N_1788,N_1534);
nor U3128 (N_3128,N_2459,N_1278);
xor U3129 (N_3129,N_1963,N_1808);
nand U3130 (N_3130,N_1802,N_2059);
or U3131 (N_3131,N_1585,N_1355);
nor U3132 (N_3132,N_2011,N_1522);
xor U3133 (N_3133,N_2430,N_2021);
and U3134 (N_3134,N_1799,N_2092);
or U3135 (N_3135,N_1977,N_1330);
nor U3136 (N_3136,N_1330,N_1352);
nand U3137 (N_3137,N_2171,N_1621);
nor U3138 (N_3138,N_2091,N_2336);
and U3139 (N_3139,N_2497,N_1508);
or U3140 (N_3140,N_2045,N_2128);
nand U3141 (N_3141,N_2255,N_1325);
and U3142 (N_3142,N_1325,N_1902);
and U3143 (N_3143,N_1836,N_1534);
and U3144 (N_3144,N_1754,N_1604);
nor U3145 (N_3145,N_2460,N_1270);
xnor U3146 (N_3146,N_1732,N_2039);
nor U3147 (N_3147,N_1482,N_1400);
and U3148 (N_3148,N_1740,N_1405);
and U3149 (N_3149,N_1547,N_1318);
nor U3150 (N_3150,N_2032,N_1690);
and U3151 (N_3151,N_2009,N_1752);
xor U3152 (N_3152,N_1530,N_1285);
xnor U3153 (N_3153,N_2160,N_2258);
nor U3154 (N_3154,N_2292,N_1464);
xnor U3155 (N_3155,N_2219,N_1842);
or U3156 (N_3156,N_1682,N_2040);
or U3157 (N_3157,N_1553,N_2351);
nor U3158 (N_3158,N_2359,N_1713);
nand U3159 (N_3159,N_1896,N_2437);
and U3160 (N_3160,N_2331,N_2160);
and U3161 (N_3161,N_2359,N_2066);
or U3162 (N_3162,N_1959,N_2190);
or U3163 (N_3163,N_2105,N_1969);
or U3164 (N_3164,N_1330,N_1481);
and U3165 (N_3165,N_2499,N_1785);
and U3166 (N_3166,N_2264,N_2276);
nand U3167 (N_3167,N_2398,N_1606);
xnor U3168 (N_3168,N_2114,N_2028);
or U3169 (N_3169,N_1555,N_2187);
and U3170 (N_3170,N_1402,N_2369);
and U3171 (N_3171,N_2098,N_2034);
xor U3172 (N_3172,N_2216,N_2215);
and U3173 (N_3173,N_2059,N_2275);
and U3174 (N_3174,N_2486,N_2482);
or U3175 (N_3175,N_2242,N_1642);
nor U3176 (N_3176,N_2446,N_1440);
and U3177 (N_3177,N_1942,N_1826);
nor U3178 (N_3178,N_1687,N_1592);
nand U3179 (N_3179,N_2467,N_2055);
nor U3180 (N_3180,N_1336,N_1526);
and U3181 (N_3181,N_2083,N_1279);
nor U3182 (N_3182,N_1371,N_1817);
nor U3183 (N_3183,N_2118,N_1823);
xnor U3184 (N_3184,N_2245,N_1941);
or U3185 (N_3185,N_1790,N_2264);
and U3186 (N_3186,N_1258,N_1382);
or U3187 (N_3187,N_1410,N_1786);
or U3188 (N_3188,N_1674,N_1957);
and U3189 (N_3189,N_1415,N_1279);
or U3190 (N_3190,N_1936,N_1285);
xor U3191 (N_3191,N_2290,N_1419);
nor U3192 (N_3192,N_2386,N_1580);
nor U3193 (N_3193,N_1981,N_1696);
nand U3194 (N_3194,N_2277,N_1997);
or U3195 (N_3195,N_1891,N_1440);
nor U3196 (N_3196,N_1453,N_2075);
and U3197 (N_3197,N_2268,N_2071);
nand U3198 (N_3198,N_1522,N_2117);
nor U3199 (N_3199,N_2069,N_2414);
nand U3200 (N_3200,N_1420,N_1870);
nor U3201 (N_3201,N_1408,N_1908);
or U3202 (N_3202,N_2107,N_2166);
xor U3203 (N_3203,N_2305,N_2365);
or U3204 (N_3204,N_1633,N_2215);
xor U3205 (N_3205,N_2347,N_1509);
xor U3206 (N_3206,N_1913,N_1386);
or U3207 (N_3207,N_1627,N_1659);
or U3208 (N_3208,N_1266,N_2482);
or U3209 (N_3209,N_2096,N_2353);
nand U3210 (N_3210,N_1374,N_2220);
or U3211 (N_3211,N_1583,N_1779);
and U3212 (N_3212,N_1395,N_2143);
or U3213 (N_3213,N_1862,N_2247);
xor U3214 (N_3214,N_1615,N_1535);
xor U3215 (N_3215,N_1747,N_2238);
or U3216 (N_3216,N_1930,N_1861);
or U3217 (N_3217,N_2174,N_2199);
and U3218 (N_3218,N_2197,N_1649);
and U3219 (N_3219,N_1774,N_1562);
and U3220 (N_3220,N_2445,N_2297);
nand U3221 (N_3221,N_2128,N_2459);
nand U3222 (N_3222,N_1973,N_1940);
xnor U3223 (N_3223,N_2126,N_2467);
and U3224 (N_3224,N_2239,N_2414);
or U3225 (N_3225,N_2260,N_1262);
or U3226 (N_3226,N_2139,N_2295);
xor U3227 (N_3227,N_2172,N_2470);
nand U3228 (N_3228,N_2214,N_1528);
or U3229 (N_3229,N_1789,N_2182);
nor U3230 (N_3230,N_2204,N_2209);
and U3231 (N_3231,N_1347,N_1548);
or U3232 (N_3232,N_2181,N_1931);
or U3233 (N_3233,N_2398,N_2074);
nor U3234 (N_3234,N_1410,N_1507);
xnor U3235 (N_3235,N_1283,N_1799);
or U3236 (N_3236,N_1930,N_1594);
nand U3237 (N_3237,N_1689,N_1949);
or U3238 (N_3238,N_1411,N_1360);
and U3239 (N_3239,N_2363,N_2055);
nand U3240 (N_3240,N_2239,N_2463);
and U3241 (N_3241,N_1307,N_1842);
xor U3242 (N_3242,N_2126,N_1490);
nor U3243 (N_3243,N_1392,N_1997);
or U3244 (N_3244,N_1944,N_2399);
xnor U3245 (N_3245,N_1941,N_2186);
or U3246 (N_3246,N_2497,N_1928);
or U3247 (N_3247,N_1871,N_1569);
and U3248 (N_3248,N_1803,N_1354);
nand U3249 (N_3249,N_2041,N_1499);
xor U3250 (N_3250,N_1565,N_1376);
xor U3251 (N_3251,N_1495,N_2171);
nor U3252 (N_3252,N_2042,N_1438);
nor U3253 (N_3253,N_1909,N_1337);
xnor U3254 (N_3254,N_1637,N_2460);
or U3255 (N_3255,N_2080,N_1645);
xnor U3256 (N_3256,N_1393,N_2162);
nand U3257 (N_3257,N_2336,N_1637);
xor U3258 (N_3258,N_1862,N_2438);
nand U3259 (N_3259,N_1856,N_1597);
nand U3260 (N_3260,N_1287,N_2473);
nand U3261 (N_3261,N_2065,N_2435);
nor U3262 (N_3262,N_2426,N_2062);
nor U3263 (N_3263,N_1837,N_1257);
and U3264 (N_3264,N_1966,N_1271);
xnor U3265 (N_3265,N_2061,N_1898);
nor U3266 (N_3266,N_1519,N_1425);
and U3267 (N_3267,N_1773,N_2433);
and U3268 (N_3268,N_2282,N_1275);
or U3269 (N_3269,N_1843,N_1464);
nor U3270 (N_3270,N_1510,N_1326);
or U3271 (N_3271,N_2002,N_1650);
nor U3272 (N_3272,N_2109,N_1507);
and U3273 (N_3273,N_1931,N_1841);
xor U3274 (N_3274,N_1289,N_1800);
or U3275 (N_3275,N_1923,N_1467);
or U3276 (N_3276,N_2311,N_1766);
and U3277 (N_3277,N_1878,N_1511);
nand U3278 (N_3278,N_2092,N_2340);
nand U3279 (N_3279,N_1811,N_1396);
xnor U3280 (N_3280,N_2221,N_1638);
xor U3281 (N_3281,N_1523,N_1270);
nand U3282 (N_3282,N_2313,N_2044);
nand U3283 (N_3283,N_1664,N_1462);
xor U3284 (N_3284,N_1390,N_1637);
and U3285 (N_3285,N_1870,N_2202);
nand U3286 (N_3286,N_1444,N_2357);
nor U3287 (N_3287,N_1648,N_1891);
or U3288 (N_3288,N_1749,N_1624);
nand U3289 (N_3289,N_1619,N_1527);
nor U3290 (N_3290,N_2438,N_1331);
xnor U3291 (N_3291,N_1738,N_2241);
nand U3292 (N_3292,N_1829,N_1361);
or U3293 (N_3293,N_1394,N_1324);
or U3294 (N_3294,N_1636,N_1783);
or U3295 (N_3295,N_1718,N_1308);
nor U3296 (N_3296,N_1262,N_2055);
or U3297 (N_3297,N_1542,N_1702);
nand U3298 (N_3298,N_2452,N_1871);
nand U3299 (N_3299,N_1339,N_2317);
xnor U3300 (N_3300,N_2167,N_2352);
or U3301 (N_3301,N_1897,N_2240);
and U3302 (N_3302,N_2419,N_1467);
or U3303 (N_3303,N_2057,N_1981);
xnor U3304 (N_3304,N_2341,N_1286);
xor U3305 (N_3305,N_1332,N_2011);
nand U3306 (N_3306,N_1913,N_2276);
and U3307 (N_3307,N_2030,N_2494);
nor U3308 (N_3308,N_2435,N_1846);
nand U3309 (N_3309,N_2104,N_1517);
or U3310 (N_3310,N_2493,N_2427);
and U3311 (N_3311,N_1976,N_2467);
and U3312 (N_3312,N_1683,N_1989);
nor U3313 (N_3313,N_2007,N_1869);
nor U3314 (N_3314,N_2167,N_1933);
nand U3315 (N_3315,N_1864,N_1808);
nor U3316 (N_3316,N_1775,N_1460);
or U3317 (N_3317,N_2423,N_2317);
xnor U3318 (N_3318,N_1966,N_2361);
xor U3319 (N_3319,N_2247,N_1747);
xnor U3320 (N_3320,N_1385,N_1466);
or U3321 (N_3321,N_1758,N_1989);
xnor U3322 (N_3322,N_1676,N_1938);
nand U3323 (N_3323,N_1834,N_1750);
and U3324 (N_3324,N_1293,N_1337);
and U3325 (N_3325,N_2061,N_1468);
and U3326 (N_3326,N_1547,N_2283);
nor U3327 (N_3327,N_2447,N_2386);
or U3328 (N_3328,N_2103,N_1451);
nand U3329 (N_3329,N_2377,N_1299);
or U3330 (N_3330,N_2049,N_2226);
and U3331 (N_3331,N_2237,N_2096);
nor U3332 (N_3332,N_1865,N_1918);
xor U3333 (N_3333,N_1870,N_1845);
nor U3334 (N_3334,N_2082,N_2439);
nor U3335 (N_3335,N_1283,N_2071);
xnor U3336 (N_3336,N_1749,N_1971);
nand U3337 (N_3337,N_1544,N_2011);
xor U3338 (N_3338,N_2410,N_1702);
nor U3339 (N_3339,N_1829,N_2013);
and U3340 (N_3340,N_1995,N_1253);
and U3341 (N_3341,N_1723,N_2124);
nand U3342 (N_3342,N_2278,N_1537);
nand U3343 (N_3343,N_1947,N_1391);
nor U3344 (N_3344,N_1464,N_2451);
nand U3345 (N_3345,N_2096,N_1846);
nor U3346 (N_3346,N_2340,N_1489);
nand U3347 (N_3347,N_1464,N_1371);
and U3348 (N_3348,N_2208,N_2034);
nand U3349 (N_3349,N_1877,N_1459);
and U3350 (N_3350,N_2330,N_2277);
nor U3351 (N_3351,N_1908,N_1495);
and U3352 (N_3352,N_2378,N_2129);
and U3353 (N_3353,N_2220,N_1876);
xor U3354 (N_3354,N_1477,N_2383);
nor U3355 (N_3355,N_2431,N_1770);
or U3356 (N_3356,N_1581,N_2488);
nand U3357 (N_3357,N_2489,N_2162);
nor U3358 (N_3358,N_2236,N_1656);
nor U3359 (N_3359,N_2332,N_1486);
xnor U3360 (N_3360,N_2243,N_1263);
and U3361 (N_3361,N_1394,N_1712);
nand U3362 (N_3362,N_2351,N_1875);
and U3363 (N_3363,N_1955,N_1921);
and U3364 (N_3364,N_1744,N_1607);
and U3365 (N_3365,N_1865,N_1590);
and U3366 (N_3366,N_2285,N_1927);
nor U3367 (N_3367,N_1462,N_2125);
and U3368 (N_3368,N_2237,N_1808);
nor U3369 (N_3369,N_2301,N_2235);
or U3370 (N_3370,N_2337,N_1255);
nor U3371 (N_3371,N_1836,N_1657);
nor U3372 (N_3372,N_2354,N_1622);
and U3373 (N_3373,N_2003,N_2298);
or U3374 (N_3374,N_1615,N_1789);
or U3375 (N_3375,N_2314,N_1986);
xor U3376 (N_3376,N_1678,N_2160);
or U3377 (N_3377,N_1340,N_2229);
or U3378 (N_3378,N_1346,N_1506);
nand U3379 (N_3379,N_2457,N_1861);
nor U3380 (N_3380,N_2380,N_2403);
and U3381 (N_3381,N_2043,N_2179);
and U3382 (N_3382,N_1296,N_2126);
nor U3383 (N_3383,N_2375,N_2074);
or U3384 (N_3384,N_2408,N_1495);
and U3385 (N_3385,N_1498,N_2268);
and U3386 (N_3386,N_1880,N_2481);
nor U3387 (N_3387,N_2256,N_1754);
and U3388 (N_3388,N_2340,N_2087);
nor U3389 (N_3389,N_1411,N_1604);
or U3390 (N_3390,N_2195,N_2254);
xnor U3391 (N_3391,N_2038,N_1984);
xor U3392 (N_3392,N_1886,N_1759);
nor U3393 (N_3393,N_2449,N_2320);
nand U3394 (N_3394,N_2444,N_2414);
or U3395 (N_3395,N_2282,N_2372);
nand U3396 (N_3396,N_1788,N_1908);
or U3397 (N_3397,N_1835,N_1302);
nand U3398 (N_3398,N_2299,N_2370);
and U3399 (N_3399,N_1925,N_1462);
nor U3400 (N_3400,N_1848,N_2267);
and U3401 (N_3401,N_2259,N_1689);
nor U3402 (N_3402,N_1502,N_2040);
nand U3403 (N_3403,N_1798,N_2120);
nand U3404 (N_3404,N_2442,N_2208);
and U3405 (N_3405,N_1370,N_2172);
or U3406 (N_3406,N_2140,N_2434);
nand U3407 (N_3407,N_2379,N_2066);
and U3408 (N_3408,N_1480,N_1590);
nor U3409 (N_3409,N_2325,N_2465);
nor U3410 (N_3410,N_2127,N_2348);
nand U3411 (N_3411,N_2419,N_1597);
and U3412 (N_3412,N_2095,N_1595);
xor U3413 (N_3413,N_2475,N_1912);
and U3414 (N_3414,N_1832,N_1943);
xnor U3415 (N_3415,N_1687,N_2200);
or U3416 (N_3416,N_1574,N_2238);
and U3417 (N_3417,N_2249,N_2124);
nor U3418 (N_3418,N_2178,N_1834);
nor U3419 (N_3419,N_2213,N_2140);
xnor U3420 (N_3420,N_2320,N_1829);
or U3421 (N_3421,N_1476,N_1897);
nor U3422 (N_3422,N_2497,N_1855);
and U3423 (N_3423,N_2462,N_1867);
and U3424 (N_3424,N_2039,N_2496);
and U3425 (N_3425,N_1985,N_1736);
nor U3426 (N_3426,N_2308,N_1355);
xnor U3427 (N_3427,N_2392,N_2202);
xnor U3428 (N_3428,N_1433,N_1376);
xnor U3429 (N_3429,N_1274,N_1420);
and U3430 (N_3430,N_1583,N_1942);
or U3431 (N_3431,N_2168,N_1770);
or U3432 (N_3432,N_1278,N_1515);
nor U3433 (N_3433,N_2063,N_2099);
and U3434 (N_3434,N_1667,N_1254);
or U3435 (N_3435,N_1782,N_2185);
nor U3436 (N_3436,N_2208,N_2358);
nor U3437 (N_3437,N_1985,N_2246);
nor U3438 (N_3438,N_1649,N_1793);
xor U3439 (N_3439,N_1525,N_1985);
nand U3440 (N_3440,N_2431,N_2334);
xor U3441 (N_3441,N_1295,N_1779);
and U3442 (N_3442,N_1805,N_1997);
nand U3443 (N_3443,N_1266,N_2135);
xnor U3444 (N_3444,N_1402,N_2446);
and U3445 (N_3445,N_2299,N_2261);
or U3446 (N_3446,N_2458,N_2258);
nand U3447 (N_3447,N_2287,N_2333);
nor U3448 (N_3448,N_2330,N_1950);
nand U3449 (N_3449,N_1632,N_2232);
nor U3450 (N_3450,N_2079,N_1833);
nand U3451 (N_3451,N_1523,N_1469);
xnor U3452 (N_3452,N_2420,N_2100);
or U3453 (N_3453,N_2195,N_2006);
and U3454 (N_3454,N_1562,N_1976);
or U3455 (N_3455,N_1891,N_2265);
or U3456 (N_3456,N_1686,N_1823);
nor U3457 (N_3457,N_1538,N_2105);
xor U3458 (N_3458,N_1336,N_1603);
nand U3459 (N_3459,N_2430,N_2040);
xor U3460 (N_3460,N_2246,N_2305);
nor U3461 (N_3461,N_1503,N_1860);
and U3462 (N_3462,N_2078,N_2401);
nand U3463 (N_3463,N_2221,N_1647);
or U3464 (N_3464,N_2107,N_1761);
or U3465 (N_3465,N_2074,N_1932);
or U3466 (N_3466,N_1996,N_1979);
nor U3467 (N_3467,N_1935,N_2340);
xnor U3468 (N_3468,N_1743,N_1364);
xnor U3469 (N_3469,N_1945,N_1703);
xor U3470 (N_3470,N_1827,N_1883);
or U3471 (N_3471,N_2351,N_2149);
nand U3472 (N_3472,N_1603,N_1920);
nor U3473 (N_3473,N_1583,N_2385);
xnor U3474 (N_3474,N_1368,N_2121);
nor U3475 (N_3475,N_1686,N_2291);
nand U3476 (N_3476,N_1671,N_1845);
or U3477 (N_3477,N_1536,N_2276);
and U3478 (N_3478,N_1978,N_1318);
nor U3479 (N_3479,N_1965,N_2302);
nor U3480 (N_3480,N_1915,N_2197);
xnor U3481 (N_3481,N_2326,N_1384);
xor U3482 (N_3482,N_2400,N_1265);
nand U3483 (N_3483,N_1393,N_1664);
and U3484 (N_3484,N_2461,N_2321);
nand U3485 (N_3485,N_1418,N_1839);
and U3486 (N_3486,N_1981,N_1321);
xor U3487 (N_3487,N_1492,N_2146);
nand U3488 (N_3488,N_1925,N_1425);
xor U3489 (N_3489,N_1344,N_1951);
and U3490 (N_3490,N_1658,N_2301);
xor U3491 (N_3491,N_1489,N_2224);
nand U3492 (N_3492,N_1354,N_2346);
or U3493 (N_3493,N_2215,N_1485);
nand U3494 (N_3494,N_2115,N_2326);
nor U3495 (N_3495,N_1352,N_2048);
or U3496 (N_3496,N_2369,N_1994);
and U3497 (N_3497,N_2129,N_2454);
xor U3498 (N_3498,N_1939,N_1882);
nor U3499 (N_3499,N_2396,N_2344);
and U3500 (N_3500,N_2283,N_1752);
nor U3501 (N_3501,N_2117,N_2076);
and U3502 (N_3502,N_1781,N_1414);
or U3503 (N_3503,N_2164,N_2466);
or U3504 (N_3504,N_2186,N_1784);
nor U3505 (N_3505,N_2231,N_1913);
or U3506 (N_3506,N_2464,N_2330);
nor U3507 (N_3507,N_2080,N_2435);
or U3508 (N_3508,N_1440,N_1768);
nor U3509 (N_3509,N_1394,N_1546);
xor U3510 (N_3510,N_2455,N_1945);
and U3511 (N_3511,N_1480,N_1364);
xor U3512 (N_3512,N_1495,N_1312);
nor U3513 (N_3513,N_1961,N_1755);
nand U3514 (N_3514,N_1664,N_2234);
or U3515 (N_3515,N_1327,N_1332);
nand U3516 (N_3516,N_1354,N_2051);
nor U3517 (N_3517,N_1505,N_2475);
and U3518 (N_3518,N_1444,N_2305);
and U3519 (N_3519,N_1489,N_1954);
and U3520 (N_3520,N_1752,N_1431);
or U3521 (N_3521,N_2070,N_2479);
nor U3522 (N_3522,N_1493,N_1787);
nor U3523 (N_3523,N_2229,N_2010);
nor U3524 (N_3524,N_1403,N_2330);
or U3525 (N_3525,N_1995,N_2205);
nor U3526 (N_3526,N_2340,N_2044);
xnor U3527 (N_3527,N_1408,N_2159);
xnor U3528 (N_3528,N_2330,N_1817);
nor U3529 (N_3529,N_2087,N_2305);
nor U3530 (N_3530,N_1377,N_1604);
xnor U3531 (N_3531,N_1740,N_1486);
xor U3532 (N_3532,N_1537,N_1671);
nand U3533 (N_3533,N_1925,N_1451);
xnor U3534 (N_3534,N_1592,N_2337);
nand U3535 (N_3535,N_1469,N_1518);
or U3536 (N_3536,N_2300,N_1304);
or U3537 (N_3537,N_2480,N_1356);
and U3538 (N_3538,N_2265,N_1652);
and U3539 (N_3539,N_1842,N_2163);
nor U3540 (N_3540,N_1458,N_2099);
nand U3541 (N_3541,N_2016,N_2449);
nor U3542 (N_3542,N_1533,N_1433);
and U3543 (N_3543,N_1425,N_1839);
or U3544 (N_3544,N_1956,N_1310);
nand U3545 (N_3545,N_1668,N_1447);
nor U3546 (N_3546,N_2132,N_1394);
nor U3547 (N_3547,N_2306,N_1331);
and U3548 (N_3548,N_1982,N_1588);
xnor U3549 (N_3549,N_1617,N_2357);
nor U3550 (N_3550,N_1973,N_1816);
or U3551 (N_3551,N_2034,N_2447);
xnor U3552 (N_3552,N_1653,N_2107);
nor U3553 (N_3553,N_1644,N_2301);
nor U3554 (N_3554,N_2216,N_2290);
and U3555 (N_3555,N_1682,N_2480);
nand U3556 (N_3556,N_1360,N_1340);
nor U3557 (N_3557,N_2135,N_1659);
or U3558 (N_3558,N_2035,N_1615);
nand U3559 (N_3559,N_1781,N_1906);
nand U3560 (N_3560,N_1657,N_1253);
nand U3561 (N_3561,N_2138,N_2279);
and U3562 (N_3562,N_1711,N_1726);
xor U3563 (N_3563,N_1608,N_2321);
xor U3564 (N_3564,N_2130,N_2059);
nand U3565 (N_3565,N_2298,N_2388);
nand U3566 (N_3566,N_2403,N_1468);
and U3567 (N_3567,N_1952,N_2294);
and U3568 (N_3568,N_1408,N_2152);
or U3569 (N_3569,N_2088,N_2007);
xnor U3570 (N_3570,N_1766,N_1279);
nand U3571 (N_3571,N_2281,N_2296);
or U3572 (N_3572,N_2076,N_2099);
xor U3573 (N_3573,N_1423,N_1878);
and U3574 (N_3574,N_1953,N_1840);
nor U3575 (N_3575,N_1931,N_2301);
or U3576 (N_3576,N_2019,N_1394);
xnor U3577 (N_3577,N_1850,N_2361);
nand U3578 (N_3578,N_1504,N_1833);
nand U3579 (N_3579,N_1821,N_1508);
nor U3580 (N_3580,N_2101,N_1993);
nand U3581 (N_3581,N_1497,N_2107);
and U3582 (N_3582,N_1526,N_1988);
nor U3583 (N_3583,N_1966,N_1889);
nor U3584 (N_3584,N_1448,N_1344);
xor U3585 (N_3585,N_1469,N_1951);
or U3586 (N_3586,N_1341,N_2036);
nand U3587 (N_3587,N_1541,N_1357);
nand U3588 (N_3588,N_1712,N_1722);
nand U3589 (N_3589,N_1880,N_2223);
and U3590 (N_3590,N_2019,N_1517);
xnor U3591 (N_3591,N_2191,N_1318);
xor U3592 (N_3592,N_1371,N_1882);
xnor U3593 (N_3593,N_2453,N_1325);
nor U3594 (N_3594,N_1640,N_1746);
nand U3595 (N_3595,N_2461,N_1677);
or U3596 (N_3596,N_1291,N_1802);
nor U3597 (N_3597,N_1514,N_1455);
and U3598 (N_3598,N_1257,N_1339);
and U3599 (N_3599,N_1508,N_2265);
nor U3600 (N_3600,N_1583,N_1313);
or U3601 (N_3601,N_1376,N_1538);
nand U3602 (N_3602,N_1308,N_1480);
or U3603 (N_3603,N_1746,N_1480);
nand U3604 (N_3604,N_2497,N_1846);
and U3605 (N_3605,N_1882,N_1575);
nor U3606 (N_3606,N_2059,N_1992);
nor U3607 (N_3607,N_2360,N_1571);
nand U3608 (N_3608,N_2292,N_1515);
nand U3609 (N_3609,N_1868,N_2059);
and U3610 (N_3610,N_1838,N_1514);
and U3611 (N_3611,N_1498,N_2295);
or U3612 (N_3612,N_1881,N_1831);
or U3613 (N_3613,N_2077,N_2381);
nor U3614 (N_3614,N_1705,N_1808);
nand U3615 (N_3615,N_2165,N_2266);
and U3616 (N_3616,N_1711,N_1980);
nand U3617 (N_3617,N_1542,N_1977);
nand U3618 (N_3618,N_2340,N_2339);
xor U3619 (N_3619,N_1946,N_1869);
nand U3620 (N_3620,N_1662,N_1757);
or U3621 (N_3621,N_1406,N_1801);
and U3622 (N_3622,N_2285,N_2404);
or U3623 (N_3623,N_1433,N_1803);
nand U3624 (N_3624,N_1362,N_1366);
nand U3625 (N_3625,N_2078,N_2479);
nand U3626 (N_3626,N_2343,N_2208);
nor U3627 (N_3627,N_1590,N_2404);
and U3628 (N_3628,N_2420,N_1429);
xor U3629 (N_3629,N_1762,N_2259);
and U3630 (N_3630,N_2028,N_1665);
nand U3631 (N_3631,N_1499,N_1275);
nor U3632 (N_3632,N_1936,N_1615);
and U3633 (N_3633,N_1726,N_1799);
nor U3634 (N_3634,N_1423,N_1879);
nand U3635 (N_3635,N_2434,N_1469);
nor U3636 (N_3636,N_1345,N_1482);
nor U3637 (N_3637,N_2069,N_2322);
nand U3638 (N_3638,N_2143,N_1302);
and U3639 (N_3639,N_2138,N_2010);
xnor U3640 (N_3640,N_2317,N_1369);
xnor U3641 (N_3641,N_1815,N_2083);
xor U3642 (N_3642,N_1960,N_2036);
nand U3643 (N_3643,N_1726,N_2357);
or U3644 (N_3644,N_1661,N_1602);
nand U3645 (N_3645,N_1423,N_1250);
nor U3646 (N_3646,N_2081,N_2066);
nand U3647 (N_3647,N_1966,N_1887);
and U3648 (N_3648,N_2444,N_2149);
nor U3649 (N_3649,N_2356,N_1373);
nor U3650 (N_3650,N_2270,N_1614);
nor U3651 (N_3651,N_1485,N_1447);
and U3652 (N_3652,N_2005,N_1819);
and U3653 (N_3653,N_2052,N_1698);
or U3654 (N_3654,N_1930,N_1395);
nor U3655 (N_3655,N_1457,N_2302);
nand U3656 (N_3656,N_1469,N_2098);
nand U3657 (N_3657,N_1693,N_2492);
xor U3658 (N_3658,N_1549,N_1814);
or U3659 (N_3659,N_1969,N_1925);
and U3660 (N_3660,N_1399,N_2096);
and U3661 (N_3661,N_2057,N_2275);
nor U3662 (N_3662,N_1715,N_1376);
nand U3663 (N_3663,N_1532,N_1707);
or U3664 (N_3664,N_2198,N_1377);
nand U3665 (N_3665,N_2250,N_1292);
and U3666 (N_3666,N_1620,N_2375);
xnor U3667 (N_3667,N_1820,N_1994);
nand U3668 (N_3668,N_1745,N_2303);
nor U3669 (N_3669,N_1382,N_1500);
nand U3670 (N_3670,N_2027,N_1639);
nand U3671 (N_3671,N_1622,N_2296);
or U3672 (N_3672,N_1412,N_1818);
xor U3673 (N_3673,N_2224,N_2128);
nor U3674 (N_3674,N_2297,N_1983);
xnor U3675 (N_3675,N_2133,N_1520);
xnor U3676 (N_3676,N_1848,N_2099);
nand U3677 (N_3677,N_2325,N_2370);
nand U3678 (N_3678,N_1882,N_2023);
or U3679 (N_3679,N_1632,N_1542);
and U3680 (N_3680,N_2248,N_1531);
nor U3681 (N_3681,N_1553,N_2174);
and U3682 (N_3682,N_1741,N_1598);
or U3683 (N_3683,N_1263,N_1311);
nand U3684 (N_3684,N_2025,N_1905);
nand U3685 (N_3685,N_1532,N_1893);
nand U3686 (N_3686,N_2295,N_2291);
xor U3687 (N_3687,N_1950,N_1663);
nor U3688 (N_3688,N_2060,N_1517);
and U3689 (N_3689,N_1557,N_1825);
nand U3690 (N_3690,N_1942,N_2493);
nor U3691 (N_3691,N_1929,N_1855);
nor U3692 (N_3692,N_1594,N_1760);
and U3693 (N_3693,N_1350,N_2353);
xnor U3694 (N_3694,N_1301,N_2370);
nor U3695 (N_3695,N_2354,N_1528);
xor U3696 (N_3696,N_1614,N_2213);
xnor U3697 (N_3697,N_1432,N_2115);
or U3698 (N_3698,N_2300,N_2014);
and U3699 (N_3699,N_1734,N_1789);
nor U3700 (N_3700,N_1372,N_1296);
nor U3701 (N_3701,N_1856,N_2499);
nor U3702 (N_3702,N_1388,N_1666);
xnor U3703 (N_3703,N_2495,N_1953);
nand U3704 (N_3704,N_1875,N_1559);
or U3705 (N_3705,N_1800,N_1494);
or U3706 (N_3706,N_2426,N_2385);
nor U3707 (N_3707,N_2019,N_1796);
or U3708 (N_3708,N_2115,N_2195);
nor U3709 (N_3709,N_1456,N_1916);
nand U3710 (N_3710,N_1950,N_2479);
and U3711 (N_3711,N_2363,N_1898);
and U3712 (N_3712,N_2378,N_2348);
xor U3713 (N_3713,N_1597,N_1561);
or U3714 (N_3714,N_1603,N_1787);
and U3715 (N_3715,N_2021,N_1625);
xnor U3716 (N_3716,N_1735,N_2213);
nand U3717 (N_3717,N_1698,N_1417);
nor U3718 (N_3718,N_1844,N_1556);
xor U3719 (N_3719,N_2338,N_1479);
or U3720 (N_3720,N_1303,N_1535);
or U3721 (N_3721,N_2357,N_2126);
and U3722 (N_3722,N_2082,N_2118);
xor U3723 (N_3723,N_2151,N_2275);
and U3724 (N_3724,N_2401,N_2127);
nor U3725 (N_3725,N_2359,N_1712);
nor U3726 (N_3726,N_2433,N_1718);
or U3727 (N_3727,N_1950,N_2354);
or U3728 (N_3728,N_1530,N_2419);
nand U3729 (N_3729,N_1789,N_1896);
and U3730 (N_3730,N_2005,N_1999);
xnor U3731 (N_3731,N_2450,N_2005);
and U3732 (N_3732,N_1664,N_1854);
xnor U3733 (N_3733,N_1295,N_1789);
nand U3734 (N_3734,N_2356,N_1870);
nand U3735 (N_3735,N_2069,N_1400);
and U3736 (N_3736,N_1589,N_2398);
nor U3737 (N_3737,N_2301,N_2420);
or U3738 (N_3738,N_2489,N_2436);
or U3739 (N_3739,N_1809,N_2223);
and U3740 (N_3740,N_2378,N_1533);
nor U3741 (N_3741,N_1928,N_2106);
and U3742 (N_3742,N_1428,N_2246);
nand U3743 (N_3743,N_2045,N_2003);
and U3744 (N_3744,N_2407,N_2048);
nor U3745 (N_3745,N_1804,N_1886);
or U3746 (N_3746,N_1550,N_1404);
and U3747 (N_3747,N_1921,N_1561);
nor U3748 (N_3748,N_2145,N_2308);
xnor U3749 (N_3749,N_1966,N_2172);
or U3750 (N_3750,N_2941,N_3351);
or U3751 (N_3751,N_3722,N_3720);
and U3752 (N_3752,N_2986,N_3008);
nand U3753 (N_3753,N_2922,N_2630);
nor U3754 (N_3754,N_3739,N_3118);
xnor U3755 (N_3755,N_3053,N_3184);
or U3756 (N_3756,N_3014,N_2844);
xor U3757 (N_3757,N_2567,N_2656);
nand U3758 (N_3758,N_3115,N_3627);
xnor U3759 (N_3759,N_3715,N_2849);
nand U3760 (N_3760,N_3382,N_3680);
or U3761 (N_3761,N_2625,N_2904);
or U3762 (N_3762,N_3272,N_3313);
or U3763 (N_3763,N_3349,N_3005);
nand U3764 (N_3764,N_3591,N_2639);
nand U3765 (N_3765,N_3575,N_2736);
and U3766 (N_3766,N_3708,N_3096);
nand U3767 (N_3767,N_3002,N_3617);
xnor U3768 (N_3768,N_3215,N_2704);
or U3769 (N_3769,N_3003,N_3194);
nand U3770 (N_3770,N_3078,N_3599);
or U3771 (N_3771,N_2501,N_3616);
and U3772 (N_3772,N_2506,N_2718);
nor U3773 (N_3773,N_2852,N_3332);
nor U3774 (N_3774,N_3701,N_3094);
and U3775 (N_3775,N_3516,N_3678);
or U3776 (N_3776,N_2798,N_2847);
nor U3777 (N_3777,N_2604,N_3267);
xor U3778 (N_3778,N_2944,N_3620);
nor U3779 (N_3779,N_3522,N_3592);
nor U3780 (N_3780,N_3360,N_3235);
xor U3781 (N_3781,N_2985,N_3697);
and U3782 (N_3782,N_3413,N_2565);
and U3783 (N_3783,N_2856,N_3232);
nand U3784 (N_3784,N_3135,N_3435);
nand U3785 (N_3785,N_3706,N_3363);
nand U3786 (N_3786,N_3148,N_3411);
xor U3787 (N_3787,N_2575,N_3454);
nor U3788 (N_3788,N_3379,N_2992);
or U3789 (N_3789,N_2942,N_2678);
xor U3790 (N_3790,N_3259,N_3529);
nor U3791 (N_3791,N_2843,N_3725);
or U3792 (N_3792,N_3694,N_3271);
nand U3793 (N_3793,N_3731,N_2806);
xnor U3794 (N_3794,N_3047,N_3388);
xnor U3795 (N_3795,N_2832,N_3227);
nand U3796 (N_3796,N_2618,N_2660);
or U3797 (N_3797,N_2668,N_3239);
nor U3798 (N_3798,N_3582,N_3427);
nor U3799 (N_3799,N_2608,N_3221);
nand U3800 (N_3800,N_2611,N_3415);
or U3801 (N_3801,N_3581,N_2773);
and U3802 (N_3802,N_2570,N_2616);
nand U3803 (N_3803,N_3493,N_3640);
xnor U3804 (N_3804,N_3525,N_2599);
xnor U3805 (N_3805,N_3317,N_2670);
nor U3806 (N_3806,N_3405,N_2958);
nand U3807 (N_3807,N_2631,N_3338);
nand U3808 (N_3808,N_3196,N_2830);
nor U3809 (N_3809,N_3636,N_2528);
xor U3810 (N_3810,N_3433,N_3623);
nand U3811 (N_3811,N_3646,N_3288);
nor U3812 (N_3812,N_2551,N_2790);
nor U3813 (N_3813,N_3690,N_2938);
nand U3814 (N_3814,N_3176,N_3450);
nor U3815 (N_3815,N_3074,N_2868);
and U3816 (N_3816,N_3589,N_2937);
or U3817 (N_3817,N_3459,N_2785);
or U3818 (N_3818,N_2640,N_2719);
and U3819 (N_3819,N_2580,N_3116);
nor U3820 (N_3820,N_3558,N_3654);
and U3821 (N_3821,N_3630,N_3736);
and U3822 (N_3822,N_3492,N_2762);
nand U3823 (N_3823,N_2726,N_3498);
and U3824 (N_3824,N_3426,N_2651);
or U3825 (N_3825,N_3605,N_3689);
xnor U3826 (N_3826,N_3716,N_3178);
nor U3827 (N_3827,N_2817,N_3126);
xnor U3828 (N_3828,N_3398,N_3536);
nor U3829 (N_3829,N_2896,N_3099);
or U3830 (N_3830,N_3579,N_3102);
nand U3831 (N_3831,N_3468,N_3628);
nand U3832 (N_3832,N_3298,N_3049);
nor U3833 (N_3833,N_2511,N_3161);
nand U3834 (N_3834,N_3286,N_3391);
xor U3835 (N_3835,N_2968,N_3670);
and U3836 (N_3836,N_2815,N_2867);
nand U3837 (N_3837,N_2561,N_3542);
and U3838 (N_3838,N_2783,N_3594);
nand U3839 (N_3839,N_3299,N_2840);
nand U3840 (N_3840,N_2556,N_3149);
and U3841 (N_3841,N_2666,N_2572);
xor U3842 (N_3842,N_2954,N_3384);
or U3843 (N_3843,N_3142,N_2715);
and U3844 (N_3844,N_3662,N_3367);
nor U3845 (N_3845,N_2881,N_3475);
nand U3846 (N_3846,N_3330,N_3552);
xor U3847 (N_3847,N_3671,N_3264);
and U3848 (N_3848,N_3257,N_3746);
xnor U3849 (N_3849,N_3738,N_3399);
or U3850 (N_3850,N_2716,N_2636);
or U3851 (N_3851,N_3369,N_3060);
nand U3852 (N_3852,N_3439,N_3103);
nand U3853 (N_3853,N_2516,N_3295);
and U3854 (N_3854,N_2967,N_2923);
and U3855 (N_3855,N_3396,N_3741);
nor U3856 (N_3856,N_3555,N_2831);
or U3857 (N_3857,N_2707,N_2703);
nor U3858 (N_3858,N_2796,N_2977);
nand U3859 (N_3859,N_2953,N_2804);
and U3860 (N_3860,N_2519,N_3704);
or U3861 (N_3861,N_3222,N_3310);
and U3862 (N_3862,N_2803,N_2858);
xnor U3863 (N_3863,N_3467,N_2998);
nand U3864 (N_3864,N_3560,N_2795);
nand U3865 (N_3865,N_3346,N_2892);
nand U3866 (N_3866,N_3596,N_3514);
nor U3867 (N_3867,N_3262,N_3693);
and U3868 (N_3868,N_3568,N_2589);
nand U3869 (N_3869,N_3425,N_3181);
nand U3870 (N_3870,N_2711,N_3269);
nand U3871 (N_3871,N_2690,N_2752);
and U3872 (N_3872,N_3653,N_3121);
and U3873 (N_3873,N_3124,N_2895);
xnor U3874 (N_3874,N_3389,N_2946);
nand U3875 (N_3875,N_3013,N_3160);
nor U3876 (N_3876,N_3319,N_3445);
nand U3877 (N_3877,N_3026,N_3559);
xnor U3878 (N_3878,N_2588,N_2526);
nor U3879 (N_3879,N_3155,N_3647);
and U3880 (N_3880,N_2842,N_2947);
xor U3881 (N_3881,N_2996,N_2983);
nand U3882 (N_3882,N_3683,N_3526);
or U3883 (N_3883,N_3104,N_2874);
and U3884 (N_3884,N_2687,N_2828);
and U3885 (N_3885,N_2808,N_3436);
xor U3886 (N_3886,N_3076,N_3110);
nand U3887 (N_3887,N_2869,N_2834);
nor U3888 (N_3888,N_2778,N_3420);
nor U3889 (N_3889,N_3549,N_3335);
nand U3890 (N_3890,N_2979,N_3331);
nand U3891 (N_3891,N_2697,N_2753);
xnor U3892 (N_3892,N_2652,N_2745);
nand U3893 (N_3893,N_3038,N_2779);
or U3894 (N_3894,N_3441,N_2851);
nand U3895 (N_3895,N_3687,N_2734);
xor U3896 (N_3896,N_3228,N_3661);
or U3897 (N_3897,N_3337,N_3077);
nand U3898 (N_3898,N_3659,N_3730);
nand U3899 (N_3899,N_3012,N_3528);
xnor U3900 (N_3900,N_2788,N_2601);
nor U3901 (N_3901,N_3655,N_2512);
or U3902 (N_3902,N_3125,N_3300);
nand U3903 (N_3903,N_2612,N_2786);
nand U3904 (N_3904,N_2645,N_3442);
nor U3905 (N_3905,N_3029,N_3376);
nand U3906 (N_3906,N_3209,N_3144);
nor U3907 (N_3907,N_2936,N_2929);
nand U3908 (N_3908,N_2820,N_3595);
and U3909 (N_3909,N_3684,N_3251);
nor U3910 (N_3910,N_3705,N_2861);
nand U3911 (N_3911,N_2665,N_3042);
or U3912 (N_3912,N_2981,N_2533);
xor U3913 (N_3913,N_3546,N_3487);
nor U3914 (N_3914,N_3089,N_2772);
and U3915 (N_3915,N_2702,N_3385);
or U3916 (N_3916,N_3061,N_3000);
nor U3917 (N_3917,N_3354,N_3258);
or U3918 (N_3918,N_2774,N_2603);
nand U3919 (N_3919,N_3580,N_3745);
or U3920 (N_3920,N_2579,N_3117);
nor U3921 (N_3921,N_3033,N_3747);
xor U3922 (N_3922,N_2883,N_2617);
xnor U3923 (N_3923,N_2569,N_2576);
nand U3924 (N_3924,N_3372,N_3368);
xor U3925 (N_3925,N_2595,N_3663);
nand U3926 (N_3926,N_3018,N_3151);
xnor U3927 (N_3927,N_2964,N_3688);
nor U3928 (N_3928,N_2848,N_3597);
nand U3929 (N_3929,N_3519,N_3179);
xor U3930 (N_3930,N_3073,N_3028);
xor U3931 (N_3931,N_3416,N_2724);
or U3932 (N_3932,N_3048,N_3022);
or U3933 (N_3933,N_2710,N_2807);
nand U3934 (N_3934,N_2673,N_3509);
nand U3935 (N_3935,N_2984,N_3123);
nand U3936 (N_3936,N_2628,N_2793);
nand U3937 (N_3937,N_2777,N_3211);
or U3938 (N_3938,N_3583,N_3213);
nor U3939 (N_3939,N_3248,N_2517);
and U3940 (N_3940,N_3703,N_3530);
nor U3941 (N_3941,N_3674,N_2521);
or U3942 (N_3942,N_3316,N_3034);
nor U3943 (N_3943,N_2523,N_3254);
and U3944 (N_3944,N_2691,N_3292);
nor U3945 (N_3945,N_2649,N_2700);
and U3946 (N_3946,N_2505,N_2963);
or U3947 (N_3947,N_3609,N_3234);
and U3948 (N_3948,N_3205,N_2717);
nand U3949 (N_3949,N_3285,N_2677);
xnor U3950 (N_3950,N_3284,N_3587);
and U3951 (N_3951,N_2880,N_2877);
and U3952 (N_3952,N_2835,N_3474);
nor U3953 (N_3953,N_3735,N_3280);
and U3954 (N_3954,N_2810,N_2747);
or U3955 (N_3955,N_2916,N_2699);
xnor U3956 (N_3956,N_3287,N_2590);
nor U3957 (N_3957,N_2841,N_2838);
and U3958 (N_3958,N_2764,N_2598);
nor U3959 (N_3959,N_3080,N_3187);
or U3960 (N_3960,N_3698,N_2761);
and U3961 (N_3961,N_2948,N_3208);
and U3962 (N_3962,N_2573,N_2749);
nor U3963 (N_3963,N_3195,N_2926);
or U3964 (N_3964,N_3244,N_3744);
nand U3965 (N_3965,N_3431,N_2875);
and U3966 (N_3966,N_3613,N_2889);
and U3967 (N_3967,N_3618,N_2574);
nor U3968 (N_3968,N_2729,N_3226);
and U3969 (N_3969,N_3365,N_3057);
or U3970 (N_3970,N_3165,N_3570);
xor U3971 (N_3971,N_2596,N_2766);
or U3972 (N_3972,N_3266,N_2776);
or U3973 (N_3973,N_3322,N_2814);
nor U3974 (N_3974,N_2741,N_2522);
xor U3975 (N_3975,N_2643,N_3036);
nor U3976 (N_3976,N_3109,N_2970);
nand U3977 (N_3977,N_2903,N_3107);
and U3978 (N_3978,N_2727,N_2988);
or U3979 (N_3979,N_3604,N_3069);
or U3980 (N_3980,N_3006,N_3629);
and U3981 (N_3981,N_3333,N_2581);
nand U3982 (N_3982,N_3001,N_3482);
nor U3983 (N_3983,N_3672,N_3634);
nor U3984 (N_3984,N_3488,N_2768);
xor U3985 (N_3985,N_3210,N_3650);
nand U3986 (N_3986,N_2965,N_3245);
xor U3987 (N_3987,N_3016,N_3146);
xor U3988 (N_3988,N_3041,N_3255);
nor U3989 (N_3989,N_3658,N_3410);
nand U3990 (N_3990,N_3071,N_3418);
xnor U3991 (N_3991,N_3397,N_3216);
nand U3992 (N_3992,N_3377,N_2756);
nand U3993 (N_3993,N_2547,N_2638);
and U3994 (N_3994,N_3289,N_3573);
and U3995 (N_3995,N_3302,N_2751);
xnor U3996 (N_3996,N_3510,N_3644);
nand U3997 (N_3997,N_3656,N_3572);
and U3998 (N_3998,N_3476,N_3557);
nor U3999 (N_3999,N_3461,N_3037);
nand U4000 (N_4000,N_3380,N_3409);
nand U4001 (N_4001,N_3748,N_2543);
and U4002 (N_4002,N_2921,N_2605);
xnor U4003 (N_4003,N_2646,N_2966);
and U4004 (N_4004,N_3406,N_3483);
and U4005 (N_4005,N_2560,N_3236);
or U4006 (N_4006,N_3578,N_3127);
xor U4007 (N_4007,N_2865,N_2924);
and U4008 (N_4008,N_3218,N_3277);
nand U4009 (N_4009,N_3502,N_3719);
nor U4010 (N_4010,N_2955,N_3352);
nand U4011 (N_4011,N_2683,N_2906);
and U4012 (N_4012,N_3050,N_3101);
nand U4013 (N_4013,N_2928,N_2976);
xor U4014 (N_4014,N_2959,N_3699);
and U4015 (N_4015,N_3565,N_3129);
and U4016 (N_4016,N_3009,N_2680);
or U4017 (N_4017,N_3742,N_3306);
and U4018 (N_4018,N_3532,N_3343);
nand U4019 (N_4019,N_3702,N_3374);
and U4020 (N_4020,N_3553,N_2635);
nor U4021 (N_4021,N_2733,N_3035);
nand U4022 (N_4022,N_2689,N_2546);
nor U4023 (N_4023,N_3717,N_3192);
and U4024 (N_4024,N_3220,N_3606);
or U4025 (N_4025,N_3154,N_3268);
nand U4026 (N_4026,N_2917,N_3438);
nand U4027 (N_4027,N_2593,N_3090);
nand U4028 (N_4028,N_3068,N_3669);
nand U4029 (N_4029,N_3347,N_2520);
xor U4030 (N_4030,N_3729,N_3190);
or U4031 (N_4031,N_2824,N_3443);
or U4032 (N_4032,N_3430,N_2909);
or U4033 (N_4033,N_3540,N_2813);
nor U4034 (N_4034,N_2913,N_3362);
or U4035 (N_4035,N_2943,N_3603);
or U4036 (N_4036,N_3726,N_3357);
nor U4037 (N_4037,N_2657,N_2633);
nand U4038 (N_4038,N_2969,N_3537);
nand U4039 (N_4039,N_3243,N_2587);
or U4040 (N_4040,N_3153,N_3469);
and U4041 (N_4041,N_3229,N_2620);
or U4042 (N_4042,N_2544,N_3095);
nor U4043 (N_4043,N_3639,N_2672);
and U4044 (N_4044,N_3711,N_3152);
nor U4045 (N_4045,N_2632,N_3324);
or U4046 (N_4046,N_3561,N_2582);
or U4047 (N_4047,N_3169,N_3189);
xor U4048 (N_4048,N_3489,N_3733);
nor U4049 (N_4049,N_3308,N_3204);
nor U4050 (N_4050,N_3700,N_3444);
or U4051 (N_4051,N_3247,N_2527);
and U4052 (N_4052,N_2583,N_3585);
or U4053 (N_4053,N_3366,N_3675);
nand U4054 (N_4054,N_3010,N_3025);
and U4055 (N_4055,N_3685,N_3651);
nor U4056 (N_4056,N_2585,N_3138);
xnor U4057 (N_4057,N_3100,N_2685);
xor U4058 (N_4058,N_2907,N_2952);
nor U4059 (N_4059,N_3088,N_3341);
xor U4060 (N_4060,N_2694,N_2562);
nor U4061 (N_4061,N_3633,N_2811);
nand U4062 (N_4062,N_2584,N_3166);
and U4063 (N_4063,N_2524,N_3682);
and U4064 (N_4064,N_2894,N_3665);
nor U4065 (N_4065,N_2782,N_2825);
and U4066 (N_4066,N_2648,N_3162);
nor U4067 (N_4067,N_3163,N_3242);
or U4068 (N_4068,N_3032,N_3350);
and U4069 (N_4069,N_2578,N_2600);
xnor U4070 (N_4070,N_2821,N_3424);
and U4071 (N_4071,N_3541,N_3608);
xor U4072 (N_4072,N_2586,N_3261);
nand U4073 (N_4073,N_2539,N_2708);
and U4074 (N_4074,N_2723,N_2541);
xnor U4075 (N_4075,N_2614,N_2644);
and U4076 (N_4076,N_2899,N_3020);
xor U4077 (N_4077,N_3311,N_3143);
nor U4078 (N_4078,N_3188,N_2681);
nor U4079 (N_4079,N_2664,N_3172);
nor U4080 (N_4080,N_2927,N_2552);
or U4081 (N_4081,N_3710,N_3323);
and U4082 (N_4082,N_3191,N_3206);
and U4083 (N_4083,N_2931,N_3743);
and U4084 (N_4084,N_2525,N_3707);
nor U4085 (N_4085,N_3563,N_2871);
or U4086 (N_4086,N_2770,N_2566);
nor U4087 (N_4087,N_2901,N_3063);
nand U4088 (N_4088,N_2994,N_3641);
nand U4089 (N_4089,N_3329,N_3457);
nand U4090 (N_4090,N_3574,N_2792);
nor U4091 (N_4091,N_3233,N_3404);
xor U4092 (N_4092,N_3512,N_3611);
and U4093 (N_4093,N_2900,N_3019);
nand U4094 (N_4094,N_3480,N_3390);
or U4095 (N_4095,N_3576,N_2767);
and U4096 (N_4096,N_2571,N_3186);
xnor U4097 (N_4097,N_3477,N_3249);
or U4098 (N_4098,N_3538,N_3217);
and U4099 (N_4099,N_3534,N_3447);
nand U4100 (N_4100,N_3645,N_3638);
or U4101 (N_4101,N_3676,N_2987);
nor U4102 (N_4102,N_2655,N_2930);
or U4103 (N_4103,N_3531,N_2623);
nand U4104 (N_4104,N_3626,N_3021);
nor U4105 (N_4105,N_3696,N_3031);
xor U4106 (N_4106,N_2549,N_2757);
and U4107 (N_4107,N_3307,N_2893);
nor U4108 (N_4108,N_3072,N_3494);
nand U4109 (N_4109,N_3275,N_3207);
xnor U4110 (N_4110,N_2925,N_3417);
xnor U4111 (N_4111,N_3648,N_2982);
nand U4112 (N_4112,N_3223,N_2692);
nor U4113 (N_4113,N_3724,N_2859);
xnor U4114 (N_4114,N_3133,N_2558);
and U4115 (N_4115,N_2740,N_2918);
or U4116 (N_4116,N_2701,N_3429);
nor U4117 (N_4117,N_3533,N_3296);
and U4118 (N_4118,N_3497,N_2529);
nor U4119 (N_4119,N_2554,N_3201);
and U4120 (N_4120,N_2728,N_3464);
nor U4121 (N_4121,N_3158,N_3523);
or U4122 (N_4122,N_2693,N_2744);
or U4123 (N_4123,N_3407,N_2746);
nand U4124 (N_4124,N_3359,N_2816);
or U4125 (N_4125,N_2837,N_2833);
and U4126 (N_4126,N_3513,N_3402);
nor U4127 (N_4127,N_2939,N_3607);
and U4128 (N_4128,N_3056,N_3139);
nor U4129 (N_4129,N_2667,N_2731);
or U4130 (N_4130,N_2679,N_3046);
and U4131 (N_4131,N_2940,N_2607);
xor U4132 (N_4132,N_3087,N_2675);
or U4133 (N_4133,N_3130,N_3219);
nor U4134 (N_4134,N_2932,N_2765);
xnor U4135 (N_4135,N_2577,N_3619);
xor U4136 (N_4136,N_2564,N_3471);
or U4137 (N_4137,N_2621,N_2502);
nor U4138 (N_4138,N_2999,N_3007);
and U4139 (N_4139,N_3569,N_3168);
or U4140 (N_4140,N_2863,N_2737);
and U4141 (N_4141,N_3419,N_2706);
or U4142 (N_4142,N_3577,N_2622);
nand U4143 (N_4143,N_2759,N_3486);
nor U4144 (N_4144,N_2763,N_3175);
nand U4145 (N_4145,N_3612,N_2642);
nor U4146 (N_4146,N_3150,N_2908);
nor U4147 (N_4147,N_3539,N_3455);
xnor U4148 (N_4148,N_3465,N_3470);
nor U4149 (N_4149,N_3673,N_3462);
or U4150 (N_4150,N_2972,N_3119);
or U4151 (N_4151,N_2771,N_3463);
nor U4152 (N_4152,N_2853,N_3017);
nor U4153 (N_4153,N_3253,N_2990);
nor U4154 (N_4154,N_3180,N_3432);
nor U4155 (N_4155,N_3473,N_3065);
xnor U4156 (N_4156,N_3624,N_3260);
xor U4157 (N_4157,N_3400,N_3423);
nor U4158 (N_4158,N_2548,N_2855);
and U4159 (N_4159,N_3543,N_2658);
and U4160 (N_4160,N_3097,N_2659);
nor U4161 (N_4161,N_2780,N_2873);
nor U4162 (N_4162,N_3734,N_2735);
or U4163 (N_4163,N_2615,N_3452);
and U4164 (N_4164,N_2854,N_2503);
nand U4165 (N_4165,N_2886,N_2870);
or U4166 (N_4166,N_3506,N_3305);
nor U4167 (N_4167,N_3664,N_2879);
nor U4168 (N_4168,N_2902,N_3600);
nand U4169 (N_4169,N_3145,N_3395);
or U4170 (N_4170,N_3082,N_3631);
xor U4171 (N_4171,N_3458,N_3108);
and U4172 (N_4172,N_3064,N_2713);
nand U4173 (N_4173,N_3503,N_3274);
and U4174 (N_4174,N_3182,N_3011);
and U4175 (N_4175,N_3668,N_2538);
or U4176 (N_4176,N_2975,N_3281);
and U4177 (N_4177,N_3045,N_2637);
xnor U4178 (N_4178,N_2755,N_2602);
nor U4179 (N_4179,N_2641,N_2629);
nor U4180 (N_4180,N_3713,N_3456);
nand U4181 (N_4181,N_3667,N_2836);
nor U4182 (N_4182,N_3590,N_3086);
or U4183 (N_4183,N_3290,N_3714);
nor U4184 (N_4184,N_2910,N_3584);
nand U4185 (N_4185,N_3136,N_3325);
nand U4186 (N_4186,N_2695,N_3067);
nor U4187 (N_4187,N_2957,N_2559);
or U4188 (N_4188,N_3601,N_3058);
or U4189 (N_4189,N_3098,N_2915);
and U4190 (N_4190,N_3054,N_3070);
nor U4191 (N_4191,N_2722,N_3387);
xnor U4192 (N_4192,N_3521,N_2542);
and U4193 (N_4193,N_3083,N_3052);
xnor U4194 (N_4194,N_3320,N_2920);
or U4195 (N_4195,N_2890,N_3203);
nor U4196 (N_4196,N_2775,N_3508);
and U4197 (N_4197,N_2897,N_2518);
nand U4198 (N_4198,N_3602,N_2878);
nand U4199 (N_4199,N_2748,N_3265);
nor U4200 (N_4200,N_2669,N_3283);
xnor U4201 (N_4201,N_3079,N_3712);
nor U4202 (N_4202,N_3282,N_3434);
xnor U4203 (N_4203,N_2557,N_2812);
nand U4204 (N_4204,N_3309,N_2933);
and U4205 (N_4205,N_3586,N_3453);
or U4206 (N_4206,N_3392,N_3515);
xnor U4207 (N_4207,N_2973,N_2784);
nor U4208 (N_4208,N_2545,N_3547);
nand U4209 (N_4209,N_3635,N_3460);
and U4210 (N_4210,N_2592,N_2978);
xnor U4211 (N_4211,N_3212,N_2536);
nor U4212 (N_4212,N_2619,N_3024);
nor U4213 (N_4213,N_3535,N_3496);
and U4214 (N_4214,N_3106,N_3159);
xnor U4215 (N_4215,N_3193,N_2725);
xor U4216 (N_4216,N_3484,N_2531);
nor U4217 (N_4217,N_2884,N_3749);
or U4218 (N_4218,N_3173,N_2787);
nand U4219 (N_4219,N_3240,N_2540);
and U4220 (N_4220,N_3170,N_3621);
xor U4221 (N_4221,N_2872,N_3263);
nor U4222 (N_4222,N_2991,N_3598);
nor U4223 (N_4223,N_2627,N_2857);
or U4224 (N_4224,N_2591,N_2654);
or U4225 (N_4225,N_3030,N_2597);
and U4226 (N_4226,N_2661,N_3566);
or U4227 (N_4227,N_2609,N_2534);
nand U4228 (N_4228,N_3686,N_3081);
nor U4229 (N_4229,N_3174,N_3564);
and U4230 (N_4230,N_2535,N_3383);
and U4231 (N_4231,N_3093,N_3214);
nand U4232 (N_4232,N_2989,N_2742);
or U4233 (N_4233,N_3241,N_3371);
nor U4234 (N_4234,N_2709,N_3556);
nand U4235 (N_4235,N_3625,N_2914);
xor U4236 (N_4236,N_3339,N_3643);
nand U4237 (N_4237,N_3622,N_3428);
nor U4238 (N_4238,N_3128,N_2739);
and U4239 (N_4239,N_3593,N_3167);
xnor U4240 (N_4240,N_3238,N_2882);
xnor U4241 (N_4241,N_3111,N_3520);
and U4242 (N_4242,N_3326,N_3479);
nor U4243 (N_4243,N_3615,N_3224);
nor U4244 (N_4244,N_3562,N_3481);
nor U4245 (N_4245,N_2532,N_2568);
nand U4246 (N_4246,N_2550,N_3527);
xnor U4247 (N_4247,N_3408,N_2885);
xor U4248 (N_4248,N_3185,N_3112);
or U4249 (N_4249,N_3164,N_3544);
nor U4250 (N_4250,N_2826,N_3403);
xnor U4251 (N_4251,N_3198,N_2945);
or U4252 (N_4252,N_3340,N_3375);
xnor U4253 (N_4253,N_2769,N_3373);
and U4254 (N_4254,N_3023,N_2705);
nor U4255 (N_4255,N_2995,N_2634);
nor U4256 (N_4256,N_3381,N_2606);
or U4257 (N_4257,N_2510,N_2721);
nor U4258 (N_4258,N_2822,N_3301);
nand U4259 (N_4259,N_3004,N_3059);
nand U4260 (N_4260,N_3062,N_2971);
xor U4261 (N_4261,N_2688,N_2730);
or U4262 (N_4262,N_3237,N_2760);
nor U4263 (N_4263,N_2980,N_2509);
or U4264 (N_4264,N_2513,N_3171);
or U4265 (N_4265,N_3681,N_2860);
or U4266 (N_4266,N_3472,N_2750);
or U4267 (N_4267,N_3276,N_2956);
or U4268 (N_4268,N_2912,N_3356);
and U4269 (N_4269,N_2686,N_3637);
xnor U4270 (N_4270,N_3131,N_3015);
nor U4271 (N_4271,N_3511,N_3140);
or U4272 (N_4272,N_2508,N_2818);
nor U4273 (N_4273,N_3437,N_3737);
nor U4274 (N_4274,N_3355,N_3666);
nor U4275 (N_4275,N_3353,N_3740);
and U4276 (N_4276,N_2537,N_3293);
and U4277 (N_4277,N_2866,N_2613);
or U4278 (N_4278,N_2684,N_3252);
or U4279 (N_4279,N_3679,N_2743);
nor U4280 (N_4280,N_2507,N_3394);
nand U4281 (N_4281,N_2960,N_2653);
nor U4282 (N_4282,N_3545,N_3345);
nand U4283 (N_4283,N_2738,N_3327);
and U4284 (N_4284,N_3315,N_2919);
nor U4285 (N_4285,N_2682,N_3386);
and U4286 (N_4286,N_2839,N_2650);
nor U4287 (N_4287,N_3304,N_3044);
and U4288 (N_4288,N_3055,N_2758);
xor U4289 (N_4289,N_3312,N_2802);
xor U4290 (N_4290,N_3156,N_3550);
nand U4291 (N_4291,N_3610,N_2962);
nand U4292 (N_4292,N_3027,N_3657);
xor U4293 (N_4293,N_2911,N_3449);
nor U4294 (N_4294,N_2809,N_3230);
xor U4295 (N_4295,N_2950,N_3183);
nor U4296 (N_4296,N_2898,N_3279);
nand U4297 (N_4297,N_3348,N_3401);
nand U4298 (N_4298,N_2732,N_3137);
or U4299 (N_4299,N_2876,N_2563);
nor U4300 (N_4300,N_3571,N_2626);
and U4301 (N_4301,N_3134,N_3336);
and U4302 (N_4302,N_3446,N_3490);
nor U4303 (N_4303,N_2845,N_2850);
xor U4304 (N_4304,N_3728,N_3051);
nor U4305 (N_4305,N_2714,N_2504);
xor U4306 (N_4306,N_3478,N_2997);
xnor U4307 (N_4307,N_3364,N_2676);
or U4308 (N_4308,N_3328,N_2951);
nand U4309 (N_4309,N_2797,N_2791);
nor U4310 (N_4310,N_2949,N_2905);
nand U4311 (N_4311,N_2829,N_2961);
nand U4312 (N_4312,N_3649,N_3414);
and U4313 (N_4313,N_3501,N_3554);
xnor U4314 (N_4314,N_2789,N_2624);
nand U4315 (N_4315,N_3358,N_2663);
xor U4316 (N_4316,N_2819,N_3695);
nand U4317 (N_4317,N_2500,N_2514);
and U4318 (N_4318,N_2800,N_3660);
nor U4319 (N_4319,N_3642,N_2674);
and U4320 (N_4320,N_3551,N_3040);
nand U4321 (N_4321,N_3157,N_3085);
xnor U4322 (N_4322,N_3200,N_2794);
or U4323 (N_4323,N_3303,N_3092);
or U4324 (N_4324,N_3451,N_3499);
nand U4325 (N_4325,N_2823,N_2671);
or U4326 (N_4326,N_3225,N_3114);
nand U4327 (N_4327,N_3177,N_2515);
nand U4328 (N_4328,N_3091,N_3485);
or U4329 (N_4329,N_3495,N_3256);
or U4330 (N_4330,N_3105,N_3440);
and U4331 (N_4331,N_3548,N_2698);
nand U4332 (N_4332,N_2610,N_2935);
and U4333 (N_4333,N_2934,N_3294);
nand U4334 (N_4334,N_2864,N_3122);
nand U4335 (N_4335,N_3334,N_2647);
xor U4336 (N_4336,N_3507,N_3517);
nor U4337 (N_4337,N_3147,N_3113);
or U4338 (N_4338,N_3588,N_3448);
or U4339 (N_4339,N_2720,N_3732);
nand U4340 (N_4340,N_2594,N_2887);
and U4341 (N_4341,N_3344,N_3692);
nand U4342 (N_4342,N_2827,N_3505);
and U4343 (N_4343,N_3297,N_3727);
xor U4344 (N_4344,N_2696,N_3342);
nor U4345 (N_4345,N_3066,N_2712);
and U4346 (N_4346,N_2974,N_3652);
nand U4347 (N_4347,N_3361,N_3421);
and U4348 (N_4348,N_3120,N_2530);
or U4349 (N_4349,N_3202,N_3567);
xnor U4350 (N_4350,N_2891,N_3321);
nand U4351 (N_4351,N_3466,N_3412);
nand U4352 (N_4352,N_3132,N_3197);
or U4353 (N_4353,N_3291,N_3518);
xor U4354 (N_4354,N_2846,N_3246);
xnor U4355 (N_4355,N_3084,N_2754);
or U4356 (N_4356,N_2993,N_2888);
xnor U4357 (N_4357,N_2662,N_3075);
nor U4358 (N_4358,N_3709,N_2801);
xnor U4359 (N_4359,N_3500,N_3677);
or U4360 (N_4360,N_3141,N_2799);
and U4361 (N_4361,N_2781,N_3504);
and U4362 (N_4362,N_3393,N_3718);
nand U4363 (N_4363,N_2805,N_3632);
and U4364 (N_4364,N_3721,N_3314);
xor U4365 (N_4365,N_3614,N_3199);
xnor U4366 (N_4366,N_3491,N_2555);
and U4367 (N_4367,N_3422,N_2553);
and U4368 (N_4368,N_3370,N_3039);
nor U4369 (N_4369,N_3250,N_3231);
and U4370 (N_4370,N_3378,N_2862);
or U4371 (N_4371,N_3318,N_3723);
or U4372 (N_4372,N_3270,N_3043);
xnor U4373 (N_4373,N_3691,N_3278);
xor U4374 (N_4374,N_3524,N_3273);
nand U4375 (N_4375,N_2743,N_2758);
or U4376 (N_4376,N_3734,N_3031);
xor U4377 (N_4377,N_3319,N_2834);
and U4378 (N_4378,N_2506,N_2954);
and U4379 (N_4379,N_2811,N_2875);
nor U4380 (N_4380,N_2845,N_2995);
xor U4381 (N_4381,N_3673,N_3459);
nand U4382 (N_4382,N_2992,N_3354);
nand U4383 (N_4383,N_3665,N_3511);
nand U4384 (N_4384,N_3420,N_2774);
nor U4385 (N_4385,N_3161,N_3086);
nor U4386 (N_4386,N_3426,N_3684);
nor U4387 (N_4387,N_3502,N_2693);
nor U4388 (N_4388,N_3310,N_3225);
nand U4389 (N_4389,N_2604,N_3399);
or U4390 (N_4390,N_2531,N_3394);
xor U4391 (N_4391,N_3557,N_3090);
and U4392 (N_4392,N_2581,N_3445);
or U4393 (N_4393,N_3137,N_3180);
nand U4394 (N_4394,N_2551,N_3272);
and U4395 (N_4395,N_3271,N_3007);
and U4396 (N_4396,N_2631,N_2714);
nand U4397 (N_4397,N_2722,N_3384);
or U4398 (N_4398,N_3020,N_2607);
and U4399 (N_4399,N_3321,N_3604);
or U4400 (N_4400,N_2962,N_2957);
nor U4401 (N_4401,N_3716,N_2513);
or U4402 (N_4402,N_3741,N_2898);
nand U4403 (N_4403,N_3737,N_3582);
and U4404 (N_4404,N_2601,N_2505);
xor U4405 (N_4405,N_2867,N_2695);
and U4406 (N_4406,N_2614,N_2995);
or U4407 (N_4407,N_3280,N_3198);
or U4408 (N_4408,N_3324,N_3120);
xor U4409 (N_4409,N_3719,N_3214);
nand U4410 (N_4410,N_2814,N_3683);
and U4411 (N_4411,N_3674,N_3516);
nand U4412 (N_4412,N_3219,N_3387);
nor U4413 (N_4413,N_3283,N_2795);
nor U4414 (N_4414,N_3427,N_3249);
xor U4415 (N_4415,N_3473,N_3458);
nor U4416 (N_4416,N_3115,N_3000);
xnor U4417 (N_4417,N_2761,N_2697);
and U4418 (N_4418,N_3221,N_2724);
xnor U4419 (N_4419,N_3166,N_3438);
nand U4420 (N_4420,N_2581,N_2940);
and U4421 (N_4421,N_3037,N_3023);
xor U4422 (N_4422,N_3242,N_3092);
xor U4423 (N_4423,N_3650,N_2988);
xor U4424 (N_4424,N_3013,N_2640);
xor U4425 (N_4425,N_3332,N_3546);
xnor U4426 (N_4426,N_3149,N_3473);
nor U4427 (N_4427,N_3300,N_2539);
xnor U4428 (N_4428,N_2828,N_3304);
and U4429 (N_4429,N_3610,N_3727);
nor U4430 (N_4430,N_2712,N_2897);
or U4431 (N_4431,N_3684,N_3413);
or U4432 (N_4432,N_2621,N_2864);
or U4433 (N_4433,N_2986,N_2950);
nand U4434 (N_4434,N_2703,N_3065);
nor U4435 (N_4435,N_2833,N_3323);
and U4436 (N_4436,N_3261,N_3070);
and U4437 (N_4437,N_3167,N_2685);
and U4438 (N_4438,N_3704,N_3571);
nor U4439 (N_4439,N_3038,N_2894);
xor U4440 (N_4440,N_2597,N_3719);
xnor U4441 (N_4441,N_3581,N_2929);
or U4442 (N_4442,N_3005,N_3272);
or U4443 (N_4443,N_2943,N_2561);
or U4444 (N_4444,N_3605,N_2548);
and U4445 (N_4445,N_2972,N_3699);
nor U4446 (N_4446,N_3073,N_3585);
or U4447 (N_4447,N_3107,N_3505);
nor U4448 (N_4448,N_3283,N_3598);
or U4449 (N_4449,N_2531,N_2941);
nand U4450 (N_4450,N_3111,N_2928);
or U4451 (N_4451,N_3385,N_3736);
nor U4452 (N_4452,N_3675,N_3534);
nor U4453 (N_4453,N_3105,N_3395);
xnor U4454 (N_4454,N_3618,N_2606);
nand U4455 (N_4455,N_2605,N_2903);
or U4456 (N_4456,N_3174,N_3040);
or U4457 (N_4457,N_3467,N_2539);
xnor U4458 (N_4458,N_3481,N_2930);
nand U4459 (N_4459,N_2589,N_3251);
nor U4460 (N_4460,N_2529,N_2606);
nand U4461 (N_4461,N_3570,N_3443);
or U4462 (N_4462,N_2569,N_3138);
or U4463 (N_4463,N_2768,N_3584);
or U4464 (N_4464,N_3172,N_3645);
xnor U4465 (N_4465,N_3441,N_3584);
nand U4466 (N_4466,N_2971,N_2621);
xnor U4467 (N_4467,N_3499,N_2915);
and U4468 (N_4468,N_2821,N_2878);
and U4469 (N_4469,N_3608,N_2504);
xnor U4470 (N_4470,N_3729,N_3475);
and U4471 (N_4471,N_2589,N_3085);
or U4472 (N_4472,N_2859,N_2943);
or U4473 (N_4473,N_2591,N_3447);
nand U4474 (N_4474,N_2674,N_3555);
nand U4475 (N_4475,N_3257,N_3723);
nand U4476 (N_4476,N_2746,N_2689);
or U4477 (N_4477,N_2679,N_3174);
nor U4478 (N_4478,N_3731,N_3482);
nand U4479 (N_4479,N_3360,N_3231);
or U4480 (N_4480,N_3103,N_3464);
xnor U4481 (N_4481,N_3571,N_2591);
or U4482 (N_4482,N_2523,N_2994);
and U4483 (N_4483,N_3068,N_3256);
and U4484 (N_4484,N_3364,N_3686);
nor U4485 (N_4485,N_2675,N_3184);
nand U4486 (N_4486,N_2967,N_3114);
or U4487 (N_4487,N_3005,N_3640);
nor U4488 (N_4488,N_3061,N_2600);
xor U4489 (N_4489,N_3656,N_3151);
nand U4490 (N_4490,N_3444,N_3262);
and U4491 (N_4491,N_2552,N_3039);
or U4492 (N_4492,N_2627,N_3387);
nand U4493 (N_4493,N_2504,N_3477);
and U4494 (N_4494,N_3653,N_3334);
or U4495 (N_4495,N_2821,N_2882);
nor U4496 (N_4496,N_3623,N_3594);
nand U4497 (N_4497,N_3046,N_3167);
xor U4498 (N_4498,N_3387,N_3473);
xnor U4499 (N_4499,N_2563,N_3465);
and U4500 (N_4500,N_2745,N_2505);
and U4501 (N_4501,N_3361,N_3118);
nor U4502 (N_4502,N_3411,N_2694);
nor U4503 (N_4503,N_3621,N_2545);
xnor U4504 (N_4504,N_2748,N_3744);
nor U4505 (N_4505,N_2805,N_2840);
nand U4506 (N_4506,N_3303,N_2581);
nor U4507 (N_4507,N_3639,N_3748);
and U4508 (N_4508,N_2918,N_2971);
nand U4509 (N_4509,N_3030,N_2922);
xor U4510 (N_4510,N_3259,N_3294);
nor U4511 (N_4511,N_3738,N_3267);
xor U4512 (N_4512,N_3297,N_2624);
and U4513 (N_4513,N_2586,N_3588);
nor U4514 (N_4514,N_3447,N_2644);
or U4515 (N_4515,N_2719,N_2608);
xnor U4516 (N_4516,N_2832,N_3489);
nor U4517 (N_4517,N_3374,N_3353);
xnor U4518 (N_4518,N_3452,N_3563);
nand U4519 (N_4519,N_3208,N_3484);
nand U4520 (N_4520,N_2640,N_2693);
and U4521 (N_4521,N_2600,N_3671);
and U4522 (N_4522,N_2816,N_3340);
or U4523 (N_4523,N_3403,N_3412);
nor U4524 (N_4524,N_2798,N_3366);
or U4525 (N_4525,N_3114,N_3495);
nor U4526 (N_4526,N_3057,N_3727);
nand U4527 (N_4527,N_3422,N_3198);
or U4528 (N_4528,N_2908,N_3065);
nand U4529 (N_4529,N_3141,N_3599);
nor U4530 (N_4530,N_2698,N_3059);
or U4531 (N_4531,N_3259,N_3585);
xor U4532 (N_4532,N_2739,N_2807);
nor U4533 (N_4533,N_3531,N_2948);
or U4534 (N_4534,N_2655,N_2808);
xnor U4535 (N_4535,N_3116,N_3416);
and U4536 (N_4536,N_3099,N_3529);
or U4537 (N_4537,N_3180,N_2543);
and U4538 (N_4538,N_3389,N_2753);
nand U4539 (N_4539,N_3485,N_2893);
nand U4540 (N_4540,N_2698,N_2887);
and U4541 (N_4541,N_2732,N_3481);
nand U4542 (N_4542,N_3502,N_3009);
or U4543 (N_4543,N_2868,N_3062);
or U4544 (N_4544,N_2884,N_2799);
nand U4545 (N_4545,N_3650,N_3703);
or U4546 (N_4546,N_3081,N_3163);
xnor U4547 (N_4547,N_3516,N_3702);
nand U4548 (N_4548,N_2767,N_2643);
nand U4549 (N_4549,N_3157,N_3091);
and U4550 (N_4550,N_3329,N_3014);
and U4551 (N_4551,N_2724,N_2746);
nand U4552 (N_4552,N_3007,N_3164);
nor U4553 (N_4553,N_2589,N_2899);
nand U4554 (N_4554,N_3373,N_3107);
or U4555 (N_4555,N_3076,N_2506);
nor U4556 (N_4556,N_2723,N_3242);
nor U4557 (N_4557,N_3327,N_2829);
or U4558 (N_4558,N_3653,N_3306);
nor U4559 (N_4559,N_3469,N_2783);
xnor U4560 (N_4560,N_2568,N_3239);
nand U4561 (N_4561,N_3245,N_2616);
nor U4562 (N_4562,N_2698,N_2833);
nor U4563 (N_4563,N_3747,N_3285);
and U4564 (N_4564,N_2898,N_3143);
xor U4565 (N_4565,N_3232,N_3339);
xor U4566 (N_4566,N_3122,N_3193);
nor U4567 (N_4567,N_3127,N_3429);
or U4568 (N_4568,N_3083,N_3491);
or U4569 (N_4569,N_3278,N_3736);
and U4570 (N_4570,N_3313,N_2790);
xor U4571 (N_4571,N_3586,N_3242);
or U4572 (N_4572,N_2625,N_2646);
xor U4573 (N_4573,N_2757,N_3578);
nand U4574 (N_4574,N_3688,N_3193);
or U4575 (N_4575,N_2748,N_3377);
or U4576 (N_4576,N_2590,N_3233);
nor U4577 (N_4577,N_3432,N_3553);
xnor U4578 (N_4578,N_2922,N_3456);
and U4579 (N_4579,N_3720,N_3053);
or U4580 (N_4580,N_3549,N_3443);
and U4581 (N_4581,N_3054,N_3581);
nor U4582 (N_4582,N_3384,N_3619);
xnor U4583 (N_4583,N_3176,N_3383);
xor U4584 (N_4584,N_2948,N_3194);
xor U4585 (N_4585,N_2947,N_3461);
nor U4586 (N_4586,N_3481,N_3070);
or U4587 (N_4587,N_3067,N_2649);
nor U4588 (N_4588,N_3671,N_2957);
nor U4589 (N_4589,N_3262,N_3079);
or U4590 (N_4590,N_3534,N_3066);
or U4591 (N_4591,N_3649,N_2824);
or U4592 (N_4592,N_3402,N_2696);
or U4593 (N_4593,N_2795,N_3212);
nor U4594 (N_4594,N_3230,N_3273);
nor U4595 (N_4595,N_3143,N_2652);
nor U4596 (N_4596,N_2697,N_3006);
or U4597 (N_4597,N_3562,N_3712);
or U4598 (N_4598,N_2925,N_2724);
nand U4599 (N_4599,N_2855,N_3094);
xnor U4600 (N_4600,N_2997,N_2747);
nand U4601 (N_4601,N_3540,N_2588);
nor U4602 (N_4602,N_3126,N_3666);
and U4603 (N_4603,N_3104,N_2912);
xor U4604 (N_4604,N_3430,N_2723);
nor U4605 (N_4605,N_3090,N_2873);
nor U4606 (N_4606,N_2587,N_2620);
or U4607 (N_4607,N_3165,N_2835);
xnor U4608 (N_4608,N_2549,N_3612);
or U4609 (N_4609,N_3343,N_3322);
or U4610 (N_4610,N_2674,N_2796);
and U4611 (N_4611,N_2656,N_2866);
and U4612 (N_4612,N_3454,N_3359);
and U4613 (N_4613,N_2658,N_3040);
nand U4614 (N_4614,N_3204,N_3190);
xor U4615 (N_4615,N_2761,N_2557);
xnor U4616 (N_4616,N_2631,N_3611);
and U4617 (N_4617,N_2663,N_3202);
and U4618 (N_4618,N_3533,N_3048);
or U4619 (N_4619,N_3599,N_2832);
or U4620 (N_4620,N_3110,N_3567);
nor U4621 (N_4621,N_2663,N_2887);
nand U4622 (N_4622,N_3732,N_2960);
and U4623 (N_4623,N_3637,N_3462);
nor U4624 (N_4624,N_3103,N_2891);
nor U4625 (N_4625,N_3175,N_3533);
nand U4626 (N_4626,N_2668,N_3173);
or U4627 (N_4627,N_2581,N_3137);
xor U4628 (N_4628,N_3264,N_3506);
nor U4629 (N_4629,N_3075,N_2648);
or U4630 (N_4630,N_3419,N_3681);
nand U4631 (N_4631,N_3230,N_2963);
or U4632 (N_4632,N_3352,N_3106);
and U4633 (N_4633,N_2769,N_2863);
nor U4634 (N_4634,N_2924,N_2921);
and U4635 (N_4635,N_2546,N_3404);
xnor U4636 (N_4636,N_3192,N_2986);
nor U4637 (N_4637,N_3623,N_3088);
nand U4638 (N_4638,N_3359,N_2835);
and U4639 (N_4639,N_2676,N_3570);
nand U4640 (N_4640,N_2716,N_3569);
xnor U4641 (N_4641,N_2672,N_3123);
nand U4642 (N_4642,N_3159,N_3003);
xnor U4643 (N_4643,N_3391,N_3528);
nand U4644 (N_4644,N_2619,N_2530);
nor U4645 (N_4645,N_3264,N_3551);
nor U4646 (N_4646,N_2574,N_3644);
and U4647 (N_4647,N_2605,N_2838);
and U4648 (N_4648,N_2701,N_3704);
nor U4649 (N_4649,N_3147,N_2773);
and U4650 (N_4650,N_3020,N_2862);
xor U4651 (N_4651,N_2675,N_2783);
nand U4652 (N_4652,N_2951,N_3298);
nor U4653 (N_4653,N_3030,N_3557);
xor U4654 (N_4654,N_2705,N_2911);
xor U4655 (N_4655,N_3568,N_2635);
nand U4656 (N_4656,N_3745,N_3256);
and U4657 (N_4657,N_2697,N_3193);
xnor U4658 (N_4658,N_3379,N_2657);
nand U4659 (N_4659,N_2807,N_3596);
xnor U4660 (N_4660,N_3142,N_2580);
nand U4661 (N_4661,N_2588,N_2927);
or U4662 (N_4662,N_3043,N_2657);
xnor U4663 (N_4663,N_3104,N_3345);
nor U4664 (N_4664,N_2562,N_3498);
nor U4665 (N_4665,N_3550,N_2865);
nor U4666 (N_4666,N_2617,N_2695);
or U4667 (N_4667,N_3250,N_3285);
xor U4668 (N_4668,N_2584,N_3498);
xnor U4669 (N_4669,N_2896,N_3043);
and U4670 (N_4670,N_3593,N_2871);
and U4671 (N_4671,N_2584,N_2917);
nand U4672 (N_4672,N_2743,N_3464);
and U4673 (N_4673,N_2813,N_2976);
and U4674 (N_4674,N_2955,N_3070);
nand U4675 (N_4675,N_3349,N_2655);
or U4676 (N_4676,N_2968,N_3357);
nand U4677 (N_4677,N_3653,N_2788);
nand U4678 (N_4678,N_2792,N_3630);
and U4679 (N_4679,N_3307,N_3659);
nor U4680 (N_4680,N_3553,N_3137);
and U4681 (N_4681,N_2545,N_3128);
nor U4682 (N_4682,N_3011,N_3575);
and U4683 (N_4683,N_2680,N_2915);
and U4684 (N_4684,N_3652,N_2992);
and U4685 (N_4685,N_3570,N_2536);
or U4686 (N_4686,N_2718,N_3594);
or U4687 (N_4687,N_2922,N_3557);
or U4688 (N_4688,N_2982,N_3403);
nor U4689 (N_4689,N_2921,N_3358);
or U4690 (N_4690,N_3159,N_2831);
nor U4691 (N_4691,N_3608,N_3047);
nand U4692 (N_4692,N_3029,N_3469);
nor U4693 (N_4693,N_3337,N_2603);
nand U4694 (N_4694,N_3430,N_3449);
xnor U4695 (N_4695,N_3093,N_2787);
nor U4696 (N_4696,N_2741,N_3048);
and U4697 (N_4697,N_3736,N_3342);
or U4698 (N_4698,N_3079,N_2782);
and U4699 (N_4699,N_3203,N_3343);
and U4700 (N_4700,N_2541,N_3333);
nor U4701 (N_4701,N_2680,N_2991);
and U4702 (N_4702,N_3261,N_2933);
nand U4703 (N_4703,N_3655,N_3001);
or U4704 (N_4704,N_2685,N_2732);
xor U4705 (N_4705,N_3139,N_3418);
xor U4706 (N_4706,N_3223,N_2582);
nand U4707 (N_4707,N_3699,N_3663);
xnor U4708 (N_4708,N_3557,N_2832);
xor U4709 (N_4709,N_2877,N_3282);
nand U4710 (N_4710,N_3611,N_3458);
xnor U4711 (N_4711,N_2722,N_2981);
nor U4712 (N_4712,N_2818,N_2806);
xnor U4713 (N_4713,N_2569,N_2809);
nor U4714 (N_4714,N_3064,N_3573);
xnor U4715 (N_4715,N_3412,N_3338);
nand U4716 (N_4716,N_2531,N_3440);
or U4717 (N_4717,N_2764,N_2950);
and U4718 (N_4718,N_3178,N_3383);
nor U4719 (N_4719,N_3008,N_2869);
or U4720 (N_4720,N_3158,N_2573);
xnor U4721 (N_4721,N_3631,N_3748);
xnor U4722 (N_4722,N_2999,N_2611);
or U4723 (N_4723,N_3143,N_2522);
or U4724 (N_4724,N_2714,N_3242);
and U4725 (N_4725,N_2644,N_3297);
xnor U4726 (N_4726,N_3603,N_2775);
or U4727 (N_4727,N_3082,N_2564);
nor U4728 (N_4728,N_3223,N_3032);
xnor U4729 (N_4729,N_3113,N_2732);
nor U4730 (N_4730,N_2503,N_3170);
or U4731 (N_4731,N_2748,N_2859);
xnor U4732 (N_4732,N_2983,N_2691);
xor U4733 (N_4733,N_3459,N_3245);
nand U4734 (N_4734,N_3105,N_3426);
and U4735 (N_4735,N_3453,N_2957);
nand U4736 (N_4736,N_2800,N_3213);
nor U4737 (N_4737,N_3538,N_3214);
nor U4738 (N_4738,N_3440,N_2864);
xor U4739 (N_4739,N_3259,N_3201);
or U4740 (N_4740,N_2655,N_3016);
nor U4741 (N_4741,N_2594,N_3281);
and U4742 (N_4742,N_2908,N_3100);
nand U4743 (N_4743,N_3305,N_3034);
and U4744 (N_4744,N_2624,N_3196);
and U4745 (N_4745,N_3312,N_3532);
nand U4746 (N_4746,N_2717,N_2569);
xor U4747 (N_4747,N_3173,N_3288);
or U4748 (N_4748,N_2656,N_3429);
and U4749 (N_4749,N_2696,N_3167);
and U4750 (N_4750,N_2985,N_3527);
xnor U4751 (N_4751,N_3412,N_3175);
xnor U4752 (N_4752,N_3125,N_2694);
or U4753 (N_4753,N_3060,N_2524);
nand U4754 (N_4754,N_3533,N_2817);
nand U4755 (N_4755,N_2729,N_2555);
or U4756 (N_4756,N_3598,N_3137);
and U4757 (N_4757,N_3523,N_3030);
or U4758 (N_4758,N_3537,N_2933);
xnor U4759 (N_4759,N_3198,N_3072);
nand U4760 (N_4760,N_2845,N_2505);
or U4761 (N_4761,N_3291,N_3513);
and U4762 (N_4762,N_3139,N_2524);
and U4763 (N_4763,N_3102,N_2909);
nand U4764 (N_4764,N_3190,N_2975);
and U4765 (N_4765,N_3608,N_3075);
or U4766 (N_4766,N_3016,N_3331);
and U4767 (N_4767,N_3703,N_2654);
xnor U4768 (N_4768,N_3118,N_3493);
nand U4769 (N_4769,N_3579,N_3442);
xnor U4770 (N_4770,N_3472,N_3605);
or U4771 (N_4771,N_2843,N_2871);
nand U4772 (N_4772,N_2602,N_3077);
or U4773 (N_4773,N_3646,N_2528);
nand U4774 (N_4774,N_2745,N_2926);
nand U4775 (N_4775,N_2877,N_3502);
xor U4776 (N_4776,N_2941,N_3058);
or U4777 (N_4777,N_2525,N_3439);
nor U4778 (N_4778,N_2863,N_3252);
and U4779 (N_4779,N_2879,N_3524);
nor U4780 (N_4780,N_3333,N_2689);
and U4781 (N_4781,N_2516,N_2832);
nand U4782 (N_4782,N_2909,N_3695);
xnor U4783 (N_4783,N_2865,N_2677);
or U4784 (N_4784,N_3320,N_3242);
and U4785 (N_4785,N_3398,N_2884);
xnor U4786 (N_4786,N_3037,N_3489);
nand U4787 (N_4787,N_2899,N_3381);
nor U4788 (N_4788,N_3590,N_3030);
xor U4789 (N_4789,N_2937,N_3153);
xor U4790 (N_4790,N_3129,N_3181);
xor U4791 (N_4791,N_3547,N_2717);
nand U4792 (N_4792,N_2758,N_2713);
nor U4793 (N_4793,N_3297,N_2697);
or U4794 (N_4794,N_3025,N_3379);
nor U4795 (N_4795,N_3166,N_2608);
and U4796 (N_4796,N_3350,N_2976);
nand U4797 (N_4797,N_2557,N_3590);
xor U4798 (N_4798,N_3617,N_3301);
xnor U4799 (N_4799,N_3662,N_2684);
or U4800 (N_4800,N_3736,N_2504);
or U4801 (N_4801,N_3204,N_3210);
nor U4802 (N_4802,N_2862,N_3280);
nor U4803 (N_4803,N_3153,N_2552);
xnor U4804 (N_4804,N_3193,N_3383);
xnor U4805 (N_4805,N_3249,N_2571);
or U4806 (N_4806,N_3029,N_3599);
nand U4807 (N_4807,N_2914,N_2873);
and U4808 (N_4808,N_3106,N_2564);
and U4809 (N_4809,N_2577,N_2943);
nor U4810 (N_4810,N_3383,N_3309);
nand U4811 (N_4811,N_3203,N_2972);
or U4812 (N_4812,N_3212,N_3570);
nor U4813 (N_4813,N_3372,N_3324);
xor U4814 (N_4814,N_3640,N_2835);
and U4815 (N_4815,N_3662,N_2557);
xor U4816 (N_4816,N_3104,N_2887);
or U4817 (N_4817,N_3160,N_3435);
and U4818 (N_4818,N_3101,N_3706);
nor U4819 (N_4819,N_2684,N_3265);
nor U4820 (N_4820,N_3568,N_3041);
xor U4821 (N_4821,N_3591,N_2846);
xor U4822 (N_4822,N_2573,N_3627);
nand U4823 (N_4823,N_3718,N_2534);
or U4824 (N_4824,N_3334,N_3129);
and U4825 (N_4825,N_2897,N_3722);
or U4826 (N_4826,N_2615,N_2967);
xor U4827 (N_4827,N_3168,N_3483);
nand U4828 (N_4828,N_3080,N_3188);
and U4829 (N_4829,N_3215,N_2958);
or U4830 (N_4830,N_3083,N_3218);
xor U4831 (N_4831,N_3205,N_3530);
nand U4832 (N_4832,N_2912,N_3530);
and U4833 (N_4833,N_2649,N_2614);
nand U4834 (N_4834,N_3638,N_2781);
xnor U4835 (N_4835,N_2806,N_3034);
nand U4836 (N_4836,N_3540,N_2685);
nor U4837 (N_4837,N_2817,N_3391);
xor U4838 (N_4838,N_3049,N_3399);
nand U4839 (N_4839,N_3623,N_3548);
or U4840 (N_4840,N_3036,N_3486);
nand U4841 (N_4841,N_2983,N_3244);
or U4842 (N_4842,N_3614,N_2876);
nand U4843 (N_4843,N_2883,N_2622);
xnor U4844 (N_4844,N_3624,N_3000);
nor U4845 (N_4845,N_2534,N_3489);
nand U4846 (N_4846,N_3367,N_3074);
nand U4847 (N_4847,N_2623,N_2553);
nor U4848 (N_4848,N_2652,N_2674);
nor U4849 (N_4849,N_2969,N_2572);
nor U4850 (N_4850,N_2700,N_3584);
or U4851 (N_4851,N_3029,N_3232);
xnor U4852 (N_4852,N_2830,N_2790);
or U4853 (N_4853,N_3258,N_2745);
or U4854 (N_4854,N_3157,N_3729);
nor U4855 (N_4855,N_2950,N_2564);
or U4856 (N_4856,N_3657,N_2561);
nand U4857 (N_4857,N_3324,N_2781);
and U4858 (N_4858,N_3741,N_3018);
or U4859 (N_4859,N_3637,N_2838);
xor U4860 (N_4860,N_3530,N_2604);
nand U4861 (N_4861,N_3535,N_2924);
or U4862 (N_4862,N_3274,N_3176);
nor U4863 (N_4863,N_2899,N_3625);
nand U4864 (N_4864,N_3539,N_3378);
or U4865 (N_4865,N_3671,N_2892);
or U4866 (N_4866,N_2698,N_3080);
xor U4867 (N_4867,N_3163,N_3320);
nand U4868 (N_4868,N_3538,N_3349);
nor U4869 (N_4869,N_2638,N_2949);
and U4870 (N_4870,N_3495,N_3142);
nand U4871 (N_4871,N_2936,N_3000);
and U4872 (N_4872,N_3344,N_2856);
xor U4873 (N_4873,N_2847,N_2997);
nand U4874 (N_4874,N_2611,N_2750);
and U4875 (N_4875,N_3457,N_2528);
xor U4876 (N_4876,N_2642,N_2690);
xor U4877 (N_4877,N_3250,N_3521);
or U4878 (N_4878,N_3414,N_3609);
nor U4879 (N_4879,N_3552,N_3346);
or U4880 (N_4880,N_3376,N_3264);
or U4881 (N_4881,N_3274,N_2849);
xor U4882 (N_4882,N_3218,N_2816);
nand U4883 (N_4883,N_3579,N_3545);
and U4884 (N_4884,N_3496,N_2658);
or U4885 (N_4885,N_3494,N_2592);
nor U4886 (N_4886,N_2890,N_2815);
or U4887 (N_4887,N_3326,N_2663);
xnor U4888 (N_4888,N_3131,N_3441);
or U4889 (N_4889,N_2577,N_3195);
nand U4890 (N_4890,N_3319,N_3491);
nand U4891 (N_4891,N_3344,N_2832);
or U4892 (N_4892,N_3170,N_2746);
nand U4893 (N_4893,N_3585,N_3474);
nand U4894 (N_4894,N_3634,N_3463);
nand U4895 (N_4895,N_3381,N_3474);
nand U4896 (N_4896,N_3150,N_2674);
nor U4897 (N_4897,N_3294,N_2786);
nand U4898 (N_4898,N_2998,N_2852);
and U4899 (N_4899,N_3452,N_3132);
nand U4900 (N_4900,N_2836,N_3098);
nor U4901 (N_4901,N_3524,N_3183);
or U4902 (N_4902,N_2538,N_3350);
nor U4903 (N_4903,N_2757,N_3098);
nor U4904 (N_4904,N_2797,N_2642);
and U4905 (N_4905,N_3322,N_2982);
and U4906 (N_4906,N_3031,N_3522);
nor U4907 (N_4907,N_3544,N_3442);
nor U4908 (N_4908,N_3479,N_3418);
and U4909 (N_4909,N_2797,N_2706);
and U4910 (N_4910,N_2540,N_2512);
nor U4911 (N_4911,N_2560,N_3421);
nor U4912 (N_4912,N_2584,N_2712);
nand U4913 (N_4913,N_3270,N_2981);
or U4914 (N_4914,N_3552,N_2793);
nand U4915 (N_4915,N_2753,N_2797);
or U4916 (N_4916,N_3067,N_2930);
or U4917 (N_4917,N_3238,N_3048);
or U4918 (N_4918,N_2606,N_2965);
xor U4919 (N_4919,N_3435,N_3675);
and U4920 (N_4920,N_3681,N_3568);
or U4921 (N_4921,N_3210,N_3193);
nand U4922 (N_4922,N_2673,N_3406);
nand U4923 (N_4923,N_2892,N_3305);
nor U4924 (N_4924,N_2995,N_2897);
nand U4925 (N_4925,N_3717,N_2656);
nor U4926 (N_4926,N_2616,N_3484);
xnor U4927 (N_4927,N_3267,N_2649);
nand U4928 (N_4928,N_3170,N_3653);
and U4929 (N_4929,N_3164,N_2605);
xor U4930 (N_4930,N_2673,N_2684);
xnor U4931 (N_4931,N_3106,N_3128);
nor U4932 (N_4932,N_2627,N_3142);
and U4933 (N_4933,N_3032,N_3215);
nor U4934 (N_4934,N_2763,N_2672);
nand U4935 (N_4935,N_3245,N_2795);
xor U4936 (N_4936,N_2676,N_3169);
and U4937 (N_4937,N_3269,N_2582);
xor U4938 (N_4938,N_3026,N_2712);
nor U4939 (N_4939,N_3721,N_3426);
or U4940 (N_4940,N_3581,N_2690);
nor U4941 (N_4941,N_2662,N_3446);
or U4942 (N_4942,N_2695,N_3631);
or U4943 (N_4943,N_2723,N_3160);
nor U4944 (N_4944,N_2920,N_3734);
nand U4945 (N_4945,N_3496,N_3485);
or U4946 (N_4946,N_2567,N_3350);
nand U4947 (N_4947,N_3436,N_3345);
or U4948 (N_4948,N_3185,N_2659);
nor U4949 (N_4949,N_2566,N_3019);
or U4950 (N_4950,N_2944,N_3310);
xnor U4951 (N_4951,N_3561,N_2854);
nor U4952 (N_4952,N_2947,N_3405);
and U4953 (N_4953,N_3695,N_3649);
nand U4954 (N_4954,N_2611,N_2890);
nor U4955 (N_4955,N_3499,N_2990);
nand U4956 (N_4956,N_2998,N_2940);
nand U4957 (N_4957,N_3401,N_3317);
or U4958 (N_4958,N_3602,N_3000);
xnor U4959 (N_4959,N_3287,N_3351);
xnor U4960 (N_4960,N_2775,N_3599);
nand U4961 (N_4961,N_3749,N_3108);
and U4962 (N_4962,N_2787,N_3418);
nand U4963 (N_4963,N_2831,N_3412);
xnor U4964 (N_4964,N_3039,N_2799);
nor U4965 (N_4965,N_3296,N_3046);
nand U4966 (N_4966,N_3205,N_3260);
and U4967 (N_4967,N_3057,N_2784);
nand U4968 (N_4968,N_3667,N_2799);
or U4969 (N_4969,N_3049,N_3520);
xor U4970 (N_4970,N_3496,N_2735);
nand U4971 (N_4971,N_3720,N_2624);
nor U4972 (N_4972,N_2809,N_2734);
nand U4973 (N_4973,N_3521,N_3079);
nor U4974 (N_4974,N_3396,N_3665);
or U4975 (N_4975,N_2962,N_3707);
xor U4976 (N_4976,N_3463,N_3003);
nand U4977 (N_4977,N_2906,N_2703);
or U4978 (N_4978,N_3652,N_3340);
or U4979 (N_4979,N_3447,N_3448);
xnor U4980 (N_4980,N_3419,N_3527);
or U4981 (N_4981,N_3717,N_3329);
nor U4982 (N_4982,N_3667,N_2759);
and U4983 (N_4983,N_3225,N_3523);
xnor U4984 (N_4984,N_2835,N_3497);
xor U4985 (N_4985,N_3382,N_3498);
or U4986 (N_4986,N_3692,N_3634);
nor U4987 (N_4987,N_2801,N_3367);
nand U4988 (N_4988,N_3545,N_2762);
nand U4989 (N_4989,N_2523,N_3361);
nor U4990 (N_4990,N_3744,N_2824);
xnor U4991 (N_4991,N_3112,N_3486);
and U4992 (N_4992,N_3538,N_2643);
nor U4993 (N_4993,N_3164,N_3695);
xor U4994 (N_4994,N_2725,N_3410);
xor U4995 (N_4995,N_3162,N_3279);
nand U4996 (N_4996,N_3408,N_3487);
and U4997 (N_4997,N_3555,N_2772);
and U4998 (N_4998,N_3589,N_2792);
and U4999 (N_4999,N_2537,N_3129);
nor U5000 (N_5000,N_4216,N_4495);
nand U5001 (N_5001,N_4866,N_3963);
and U5002 (N_5002,N_4985,N_4843);
and U5003 (N_5003,N_4473,N_3934);
nor U5004 (N_5004,N_4362,N_4978);
xnor U5005 (N_5005,N_4748,N_4011);
or U5006 (N_5006,N_3806,N_4123);
nand U5007 (N_5007,N_3971,N_4348);
nand U5008 (N_5008,N_4766,N_4304);
and U5009 (N_5009,N_4772,N_4644);
or U5010 (N_5010,N_4100,N_3756);
and U5011 (N_5011,N_4835,N_3938);
xnor U5012 (N_5012,N_4744,N_4285);
or U5013 (N_5013,N_3751,N_4196);
nor U5014 (N_5014,N_4399,N_3845);
and U5015 (N_5015,N_3814,N_4230);
xnor U5016 (N_5016,N_4208,N_3798);
nand U5017 (N_5017,N_3995,N_3973);
and U5018 (N_5018,N_4541,N_4825);
xor U5019 (N_5019,N_4195,N_4253);
or U5020 (N_5020,N_4725,N_4817);
or U5021 (N_5021,N_4366,N_4865);
xor U5022 (N_5022,N_4297,N_3812);
xnor U5023 (N_5023,N_4104,N_4702);
xnor U5024 (N_5024,N_3854,N_3948);
or U5025 (N_5025,N_3771,N_4331);
xor U5026 (N_5026,N_3828,N_4176);
nand U5027 (N_5027,N_4819,N_4309);
xor U5028 (N_5028,N_4977,N_4501);
and U5029 (N_5029,N_4633,N_3762);
and U5030 (N_5030,N_4875,N_4869);
nand U5031 (N_5031,N_4169,N_4719);
and U5032 (N_5032,N_4642,N_4911);
and U5033 (N_5033,N_4530,N_4679);
and U5034 (N_5034,N_4701,N_4528);
or U5035 (N_5035,N_4481,N_4807);
nor U5036 (N_5036,N_4155,N_4874);
or U5037 (N_5037,N_3778,N_4082);
and U5038 (N_5038,N_4885,N_3989);
and U5039 (N_5039,N_4424,N_4578);
nand U5040 (N_5040,N_4929,N_4747);
and U5041 (N_5041,N_4496,N_4686);
nand U5042 (N_5042,N_4832,N_4147);
xor U5043 (N_5043,N_4326,N_4849);
or U5044 (N_5044,N_4788,N_4654);
or U5045 (N_5045,N_4862,N_4574);
nand U5046 (N_5046,N_4806,N_4171);
xor U5047 (N_5047,N_4863,N_4181);
or U5048 (N_5048,N_4880,N_3884);
nand U5049 (N_5049,N_4466,N_4061);
and U5050 (N_5050,N_4520,N_4937);
and U5051 (N_5051,N_3876,N_4507);
nand U5052 (N_5052,N_4342,N_4969);
nand U5053 (N_5053,N_4858,N_4096);
or U5054 (N_5054,N_4666,N_4314);
and U5055 (N_5055,N_3839,N_4135);
nand U5056 (N_5056,N_3918,N_3920);
nor U5057 (N_5057,N_4222,N_3803);
nor U5058 (N_5058,N_4197,N_4095);
nand U5059 (N_5059,N_3895,N_4349);
nand U5060 (N_5060,N_4044,N_4795);
and U5061 (N_5061,N_4796,N_3793);
nand U5062 (N_5062,N_4895,N_4925);
and U5063 (N_5063,N_4791,N_3997);
or U5064 (N_5064,N_4370,N_4357);
or U5065 (N_5065,N_4514,N_4535);
and U5066 (N_5066,N_4598,N_4251);
nor U5067 (N_5067,N_4497,N_4793);
nor U5068 (N_5068,N_4846,N_4143);
nand U5069 (N_5069,N_4469,N_3979);
and U5070 (N_5070,N_4632,N_4465);
or U5071 (N_5071,N_4160,N_4560);
nand U5072 (N_5072,N_4960,N_3908);
or U5073 (N_5073,N_4919,N_4103);
nand U5074 (N_5074,N_4641,N_4760);
or U5075 (N_5075,N_4844,N_4539);
nand U5076 (N_5076,N_3942,N_4516);
nand U5077 (N_5077,N_3850,N_4831);
and U5078 (N_5078,N_4891,N_4042);
nand U5079 (N_5079,N_4274,N_4966);
nor U5080 (N_5080,N_4026,N_4391);
nand U5081 (N_5081,N_4752,N_4323);
and U5082 (N_5082,N_4470,N_4444);
nand U5083 (N_5083,N_4199,N_4436);
and U5084 (N_5084,N_4125,N_4649);
and U5085 (N_5085,N_4313,N_4939);
xnor U5086 (N_5086,N_3788,N_4665);
and U5087 (N_5087,N_4588,N_3841);
and U5088 (N_5088,N_4212,N_4322);
nor U5089 (N_5089,N_4689,N_4412);
nand U5090 (N_5090,N_3860,N_3919);
nand U5091 (N_5091,N_4664,N_3927);
xor U5092 (N_5092,N_4359,N_4965);
or U5093 (N_5093,N_4280,N_4685);
nand U5094 (N_5094,N_4585,N_4903);
nor U5095 (N_5095,N_4784,N_4250);
xnor U5096 (N_5096,N_4630,N_4433);
nor U5097 (N_5097,N_4119,N_4422);
nand U5098 (N_5098,N_4850,N_4316);
and U5099 (N_5099,N_4127,N_4211);
xnor U5100 (N_5100,N_4158,N_4434);
and U5101 (N_5101,N_4876,N_4474);
nor U5102 (N_5102,N_4833,N_4615);
nor U5103 (N_5103,N_4106,N_4109);
nand U5104 (N_5104,N_4695,N_4607);
xor U5105 (N_5105,N_3846,N_4975);
nand U5106 (N_5106,N_3880,N_4710);
or U5107 (N_5107,N_4418,N_4750);
xnor U5108 (N_5108,N_4899,N_4781);
and U5109 (N_5109,N_4035,N_3848);
or U5110 (N_5110,N_3832,N_4526);
xor U5111 (N_5111,N_4332,N_4740);
or U5112 (N_5112,N_3898,N_3835);
nor U5113 (N_5113,N_4311,N_4463);
xnor U5114 (N_5114,N_4484,N_4693);
and U5115 (N_5115,N_3914,N_4848);
nand U5116 (N_5116,N_4694,N_4471);
xor U5117 (N_5117,N_4955,N_4092);
nor U5118 (N_5118,N_4478,N_4651);
or U5119 (N_5119,N_4636,N_4838);
nand U5120 (N_5120,N_4543,N_4295);
and U5121 (N_5121,N_4797,N_4063);
and U5122 (N_5122,N_4732,N_4390);
xnor U5123 (N_5123,N_3802,N_4043);
or U5124 (N_5124,N_4967,N_4048);
nor U5125 (N_5125,N_4328,N_3752);
nand U5126 (N_5126,N_4924,N_4202);
nor U5127 (N_5127,N_4555,N_4237);
nand U5128 (N_5128,N_4745,N_4896);
xor U5129 (N_5129,N_4265,N_4724);
and U5130 (N_5130,N_3950,N_4175);
nand U5131 (N_5131,N_4993,N_4172);
and U5132 (N_5132,N_3833,N_3951);
nor U5133 (N_5133,N_3799,N_4234);
and U5134 (N_5134,N_4217,N_4137);
xor U5135 (N_5135,N_4413,N_4922);
xor U5136 (N_5136,N_4089,N_4868);
nor U5137 (N_5137,N_4557,N_4601);
and U5138 (N_5138,N_4226,N_4883);
and U5139 (N_5139,N_4565,N_4558);
nand U5140 (N_5140,N_4834,N_4957);
nand U5141 (N_5141,N_4626,N_4245);
xor U5142 (N_5142,N_4178,N_4236);
xor U5143 (N_5143,N_4718,N_4948);
xor U5144 (N_5144,N_4402,N_4839);
and U5145 (N_5145,N_3838,N_4472);
xor U5146 (N_5146,N_3954,N_4705);
xnor U5147 (N_5147,N_4900,N_4121);
nor U5148 (N_5148,N_3889,N_4249);
nand U5149 (N_5149,N_4406,N_4204);
nand U5150 (N_5150,N_3968,N_4681);
and U5151 (N_5151,N_4403,N_4811);
or U5152 (N_5152,N_4527,N_3953);
and U5153 (N_5153,N_4270,N_4301);
and U5154 (N_5154,N_4517,N_4003);
xor U5155 (N_5155,N_4462,N_4404);
nor U5156 (N_5156,N_3892,N_3776);
xnor U5157 (N_5157,N_4799,N_4684);
nand U5158 (N_5158,N_4656,N_4427);
nand U5159 (N_5159,N_3998,N_4266);
and U5160 (N_5160,N_4166,N_4736);
or U5161 (N_5161,N_4031,N_4284);
xnor U5162 (N_5162,N_4142,N_4170);
nor U5163 (N_5163,N_4518,N_4450);
nor U5164 (N_5164,N_4243,N_4131);
xor U5165 (N_5165,N_3900,N_3881);
and U5166 (N_5166,N_4203,N_4151);
or U5167 (N_5167,N_3780,N_3956);
nor U5168 (N_5168,N_3890,N_4224);
nor U5169 (N_5169,N_3753,N_4079);
or U5170 (N_5170,N_4376,N_3772);
xnor U5171 (N_5171,N_4532,N_4392);
nor U5172 (N_5172,N_4602,N_4809);
nand U5173 (N_5173,N_4380,N_4675);
nand U5174 (N_5174,N_4296,N_4460);
xor U5175 (N_5175,N_4647,N_4767);
xor U5176 (N_5176,N_4864,N_4974);
nor U5177 (N_5177,N_4521,N_4979);
or U5178 (N_5178,N_4918,N_3894);
nand U5179 (N_5179,N_4101,N_4416);
nand U5180 (N_5180,N_4374,N_4639);
nor U5181 (N_5181,N_4032,N_4655);
nand U5182 (N_5182,N_4408,N_3888);
nand U5183 (N_5183,N_3988,N_3755);
or U5184 (N_5184,N_3796,N_4298);
and U5185 (N_5185,N_4777,N_4591);
and U5186 (N_5186,N_4334,N_4491);
xnor U5187 (N_5187,N_4996,N_4814);
and U5188 (N_5188,N_4012,N_3815);
nor U5189 (N_5189,N_4477,N_4504);
xor U5190 (N_5190,N_4587,N_4581);
and U5191 (N_5191,N_4346,N_4947);
xor U5192 (N_5192,N_4486,N_4753);
nand U5193 (N_5193,N_4935,N_4882);
or U5194 (N_5194,N_4837,N_3999);
nand U5195 (N_5195,N_4091,N_4836);
and U5196 (N_5196,N_4361,N_4708);
and U5197 (N_5197,N_4625,N_3991);
and U5198 (N_5198,N_4480,N_4716);
nor U5199 (N_5199,N_3917,N_4191);
or U5200 (N_5200,N_3960,N_3872);
and U5201 (N_5201,N_4494,N_3840);
or U5202 (N_5202,N_4488,N_4529);
or U5203 (N_5203,N_4897,N_4859);
or U5204 (N_5204,N_3777,N_4886);
or U5205 (N_5205,N_4333,N_4085);
xor U5206 (N_5206,N_4546,N_4372);
nand U5207 (N_5207,N_3750,N_4431);
nand U5208 (N_5208,N_3873,N_4273);
and U5209 (N_5209,N_4768,N_4168);
and U5210 (N_5210,N_3763,N_4021);
xor U5211 (N_5211,N_4759,N_4099);
nor U5212 (N_5212,N_4713,N_4051);
nand U5213 (N_5213,N_4714,N_4064);
xor U5214 (N_5214,N_3851,N_4324);
nand U5215 (N_5215,N_4210,N_4873);
nor U5216 (N_5216,N_3924,N_4735);
nor U5217 (N_5217,N_3984,N_4658);
nand U5218 (N_5218,N_4177,N_4762);
xor U5219 (N_5219,N_4934,N_3844);
and U5220 (N_5220,N_3864,N_4786);
and U5221 (N_5221,N_4163,N_4648);
and U5222 (N_5222,N_4417,N_4743);
xnor U5223 (N_5223,N_4164,N_4697);
nor U5224 (N_5224,N_4257,N_4022);
nor U5225 (N_5225,N_4017,N_3817);
or U5226 (N_5226,N_4783,N_4442);
and U5227 (N_5227,N_4650,N_4126);
and U5228 (N_5228,N_3935,N_4419);
or U5229 (N_5229,N_3760,N_4592);
nor U5230 (N_5230,N_3822,N_4387);
and U5231 (N_5231,N_4200,N_4822);
and U5232 (N_5232,N_4148,N_4992);
nor U5233 (N_5233,N_4242,N_3930);
and U5234 (N_5234,N_4668,N_4940);
xor U5235 (N_5235,N_4890,N_4072);
xnor U5236 (N_5236,N_4277,N_3794);
nand U5237 (N_5237,N_4995,N_4667);
nor U5238 (N_5238,N_3855,N_3878);
nor U5239 (N_5239,N_4721,N_4606);
and U5240 (N_5240,N_4964,N_4040);
nand U5241 (N_5241,N_3945,N_3885);
nor U5242 (N_5242,N_4821,N_4379);
nand U5243 (N_5243,N_4938,N_4004);
and U5244 (N_5244,N_3931,N_3783);
nor U5245 (N_5245,N_4122,N_4782);
or U5246 (N_5246,N_4002,N_3964);
xnor U5247 (N_5247,N_4916,N_4299);
xnor U5248 (N_5248,N_4439,N_4174);
nor U5249 (N_5249,N_3940,N_3893);
xor U5250 (N_5250,N_4382,N_4842);
nand U5251 (N_5251,N_3868,N_4385);
or U5252 (N_5252,N_3903,N_4162);
nor U5253 (N_5253,N_4206,N_3768);
nand U5254 (N_5254,N_4437,N_4941);
nand U5255 (N_5255,N_3980,N_3784);
nor U5256 (N_5256,N_4586,N_4047);
nor U5257 (N_5257,N_4942,N_4464);
or U5258 (N_5258,N_4094,N_4423);
and U5259 (N_5259,N_3757,N_4828);
or U5260 (N_5260,N_4726,N_4909);
nand U5261 (N_5261,N_4114,N_4503);
nand U5262 (N_5262,N_4677,N_4000);
and U5263 (N_5263,N_4110,N_4787);
and U5264 (N_5264,N_4401,N_4027);
and U5265 (N_5265,N_4383,N_3972);
xnor U5266 (N_5266,N_4902,N_4506);
nor U5267 (N_5267,N_4608,N_4728);
nand U5268 (N_5268,N_4595,N_3819);
and U5269 (N_5269,N_4081,N_4049);
xor U5270 (N_5270,N_4435,N_4888);
nor U5271 (N_5271,N_4189,N_4640);
and U5272 (N_5272,N_4467,N_3759);
nor U5273 (N_5273,N_4704,N_4033);
and U5274 (N_5274,N_3852,N_4232);
nor U5275 (N_5275,N_4764,N_4623);
nor U5276 (N_5276,N_4548,N_4415);
nand U5277 (N_5277,N_4712,N_4145);
nor U5278 (N_5278,N_4926,N_4247);
or U5279 (N_5279,N_3787,N_3769);
xnor U5280 (N_5280,N_3804,N_4855);
or U5281 (N_5281,N_4421,N_4987);
and U5282 (N_5282,N_4563,N_4830);
xnor U5283 (N_5283,N_4059,N_4140);
nand U5284 (N_5284,N_4396,N_4510);
xor U5285 (N_5285,N_4998,N_3867);
or U5286 (N_5286,N_4258,N_4989);
nand U5287 (N_5287,N_3816,N_4534);
or U5288 (N_5288,N_3843,N_4330);
or U5289 (N_5289,N_4877,N_4617);
xnor U5290 (N_5290,N_4511,N_3791);
and U5291 (N_5291,N_4898,N_4915);
or U5292 (N_5292,N_4997,N_4146);
xnor U5293 (N_5293,N_4933,N_4816);
and U5294 (N_5294,N_4192,N_4315);
xnor U5295 (N_5295,N_4347,N_4225);
xnor U5296 (N_5296,N_4046,N_4156);
nand U5297 (N_5297,N_4884,N_4559);
xor U5298 (N_5298,N_4432,N_4860);
xor U5299 (N_5299,N_4183,N_4050);
and U5300 (N_5300,N_4167,N_4575);
nand U5301 (N_5301,N_3773,N_4931);
nand U5302 (N_5302,N_4010,N_4871);
or U5303 (N_5303,N_4275,N_3910);
and U5304 (N_5304,N_4209,N_4893);
xor U5305 (N_5305,N_4981,N_4138);
xnor U5306 (N_5306,N_4154,N_4075);
and U5307 (N_5307,N_4930,N_4986);
and U5308 (N_5308,N_4566,N_4589);
xor U5309 (N_5309,N_4643,N_4205);
xor U5310 (N_5310,N_4824,N_4680);
nor U5311 (N_5311,N_3807,N_3825);
xor U5312 (N_5312,N_4238,N_4182);
nor U5313 (N_5313,N_4827,N_4709);
xor U5314 (N_5314,N_4455,N_4845);
or U5315 (N_5315,N_4340,N_3899);
nor U5316 (N_5316,N_3823,N_4776);
nor U5317 (N_5317,N_4310,N_4308);
xnor U5318 (N_5318,N_4620,N_4739);
or U5319 (N_5319,N_4599,N_4678);
nor U5320 (N_5320,N_3758,N_4971);
nor U5321 (N_5321,N_4134,N_3949);
and U5322 (N_5322,N_3785,N_4687);
xor U5323 (N_5323,N_3958,N_4813);
xnor U5324 (N_5324,N_4983,N_4117);
and U5325 (N_5325,N_4388,N_3859);
or U5326 (N_5326,N_4228,N_4512);
and U5327 (N_5327,N_4577,N_4276);
nor U5328 (N_5328,N_4373,N_4515);
xor U5329 (N_5329,N_4287,N_4812);
and U5330 (N_5330,N_4912,N_4005);
xnor U5331 (N_5331,N_4272,N_4271);
and U5332 (N_5332,N_4722,N_3905);
xnor U5333 (N_5333,N_3865,N_3926);
or U5334 (N_5334,N_4857,N_4461);
xnor U5335 (N_5335,N_4384,N_3826);
and U5336 (N_5336,N_4988,N_4235);
nor U5337 (N_5337,N_4364,N_4339);
or U5338 (N_5338,N_4561,N_4624);
and U5339 (N_5339,N_3863,N_4778);
or U5340 (N_5340,N_4319,N_4800);
and U5341 (N_5341,N_4213,N_4706);
xnor U5342 (N_5342,N_4653,N_4219);
nor U5343 (N_5343,N_4723,N_4030);
and U5344 (N_5344,N_4944,N_4962);
xnor U5345 (N_5345,N_3824,N_4758);
nor U5346 (N_5346,N_4847,N_4377);
nor U5347 (N_5347,N_4594,N_3925);
nor U5348 (N_5348,N_4805,N_3976);
nor U5349 (N_5349,N_4028,N_3974);
and U5350 (N_5350,N_3808,N_4547);
xnor U5351 (N_5351,N_4984,N_4593);
or U5352 (N_5352,N_3982,N_4283);
and U5353 (N_5353,N_4892,N_4785);
nand U5354 (N_5354,N_4045,N_4479);
nor U5355 (N_5355,N_4553,N_4731);
nand U5356 (N_5356,N_4792,N_4227);
xnor U5357 (N_5357,N_3818,N_3767);
xor U5358 (N_5358,N_3975,N_3830);
and U5359 (N_5359,N_4150,N_3955);
xnor U5360 (N_5360,N_4889,N_4129);
nand U5361 (N_5361,N_4808,N_3786);
xor U5362 (N_5362,N_4352,N_3766);
or U5363 (N_5363,N_3936,N_4982);
nor U5364 (N_5364,N_4703,N_4286);
nor U5365 (N_5365,N_4818,N_4300);
nor U5366 (N_5366,N_4688,N_4771);
xor U5367 (N_5367,N_3883,N_4956);
xnor U5368 (N_5368,N_3874,N_4698);
or U5369 (N_5369,N_4621,N_3990);
nand U5370 (N_5370,N_4070,N_4670);
xor U5371 (N_5371,N_3907,N_4928);
or U5372 (N_5372,N_3882,N_4854);
nor U5373 (N_5373,N_4755,N_4810);
nand U5374 (N_5374,N_4262,N_4756);
nor U5375 (N_5375,N_3837,N_4240);
or U5376 (N_5376,N_4562,N_4738);
and U5377 (N_5377,N_4305,N_3932);
and U5378 (N_5378,N_4088,N_4634);
xnor U5379 (N_5379,N_4958,N_3805);
or U5380 (N_5380,N_4492,N_3779);
xor U5381 (N_5381,N_4108,N_4550);
and U5382 (N_5382,N_4329,N_4959);
and U5383 (N_5383,N_4306,N_4907);
and U5384 (N_5384,N_4618,N_4152);
or U5385 (N_5385,N_4256,N_4102);
and U5386 (N_5386,N_4921,N_4531);
or U5387 (N_5387,N_4963,N_4097);
and U5388 (N_5388,N_4368,N_4278);
xnor U5389 (N_5389,N_4446,N_4006);
nor U5390 (N_5390,N_4034,N_4917);
or U5391 (N_5391,N_4699,N_4394);
and U5392 (N_5392,N_3912,N_4303);
nor U5393 (N_5393,N_4980,N_4801);
and U5394 (N_5394,N_4090,N_4073);
nand U5395 (N_5395,N_4335,N_3970);
and U5396 (N_5396,N_3929,N_3901);
nand U5397 (N_5397,N_4248,N_4609);
nand U5398 (N_5398,N_4290,N_4727);
xor U5399 (N_5399,N_4596,N_4438);
nor U5400 (N_5400,N_3857,N_4545);
nand U5401 (N_5401,N_4337,N_3981);
xnor U5402 (N_5402,N_4386,N_4500);
or U5403 (N_5403,N_3891,N_4887);
nor U5404 (N_5404,N_4733,N_4001);
xnor U5405 (N_5405,N_4533,N_4954);
or U5406 (N_5406,N_4360,N_4829);
nor U5407 (N_5407,N_4815,N_3811);
nand U5408 (N_5408,N_4338,N_4690);
or U5409 (N_5409,N_3962,N_4268);
or U5410 (N_5410,N_3858,N_4552);
and U5411 (N_5411,N_3829,N_4780);
or U5412 (N_5412,N_3915,N_4638);
xnor U5413 (N_5413,N_4645,N_4619);
xor U5414 (N_5414,N_4062,N_4950);
nand U5415 (N_5415,N_4254,N_4878);
nor U5416 (N_5416,N_3941,N_4537);
nor U5417 (N_5417,N_4389,N_3765);
and U5418 (N_5418,N_4223,N_4584);
nand U5419 (N_5419,N_3849,N_4024);
or U5420 (N_5420,N_4672,N_4908);
and U5421 (N_5421,N_4207,N_3875);
nand U5422 (N_5422,N_4186,N_4751);
xnor U5423 (N_5423,N_4614,N_4054);
nor U5424 (N_5424,N_4336,N_4105);
nor U5425 (N_5425,N_4066,N_4676);
nor U5426 (N_5426,N_4779,N_4369);
and U5427 (N_5427,N_4113,N_4970);
nand U5428 (N_5428,N_3754,N_4635);
or U5429 (N_5429,N_4525,N_4008);
nor U5430 (N_5430,N_4674,N_4184);
or U5431 (N_5431,N_4583,N_4426);
and U5432 (N_5432,N_4325,N_4130);
or U5433 (N_5433,N_4407,N_4294);
and U5434 (N_5434,N_4239,N_4057);
nor U5435 (N_5435,N_3810,N_4261);
nand U5436 (N_5436,N_4913,N_4972);
nand U5437 (N_5437,N_4393,N_4973);
nor U5438 (N_5438,N_4905,N_3923);
or U5439 (N_5439,N_3946,N_4267);
nand U5440 (N_5440,N_4746,N_4132);
or U5441 (N_5441,N_3977,N_4524);
nor U5442 (N_5442,N_4078,N_4058);
nor U5443 (N_5443,N_4646,N_4020);
xnor U5444 (N_5444,N_4519,N_4741);
nand U5445 (N_5445,N_3809,N_4263);
xnor U5446 (N_5446,N_4165,N_4600);
nor U5447 (N_5447,N_4037,N_3870);
nand U5448 (N_5448,N_4029,N_4356);
and U5449 (N_5449,N_4111,N_4794);
or U5450 (N_5450,N_4683,N_4445);
or U5451 (N_5451,N_4136,N_4489);
nand U5452 (N_5452,N_4945,N_4400);
nand U5453 (N_5453,N_4293,N_4569);
xor U5454 (N_5454,N_4867,N_4080);
xnor U5455 (N_5455,N_4367,N_3909);
or U5456 (N_5456,N_4409,N_3820);
nand U5457 (N_5457,N_4682,N_4657);
nand U5458 (N_5458,N_3792,N_4802);
and U5459 (N_5459,N_4804,N_4904);
or U5460 (N_5460,N_3821,N_3853);
xor U5461 (N_5461,N_3827,N_3801);
xor U5462 (N_5462,N_4269,N_3897);
and U5463 (N_5463,N_4468,N_3774);
or U5464 (N_5464,N_4425,N_4637);
nand U5465 (N_5465,N_4861,N_4579);
or U5466 (N_5466,N_4729,N_3813);
and U5467 (N_5467,N_4180,N_3781);
or U5468 (N_5468,N_4659,N_4055);
or U5469 (N_5469,N_4023,N_4214);
and U5470 (N_5470,N_4700,N_4039);
nor U5471 (N_5471,N_4483,N_4513);
and U5472 (N_5472,N_4961,N_3966);
xnor U5473 (N_5473,N_4014,N_4789);
or U5474 (N_5474,N_3913,N_4823);
nor U5475 (N_5475,N_4482,N_4536);
nor U5476 (N_5476,N_4093,N_4149);
xor U5477 (N_5477,N_4429,N_4341);
xor U5478 (N_5478,N_3869,N_4065);
and U5479 (N_5479,N_4879,N_4611);
or U5480 (N_5480,N_4628,N_4949);
xnor U5481 (N_5481,N_4840,N_4790);
and U5482 (N_5482,N_4307,N_4894);
or U5483 (N_5483,N_3877,N_4264);
nand U5484 (N_5484,N_4803,N_4321);
xnor U5485 (N_5485,N_3775,N_4255);
nand U5486 (N_5486,N_4604,N_3795);
and U5487 (N_5487,N_4720,N_4673);
xor U5488 (N_5488,N_4198,N_4449);
nand U5489 (N_5489,N_4540,N_4717);
and U5490 (N_5490,N_4355,N_4820);
nor U5491 (N_5491,N_4144,N_4025);
xnor U5492 (N_5492,N_4910,N_3896);
nor U5493 (N_5493,N_4943,N_4318);
nand U5494 (N_5494,N_4568,N_4652);
nand U5495 (N_5495,N_4730,N_4187);
and U5496 (N_5496,N_4289,N_4053);
nand U5497 (N_5497,N_4009,N_4071);
nand U5498 (N_5498,N_3836,N_4179);
and U5499 (N_5499,N_4443,N_4139);
or U5500 (N_5500,N_4086,N_4398);
or U5501 (N_5501,N_4734,N_4320);
nor U5502 (N_5502,N_4233,N_4508);
nor U5503 (N_5503,N_4302,N_4414);
xor U5504 (N_5504,N_4556,N_4188);
and U5505 (N_5505,N_4194,N_4523);
nor U5506 (N_5506,N_3983,N_4502);
xnor U5507 (N_5507,N_4671,N_4953);
and U5508 (N_5508,N_3879,N_3944);
nand U5509 (N_5509,N_4629,N_4952);
xnor U5510 (N_5510,N_4661,N_4757);
xor U5511 (N_5511,N_4153,N_4067);
xor U5512 (N_5512,N_4448,N_4410);
nor U5513 (N_5513,N_4076,N_4378);
or U5514 (N_5514,N_4395,N_4036);
xor U5515 (N_5515,N_4570,N_4549);
xor U5516 (N_5516,N_4851,N_4411);
or U5517 (N_5517,N_4038,N_4260);
and U5518 (N_5518,N_4292,N_4068);
or U5519 (N_5519,N_3916,N_3921);
nand U5520 (N_5520,N_3939,N_4259);
or U5521 (N_5521,N_4493,N_3922);
nand U5522 (N_5522,N_4554,N_3902);
nand U5523 (N_5523,N_4098,N_4441);
nor U5524 (N_5524,N_3961,N_4551);
and U5525 (N_5525,N_4018,N_4007);
xor U5526 (N_5526,N_4932,N_4737);
xnor U5527 (N_5527,N_3831,N_4190);
nor U5528 (N_5528,N_4770,N_4215);
or U5529 (N_5529,N_4327,N_4381);
nor U5530 (N_5530,N_3789,N_4841);
nor U5531 (N_5531,N_3959,N_3847);
nand U5532 (N_5532,N_4990,N_4826);
or U5533 (N_5533,N_3770,N_4692);
or U5534 (N_5534,N_4707,N_4711);
nand U5535 (N_5535,N_4610,N_4282);
xnor U5536 (N_5536,N_4691,N_3911);
and U5537 (N_5537,N_4087,N_4765);
xnor U5538 (N_5538,N_4798,N_4773);
or U5539 (N_5539,N_4505,N_4405);
nand U5540 (N_5540,N_4976,N_4041);
nand U5541 (N_5541,N_4923,N_4490);
nor U5542 (N_5542,N_3886,N_4576);
xor U5543 (N_5543,N_4509,N_3871);
xor U5544 (N_5544,N_4288,N_4371);
nand U5545 (N_5545,N_4452,N_4013);
nand U5546 (N_5546,N_4358,N_4696);
nor U5547 (N_5547,N_3842,N_4159);
xor U5548 (N_5548,N_4116,N_4279);
nor U5549 (N_5549,N_4453,N_4603);
or U5550 (N_5550,N_4968,N_4185);
xnor U5551 (N_5551,N_4580,N_4572);
nor U5552 (N_5552,N_3993,N_4084);
nor U5553 (N_5553,N_3861,N_4920);
nand U5554 (N_5554,N_4991,N_3992);
xor U5555 (N_5555,N_4120,N_4281);
nor U5556 (N_5556,N_4906,N_3943);
nand U5557 (N_5557,N_4458,N_3978);
nand U5558 (N_5558,N_4241,N_4083);
nor U5559 (N_5559,N_4133,N_4456);
xor U5560 (N_5560,N_4077,N_4015);
and U5561 (N_5561,N_4475,N_3887);
and U5562 (N_5562,N_4573,N_4244);
or U5563 (N_5563,N_4498,N_4669);
nor U5564 (N_5564,N_4345,N_4420);
or U5565 (N_5565,N_4440,N_3856);
or U5566 (N_5566,N_3965,N_4201);
nor U5567 (N_5567,N_4754,N_4128);
and U5568 (N_5568,N_4597,N_4107);
nor U5569 (N_5569,N_4447,N_4019);
nand U5570 (N_5570,N_4775,N_4715);
nor U5571 (N_5571,N_4060,N_4763);
xor U5572 (N_5572,N_3904,N_3987);
nand U5573 (N_5573,N_3797,N_4375);
xnor U5574 (N_5574,N_4220,N_3834);
nor U5575 (N_5575,N_4193,N_4343);
or U5576 (N_5576,N_4430,N_4622);
or U5577 (N_5577,N_4457,N_4124);
or U5578 (N_5578,N_3906,N_4853);
and U5579 (N_5579,N_3969,N_4872);
nand U5580 (N_5580,N_3957,N_4901);
nand U5581 (N_5581,N_3952,N_4365);
or U5582 (N_5582,N_4605,N_4522);
xnor U5583 (N_5583,N_4946,N_4218);
or U5584 (N_5584,N_4999,N_4016);
xnor U5585 (N_5585,N_4612,N_4582);
and U5586 (N_5586,N_4141,N_4056);
or U5587 (N_5587,N_4852,N_3928);
or U5588 (N_5588,N_4291,N_3986);
nand U5589 (N_5589,N_4761,N_4660);
nor U5590 (N_5590,N_4459,N_4317);
and U5591 (N_5591,N_4994,N_4631);
nand U5592 (N_5592,N_4353,N_4774);
nor U5593 (N_5593,N_4856,N_4157);
nor U5594 (N_5594,N_4914,N_4542);
and U5595 (N_5595,N_4052,N_4112);
xor U5596 (N_5596,N_4571,N_4613);
nor U5597 (N_5597,N_4161,N_4544);
nand U5598 (N_5598,N_4173,N_3994);
and U5599 (N_5599,N_3761,N_4881);
or U5600 (N_5600,N_4662,N_3800);
or U5601 (N_5601,N_4451,N_4246);
nor U5602 (N_5602,N_4590,N_4487);
nor U5603 (N_5603,N_3996,N_4428);
nand U5604 (N_5604,N_4627,N_4951);
nor U5605 (N_5605,N_4397,N_3782);
and U5606 (N_5606,N_4354,N_4936);
xor U5607 (N_5607,N_4663,N_4742);
or U5608 (N_5608,N_4485,N_4454);
or U5609 (N_5609,N_3967,N_4118);
nor U5610 (N_5610,N_4616,N_4927);
nand U5611 (N_5611,N_4749,N_4351);
and U5612 (N_5612,N_4229,N_4567);
xor U5613 (N_5613,N_4363,N_3790);
nand U5614 (N_5614,N_3764,N_3937);
nor U5615 (N_5615,N_3862,N_4252);
nand U5616 (N_5616,N_4538,N_4499);
and U5617 (N_5617,N_4221,N_4870);
nand U5618 (N_5618,N_4312,N_4564);
nor U5619 (N_5619,N_3866,N_4344);
nor U5620 (N_5620,N_3933,N_4350);
xnor U5621 (N_5621,N_3947,N_4074);
nor U5622 (N_5622,N_4069,N_4115);
xnor U5623 (N_5623,N_4231,N_4476);
xnor U5624 (N_5624,N_4769,N_3985);
or U5625 (N_5625,N_4382,N_4046);
xor U5626 (N_5626,N_4680,N_3847);
or U5627 (N_5627,N_4653,N_4391);
xnor U5628 (N_5628,N_4068,N_4531);
xnor U5629 (N_5629,N_4087,N_4555);
xor U5630 (N_5630,N_4619,N_4627);
nor U5631 (N_5631,N_4004,N_4462);
nor U5632 (N_5632,N_4621,N_4443);
xor U5633 (N_5633,N_3759,N_3985);
nor U5634 (N_5634,N_4625,N_4913);
nor U5635 (N_5635,N_3902,N_4865);
nand U5636 (N_5636,N_4108,N_4018);
nand U5637 (N_5637,N_4453,N_4410);
xnor U5638 (N_5638,N_4806,N_4941);
or U5639 (N_5639,N_4828,N_4719);
or U5640 (N_5640,N_4799,N_4647);
and U5641 (N_5641,N_4345,N_4535);
or U5642 (N_5642,N_4575,N_4060);
nand U5643 (N_5643,N_3769,N_4544);
nand U5644 (N_5644,N_4270,N_4468);
xor U5645 (N_5645,N_4569,N_4312);
and U5646 (N_5646,N_4085,N_4077);
or U5647 (N_5647,N_3883,N_4254);
xnor U5648 (N_5648,N_4747,N_4780);
xnor U5649 (N_5649,N_4861,N_4809);
nor U5650 (N_5650,N_4939,N_4052);
nor U5651 (N_5651,N_3895,N_4631);
nor U5652 (N_5652,N_3752,N_4211);
nand U5653 (N_5653,N_4797,N_4286);
nand U5654 (N_5654,N_4082,N_4595);
and U5655 (N_5655,N_4413,N_4356);
nand U5656 (N_5656,N_4976,N_4575);
or U5657 (N_5657,N_4841,N_4865);
xor U5658 (N_5658,N_4685,N_4556);
xor U5659 (N_5659,N_3817,N_4690);
xor U5660 (N_5660,N_4250,N_4347);
nor U5661 (N_5661,N_4230,N_4503);
and U5662 (N_5662,N_4628,N_4046);
and U5663 (N_5663,N_3818,N_4139);
xor U5664 (N_5664,N_4111,N_4290);
and U5665 (N_5665,N_4888,N_3922);
or U5666 (N_5666,N_3848,N_4018);
xnor U5667 (N_5667,N_4458,N_4203);
nor U5668 (N_5668,N_4117,N_4071);
or U5669 (N_5669,N_4726,N_4418);
xnor U5670 (N_5670,N_3792,N_4758);
and U5671 (N_5671,N_4266,N_4319);
nor U5672 (N_5672,N_4573,N_4949);
nor U5673 (N_5673,N_3779,N_3926);
nor U5674 (N_5674,N_4360,N_3930);
or U5675 (N_5675,N_4437,N_4481);
or U5676 (N_5676,N_4582,N_4717);
nand U5677 (N_5677,N_4260,N_4686);
or U5678 (N_5678,N_4490,N_4743);
or U5679 (N_5679,N_4210,N_4469);
nand U5680 (N_5680,N_3871,N_4627);
and U5681 (N_5681,N_4487,N_4472);
or U5682 (N_5682,N_4962,N_3937);
or U5683 (N_5683,N_4506,N_4822);
xor U5684 (N_5684,N_4671,N_4928);
xnor U5685 (N_5685,N_4417,N_4529);
and U5686 (N_5686,N_3902,N_3864);
xnor U5687 (N_5687,N_3958,N_4693);
and U5688 (N_5688,N_4397,N_4692);
nor U5689 (N_5689,N_4290,N_3947);
xor U5690 (N_5690,N_3932,N_4206);
and U5691 (N_5691,N_3762,N_4954);
or U5692 (N_5692,N_4087,N_4945);
or U5693 (N_5693,N_4718,N_4172);
nor U5694 (N_5694,N_4524,N_4952);
xnor U5695 (N_5695,N_4718,N_4380);
xnor U5696 (N_5696,N_4862,N_4330);
or U5697 (N_5697,N_4544,N_4568);
nor U5698 (N_5698,N_3789,N_4647);
and U5699 (N_5699,N_4295,N_4757);
and U5700 (N_5700,N_3753,N_4624);
or U5701 (N_5701,N_4026,N_4313);
xor U5702 (N_5702,N_4038,N_4785);
xor U5703 (N_5703,N_4665,N_4477);
and U5704 (N_5704,N_4613,N_4014);
or U5705 (N_5705,N_3753,N_4008);
xnor U5706 (N_5706,N_4469,N_3964);
nor U5707 (N_5707,N_3969,N_4998);
nor U5708 (N_5708,N_4246,N_3998);
or U5709 (N_5709,N_3919,N_4142);
nand U5710 (N_5710,N_4097,N_4491);
nand U5711 (N_5711,N_4728,N_4743);
or U5712 (N_5712,N_4631,N_4825);
nor U5713 (N_5713,N_4825,N_4318);
xor U5714 (N_5714,N_4555,N_4903);
xnor U5715 (N_5715,N_4843,N_4294);
xnor U5716 (N_5716,N_3933,N_4015);
xor U5717 (N_5717,N_4676,N_4568);
or U5718 (N_5718,N_4156,N_4769);
and U5719 (N_5719,N_4471,N_4070);
nand U5720 (N_5720,N_3934,N_4822);
and U5721 (N_5721,N_4949,N_4697);
xor U5722 (N_5722,N_3774,N_3935);
xor U5723 (N_5723,N_4189,N_3822);
nand U5724 (N_5724,N_4770,N_4374);
xnor U5725 (N_5725,N_4487,N_4290);
nor U5726 (N_5726,N_4716,N_4535);
nor U5727 (N_5727,N_4083,N_3866);
nor U5728 (N_5728,N_4969,N_4373);
and U5729 (N_5729,N_4739,N_4598);
xnor U5730 (N_5730,N_4301,N_4202);
nand U5731 (N_5731,N_4930,N_3888);
and U5732 (N_5732,N_4421,N_4546);
and U5733 (N_5733,N_4814,N_4270);
or U5734 (N_5734,N_4899,N_4809);
nor U5735 (N_5735,N_3774,N_3922);
xor U5736 (N_5736,N_4580,N_3888);
xor U5737 (N_5737,N_4877,N_4799);
nor U5738 (N_5738,N_3770,N_4840);
or U5739 (N_5739,N_4209,N_4033);
xor U5740 (N_5740,N_4509,N_3996);
nand U5741 (N_5741,N_4596,N_4212);
xor U5742 (N_5742,N_3949,N_4983);
and U5743 (N_5743,N_4430,N_4043);
or U5744 (N_5744,N_3967,N_4392);
xnor U5745 (N_5745,N_4074,N_4591);
or U5746 (N_5746,N_4169,N_4115);
and U5747 (N_5747,N_4719,N_4622);
nand U5748 (N_5748,N_4396,N_4274);
nor U5749 (N_5749,N_3977,N_3770);
and U5750 (N_5750,N_4011,N_4759);
and U5751 (N_5751,N_4591,N_3901);
xnor U5752 (N_5752,N_4338,N_4576);
xnor U5753 (N_5753,N_3874,N_4841);
or U5754 (N_5754,N_4022,N_4245);
or U5755 (N_5755,N_4267,N_4206);
nand U5756 (N_5756,N_4670,N_3751);
xnor U5757 (N_5757,N_4601,N_3795);
or U5758 (N_5758,N_3909,N_4970);
and U5759 (N_5759,N_4325,N_4029);
nand U5760 (N_5760,N_4745,N_4824);
nor U5761 (N_5761,N_4152,N_3790);
and U5762 (N_5762,N_3842,N_4559);
and U5763 (N_5763,N_4888,N_4811);
nand U5764 (N_5764,N_4109,N_4899);
xor U5765 (N_5765,N_4483,N_3966);
and U5766 (N_5766,N_4117,N_3972);
or U5767 (N_5767,N_3761,N_4756);
or U5768 (N_5768,N_4659,N_4200);
nor U5769 (N_5769,N_4300,N_4108);
or U5770 (N_5770,N_4195,N_4025);
nor U5771 (N_5771,N_4706,N_3754);
nand U5772 (N_5772,N_4354,N_4394);
or U5773 (N_5773,N_4658,N_4959);
nand U5774 (N_5774,N_3922,N_4982);
xor U5775 (N_5775,N_3909,N_4804);
nand U5776 (N_5776,N_3834,N_4997);
nor U5777 (N_5777,N_4208,N_4547);
xnor U5778 (N_5778,N_4421,N_3913);
xor U5779 (N_5779,N_4172,N_4346);
and U5780 (N_5780,N_4042,N_4857);
xnor U5781 (N_5781,N_4962,N_4440);
and U5782 (N_5782,N_4558,N_4569);
nand U5783 (N_5783,N_4151,N_4571);
nand U5784 (N_5784,N_4871,N_4360);
or U5785 (N_5785,N_4903,N_4691);
nand U5786 (N_5786,N_4731,N_4543);
nor U5787 (N_5787,N_4175,N_4019);
nor U5788 (N_5788,N_3812,N_4126);
and U5789 (N_5789,N_4942,N_4301);
nor U5790 (N_5790,N_4416,N_4029);
xor U5791 (N_5791,N_4994,N_4147);
or U5792 (N_5792,N_4948,N_3965);
nand U5793 (N_5793,N_3987,N_4353);
nor U5794 (N_5794,N_4074,N_4371);
or U5795 (N_5795,N_3756,N_3980);
and U5796 (N_5796,N_3791,N_4225);
xor U5797 (N_5797,N_4586,N_4306);
and U5798 (N_5798,N_4319,N_4262);
and U5799 (N_5799,N_4509,N_3990);
nor U5800 (N_5800,N_3956,N_4128);
or U5801 (N_5801,N_4696,N_4963);
nor U5802 (N_5802,N_3964,N_4636);
nand U5803 (N_5803,N_4351,N_4555);
or U5804 (N_5804,N_4465,N_4590);
nor U5805 (N_5805,N_4496,N_4310);
xnor U5806 (N_5806,N_4153,N_4037);
and U5807 (N_5807,N_4253,N_3758);
xnor U5808 (N_5808,N_4369,N_4430);
nand U5809 (N_5809,N_3972,N_4764);
nor U5810 (N_5810,N_4985,N_4707);
nand U5811 (N_5811,N_4737,N_3826);
or U5812 (N_5812,N_4935,N_4244);
xor U5813 (N_5813,N_3811,N_4916);
xnor U5814 (N_5814,N_4306,N_4215);
nand U5815 (N_5815,N_4698,N_4005);
nand U5816 (N_5816,N_4278,N_4947);
or U5817 (N_5817,N_4949,N_3902);
or U5818 (N_5818,N_3816,N_4440);
and U5819 (N_5819,N_4093,N_3824);
and U5820 (N_5820,N_4883,N_4786);
or U5821 (N_5821,N_3804,N_3811);
xnor U5822 (N_5822,N_4656,N_3945);
or U5823 (N_5823,N_4582,N_4485);
or U5824 (N_5824,N_3931,N_4381);
xnor U5825 (N_5825,N_4037,N_4442);
xor U5826 (N_5826,N_4242,N_4515);
xor U5827 (N_5827,N_4895,N_4112);
xnor U5828 (N_5828,N_4824,N_4634);
nand U5829 (N_5829,N_4134,N_3775);
nor U5830 (N_5830,N_4840,N_4209);
xor U5831 (N_5831,N_4637,N_4234);
and U5832 (N_5832,N_4447,N_3851);
xnor U5833 (N_5833,N_3998,N_4985);
xor U5834 (N_5834,N_4339,N_4014);
nand U5835 (N_5835,N_4926,N_4658);
or U5836 (N_5836,N_4206,N_4435);
and U5837 (N_5837,N_4673,N_4445);
nand U5838 (N_5838,N_4699,N_4427);
or U5839 (N_5839,N_4406,N_4602);
xor U5840 (N_5840,N_4989,N_4845);
nand U5841 (N_5841,N_4854,N_4006);
nor U5842 (N_5842,N_4209,N_4922);
or U5843 (N_5843,N_3875,N_4156);
xnor U5844 (N_5844,N_3921,N_4313);
and U5845 (N_5845,N_4545,N_3810);
nand U5846 (N_5846,N_4225,N_4639);
and U5847 (N_5847,N_4095,N_4282);
nor U5848 (N_5848,N_4453,N_3755);
nand U5849 (N_5849,N_4656,N_3774);
xnor U5850 (N_5850,N_3936,N_3838);
or U5851 (N_5851,N_4819,N_4374);
or U5852 (N_5852,N_4374,N_4182);
xor U5853 (N_5853,N_4728,N_3858);
nand U5854 (N_5854,N_4681,N_4523);
or U5855 (N_5855,N_4194,N_3852);
xnor U5856 (N_5856,N_4712,N_4423);
nand U5857 (N_5857,N_4317,N_4698);
nor U5858 (N_5858,N_4077,N_4425);
and U5859 (N_5859,N_4207,N_4406);
xnor U5860 (N_5860,N_3833,N_4633);
nor U5861 (N_5861,N_4026,N_4989);
nor U5862 (N_5862,N_4587,N_3823);
and U5863 (N_5863,N_4236,N_3877);
and U5864 (N_5864,N_4915,N_4104);
nand U5865 (N_5865,N_3976,N_3751);
nor U5866 (N_5866,N_3956,N_3934);
and U5867 (N_5867,N_3759,N_4218);
xor U5868 (N_5868,N_4043,N_4217);
and U5869 (N_5869,N_4021,N_4660);
nand U5870 (N_5870,N_3979,N_4750);
and U5871 (N_5871,N_4716,N_4747);
nor U5872 (N_5872,N_3916,N_4675);
nand U5873 (N_5873,N_4072,N_4473);
or U5874 (N_5874,N_4812,N_4717);
xnor U5875 (N_5875,N_4293,N_3856);
nor U5876 (N_5876,N_3769,N_4113);
nor U5877 (N_5877,N_4233,N_4515);
xnor U5878 (N_5878,N_4908,N_4832);
nand U5879 (N_5879,N_4094,N_3933);
or U5880 (N_5880,N_4428,N_4998);
and U5881 (N_5881,N_4696,N_4029);
and U5882 (N_5882,N_4224,N_3835);
xor U5883 (N_5883,N_4523,N_4768);
or U5884 (N_5884,N_4677,N_4216);
nor U5885 (N_5885,N_4010,N_4703);
nand U5886 (N_5886,N_4646,N_3828);
and U5887 (N_5887,N_4062,N_4315);
or U5888 (N_5888,N_4577,N_4574);
nor U5889 (N_5889,N_4805,N_4190);
xor U5890 (N_5890,N_3868,N_4411);
and U5891 (N_5891,N_4562,N_3973);
nor U5892 (N_5892,N_4554,N_3924);
or U5893 (N_5893,N_4737,N_4380);
xor U5894 (N_5894,N_4709,N_4894);
and U5895 (N_5895,N_3916,N_3910);
and U5896 (N_5896,N_4603,N_3948);
nor U5897 (N_5897,N_4778,N_4073);
or U5898 (N_5898,N_4247,N_3946);
and U5899 (N_5899,N_4317,N_4522);
xor U5900 (N_5900,N_4856,N_3874);
nor U5901 (N_5901,N_3806,N_4977);
xnor U5902 (N_5902,N_4641,N_4085);
xor U5903 (N_5903,N_4160,N_4484);
nand U5904 (N_5904,N_4494,N_4190);
or U5905 (N_5905,N_4284,N_4594);
nor U5906 (N_5906,N_4550,N_3989);
and U5907 (N_5907,N_4414,N_4785);
nand U5908 (N_5908,N_3799,N_3771);
nand U5909 (N_5909,N_4522,N_4308);
xor U5910 (N_5910,N_3965,N_3884);
or U5911 (N_5911,N_4100,N_4499);
xor U5912 (N_5912,N_3896,N_3759);
or U5913 (N_5913,N_4808,N_4946);
xnor U5914 (N_5914,N_4131,N_4364);
xor U5915 (N_5915,N_4094,N_3994);
and U5916 (N_5916,N_3772,N_4115);
nand U5917 (N_5917,N_4166,N_4239);
nand U5918 (N_5918,N_4486,N_4897);
xor U5919 (N_5919,N_4584,N_4207);
or U5920 (N_5920,N_4282,N_4832);
nor U5921 (N_5921,N_4551,N_4323);
and U5922 (N_5922,N_3847,N_4667);
nor U5923 (N_5923,N_4058,N_4845);
nor U5924 (N_5924,N_4501,N_4482);
nand U5925 (N_5925,N_4215,N_3811);
xnor U5926 (N_5926,N_4091,N_4291);
xor U5927 (N_5927,N_4467,N_4525);
nand U5928 (N_5928,N_4341,N_4954);
xor U5929 (N_5929,N_4610,N_4373);
and U5930 (N_5930,N_4826,N_3866);
nor U5931 (N_5931,N_3825,N_4497);
nand U5932 (N_5932,N_4748,N_4816);
nand U5933 (N_5933,N_4467,N_3812);
or U5934 (N_5934,N_3852,N_4493);
and U5935 (N_5935,N_3859,N_4465);
nor U5936 (N_5936,N_4482,N_3983);
nand U5937 (N_5937,N_4102,N_4536);
nand U5938 (N_5938,N_4726,N_4389);
nor U5939 (N_5939,N_4047,N_4936);
or U5940 (N_5940,N_4832,N_3989);
nor U5941 (N_5941,N_3928,N_4243);
xnor U5942 (N_5942,N_4174,N_4870);
and U5943 (N_5943,N_4312,N_4916);
or U5944 (N_5944,N_4818,N_4843);
and U5945 (N_5945,N_4853,N_4223);
or U5946 (N_5946,N_4123,N_3962);
nand U5947 (N_5947,N_4974,N_4920);
xor U5948 (N_5948,N_4317,N_4403);
xnor U5949 (N_5949,N_4210,N_4376);
xor U5950 (N_5950,N_4872,N_4272);
nand U5951 (N_5951,N_4639,N_4898);
and U5952 (N_5952,N_3986,N_4745);
nand U5953 (N_5953,N_4158,N_4291);
nand U5954 (N_5954,N_4263,N_4209);
xnor U5955 (N_5955,N_4457,N_4605);
and U5956 (N_5956,N_3863,N_3958);
nor U5957 (N_5957,N_3834,N_4346);
xnor U5958 (N_5958,N_4524,N_3976);
nor U5959 (N_5959,N_4147,N_4583);
and U5960 (N_5960,N_4920,N_4147);
xnor U5961 (N_5961,N_4410,N_4556);
nor U5962 (N_5962,N_3980,N_4307);
nand U5963 (N_5963,N_4220,N_3812);
nor U5964 (N_5964,N_3808,N_4449);
and U5965 (N_5965,N_4462,N_4697);
xnor U5966 (N_5966,N_4215,N_4910);
nand U5967 (N_5967,N_4127,N_4073);
nand U5968 (N_5968,N_4480,N_4294);
nor U5969 (N_5969,N_4031,N_4763);
nand U5970 (N_5970,N_4226,N_4255);
or U5971 (N_5971,N_4624,N_4977);
nor U5972 (N_5972,N_3917,N_4768);
and U5973 (N_5973,N_4493,N_4591);
xor U5974 (N_5974,N_4549,N_4935);
and U5975 (N_5975,N_4331,N_4452);
xnor U5976 (N_5976,N_3806,N_4186);
nor U5977 (N_5977,N_4533,N_4562);
nand U5978 (N_5978,N_4312,N_4688);
xor U5979 (N_5979,N_4959,N_4072);
or U5980 (N_5980,N_4410,N_4023);
nand U5981 (N_5981,N_4894,N_4016);
nand U5982 (N_5982,N_4458,N_4687);
nor U5983 (N_5983,N_4641,N_3807);
nand U5984 (N_5984,N_4459,N_3790);
xnor U5985 (N_5985,N_4814,N_4003);
nor U5986 (N_5986,N_4818,N_4272);
or U5987 (N_5987,N_4773,N_3906);
xnor U5988 (N_5988,N_3942,N_4597);
xnor U5989 (N_5989,N_4789,N_4286);
and U5990 (N_5990,N_4552,N_4792);
and U5991 (N_5991,N_4308,N_3801);
xor U5992 (N_5992,N_3909,N_4749);
nor U5993 (N_5993,N_4793,N_3795);
xor U5994 (N_5994,N_4535,N_4343);
or U5995 (N_5995,N_4845,N_4549);
or U5996 (N_5996,N_4232,N_4217);
nor U5997 (N_5997,N_4528,N_4498);
nor U5998 (N_5998,N_4189,N_4568);
or U5999 (N_5999,N_4585,N_3981);
and U6000 (N_6000,N_4877,N_4533);
nor U6001 (N_6001,N_4208,N_4603);
nand U6002 (N_6002,N_4934,N_4172);
nor U6003 (N_6003,N_4879,N_3910);
nand U6004 (N_6004,N_4664,N_4447);
nor U6005 (N_6005,N_4693,N_4101);
xnor U6006 (N_6006,N_4129,N_3930);
nor U6007 (N_6007,N_4235,N_4873);
xnor U6008 (N_6008,N_4809,N_4992);
or U6009 (N_6009,N_3821,N_4848);
and U6010 (N_6010,N_4202,N_3866);
nand U6011 (N_6011,N_4773,N_3813);
xor U6012 (N_6012,N_4825,N_4179);
nor U6013 (N_6013,N_4322,N_4649);
and U6014 (N_6014,N_4725,N_4248);
nand U6015 (N_6015,N_4830,N_4966);
nor U6016 (N_6016,N_4150,N_4100);
and U6017 (N_6017,N_4345,N_4520);
nor U6018 (N_6018,N_3900,N_4747);
nor U6019 (N_6019,N_4570,N_4099);
and U6020 (N_6020,N_3909,N_4675);
nor U6021 (N_6021,N_4800,N_3812);
and U6022 (N_6022,N_4951,N_3820);
nand U6023 (N_6023,N_3987,N_4939);
or U6024 (N_6024,N_4672,N_4531);
nor U6025 (N_6025,N_4915,N_4068);
xnor U6026 (N_6026,N_4751,N_4319);
xor U6027 (N_6027,N_4132,N_4120);
nand U6028 (N_6028,N_4911,N_4395);
xor U6029 (N_6029,N_4372,N_4853);
nand U6030 (N_6030,N_3980,N_4760);
nand U6031 (N_6031,N_4718,N_4859);
and U6032 (N_6032,N_4659,N_4709);
and U6033 (N_6033,N_4802,N_3856);
nand U6034 (N_6034,N_3947,N_4879);
xor U6035 (N_6035,N_4101,N_4497);
nor U6036 (N_6036,N_3865,N_4452);
and U6037 (N_6037,N_4638,N_4458);
nand U6038 (N_6038,N_4455,N_3964);
nor U6039 (N_6039,N_4155,N_4733);
xnor U6040 (N_6040,N_4588,N_3755);
nand U6041 (N_6041,N_4512,N_4964);
or U6042 (N_6042,N_4716,N_4197);
nor U6043 (N_6043,N_3835,N_4725);
nand U6044 (N_6044,N_4165,N_3870);
nand U6045 (N_6045,N_4138,N_4148);
or U6046 (N_6046,N_4331,N_3805);
xnor U6047 (N_6047,N_4169,N_3920);
xor U6048 (N_6048,N_4470,N_4930);
nand U6049 (N_6049,N_4964,N_4748);
nand U6050 (N_6050,N_4330,N_4164);
or U6051 (N_6051,N_4206,N_4543);
nor U6052 (N_6052,N_3829,N_4315);
or U6053 (N_6053,N_4871,N_3793);
nor U6054 (N_6054,N_4958,N_4095);
nor U6055 (N_6055,N_4596,N_4876);
nor U6056 (N_6056,N_3983,N_4461);
nor U6057 (N_6057,N_4344,N_4574);
nand U6058 (N_6058,N_3839,N_4195);
and U6059 (N_6059,N_3934,N_4616);
and U6060 (N_6060,N_4698,N_4384);
nand U6061 (N_6061,N_4179,N_4817);
and U6062 (N_6062,N_4347,N_3881);
or U6063 (N_6063,N_4446,N_4157);
and U6064 (N_6064,N_4654,N_4469);
nor U6065 (N_6065,N_3978,N_4749);
nor U6066 (N_6066,N_4755,N_4664);
and U6067 (N_6067,N_3798,N_4797);
xor U6068 (N_6068,N_4596,N_3870);
nor U6069 (N_6069,N_3988,N_4101);
and U6070 (N_6070,N_4134,N_4074);
nand U6071 (N_6071,N_4051,N_4263);
or U6072 (N_6072,N_4322,N_4259);
xor U6073 (N_6073,N_4789,N_3867);
nand U6074 (N_6074,N_4993,N_4502);
nand U6075 (N_6075,N_3860,N_4602);
or U6076 (N_6076,N_3819,N_3939);
and U6077 (N_6077,N_4490,N_3868);
nand U6078 (N_6078,N_4060,N_4552);
nor U6079 (N_6079,N_4257,N_3755);
nand U6080 (N_6080,N_4015,N_3758);
and U6081 (N_6081,N_4260,N_4545);
nand U6082 (N_6082,N_3952,N_4001);
and U6083 (N_6083,N_4978,N_4612);
xnor U6084 (N_6084,N_4161,N_4201);
and U6085 (N_6085,N_4581,N_4998);
nor U6086 (N_6086,N_4653,N_4919);
and U6087 (N_6087,N_4595,N_3781);
and U6088 (N_6088,N_4920,N_4248);
or U6089 (N_6089,N_4068,N_4596);
xor U6090 (N_6090,N_3965,N_4882);
or U6091 (N_6091,N_4106,N_4427);
or U6092 (N_6092,N_4720,N_4375);
nand U6093 (N_6093,N_3835,N_4842);
xnor U6094 (N_6094,N_4352,N_4286);
xor U6095 (N_6095,N_3878,N_3988);
nor U6096 (N_6096,N_4445,N_4648);
nand U6097 (N_6097,N_4150,N_3831);
and U6098 (N_6098,N_4494,N_4277);
nand U6099 (N_6099,N_4242,N_4341);
and U6100 (N_6100,N_4493,N_4203);
or U6101 (N_6101,N_4938,N_3989);
or U6102 (N_6102,N_4008,N_4337);
nor U6103 (N_6103,N_4057,N_4040);
xnor U6104 (N_6104,N_4711,N_4339);
and U6105 (N_6105,N_4517,N_3992);
or U6106 (N_6106,N_3882,N_4077);
nor U6107 (N_6107,N_4158,N_4564);
nand U6108 (N_6108,N_4131,N_4988);
nor U6109 (N_6109,N_4503,N_3761);
nor U6110 (N_6110,N_4626,N_3953);
and U6111 (N_6111,N_4024,N_4283);
or U6112 (N_6112,N_4330,N_4948);
or U6113 (N_6113,N_4104,N_4161);
xnor U6114 (N_6114,N_4157,N_3843);
nor U6115 (N_6115,N_3843,N_4741);
xor U6116 (N_6116,N_4916,N_3952);
nand U6117 (N_6117,N_3755,N_4454);
xnor U6118 (N_6118,N_4906,N_3781);
or U6119 (N_6119,N_4335,N_4389);
or U6120 (N_6120,N_3789,N_4884);
nand U6121 (N_6121,N_3922,N_4808);
and U6122 (N_6122,N_4422,N_3830);
nand U6123 (N_6123,N_4741,N_4009);
nand U6124 (N_6124,N_4929,N_4935);
nor U6125 (N_6125,N_4751,N_4914);
xnor U6126 (N_6126,N_4960,N_4477);
xnor U6127 (N_6127,N_3865,N_4585);
nor U6128 (N_6128,N_4911,N_4708);
nand U6129 (N_6129,N_4790,N_4054);
nor U6130 (N_6130,N_4791,N_4499);
xor U6131 (N_6131,N_4381,N_4959);
and U6132 (N_6132,N_4943,N_4392);
or U6133 (N_6133,N_4116,N_4492);
nor U6134 (N_6134,N_4574,N_4404);
xor U6135 (N_6135,N_4675,N_4541);
and U6136 (N_6136,N_3754,N_4733);
and U6137 (N_6137,N_4446,N_4073);
xnor U6138 (N_6138,N_4251,N_4548);
nand U6139 (N_6139,N_4213,N_4773);
nand U6140 (N_6140,N_4447,N_4963);
nand U6141 (N_6141,N_3940,N_4671);
and U6142 (N_6142,N_4922,N_4143);
xor U6143 (N_6143,N_4980,N_4850);
xor U6144 (N_6144,N_3822,N_4839);
and U6145 (N_6145,N_4205,N_4746);
nor U6146 (N_6146,N_4073,N_4853);
xnor U6147 (N_6147,N_4440,N_4044);
and U6148 (N_6148,N_3763,N_4479);
nor U6149 (N_6149,N_4791,N_3867);
nor U6150 (N_6150,N_4234,N_4733);
nor U6151 (N_6151,N_4370,N_4355);
and U6152 (N_6152,N_4964,N_3930);
nor U6153 (N_6153,N_4369,N_4888);
or U6154 (N_6154,N_4966,N_4500);
xnor U6155 (N_6155,N_4470,N_3788);
nor U6156 (N_6156,N_4248,N_4475);
nor U6157 (N_6157,N_4138,N_4723);
or U6158 (N_6158,N_4010,N_4322);
or U6159 (N_6159,N_4823,N_4910);
xnor U6160 (N_6160,N_4362,N_4569);
xor U6161 (N_6161,N_4326,N_4451);
nand U6162 (N_6162,N_4421,N_4389);
nor U6163 (N_6163,N_4442,N_4315);
or U6164 (N_6164,N_4901,N_4089);
and U6165 (N_6165,N_4187,N_4194);
xnor U6166 (N_6166,N_4739,N_4658);
or U6167 (N_6167,N_4433,N_4839);
nand U6168 (N_6168,N_3876,N_4315);
and U6169 (N_6169,N_3801,N_4544);
nand U6170 (N_6170,N_4644,N_4301);
and U6171 (N_6171,N_4498,N_4737);
nor U6172 (N_6172,N_4032,N_3798);
and U6173 (N_6173,N_4598,N_3757);
or U6174 (N_6174,N_4553,N_4078);
nand U6175 (N_6175,N_4532,N_4035);
nand U6176 (N_6176,N_4141,N_4930);
nor U6177 (N_6177,N_4854,N_4038);
nor U6178 (N_6178,N_4505,N_3968);
nand U6179 (N_6179,N_4215,N_4643);
xnor U6180 (N_6180,N_4495,N_3797);
or U6181 (N_6181,N_3766,N_3933);
xor U6182 (N_6182,N_4331,N_4561);
and U6183 (N_6183,N_4329,N_4228);
xnor U6184 (N_6184,N_4219,N_4223);
and U6185 (N_6185,N_4232,N_4543);
nor U6186 (N_6186,N_4556,N_4908);
nand U6187 (N_6187,N_4295,N_4363);
or U6188 (N_6188,N_4289,N_3922);
or U6189 (N_6189,N_4141,N_3933);
xor U6190 (N_6190,N_4017,N_4325);
nand U6191 (N_6191,N_4332,N_4726);
nor U6192 (N_6192,N_4477,N_4974);
nor U6193 (N_6193,N_4610,N_4396);
nand U6194 (N_6194,N_4282,N_4200);
nand U6195 (N_6195,N_3950,N_4220);
nand U6196 (N_6196,N_4308,N_4767);
or U6197 (N_6197,N_4127,N_4602);
nand U6198 (N_6198,N_4967,N_4000);
xor U6199 (N_6199,N_4661,N_4578);
nor U6200 (N_6200,N_4718,N_4265);
and U6201 (N_6201,N_4218,N_4826);
nor U6202 (N_6202,N_3920,N_4483);
and U6203 (N_6203,N_4555,N_4394);
xor U6204 (N_6204,N_3989,N_4203);
or U6205 (N_6205,N_4110,N_4422);
nor U6206 (N_6206,N_4958,N_4330);
and U6207 (N_6207,N_4514,N_4342);
and U6208 (N_6208,N_4492,N_4380);
and U6209 (N_6209,N_4441,N_4409);
nand U6210 (N_6210,N_3978,N_4774);
xnor U6211 (N_6211,N_4566,N_4837);
nand U6212 (N_6212,N_4700,N_3788);
and U6213 (N_6213,N_3855,N_4463);
xnor U6214 (N_6214,N_4934,N_4227);
and U6215 (N_6215,N_4860,N_4679);
nor U6216 (N_6216,N_4883,N_4495);
nand U6217 (N_6217,N_4083,N_4687);
xor U6218 (N_6218,N_4464,N_4513);
nand U6219 (N_6219,N_4738,N_4351);
xnor U6220 (N_6220,N_3850,N_3779);
and U6221 (N_6221,N_4965,N_4171);
nor U6222 (N_6222,N_4253,N_4126);
or U6223 (N_6223,N_4768,N_4141);
xnor U6224 (N_6224,N_4742,N_4977);
nor U6225 (N_6225,N_4842,N_4992);
nor U6226 (N_6226,N_4047,N_4844);
xor U6227 (N_6227,N_3857,N_4742);
nor U6228 (N_6228,N_4693,N_4876);
xnor U6229 (N_6229,N_4325,N_3969);
xor U6230 (N_6230,N_4957,N_4476);
nand U6231 (N_6231,N_4617,N_4598);
xnor U6232 (N_6232,N_4646,N_4334);
or U6233 (N_6233,N_3810,N_3837);
nand U6234 (N_6234,N_4648,N_3828);
or U6235 (N_6235,N_4511,N_4598);
or U6236 (N_6236,N_4753,N_4662);
nor U6237 (N_6237,N_4222,N_4878);
nor U6238 (N_6238,N_4595,N_3879);
and U6239 (N_6239,N_4765,N_4527);
xor U6240 (N_6240,N_4390,N_4877);
nand U6241 (N_6241,N_4870,N_4882);
xor U6242 (N_6242,N_4094,N_4064);
nand U6243 (N_6243,N_4453,N_4667);
xor U6244 (N_6244,N_4980,N_4261);
nand U6245 (N_6245,N_4997,N_4878);
and U6246 (N_6246,N_4655,N_4017);
nor U6247 (N_6247,N_4959,N_4530);
xor U6248 (N_6248,N_3799,N_3757);
xnor U6249 (N_6249,N_4586,N_4432);
or U6250 (N_6250,N_5991,N_5431);
nor U6251 (N_6251,N_6156,N_5376);
and U6252 (N_6252,N_5496,N_6119);
or U6253 (N_6253,N_5081,N_5167);
nor U6254 (N_6254,N_5780,N_5965);
xnor U6255 (N_6255,N_5914,N_6182);
nand U6256 (N_6256,N_6009,N_5162);
or U6257 (N_6257,N_5428,N_5394);
and U6258 (N_6258,N_5146,N_6231);
and U6259 (N_6259,N_5970,N_5193);
and U6260 (N_6260,N_5282,N_6089);
and U6261 (N_6261,N_5690,N_5044);
or U6262 (N_6262,N_5020,N_5318);
xor U6263 (N_6263,N_5570,N_6055);
or U6264 (N_6264,N_5753,N_5077);
and U6265 (N_6265,N_5601,N_5072);
and U6266 (N_6266,N_5211,N_5281);
and U6267 (N_6267,N_6073,N_5485);
nand U6268 (N_6268,N_5385,N_6022);
nand U6269 (N_6269,N_5721,N_5210);
or U6270 (N_6270,N_6214,N_5479);
or U6271 (N_6271,N_5748,N_5616);
nand U6272 (N_6272,N_5239,N_5252);
xor U6273 (N_6273,N_6130,N_5164);
xor U6274 (N_6274,N_5054,N_6082);
xor U6275 (N_6275,N_5157,N_5313);
and U6276 (N_6276,N_5108,N_6035);
nand U6277 (N_6277,N_5097,N_6065);
and U6278 (N_6278,N_5585,N_5664);
and U6279 (N_6279,N_5076,N_5047);
nand U6280 (N_6280,N_5170,N_5336);
and U6281 (N_6281,N_5316,N_6056);
nand U6282 (N_6282,N_6019,N_5544);
nor U6283 (N_6283,N_5499,N_5326);
and U6284 (N_6284,N_5728,N_5695);
and U6285 (N_6285,N_6144,N_5540);
xor U6286 (N_6286,N_5660,N_5738);
xor U6287 (N_6287,N_5986,N_5899);
or U6288 (N_6288,N_5090,N_5073);
or U6289 (N_6289,N_6034,N_6048);
xor U6290 (N_6290,N_5174,N_5907);
and U6291 (N_6291,N_5468,N_5953);
and U6292 (N_6292,N_6099,N_5353);
nand U6293 (N_6293,N_6139,N_5286);
xor U6294 (N_6294,N_6216,N_5471);
xor U6295 (N_6295,N_5079,N_5637);
and U6296 (N_6296,N_5181,N_6206);
and U6297 (N_6297,N_5040,N_5216);
and U6298 (N_6298,N_5103,N_5696);
xnor U6299 (N_6299,N_5543,N_5250);
xor U6300 (N_6300,N_5848,N_6087);
and U6301 (N_6301,N_5602,N_5561);
xnor U6302 (N_6302,N_5635,N_5667);
nand U6303 (N_6303,N_5041,N_5045);
and U6304 (N_6304,N_5972,N_5930);
and U6305 (N_6305,N_5547,N_5135);
nand U6306 (N_6306,N_6166,N_6049);
or U6307 (N_6307,N_5746,N_5118);
xor U6308 (N_6308,N_5777,N_5159);
nand U6309 (N_6309,N_6234,N_6064);
nand U6310 (N_6310,N_5994,N_5199);
nand U6311 (N_6311,N_6159,N_5673);
xnor U6312 (N_6312,N_6249,N_6208);
and U6313 (N_6313,N_5367,N_5620);
or U6314 (N_6314,N_5618,N_5904);
or U6315 (N_6315,N_5888,N_5507);
and U6316 (N_6316,N_5574,N_5990);
nand U6317 (N_6317,N_5708,N_5098);
nand U6318 (N_6318,N_5617,N_5249);
nor U6319 (N_6319,N_5232,N_5137);
nor U6320 (N_6320,N_5508,N_6026);
or U6321 (N_6321,N_5973,N_5562);
nand U6322 (N_6322,N_6017,N_6225);
xor U6323 (N_6323,N_6097,N_5225);
or U6324 (N_6324,N_5466,N_5450);
xnor U6325 (N_6325,N_5587,N_5614);
nor U6326 (N_6326,N_5010,N_5091);
nor U6327 (N_6327,N_5224,N_5947);
and U6328 (N_6328,N_6115,N_6143);
xnor U6329 (N_6329,N_6021,N_5887);
or U6330 (N_6330,N_5593,N_6188);
and U6331 (N_6331,N_6190,N_6107);
nand U6332 (N_6332,N_6239,N_5788);
and U6333 (N_6333,N_5104,N_5112);
nor U6334 (N_6334,N_5706,N_6170);
or U6335 (N_6335,N_5577,N_6062);
or U6336 (N_6336,N_5084,N_5329);
xor U6337 (N_6337,N_5530,N_5056);
xnor U6338 (N_6338,N_5130,N_5343);
nor U6339 (N_6339,N_5865,N_5554);
xnor U6340 (N_6340,N_6078,N_5787);
or U6341 (N_6341,N_5327,N_6189);
nor U6342 (N_6342,N_5911,N_5944);
xnor U6343 (N_6343,N_5219,N_5548);
or U6344 (N_6344,N_5491,N_5426);
nor U6345 (N_6345,N_5589,N_5458);
nor U6346 (N_6346,N_5785,N_5852);
xor U6347 (N_6347,N_5786,N_5303);
and U6348 (N_6348,N_5568,N_5226);
and U6349 (N_6349,N_5029,N_5808);
or U6350 (N_6350,N_6212,N_5334);
nand U6351 (N_6351,N_6007,N_6210);
xor U6352 (N_6352,N_5014,N_5338);
nand U6353 (N_6353,N_5378,N_5348);
and U6354 (N_6354,N_5743,N_5525);
nor U6355 (N_6355,N_5682,N_6185);
nand U6356 (N_6356,N_5576,N_5939);
nor U6357 (N_6357,N_5908,N_5946);
or U6358 (N_6358,N_5846,N_5950);
or U6359 (N_6359,N_5532,N_5732);
nor U6360 (N_6360,N_5075,N_5173);
nand U6361 (N_6361,N_5534,N_6042);
nor U6362 (N_6362,N_5957,N_5228);
and U6363 (N_6363,N_5653,N_6142);
nor U6364 (N_6364,N_5258,N_5046);
xor U6365 (N_6365,N_5767,N_5280);
xor U6366 (N_6366,N_6134,N_5154);
nand U6367 (N_6367,N_6132,N_5579);
xnor U6368 (N_6368,N_5565,N_5409);
or U6369 (N_6369,N_6108,N_5429);
nor U6370 (N_6370,N_5514,N_5215);
and U6371 (N_6371,N_5423,N_5051);
or U6372 (N_6372,N_5897,N_5415);
xnor U6373 (N_6373,N_5257,N_5920);
nand U6374 (N_6374,N_5085,N_5034);
nand U6375 (N_6375,N_5681,N_5190);
xor U6376 (N_6376,N_5838,N_5810);
nand U6377 (N_6377,N_5275,N_5149);
nand U6378 (N_6378,N_6030,N_5581);
nand U6379 (N_6379,N_5985,N_6196);
nand U6380 (N_6380,N_6104,N_5791);
nor U6381 (N_6381,N_5442,N_5651);
and U6382 (N_6382,N_5597,N_6066);
or U6383 (N_6383,N_5679,N_5397);
xor U6384 (N_6384,N_6197,N_5606);
or U6385 (N_6385,N_5332,N_5320);
xor U6386 (N_6386,N_6113,N_5274);
nor U6387 (N_6387,N_5523,N_6095);
and U6388 (N_6388,N_5110,N_5634);
xnor U6389 (N_6389,N_5136,N_5652);
xor U6390 (N_6390,N_5234,N_5358);
or U6391 (N_6391,N_5567,N_5424);
xor U6392 (N_6392,N_5206,N_5015);
nand U6393 (N_6393,N_5750,N_6105);
nor U6394 (N_6394,N_5408,N_5940);
nor U6395 (N_6395,N_5421,N_6195);
xor U6396 (N_6396,N_6077,N_5043);
or U6397 (N_6397,N_5636,N_5484);
nand U6398 (N_6398,N_5997,N_5214);
nand U6399 (N_6399,N_5179,N_5493);
and U6400 (N_6400,N_5734,N_6235);
xor U6401 (N_6401,N_5209,N_5727);
or U6402 (N_6402,N_5125,N_6246);
or U6403 (N_6403,N_5453,N_6238);
or U6404 (N_6404,N_5022,N_6059);
and U6405 (N_6405,N_5642,N_6191);
xnor U6406 (N_6406,N_6070,N_5893);
nor U6407 (N_6407,N_5552,N_5140);
nand U6408 (N_6408,N_6145,N_5454);
nor U6409 (N_6409,N_5126,N_6111);
nor U6410 (N_6410,N_5811,N_5194);
xnor U6411 (N_6411,N_5685,N_5122);
xor U6412 (N_6412,N_5178,N_5781);
and U6413 (N_6413,N_5680,N_6240);
xor U6414 (N_6414,N_5891,N_5663);
xnor U6415 (N_6415,N_6069,N_6129);
or U6416 (N_6416,N_5900,N_5903);
nor U6417 (N_6417,N_6008,N_5074);
or U6418 (N_6418,N_5177,N_6037);
nand U6419 (N_6419,N_5856,N_5227);
nor U6420 (N_6420,N_5447,N_5153);
or U6421 (N_6421,N_5482,N_5360);
nor U6422 (N_6422,N_6093,N_6175);
nand U6423 (N_6423,N_5065,N_5535);
xnor U6424 (N_6424,N_5335,N_5693);
nand U6425 (N_6425,N_5236,N_5765);
and U6426 (N_6426,N_5952,N_5533);
xnor U6427 (N_6427,N_5124,N_6112);
xnor U6428 (N_6428,N_6029,N_5080);
and U6429 (N_6429,N_6213,N_5351);
nor U6430 (N_6430,N_5158,N_6202);
nand U6431 (N_6431,N_5676,N_6123);
and U6432 (N_6432,N_6006,N_5038);
and U6433 (N_6433,N_6052,N_5915);
nor U6434 (N_6434,N_5263,N_5648);
xor U6435 (N_6435,N_5834,N_5621);
or U6436 (N_6436,N_5129,N_6218);
nand U6437 (N_6437,N_6098,N_5488);
and U6438 (N_6438,N_5747,N_6102);
nor U6439 (N_6439,N_5912,N_6031);
nor U6440 (N_6440,N_5465,N_5866);
xnor U6441 (N_6441,N_5926,N_6161);
and U6442 (N_6442,N_5945,N_5923);
xor U6443 (N_6443,N_5391,N_5063);
and U6444 (N_6444,N_5495,N_6199);
nand U6445 (N_6445,N_5261,N_5011);
and U6446 (N_6446,N_5062,N_5744);
or U6447 (N_6447,N_5251,N_5240);
nand U6448 (N_6448,N_5133,N_6036);
nand U6449 (N_6449,N_6046,N_5427);
and U6450 (N_6450,N_5455,N_5055);
or U6451 (N_6451,N_6223,N_5436);
and U6452 (N_6452,N_5520,N_5752);
nand U6453 (N_6453,N_5069,N_6044);
nand U6454 (N_6454,N_5524,N_5438);
and U6455 (N_6455,N_5483,N_5884);
xnor U6456 (N_6456,N_6000,N_6171);
nand U6457 (N_6457,N_5967,N_5880);
xor U6458 (N_6458,N_5982,N_5612);
or U6459 (N_6459,N_6138,N_5476);
nand U6460 (N_6460,N_5247,N_5502);
nand U6461 (N_6461,N_6016,N_6174);
and U6462 (N_6462,N_5528,N_5630);
or U6463 (N_6463,N_5718,N_5832);
or U6464 (N_6464,N_5383,N_5874);
and U6465 (N_6465,N_6229,N_5615);
nand U6466 (N_6466,N_5737,N_5035);
xor U6467 (N_6467,N_6023,N_5805);
or U6468 (N_6468,N_6237,N_5143);
nor U6469 (N_6469,N_5312,N_5961);
xnor U6470 (N_6470,N_5202,N_5778);
xnor U6471 (N_6471,N_5345,N_6118);
nor U6472 (N_6472,N_5729,N_5704);
xnor U6473 (N_6473,N_5404,N_6110);
and U6474 (N_6474,N_5835,N_5701);
nand U6475 (N_6475,N_5283,N_5083);
xor U6476 (N_6476,N_5699,N_5825);
or U6477 (N_6477,N_5941,N_5824);
nor U6478 (N_6478,N_5613,N_5434);
nor U6479 (N_6479,N_5890,N_5025);
and U6480 (N_6480,N_5864,N_5595);
nor U6481 (N_6481,N_5019,N_5183);
and U6482 (N_6482,N_6241,N_5922);
nand U6483 (N_6483,N_5583,N_5441);
nand U6484 (N_6484,N_5851,N_6163);
nor U6485 (N_6485,N_6053,N_5871);
nand U6486 (N_6486,N_5220,N_5398);
nor U6487 (N_6487,N_5382,N_5392);
or U6488 (N_6488,N_5764,N_5669);
xor U6489 (N_6489,N_5371,N_5407);
xor U6490 (N_6490,N_5992,N_6043);
nor U6491 (N_6491,N_5793,N_6060);
nor U6492 (N_6492,N_5831,N_5598);
nor U6493 (N_6493,N_5882,N_5486);
xnor U6494 (N_6494,N_5356,N_5932);
and U6495 (N_6495,N_5766,N_5668);
and U6496 (N_6496,N_6244,N_5694);
nor U6497 (N_6497,N_5803,N_6032);
nand U6498 (N_6498,N_5078,N_5710);
or U6499 (N_6499,N_5412,N_5213);
xor U6500 (N_6500,N_5981,N_6160);
xor U6501 (N_6501,N_5132,N_5867);
or U6502 (N_6502,N_5850,N_5958);
xor U6503 (N_6503,N_6205,N_5588);
and U6504 (N_6504,N_5841,N_5641);
and U6505 (N_6505,N_5317,N_5352);
nand U6506 (N_6506,N_5948,N_5467);
nor U6507 (N_6507,N_6230,N_5205);
nor U6508 (N_6508,N_6247,N_5008);
and U6509 (N_6509,N_5714,N_5323);
or U6510 (N_6510,N_5337,N_5272);
xor U6511 (N_6511,N_5067,N_6176);
or U6512 (N_6512,N_5724,N_6040);
and U6513 (N_6513,N_6106,N_5715);
and U6514 (N_6514,N_5417,N_6221);
nand U6515 (N_6515,N_6135,N_6187);
nor U6516 (N_6516,N_5270,N_6180);
and U6517 (N_6517,N_5949,N_5716);
nand U6518 (N_6518,N_5559,N_5754);
nor U6519 (N_6519,N_5684,N_5366);
and U6520 (N_6520,N_5999,N_5030);
nor U6521 (N_6521,N_5119,N_5445);
nand U6522 (N_6522,N_5643,N_5580);
nor U6523 (N_6523,N_5156,N_5023);
nor U6524 (N_6524,N_5107,N_5388);
nor U6525 (N_6525,N_5207,N_5756);
nor U6526 (N_6526,N_6172,N_5487);
xnor U6527 (N_6527,N_5840,N_5142);
nor U6528 (N_6528,N_5736,N_5235);
and U6529 (N_6529,N_5713,N_6122);
nand U6530 (N_6530,N_6233,N_5833);
and U6531 (N_6531,N_5647,N_6165);
nand U6532 (N_6532,N_5931,N_5527);
nor U6533 (N_6533,N_5089,N_5632);
nand U6534 (N_6534,N_5644,N_5863);
and U6535 (N_6535,N_5373,N_6215);
or U6536 (N_6536,N_6146,N_5481);
and U6537 (N_6537,N_5549,N_5700);
or U6538 (N_6538,N_5384,N_6020);
and U6539 (N_6539,N_5459,N_5698);
nor U6540 (N_6540,N_5599,N_5818);
xor U6541 (N_6541,N_5814,N_6167);
or U6542 (N_6542,N_5705,N_5114);
nor U6543 (N_6543,N_6245,N_5497);
xnor U6544 (N_6544,N_5742,N_5927);
xor U6545 (N_6545,N_5809,N_5460);
and U6546 (N_6546,N_5921,N_5860);
nor U6547 (N_6547,N_5042,N_6155);
xnor U6548 (N_6548,N_5896,N_5422);
and U6549 (N_6549,N_5248,N_6074);
nand U6550 (N_6550,N_5002,N_5357);
and U6551 (N_6551,N_5013,N_5806);
or U6552 (N_6552,N_5197,N_5295);
or U6553 (N_6553,N_5800,N_5299);
and U6554 (N_6554,N_5432,N_5403);
and U6555 (N_6555,N_6068,N_5522);
nor U6556 (N_6556,N_5291,N_5186);
and U6557 (N_6557,N_5526,N_5416);
and U6558 (N_6558,N_5399,N_5976);
or U6559 (N_6559,N_6096,N_6173);
or U6560 (N_6560,N_6061,N_5324);
nor U6561 (N_6561,N_5285,N_5298);
nand U6562 (N_6562,N_5823,N_5152);
xnor U6563 (N_6563,N_5719,N_5380);
and U6564 (N_6564,N_5688,N_5007);
or U6565 (N_6565,N_5649,N_5331);
nand U6566 (N_6566,N_5284,N_5645);
and U6567 (N_6567,N_5917,N_5938);
or U6568 (N_6568,N_5032,N_5254);
and U6569 (N_6569,N_5000,N_5740);
nand U6570 (N_6570,N_5231,N_6204);
and U6571 (N_6571,N_5026,N_5692);
xnor U6572 (N_6572,N_5596,N_6057);
nand U6573 (N_6573,N_5771,N_5273);
xor U6574 (N_6574,N_6125,N_5913);
xor U6575 (N_6575,N_5379,N_5310);
nand U6576 (N_6576,N_5521,N_5293);
and U6577 (N_6577,N_5396,N_5775);
nor U6578 (N_6578,N_5974,N_5905);
xor U6579 (N_6579,N_5354,N_6140);
xnor U6580 (N_6580,N_5813,N_6164);
and U6581 (N_6581,N_6085,N_5996);
nand U6582 (N_6582,N_6075,N_5212);
and U6583 (N_6583,N_6072,N_5503);
nand U6584 (N_6584,N_5687,N_5309);
nor U6585 (N_6585,N_6114,N_5362);
nor U6586 (N_6586,N_5571,N_5797);
nor U6587 (N_6587,N_5150,N_5609);
or U6588 (N_6588,N_5009,N_5463);
nand U6589 (N_6589,N_5333,N_5650);
nor U6590 (N_6590,N_5113,N_6038);
or U6591 (N_6591,N_5768,N_5555);
nand U6592 (N_6592,N_5519,N_5859);
nor U6593 (N_6593,N_5873,N_6224);
or U6594 (N_6594,N_5906,N_6203);
nor U6595 (N_6595,N_5444,N_5822);
xnor U6596 (N_6596,N_5141,N_5148);
or U6597 (N_6597,N_5208,N_5155);
or U6598 (N_6598,N_5633,N_5256);
nor U6599 (N_6599,N_5259,N_5784);
nand U6600 (N_6600,N_5279,N_5629);
nor U6601 (N_6601,N_5498,N_5457);
or U6602 (N_6602,N_5064,N_5798);
and U6603 (N_6603,N_5192,N_5659);
and U6604 (N_6604,N_5536,N_5049);
nor U6605 (N_6605,N_6024,N_5600);
nor U6606 (N_6606,N_5779,N_6033);
and U6607 (N_6607,N_5440,N_5500);
xnor U6608 (N_6608,N_6011,N_5703);
nor U6609 (N_6609,N_5792,N_5815);
nand U6610 (N_6610,N_5021,N_5959);
xor U6611 (N_6611,N_5977,N_5807);
nand U6612 (N_6612,N_5733,N_5246);
nand U6613 (N_6613,N_6025,N_5889);
xor U6614 (N_6614,N_5862,N_5387);
xor U6615 (N_6615,N_5829,N_5638);
nand U6616 (N_6616,N_6116,N_5052);
and U6617 (N_6617,N_5709,N_5879);
nor U6618 (N_6618,N_6100,N_5826);
nand U6619 (N_6619,N_6124,N_5475);
and U6620 (N_6620,N_5674,N_5330);
xor U6621 (N_6621,N_5004,N_5131);
and U6622 (N_6622,N_6131,N_6222);
nor U6623 (N_6623,N_5300,N_6178);
nand U6624 (N_6624,N_5204,N_5461);
nand U6625 (N_6625,N_5513,N_5265);
and U6626 (N_6626,N_5165,N_5368);
nand U6627 (N_6627,N_5820,N_5790);
nor U6628 (N_6628,N_5071,N_5314);
and U6629 (N_6629,N_5722,N_5059);
xnor U6630 (N_6630,N_5799,N_5640);
and U6631 (N_6631,N_5933,N_5405);
xor U6632 (N_6632,N_5169,N_5504);
xnor U6633 (N_6633,N_5802,N_5842);
or U6634 (N_6634,N_5639,N_6152);
or U6635 (N_6635,N_5956,N_5963);
xnor U6636 (N_6636,N_5229,N_6058);
nand U6637 (N_6637,N_6005,N_5839);
nand U6638 (N_6638,N_5628,N_5086);
nand U6639 (N_6639,N_5557,N_5127);
nor U6640 (N_6640,N_5936,N_5849);
and U6641 (N_6641,N_5876,N_6243);
and U6642 (N_6642,N_5033,N_5707);
nor U6643 (N_6643,N_5553,N_5419);
nand U6644 (N_6644,N_5610,N_5328);
nand U6645 (N_6645,N_5494,N_5783);
or U6646 (N_6646,N_5881,N_5449);
or U6647 (N_6647,N_6018,N_5902);
nand U6648 (N_6648,N_5723,N_5319);
nor U6649 (N_6649,N_5712,N_5370);
nand U6650 (N_6650,N_5539,N_5594);
xnor U6651 (N_6651,N_5016,N_6079);
xor U6652 (N_6652,N_5187,N_5960);
or U6653 (N_6653,N_5448,N_6136);
xnor U6654 (N_6654,N_5726,N_5109);
nor U6655 (N_6655,N_5678,N_5350);
xnor U6656 (N_6656,N_5545,N_6183);
and U6657 (N_6657,N_6090,N_6083);
nor U6658 (N_6658,N_6003,N_5776);
xnor U6659 (N_6659,N_5469,N_5837);
nor U6660 (N_6660,N_5222,N_5804);
or U6661 (N_6661,N_6126,N_5393);
or U6662 (N_6662,N_6028,N_5301);
and U6663 (N_6663,N_5420,N_5918);
xnor U6664 (N_6664,N_6054,N_5541);
nor U6665 (N_6665,N_5462,N_6101);
nand U6666 (N_6666,N_6201,N_6200);
and U6667 (N_6667,N_5017,N_6162);
or U6668 (N_6668,N_5836,N_6091);
and U6669 (N_6669,N_5556,N_5238);
nand U6670 (N_6670,N_5245,N_5018);
xor U6671 (N_6671,N_5509,N_5794);
nor U6672 (N_6672,N_5100,N_5147);
nand U6673 (N_6673,N_5414,N_5550);
xor U6674 (N_6674,N_6010,N_5359);
xor U6675 (N_6675,N_6050,N_5340);
or U6676 (N_6676,N_5188,N_5296);
nand U6677 (N_6677,N_5492,N_6151);
or U6678 (N_6678,N_5289,N_5789);
or U6679 (N_6679,N_5877,N_5591);
and U6680 (N_6680,N_5819,N_5121);
nand U6681 (N_6681,N_5817,N_5066);
or U6682 (N_6682,N_5725,N_5344);
or U6683 (N_6683,N_5929,N_5998);
or U6684 (N_6684,N_5474,N_6141);
and U6685 (N_6685,N_5406,N_5191);
or U6686 (N_6686,N_5386,N_5885);
xor U6687 (N_6687,N_5894,N_5763);
nor U6688 (N_6688,N_6207,N_5654);
nor U6689 (N_6689,N_6067,N_6133);
nand U6690 (N_6690,N_6027,N_5518);
nand U6691 (N_6691,N_5774,N_5269);
and U6692 (N_6692,N_5830,N_5816);
or U6693 (N_6693,N_6184,N_5276);
or U6694 (N_6694,N_5425,N_5909);
xnor U6695 (N_6695,N_5308,N_5243);
xnor U6696 (N_6696,N_5966,N_5171);
nand U6697 (N_6697,N_5346,N_5070);
or U6698 (N_6698,N_5755,N_5145);
nand U6699 (N_6699,N_5878,N_5590);
nor U6700 (N_6700,N_5511,N_6002);
and U6701 (N_6701,N_5375,N_5489);
or U6702 (N_6702,N_5266,N_5968);
or U6703 (N_6703,N_5363,N_5762);
nand U6704 (N_6704,N_5542,N_5657);
nor U6705 (N_6705,N_6193,N_5772);
nor U6706 (N_6706,N_5843,N_5437);
and U6707 (N_6707,N_5531,N_5666);
or U6708 (N_6708,N_5185,N_5166);
and U6709 (N_6709,N_5604,N_5369);
nand U6710 (N_6710,N_5720,N_5292);
xnor U6711 (N_6711,N_6192,N_5951);
xnor U6712 (N_6712,N_6150,N_5847);
and U6713 (N_6713,N_5573,N_5037);
nor U6714 (N_6714,N_5954,N_5161);
nand U6715 (N_6715,N_5886,N_5578);
or U6716 (N_6716,N_6186,N_5201);
nor U6717 (N_6717,N_5082,N_5264);
nand U6718 (N_6718,N_5758,N_5984);
nor U6719 (N_6719,N_5626,N_6121);
and U6720 (N_6720,N_5061,N_6088);
xor U6721 (N_6721,N_5658,N_5760);
nand U6722 (N_6722,N_5381,N_5625);
nand U6723 (N_6723,N_5569,N_6158);
nand U6724 (N_6724,N_5175,N_5277);
and U6725 (N_6725,N_5517,N_5347);
nor U6726 (N_6726,N_5869,N_5980);
nor U6727 (N_6727,N_5176,N_5608);
or U6728 (N_6728,N_5564,N_5853);
nor U6729 (N_6729,N_5267,N_5389);
nor U6730 (N_6730,N_6047,N_5962);
nand U6731 (N_6731,N_5670,N_5028);
or U6732 (N_6732,N_5123,N_5230);
and U6733 (N_6733,N_5268,N_5942);
xor U6734 (N_6734,N_5558,N_5955);
nand U6735 (N_6735,N_5844,N_5689);
nor U6736 (N_6736,N_6063,N_6084);
xor U6737 (N_6737,N_5096,N_5686);
or U6738 (N_6738,N_5410,N_5586);
xnor U6739 (N_6739,N_5087,N_5611);
and U6740 (N_6740,N_6169,N_5305);
nand U6741 (N_6741,N_5702,N_6076);
nand U6742 (N_6742,N_5671,N_5306);
nand U6743 (N_6743,N_5761,N_6013);
nor U6744 (N_6744,N_5582,N_5180);
nand U6745 (N_6745,N_5901,N_5655);
nand U6746 (N_6746,N_5402,N_5472);
and U6747 (N_6747,N_5058,N_5464);
nand U6748 (N_6748,N_6227,N_5711);
xnor U6749 (N_6749,N_5241,N_5253);
and U6750 (N_6750,N_5584,N_5036);
and U6751 (N_6751,N_5144,N_5451);
and U6752 (N_6752,N_5983,N_6154);
xnor U6753 (N_6753,N_5995,N_6220);
xnor U6754 (N_6754,N_5372,N_5297);
nor U6755 (N_6755,N_5341,N_5661);
or U6756 (N_6756,N_5516,N_5242);
nor U6757 (N_6757,N_5505,N_5934);
and U6758 (N_6758,N_5088,N_5151);
nor U6759 (N_6759,N_5937,N_6179);
or U6760 (N_6760,N_6051,N_5395);
nor U6761 (N_6761,N_5218,N_5631);
xnor U6762 (N_6762,N_5857,N_5827);
and U6763 (N_6763,N_5575,N_5390);
nand U6764 (N_6764,N_5005,N_5782);
or U6765 (N_6765,N_5677,N_5138);
or U6766 (N_6766,N_5128,N_5217);
nand U6767 (N_6767,N_5935,N_5529);
and U6768 (N_6768,N_6045,N_5855);
xnor U6769 (N_6769,N_5200,N_5024);
xnor U6770 (N_6770,N_5134,N_5751);
and U6771 (N_6771,N_5311,N_6209);
or U6772 (N_6772,N_5342,N_6120);
nor U6773 (N_6773,N_6109,N_5233);
and U6774 (N_6774,N_5271,N_5478);
nand U6775 (N_6775,N_5928,N_5895);
nor U6776 (N_6776,N_5624,N_5473);
xnor U6777 (N_6777,N_5287,N_6103);
nor U6778 (N_6778,N_5662,N_5515);
xnor U6779 (N_6779,N_5223,N_5443);
or U6780 (N_6780,N_5101,N_6168);
nor U6781 (N_6781,N_5490,N_5560);
nor U6782 (N_6782,N_5111,N_5745);
nand U6783 (N_6783,N_5189,N_6137);
nor U6784 (N_6784,N_5861,N_5987);
nand U6785 (N_6785,N_5433,N_5115);
xnor U6786 (N_6786,N_5537,N_5446);
and U6787 (N_6787,N_6001,N_5538);
and U6788 (N_6788,N_5068,N_5120);
xor U6789 (N_6789,N_5975,N_5697);
and U6790 (N_6790,N_5892,N_5411);
nor U6791 (N_6791,N_6128,N_5057);
nor U6792 (N_6792,N_6071,N_5094);
nor U6793 (N_6793,N_5656,N_6148);
xnor U6794 (N_6794,N_5006,N_5288);
or U6795 (N_6795,N_5510,N_5117);
nand U6796 (N_6796,N_5260,N_6177);
or U6797 (N_6797,N_6014,N_5969);
nand U6798 (N_6798,N_6080,N_5943);
and U6799 (N_6799,N_5619,N_5039);
xnor U6800 (N_6800,N_5769,N_5675);
or U6801 (N_6801,N_5322,N_5092);
nor U6802 (N_6802,N_6211,N_5244);
nand U6803 (N_6803,N_5919,N_5623);
and U6804 (N_6804,N_5470,N_5304);
xnor U6805 (N_6805,N_5321,N_5563);
nor U6806 (N_6806,N_6081,N_5374);
xnor U6807 (N_6807,N_5456,N_5452);
xor U6808 (N_6808,N_5315,N_5400);
nor U6809 (N_6809,N_5139,N_5506);
nor U6810 (N_6810,N_5435,N_5607);
nor U6811 (N_6811,N_5290,N_5672);
nor U6812 (N_6812,N_5858,N_6198);
and U6813 (N_6813,N_5731,N_5095);
nor U6814 (N_6814,N_5116,N_6086);
or U6815 (N_6815,N_5989,N_5741);
nor U6816 (N_6816,N_5910,N_5361);
and U6817 (N_6817,N_5048,N_5717);
xor U6818 (N_6818,N_5195,N_5979);
or U6819 (N_6819,N_5898,N_5872);
xor U6820 (N_6820,N_6232,N_5883);
and U6821 (N_6821,N_5262,N_5501);
and U6822 (N_6822,N_6228,N_5845);
or U6823 (N_6823,N_5691,N_5875);
nor U6824 (N_6824,N_5430,N_5339);
nor U6825 (N_6825,N_5854,N_5770);
and U6826 (N_6826,N_6117,N_5665);
xnor U6827 (N_6827,N_5480,N_5993);
or U6828 (N_6828,N_5868,N_5801);
and U6829 (N_6829,N_5413,N_5812);
or U6830 (N_6830,N_5182,N_5294);
and U6831 (N_6831,N_5739,N_5237);
nor U6832 (N_6832,N_5646,N_5198);
nand U6833 (N_6833,N_6236,N_6157);
nand U6834 (N_6834,N_5278,N_5735);
nand U6835 (N_6835,N_6094,N_5828);
or U6836 (N_6836,N_5551,N_5603);
and U6837 (N_6837,N_5307,N_6219);
and U6838 (N_6838,N_5003,N_6127);
and U6839 (N_6839,N_5102,N_5796);
xor U6840 (N_6840,N_5012,N_6039);
or U6841 (N_6841,N_5964,N_5916);
nand U6842 (N_6842,N_5184,N_6194);
xor U6843 (N_6843,N_5988,N_5683);
xor U6844 (N_6844,N_5203,N_5001);
nor U6845 (N_6845,N_5401,N_6149);
nand U6846 (N_6846,N_6147,N_5622);
or U6847 (N_6847,N_5757,N_6217);
xnor U6848 (N_6848,N_5592,N_5255);
xnor U6849 (N_6849,N_5349,N_5749);
xnor U6850 (N_6850,N_6181,N_5196);
or U6851 (N_6851,N_5031,N_5172);
or U6852 (N_6852,N_5439,N_5418);
or U6853 (N_6853,N_5163,N_5099);
nand U6854 (N_6854,N_5365,N_5302);
nand U6855 (N_6855,N_6041,N_6092);
and U6856 (N_6856,N_5870,N_5160);
nor U6857 (N_6857,N_5730,N_5050);
xor U6858 (N_6858,N_5325,N_5477);
or U6859 (N_6859,N_5364,N_5027);
and U6860 (N_6860,N_5566,N_6248);
nor U6861 (N_6861,N_6153,N_5355);
nand U6862 (N_6862,N_5773,N_5546);
nor U6863 (N_6863,N_5978,N_5105);
nor U6864 (N_6864,N_5795,N_5924);
nor U6865 (N_6865,N_6004,N_5605);
xor U6866 (N_6866,N_6226,N_6242);
xnor U6867 (N_6867,N_5053,N_5168);
and U6868 (N_6868,N_6015,N_5572);
and U6869 (N_6869,N_5971,N_6012);
or U6870 (N_6870,N_5627,N_5221);
or U6871 (N_6871,N_5759,N_5060);
or U6872 (N_6872,N_5106,N_5093);
xnor U6873 (N_6873,N_5821,N_5377);
nor U6874 (N_6874,N_5512,N_5925);
nor U6875 (N_6875,N_6102,N_5253);
nor U6876 (N_6876,N_6014,N_5445);
or U6877 (N_6877,N_5440,N_5493);
xnor U6878 (N_6878,N_5937,N_5985);
and U6879 (N_6879,N_6223,N_6106);
nand U6880 (N_6880,N_5817,N_5084);
or U6881 (N_6881,N_6106,N_5295);
nand U6882 (N_6882,N_5265,N_5780);
xor U6883 (N_6883,N_5985,N_5815);
and U6884 (N_6884,N_5215,N_5015);
and U6885 (N_6885,N_5992,N_5518);
nand U6886 (N_6886,N_5303,N_5803);
nor U6887 (N_6887,N_5060,N_5063);
xnor U6888 (N_6888,N_5506,N_5464);
and U6889 (N_6889,N_5907,N_6249);
nor U6890 (N_6890,N_5852,N_5824);
and U6891 (N_6891,N_5978,N_5098);
and U6892 (N_6892,N_5184,N_5943);
and U6893 (N_6893,N_5253,N_5205);
nand U6894 (N_6894,N_5753,N_6130);
xnor U6895 (N_6895,N_5432,N_5730);
xnor U6896 (N_6896,N_5048,N_6174);
nor U6897 (N_6897,N_5670,N_5402);
nor U6898 (N_6898,N_5268,N_6204);
and U6899 (N_6899,N_5331,N_5318);
nor U6900 (N_6900,N_5253,N_5482);
or U6901 (N_6901,N_5380,N_5015);
xor U6902 (N_6902,N_5233,N_6086);
xnor U6903 (N_6903,N_5932,N_5589);
and U6904 (N_6904,N_5402,N_6039);
xnor U6905 (N_6905,N_6222,N_5331);
or U6906 (N_6906,N_5625,N_5252);
nor U6907 (N_6907,N_5206,N_5820);
and U6908 (N_6908,N_5989,N_5077);
nor U6909 (N_6909,N_5887,N_5051);
and U6910 (N_6910,N_5034,N_5070);
nor U6911 (N_6911,N_6210,N_5945);
nor U6912 (N_6912,N_5859,N_5792);
nor U6913 (N_6913,N_5807,N_5226);
nor U6914 (N_6914,N_6229,N_5192);
nand U6915 (N_6915,N_5083,N_6092);
nor U6916 (N_6916,N_5370,N_5179);
xnor U6917 (N_6917,N_6068,N_5356);
or U6918 (N_6918,N_5134,N_5512);
and U6919 (N_6919,N_5335,N_5442);
nand U6920 (N_6920,N_5663,N_5491);
and U6921 (N_6921,N_5928,N_5260);
nand U6922 (N_6922,N_5084,N_5682);
nand U6923 (N_6923,N_5069,N_5914);
nor U6924 (N_6924,N_5708,N_5327);
nand U6925 (N_6925,N_5938,N_5666);
xor U6926 (N_6926,N_5425,N_5605);
xnor U6927 (N_6927,N_5885,N_6213);
or U6928 (N_6928,N_5453,N_5320);
xor U6929 (N_6929,N_6012,N_6157);
nor U6930 (N_6930,N_5651,N_6147);
and U6931 (N_6931,N_5114,N_5319);
nor U6932 (N_6932,N_5727,N_5688);
xor U6933 (N_6933,N_5337,N_5176);
nor U6934 (N_6934,N_5443,N_5477);
nor U6935 (N_6935,N_5285,N_6192);
nand U6936 (N_6936,N_5350,N_5961);
xor U6937 (N_6937,N_5160,N_5100);
xor U6938 (N_6938,N_5018,N_6109);
xnor U6939 (N_6939,N_5258,N_5765);
nand U6940 (N_6940,N_5192,N_5479);
nor U6941 (N_6941,N_5168,N_5676);
nor U6942 (N_6942,N_5597,N_5593);
and U6943 (N_6943,N_5476,N_5113);
xnor U6944 (N_6944,N_5613,N_5707);
xor U6945 (N_6945,N_5180,N_5524);
nand U6946 (N_6946,N_5154,N_6183);
xor U6947 (N_6947,N_6224,N_5148);
xnor U6948 (N_6948,N_5903,N_6085);
and U6949 (N_6949,N_6014,N_5554);
nor U6950 (N_6950,N_6094,N_6138);
or U6951 (N_6951,N_5924,N_6068);
or U6952 (N_6952,N_5427,N_5454);
nor U6953 (N_6953,N_6010,N_5003);
nand U6954 (N_6954,N_6148,N_6209);
nor U6955 (N_6955,N_5693,N_5537);
nand U6956 (N_6956,N_5696,N_5524);
or U6957 (N_6957,N_5386,N_5992);
and U6958 (N_6958,N_5660,N_5626);
nand U6959 (N_6959,N_5700,N_5818);
nand U6960 (N_6960,N_5210,N_5966);
nand U6961 (N_6961,N_5641,N_5898);
xnor U6962 (N_6962,N_6131,N_5143);
xnor U6963 (N_6963,N_5344,N_6154);
and U6964 (N_6964,N_6072,N_5157);
or U6965 (N_6965,N_5220,N_5888);
and U6966 (N_6966,N_5417,N_6030);
or U6967 (N_6967,N_5137,N_6179);
nand U6968 (N_6968,N_5636,N_5113);
nand U6969 (N_6969,N_5747,N_5132);
nand U6970 (N_6970,N_5534,N_5761);
and U6971 (N_6971,N_6076,N_6194);
nor U6972 (N_6972,N_5894,N_5851);
xnor U6973 (N_6973,N_5265,N_5469);
or U6974 (N_6974,N_5697,N_5193);
nand U6975 (N_6975,N_5342,N_5722);
xnor U6976 (N_6976,N_5463,N_5313);
and U6977 (N_6977,N_5897,N_6014);
xor U6978 (N_6978,N_5687,N_5004);
nor U6979 (N_6979,N_6231,N_5363);
and U6980 (N_6980,N_6205,N_5423);
nor U6981 (N_6981,N_5795,N_5031);
and U6982 (N_6982,N_5087,N_5267);
xnor U6983 (N_6983,N_5400,N_5245);
nor U6984 (N_6984,N_5999,N_5648);
xnor U6985 (N_6985,N_5637,N_5050);
xnor U6986 (N_6986,N_5261,N_5368);
xnor U6987 (N_6987,N_5590,N_6235);
nor U6988 (N_6988,N_5210,N_5663);
nor U6989 (N_6989,N_5257,N_6038);
nor U6990 (N_6990,N_5238,N_6217);
nand U6991 (N_6991,N_5317,N_5915);
nor U6992 (N_6992,N_5641,N_5305);
nand U6993 (N_6993,N_6129,N_5766);
and U6994 (N_6994,N_5591,N_6041);
nor U6995 (N_6995,N_5817,N_5070);
nand U6996 (N_6996,N_5373,N_5116);
nand U6997 (N_6997,N_5015,N_6204);
and U6998 (N_6998,N_5908,N_5925);
nand U6999 (N_6999,N_5036,N_5740);
or U7000 (N_7000,N_5393,N_5430);
xor U7001 (N_7001,N_5800,N_5054);
xnor U7002 (N_7002,N_5597,N_5169);
xnor U7003 (N_7003,N_5574,N_5671);
and U7004 (N_7004,N_6190,N_5872);
nand U7005 (N_7005,N_5911,N_5524);
nor U7006 (N_7006,N_5009,N_5744);
and U7007 (N_7007,N_6210,N_5324);
xor U7008 (N_7008,N_6234,N_5886);
nor U7009 (N_7009,N_5436,N_5234);
nor U7010 (N_7010,N_5862,N_5562);
nor U7011 (N_7011,N_6029,N_5464);
nand U7012 (N_7012,N_5034,N_6005);
nor U7013 (N_7013,N_5654,N_5992);
nand U7014 (N_7014,N_6190,N_5123);
and U7015 (N_7015,N_5536,N_5976);
nand U7016 (N_7016,N_6084,N_5170);
and U7017 (N_7017,N_6093,N_6238);
xnor U7018 (N_7018,N_5942,N_5410);
and U7019 (N_7019,N_6176,N_5780);
nor U7020 (N_7020,N_5500,N_5394);
xor U7021 (N_7021,N_5801,N_5462);
nor U7022 (N_7022,N_5079,N_5653);
nand U7023 (N_7023,N_5710,N_5937);
xnor U7024 (N_7024,N_5951,N_5978);
nor U7025 (N_7025,N_5514,N_5897);
nor U7026 (N_7026,N_5571,N_5052);
nand U7027 (N_7027,N_5834,N_5669);
nor U7028 (N_7028,N_5767,N_6027);
and U7029 (N_7029,N_5421,N_5153);
and U7030 (N_7030,N_6227,N_5788);
nand U7031 (N_7031,N_5500,N_5324);
xnor U7032 (N_7032,N_5218,N_5791);
or U7033 (N_7033,N_5711,N_5219);
xnor U7034 (N_7034,N_6106,N_5475);
and U7035 (N_7035,N_5491,N_5594);
or U7036 (N_7036,N_5702,N_5209);
nand U7037 (N_7037,N_5842,N_5584);
and U7038 (N_7038,N_5286,N_6102);
and U7039 (N_7039,N_6068,N_5488);
nand U7040 (N_7040,N_5848,N_5585);
nor U7041 (N_7041,N_6182,N_5409);
nand U7042 (N_7042,N_5595,N_5608);
nor U7043 (N_7043,N_5664,N_5636);
nand U7044 (N_7044,N_5705,N_5948);
or U7045 (N_7045,N_5978,N_5300);
nor U7046 (N_7046,N_5760,N_5803);
and U7047 (N_7047,N_5112,N_6181);
and U7048 (N_7048,N_5313,N_5454);
xor U7049 (N_7049,N_5054,N_5981);
or U7050 (N_7050,N_5004,N_6114);
or U7051 (N_7051,N_6198,N_5063);
xor U7052 (N_7052,N_5313,N_5385);
nor U7053 (N_7053,N_5599,N_5022);
nor U7054 (N_7054,N_5235,N_5450);
or U7055 (N_7055,N_5257,N_6141);
nand U7056 (N_7056,N_5962,N_6104);
and U7057 (N_7057,N_5752,N_5367);
nor U7058 (N_7058,N_6218,N_5250);
xor U7059 (N_7059,N_5840,N_5564);
xnor U7060 (N_7060,N_5684,N_5769);
and U7061 (N_7061,N_5410,N_6101);
xor U7062 (N_7062,N_5233,N_5380);
and U7063 (N_7063,N_5192,N_5270);
and U7064 (N_7064,N_5748,N_6228);
nand U7065 (N_7065,N_5022,N_5707);
nor U7066 (N_7066,N_6148,N_5809);
xor U7067 (N_7067,N_5830,N_6078);
nor U7068 (N_7068,N_5386,N_6239);
and U7069 (N_7069,N_6222,N_5644);
xor U7070 (N_7070,N_5006,N_5039);
or U7071 (N_7071,N_6177,N_6171);
nand U7072 (N_7072,N_5838,N_5813);
nor U7073 (N_7073,N_5339,N_5222);
nand U7074 (N_7074,N_5658,N_5114);
nor U7075 (N_7075,N_5827,N_5983);
and U7076 (N_7076,N_5127,N_5014);
and U7077 (N_7077,N_5141,N_5193);
nor U7078 (N_7078,N_5510,N_6114);
xnor U7079 (N_7079,N_6054,N_5443);
or U7080 (N_7080,N_5435,N_5564);
and U7081 (N_7081,N_6117,N_5649);
or U7082 (N_7082,N_5030,N_5944);
or U7083 (N_7083,N_5337,N_5627);
and U7084 (N_7084,N_5657,N_5424);
nand U7085 (N_7085,N_5509,N_5040);
nand U7086 (N_7086,N_5067,N_5004);
and U7087 (N_7087,N_5665,N_5712);
nor U7088 (N_7088,N_5273,N_5311);
and U7089 (N_7089,N_5604,N_5635);
nor U7090 (N_7090,N_5164,N_5271);
and U7091 (N_7091,N_6022,N_5291);
and U7092 (N_7092,N_5001,N_5833);
and U7093 (N_7093,N_5996,N_5051);
or U7094 (N_7094,N_5428,N_5608);
nand U7095 (N_7095,N_5371,N_5157);
xor U7096 (N_7096,N_5987,N_6129);
xor U7097 (N_7097,N_6211,N_6089);
or U7098 (N_7098,N_5482,N_5195);
xnor U7099 (N_7099,N_5565,N_5342);
nand U7100 (N_7100,N_5207,N_6100);
nor U7101 (N_7101,N_5278,N_5445);
or U7102 (N_7102,N_6137,N_6132);
and U7103 (N_7103,N_5012,N_5719);
nor U7104 (N_7104,N_5996,N_5575);
or U7105 (N_7105,N_5445,N_5974);
xnor U7106 (N_7106,N_5414,N_5674);
and U7107 (N_7107,N_5345,N_5356);
nor U7108 (N_7108,N_5460,N_6117);
xor U7109 (N_7109,N_5257,N_5331);
nor U7110 (N_7110,N_6205,N_5639);
or U7111 (N_7111,N_6128,N_5692);
nand U7112 (N_7112,N_5504,N_6138);
nand U7113 (N_7113,N_5541,N_5778);
and U7114 (N_7114,N_5558,N_5521);
nand U7115 (N_7115,N_5594,N_5084);
nand U7116 (N_7116,N_5441,N_5423);
and U7117 (N_7117,N_5266,N_5558);
nor U7118 (N_7118,N_5394,N_5521);
and U7119 (N_7119,N_5512,N_5962);
or U7120 (N_7120,N_5938,N_6249);
nand U7121 (N_7121,N_5353,N_5723);
xor U7122 (N_7122,N_5108,N_5766);
nor U7123 (N_7123,N_5237,N_5573);
and U7124 (N_7124,N_5506,N_6154);
nor U7125 (N_7125,N_5884,N_5578);
nor U7126 (N_7126,N_5321,N_5212);
xnor U7127 (N_7127,N_5982,N_6161);
or U7128 (N_7128,N_5021,N_5746);
nand U7129 (N_7129,N_5504,N_5955);
and U7130 (N_7130,N_5997,N_5848);
nand U7131 (N_7131,N_6218,N_5360);
and U7132 (N_7132,N_5362,N_5346);
xor U7133 (N_7133,N_5752,N_5958);
nor U7134 (N_7134,N_6050,N_5053);
or U7135 (N_7135,N_6034,N_5637);
xor U7136 (N_7136,N_5688,N_6111);
or U7137 (N_7137,N_5357,N_5671);
nand U7138 (N_7138,N_6031,N_5913);
nor U7139 (N_7139,N_5465,N_5978);
xnor U7140 (N_7140,N_5384,N_5102);
xnor U7141 (N_7141,N_5289,N_6031);
xnor U7142 (N_7142,N_5724,N_5420);
or U7143 (N_7143,N_6065,N_6172);
xnor U7144 (N_7144,N_5176,N_5344);
or U7145 (N_7145,N_5021,N_5601);
xnor U7146 (N_7146,N_6056,N_5777);
or U7147 (N_7147,N_6097,N_5963);
or U7148 (N_7148,N_5305,N_5164);
nand U7149 (N_7149,N_5180,N_5256);
nand U7150 (N_7150,N_5525,N_6159);
nand U7151 (N_7151,N_6096,N_5627);
nor U7152 (N_7152,N_5086,N_5433);
nand U7153 (N_7153,N_5609,N_5176);
nand U7154 (N_7154,N_5906,N_5643);
nor U7155 (N_7155,N_5235,N_5924);
nor U7156 (N_7156,N_5453,N_6069);
nand U7157 (N_7157,N_6180,N_5259);
and U7158 (N_7158,N_5159,N_5747);
xnor U7159 (N_7159,N_5349,N_5776);
nand U7160 (N_7160,N_6098,N_5875);
nor U7161 (N_7161,N_5807,N_6061);
and U7162 (N_7162,N_6209,N_5550);
or U7163 (N_7163,N_5057,N_5823);
nor U7164 (N_7164,N_5775,N_5334);
or U7165 (N_7165,N_5325,N_6014);
and U7166 (N_7166,N_5056,N_5898);
nand U7167 (N_7167,N_5122,N_5576);
nor U7168 (N_7168,N_5847,N_5157);
or U7169 (N_7169,N_5182,N_5422);
and U7170 (N_7170,N_6008,N_6038);
and U7171 (N_7171,N_5784,N_6244);
nand U7172 (N_7172,N_5238,N_5542);
nand U7173 (N_7173,N_5092,N_5688);
nand U7174 (N_7174,N_5585,N_6224);
nor U7175 (N_7175,N_5013,N_5004);
nand U7176 (N_7176,N_5934,N_6239);
and U7177 (N_7177,N_5087,N_5663);
and U7178 (N_7178,N_6220,N_5090);
nor U7179 (N_7179,N_5990,N_5897);
nor U7180 (N_7180,N_5328,N_6147);
nand U7181 (N_7181,N_5651,N_5537);
nand U7182 (N_7182,N_5112,N_5388);
or U7183 (N_7183,N_5293,N_5673);
and U7184 (N_7184,N_5520,N_5158);
and U7185 (N_7185,N_5667,N_5470);
nor U7186 (N_7186,N_5417,N_5275);
nor U7187 (N_7187,N_6114,N_5609);
xnor U7188 (N_7188,N_5362,N_5021);
xnor U7189 (N_7189,N_6143,N_5217);
or U7190 (N_7190,N_5385,N_5474);
nand U7191 (N_7191,N_5221,N_6194);
or U7192 (N_7192,N_5063,N_5810);
nand U7193 (N_7193,N_5559,N_5657);
xnor U7194 (N_7194,N_5155,N_5106);
nand U7195 (N_7195,N_5409,N_5737);
or U7196 (N_7196,N_6206,N_6089);
xnor U7197 (N_7197,N_5058,N_5286);
nand U7198 (N_7198,N_5019,N_5057);
nor U7199 (N_7199,N_5944,N_6098);
nor U7200 (N_7200,N_5148,N_5822);
or U7201 (N_7201,N_5131,N_5716);
nor U7202 (N_7202,N_6146,N_5094);
or U7203 (N_7203,N_5565,N_6199);
nand U7204 (N_7204,N_5827,N_5088);
nand U7205 (N_7205,N_5194,N_5594);
nand U7206 (N_7206,N_6144,N_5993);
xor U7207 (N_7207,N_5414,N_5614);
nor U7208 (N_7208,N_6084,N_5655);
xor U7209 (N_7209,N_5300,N_5998);
and U7210 (N_7210,N_5254,N_5622);
nor U7211 (N_7211,N_5171,N_5927);
or U7212 (N_7212,N_5569,N_5091);
or U7213 (N_7213,N_5652,N_5680);
nand U7214 (N_7214,N_6101,N_5732);
or U7215 (N_7215,N_6070,N_5569);
and U7216 (N_7216,N_5666,N_5556);
xor U7217 (N_7217,N_5107,N_5093);
xor U7218 (N_7218,N_6137,N_6231);
nand U7219 (N_7219,N_5880,N_5670);
or U7220 (N_7220,N_5656,N_5720);
and U7221 (N_7221,N_5973,N_5809);
or U7222 (N_7222,N_5902,N_6156);
and U7223 (N_7223,N_5744,N_5704);
and U7224 (N_7224,N_5112,N_5713);
nand U7225 (N_7225,N_5678,N_6032);
or U7226 (N_7226,N_5270,N_6110);
xor U7227 (N_7227,N_5291,N_5930);
xnor U7228 (N_7228,N_5184,N_6026);
nor U7229 (N_7229,N_5391,N_5899);
nor U7230 (N_7230,N_5312,N_5911);
nor U7231 (N_7231,N_6013,N_5714);
or U7232 (N_7232,N_5617,N_6102);
xor U7233 (N_7233,N_5646,N_5938);
nand U7234 (N_7234,N_5586,N_5200);
or U7235 (N_7235,N_5142,N_5008);
nor U7236 (N_7236,N_5793,N_5600);
nand U7237 (N_7237,N_5504,N_5712);
and U7238 (N_7238,N_5690,N_5438);
and U7239 (N_7239,N_5301,N_5182);
xnor U7240 (N_7240,N_6221,N_5439);
nor U7241 (N_7241,N_5312,N_6101);
or U7242 (N_7242,N_6052,N_6096);
or U7243 (N_7243,N_5627,N_5445);
nor U7244 (N_7244,N_5619,N_5818);
nand U7245 (N_7245,N_5182,N_5771);
and U7246 (N_7246,N_5462,N_5993);
nand U7247 (N_7247,N_5851,N_5126);
or U7248 (N_7248,N_5540,N_6105);
nand U7249 (N_7249,N_5211,N_5424);
nand U7250 (N_7250,N_5915,N_5823);
xor U7251 (N_7251,N_6165,N_6024);
and U7252 (N_7252,N_5454,N_6167);
and U7253 (N_7253,N_5701,N_5645);
and U7254 (N_7254,N_5762,N_5289);
or U7255 (N_7255,N_5597,N_5178);
and U7256 (N_7256,N_6192,N_6210);
xnor U7257 (N_7257,N_5532,N_5897);
nor U7258 (N_7258,N_5968,N_6050);
nor U7259 (N_7259,N_5610,N_5056);
nor U7260 (N_7260,N_5831,N_5607);
and U7261 (N_7261,N_5544,N_5672);
and U7262 (N_7262,N_5989,N_5781);
or U7263 (N_7263,N_5081,N_5390);
nor U7264 (N_7264,N_5868,N_6236);
and U7265 (N_7265,N_5468,N_5813);
nor U7266 (N_7266,N_6180,N_6015);
xnor U7267 (N_7267,N_6153,N_5284);
nand U7268 (N_7268,N_6188,N_6215);
and U7269 (N_7269,N_5061,N_5204);
nor U7270 (N_7270,N_5983,N_6230);
and U7271 (N_7271,N_6225,N_6155);
xnor U7272 (N_7272,N_5485,N_5973);
nor U7273 (N_7273,N_5809,N_5910);
nand U7274 (N_7274,N_5275,N_5881);
and U7275 (N_7275,N_5911,N_5229);
nand U7276 (N_7276,N_5801,N_5624);
xnor U7277 (N_7277,N_5980,N_5604);
nand U7278 (N_7278,N_6090,N_6215);
xor U7279 (N_7279,N_6081,N_6187);
nand U7280 (N_7280,N_5838,N_5590);
nand U7281 (N_7281,N_6071,N_5496);
or U7282 (N_7282,N_5251,N_5724);
or U7283 (N_7283,N_5889,N_5017);
and U7284 (N_7284,N_5987,N_6171);
and U7285 (N_7285,N_5956,N_6215);
nor U7286 (N_7286,N_5898,N_5900);
nor U7287 (N_7287,N_5163,N_5862);
and U7288 (N_7288,N_5679,N_5469);
nand U7289 (N_7289,N_5809,N_5025);
xnor U7290 (N_7290,N_5973,N_5390);
nand U7291 (N_7291,N_5689,N_5009);
or U7292 (N_7292,N_5408,N_5469);
and U7293 (N_7293,N_6192,N_6044);
or U7294 (N_7294,N_5590,N_6225);
nand U7295 (N_7295,N_5792,N_5857);
nand U7296 (N_7296,N_5860,N_6193);
nor U7297 (N_7297,N_6043,N_5426);
and U7298 (N_7298,N_5924,N_5307);
and U7299 (N_7299,N_5298,N_5418);
and U7300 (N_7300,N_5349,N_5816);
and U7301 (N_7301,N_5680,N_6122);
nand U7302 (N_7302,N_5544,N_5771);
nor U7303 (N_7303,N_5989,N_5212);
nor U7304 (N_7304,N_5738,N_6198);
xor U7305 (N_7305,N_5931,N_6125);
and U7306 (N_7306,N_5764,N_6093);
nand U7307 (N_7307,N_5551,N_5496);
nor U7308 (N_7308,N_5609,N_6030);
and U7309 (N_7309,N_5342,N_5351);
nor U7310 (N_7310,N_5497,N_6140);
nor U7311 (N_7311,N_5804,N_6162);
and U7312 (N_7312,N_5347,N_5918);
xor U7313 (N_7313,N_5037,N_5624);
and U7314 (N_7314,N_5018,N_6090);
nand U7315 (N_7315,N_6073,N_5250);
and U7316 (N_7316,N_6200,N_5346);
nor U7317 (N_7317,N_5468,N_5833);
and U7318 (N_7318,N_5489,N_5907);
nand U7319 (N_7319,N_5979,N_5968);
nor U7320 (N_7320,N_5198,N_5785);
nor U7321 (N_7321,N_5824,N_5828);
xor U7322 (N_7322,N_6098,N_6000);
nor U7323 (N_7323,N_6064,N_5154);
nor U7324 (N_7324,N_6074,N_5541);
nand U7325 (N_7325,N_5409,N_5837);
xor U7326 (N_7326,N_5895,N_5062);
nor U7327 (N_7327,N_5236,N_6148);
and U7328 (N_7328,N_5733,N_5235);
nand U7329 (N_7329,N_6026,N_6076);
xnor U7330 (N_7330,N_5818,N_6021);
and U7331 (N_7331,N_6048,N_5899);
xnor U7332 (N_7332,N_6124,N_5981);
or U7333 (N_7333,N_5482,N_6050);
or U7334 (N_7334,N_5639,N_5204);
nand U7335 (N_7335,N_5621,N_5526);
or U7336 (N_7336,N_5104,N_5449);
or U7337 (N_7337,N_5035,N_5357);
and U7338 (N_7338,N_5927,N_5912);
nor U7339 (N_7339,N_5556,N_5107);
and U7340 (N_7340,N_5853,N_5862);
or U7341 (N_7341,N_5116,N_5042);
nor U7342 (N_7342,N_5067,N_6219);
and U7343 (N_7343,N_5039,N_6234);
or U7344 (N_7344,N_5742,N_5358);
xnor U7345 (N_7345,N_5724,N_5854);
xnor U7346 (N_7346,N_5197,N_5852);
xnor U7347 (N_7347,N_5451,N_5535);
and U7348 (N_7348,N_5943,N_5809);
and U7349 (N_7349,N_5055,N_5987);
and U7350 (N_7350,N_5132,N_5588);
xnor U7351 (N_7351,N_5846,N_5816);
or U7352 (N_7352,N_5202,N_5730);
nand U7353 (N_7353,N_5491,N_5504);
or U7354 (N_7354,N_5350,N_5436);
and U7355 (N_7355,N_5306,N_5800);
and U7356 (N_7356,N_5427,N_5283);
nor U7357 (N_7357,N_5635,N_6082);
nand U7358 (N_7358,N_5147,N_5744);
xor U7359 (N_7359,N_5592,N_5227);
or U7360 (N_7360,N_5392,N_5694);
or U7361 (N_7361,N_6124,N_5745);
or U7362 (N_7362,N_5460,N_6036);
or U7363 (N_7363,N_5541,N_5312);
nand U7364 (N_7364,N_5179,N_5467);
or U7365 (N_7365,N_5752,N_5868);
nand U7366 (N_7366,N_5561,N_5470);
or U7367 (N_7367,N_5078,N_5834);
or U7368 (N_7368,N_5570,N_5627);
nand U7369 (N_7369,N_5454,N_5479);
nand U7370 (N_7370,N_5984,N_5456);
or U7371 (N_7371,N_5559,N_5564);
nand U7372 (N_7372,N_5115,N_5366);
and U7373 (N_7373,N_5297,N_5963);
or U7374 (N_7374,N_6210,N_5172);
nand U7375 (N_7375,N_5323,N_6145);
nor U7376 (N_7376,N_5621,N_5590);
or U7377 (N_7377,N_5906,N_5136);
nand U7378 (N_7378,N_5021,N_5848);
nand U7379 (N_7379,N_6221,N_5105);
xor U7380 (N_7380,N_5581,N_6143);
or U7381 (N_7381,N_5656,N_5810);
nor U7382 (N_7382,N_5731,N_6039);
and U7383 (N_7383,N_5653,N_6022);
and U7384 (N_7384,N_5336,N_6052);
nor U7385 (N_7385,N_5613,N_6245);
or U7386 (N_7386,N_5021,N_5139);
xnor U7387 (N_7387,N_6131,N_5816);
nor U7388 (N_7388,N_5838,N_5435);
or U7389 (N_7389,N_6214,N_5775);
and U7390 (N_7390,N_5410,N_5707);
nor U7391 (N_7391,N_5121,N_5176);
nor U7392 (N_7392,N_5535,N_5358);
xnor U7393 (N_7393,N_5668,N_5377);
nor U7394 (N_7394,N_5286,N_5498);
and U7395 (N_7395,N_5221,N_5519);
or U7396 (N_7396,N_5693,N_5135);
or U7397 (N_7397,N_6053,N_5933);
and U7398 (N_7398,N_5522,N_5597);
nand U7399 (N_7399,N_5010,N_5828);
nand U7400 (N_7400,N_5407,N_6087);
xor U7401 (N_7401,N_5657,N_5561);
or U7402 (N_7402,N_5845,N_5107);
or U7403 (N_7403,N_6129,N_6152);
xnor U7404 (N_7404,N_5240,N_5520);
xnor U7405 (N_7405,N_5933,N_5989);
and U7406 (N_7406,N_5662,N_5293);
nand U7407 (N_7407,N_5806,N_5053);
nor U7408 (N_7408,N_5923,N_6203);
nand U7409 (N_7409,N_6145,N_5856);
nand U7410 (N_7410,N_5997,N_5730);
and U7411 (N_7411,N_5373,N_6107);
and U7412 (N_7412,N_5164,N_5055);
nor U7413 (N_7413,N_5195,N_5755);
xnor U7414 (N_7414,N_6221,N_5288);
and U7415 (N_7415,N_5387,N_5990);
nand U7416 (N_7416,N_5777,N_6093);
nor U7417 (N_7417,N_6030,N_5846);
nor U7418 (N_7418,N_5200,N_5138);
nand U7419 (N_7419,N_6093,N_5952);
or U7420 (N_7420,N_5689,N_5589);
or U7421 (N_7421,N_5729,N_5773);
nor U7422 (N_7422,N_6247,N_6073);
nand U7423 (N_7423,N_5072,N_5056);
and U7424 (N_7424,N_6082,N_5114);
or U7425 (N_7425,N_5272,N_5574);
nand U7426 (N_7426,N_5447,N_5333);
or U7427 (N_7427,N_5942,N_6177);
and U7428 (N_7428,N_6067,N_5083);
and U7429 (N_7429,N_5068,N_5780);
nand U7430 (N_7430,N_5109,N_5907);
and U7431 (N_7431,N_5870,N_5719);
xor U7432 (N_7432,N_5956,N_5895);
and U7433 (N_7433,N_5927,N_5802);
xnor U7434 (N_7434,N_5897,N_5376);
or U7435 (N_7435,N_5466,N_5032);
nand U7436 (N_7436,N_5678,N_5073);
or U7437 (N_7437,N_5946,N_6076);
nand U7438 (N_7438,N_5393,N_5765);
and U7439 (N_7439,N_5670,N_5190);
nor U7440 (N_7440,N_5495,N_5053);
nand U7441 (N_7441,N_6140,N_5832);
nand U7442 (N_7442,N_6219,N_5890);
and U7443 (N_7443,N_5919,N_5429);
nand U7444 (N_7444,N_5033,N_5994);
or U7445 (N_7445,N_6200,N_5972);
and U7446 (N_7446,N_6019,N_5046);
nand U7447 (N_7447,N_5839,N_5807);
nand U7448 (N_7448,N_5103,N_6235);
and U7449 (N_7449,N_5971,N_5454);
nand U7450 (N_7450,N_5619,N_6051);
nand U7451 (N_7451,N_5126,N_6154);
nor U7452 (N_7452,N_5087,N_5933);
or U7453 (N_7453,N_5669,N_5020);
and U7454 (N_7454,N_5799,N_6082);
nor U7455 (N_7455,N_6004,N_5422);
and U7456 (N_7456,N_5017,N_5660);
nand U7457 (N_7457,N_5604,N_5581);
and U7458 (N_7458,N_5615,N_5466);
and U7459 (N_7459,N_5064,N_5212);
and U7460 (N_7460,N_5565,N_5304);
nor U7461 (N_7461,N_5904,N_5377);
and U7462 (N_7462,N_5312,N_5031);
and U7463 (N_7463,N_5834,N_6192);
or U7464 (N_7464,N_5168,N_5605);
xnor U7465 (N_7465,N_5837,N_6119);
nor U7466 (N_7466,N_5148,N_6083);
nor U7467 (N_7467,N_6060,N_5771);
and U7468 (N_7468,N_5003,N_5919);
nand U7469 (N_7469,N_5083,N_5180);
nand U7470 (N_7470,N_6176,N_5936);
nor U7471 (N_7471,N_5909,N_5967);
and U7472 (N_7472,N_6137,N_6062);
nor U7473 (N_7473,N_5370,N_5479);
and U7474 (N_7474,N_5204,N_5427);
xnor U7475 (N_7475,N_5309,N_5897);
xnor U7476 (N_7476,N_5045,N_5896);
or U7477 (N_7477,N_5741,N_5603);
nor U7478 (N_7478,N_5965,N_5092);
nand U7479 (N_7479,N_5722,N_5664);
or U7480 (N_7480,N_6197,N_5785);
nor U7481 (N_7481,N_5934,N_5180);
and U7482 (N_7482,N_5585,N_6227);
nand U7483 (N_7483,N_5854,N_5591);
xnor U7484 (N_7484,N_5618,N_5691);
and U7485 (N_7485,N_5286,N_6085);
or U7486 (N_7486,N_5935,N_6112);
or U7487 (N_7487,N_5818,N_5568);
and U7488 (N_7488,N_5413,N_5754);
xnor U7489 (N_7489,N_5317,N_5367);
or U7490 (N_7490,N_5102,N_6042);
nand U7491 (N_7491,N_5427,N_6114);
and U7492 (N_7492,N_5590,N_5924);
nor U7493 (N_7493,N_5412,N_6007);
nand U7494 (N_7494,N_5385,N_5191);
and U7495 (N_7495,N_5381,N_6078);
nand U7496 (N_7496,N_5651,N_5449);
xor U7497 (N_7497,N_5862,N_6127);
and U7498 (N_7498,N_6083,N_5164);
xor U7499 (N_7499,N_5090,N_6071);
xor U7500 (N_7500,N_7241,N_6688);
or U7501 (N_7501,N_7192,N_7492);
nand U7502 (N_7502,N_7057,N_7391);
nand U7503 (N_7503,N_6697,N_6947);
nor U7504 (N_7504,N_7307,N_7035);
or U7505 (N_7505,N_6499,N_6591);
xor U7506 (N_7506,N_7411,N_6577);
and U7507 (N_7507,N_6358,N_6425);
xnor U7508 (N_7508,N_6286,N_7060);
nor U7509 (N_7509,N_7022,N_6494);
nand U7510 (N_7510,N_6567,N_7319);
and U7511 (N_7511,N_6768,N_6620);
nand U7512 (N_7512,N_7385,N_7376);
nand U7513 (N_7513,N_7250,N_7470);
xnor U7514 (N_7514,N_6710,N_7291);
and U7515 (N_7515,N_6434,N_7464);
xor U7516 (N_7516,N_6338,N_6738);
nand U7517 (N_7517,N_7432,N_6865);
and U7518 (N_7518,N_6760,N_7354);
xor U7519 (N_7519,N_7176,N_7325);
xnor U7520 (N_7520,N_6344,N_6551);
nand U7521 (N_7521,N_6655,N_6307);
and U7522 (N_7522,N_7439,N_7284);
xnor U7523 (N_7523,N_7412,N_6519);
nor U7524 (N_7524,N_6582,N_7332);
nand U7525 (N_7525,N_7251,N_6848);
nand U7526 (N_7526,N_7457,N_7487);
nor U7527 (N_7527,N_7100,N_7488);
and U7528 (N_7528,N_6896,N_6803);
nand U7529 (N_7529,N_7358,N_7016);
nor U7530 (N_7530,N_6790,N_7047);
and U7531 (N_7531,N_6492,N_6424);
nand U7532 (N_7532,N_6703,N_6621);
nor U7533 (N_7533,N_6256,N_6983);
and U7534 (N_7534,N_6742,N_6676);
nand U7535 (N_7535,N_6780,N_7223);
or U7536 (N_7536,N_7407,N_7215);
and U7537 (N_7537,N_6337,N_7165);
nand U7538 (N_7538,N_7114,N_7294);
xor U7539 (N_7539,N_6754,N_7170);
xnor U7540 (N_7540,N_6900,N_6430);
and U7541 (N_7541,N_6648,N_6733);
nand U7542 (N_7542,N_6299,N_6277);
or U7543 (N_7543,N_7304,N_7327);
and U7544 (N_7544,N_7097,N_6287);
nand U7545 (N_7545,N_6909,N_6642);
nand U7546 (N_7546,N_6258,N_6651);
or U7547 (N_7547,N_6535,N_6480);
and U7548 (N_7548,N_6934,N_6352);
xor U7549 (N_7549,N_6894,N_6407);
nor U7550 (N_7550,N_7220,N_6594);
or U7551 (N_7551,N_6883,N_6601);
and U7552 (N_7552,N_6390,N_7103);
nand U7553 (N_7553,N_7036,N_7217);
nor U7554 (N_7554,N_6922,N_6412);
xnor U7555 (N_7555,N_6952,N_6614);
xnor U7556 (N_7556,N_6626,N_7414);
xnor U7557 (N_7557,N_7127,N_6787);
and U7558 (N_7558,N_6300,N_7038);
nor U7559 (N_7559,N_6808,N_6441);
nor U7560 (N_7560,N_6255,N_7473);
or U7561 (N_7561,N_7151,N_6931);
or U7562 (N_7562,N_6397,N_6961);
and U7563 (N_7563,N_7401,N_7474);
and U7564 (N_7564,N_6758,N_7078);
nor U7565 (N_7565,N_7377,N_6455);
nand U7566 (N_7566,N_6964,N_6264);
or U7567 (N_7567,N_7044,N_7096);
nor U7568 (N_7568,N_7454,N_6654);
and U7569 (N_7569,N_6868,N_7183);
and U7570 (N_7570,N_7074,N_7123);
and U7571 (N_7571,N_7013,N_6580);
and U7572 (N_7572,N_7417,N_6978);
nand U7573 (N_7573,N_7026,N_6731);
and U7574 (N_7574,N_6290,N_6971);
nand U7575 (N_7575,N_6788,N_7300);
and U7576 (N_7576,N_7196,N_6418);
and U7577 (N_7577,N_7471,N_6717);
nand U7578 (N_7578,N_6857,N_6377);
or U7579 (N_7579,N_7384,N_6454);
and U7580 (N_7580,N_6420,N_6432);
and U7581 (N_7581,N_6289,N_6734);
nor U7582 (N_7582,N_6773,N_6263);
or U7583 (N_7583,N_6340,N_6834);
nand U7584 (N_7584,N_6638,N_7476);
nor U7585 (N_7585,N_7469,N_7484);
or U7586 (N_7586,N_6807,N_6702);
or U7587 (N_7587,N_6810,N_6438);
and U7588 (N_7588,N_6360,N_6715);
xnor U7589 (N_7589,N_7226,N_6720);
xor U7590 (N_7590,N_6907,N_6914);
nor U7591 (N_7591,N_6942,N_7191);
nor U7592 (N_7592,N_6837,N_7399);
or U7593 (N_7593,N_6872,N_7054);
and U7594 (N_7594,N_6449,N_7477);
or U7595 (N_7595,N_6730,N_6437);
nand U7596 (N_7596,N_7310,N_7283);
nand U7597 (N_7597,N_6483,N_7208);
or U7598 (N_7598,N_6252,N_7059);
and U7599 (N_7599,N_6926,N_6280);
nand U7600 (N_7600,N_7328,N_6747);
xor U7601 (N_7601,N_6472,N_6291);
nor U7602 (N_7602,N_7426,N_6635);
xnor U7603 (N_7603,N_7298,N_7353);
xor U7604 (N_7604,N_6431,N_7169);
nand U7605 (N_7605,N_6276,N_7380);
and U7606 (N_7606,N_7105,N_7340);
nor U7607 (N_7607,N_6955,N_7289);
xnor U7608 (N_7608,N_7039,N_6871);
and U7609 (N_7609,N_6728,N_7005);
nor U7610 (N_7610,N_6849,N_6295);
xor U7611 (N_7611,N_6321,N_6714);
nand U7612 (N_7612,N_6481,N_6991);
xnor U7613 (N_7613,N_7404,N_6799);
xnor U7614 (N_7614,N_7315,N_6313);
nor U7615 (N_7615,N_7428,N_6466);
nand U7616 (N_7616,N_6963,N_7436);
xor U7617 (N_7617,N_7356,N_6504);
or U7618 (N_7618,N_6285,N_7027);
and U7619 (N_7619,N_6716,N_6643);
xnor U7620 (N_7620,N_6552,N_6405);
nand U7621 (N_7621,N_6759,N_7425);
xnor U7622 (N_7622,N_6673,N_7366);
nor U7623 (N_7623,N_6801,N_6330);
and U7624 (N_7624,N_6969,N_6452);
or U7625 (N_7625,N_6569,N_7440);
and U7626 (N_7626,N_7434,N_7453);
nor U7627 (N_7627,N_6895,N_6615);
nand U7628 (N_7628,N_6924,N_7085);
xnor U7629 (N_7629,N_6393,N_7086);
xor U7630 (N_7630,N_7032,N_6435);
and U7631 (N_7631,N_7478,N_7280);
and U7632 (N_7632,N_7331,N_7224);
nand U7633 (N_7633,N_7371,N_7024);
xnor U7634 (N_7634,N_6553,N_6928);
and U7635 (N_7635,N_7347,N_6973);
and U7636 (N_7636,N_6279,N_6404);
and U7637 (N_7637,N_6274,N_7333);
nand U7638 (N_7638,N_7359,N_7372);
nand U7639 (N_7639,N_7137,N_6361);
nor U7640 (N_7640,N_6858,N_6736);
or U7641 (N_7641,N_6305,N_6386);
nand U7642 (N_7642,N_6378,N_6260);
nor U7643 (N_7643,N_6881,N_7465);
nor U7644 (N_7644,N_7066,N_7423);
nand U7645 (N_7645,N_6892,N_7240);
xor U7646 (N_7646,N_7007,N_7205);
or U7647 (N_7647,N_6254,N_7337);
nor U7648 (N_7648,N_7209,N_6828);
nand U7649 (N_7649,N_6270,N_7132);
or U7650 (N_7650,N_6605,N_6656);
xnor U7651 (N_7651,N_6689,N_7180);
and U7652 (N_7652,N_7216,N_7444);
or U7653 (N_7653,N_6525,N_6941);
nand U7654 (N_7654,N_6319,N_6613);
xnor U7655 (N_7655,N_6867,N_6541);
nand U7656 (N_7656,N_7301,N_6379);
xor U7657 (N_7657,N_7125,N_6984);
and U7658 (N_7658,N_6999,N_6584);
xor U7659 (N_7659,N_7142,N_6815);
or U7660 (N_7660,N_6581,N_6311);
nor U7661 (N_7661,N_6681,N_6987);
nor U7662 (N_7662,N_7480,N_7239);
xor U7663 (N_7663,N_7313,N_6953);
nor U7664 (N_7664,N_6817,N_6485);
xor U7665 (N_7665,N_6832,N_6554);
and U7666 (N_7666,N_6528,N_6746);
or U7667 (N_7667,N_7056,N_6958);
xnor U7668 (N_7668,N_7058,N_6380);
nand U7669 (N_7669,N_7257,N_6735);
nor U7670 (N_7670,N_6427,N_6726);
nand U7671 (N_7671,N_6335,N_6923);
xor U7672 (N_7672,N_6444,N_7211);
or U7673 (N_7673,N_7475,N_6328);
or U7674 (N_7674,N_6901,N_6644);
nor U7675 (N_7675,N_7387,N_6312);
nand U7676 (N_7676,N_6765,N_7050);
nor U7677 (N_7677,N_7030,N_7431);
nand U7678 (N_7678,N_6536,N_7258);
and U7679 (N_7679,N_6318,N_6320);
or U7680 (N_7680,N_6273,N_7194);
xor U7681 (N_7681,N_7247,N_6473);
nor U7682 (N_7682,N_7441,N_6779);
and U7683 (N_7683,N_6331,N_7330);
nor U7684 (N_7684,N_6829,N_6253);
nor U7685 (N_7685,N_6529,N_6575);
xor U7686 (N_7686,N_6645,N_7438);
and U7687 (N_7687,N_7177,N_6686);
and U7688 (N_7688,N_6721,N_6636);
xor U7689 (N_7689,N_7343,N_7246);
nor U7690 (N_7690,N_6699,N_7134);
nor U7691 (N_7691,N_6884,N_6446);
or U7692 (N_7692,N_7034,N_6532);
and U7693 (N_7693,N_7272,N_6513);
and U7694 (N_7694,N_7167,N_7214);
nand U7695 (N_7695,N_6346,N_7419);
nor U7696 (N_7696,N_6469,N_7120);
nand U7697 (N_7697,N_7263,N_7067);
xnor U7698 (N_7698,N_6394,N_6869);
or U7699 (N_7699,N_7275,N_6985);
or U7700 (N_7700,N_7421,N_7140);
or U7701 (N_7701,N_6911,N_6744);
nor U7702 (N_7702,N_6443,N_7261);
and U7703 (N_7703,N_7163,N_6861);
or U7704 (N_7704,N_6606,N_6351);
nor U7705 (N_7705,N_7029,N_7264);
and U7706 (N_7706,N_6675,N_6692);
nand U7707 (N_7707,N_6448,N_6946);
or U7708 (N_7708,N_7020,N_6793);
nand U7709 (N_7709,N_6570,N_7302);
nand U7710 (N_7710,N_6453,N_7292);
nor U7711 (N_7711,N_7023,N_6853);
nand U7712 (N_7712,N_7445,N_6559);
nand U7713 (N_7713,N_6657,N_6595);
nor U7714 (N_7714,N_7461,N_7447);
nand U7715 (N_7715,N_6622,N_7221);
xor U7716 (N_7716,N_6557,N_6830);
nor U7717 (N_7717,N_6477,N_7113);
nor U7718 (N_7718,N_6538,N_6677);
nor U7719 (N_7719,N_6791,N_7061);
xor U7720 (N_7720,N_6356,N_6745);
nand U7721 (N_7721,N_6265,N_6332);
nand U7722 (N_7722,N_6683,N_6893);
and U7723 (N_7723,N_6457,N_6399);
xnor U7724 (N_7724,N_7168,N_6566);
nor U7725 (N_7725,N_7228,N_6724);
xor U7726 (N_7726,N_6609,N_6740);
nor U7727 (N_7727,N_6695,N_6863);
nor U7728 (N_7728,N_7346,N_7269);
nor U7729 (N_7729,N_7468,N_7348);
nand U7730 (N_7730,N_6732,N_7293);
nand U7731 (N_7731,N_7197,N_7006);
nor U7732 (N_7732,N_6616,N_6889);
xor U7733 (N_7733,N_6451,N_6339);
nand U7734 (N_7734,N_6384,N_6269);
nand U7735 (N_7735,N_7463,N_6669);
and U7736 (N_7736,N_6981,N_7479);
or U7737 (N_7737,N_7102,N_6467);
nor U7738 (N_7738,N_6599,N_7104);
nor U7739 (N_7739,N_7010,N_7203);
nand U7740 (N_7740,N_6365,N_6992);
or U7741 (N_7741,N_6891,N_6366);
and U7742 (N_7742,N_6854,N_6342);
nand U7743 (N_7743,N_7200,N_7312);
xnor U7744 (N_7744,N_6661,N_6476);
xor U7745 (N_7745,N_7450,N_6388);
nor U7746 (N_7746,N_6370,N_6488);
or U7747 (N_7747,N_6461,N_7236);
nor U7748 (N_7748,N_6664,N_7396);
and U7749 (N_7749,N_6850,N_7318);
nor U7750 (N_7750,N_7198,N_6727);
xnor U7751 (N_7751,N_6995,N_6348);
xor U7752 (N_7752,N_6826,N_6521);
or U7753 (N_7753,N_6560,N_6387);
nand U7754 (N_7754,N_6296,N_7344);
nor U7755 (N_7755,N_6628,N_6633);
xor U7756 (N_7756,N_6306,N_6442);
and U7757 (N_7757,N_6814,N_6842);
xnor U7758 (N_7758,N_7147,N_6267);
nor U7759 (N_7759,N_6956,N_7055);
and U7760 (N_7760,N_6761,N_7083);
and U7761 (N_7761,N_6988,N_6663);
nand U7762 (N_7762,N_6887,N_6957);
nor U7763 (N_7763,N_7043,N_7281);
xnor U7764 (N_7764,N_6960,N_6281);
nor U7765 (N_7765,N_7213,N_7124);
xnor U7766 (N_7766,N_6766,N_6250);
nor U7767 (N_7767,N_7162,N_6840);
xnor U7768 (N_7768,N_6283,N_6798);
xnor U7769 (N_7769,N_7430,N_7388);
nand U7770 (N_7770,N_7279,N_7107);
and U7771 (N_7771,N_6414,N_7004);
nor U7772 (N_7772,N_7225,N_7278);
nand U7773 (N_7773,N_6403,N_7070);
or U7774 (N_7774,N_6796,N_6308);
nand U7775 (N_7775,N_7449,N_7111);
nand U7776 (N_7776,N_6870,N_7028);
nand U7777 (N_7777,N_7156,N_7260);
nor U7778 (N_7778,N_7497,N_6514);
xnor U7779 (N_7779,N_6395,N_7459);
or U7780 (N_7780,N_6345,N_7413);
and U7781 (N_7781,N_6336,N_7185);
or U7782 (N_7782,N_6972,N_7046);
or U7783 (N_7783,N_6847,N_6712);
nor U7784 (N_7784,N_6563,N_6813);
or U7785 (N_7785,N_7173,N_6792);
nor U7786 (N_7786,N_7234,N_6709);
nor U7787 (N_7787,N_6593,N_6753);
or U7788 (N_7788,N_6932,N_7429);
or U7789 (N_7789,N_6687,N_6827);
and U7790 (N_7790,N_7122,N_6315);
xnor U7791 (N_7791,N_7481,N_6350);
nor U7792 (N_7792,N_6925,N_6439);
and U7793 (N_7793,N_6498,N_7498);
xnor U7794 (N_7794,N_6693,N_6800);
or U7795 (N_7795,N_6505,N_6284);
nand U7796 (N_7796,N_7222,N_6371);
nand U7797 (N_7797,N_7121,N_6588);
nand U7798 (N_7798,N_7448,N_6920);
or U7799 (N_7799,N_6516,N_6561);
or U7800 (N_7800,N_6764,N_6293);
xnor U7801 (N_7801,N_7187,N_6470);
and U7802 (N_7802,N_6706,N_6515);
nor U7803 (N_7803,N_6708,N_7141);
and U7804 (N_7804,N_6372,N_7095);
xnor U7805 (N_7805,N_7231,N_7323);
xnor U7806 (N_7806,N_7357,N_6718);
or U7807 (N_7807,N_6422,N_7424);
xor U7808 (N_7808,N_6450,N_6625);
or U7809 (N_7809,N_7071,N_7227);
or U7810 (N_7810,N_6824,N_7415);
and U7811 (N_7811,N_6292,N_6927);
nand U7812 (N_7812,N_6782,N_6259);
or U7813 (N_7813,N_6748,N_7073);
nor U7814 (N_7814,N_7229,N_6326);
xor U7815 (N_7815,N_7131,N_6685);
nand U7816 (N_7816,N_7206,N_7255);
xor U7817 (N_7817,N_7063,N_6413);
and U7818 (N_7818,N_6885,N_6755);
and U7819 (N_7819,N_6771,N_7322);
nor U7820 (N_7820,N_7375,N_7287);
nand U7821 (N_7821,N_6409,N_7108);
nor U7822 (N_7822,N_6478,N_6507);
nand U7823 (N_7823,N_7379,N_6659);
and U7824 (N_7824,N_6596,N_6542);
or U7825 (N_7825,N_6583,N_6977);
or U7826 (N_7826,N_7150,N_7017);
nor U7827 (N_7827,N_7299,N_6534);
nand U7828 (N_7828,N_6862,N_6989);
nor U7829 (N_7829,N_6266,N_6341);
and U7830 (N_7830,N_7045,N_6767);
or U7831 (N_7831,N_6608,N_7277);
and U7832 (N_7832,N_6607,N_6866);
or U7833 (N_7833,N_7119,N_7079);
xnor U7834 (N_7834,N_7297,N_7362);
nand U7835 (N_7835,N_6524,N_7336);
xnor U7836 (N_7836,N_6354,N_7199);
and U7837 (N_7837,N_6774,N_6310);
nor U7838 (N_7838,N_6951,N_6831);
nor U7839 (N_7839,N_6789,N_6667);
or U7840 (N_7840,N_6489,N_6839);
or U7841 (N_7841,N_6589,N_6324);
nand U7842 (N_7842,N_6979,N_7406);
nand U7843 (N_7843,N_6304,N_7329);
nand U7844 (N_7844,N_7311,N_7326);
or U7845 (N_7845,N_6410,N_7068);
or U7846 (N_7846,N_6484,N_7166);
and U7847 (N_7847,N_7159,N_7296);
xor U7848 (N_7848,N_6913,N_6502);
xnor U7849 (N_7849,N_6713,N_6509);
nand U7850 (N_7850,N_6739,N_6882);
and U7851 (N_7851,N_6333,N_7365);
xor U7852 (N_7852,N_6316,N_7018);
nand U7853 (N_7853,N_7395,N_6804);
nand U7854 (N_7854,N_7427,N_6428);
xnor U7855 (N_7855,N_7352,N_6805);
xor U7856 (N_7856,N_6411,N_6684);
or U7857 (N_7857,N_7037,N_6943);
xor U7858 (N_7858,N_6844,N_7249);
nor U7859 (N_7859,N_6347,N_7181);
and U7860 (N_7860,N_7065,N_7485);
or U7861 (N_7861,N_6875,N_7253);
xnor U7862 (N_7862,N_6612,N_6543);
nand U7863 (N_7863,N_6694,N_6497);
xnor U7864 (N_7864,N_6629,N_7295);
or U7865 (N_7865,N_6298,N_7233);
xor U7866 (N_7866,N_7069,N_7155);
nand U7867 (N_7867,N_6468,N_6729);
nand U7868 (N_7868,N_6864,N_7252);
nand U7869 (N_7869,N_7491,N_7410);
nor U7870 (N_7870,N_7174,N_6375);
nor U7871 (N_7871,N_7153,N_6835);
and U7872 (N_7872,N_6322,N_6303);
nor U7873 (N_7873,N_6619,N_6539);
nor U7874 (N_7874,N_6775,N_7386);
nand U7875 (N_7875,N_6772,N_6398);
nand U7876 (N_7876,N_6937,N_7072);
nor U7877 (N_7877,N_6627,N_6520);
nor U7878 (N_7878,N_7433,N_6314);
nor U7879 (N_7879,N_7402,N_7370);
nand U7880 (N_7880,N_6503,N_7256);
or U7881 (N_7881,N_7171,N_7207);
or U7882 (N_7882,N_7446,N_6373);
nand U7883 (N_7883,N_7400,N_7305);
or U7884 (N_7884,N_7160,N_6423);
and U7885 (N_7885,N_6776,N_6278);
nor U7886 (N_7886,N_7466,N_6898);
nor U7887 (N_7887,N_7052,N_7314);
xnor U7888 (N_7888,N_6757,N_7369);
nand U7889 (N_7889,N_6944,N_7266);
nor U7890 (N_7890,N_6940,N_6906);
xor U7891 (N_7891,N_7398,N_6672);
and U7892 (N_7892,N_6573,N_6666);
nand U7893 (N_7893,N_7143,N_7130);
or U7894 (N_7894,N_6751,N_7094);
nand U7895 (N_7895,N_7361,N_6391);
or U7896 (N_7896,N_6618,N_7349);
nor U7897 (N_7897,N_6549,N_6938);
and U7898 (N_7898,N_6576,N_7285);
or U7899 (N_7899,N_6701,N_7378);
nand U7900 (N_7900,N_6462,N_6678);
nor U7901 (N_7901,N_7040,N_6668);
or U7902 (N_7902,N_6841,N_7368);
and U7903 (N_7903,N_6610,N_6976);
and U7904 (N_7904,N_7238,N_7182);
and U7905 (N_7905,N_7483,N_6851);
nand U7906 (N_7906,N_7129,N_6919);
or U7907 (N_7907,N_6876,N_7077);
and U7908 (N_7908,N_6811,N_7242);
xor U7909 (N_7909,N_7091,N_6674);
and U7910 (N_7910,N_6617,N_7495);
and U7911 (N_7911,N_6374,N_6297);
and U7912 (N_7912,N_6750,N_7321);
or U7913 (N_7913,N_6406,N_7409);
and U7914 (N_7914,N_6743,N_7053);
xnor U7915 (N_7915,N_7075,N_6275);
and U7916 (N_7916,N_6860,N_6630);
or U7917 (N_7917,N_7193,N_6998);
xor U7918 (N_7918,N_7342,N_6624);
or U7919 (N_7919,N_7009,N_6517);
nor U7920 (N_7920,N_6475,N_7076);
xnor U7921 (N_7921,N_6641,N_7408);
xnor U7922 (N_7922,N_7355,N_7397);
nor U7923 (N_7923,N_6261,N_6385);
and U7924 (N_7924,N_6571,N_7099);
or U7925 (N_7925,N_7364,N_6527);
nand U7926 (N_7926,N_6741,N_7262);
and U7927 (N_7927,N_7276,N_6592);
nand U7928 (N_7928,N_6996,N_7462);
nand U7929 (N_7929,N_7403,N_6873);
and U7930 (N_7930,N_7317,N_6433);
or U7931 (N_7931,N_7031,N_7392);
and U7932 (N_7932,N_6474,N_6994);
nor U7933 (N_7933,N_6939,N_6878);
nor U7934 (N_7934,N_6819,N_6763);
and U7935 (N_7935,N_7288,N_6417);
nor U7936 (N_7936,N_6558,N_7308);
nor U7937 (N_7937,N_7303,N_6719);
nor U7938 (N_7938,N_6631,N_7338);
xnor U7939 (N_7939,N_6491,N_6334);
xnor U7940 (N_7940,N_7456,N_6353);
nor U7941 (N_7941,N_6646,N_6637);
nand U7942 (N_7942,N_6396,N_6945);
xnor U7943 (N_7943,N_7394,N_6846);
or U7944 (N_7944,N_6650,N_6822);
nor U7945 (N_7945,N_7270,N_7245);
nand U7946 (N_7946,N_6632,N_6647);
nand U7947 (N_7947,N_7145,N_6268);
or U7948 (N_7948,N_7081,N_6522);
nand U7949 (N_7949,N_7115,N_6935);
and U7950 (N_7950,N_6518,N_6806);
nand U7951 (N_7951,N_6970,N_7244);
nor U7952 (N_7952,N_7008,N_7273);
nor U7953 (N_7953,N_6288,N_7493);
or U7954 (N_7954,N_6680,N_6362);
nor U7955 (N_7955,N_6262,N_7443);
or U7956 (N_7956,N_6369,N_7161);
or U7957 (N_7957,N_7033,N_7092);
nand U7958 (N_7958,N_6662,N_6812);
xnor U7959 (N_7959,N_7286,N_6968);
nand U7960 (N_7960,N_7179,N_7467);
xnor U7961 (N_7961,N_7494,N_7000);
or U7962 (N_7962,N_6691,N_6954);
nand U7963 (N_7963,N_6343,N_7116);
nor U7964 (N_7964,N_6421,N_7204);
nand U7965 (N_7965,N_6856,N_6349);
xnor U7966 (N_7966,N_7267,N_7049);
and U7967 (N_7967,N_6905,N_7218);
and U7968 (N_7968,N_7080,N_6690);
nor U7969 (N_7969,N_7486,N_7499);
nand U7970 (N_7970,N_7232,N_6586);
xor U7971 (N_7971,N_6402,N_6456);
or U7972 (N_7972,N_7437,N_6783);
nor U7973 (N_7973,N_7363,N_7243);
or U7974 (N_7974,N_7381,N_6556);
or U7975 (N_7975,N_7345,N_6722);
xnor U7976 (N_7976,N_6910,N_6912);
nand U7977 (N_7977,N_6671,N_7389);
nand U7978 (N_7978,N_6816,N_6965);
and U7979 (N_7979,N_7133,N_6464);
nand U7980 (N_7980,N_7003,N_6917);
nor U7981 (N_7981,N_7309,N_6725);
or U7982 (N_7982,N_7335,N_7090);
nand U7983 (N_7983,N_6309,N_6392);
nor U7984 (N_7984,N_6833,N_6459);
or U7985 (N_7985,N_6465,N_6665);
or U7986 (N_7986,N_7316,N_6508);
and U7987 (N_7987,N_7442,N_7383);
nor U7988 (N_7988,N_7062,N_7148);
xnor U7989 (N_7989,N_7489,N_6975);
nor U7990 (N_7990,N_6482,N_7189);
or U7991 (N_7991,N_6426,N_7126);
or U7992 (N_7992,N_7164,N_6447);
or U7993 (N_7993,N_6936,N_6859);
or U7994 (N_7994,N_6962,N_6902);
xor U7995 (N_7995,N_6921,N_6933);
nand U7996 (N_7996,N_6251,N_6825);
nor U7997 (N_7997,N_6929,N_7118);
xor U7998 (N_7998,N_6982,N_6323);
or U7999 (N_7999,N_7341,N_7393);
or U8000 (N_8000,N_6325,N_6623);
nand U8001 (N_8001,N_6546,N_6572);
nor U8002 (N_8002,N_6704,N_7382);
nor U8003 (N_8003,N_7339,N_6317);
nor U8004 (N_8004,N_7184,N_6852);
nor U8005 (N_8005,N_6537,N_6698);
nor U8006 (N_8006,N_6530,N_6598);
and U8007 (N_8007,N_6752,N_6794);
and U8008 (N_8008,N_6652,N_6781);
or U8009 (N_8009,N_7458,N_6587);
or U8010 (N_8010,N_6400,N_7248);
nand U8011 (N_8011,N_6578,N_6544);
or U8012 (N_8012,N_6408,N_6821);
or U8013 (N_8013,N_7087,N_6548);
nand U8014 (N_8014,N_7268,N_6496);
nor U8015 (N_8015,N_6762,N_6918);
nor U8016 (N_8016,N_6795,N_6500);
nor U8017 (N_8017,N_6899,N_7139);
nor U8018 (N_8018,N_7089,N_6890);
nor U8019 (N_8019,N_7195,N_6877);
nor U8020 (N_8020,N_6679,N_7138);
nor U8021 (N_8021,N_7435,N_6980);
or U8022 (N_8022,N_7351,N_6574);
or U8023 (N_8023,N_6376,N_7350);
or U8024 (N_8024,N_7175,N_7452);
nor U8025 (N_8025,N_6471,N_6836);
xor U8026 (N_8026,N_7254,N_6990);
xor U8027 (N_8027,N_6600,N_7420);
nand U8028 (N_8028,N_7011,N_7451);
xnor U8029 (N_8029,N_6797,N_6974);
nor U8030 (N_8030,N_7405,N_6705);
or U8031 (N_8031,N_7290,N_6355);
or U8032 (N_8032,N_6639,N_6531);
or U8033 (N_8033,N_6784,N_6930);
nand U8034 (N_8034,N_7021,N_6383);
xor U8035 (N_8035,N_6329,N_7360);
xor U8036 (N_8036,N_7082,N_6429);
nand U8037 (N_8037,N_6823,N_6845);
and U8038 (N_8038,N_7093,N_7422);
and U8039 (N_8039,N_6967,N_6565);
nor U8040 (N_8040,N_6604,N_6523);
nand U8041 (N_8041,N_6257,N_6294);
nor U8042 (N_8042,N_7455,N_6707);
nand U8043 (N_8043,N_6440,N_6368);
and U8044 (N_8044,N_7178,N_7012);
nand U8045 (N_8045,N_7144,N_6653);
nand U8046 (N_8046,N_7042,N_7136);
or U8047 (N_8047,N_7186,N_7001);
or U8048 (N_8048,N_6416,N_7015);
nand U8049 (N_8049,N_6282,N_7064);
nand U8050 (N_8050,N_7282,N_6649);
nand U8051 (N_8051,N_6564,N_7048);
or U8052 (N_8052,N_6820,N_6562);
xor U8053 (N_8053,N_6436,N_6302);
nand U8054 (N_8054,N_6506,N_6585);
nand U8055 (N_8055,N_6658,N_6511);
or U8056 (N_8056,N_6389,N_6640);
or U8057 (N_8057,N_7416,N_6359);
xor U8058 (N_8058,N_7212,N_6915);
nand U8059 (N_8059,N_6579,N_6495);
or U8060 (N_8060,N_7106,N_7146);
xnor U8061 (N_8061,N_7101,N_6888);
and U8062 (N_8062,N_6737,N_7041);
or U8063 (N_8063,N_6555,N_6550);
nor U8064 (N_8064,N_6696,N_6904);
nor U8065 (N_8065,N_6880,N_7002);
and U8066 (N_8066,N_7306,N_6756);
nand U8067 (N_8067,N_6401,N_6897);
or U8068 (N_8068,N_7154,N_6723);
or U8069 (N_8069,N_7117,N_6843);
nand U8070 (N_8070,N_7025,N_7109);
or U8071 (N_8071,N_6959,N_7237);
xnor U8072 (N_8072,N_6993,N_6301);
and U8073 (N_8073,N_6770,N_6526);
nand U8074 (N_8074,N_7172,N_6363);
nand U8075 (N_8075,N_7230,N_6512);
and U8076 (N_8076,N_6948,N_6568);
nor U8077 (N_8077,N_6364,N_7098);
or U8078 (N_8078,N_6602,N_6749);
xor U8079 (N_8079,N_6445,N_7390);
and U8080 (N_8080,N_7235,N_7324);
and U8081 (N_8081,N_6682,N_6590);
nand U8082 (N_8082,N_6533,N_6777);
or U8083 (N_8083,N_7418,N_6986);
or U8084 (N_8084,N_6597,N_6886);
nand U8085 (N_8085,N_6660,N_6510);
and U8086 (N_8086,N_6700,N_6949);
and U8087 (N_8087,N_6785,N_6603);
and U8088 (N_8088,N_7112,N_7472);
and U8089 (N_8089,N_6357,N_6903);
or U8090 (N_8090,N_6838,N_6778);
nand U8091 (N_8091,N_6271,N_6711);
and U8092 (N_8092,N_6540,N_6818);
nand U8093 (N_8093,N_6786,N_6486);
nand U8094 (N_8094,N_6879,N_7158);
nand U8095 (N_8095,N_7157,N_6501);
or U8096 (N_8096,N_6916,N_7259);
xor U8097 (N_8097,N_6611,N_7460);
nand U8098 (N_8098,N_6419,N_7152);
or U8099 (N_8099,N_7320,N_7490);
or U8100 (N_8100,N_6966,N_6458);
nor U8101 (N_8101,N_6415,N_6908);
nor U8102 (N_8102,N_6272,N_7265);
or U8103 (N_8103,N_7019,N_7088);
nor U8104 (N_8104,N_6769,N_6545);
nand U8105 (N_8105,N_7496,N_7334);
and U8106 (N_8106,N_6634,N_6547);
or U8107 (N_8107,N_6479,N_7367);
xnor U8108 (N_8108,N_6493,N_6490);
xor U8109 (N_8109,N_6809,N_6874);
and U8110 (N_8110,N_7219,N_6463);
or U8111 (N_8111,N_6802,N_7271);
nand U8112 (N_8112,N_7190,N_7128);
nand U8113 (N_8113,N_7373,N_6367);
and U8114 (N_8114,N_7110,N_6670);
nor U8115 (N_8115,N_7374,N_7149);
and U8116 (N_8116,N_7084,N_6950);
or U8117 (N_8117,N_6997,N_7202);
or U8118 (N_8118,N_6460,N_6855);
or U8119 (N_8119,N_7188,N_6381);
and U8120 (N_8120,N_6487,N_7482);
nor U8121 (N_8121,N_7274,N_7135);
nor U8122 (N_8122,N_7014,N_7201);
or U8123 (N_8123,N_7210,N_7051);
or U8124 (N_8124,N_6327,N_6382);
xor U8125 (N_8125,N_7438,N_6406);
and U8126 (N_8126,N_6526,N_6903);
nor U8127 (N_8127,N_7460,N_7266);
nor U8128 (N_8128,N_6875,N_7439);
and U8129 (N_8129,N_7399,N_6864);
and U8130 (N_8130,N_6268,N_7276);
xnor U8131 (N_8131,N_7303,N_7232);
or U8132 (N_8132,N_7058,N_6901);
and U8133 (N_8133,N_6998,N_6589);
and U8134 (N_8134,N_6252,N_6572);
nand U8135 (N_8135,N_6944,N_6439);
and U8136 (N_8136,N_6637,N_7267);
nor U8137 (N_8137,N_6681,N_6661);
and U8138 (N_8138,N_7285,N_7028);
nand U8139 (N_8139,N_7259,N_6352);
nor U8140 (N_8140,N_6611,N_6574);
nor U8141 (N_8141,N_6613,N_7299);
and U8142 (N_8142,N_6991,N_7052);
nor U8143 (N_8143,N_6980,N_7187);
and U8144 (N_8144,N_6937,N_6967);
nor U8145 (N_8145,N_6430,N_6691);
nor U8146 (N_8146,N_6318,N_6770);
or U8147 (N_8147,N_6541,N_6849);
nand U8148 (N_8148,N_7458,N_6694);
nand U8149 (N_8149,N_7361,N_6357);
or U8150 (N_8150,N_6946,N_7167);
nor U8151 (N_8151,N_6568,N_6782);
xor U8152 (N_8152,N_6330,N_6295);
or U8153 (N_8153,N_6908,N_7447);
xor U8154 (N_8154,N_7029,N_6323);
nor U8155 (N_8155,N_6504,N_6626);
nor U8156 (N_8156,N_6758,N_7134);
xor U8157 (N_8157,N_6440,N_7490);
or U8158 (N_8158,N_6858,N_6526);
nor U8159 (N_8159,N_7486,N_6820);
nor U8160 (N_8160,N_6581,N_7187);
xnor U8161 (N_8161,N_7114,N_6704);
xnor U8162 (N_8162,N_7125,N_6901);
or U8163 (N_8163,N_6296,N_6437);
or U8164 (N_8164,N_6838,N_6259);
and U8165 (N_8165,N_7141,N_7369);
nand U8166 (N_8166,N_6602,N_6761);
and U8167 (N_8167,N_6977,N_6965);
or U8168 (N_8168,N_6585,N_7393);
nor U8169 (N_8169,N_6258,N_6859);
nand U8170 (N_8170,N_7398,N_6947);
nor U8171 (N_8171,N_6638,N_6931);
nor U8172 (N_8172,N_7441,N_6571);
xnor U8173 (N_8173,N_7079,N_6383);
nand U8174 (N_8174,N_6617,N_7219);
nor U8175 (N_8175,N_7331,N_6777);
xnor U8176 (N_8176,N_6836,N_7249);
nor U8177 (N_8177,N_6979,N_7429);
nand U8178 (N_8178,N_6510,N_7375);
or U8179 (N_8179,N_7351,N_6875);
nor U8180 (N_8180,N_6482,N_6743);
and U8181 (N_8181,N_6444,N_7008);
and U8182 (N_8182,N_7087,N_7297);
or U8183 (N_8183,N_6258,N_6275);
nor U8184 (N_8184,N_6624,N_7212);
xnor U8185 (N_8185,N_6527,N_7422);
xor U8186 (N_8186,N_7219,N_6931);
or U8187 (N_8187,N_7187,N_6311);
nand U8188 (N_8188,N_6608,N_7365);
nor U8189 (N_8189,N_6273,N_7251);
xor U8190 (N_8190,N_6695,N_7333);
and U8191 (N_8191,N_7228,N_7156);
nand U8192 (N_8192,N_6784,N_7485);
nand U8193 (N_8193,N_7427,N_7387);
xnor U8194 (N_8194,N_6938,N_7296);
nor U8195 (N_8195,N_7178,N_6986);
or U8196 (N_8196,N_6742,N_6327);
nand U8197 (N_8197,N_6421,N_6393);
nor U8198 (N_8198,N_6959,N_6500);
xor U8199 (N_8199,N_6474,N_7323);
and U8200 (N_8200,N_6975,N_6579);
nor U8201 (N_8201,N_7279,N_6825);
or U8202 (N_8202,N_6583,N_7208);
nand U8203 (N_8203,N_6890,N_7383);
xnor U8204 (N_8204,N_6878,N_6909);
and U8205 (N_8205,N_7230,N_6433);
nand U8206 (N_8206,N_6472,N_6922);
xnor U8207 (N_8207,N_6513,N_7126);
nand U8208 (N_8208,N_7264,N_6586);
nand U8209 (N_8209,N_7178,N_6980);
nor U8210 (N_8210,N_6893,N_7021);
xnor U8211 (N_8211,N_7118,N_6313);
nand U8212 (N_8212,N_7142,N_7335);
and U8213 (N_8213,N_6975,N_6729);
nor U8214 (N_8214,N_7484,N_7431);
and U8215 (N_8215,N_6450,N_6655);
nor U8216 (N_8216,N_6957,N_6338);
nor U8217 (N_8217,N_6422,N_6643);
nand U8218 (N_8218,N_6635,N_6497);
xor U8219 (N_8219,N_7325,N_7172);
nor U8220 (N_8220,N_6804,N_7427);
xor U8221 (N_8221,N_7261,N_6857);
nor U8222 (N_8222,N_6751,N_6654);
and U8223 (N_8223,N_6683,N_6657);
xnor U8224 (N_8224,N_6688,N_6526);
or U8225 (N_8225,N_6607,N_6699);
xor U8226 (N_8226,N_7208,N_6650);
or U8227 (N_8227,N_6424,N_6629);
or U8228 (N_8228,N_7091,N_6720);
nor U8229 (N_8229,N_6522,N_6825);
nor U8230 (N_8230,N_7304,N_6488);
and U8231 (N_8231,N_6969,N_7391);
nor U8232 (N_8232,N_6674,N_7019);
nand U8233 (N_8233,N_7355,N_6391);
xnor U8234 (N_8234,N_7042,N_6634);
and U8235 (N_8235,N_7388,N_6307);
nand U8236 (N_8236,N_7126,N_7420);
nor U8237 (N_8237,N_6274,N_7137);
nor U8238 (N_8238,N_7321,N_6400);
xor U8239 (N_8239,N_7082,N_6609);
nand U8240 (N_8240,N_6373,N_6764);
nand U8241 (N_8241,N_7270,N_6308);
or U8242 (N_8242,N_7152,N_7167);
nor U8243 (N_8243,N_6834,N_6532);
or U8244 (N_8244,N_6436,N_7351);
and U8245 (N_8245,N_6710,N_6963);
or U8246 (N_8246,N_6649,N_6716);
or U8247 (N_8247,N_6933,N_6551);
nor U8248 (N_8248,N_6296,N_7448);
and U8249 (N_8249,N_7228,N_7465);
or U8250 (N_8250,N_7374,N_6994);
and U8251 (N_8251,N_7109,N_7493);
nand U8252 (N_8252,N_6560,N_6366);
nor U8253 (N_8253,N_6809,N_6418);
xnor U8254 (N_8254,N_6835,N_6254);
or U8255 (N_8255,N_6257,N_6329);
nand U8256 (N_8256,N_6802,N_7166);
nand U8257 (N_8257,N_6287,N_7087);
nor U8258 (N_8258,N_7250,N_7410);
nor U8259 (N_8259,N_7383,N_7110);
and U8260 (N_8260,N_6389,N_6533);
xnor U8261 (N_8261,N_6925,N_7477);
nand U8262 (N_8262,N_6786,N_7485);
and U8263 (N_8263,N_7330,N_6755);
or U8264 (N_8264,N_6335,N_7064);
and U8265 (N_8265,N_7215,N_6284);
and U8266 (N_8266,N_6677,N_7072);
xnor U8267 (N_8267,N_6922,N_6593);
nand U8268 (N_8268,N_6713,N_6601);
and U8269 (N_8269,N_6522,N_6421);
nor U8270 (N_8270,N_6607,N_6531);
nand U8271 (N_8271,N_6623,N_6347);
and U8272 (N_8272,N_7498,N_6952);
or U8273 (N_8273,N_6569,N_7260);
xnor U8274 (N_8274,N_6842,N_6258);
nor U8275 (N_8275,N_6416,N_7345);
or U8276 (N_8276,N_6685,N_6775);
and U8277 (N_8277,N_6990,N_6811);
and U8278 (N_8278,N_7446,N_7225);
or U8279 (N_8279,N_6422,N_7085);
nand U8280 (N_8280,N_6849,N_6390);
or U8281 (N_8281,N_6866,N_6513);
or U8282 (N_8282,N_6604,N_6713);
nor U8283 (N_8283,N_7018,N_6521);
xor U8284 (N_8284,N_6272,N_7286);
and U8285 (N_8285,N_6668,N_7017);
nor U8286 (N_8286,N_7248,N_6992);
nor U8287 (N_8287,N_6883,N_7125);
nand U8288 (N_8288,N_6310,N_6548);
nor U8289 (N_8289,N_7071,N_6283);
or U8290 (N_8290,N_7231,N_7434);
and U8291 (N_8291,N_6328,N_7021);
nand U8292 (N_8292,N_7248,N_7268);
and U8293 (N_8293,N_6366,N_7113);
nand U8294 (N_8294,N_6275,N_7203);
nor U8295 (N_8295,N_6520,N_6871);
nand U8296 (N_8296,N_6895,N_7155);
nor U8297 (N_8297,N_7250,N_6618);
nor U8298 (N_8298,N_7287,N_6340);
and U8299 (N_8299,N_6828,N_6505);
and U8300 (N_8300,N_7211,N_6532);
xor U8301 (N_8301,N_6407,N_6986);
nand U8302 (N_8302,N_7184,N_6362);
and U8303 (N_8303,N_7261,N_6783);
or U8304 (N_8304,N_7366,N_6647);
and U8305 (N_8305,N_6877,N_7003);
or U8306 (N_8306,N_6890,N_6970);
and U8307 (N_8307,N_7206,N_6250);
nor U8308 (N_8308,N_6878,N_7448);
nand U8309 (N_8309,N_6725,N_7272);
and U8310 (N_8310,N_7487,N_6631);
xor U8311 (N_8311,N_7448,N_7181);
nor U8312 (N_8312,N_7330,N_7438);
or U8313 (N_8313,N_6354,N_7342);
nor U8314 (N_8314,N_7023,N_6536);
xnor U8315 (N_8315,N_7396,N_6292);
and U8316 (N_8316,N_7117,N_7114);
nand U8317 (N_8317,N_6657,N_6978);
and U8318 (N_8318,N_7475,N_6375);
xnor U8319 (N_8319,N_7382,N_6385);
nor U8320 (N_8320,N_6759,N_6494);
or U8321 (N_8321,N_6394,N_6267);
and U8322 (N_8322,N_7316,N_7177);
nor U8323 (N_8323,N_6912,N_6965);
xor U8324 (N_8324,N_7161,N_7254);
nor U8325 (N_8325,N_7378,N_7349);
xnor U8326 (N_8326,N_7258,N_7415);
nor U8327 (N_8327,N_6708,N_6443);
xnor U8328 (N_8328,N_7330,N_6371);
xnor U8329 (N_8329,N_6828,N_6914);
xor U8330 (N_8330,N_7482,N_6704);
or U8331 (N_8331,N_7431,N_7233);
xnor U8332 (N_8332,N_6882,N_6774);
xnor U8333 (N_8333,N_6593,N_6745);
xnor U8334 (N_8334,N_7265,N_7424);
nand U8335 (N_8335,N_7459,N_6254);
nand U8336 (N_8336,N_7206,N_7091);
xnor U8337 (N_8337,N_6859,N_7173);
nor U8338 (N_8338,N_6976,N_7466);
xor U8339 (N_8339,N_6583,N_6630);
and U8340 (N_8340,N_6964,N_6460);
xor U8341 (N_8341,N_6716,N_7377);
nand U8342 (N_8342,N_7026,N_7480);
or U8343 (N_8343,N_6540,N_6601);
xor U8344 (N_8344,N_6439,N_7345);
and U8345 (N_8345,N_7186,N_7250);
nor U8346 (N_8346,N_6663,N_6683);
nand U8347 (N_8347,N_7070,N_7092);
and U8348 (N_8348,N_6377,N_7287);
xor U8349 (N_8349,N_6910,N_6794);
and U8350 (N_8350,N_7412,N_7443);
and U8351 (N_8351,N_7021,N_6927);
or U8352 (N_8352,N_6950,N_7206);
nand U8353 (N_8353,N_6687,N_7246);
and U8354 (N_8354,N_6314,N_6717);
or U8355 (N_8355,N_7385,N_6628);
or U8356 (N_8356,N_7044,N_6400);
or U8357 (N_8357,N_6330,N_6329);
nor U8358 (N_8358,N_6313,N_6665);
or U8359 (N_8359,N_7428,N_7405);
or U8360 (N_8360,N_7013,N_6615);
or U8361 (N_8361,N_7103,N_7481);
or U8362 (N_8362,N_7184,N_7248);
nor U8363 (N_8363,N_6995,N_7211);
nand U8364 (N_8364,N_7330,N_6938);
and U8365 (N_8365,N_7190,N_7397);
nand U8366 (N_8366,N_7279,N_6793);
xor U8367 (N_8367,N_6348,N_6763);
xnor U8368 (N_8368,N_6566,N_6730);
or U8369 (N_8369,N_7235,N_6419);
nand U8370 (N_8370,N_7233,N_6582);
or U8371 (N_8371,N_6770,N_7151);
or U8372 (N_8372,N_6940,N_6936);
nor U8373 (N_8373,N_6896,N_7484);
and U8374 (N_8374,N_6397,N_7242);
nor U8375 (N_8375,N_6556,N_6404);
and U8376 (N_8376,N_7407,N_7059);
and U8377 (N_8377,N_7341,N_7022);
nor U8378 (N_8378,N_7335,N_6619);
or U8379 (N_8379,N_7125,N_6473);
nand U8380 (N_8380,N_6537,N_7023);
nand U8381 (N_8381,N_7340,N_7401);
or U8382 (N_8382,N_7092,N_6534);
xor U8383 (N_8383,N_6328,N_6670);
xnor U8384 (N_8384,N_7197,N_6395);
and U8385 (N_8385,N_6727,N_7318);
nor U8386 (N_8386,N_7258,N_6810);
and U8387 (N_8387,N_6897,N_7430);
and U8388 (N_8388,N_6635,N_7294);
and U8389 (N_8389,N_6488,N_6446);
xor U8390 (N_8390,N_6842,N_7377);
and U8391 (N_8391,N_6925,N_6676);
or U8392 (N_8392,N_7049,N_6326);
xor U8393 (N_8393,N_7003,N_6644);
xor U8394 (N_8394,N_6913,N_6592);
and U8395 (N_8395,N_6682,N_6710);
nor U8396 (N_8396,N_7153,N_6675);
or U8397 (N_8397,N_7350,N_6480);
and U8398 (N_8398,N_6350,N_7076);
nand U8399 (N_8399,N_6889,N_7144);
nor U8400 (N_8400,N_6402,N_7085);
nor U8401 (N_8401,N_6735,N_6384);
nor U8402 (N_8402,N_6659,N_6957);
or U8403 (N_8403,N_6713,N_7495);
nor U8404 (N_8404,N_6324,N_7276);
nor U8405 (N_8405,N_7039,N_6377);
xor U8406 (N_8406,N_6330,N_7499);
xnor U8407 (N_8407,N_6732,N_6316);
xor U8408 (N_8408,N_7317,N_6595);
and U8409 (N_8409,N_6828,N_7288);
nor U8410 (N_8410,N_6995,N_6667);
nor U8411 (N_8411,N_6353,N_7014);
nor U8412 (N_8412,N_6471,N_6254);
nand U8413 (N_8413,N_7279,N_6877);
or U8414 (N_8414,N_6803,N_7159);
or U8415 (N_8415,N_7499,N_7082);
nand U8416 (N_8416,N_6383,N_6326);
and U8417 (N_8417,N_6412,N_6345);
and U8418 (N_8418,N_7292,N_7287);
nand U8419 (N_8419,N_6912,N_6309);
nor U8420 (N_8420,N_7220,N_6891);
xor U8421 (N_8421,N_7002,N_7067);
nor U8422 (N_8422,N_6818,N_7411);
and U8423 (N_8423,N_6873,N_7135);
or U8424 (N_8424,N_6614,N_6386);
and U8425 (N_8425,N_6649,N_7383);
xnor U8426 (N_8426,N_6721,N_6459);
and U8427 (N_8427,N_7354,N_6334);
or U8428 (N_8428,N_7299,N_7358);
xnor U8429 (N_8429,N_6264,N_6812);
xor U8430 (N_8430,N_6613,N_7251);
xnor U8431 (N_8431,N_6866,N_6459);
nor U8432 (N_8432,N_6629,N_7318);
or U8433 (N_8433,N_6940,N_7083);
xor U8434 (N_8434,N_7050,N_6419);
nand U8435 (N_8435,N_6508,N_7138);
and U8436 (N_8436,N_6525,N_6981);
or U8437 (N_8437,N_6967,N_6627);
xnor U8438 (N_8438,N_6500,N_6321);
nor U8439 (N_8439,N_6403,N_6534);
nor U8440 (N_8440,N_6765,N_6890);
and U8441 (N_8441,N_7450,N_6580);
or U8442 (N_8442,N_7241,N_6591);
or U8443 (N_8443,N_6540,N_6470);
xor U8444 (N_8444,N_7173,N_6397);
nor U8445 (N_8445,N_7264,N_7140);
or U8446 (N_8446,N_7489,N_7226);
xnor U8447 (N_8447,N_6774,N_7291);
and U8448 (N_8448,N_6970,N_6559);
nand U8449 (N_8449,N_6804,N_7187);
or U8450 (N_8450,N_7364,N_6423);
and U8451 (N_8451,N_6987,N_6561);
nand U8452 (N_8452,N_6478,N_7338);
and U8453 (N_8453,N_6316,N_7427);
nand U8454 (N_8454,N_7122,N_6549);
xor U8455 (N_8455,N_6336,N_6646);
xor U8456 (N_8456,N_6573,N_7415);
xor U8457 (N_8457,N_6703,N_6831);
nand U8458 (N_8458,N_7278,N_6651);
and U8459 (N_8459,N_6724,N_6570);
xor U8460 (N_8460,N_7365,N_7457);
or U8461 (N_8461,N_6931,N_7194);
nor U8462 (N_8462,N_6795,N_6702);
nand U8463 (N_8463,N_6730,N_6660);
nand U8464 (N_8464,N_6580,N_7259);
and U8465 (N_8465,N_6783,N_6858);
and U8466 (N_8466,N_6647,N_6264);
nand U8467 (N_8467,N_6389,N_6419);
nor U8468 (N_8468,N_7195,N_7186);
nor U8469 (N_8469,N_6804,N_7039);
nor U8470 (N_8470,N_6362,N_6604);
nand U8471 (N_8471,N_7310,N_7372);
xnor U8472 (N_8472,N_7189,N_7064);
or U8473 (N_8473,N_6446,N_6274);
nand U8474 (N_8474,N_7144,N_7376);
xor U8475 (N_8475,N_6857,N_6781);
and U8476 (N_8476,N_7214,N_6488);
nor U8477 (N_8477,N_6693,N_6289);
nand U8478 (N_8478,N_7235,N_6803);
xor U8479 (N_8479,N_7308,N_7380);
and U8480 (N_8480,N_7059,N_7231);
xnor U8481 (N_8481,N_6404,N_7171);
nand U8482 (N_8482,N_7384,N_7310);
xor U8483 (N_8483,N_6567,N_6392);
and U8484 (N_8484,N_7244,N_6629);
or U8485 (N_8485,N_7208,N_6263);
nand U8486 (N_8486,N_7318,N_6660);
or U8487 (N_8487,N_6984,N_6774);
and U8488 (N_8488,N_6391,N_7497);
and U8489 (N_8489,N_6918,N_6801);
or U8490 (N_8490,N_7249,N_6768);
nor U8491 (N_8491,N_6256,N_7040);
or U8492 (N_8492,N_7436,N_6411);
and U8493 (N_8493,N_7443,N_6532);
or U8494 (N_8494,N_6573,N_6272);
nor U8495 (N_8495,N_6390,N_6659);
nand U8496 (N_8496,N_7175,N_6945);
nor U8497 (N_8497,N_7100,N_7278);
and U8498 (N_8498,N_7106,N_7469);
nand U8499 (N_8499,N_7344,N_7095);
and U8500 (N_8500,N_6937,N_7414);
xnor U8501 (N_8501,N_7030,N_6626);
or U8502 (N_8502,N_7218,N_6573);
and U8503 (N_8503,N_7434,N_6705);
nand U8504 (N_8504,N_6717,N_7495);
and U8505 (N_8505,N_6992,N_6312);
nand U8506 (N_8506,N_7439,N_6437);
and U8507 (N_8507,N_7302,N_6585);
or U8508 (N_8508,N_7239,N_6937);
nor U8509 (N_8509,N_7383,N_6504);
xnor U8510 (N_8510,N_7033,N_6805);
nor U8511 (N_8511,N_6254,N_6939);
nor U8512 (N_8512,N_6769,N_6479);
xnor U8513 (N_8513,N_6966,N_6913);
xnor U8514 (N_8514,N_6499,N_6728);
or U8515 (N_8515,N_6671,N_6673);
or U8516 (N_8516,N_7217,N_6419);
nand U8517 (N_8517,N_7245,N_6397);
or U8518 (N_8518,N_7397,N_6644);
or U8519 (N_8519,N_7113,N_6996);
nor U8520 (N_8520,N_6397,N_6273);
xor U8521 (N_8521,N_6661,N_7296);
nor U8522 (N_8522,N_7221,N_6994);
nor U8523 (N_8523,N_6621,N_6467);
nor U8524 (N_8524,N_6953,N_7150);
and U8525 (N_8525,N_6493,N_6782);
nand U8526 (N_8526,N_6543,N_6335);
nand U8527 (N_8527,N_6570,N_6996);
nor U8528 (N_8528,N_6705,N_6574);
nand U8529 (N_8529,N_6504,N_6972);
nand U8530 (N_8530,N_7419,N_7037);
or U8531 (N_8531,N_6712,N_6928);
or U8532 (N_8532,N_6465,N_7238);
and U8533 (N_8533,N_6718,N_7344);
xor U8534 (N_8534,N_7478,N_7060);
xnor U8535 (N_8535,N_6925,N_7148);
and U8536 (N_8536,N_6649,N_6579);
xnor U8537 (N_8537,N_6611,N_6588);
nand U8538 (N_8538,N_6881,N_6556);
xor U8539 (N_8539,N_7112,N_6618);
xnor U8540 (N_8540,N_6616,N_7408);
or U8541 (N_8541,N_7434,N_6883);
xor U8542 (N_8542,N_6781,N_6459);
nand U8543 (N_8543,N_6856,N_6925);
nor U8544 (N_8544,N_6473,N_6867);
nand U8545 (N_8545,N_7396,N_6760);
or U8546 (N_8546,N_6488,N_7432);
nor U8547 (N_8547,N_6518,N_7453);
nand U8548 (N_8548,N_7451,N_6670);
nand U8549 (N_8549,N_6447,N_6483);
and U8550 (N_8550,N_6884,N_6622);
xor U8551 (N_8551,N_7037,N_6588);
or U8552 (N_8552,N_7178,N_7034);
xor U8553 (N_8553,N_6516,N_6702);
xor U8554 (N_8554,N_6937,N_6437);
nand U8555 (N_8555,N_6635,N_7021);
or U8556 (N_8556,N_7302,N_6620);
and U8557 (N_8557,N_6836,N_6418);
xnor U8558 (N_8558,N_6274,N_6693);
or U8559 (N_8559,N_7208,N_6717);
or U8560 (N_8560,N_6829,N_7089);
nand U8561 (N_8561,N_7071,N_6553);
and U8562 (N_8562,N_6622,N_7104);
nor U8563 (N_8563,N_6256,N_6435);
xor U8564 (N_8564,N_6495,N_7396);
nor U8565 (N_8565,N_7014,N_7298);
nand U8566 (N_8566,N_6321,N_6769);
and U8567 (N_8567,N_6980,N_6954);
and U8568 (N_8568,N_7389,N_7273);
nor U8569 (N_8569,N_6752,N_6804);
or U8570 (N_8570,N_6306,N_7296);
xor U8571 (N_8571,N_7117,N_6610);
nand U8572 (N_8572,N_6418,N_6511);
or U8573 (N_8573,N_6961,N_6790);
and U8574 (N_8574,N_7223,N_7068);
nand U8575 (N_8575,N_6579,N_6687);
nor U8576 (N_8576,N_7394,N_6705);
xnor U8577 (N_8577,N_6997,N_6509);
xnor U8578 (N_8578,N_6473,N_7407);
or U8579 (N_8579,N_6435,N_6295);
xor U8580 (N_8580,N_7035,N_7487);
nor U8581 (N_8581,N_7055,N_6904);
xor U8582 (N_8582,N_7199,N_7437);
nand U8583 (N_8583,N_7299,N_6566);
and U8584 (N_8584,N_7493,N_7131);
xnor U8585 (N_8585,N_6886,N_7257);
xor U8586 (N_8586,N_7367,N_6606);
and U8587 (N_8587,N_7056,N_7090);
and U8588 (N_8588,N_6695,N_6885);
nand U8589 (N_8589,N_6726,N_7325);
xor U8590 (N_8590,N_7499,N_7420);
nand U8591 (N_8591,N_6644,N_6610);
nand U8592 (N_8592,N_6356,N_6855);
or U8593 (N_8593,N_6866,N_7347);
nor U8594 (N_8594,N_7143,N_6460);
nor U8595 (N_8595,N_6692,N_6999);
and U8596 (N_8596,N_6638,N_7030);
and U8597 (N_8597,N_6822,N_6702);
or U8598 (N_8598,N_7358,N_7263);
xnor U8599 (N_8599,N_6695,N_6796);
xor U8600 (N_8600,N_7115,N_6865);
nor U8601 (N_8601,N_6338,N_7392);
nand U8602 (N_8602,N_6493,N_7198);
xnor U8603 (N_8603,N_6751,N_6332);
and U8604 (N_8604,N_6582,N_7133);
and U8605 (N_8605,N_6894,N_6616);
nand U8606 (N_8606,N_6436,N_7042);
nor U8607 (N_8607,N_7374,N_7341);
and U8608 (N_8608,N_6523,N_6819);
nand U8609 (N_8609,N_6261,N_6501);
or U8610 (N_8610,N_7037,N_6382);
nand U8611 (N_8611,N_6336,N_7068);
xor U8612 (N_8612,N_6431,N_6766);
xor U8613 (N_8613,N_6881,N_7418);
nand U8614 (N_8614,N_7081,N_6706);
nand U8615 (N_8615,N_6808,N_7323);
or U8616 (N_8616,N_6699,N_6895);
nor U8617 (N_8617,N_6817,N_7423);
xor U8618 (N_8618,N_6858,N_6630);
nand U8619 (N_8619,N_6964,N_7063);
or U8620 (N_8620,N_7323,N_6732);
xnor U8621 (N_8621,N_6273,N_7170);
nor U8622 (N_8622,N_6326,N_6601);
nand U8623 (N_8623,N_7326,N_6879);
and U8624 (N_8624,N_7018,N_6442);
or U8625 (N_8625,N_6572,N_7054);
and U8626 (N_8626,N_7253,N_6560);
and U8627 (N_8627,N_7415,N_6679);
or U8628 (N_8628,N_7312,N_7063);
nor U8629 (N_8629,N_7315,N_6407);
or U8630 (N_8630,N_7179,N_6481);
nand U8631 (N_8631,N_7100,N_6304);
nand U8632 (N_8632,N_7372,N_6571);
or U8633 (N_8633,N_7190,N_6294);
xor U8634 (N_8634,N_6480,N_6677);
xor U8635 (N_8635,N_7486,N_6866);
xnor U8636 (N_8636,N_7250,N_7359);
nand U8637 (N_8637,N_7337,N_7272);
nor U8638 (N_8638,N_6649,N_7376);
xnor U8639 (N_8639,N_6278,N_7269);
nand U8640 (N_8640,N_6406,N_7403);
and U8641 (N_8641,N_6294,N_7110);
nand U8642 (N_8642,N_6253,N_6580);
xor U8643 (N_8643,N_6856,N_7294);
or U8644 (N_8644,N_6955,N_6460);
nand U8645 (N_8645,N_6764,N_7228);
xor U8646 (N_8646,N_7460,N_7478);
and U8647 (N_8647,N_7230,N_6709);
xor U8648 (N_8648,N_6702,N_6758);
or U8649 (N_8649,N_7401,N_7493);
and U8650 (N_8650,N_6770,N_7233);
nor U8651 (N_8651,N_6708,N_6536);
nand U8652 (N_8652,N_6617,N_7042);
or U8653 (N_8653,N_7007,N_6469);
nor U8654 (N_8654,N_7268,N_6949);
nand U8655 (N_8655,N_7416,N_6399);
nand U8656 (N_8656,N_7124,N_7267);
nor U8657 (N_8657,N_6454,N_7325);
xnor U8658 (N_8658,N_6251,N_7346);
nand U8659 (N_8659,N_7001,N_7345);
xnor U8660 (N_8660,N_7134,N_6458);
xnor U8661 (N_8661,N_6286,N_6377);
nand U8662 (N_8662,N_6588,N_7402);
and U8663 (N_8663,N_6434,N_6963);
or U8664 (N_8664,N_7336,N_6885);
and U8665 (N_8665,N_6357,N_7052);
or U8666 (N_8666,N_6643,N_6439);
xor U8667 (N_8667,N_6809,N_6533);
xor U8668 (N_8668,N_7044,N_6418);
and U8669 (N_8669,N_6899,N_7217);
nor U8670 (N_8670,N_7305,N_7278);
and U8671 (N_8671,N_6755,N_7035);
nand U8672 (N_8672,N_6368,N_7093);
xor U8673 (N_8673,N_6260,N_6550);
nor U8674 (N_8674,N_7064,N_6779);
nand U8675 (N_8675,N_6461,N_7372);
or U8676 (N_8676,N_6470,N_6621);
nor U8677 (N_8677,N_6489,N_7479);
nand U8678 (N_8678,N_7224,N_7391);
nor U8679 (N_8679,N_7058,N_6700);
xor U8680 (N_8680,N_7310,N_7266);
or U8681 (N_8681,N_6697,N_7458);
nor U8682 (N_8682,N_7375,N_7125);
and U8683 (N_8683,N_7319,N_6460);
nor U8684 (N_8684,N_7003,N_7189);
nand U8685 (N_8685,N_7493,N_6820);
xor U8686 (N_8686,N_6644,N_6808);
xnor U8687 (N_8687,N_7332,N_7197);
xor U8688 (N_8688,N_7450,N_6487);
and U8689 (N_8689,N_6873,N_7134);
nand U8690 (N_8690,N_7087,N_6311);
or U8691 (N_8691,N_6955,N_6865);
nand U8692 (N_8692,N_6477,N_7141);
and U8693 (N_8693,N_6658,N_7108);
xor U8694 (N_8694,N_6461,N_7232);
xor U8695 (N_8695,N_7247,N_7373);
or U8696 (N_8696,N_6844,N_6684);
or U8697 (N_8697,N_6948,N_7264);
nor U8698 (N_8698,N_6720,N_6364);
nand U8699 (N_8699,N_6408,N_7330);
or U8700 (N_8700,N_6314,N_6557);
or U8701 (N_8701,N_6474,N_6899);
nor U8702 (N_8702,N_6270,N_7081);
xnor U8703 (N_8703,N_6464,N_6419);
nand U8704 (N_8704,N_6310,N_6281);
xor U8705 (N_8705,N_6929,N_6320);
nor U8706 (N_8706,N_7217,N_6826);
or U8707 (N_8707,N_6825,N_6346);
nor U8708 (N_8708,N_6834,N_7145);
xnor U8709 (N_8709,N_6575,N_6401);
or U8710 (N_8710,N_7019,N_6291);
nand U8711 (N_8711,N_6668,N_7282);
or U8712 (N_8712,N_7066,N_7188);
xor U8713 (N_8713,N_7142,N_6548);
or U8714 (N_8714,N_6985,N_6425);
xor U8715 (N_8715,N_6810,N_7450);
or U8716 (N_8716,N_6830,N_6488);
nand U8717 (N_8717,N_6646,N_7145);
xor U8718 (N_8718,N_6506,N_6720);
xor U8719 (N_8719,N_6586,N_7055);
or U8720 (N_8720,N_7096,N_6955);
nand U8721 (N_8721,N_7226,N_6292);
or U8722 (N_8722,N_7316,N_7203);
or U8723 (N_8723,N_6581,N_7189);
and U8724 (N_8724,N_6898,N_7337);
nor U8725 (N_8725,N_7397,N_6546);
or U8726 (N_8726,N_6913,N_6550);
nand U8727 (N_8727,N_6714,N_6946);
nand U8728 (N_8728,N_7209,N_6434);
and U8729 (N_8729,N_7140,N_7243);
nand U8730 (N_8730,N_7199,N_6392);
and U8731 (N_8731,N_6559,N_6303);
xor U8732 (N_8732,N_6410,N_6669);
nand U8733 (N_8733,N_7481,N_7492);
or U8734 (N_8734,N_6561,N_7228);
xor U8735 (N_8735,N_6344,N_7197);
and U8736 (N_8736,N_6884,N_6256);
nor U8737 (N_8737,N_7365,N_6280);
nor U8738 (N_8738,N_7312,N_6478);
xnor U8739 (N_8739,N_7221,N_7021);
xnor U8740 (N_8740,N_7067,N_6545);
nor U8741 (N_8741,N_6446,N_6776);
nor U8742 (N_8742,N_7035,N_6815);
xor U8743 (N_8743,N_7435,N_7357);
nand U8744 (N_8744,N_6772,N_7094);
and U8745 (N_8745,N_6346,N_6909);
or U8746 (N_8746,N_7052,N_7134);
and U8747 (N_8747,N_6280,N_7098);
nand U8748 (N_8748,N_6881,N_6707);
xnor U8749 (N_8749,N_7399,N_7370);
or U8750 (N_8750,N_8736,N_7895);
nor U8751 (N_8751,N_8096,N_8403);
and U8752 (N_8752,N_8019,N_8347);
xnor U8753 (N_8753,N_7504,N_8581);
nor U8754 (N_8754,N_8430,N_7742);
and U8755 (N_8755,N_7637,N_8364);
nand U8756 (N_8756,N_8421,N_8393);
xor U8757 (N_8757,N_7990,N_7976);
and U8758 (N_8758,N_8638,N_8556);
or U8759 (N_8759,N_7739,N_7508);
xor U8760 (N_8760,N_8548,N_8157);
nor U8761 (N_8761,N_8398,N_8708);
nand U8762 (N_8762,N_8582,N_8433);
and U8763 (N_8763,N_7845,N_7623);
or U8764 (N_8764,N_8272,N_8574);
and U8765 (N_8765,N_8667,N_8693);
nor U8766 (N_8766,N_7756,N_8061);
and U8767 (N_8767,N_7596,N_8731);
and U8768 (N_8768,N_7560,N_7527);
and U8769 (N_8769,N_7725,N_7803);
or U8770 (N_8770,N_8609,N_7599);
nand U8771 (N_8771,N_8559,N_8400);
nand U8772 (N_8772,N_7606,N_7751);
nor U8773 (N_8773,N_8237,N_8102);
nand U8774 (N_8774,N_8217,N_8098);
nor U8775 (N_8775,N_7771,N_8128);
nor U8776 (N_8776,N_8070,N_7899);
nor U8777 (N_8777,N_8447,N_8535);
or U8778 (N_8778,N_7592,N_7589);
or U8779 (N_8779,N_8345,N_8058);
or U8780 (N_8780,N_7620,N_8629);
and U8781 (N_8781,N_7965,N_8044);
and U8782 (N_8782,N_7854,N_8442);
xnor U8783 (N_8783,N_7827,N_7883);
nand U8784 (N_8784,N_8072,N_8225);
nand U8785 (N_8785,N_7544,N_7554);
xnor U8786 (N_8786,N_7992,N_8627);
xnor U8787 (N_8787,N_8181,N_8579);
nor U8788 (N_8788,N_8562,N_8317);
or U8789 (N_8789,N_7839,N_7962);
and U8790 (N_8790,N_8195,N_8684);
nor U8791 (N_8791,N_8606,N_7915);
nand U8792 (N_8792,N_7831,N_7678);
nor U8793 (N_8793,N_7891,N_7706);
and U8794 (N_8794,N_7900,N_8445);
and U8795 (N_8795,N_7963,N_7598);
nand U8796 (N_8796,N_8049,N_8645);
nand U8797 (N_8797,N_8482,N_8372);
nor U8798 (N_8798,N_7987,N_8135);
and U8799 (N_8799,N_7846,N_8504);
or U8800 (N_8800,N_8005,N_8122);
or U8801 (N_8801,N_8196,N_7522);
and U8802 (N_8802,N_8382,N_7741);
or U8803 (N_8803,N_8668,N_8286);
and U8804 (N_8804,N_8730,N_8238);
nor U8805 (N_8805,N_7667,N_8468);
xor U8806 (N_8806,N_8654,N_7828);
nand U8807 (N_8807,N_7796,N_8282);
and U8808 (N_8808,N_7849,N_8264);
xnor U8809 (N_8809,N_7959,N_8322);
xnor U8810 (N_8810,N_8180,N_8614);
or U8811 (N_8811,N_7823,N_7769);
nand U8812 (N_8812,N_7572,N_7733);
nor U8813 (N_8813,N_8649,N_7552);
xor U8814 (N_8814,N_8304,N_7998);
and U8815 (N_8815,N_8594,N_8192);
nor U8816 (N_8816,N_8633,N_8546);
nand U8817 (N_8817,N_8586,N_8306);
and U8818 (N_8818,N_8414,N_8167);
nor U8819 (N_8819,N_8391,N_8675);
nand U8820 (N_8820,N_8682,N_8143);
nor U8821 (N_8821,N_7717,N_7996);
or U8822 (N_8822,N_7541,N_8169);
nand U8823 (N_8823,N_7933,N_8437);
xor U8824 (N_8824,N_7688,N_7981);
xor U8825 (N_8825,N_8734,N_7927);
xnor U8826 (N_8826,N_8114,N_8302);
xor U8827 (N_8827,N_7521,N_8230);
and U8828 (N_8828,N_8462,N_8413);
nor U8829 (N_8829,N_8250,N_8215);
and U8830 (N_8830,N_8045,N_7893);
nand U8831 (N_8831,N_8340,N_8380);
nor U8832 (N_8832,N_8125,N_8078);
xor U8833 (N_8833,N_7906,N_8453);
and U8834 (N_8834,N_8490,N_8310);
or U8835 (N_8835,N_8343,N_7975);
xnor U8836 (N_8836,N_8141,N_8431);
or U8837 (N_8837,N_7749,N_8567);
and U8838 (N_8838,N_7876,N_8226);
or U8839 (N_8839,N_7629,N_7511);
xor U8840 (N_8840,N_8186,N_8625);
or U8841 (N_8841,N_7590,N_7857);
nand U8842 (N_8842,N_7916,N_8362);
xnor U8843 (N_8843,N_7600,N_7533);
xor U8844 (N_8844,N_8580,N_8295);
and U8845 (N_8845,N_7738,N_8725);
or U8846 (N_8846,N_7797,N_7616);
nand U8847 (N_8847,N_8223,N_8626);
and U8848 (N_8848,N_8419,N_7559);
nand U8849 (N_8849,N_7698,N_8274);
and U8850 (N_8850,N_7786,N_8155);
nand U8851 (N_8851,N_8551,N_7960);
xnor U8852 (N_8852,N_7730,N_8086);
or U8853 (N_8853,N_8288,N_8020);
xnor U8854 (N_8854,N_8188,N_8202);
nor U8855 (N_8855,N_8370,N_7978);
xnor U8856 (N_8856,N_7753,N_7806);
nor U8857 (N_8857,N_8591,N_8093);
nand U8858 (N_8858,N_8030,N_7718);
or U8859 (N_8859,N_8227,N_8129);
and U8860 (N_8860,N_8666,N_7687);
nor U8861 (N_8861,N_7826,N_8022);
or U8862 (N_8862,N_8236,N_7999);
xor U8863 (N_8863,N_7563,N_8262);
and U8864 (N_8864,N_8588,N_7997);
nand U8865 (N_8865,N_7701,N_7516);
nand U8866 (N_8866,N_8278,N_8210);
nand U8867 (N_8867,N_7611,N_7682);
nand U8868 (N_8868,N_8385,N_7938);
xor U8869 (N_8869,N_8472,N_8745);
or U8870 (N_8870,N_8464,N_8620);
nor U8871 (N_8871,N_8441,N_8144);
nor U8872 (N_8872,N_8444,N_7856);
or U8873 (N_8873,N_7634,N_7932);
nor U8874 (N_8874,N_8348,N_8240);
nor U8875 (N_8875,N_8248,N_7517);
nor U8876 (N_8876,N_8516,N_8099);
and U8877 (N_8877,N_8432,N_8721);
nand U8878 (N_8878,N_8450,N_7569);
nand U8879 (N_8879,N_8571,N_8583);
nor U8880 (N_8880,N_8212,N_8601);
nor U8881 (N_8881,N_8235,N_7736);
and U8882 (N_8882,N_8694,N_8742);
xor U8883 (N_8883,N_8687,N_8705);
xnor U8884 (N_8884,N_8040,N_8471);
and U8885 (N_8885,N_8252,N_7781);
nor U8886 (N_8886,N_8069,N_8035);
xnor U8887 (N_8887,N_8232,N_8715);
nand U8888 (N_8888,N_7625,N_7822);
nand U8889 (N_8889,N_7852,N_8531);
and U8890 (N_8890,N_8048,N_7529);
xor U8891 (N_8891,N_8162,N_7809);
nor U8892 (N_8892,N_8136,N_7649);
nor U8893 (N_8893,N_8205,N_7807);
nand U8894 (N_8894,N_8229,N_7602);
and U8895 (N_8895,N_8090,N_8085);
and U8896 (N_8896,N_8153,N_7875);
nor U8897 (N_8897,N_8643,N_7984);
xnor U8898 (N_8898,N_7972,N_8368);
and U8899 (N_8899,N_8637,N_7628);
or U8900 (N_8900,N_7608,N_7789);
and U8901 (N_8901,N_8358,N_8405);
or U8902 (N_8902,N_8323,N_8263);
xor U8903 (N_8903,N_7791,N_7673);
nor U8904 (N_8904,N_7581,N_8700);
xnor U8905 (N_8905,N_7524,N_8463);
nor U8906 (N_8906,N_8289,N_8677);
and U8907 (N_8907,N_8259,N_8004);
xor U8908 (N_8908,N_8321,N_7676);
nand U8909 (N_8909,N_8046,N_8602);
nand U8910 (N_8910,N_7635,N_7532);
nor U8911 (N_8911,N_8554,N_8273);
nand U8912 (N_8912,N_7873,N_8543);
or U8913 (N_8913,N_7994,N_8454);
or U8914 (N_8914,N_7523,N_7703);
xor U8915 (N_8915,N_8469,N_7579);
and U8916 (N_8916,N_7993,N_8507);
or U8917 (N_8917,N_8103,N_8168);
and U8918 (N_8918,N_8130,N_7770);
nor U8919 (N_8919,N_7660,N_8477);
nand U8920 (N_8920,N_8569,N_7768);
and U8921 (N_8921,N_8200,N_7897);
nor U8922 (N_8922,N_8294,N_8110);
and U8923 (N_8923,N_8506,N_8006);
and U8924 (N_8924,N_8656,N_7662);
nor U8925 (N_8925,N_8537,N_7652);
or U8926 (N_8926,N_8500,N_8642);
xnor U8927 (N_8927,N_8622,N_8108);
nor U8928 (N_8928,N_7626,N_8630);
or U8929 (N_8929,N_8100,N_7661);
xor U8930 (N_8930,N_7841,N_8529);
nand U8931 (N_8931,N_8170,N_8261);
nor U8932 (N_8932,N_7737,N_8713);
nor U8933 (N_8933,N_8652,N_8399);
xor U8934 (N_8934,N_8644,N_7665);
and U8935 (N_8935,N_7712,N_8679);
nor U8936 (N_8936,N_8239,N_8617);
nand U8937 (N_8937,N_8723,N_7958);
nor U8938 (N_8938,N_7840,N_7956);
nand U8939 (N_8939,N_8204,N_8412);
or U8940 (N_8940,N_8118,N_8467);
nand U8941 (N_8941,N_7886,N_8635);
and U8942 (N_8942,N_8255,N_8658);
xnor U8943 (N_8943,N_7709,N_7744);
and U8944 (N_8944,N_8619,N_8676);
and U8945 (N_8945,N_7758,N_8185);
xnor U8946 (N_8946,N_8147,N_7947);
or U8947 (N_8947,N_8628,N_7808);
nand U8948 (N_8948,N_7639,N_7872);
nor U8949 (N_8949,N_8246,N_7834);
nor U8950 (N_8950,N_8231,N_8401);
xnor U8951 (N_8951,N_8727,N_8697);
nand U8952 (N_8952,N_7812,N_8079);
nand U8953 (N_8953,N_8435,N_8530);
nor U8954 (N_8954,N_8095,N_8423);
xnor U8955 (N_8955,N_8308,N_7892);
nand U8956 (N_8956,N_7862,N_8293);
and U8957 (N_8957,N_7539,N_8316);
or U8958 (N_8958,N_7503,N_8520);
or U8959 (N_8959,N_8363,N_8305);
and U8960 (N_8960,N_8459,N_7815);
or U8961 (N_8961,N_8523,N_8335);
nand U8962 (N_8962,N_8489,N_7818);
nor U8963 (N_8963,N_7939,N_8220);
or U8964 (N_8964,N_8208,N_8497);
nand U8965 (N_8965,N_8493,N_8296);
and U8966 (N_8966,N_8427,N_7550);
nor U8967 (N_8967,N_7804,N_7684);
nand U8968 (N_8968,N_8549,N_8092);
or U8969 (N_8969,N_7842,N_8517);
or U8970 (N_8970,N_8669,N_7868);
nor U8971 (N_8971,N_8483,N_8383);
or U8972 (N_8972,N_7943,N_8542);
or U8973 (N_8973,N_8689,N_8314);
nand U8974 (N_8974,N_8501,N_7750);
nor U8975 (N_8975,N_8164,N_7869);
or U8976 (N_8976,N_8729,N_7545);
nand U8977 (N_8977,N_8244,N_7754);
and U8978 (N_8978,N_8661,N_7685);
or U8979 (N_8979,N_8201,N_7967);
and U8980 (N_8980,N_7775,N_8392);
or U8981 (N_8981,N_7578,N_8320);
nand U8982 (N_8982,N_7830,N_8119);
nand U8983 (N_8983,N_8234,N_7763);
xnor U8984 (N_8984,N_7946,N_8662);
nand U8985 (N_8985,N_8254,N_7735);
xnor U8986 (N_8986,N_8408,N_7704);
nand U8987 (N_8987,N_8284,N_8023);
or U8988 (N_8988,N_7716,N_8175);
or U8989 (N_8989,N_8338,N_8015);
and U8990 (N_8990,N_8659,N_8053);
nor U8991 (N_8991,N_8416,N_8183);
nand U8992 (N_8992,N_8371,N_8142);
nor U8993 (N_8993,N_8434,N_8714);
xnor U8994 (N_8994,N_8233,N_7914);
or U8995 (N_8995,N_7817,N_8508);
and U8996 (N_8996,N_7568,N_7923);
or U8997 (N_8997,N_7924,N_8216);
nor U8998 (N_8998,N_8054,N_7778);
and U8999 (N_8999,N_8566,N_8378);
or U9000 (N_9000,N_8319,N_8356);
nand U9001 (N_9001,N_7723,N_8716);
nor U9002 (N_9002,N_7597,N_7566);
nor U9003 (N_9003,N_7612,N_8366);
and U9004 (N_9004,N_7564,N_7957);
or U9005 (N_9005,N_8440,N_8138);
xnor U9006 (N_9006,N_7764,N_8166);
xor U9007 (N_9007,N_7885,N_8214);
and U9008 (N_9008,N_7908,N_7707);
and U9009 (N_9009,N_7903,N_8140);
xnor U9010 (N_9010,N_7968,N_8448);
or U9011 (N_9011,N_8369,N_7982);
nor U9012 (N_9012,N_7889,N_7510);
and U9013 (N_9013,N_8123,N_8722);
nand U9014 (N_9014,N_7672,N_7874);
nor U9015 (N_9015,N_8397,N_7647);
nand U9016 (N_9016,N_8595,N_8012);
nand U9017 (N_9017,N_7528,N_8080);
nor U9018 (N_9018,N_8124,N_8218);
and U9019 (N_9019,N_7585,N_8115);
xnor U9020 (N_9020,N_8406,N_8299);
nand U9021 (N_9021,N_8749,N_8597);
or U9022 (N_9022,N_7573,N_8060);
xor U9023 (N_9023,N_8038,N_8577);
nor U9024 (N_9024,N_7586,N_7917);
and U9025 (N_9025,N_7871,N_8156);
or U9026 (N_9026,N_7991,N_8065);
xnor U9027 (N_9027,N_7505,N_7697);
xor U9028 (N_9028,N_8094,N_8573);
xnor U9029 (N_9029,N_7980,N_8071);
nor U9030 (N_9030,N_7713,N_8486);
and U9031 (N_9031,N_7593,N_8088);
nor U9032 (N_9032,N_8528,N_8703);
nand U9033 (N_9033,N_8672,N_7913);
or U9034 (N_9034,N_8512,N_7727);
xnor U9035 (N_9035,N_8283,N_8636);
nor U9036 (N_9036,N_8541,N_7636);
nor U9037 (N_9037,N_7577,N_7877);
nand U9038 (N_9038,N_8021,N_7543);
nand U9039 (N_9039,N_7853,N_8726);
and U9040 (N_9040,N_8592,N_8439);
nand U9041 (N_9041,N_7576,N_7832);
xnor U9042 (N_9042,N_7855,N_7512);
or U9043 (N_9043,N_7624,N_7920);
or U9044 (N_9044,N_8076,N_7757);
nor U9045 (N_9045,N_7863,N_7941);
nor U9046 (N_9046,N_7642,N_7617);
xor U9047 (N_9047,N_8488,N_8275);
or U9048 (N_9048,N_7731,N_7691);
xor U9049 (N_9049,N_7977,N_7674);
xor U9050 (N_9050,N_8353,N_8698);
xor U9051 (N_9051,N_7810,N_7940);
xnor U9052 (N_9052,N_7971,N_8010);
or U9053 (N_9053,N_8066,N_7724);
nand U9054 (N_9054,N_7772,N_8671);
nor U9055 (N_9055,N_7621,N_8741);
nor U9056 (N_9056,N_8688,N_8148);
nor U9057 (N_9057,N_7907,N_8270);
nor U9058 (N_9058,N_7710,N_8585);
or U9059 (N_9059,N_7765,N_8470);
nor U9060 (N_9060,N_8707,N_8309);
or U9061 (N_9061,N_7798,N_8436);
xnor U9062 (N_9062,N_8509,N_8267);
xnor U9063 (N_9063,N_7773,N_8561);
and U9064 (N_9064,N_8381,N_8524);
nand U9065 (N_9065,N_8499,N_8326);
xor U9066 (N_9066,N_8134,N_7955);
and U9067 (N_9067,N_8106,N_8055);
nor U9068 (N_9068,N_7513,N_8377);
and U9069 (N_9069,N_8466,N_8558);
or U9070 (N_9070,N_8639,N_8612);
or U9071 (N_9071,N_8605,N_8438);
or U9072 (N_9072,N_8357,N_8105);
nor U9073 (N_9073,N_8355,N_8449);
nand U9074 (N_9074,N_8575,N_8311);
nor U9075 (N_9075,N_8191,N_8495);
nor U9076 (N_9076,N_8075,N_8171);
xor U9077 (N_9077,N_8475,N_8396);
or U9078 (N_9078,N_8172,N_7813);
and U9079 (N_9079,N_7859,N_7861);
nand U9080 (N_9080,N_7699,N_7787);
or U9081 (N_9081,N_7632,N_8187);
nor U9082 (N_9082,N_7670,N_8387);
nor U9083 (N_9083,N_8496,N_7951);
nor U9084 (N_9084,N_8354,N_7909);
xnor U9085 (N_9085,N_7884,N_7879);
nand U9086 (N_9086,N_7515,N_8565);
and U9087 (N_9087,N_7525,N_7887);
or U9088 (N_9088,N_7680,N_8553);
nand U9089 (N_9089,N_8163,N_7575);
nand U9090 (N_9090,N_7986,N_7935);
xor U9091 (N_9091,N_8365,N_7911);
xnor U9092 (N_9092,N_8706,N_7609);
nor U9093 (N_9093,N_7784,N_8374);
nor U9094 (N_9094,N_8618,N_7562);
and U9095 (N_9095,N_7896,N_8117);
xnor U9096 (N_9096,N_8026,N_7705);
nand U9097 (N_9097,N_7549,N_7557);
or U9098 (N_9098,N_7526,N_7546);
or U9099 (N_9099,N_7979,N_7819);
nand U9100 (N_9100,N_7582,N_8315);
and U9101 (N_9101,N_7613,N_7655);
nor U9102 (N_9102,N_7567,N_8271);
xnor U9103 (N_9103,N_7501,N_8456);
and U9104 (N_9104,N_8247,N_7622);
and U9105 (N_9105,N_7881,N_7548);
nor U9106 (N_9106,N_8460,N_8428);
or U9107 (N_9107,N_7752,N_8743);
or U9108 (N_9108,N_8109,N_8131);
nor U9109 (N_9109,N_7766,N_7882);
and U9110 (N_9110,N_7919,N_8177);
nor U9111 (N_9111,N_8064,N_7627);
nor U9112 (N_9112,N_8576,N_8429);
and U9113 (N_9113,N_7767,N_7574);
and U9114 (N_9114,N_8137,N_7558);
nor U9115 (N_9115,N_8718,N_7728);
or U9116 (N_9116,N_8498,N_8532);
or U9117 (N_9117,N_8685,N_7696);
and U9118 (N_9118,N_8279,N_7851);
xnor U9119 (N_9119,N_8402,N_8113);
or U9120 (N_9120,N_8701,N_8663);
xnor U9121 (N_9121,N_8341,N_7777);
nor U9122 (N_9122,N_8557,N_8640);
nand U9123 (N_9123,N_7850,N_7902);
xor U9124 (N_9124,N_8027,N_8728);
or U9125 (N_9125,N_7610,N_7721);
and U9126 (N_9126,N_8717,N_7792);
nor U9127 (N_9127,N_8492,N_8062);
and U9128 (N_9128,N_7565,N_8257);
nor U9129 (N_9129,N_8533,N_8190);
xor U9130 (N_9130,N_8313,N_8184);
nand U9131 (N_9131,N_8199,N_8733);
nand U9132 (N_9132,N_8303,N_8481);
and U9133 (N_9133,N_7983,N_8732);
xor U9134 (N_9134,N_8121,N_8074);
nand U9135 (N_9135,N_7603,N_8158);
or U9136 (N_9136,N_8280,N_7901);
or U9137 (N_9137,N_7714,N_8328);
or U9138 (N_9138,N_8578,N_8511);
nand U9139 (N_9139,N_7934,N_8160);
nor U9140 (N_9140,N_7795,N_8047);
nand U9141 (N_9141,N_8680,N_7748);
nand U9142 (N_9142,N_8329,N_8116);
or U9143 (N_9143,N_7918,N_8545);
and U9144 (N_9144,N_7722,N_7837);
xor U9145 (N_9145,N_8318,N_8526);
nand U9146 (N_9146,N_8352,N_7537);
xor U9147 (N_9147,N_7746,N_8133);
xnor U9148 (N_9148,N_7648,N_8572);
or U9149 (N_9149,N_8446,N_8702);
xor U9150 (N_9150,N_8525,N_7607);
and U9151 (N_9151,N_7843,N_8598);
nand U9152 (N_9152,N_7518,N_7604);
xnor U9153 (N_9153,N_8484,N_8491);
nor U9154 (N_9154,N_7948,N_8394);
or U9155 (N_9155,N_8600,N_8082);
xnor U9156 (N_9156,N_8555,N_8179);
or U9157 (N_9157,N_8300,N_7708);
nand U9158 (N_9158,N_8367,N_7760);
nand U9159 (N_9159,N_7726,N_7502);
xor U9160 (N_9160,N_7780,N_8651);
or U9161 (N_9161,N_8016,N_8349);
nor U9162 (N_9162,N_8710,N_7793);
or U9163 (N_9163,N_7700,N_7618);
xor U9164 (N_9164,N_8424,N_8154);
nand U9165 (N_9165,N_8039,N_7930);
or U9166 (N_9166,N_8540,N_8127);
and U9167 (N_9167,N_8151,N_8384);
nor U9168 (N_9168,N_7534,N_8426);
nor U9169 (N_9169,N_7646,N_8513);
xor U9170 (N_9170,N_8265,N_8521);
and U9171 (N_9171,N_8473,N_7912);
nor U9172 (N_9172,N_8132,N_7776);
nor U9173 (N_9173,N_8691,N_7656);
nand U9174 (N_9174,N_8485,N_8194);
and U9175 (N_9175,N_8389,N_8312);
xor U9176 (N_9176,N_7801,N_8550);
xor U9177 (N_9177,N_8359,N_8037);
nor U9178 (N_9178,N_8111,N_8411);
and U9179 (N_9179,N_7890,N_8740);
nand U9180 (N_9180,N_8712,N_7538);
nor U9181 (N_9181,N_8159,N_8646);
nor U9182 (N_9182,N_7937,N_7694);
xor U9183 (N_9183,N_8388,N_7553);
or U9184 (N_9184,N_7945,N_8018);
and U9185 (N_9185,N_8003,N_8336);
nor U9186 (N_9186,N_8719,N_7650);
nand U9187 (N_9187,N_8126,N_7536);
xnor U9188 (N_9188,N_8258,N_7774);
xor U9189 (N_9189,N_7644,N_8041);
nand U9190 (N_9190,N_7816,N_8476);
or U9191 (N_9191,N_8251,N_7922);
nand U9192 (N_9192,N_8161,N_7734);
xnor U9193 (N_9193,N_8724,N_8692);
xor U9194 (N_9194,N_8266,N_7762);
xnor U9195 (N_9195,N_7580,N_7790);
nor U9196 (N_9196,N_8332,N_7836);
or U9197 (N_9197,N_8560,N_8505);
or U9198 (N_9198,N_7833,N_8410);
or U9199 (N_9199,N_8243,N_8461);
nor U9200 (N_9200,N_8623,N_8425);
nor U9201 (N_9201,N_7936,N_8544);
and U9202 (N_9202,N_8276,N_8634);
nand U9203 (N_9203,N_7729,N_8407);
and U9204 (N_9204,N_8683,N_7942);
nand U9205 (N_9205,N_8334,N_8091);
and U9206 (N_9206,N_7530,N_7657);
and U9207 (N_9207,N_7995,N_8443);
and U9208 (N_9208,N_8197,N_8631);
xor U9209 (N_9209,N_8748,N_8221);
nand U9210 (N_9210,N_8664,N_8145);
and U9211 (N_9211,N_7719,N_8587);
nand U9212 (N_9212,N_8011,N_7535);
nand U9213 (N_9213,N_8379,N_8599);
or U9214 (N_9214,N_8189,N_8547);
nor U9215 (N_9215,N_7785,N_8253);
nand U9216 (N_9216,N_8033,N_8043);
and U9217 (N_9217,N_8327,N_7732);
nand U9218 (N_9218,N_7905,N_7630);
nand U9219 (N_9219,N_8641,N_7556);
xnor U9220 (N_9220,N_7974,N_8590);
nor U9221 (N_9221,N_8665,N_8063);
and U9222 (N_9222,N_8346,N_7858);
nor U9223 (N_9223,N_8324,N_7638);
and U9224 (N_9224,N_8077,N_8522);
or U9225 (N_9225,N_8052,N_7782);
or U9226 (N_9226,N_7878,N_7954);
nand U9227 (N_9227,N_8260,N_8739);
nand U9228 (N_9228,N_8695,N_8285);
or U9229 (N_9229,N_8720,N_8390);
nor U9230 (N_9230,N_7643,N_8696);
or U9231 (N_9231,N_7910,N_8193);
nor U9232 (N_9232,N_8616,N_8593);
and U9233 (N_9233,N_8083,N_7988);
and U9234 (N_9234,N_8107,N_8002);
nor U9235 (N_9235,N_8301,N_7755);
nor U9236 (N_9236,N_7838,N_7659);
nor U9237 (N_9237,N_8084,N_8474);
and U9238 (N_9238,N_8699,N_8059);
or U9239 (N_9239,N_8176,N_8514);
nand U9240 (N_9240,N_7720,N_7966);
and U9241 (N_9241,N_7969,N_8036);
or U9242 (N_9242,N_8607,N_8536);
nor U9243 (N_9243,N_7571,N_7929);
nor U9244 (N_9244,N_8624,N_8650);
or U9245 (N_9245,N_8174,N_7702);
nor U9246 (N_9246,N_7964,N_7615);
nand U9247 (N_9247,N_8219,N_8744);
or U9248 (N_9248,N_7799,N_8632);
xor U9249 (N_9249,N_8350,N_8417);
nand U9250 (N_9250,N_7689,N_8452);
nor U9251 (N_9251,N_7601,N_7715);
and U9252 (N_9252,N_7926,N_7848);
nand U9253 (N_9253,N_7668,N_7692);
nand U9254 (N_9254,N_8112,N_7961);
and U9255 (N_9255,N_8360,N_8344);
or U9256 (N_9256,N_7690,N_7654);
xnor U9257 (N_9257,N_7844,N_8518);
xnor U9258 (N_9258,N_7506,N_8455);
nor U9259 (N_9259,N_8539,N_7743);
and U9260 (N_9260,N_8538,N_8330);
or U9261 (N_9261,N_8001,N_8228);
nor U9262 (N_9262,N_7805,N_8073);
nor U9263 (N_9263,N_8051,N_8203);
nor U9264 (N_9264,N_7669,N_8014);
nor U9265 (N_9265,N_8657,N_7989);
nor U9266 (N_9266,N_8104,N_8610);
nand U9267 (N_9267,N_7747,N_8101);
and U9268 (N_9268,N_7509,N_8042);
nand U9269 (N_9269,N_7658,N_8527);
nor U9270 (N_9270,N_8420,N_7653);
or U9271 (N_9271,N_8510,N_7540);
xor U9272 (N_9272,N_8149,N_8031);
and U9273 (N_9273,N_7584,N_7570);
xnor U9274 (N_9274,N_8333,N_8139);
nand U9275 (N_9275,N_7591,N_7677);
or U9276 (N_9276,N_7675,N_8615);
xor U9277 (N_9277,N_8269,N_8277);
nand U9278 (N_9278,N_8686,N_8621);
and U9279 (N_9279,N_8375,N_7587);
and U9280 (N_9280,N_8342,N_8422);
xnor U9281 (N_9281,N_8290,N_7555);
and U9282 (N_9282,N_7614,N_7888);
xor U9283 (N_9283,N_7779,N_8409);
or U9284 (N_9284,N_8673,N_7745);
or U9285 (N_9285,N_8150,N_8608);
or U9286 (N_9286,N_7663,N_7681);
xor U9287 (N_9287,N_8057,N_7811);
xnor U9288 (N_9288,N_7583,N_8711);
and U9289 (N_9289,N_7542,N_7870);
nand U9290 (N_9290,N_8660,N_8165);
and U9291 (N_9291,N_8735,N_7867);
or U9292 (N_9292,N_8465,N_8213);
or U9293 (N_9293,N_8681,N_8067);
nor U9294 (N_9294,N_8292,N_8256);
and U9295 (N_9295,N_7835,N_8207);
xor U9296 (N_9296,N_8209,N_7551);
xor U9297 (N_9297,N_8249,N_8034);
and U9298 (N_9298,N_7865,N_7640);
or U9299 (N_9299,N_7531,N_8361);
xnor U9300 (N_9300,N_8653,N_7950);
nor U9301 (N_9301,N_7944,N_7759);
or U9302 (N_9302,N_8611,N_8245);
nor U9303 (N_9303,N_7631,N_7952);
or U9304 (N_9304,N_7664,N_8291);
nand U9305 (N_9305,N_7761,N_7686);
nand U9306 (N_9306,N_7794,N_8674);
and U9307 (N_9307,N_8050,N_8479);
or U9308 (N_9308,N_7880,N_8242);
nor U9309 (N_9309,N_7953,N_7973);
and U9310 (N_9310,N_8146,N_8152);
nor U9311 (N_9311,N_8418,N_7860);
nor U9312 (N_9312,N_8013,N_8563);
or U9313 (N_9313,N_8032,N_7519);
nor U9314 (N_9314,N_8503,N_8690);
or U9315 (N_9315,N_7595,N_8589);
nand U9316 (N_9316,N_8502,N_8028);
nor U9317 (N_9317,N_7949,N_8339);
and U9318 (N_9318,N_8222,N_8007);
xor U9319 (N_9319,N_8670,N_7824);
nor U9320 (N_9320,N_7925,N_8552);
xnor U9321 (N_9321,N_7641,N_7547);
and U9322 (N_9322,N_8198,N_8738);
and U9323 (N_9323,N_8457,N_7847);
nor U9324 (N_9324,N_8415,N_8173);
xor U9325 (N_9325,N_8182,N_7788);
nor U9326 (N_9326,N_8737,N_8534);
and U9327 (N_9327,N_8480,N_8087);
nor U9328 (N_9328,N_8000,N_7605);
or U9329 (N_9329,N_8281,N_8404);
and U9330 (N_9330,N_8568,N_8458);
and U9331 (N_9331,N_8487,N_7802);
nor U9332 (N_9332,N_7866,N_8564);
nor U9333 (N_9333,N_7645,N_7825);
xnor U9334 (N_9334,N_8287,N_8613);
nand U9335 (N_9335,N_8009,N_8515);
nor U9336 (N_9336,N_7695,N_8068);
nor U9337 (N_9337,N_8647,N_7619);
or U9338 (N_9338,N_8206,N_8746);
and U9339 (N_9339,N_8024,N_8056);
and U9340 (N_9340,N_8604,N_8386);
and U9341 (N_9341,N_8029,N_8298);
nor U9342 (N_9342,N_7561,N_8570);
xor U9343 (N_9343,N_7520,N_7904);
xnor U9344 (N_9344,N_8655,N_7514);
nor U9345 (N_9345,N_8519,N_8178);
nor U9346 (N_9346,N_8603,N_7651);
nor U9347 (N_9347,N_7500,N_8089);
nand U9348 (N_9348,N_7693,N_7594);
nor U9349 (N_9349,N_7666,N_8120);
nor U9350 (N_9350,N_7985,N_8478);
nor U9351 (N_9351,N_8584,N_7928);
nor U9352 (N_9352,N_7898,N_8451);
nand U9353 (N_9353,N_8395,N_8307);
or U9354 (N_9354,N_7507,N_8648);
or U9355 (N_9355,N_7864,N_8025);
nand U9356 (N_9356,N_8709,N_7783);
nand U9357 (N_9357,N_8351,N_8224);
nor U9358 (N_9358,N_7814,N_8268);
nand U9359 (N_9359,N_8081,N_7821);
xor U9360 (N_9360,N_7894,N_8325);
nand U9361 (N_9361,N_8017,N_7711);
nor U9362 (N_9362,N_8678,N_8704);
nor U9363 (N_9363,N_8211,N_7931);
nor U9364 (N_9364,N_8241,N_8097);
and U9365 (N_9365,N_8596,N_8331);
xnor U9366 (N_9366,N_7829,N_8373);
and U9367 (N_9367,N_8376,N_7633);
xor U9368 (N_9368,N_7921,N_8337);
nor U9369 (N_9369,N_8008,N_7683);
nand U9370 (N_9370,N_7740,N_8297);
nor U9371 (N_9371,N_8494,N_8747);
or U9372 (N_9372,N_7679,N_7800);
nor U9373 (N_9373,N_7970,N_7671);
xor U9374 (N_9374,N_7588,N_7820);
nand U9375 (N_9375,N_8705,N_8408);
xnor U9376 (N_9376,N_8439,N_7880);
and U9377 (N_9377,N_7711,N_8526);
nand U9378 (N_9378,N_7538,N_8455);
nor U9379 (N_9379,N_8051,N_8436);
nand U9380 (N_9380,N_7737,N_7727);
nand U9381 (N_9381,N_8662,N_8385);
and U9382 (N_9382,N_7991,N_8495);
and U9383 (N_9383,N_8214,N_8587);
and U9384 (N_9384,N_7875,N_8162);
nand U9385 (N_9385,N_7549,N_8541);
xnor U9386 (N_9386,N_7806,N_7549);
and U9387 (N_9387,N_7711,N_8734);
nand U9388 (N_9388,N_8448,N_8667);
xnor U9389 (N_9389,N_8341,N_7914);
and U9390 (N_9390,N_7767,N_7705);
or U9391 (N_9391,N_8103,N_7734);
xnor U9392 (N_9392,N_8365,N_8376);
or U9393 (N_9393,N_8238,N_7698);
and U9394 (N_9394,N_7667,N_8673);
and U9395 (N_9395,N_8375,N_8074);
nor U9396 (N_9396,N_8680,N_8295);
or U9397 (N_9397,N_7967,N_8318);
and U9398 (N_9398,N_8612,N_7879);
nand U9399 (N_9399,N_8601,N_7761);
or U9400 (N_9400,N_8113,N_8403);
or U9401 (N_9401,N_8672,N_8450);
nor U9402 (N_9402,N_8020,N_8384);
or U9403 (N_9403,N_7811,N_7610);
nor U9404 (N_9404,N_8475,N_7549);
nand U9405 (N_9405,N_8685,N_8274);
and U9406 (N_9406,N_8342,N_7825);
xnor U9407 (N_9407,N_7605,N_8601);
and U9408 (N_9408,N_8181,N_7551);
nand U9409 (N_9409,N_7799,N_8041);
and U9410 (N_9410,N_8324,N_7561);
nand U9411 (N_9411,N_8667,N_8632);
nor U9412 (N_9412,N_8454,N_8708);
nand U9413 (N_9413,N_8545,N_8594);
nor U9414 (N_9414,N_7522,N_8520);
nand U9415 (N_9415,N_7626,N_8184);
and U9416 (N_9416,N_7568,N_7526);
or U9417 (N_9417,N_7540,N_8213);
and U9418 (N_9418,N_7620,N_8055);
or U9419 (N_9419,N_8450,N_8137);
xnor U9420 (N_9420,N_7697,N_8616);
nand U9421 (N_9421,N_8527,N_7663);
nand U9422 (N_9422,N_8740,N_8434);
xor U9423 (N_9423,N_7515,N_7878);
xor U9424 (N_9424,N_8708,N_8106);
and U9425 (N_9425,N_8236,N_8591);
nand U9426 (N_9426,N_7926,N_7734);
nor U9427 (N_9427,N_8249,N_8251);
or U9428 (N_9428,N_8398,N_8630);
xor U9429 (N_9429,N_8197,N_8511);
nand U9430 (N_9430,N_8740,N_7867);
xor U9431 (N_9431,N_7791,N_8472);
xnor U9432 (N_9432,N_8483,N_8704);
and U9433 (N_9433,N_8323,N_7870);
nand U9434 (N_9434,N_7709,N_8192);
or U9435 (N_9435,N_8055,N_7701);
nand U9436 (N_9436,N_7622,N_7944);
xnor U9437 (N_9437,N_7955,N_8537);
xor U9438 (N_9438,N_8088,N_8542);
nand U9439 (N_9439,N_8134,N_8070);
nand U9440 (N_9440,N_8185,N_7737);
nand U9441 (N_9441,N_8004,N_8231);
or U9442 (N_9442,N_8193,N_8430);
nor U9443 (N_9443,N_8617,N_7804);
nand U9444 (N_9444,N_7586,N_8372);
nand U9445 (N_9445,N_8739,N_8032);
nor U9446 (N_9446,N_7866,N_8335);
nor U9447 (N_9447,N_7942,N_8010);
and U9448 (N_9448,N_7521,N_8016);
or U9449 (N_9449,N_8709,N_8438);
and U9450 (N_9450,N_8536,N_7667);
xnor U9451 (N_9451,N_8101,N_7623);
xnor U9452 (N_9452,N_8302,N_7632);
nor U9453 (N_9453,N_7702,N_8619);
xor U9454 (N_9454,N_8391,N_7894);
or U9455 (N_9455,N_8207,N_8702);
and U9456 (N_9456,N_8715,N_8352);
nor U9457 (N_9457,N_7702,N_7817);
xor U9458 (N_9458,N_7993,N_7798);
and U9459 (N_9459,N_8343,N_8703);
nand U9460 (N_9460,N_8610,N_8408);
nand U9461 (N_9461,N_8281,N_7569);
nor U9462 (N_9462,N_8506,N_8130);
and U9463 (N_9463,N_7963,N_7673);
xor U9464 (N_9464,N_7843,N_8633);
nor U9465 (N_9465,N_8725,N_7686);
nor U9466 (N_9466,N_7808,N_8193);
and U9467 (N_9467,N_7640,N_7851);
or U9468 (N_9468,N_8576,N_7505);
xnor U9469 (N_9469,N_8444,N_8607);
and U9470 (N_9470,N_8710,N_8050);
and U9471 (N_9471,N_7593,N_8542);
or U9472 (N_9472,N_8581,N_8743);
nor U9473 (N_9473,N_8298,N_8377);
xor U9474 (N_9474,N_8170,N_7723);
xor U9475 (N_9475,N_8389,N_7890);
or U9476 (N_9476,N_7535,N_8566);
and U9477 (N_9477,N_8152,N_8657);
nor U9478 (N_9478,N_8057,N_7747);
xor U9479 (N_9479,N_8484,N_8532);
nand U9480 (N_9480,N_8592,N_8019);
nand U9481 (N_9481,N_7515,N_7843);
or U9482 (N_9482,N_8019,N_7813);
or U9483 (N_9483,N_8215,N_8350);
and U9484 (N_9484,N_8563,N_7626);
nor U9485 (N_9485,N_8286,N_8509);
nor U9486 (N_9486,N_8678,N_8467);
xnor U9487 (N_9487,N_8485,N_7683);
nand U9488 (N_9488,N_8537,N_7857);
nand U9489 (N_9489,N_7662,N_8504);
xnor U9490 (N_9490,N_7644,N_8222);
nor U9491 (N_9491,N_7999,N_8279);
and U9492 (N_9492,N_7667,N_8459);
xor U9493 (N_9493,N_8364,N_8497);
nand U9494 (N_9494,N_8313,N_8607);
and U9495 (N_9495,N_7662,N_8066);
xor U9496 (N_9496,N_8416,N_7685);
and U9497 (N_9497,N_7649,N_8335);
nor U9498 (N_9498,N_8113,N_8034);
nor U9499 (N_9499,N_7824,N_8099);
xnor U9500 (N_9500,N_7850,N_8324);
xor U9501 (N_9501,N_8393,N_8731);
nor U9502 (N_9502,N_7855,N_8564);
or U9503 (N_9503,N_8241,N_8053);
nor U9504 (N_9504,N_7535,N_8625);
nor U9505 (N_9505,N_8412,N_8738);
xor U9506 (N_9506,N_8686,N_8038);
and U9507 (N_9507,N_7582,N_7882);
and U9508 (N_9508,N_8389,N_8748);
or U9509 (N_9509,N_7528,N_7922);
or U9510 (N_9510,N_7813,N_8673);
nand U9511 (N_9511,N_8594,N_7921);
nor U9512 (N_9512,N_7569,N_8722);
or U9513 (N_9513,N_8393,N_8360);
and U9514 (N_9514,N_8026,N_8731);
and U9515 (N_9515,N_8109,N_7805);
nor U9516 (N_9516,N_8130,N_8275);
and U9517 (N_9517,N_8722,N_8376);
and U9518 (N_9518,N_8287,N_8655);
nand U9519 (N_9519,N_8331,N_8098);
or U9520 (N_9520,N_7656,N_7660);
nor U9521 (N_9521,N_7740,N_8004);
or U9522 (N_9522,N_8474,N_7550);
xnor U9523 (N_9523,N_8470,N_8650);
nor U9524 (N_9524,N_8142,N_8286);
nand U9525 (N_9525,N_8086,N_7878);
nor U9526 (N_9526,N_8066,N_8163);
nor U9527 (N_9527,N_7723,N_8555);
and U9528 (N_9528,N_8280,N_7683);
nand U9529 (N_9529,N_7634,N_7937);
and U9530 (N_9530,N_8618,N_8032);
nor U9531 (N_9531,N_7811,N_8151);
xnor U9532 (N_9532,N_7568,N_8167);
or U9533 (N_9533,N_8448,N_8491);
and U9534 (N_9534,N_8103,N_8664);
nor U9535 (N_9535,N_8084,N_7601);
or U9536 (N_9536,N_7921,N_7727);
or U9537 (N_9537,N_7617,N_8489);
nor U9538 (N_9538,N_7592,N_8306);
nand U9539 (N_9539,N_8061,N_8570);
or U9540 (N_9540,N_8608,N_7733);
nand U9541 (N_9541,N_8432,N_8371);
nor U9542 (N_9542,N_7795,N_8065);
nor U9543 (N_9543,N_8659,N_7501);
nor U9544 (N_9544,N_8680,N_8235);
xnor U9545 (N_9545,N_8319,N_8692);
and U9546 (N_9546,N_8357,N_8500);
and U9547 (N_9547,N_8328,N_8214);
and U9548 (N_9548,N_8625,N_8282);
nor U9549 (N_9549,N_7659,N_7639);
nor U9550 (N_9550,N_8502,N_7791);
nor U9551 (N_9551,N_8020,N_8576);
nand U9552 (N_9552,N_8420,N_8166);
and U9553 (N_9553,N_8588,N_8519);
and U9554 (N_9554,N_7777,N_8178);
or U9555 (N_9555,N_7664,N_7746);
and U9556 (N_9556,N_8296,N_8294);
and U9557 (N_9557,N_8560,N_7633);
nand U9558 (N_9558,N_8231,N_7686);
nand U9559 (N_9559,N_7590,N_7961);
nor U9560 (N_9560,N_8597,N_8633);
and U9561 (N_9561,N_7680,N_8006);
nand U9562 (N_9562,N_7644,N_8416);
xor U9563 (N_9563,N_7772,N_7605);
or U9564 (N_9564,N_8441,N_8301);
or U9565 (N_9565,N_8304,N_7645);
or U9566 (N_9566,N_7779,N_8450);
nand U9567 (N_9567,N_8353,N_8675);
nor U9568 (N_9568,N_7610,N_7715);
xor U9569 (N_9569,N_8087,N_8644);
nor U9570 (N_9570,N_7614,N_7931);
and U9571 (N_9571,N_8438,N_8502);
and U9572 (N_9572,N_8196,N_7932);
nand U9573 (N_9573,N_7639,N_8399);
xnor U9574 (N_9574,N_7604,N_8096);
nand U9575 (N_9575,N_8667,N_8050);
or U9576 (N_9576,N_7743,N_7915);
nor U9577 (N_9577,N_8636,N_7712);
nor U9578 (N_9578,N_7638,N_8594);
and U9579 (N_9579,N_8481,N_8180);
nand U9580 (N_9580,N_7639,N_7847);
xnor U9581 (N_9581,N_8391,N_8622);
nor U9582 (N_9582,N_8397,N_8253);
and U9583 (N_9583,N_7823,N_8187);
nor U9584 (N_9584,N_7536,N_8326);
xor U9585 (N_9585,N_7782,N_7812);
nand U9586 (N_9586,N_8565,N_8719);
nor U9587 (N_9587,N_7608,N_8441);
or U9588 (N_9588,N_8249,N_7879);
and U9589 (N_9589,N_7900,N_8442);
and U9590 (N_9590,N_7720,N_8206);
xor U9591 (N_9591,N_8100,N_8339);
nor U9592 (N_9592,N_8116,N_8345);
and U9593 (N_9593,N_8432,N_7776);
nor U9594 (N_9594,N_8505,N_7567);
xnor U9595 (N_9595,N_8380,N_8478);
nor U9596 (N_9596,N_8390,N_8733);
nand U9597 (N_9597,N_7841,N_8577);
xnor U9598 (N_9598,N_7769,N_7838);
nor U9599 (N_9599,N_8416,N_8593);
nor U9600 (N_9600,N_8317,N_8328);
nor U9601 (N_9601,N_7748,N_8001);
nand U9602 (N_9602,N_8324,N_7790);
xor U9603 (N_9603,N_8076,N_7559);
or U9604 (N_9604,N_7696,N_7542);
nand U9605 (N_9605,N_8622,N_8019);
and U9606 (N_9606,N_7693,N_7915);
xor U9607 (N_9607,N_8021,N_8332);
nor U9608 (N_9608,N_8514,N_8478);
nor U9609 (N_9609,N_8633,N_7535);
nor U9610 (N_9610,N_8683,N_8425);
and U9611 (N_9611,N_7511,N_7880);
and U9612 (N_9612,N_8276,N_8154);
nand U9613 (N_9613,N_8299,N_8538);
nand U9614 (N_9614,N_8408,N_8655);
nor U9615 (N_9615,N_8081,N_8311);
nand U9616 (N_9616,N_7612,N_7962);
xnor U9617 (N_9617,N_7686,N_8613);
nand U9618 (N_9618,N_8125,N_7755);
or U9619 (N_9619,N_8599,N_7807);
and U9620 (N_9620,N_8006,N_8514);
or U9621 (N_9621,N_8488,N_8106);
or U9622 (N_9622,N_7634,N_7521);
nor U9623 (N_9623,N_7757,N_8049);
xnor U9624 (N_9624,N_8691,N_8711);
nor U9625 (N_9625,N_8138,N_7981);
or U9626 (N_9626,N_7957,N_8404);
nor U9627 (N_9627,N_8382,N_8169);
nor U9628 (N_9628,N_7518,N_8669);
and U9629 (N_9629,N_8223,N_8740);
and U9630 (N_9630,N_8171,N_7840);
or U9631 (N_9631,N_8508,N_8194);
or U9632 (N_9632,N_8092,N_7604);
nand U9633 (N_9633,N_8549,N_8187);
nand U9634 (N_9634,N_8643,N_8276);
nand U9635 (N_9635,N_7956,N_8481);
and U9636 (N_9636,N_8163,N_7659);
nand U9637 (N_9637,N_8183,N_8749);
and U9638 (N_9638,N_8418,N_7793);
or U9639 (N_9639,N_8126,N_8355);
nand U9640 (N_9640,N_8698,N_7788);
xor U9641 (N_9641,N_7870,N_7722);
or U9642 (N_9642,N_8298,N_7961);
xor U9643 (N_9643,N_7995,N_7707);
xnor U9644 (N_9644,N_7945,N_7856);
nand U9645 (N_9645,N_8542,N_8529);
nor U9646 (N_9646,N_8247,N_7537);
nand U9647 (N_9647,N_7503,N_7623);
nor U9648 (N_9648,N_7507,N_7629);
nand U9649 (N_9649,N_8132,N_7822);
nand U9650 (N_9650,N_7638,N_7539);
or U9651 (N_9651,N_8516,N_7522);
nand U9652 (N_9652,N_8306,N_8211);
or U9653 (N_9653,N_7990,N_8356);
or U9654 (N_9654,N_7503,N_8665);
nand U9655 (N_9655,N_8702,N_8626);
xor U9656 (N_9656,N_7791,N_8666);
and U9657 (N_9657,N_8493,N_7749);
xor U9658 (N_9658,N_8610,N_8022);
nor U9659 (N_9659,N_8384,N_8340);
xor U9660 (N_9660,N_7698,N_7741);
xor U9661 (N_9661,N_8283,N_8528);
or U9662 (N_9662,N_8196,N_8259);
xor U9663 (N_9663,N_7778,N_8741);
or U9664 (N_9664,N_7541,N_8653);
and U9665 (N_9665,N_8243,N_8022);
xor U9666 (N_9666,N_8630,N_7864);
xnor U9667 (N_9667,N_7923,N_8468);
and U9668 (N_9668,N_8306,N_7755);
nand U9669 (N_9669,N_7944,N_8442);
nor U9670 (N_9670,N_8030,N_7892);
nand U9671 (N_9671,N_8670,N_7804);
xor U9672 (N_9672,N_7972,N_8166);
nor U9673 (N_9673,N_8632,N_7817);
nand U9674 (N_9674,N_8042,N_7712);
nor U9675 (N_9675,N_8675,N_8570);
nor U9676 (N_9676,N_8576,N_8701);
nor U9677 (N_9677,N_7819,N_8455);
or U9678 (N_9678,N_7761,N_7964);
xnor U9679 (N_9679,N_8445,N_8701);
and U9680 (N_9680,N_8248,N_8178);
and U9681 (N_9681,N_8386,N_7814);
xor U9682 (N_9682,N_7680,N_8663);
xor U9683 (N_9683,N_7939,N_8124);
or U9684 (N_9684,N_8009,N_8098);
nor U9685 (N_9685,N_8330,N_7702);
or U9686 (N_9686,N_8123,N_8448);
and U9687 (N_9687,N_7604,N_8383);
or U9688 (N_9688,N_8539,N_8178);
or U9689 (N_9689,N_8243,N_7827);
and U9690 (N_9690,N_8064,N_8095);
xnor U9691 (N_9691,N_8541,N_7877);
nand U9692 (N_9692,N_7845,N_8626);
nand U9693 (N_9693,N_8651,N_8649);
or U9694 (N_9694,N_7640,N_7933);
and U9695 (N_9695,N_7760,N_8490);
xnor U9696 (N_9696,N_7751,N_8574);
or U9697 (N_9697,N_8011,N_8624);
and U9698 (N_9698,N_8139,N_8602);
or U9699 (N_9699,N_8211,N_8030);
or U9700 (N_9700,N_8386,N_7530);
or U9701 (N_9701,N_8643,N_8287);
nand U9702 (N_9702,N_8698,N_7534);
and U9703 (N_9703,N_8465,N_8460);
nor U9704 (N_9704,N_8326,N_8290);
nor U9705 (N_9705,N_8283,N_8229);
or U9706 (N_9706,N_7910,N_7930);
nand U9707 (N_9707,N_8459,N_8051);
nor U9708 (N_9708,N_8289,N_8296);
and U9709 (N_9709,N_7742,N_8618);
or U9710 (N_9710,N_8415,N_7748);
or U9711 (N_9711,N_8091,N_8040);
nand U9712 (N_9712,N_7573,N_7839);
xor U9713 (N_9713,N_8507,N_7686);
xnor U9714 (N_9714,N_7931,N_7529);
and U9715 (N_9715,N_8497,N_8653);
nand U9716 (N_9716,N_7532,N_8673);
or U9717 (N_9717,N_8295,N_8711);
xnor U9718 (N_9718,N_8735,N_8162);
xnor U9719 (N_9719,N_8483,N_7570);
nand U9720 (N_9720,N_7980,N_7836);
nand U9721 (N_9721,N_8405,N_8518);
nand U9722 (N_9722,N_8166,N_8037);
or U9723 (N_9723,N_7988,N_8058);
nor U9724 (N_9724,N_8426,N_8746);
xor U9725 (N_9725,N_8538,N_8434);
xnor U9726 (N_9726,N_7687,N_8620);
or U9727 (N_9727,N_8026,N_7641);
nand U9728 (N_9728,N_8712,N_8233);
xnor U9729 (N_9729,N_8132,N_7998);
and U9730 (N_9730,N_8147,N_8487);
xor U9731 (N_9731,N_8477,N_8660);
nor U9732 (N_9732,N_7967,N_8182);
nor U9733 (N_9733,N_7544,N_8381);
xor U9734 (N_9734,N_8701,N_8053);
nor U9735 (N_9735,N_8292,N_8240);
or U9736 (N_9736,N_7850,N_8554);
or U9737 (N_9737,N_8295,N_8460);
nand U9738 (N_9738,N_8145,N_8197);
xor U9739 (N_9739,N_8419,N_8454);
nand U9740 (N_9740,N_8358,N_7884);
or U9741 (N_9741,N_8065,N_7599);
or U9742 (N_9742,N_8738,N_8709);
nor U9743 (N_9743,N_7802,N_8414);
nor U9744 (N_9744,N_8335,N_8657);
and U9745 (N_9745,N_7675,N_8399);
nand U9746 (N_9746,N_7942,N_8258);
xnor U9747 (N_9747,N_8480,N_8703);
nor U9748 (N_9748,N_7514,N_8371);
nand U9749 (N_9749,N_8540,N_7700);
or U9750 (N_9750,N_7640,N_7710);
and U9751 (N_9751,N_8154,N_8142);
xnor U9752 (N_9752,N_7587,N_8312);
nand U9753 (N_9753,N_7730,N_7778);
xnor U9754 (N_9754,N_8061,N_7826);
nor U9755 (N_9755,N_7737,N_8086);
xor U9756 (N_9756,N_8569,N_7689);
or U9757 (N_9757,N_7919,N_8043);
xor U9758 (N_9758,N_7532,N_8131);
xnor U9759 (N_9759,N_7505,N_8065);
nand U9760 (N_9760,N_8141,N_7889);
nand U9761 (N_9761,N_8745,N_7712);
and U9762 (N_9762,N_8449,N_7641);
nand U9763 (N_9763,N_8164,N_8251);
or U9764 (N_9764,N_8226,N_7501);
and U9765 (N_9765,N_8345,N_8026);
xor U9766 (N_9766,N_8198,N_7741);
nand U9767 (N_9767,N_7635,N_8488);
xor U9768 (N_9768,N_8491,N_8167);
and U9769 (N_9769,N_8351,N_8173);
xnor U9770 (N_9770,N_7527,N_8717);
and U9771 (N_9771,N_7681,N_7807);
nand U9772 (N_9772,N_8503,N_8235);
xnor U9773 (N_9773,N_7616,N_8572);
and U9774 (N_9774,N_8012,N_8494);
nand U9775 (N_9775,N_7642,N_7530);
nor U9776 (N_9776,N_8095,N_7595);
and U9777 (N_9777,N_8565,N_7692);
nor U9778 (N_9778,N_7715,N_8658);
nand U9779 (N_9779,N_7861,N_8183);
or U9780 (N_9780,N_8728,N_7834);
or U9781 (N_9781,N_8006,N_7773);
nand U9782 (N_9782,N_7802,N_7846);
or U9783 (N_9783,N_7886,N_8524);
or U9784 (N_9784,N_7562,N_7755);
nand U9785 (N_9785,N_8626,N_8022);
nor U9786 (N_9786,N_7591,N_8069);
xnor U9787 (N_9787,N_7951,N_7857);
nor U9788 (N_9788,N_7538,N_7553);
or U9789 (N_9789,N_8747,N_8505);
xnor U9790 (N_9790,N_7801,N_7753);
nor U9791 (N_9791,N_8307,N_7810);
nand U9792 (N_9792,N_8164,N_7501);
and U9793 (N_9793,N_8179,N_8130);
nor U9794 (N_9794,N_8263,N_8135);
or U9795 (N_9795,N_7868,N_8708);
nand U9796 (N_9796,N_8006,N_8181);
nand U9797 (N_9797,N_8361,N_8327);
nand U9798 (N_9798,N_8682,N_8430);
xnor U9799 (N_9799,N_7611,N_7672);
xnor U9800 (N_9800,N_8739,N_8402);
nor U9801 (N_9801,N_8446,N_7773);
xnor U9802 (N_9802,N_8626,N_8602);
and U9803 (N_9803,N_7945,N_7770);
xor U9804 (N_9804,N_7881,N_7918);
xnor U9805 (N_9805,N_8059,N_8614);
and U9806 (N_9806,N_8047,N_8248);
nand U9807 (N_9807,N_8059,N_7717);
nor U9808 (N_9808,N_8720,N_7952);
and U9809 (N_9809,N_8092,N_8263);
nor U9810 (N_9810,N_8345,N_7585);
or U9811 (N_9811,N_8583,N_8163);
xor U9812 (N_9812,N_7903,N_7592);
nand U9813 (N_9813,N_7951,N_8237);
xor U9814 (N_9814,N_8647,N_8033);
and U9815 (N_9815,N_7919,N_8356);
nand U9816 (N_9816,N_7998,N_7962);
nor U9817 (N_9817,N_8572,N_8358);
nand U9818 (N_9818,N_8552,N_8325);
and U9819 (N_9819,N_8447,N_7712);
nand U9820 (N_9820,N_8577,N_8451);
and U9821 (N_9821,N_7666,N_7856);
nor U9822 (N_9822,N_8717,N_7662);
xor U9823 (N_9823,N_7537,N_7958);
xnor U9824 (N_9824,N_8296,N_7732);
nand U9825 (N_9825,N_8124,N_8250);
nor U9826 (N_9826,N_8389,N_8007);
nand U9827 (N_9827,N_7674,N_8587);
or U9828 (N_9828,N_8150,N_8107);
xnor U9829 (N_9829,N_7999,N_8040);
nor U9830 (N_9830,N_7741,N_7630);
xor U9831 (N_9831,N_8267,N_8297);
nor U9832 (N_9832,N_8493,N_8695);
or U9833 (N_9833,N_8076,N_8606);
and U9834 (N_9834,N_7606,N_8226);
nor U9835 (N_9835,N_8401,N_8671);
or U9836 (N_9836,N_7565,N_7846);
xor U9837 (N_9837,N_8698,N_8713);
xnor U9838 (N_9838,N_8721,N_7830);
xor U9839 (N_9839,N_8446,N_8726);
or U9840 (N_9840,N_8598,N_8236);
and U9841 (N_9841,N_8588,N_8359);
nor U9842 (N_9842,N_8538,N_8476);
nand U9843 (N_9843,N_7684,N_8201);
or U9844 (N_9844,N_8474,N_8226);
or U9845 (N_9845,N_7628,N_8051);
nand U9846 (N_9846,N_8219,N_7665);
nand U9847 (N_9847,N_8672,N_7949);
nand U9848 (N_9848,N_8607,N_8089);
xor U9849 (N_9849,N_7560,N_7867);
or U9850 (N_9850,N_7508,N_8196);
and U9851 (N_9851,N_8694,N_7715);
nor U9852 (N_9852,N_8018,N_8008);
nor U9853 (N_9853,N_8524,N_7646);
xnor U9854 (N_9854,N_8004,N_8709);
xnor U9855 (N_9855,N_8255,N_8457);
or U9856 (N_9856,N_7808,N_8027);
nand U9857 (N_9857,N_8308,N_7735);
and U9858 (N_9858,N_7527,N_8159);
nor U9859 (N_9859,N_8054,N_8296);
xnor U9860 (N_9860,N_7719,N_7916);
nor U9861 (N_9861,N_7929,N_7745);
xor U9862 (N_9862,N_8547,N_8224);
and U9863 (N_9863,N_8357,N_8235);
nor U9864 (N_9864,N_7782,N_8445);
nor U9865 (N_9865,N_7880,N_8180);
nor U9866 (N_9866,N_7871,N_7820);
and U9867 (N_9867,N_7588,N_8117);
nor U9868 (N_9868,N_8038,N_7743);
xnor U9869 (N_9869,N_8480,N_7515);
nor U9870 (N_9870,N_8632,N_8507);
or U9871 (N_9871,N_7536,N_8560);
or U9872 (N_9872,N_8672,N_8001);
nor U9873 (N_9873,N_7986,N_8236);
xor U9874 (N_9874,N_7857,N_8527);
or U9875 (N_9875,N_7820,N_8502);
nand U9876 (N_9876,N_8279,N_8022);
nand U9877 (N_9877,N_8286,N_7828);
or U9878 (N_9878,N_8206,N_8532);
and U9879 (N_9879,N_8442,N_7659);
nand U9880 (N_9880,N_7520,N_7856);
and U9881 (N_9881,N_7946,N_8114);
nand U9882 (N_9882,N_8386,N_8533);
nor U9883 (N_9883,N_7735,N_7725);
nor U9884 (N_9884,N_8745,N_7689);
nor U9885 (N_9885,N_8704,N_7722);
nor U9886 (N_9886,N_7960,N_8411);
or U9887 (N_9887,N_7906,N_8645);
and U9888 (N_9888,N_7910,N_8509);
and U9889 (N_9889,N_7930,N_8135);
nand U9890 (N_9890,N_8535,N_8126);
xor U9891 (N_9891,N_8042,N_7555);
xnor U9892 (N_9892,N_7786,N_7879);
xnor U9893 (N_9893,N_8723,N_8560);
or U9894 (N_9894,N_7688,N_7622);
nand U9895 (N_9895,N_8418,N_8340);
and U9896 (N_9896,N_8606,N_7840);
nand U9897 (N_9897,N_7594,N_7624);
and U9898 (N_9898,N_7822,N_8059);
nand U9899 (N_9899,N_7741,N_8126);
and U9900 (N_9900,N_7723,N_8653);
or U9901 (N_9901,N_8369,N_8480);
nand U9902 (N_9902,N_8350,N_8695);
and U9903 (N_9903,N_8384,N_8244);
xnor U9904 (N_9904,N_8487,N_7993);
nand U9905 (N_9905,N_7727,N_8446);
nor U9906 (N_9906,N_7771,N_8196);
nand U9907 (N_9907,N_8720,N_8516);
or U9908 (N_9908,N_7530,N_8467);
nor U9909 (N_9909,N_7697,N_8068);
and U9910 (N_9910,N_8503,N_7822);
nand U9911 (N_9911,N_8438,N_8733);
nand U9912 (N_9912,N_8570,N_8272);
and U9913 (N_9913,N_8276,N_8689);
xor U9914 (N_9914,N_7670,N_7991);
xor U9915 (N_9915,N_8239,N_8019);
nor U9916 (N_9916,N_8638,N_8660);
nand U9917 (N_9917,N_7528,N_8728);
xor U9918 (N_9918,N_8264,N_8135);
nor U9919 (N_9919,N_8063,N_7937);
nand U9920 (N_9920,N_8607,N_7554);
and U9921 (N_9921,N_8501,N_8585);
and U9922 (N_9922,N_7720,N_8208);
or U9923 (N_9923,N_7616,N_7573);
or U9924 (N_9924,N_8407,N_8125);
and U9925 (N_9925,N_7752,N_8309);
and U9926 (N_9926,N_7984,N_7590);
xnor U9927 (N_9927,N_7738,N_7894);
nand U9928 (N_9928,N_8588,N_7500);
and U9929 (N_9929,N_8126,N_7543);
xnor U9930 (N_9930,N_8533,N_8501);
xor U9931 (N_9931,N_7511,N_8605);
and U9932 (N_9932,N_8295,N_8496);
nand U9933 (N_9933,N_8154,N_8592);
and U9934 (N_9934,N_8243,N_8528);
xor U9935 (N_9935,N_7552,N_8735);
xor U9936 (N_9936,N_8732,N_7650);
and U9937 (N_9937,N_8505,N_7507);
xor U9938 (N_9938,N_8034,N_8693);
and U9939 (N_9939,N_7920,N_8711);
nand U9940 (N_9940,N_8481,N_7715);
xnor U9941 (N_9941,N_8231,N_7969);
nand U9942 (N_9942,N_8263,N_8238);
xor U9943 (N_9943,N_7529,N_8628);
and U9944 (N_9944,N_8733,N_8280);
or U9945 (N_9945,N_8713,N_8512);
nor U9946 (N_9946,N_7686,N_7671);
nor U9947 (N_9947,N_8262,N_8065);
nand U9948 (N_9948,N_8434,N_7587);
xnor U9949 (N_9949,N_8329,N_7696);
and U9950 (N_9950,N_8043,N_8308);
or U9951 (N_9951,N_8742,N_8113);
xnor U9952 (N_9952,N_8049,N_7801);
xor U9953 (N_9953,N_8081,N_8475);
nor U9954 (N_9954,N_8481,N_7735);
xnor U9955 (N_9955,N_7891,N_7632);
xor U9956 (N_9956,N_7589,N_8129);
and U9957 (N_9957,N_8696,N_8694);
xnor U9958 (N_9958,N_8723,N_7632);
and U9959 (N_9959,N_7940,N_7998);
or U9960 (N_9960,N_8484,N_7570);
nand U9961 (N_9961,N_8115,N_7727);
and U9962 (N_9962,N_8220,N_8583);
or U9963 (N_9963,N_7646,N_7878);
nor U9964 (N_9964,N_8180,N_8570);
or U9965 (N_9965,N_7809,N_7913);
or U9966 (N_9966,N_8032,N_8315);
nand U9967 (N_9967,N_8411,N_8700);
and U9968 (N_9968,N_8704,N_7831);
xnor U9969 (N_9969,N_7517,N_7739);
or U9970 (N_9970,N_7557,N_7602);
and U9971 (N_9971,N_7642,N_8748);
nand U9972 (N_9972,N_7765,N_7971);
and U9973 (N_9973,N_8156,N_7990);
nor U9974 (N_9974,N_8501,N_8295);
xor U9975 (N_9975,N_7927,N_8015);
or U9976 (N_9976,N_7555,N_8457);
or U9977 (N_9977,N_8419,N_7935);
nand U9978 (N_9978,N_8249,N_8044);
or U9979 (N_9979,N_7843,N_7644);
or U9980 (N_9980,N_7714,N_8347);
and U9981 (N_9981,N_8676,N_7564);
xnor U9982 (N_9982,N_8677,N_7881);
and U9983 (N_9983,N_7756,N_7886);
and U9984 (N_9984,N_8253,N_7635);
nor U9985 (N_9985,N_7903,N_8085);
and U9986 (N_9986,N_7596,N_7661);
xnor U9987 (N_9987,N_8584,N_8592);
and U9988 (N_9988,N_8116,N_8633);
nor U9989 (N_9989,N_7974,N_7965);
nand U9990 (N_9990,N_8002,N_8684);
nor U9991 (N_9991,N_7602,N_8735);
nor U9992 (N_9992,N_7747,N_8078);
xor U9993 (N_9993,N_7993,N_7727);
xnor U9994 (N_9994,N_8182,N_7806);
xnor U9995 (N_9995,N_8502,N_8253);
or U9996 (N_9996,N_8479,N_8565);
or U9997 (N_9997,N_8316,N_7652);
and U9998 (N_9998,N_8527,N_7807);
nand U9999 (N_9999,N_7550,N_8379);
and U10000 (N_10000,N_9880,N_9565);
or U10001 (N_10001,N_9155,N_9649);
xnor U10002 (N_10002,N_9911,N_8818);
nand U10003 (N_10003,N_9326,N_9685);
nand U10004 (N_10004,N_9756,N_9855);
xor U10005 (N_10005,N_9696,N_9031);
nand U10006 (N_10006,N_9280,N_8875);
nand U10007 (N_10007,N_9513,N_9820);
nor U10008 (N_10008,N_9997,N_8861);
nor U10009 (N_10009,N_9913,N_9842);
or U10010 (N_10010,N_9009,N_9865);
and U10011 (N_10011,N_8864,N_9066);
xor U10012 (N_10012,N_9924,N_8844);
nand U10013 (N_10013,N_9753,N_8838);
nand U10014 (N_10014,N_9844,N_9364);
or U10015 (N_10015,N_8958,N_9255);
nor U10016 (N_10016,N_9692,N_9204);
and U10017 (N_10017,N_9959,N_9626);
or U10018 (N_10018,N_9270,N_9431);
or U10019 (N_10019,N_8840,N_9025);
nand U10020 (N_10020,N_9430,N_9616);
or U10021 (N_10021,N_8904,N_9879);
and U10022 (N_10022,N_8901,N_9787);
and U10023 (N_10023,N_9514,N_9015);
nand U10024 (N_10024,N_9713,N_9619);
xnor U10025 (N_10025,N_8899,N_9758);
or U10026 (N_10026,N_9931,N_9214);
nand U10027 (N_10027,N_9044,N_9733);
nand U10028 (N_10028,N_9955,N_9331);
nand U10029 (N_10029,N_9599,N_9540);
xnor U10030 (N_10030,N_9223,N_9112);
nor U10031 (N_10031,N_9466,N_9989);
or U10032 (N_10032,N_8862,N_8800);
nand U10033 (N_10033,N_9013,N_9121);
xor U10034 (N_10034,N_9423,N_9827);
and U10035 (N_10035,N_8791,N_8996);
nor U10036 (N_10036,N_9886,N_8824);
and U10037 (N_10037,N_9515,N_9607);
or U10038 (N_10038,N_8999,N_9688);
xor U10039 (N_10039,N_9935,N_9137);
xor U10040 (N_10040,N_9057,N_9504);
or U10041 (N_10041,N_9114,N_9406);
or U10042 (N_10042,N_8902,N_9287);
nand U10043 (N_10043,N_9097,N_9100);
or U10044 (N_10044,N_9077,N_9983);
or U10045 (N_10045,N_8868,N_9461);
nand U10046 (N_10046,N_9645,N_8892);
and U10047 (N_10047,N_9725,N_9408);
nand U10048 (N_10048,N_9995,N_8889);
nor U10049 (N_10049,N_8764,N_9054);
and U10050 (N_10050,N_9166,N_8780);
xor U10051 (N_10051,N_9135,N_9470);
or U10052 (N_10052,N_8926,N_9857);
or U10053 (N_10053,N_8903,N_8927);
or U10054 (N_10054,N_9948,N_9048);
and U10055 (N_10055,N_9267,N_9977);
or U10056 (N_10056,N_9835,N_8989);
xor U10057 (N_10057,N_9803,N_9847);
xnor U10058 (N_10058,N_9336,N_9691);
and U10059 (N_10059,N_9106,N_9199);
nor U10060 (N_10060,N_8888,N_8956);
nor U10061 (N_10061,N_9561,N_8964);
and U10062 (N_10062,N_8783,N_9239);
xnor U10063 (N_10063,N_9081,N_9960);
xor U10064 (N_10064,N_9392,N_9578);
xnor U10065 (N_10065,N_9181,N_9316);
and U10066 (N_10066,N_9770,N_9129);
and U10067 (N_10067,N_9714,N_9990);
or U10068 (N_10068,N_9544,N_9123);
nand U10069 (N_10069,N_9251,N_9058);
xnor U10070 (N_10070,N_8912,N_9550);
nor U10071 (N_10071,N_9889,N_9850);
nor U10072 (N_10072,N_9912,N_8962);
or U10073 (N_10073,N_9853,N_8874);
nand U10074 (N_10074,N_9689,N_9420);
nand U10075 (N_10075,N_9200,N_9528);
or U10076 (N_10076,N_9205,N_9160);
nor U10077 (N_10077,N_8819,N_9186);
nor U10078 (N_10078,N_9901,N_9868);
nand U10079 (N_10079,N_8831,N_9278);
xor U10080 (N_10080,N_9676,N_9010);
xnor U10081 (N_10081,N_8925,N_9450);
or U10082 (N_10082,N_9973,N_9875);
or U10083 (N_10083,N_9001,N_9614);
xor U10084 (N_10084,N_9076,N_8804);
and U10085 (N_10085,N_8810,N_9162);
and U10086 (N_10086,N_9272,N_8916);
and U10087 (N_10087,N_9905,N_9424);
nor U10088 (N_10088,N_9652,N_8836);
nor U10089 (N_10089,N_8794,N_9116);
and U10090 (N_10090,N_9334,N_9472);
or U10091 (N_10091,N_9932,N_8805);
nand U10092 (N_10092,N_9441,N_9506);
nand U10093 (N_10093,N_9385,N_8871);
or U10094 (N_10094,N_9344,N_9915);
nor U10095 (N_10095,N_9498,N_9546);
nor U10096 (N_10096,N_8755,N_9130);
nand U10097 (N_10097,N_9635,N_9415);
and U10098 (N_10098,N_8858,N_9740);
or U10099 (N_10099,N_8975,N_8760);
nor U10100 (N_10100,N_9159,N_8809);
or U10101 (N_10101,N_9775,N_9683);
and U10102 (N_10102,N_8779,N_9501);
and U10103 (N_10103,N_9542,N_9548);
and U10104 (N_10104,N_9341,N_9361);
nor U10105 (N_10105,N_9474,N_9521);
and U10106 (N_10106,N_9084,N_9378);
xor U10107 (N_10107,N_9185,N_9560);
nand U10108 (N_10108,N_9360,N_9197);
nor U10109 (N_10109,N_8895,N_8795);
nor U10110 (N_10110,N_9678,N_8837);
and U10111 (N_10111,N_8821,N_8785);
xor U10112 (N_10112,N_9495,N_9212);
nor U10113 (N_10113,N_8984,N_8773);
and U10114 (N_10114,N_8827,N_9016);
nand U10115 (N_10115,N_9559,N_9772);
nand U10116 (N_10116,N_8812,N_9532);
nand U10117 (N_10117,N_8883,N_9227);
or U10118 (N_10118,N_8993,N_9545);
or U10119 (N_10119,N_9762,N_9936);
or U10120 (N_10120,N_9050,N_9790);
xnor U10121 (N_10121,N_9749,N_9873);
nand U10122 (N_10122,N_9864,N_9310);
nand U10123 (N_10123,N_8762,N_8945);
nor U10124 (N_10124,N_9436,N_9355);
xor U10125 (N_10125,N_9362,N_9828);
xor U10126 (N_10126,N_9631,N_9808);
nor U10127 (N_10127,N_9851,N_9788);
nor U10128 (N_10128,N_9249,N_9105);
nand U10129 (N_10129,N_9908,N_8752);
nand U10130 (N_10130,N_9980,N_9623);
or U10131 (N_10131,N_8811,N_9982);
nand U10132 (N_10132,N_9573,N_9554);
xor U10133 (N_10133,N_9359,N_9456);
nand U10134 (N_10134,N_9486,N_9867);
or U10135 (N_10135,N_9568,N_9113);
and U10136 (N_10136,N_9226,N_9642);
nor U10137 (N_10137,N_9383,N_9816);
and U10138 (N_10138,N_9622,N_9551);
xor U10139 (N_10139,N_9286,N_9274);
and U10140 (N_10140,N_9417,N_9878);
nand U10141 (N_10141,N_9017,N_9340);
xor U10142 (N_10142,N_9373,N_9098);
xor U10143 (N_10143,N_9640,N_9686);
xor U10144 (N_10144,N_9478,N_9526);
and U10145 (N_10145,N_9072,N_9177);
and U10146 (N_10146,N_8946,N_8830);
xor U10147 (N_10147,N_9372,N_8924);
nor U10148 (N_10148,N_9539,N_9938);
nor U10149 (N_10149,N_9247,N_9133);
and U10150 (N_10150,N_9530,N_9047);
and U10151 (N_10151,N_9489,N_9475);
nor U10152 (N_10152,N_9231,N_8906);
xor U10153 (N_10153,N_9386,N_8754);
and U10154 (N_10154,N_9435,N_9188);
or U10155 (N_10155,N_9172,N_9896);
nor U10156 (N_10156,N_9687,N_9745);
nand U10157 (N_10157,N_9458,N_9497);
nor U10158 (N_10158,N_9073,N_9968);
nand U10159 (N_10159,N_9055,N_9625);
and U10160 (N_10160,N_9213,N_9252);
or U10161 (N_10161,N_9782,N_8973);
and U10162 (N_10162,N_8980,N_9301);
and U10163 (N_10163,N_9926,N_9141);
nor U10164 (N_10164,N_9706,N_9613);
and U10165 (N_10165,N_9209,N_8799);
or U10166 (N_10166,N_8898,N_9969);
or U10167 (N_10167,N_9157,N_8797);
or U10168 (N_10168,N_8822,N_9307);
nor U10169 (N_10169,N_9027,N_9246);
nor U10170 (N_10170,N_9781,N_9743);
and U10171 (N_10171,N_9894,N_8950);
and U10172 (N_10172,N_9858,N_9575);
nand U10173 (N_10173,N_9751,N_9651);
xnor U10174 (N_10174,N_8787,N_9438);
or U10175 (N_10175,N_9152,N_9170);
xnor U10176 (N_10176,N_9096,N_9732);
or U10177 (N_10177,N_9870,N_8908);
xor U10178 (N_10178,N_9812,N_9899);
xor U10179 (N_10179,N_8955,N_9991);
and U10180 (N_10180,N_9914,N_9473);
xor U10181 (N_10181,N_9907,N_9648);
nand U10182 (N_10182,N_8995,N_8774);
xor U10183 (N_10183,N_9036,N_9571);
nand U10184 (N_10184,N_9437,N_9018);
and U10185 (N_10185,N_9621,N_9293);
nand U10186 (N_10186,N_9034,N_9811);
nor U10187 (N_10187,N_9403,N_9021);
nor U10188 (N_10188,N_8941,N_9837);
nand U10189 (N_10189,N_9863,N_8772);
nand U10190 (N_10190,N_9104,N_9074);
or U10191 (N_10191,N_9306,N_9039);
or U10192 (N_10192,N_8887,N_9518);
nand U10193 (N_10193,N_9777,N_9275);
xnor U10194 (N_10194,N_9801,N_9946);
and U10195 (N_10195,N_9345,N_9471);
or U10196 (N_10196,N_9669,N_8971);
nand U10197 (N_10197,N_8765,N_9218);
xor U10198 (N_10198,N_9419,N_9264);
or U10199 (N_10199,N_8876,N_9576);
nor U10200 (N_10200,N_9253,N_8866);
nand U10201 (N_10201,N_8970,N_9229);
nand U10202 (N_10202,N_9709,N_9465);
xor U10203 (N_10203,N_9742,N_8922);
xor U10204 (N_10204,N_8803,N_8786);
and U10205 (N_10205,N_8826,N_9708);
and U10206 (N_10206,N_9407,N_9978);
nand U10207 (N_10207,N_8923,N_9078);
or U10208 (N_10208,N_9292,N_9191);
nand U10209 (N_10209,N_9825,N_9375);
nor U10210 (N_10210,N_8759,N_9603);
nand U10211 (N_10211,N_9067,N_8961);
or U10212 (N_10212,N_8942,N_9221);
or U10213 (N_10213,N_9128,N_9587);
xnor U10214 (N_10214,N_9921,N_9434);
nor U10215 (N_10215,N_9700,N_9365);
xnor U10216 (N_10216,N_9682,N_9895);
nand U10217 (N_10217,N_9444,N_9196);
and U10218 (N_10218,N_8894,N_9194);
and U10219 (N_10219,N_9809,N_9759);
and U10220 (N_10220,N_9349,N_9443);
nor U10221 (N_10221,N_9279,N_9508);
nor U10222 (N_10222,N_8778,N_9257);
xor U10223 (N_10223,N_9679,N_9477);
nor U10224 (N_10224,N_8947,N_9917);
or U10225 (N_10225,N_9059,N_9026);
and U10226 (N_10226,N_9367,N_9124);
nand U10227 (N_10227,N_9224,N_9242);
nand U10228 (N_10228,N_9299,N_9291);
nor U10229 (N_10229,N_8854,N_9315);
nand U10230 (N_10230,N_9958,N_9061);
and U10231 (N_10231,N_9999,N_9746);
nand U10232 (N_10232,N_9987,N_9111);
xnor U10233 (N_10233,N_9397,N_9722);
xnor U10234 (N_10234,N_9861,N_9677);
or U10235 (N_10235,N_9662,N_9019);
nand U10236 (N_10236,N_9402,N_9533);
and U10237 (N_10237,N_9854,N_9418);
nand U10238 (N_10238,N_9726,N_9928);
nand U10239 (N_10239,N_9260,N_8885);
nand U10240 (N_10240,N_8957,N_9366);
xnor U10241 (N_10241,N_9884,N_9201);
nand U10242 (N_10242,N_9215,N_9845);
and U10243 (N_10243,N_9618,N_9633);
or U10244 (N_10244,N_9822,N_9927);
xnor U10245 (N_10245,N_8841,N_9755);
and U10246 (N_10246,N_9943,N_9351);
nor U10247 (N_10247,N_9206,N_9643);
xnor U10248 (N_10248,N_9063,N_9778);
or U10249 (N_10249,N_9222,N_9192);
nand U10250 (N_10250,N_8900,N_9484);
nand U10251 (N_10251,N_9597,N_9799);
nand U10252 (N_10252,N_9014,N_9841);
nand U10253 (N_10253,N_9593,N_9588);
nand U10254 (N_10254,N_9939,N_9394);
nor U10255 (N_10255,N_9904,N_9338);
nor U10256 (N_10256,N_9876,N_9881);
nor U10257 (N_10257,N_9389,N_8983);
xor U10258 (N_10258,N_9296,N_9321);
or U10259 (N_10259,N_8878,N_8990);
nand U10260 (N_10260,N_8910,N_9099);
and U10261 (N_10261,N_9937,N_9922);
xor U10262 (N_10262,N_9376,N_9243);
nor U10263 (N_10263,N_9080,N_9690);
or U10264 (N_10264,N_9327,N_9404);
nand U10265 (N_10265,N_8951,N_8905);
nand U10266 (N_10266,N_9694,N_9453);
and U10267 (N_10267,N_9832,N_9273);
nand U10268 (N_10268,N_9000,N_9122);
and U10269 (N_10269,N_9079,N_9131);
or U10270 (N_10270,N_9984,N_9570);
nand U10271 (N_10271,N_9527,N_9695);
or U10272 (N_10272,N_9398,N_8969);
or U10273 (N_10273,N_9707,N_9783);
nand U10274 (N_10274,N_9298,N_9011);
nor U10275 (N_10275,N_9802,N_9507);
xnor U10276 (N_10276,N_9885,N_9193);
or U10277 (N_10277,N_9636,N_9988);
and U10278 (N_10278,N_9425,N_9796);
nor U10279 (N_10279,N_9350,N_9422);
nor U10280 (N_10280,N_8771,N_9757);
and U10281 (N_10281,N_9254,N_9346);
nor U10282 (N_10282,N_9284,N_9161);
nand U10283 (N_10283,N_9493,N_9496);
nor U10284 (N_10284,N_9940,N_8817);
xnor U10285 (N_10285,N_9673,N_9258);
or U10286 (N_10286,N_8829,N_9962);
or U10287 (N_10287,N_9312,N_8986);
and U10288 (N_10288,N_8813,N_9439);
xor U10289 (N_10289,N_9760,N_9664);
nand U10290 (N_10290,N_8845,N_9589);
nor U10291 (N_10291,N_9482,N_9354);
nor U10292 (N_10292,N_9101,N_9612);
nand U10293 (N_10293,N_9994,N_8806);
nand U10294 (N_10294,N_9236,N_9490);
nor U10295 (N_10295,N_9583,N_9950);
and U10296 (N_10296,N_9070,N_9468);
xnor U10297 (N_10297,N_8770,N_8870);
or U10298 (N_10298,N_8851,N_9516);
or U10299 (N_10299,N_8846,N_8982);
and U10300 (N_10300,N_9829,N_9405);
and U10301 (N_10301,N_9168,N_9805);
xor U10302 (N_10302,N_8976,N_9118);
xnor U10303 (N_10303,N_8850,N_9789);
xnor U10304 (N_10304,N_9303,N_9452);
nor U10305 (N_10305,N_9949,N_9448);
or U10306 (N_10306,N_9702,N_9848);
nor U10307 (N_10307,N_9182,N_9329);
or U10308 (N_10308,N_9179,N_9947);
and U10309 (N_10309,N_9125,N_9776);
or U10310 (N_10310,N_8891,N_8897);
xnor U10311 (N_10311,N_9813,N_9174);
and U10312 (N_10312,N_9323,N_9723);
or U10313 (N_10313,N_9410,N_9705);
nand U10314 (N_10314,N_9534,N_9370);
xor U10315 (N_10315,N_9283,N_9840);
xor U10316 (N_10316,N_9956,N_9297);
xnor U10317 (N_10317,N_9369,N_9720);
nand U10318 (N_10318,N_9138,N_8801);
and U10319 (N_10319,N_9040,N_9536);
nor U10320 (N_10320,N_9771,N_9409);
nor U10321 (N_10321,N_9262,N_8918);
xor U10322 (N_10322,N_9109,N_9281);
nor U10323 (N_10323,N_9210,N_9142);
and U10324 (N_10324,N_9007,N_8981);
nand U10325 (N_10325,N_9164,N_9727);
or U10326 (N_10326,N_9454,N_9225);
nand U10327 (N_10327,N_9838,N_9305);
or U10328 (N_10328,N_8929,N_9483);
xnor U10329 (N_10329,N_8880,N_8909);
nand U10330 (N_10330,N_9650,N_9088);
nand U10331 (N_10331,N_9919,N_9584);
or U10332 (N_10332,N_9862,N_9457);
or U10333 (N_10333,N_9976,N_9380);
or U10334 (N_10334,N_8940,N_9952);
xor U10335 (N_10335,N_9933,N_9357);
nor U10336 (N_10336,N_9986,N_8966);
nor U10337 (N_10337,N_9368,N_9387);
and U10338 (N_10338,N_9476,N_8849);
nor U10339 (N_10339,N_9491,N_8881);
xor U10340 (N_10340,N_9970,N_9051);
or U10341 (N_10341,N_9266,N_9150);
and U10342 (N_10342,N_8857,N_9171);
or U10343 (N_10343,N_9343,N_9395);
nand U10344 (N_10344,N_9330,N_9235);
and U10345 (N_10345,N_9006,N_8872);
or U10346 (N_10346,N_9510,N_8937);
and U10347 (N_10347,N_9308,N_9577);
xor U10348 (N_10348,N_9020,N_9324);
nand U10349 (N_10349,N_8782,N_9767);
or U10350 (N_10350,N_9769,N_9807);
nor U10351 (N_10351,N_8949,N_9866);
or U10352 (N_10352,N_9719,N_9611);
nand U10353 (N_10353,N_9462,N_9703);
nor U10354 (N_10354,N_9241,N_9728);
nor U10355 (N_10355,N_9447,N_9620);
nor U10356 (N_10356,N_9957,N_9319);
or U10357 (N_10357,N_9996,N_9897);
and U10358 (N_10358,N_9818,N_9037);
xor U10359 (N_10359,N_9035,N_9741);
xor U10360 (N_10360,N_9429,N_9208);
and U10361 (N_10361,N_9580,N_9304);
xnor U10362 (N_10362,N_9481,N_9856);
nor U10363 (N_10363,N_9601,N_9401);
and U10364 (N_10364,N_9522,N_8994);
and U10365 (N_10365,N_9377,N_9089);
and U10366 (N_10366,N_9900,N_9967);
nor U10367 (N_10367,N_9953,N_9232);
and U10368 (N_10368,N_9711,N_8865);
nor U10369 (N_10369,N_8815,N_9175);
and U10370 (N_10370,N_9892,N_9198);
xor U10371 (N_10371,N_9149,N_8758);
xor U10372 (N_10372,N_9675,N_9207);
nor U10373 (N_10373,N_9893,N_9833);
or U10374 (N_10374,N_9176,N_9399);
xnor U10375 (N_10375,N_9780,N_9916);
xnor U10376 (N_10376,N_9317,N_9632);
and U10377 (N_10377,N_8832,N_8843);
nor U10378 (N_10378,N_9396,N_9665);
or U10379 (N_10379,N_9065,N_9730);
nand U10380 (N_10380,N_8911,N_9792);
nor U10381 (N_10381,N_9023,N_9824);
or U10382 (N_10382,N_9467,N_9738);
or U10383 (N_10383,N_9716,N_9804);
or U10384 (N_10384,N_9661,N_9764);
nand U10385 (N_10385,N_9256,N_8767);
and U10386 (N_10386,N_9734,N_9511);
or U10387 (N_10387,N_9309,N_8753);
nor U10388 (N_10388,N_9641,N_9391);
or U10389 (N_10389,N_9624,N_9543);
or U10390 (N_10390,N_9183,N_9277);
nor U10391 (N_10391,N_9075,N_8777);
and U10392 (N_10392,N_9779,N_8992);
and U10393 (N_10393,N_9485,N_9032);
nor U10394 (N_10394,N_9699,N_9517);
or U10395 (N_10395,N_9891,N_9024);
nor U10396 (N_10396,N_9156,N_9068);
xor U10397 (N_10397,N_9165,N_9328);
nand U10398 (N_10398,N_8952,N_9525);
or U10399 (N_10399,N_9320,N_9930);
nor U10400 (N_10400,N_9909,N_9140);
xor U10401 (N_10401,N_9082,N_9882);
and U10402 (N_10402,N_8890,N_9028);
nand U10403 (N_10403,N_9763,N_9639);
xnor U10404 (N_10404,N_9600,N_9721);
and U10405 (N_10405,N_9233,N_9219);
and U10406 (N_10406,N_9998,N_9245);
or U10407 (N_10407,N_9671,N_9049);
nor U10408 (N_10408,N_9136,N_8944);
and U10409 (N_10409,N_9381,N_9581);
or U10410 (N_10410,N_9087,N_9095);
nor U10411 (N_10411,N_9590,N_9294);
or U10412 (N_10412,N_9564,N_9371);
or U10413 (N_10413,N_9143,N_9244);
and U10414 (N_10414,N_8938,N_8974);
or U10415 (N_10415,N_8877,N_9674);
nand U10416 (N_10416,N_9460,N_8781);
nand U10417 (N_10417,N_9502,N_9843);
nor U10418 (N_10418,N_8960,N_9314);
nor U10419 (N_10419,N_9666,N_9869);
xor U10420 (N_10420,N_9154,N_9520);
or U10421 (N_10421,N_9045,N_9322);
and U10422 (N_10422,N_8828,N_9363);
nand U10423 (N_10423,N_9718,N_8863);
xor U10424 (N_10424,N_9426,N_9390);
nand U10425 (N_10425,N_9785,N_9216);
nand U10426 (N_10426,N_9934,N_8978);
xor U10427 (N_10427,N_9617,N_9265);
or U10428 (N_10428,N_8972,N_9965);
and U10429 (N_10429,N_8979,N_9806);
and U10430 (N_10430,N_9942,N_9029);
nor U10431 (N_10431,N_9302,N_9918);
xor U10432 (N_10432,N_8948,N_9237);
nand U10433 (N_10433,N_9003,N_9290);
or U10434 (N_10434,N_9494,N_9393);
or U10435 (N_10435,N_9288,N_9127);
and U10436 (N_10436,N_9541,N_9668);
nor U10437 (N_10437,N_9910,N_9332);
and U10438 (N_10438,N_8997,N_9503);
nand U10439 (N_10439,N_9463,N_8834);
and U10440 (N_10440,N_9585,N_9964);
and U10441 (N_10441,N_9586,N_9834);
nor U10442 (N_10442,N_8928,N_9610);
or U10443 (N_10443,N_9414,N_9849);
and U10444 (N_10444,N_9602,N_9582);
nand U10445 (N_10445,N_9791,N_8879);
or U10446 (N_10446,N_9766,N_9295);
or U10447 (N_10447,N_9120,N_9289);
and U10448 (N_10448,N_9318,N_9030);
xor U10449 (N_10449,N_9421,N_8802);
nand U10450 (N_10450,N_8852,N_9469);
or U10451 (N_10451,N_9670,N_9748);
nand U10452 (N_10452,N_9374,N_9313);
nor U10453 (N_10453,N_8820,N_9117);
xnor U10454 (N_10454,N_9731,N_9230);
nand U10455 (N_10455,N_9276,N_9509);
xor U10456 (N_10456,N_8859,N_9557);
and U10457 (N_10457,N_9971,N_9754);
nand U10458 (N_10458,N_8921,N_9768);
xnor U10459 (N_10459,N_9630,N_8769);
nor U10460 (N_10460,N_9325,N_9638);
nor U10461 (N_10461,N_9961,N_9353);
nand U10462 (N_10462,N_9523,N_9038);
nor U10463 (N_10463,N_9572,N_8789);
or U10464 (N_10464,N_9005,N_9069);
xnor U10465 (N_10465,N_9086,N_9654);
or U10466 (N_10466,N_9537,N_9656);
or U10467 (N_10467,N_9180,N_9203);
or U10468 (N_10468,N_9609,N_9538);
nor U10469 (N_10469,N_9985,N_8808);
nand U10470 (N_10470,N_9459,N_8807);
and U10471 (N_10471,N_8977,N_9724);
nand U10472 (N_10472,N_9979,N_9883);
or U10473 (N_10473,N_9693,N_9449);
nor U10474 (N_10474,N_8814,N_9552);
and U10475 (N_10475,N_9604,N_9963);
xor U10476 (N_10476,N_9794,N_8790);
or U10477 (N_10477,N_9167,N_9786);
nor U10478 (N_10478,N_8914,N_9248);
xor U10479 (N_10479,N_9553,N_9144);
nand U10480 (N_10480,N_9556,N_9110);
nand U10481 (N_10481,N_8842,N_9169);
nor U10482 (N_10482,N_8792,N_9046);
and U10483 (N_10483,N_9139,N_8761);
nor U10484 (N_10484,N_9752,N_9944);
nand U10485 (N_10485,N_9596,N_9428);
xor U10486 (N_10486,N_9263,N_9132);
nand U10487 (N_10487,N_9830,N_8775);
nor U10488 (N_10488,N_9505,N_9268);
and U10489 (N_10489,N_9282,N_9102);
xnor U10490 (N_10490,N_8919,N_8847);
and U10491 (N_10491,N_9660,N_9569);
and U10492 (N_10492,N_9285,N_9945);
and U10493 (N_10493,N_9004,N_9872);
nand U10494 (N_10494,N_9697,N_9512);
nand U10495 (N_10495,N_9663,N_9815);
and U10496 (N_10496,N_9836,N_9680);
nand U10497 (N_10497,N_9091,N_9195);
or U10498 (N_10498,N_9823,N_8987);
xor U10499 (N_10499,N_9795,N_9634);
and U10500 (N_10500,N_9972,N_9531);
nand U10501 (N_10501,N_8848,N_9566);
nor U10502 (N_10502,N_9871,N_9659);
or U10503 (N_10503,N_9852,N_8931);
nor U10504 (N_10504,N_9062,N_9826);
nand U10505 (N_10505,N_8855,N_9440);
xnor U10506 (N_10506,N_9888,N_9261);
and U10507 (N_10507,N_9647,N_9335);
or U10508 (N_10508,N_9234,N_9083);
and U10509 (N_10509,N_9672,N_9579);
nor U10510 (N_10510,N_9555,N_9797);
and U10511 (N_10511,N_8776,N_8825);
or U10512 (N_10512,N_9060,N_8932);
nand U10513 (N_10513,N_9877,N_9993);
and U10514 (N_10514,N_9574,N_9598);
nor U10515 (N_10515,N_9747,N_9750);
xnor U10516 (N_10516,N_9184,N_9920);
nand U10517 (N_10517,N_9108,N_9455);
or U10518 (N_10518,N_9644,N_9148);
or U10519 (N_10519,N_9701,N_9416);
or U10520 (N_10520,N_8959,N_9710);
or U10521 (N_10521,N_8823,N_9698);
xnor U10522 (N_10522,N_9173,N_9906);
or U10523 (N_10523,N_9115,N_9189);
xnor U10524 (N_10524,N_9793,N_9761);
nand U10525 (N_10525,N_9981,N_9311);
and U10526 (N_10526,N_8917,N_9684);
nor U10527 (N_10527,N_9499,N_8967);
nand U10528 (N_10528,N_9903,N_9608);
or U10529 (N_10529,N_9859,N_8798);
and U10530 (N_10530,N_9333,N_9810);
nand U10531 (N_10531,N_9975,N_9821);
or U10532 (N_10532,N_8856,N_9146);
xor U10533 (N_10533,N_8886,N_9774);
nor U10534 (N_10534,N_8860,N_8915);
or U10535 (N_10535,N_9217,N_9041);
nand U10536 (N_10536,N_9382,N_9488);
nand U10537 (N_10537,N_8936,N_9300);
or U10538 (N_10538,N_8963,N_9653);
or U10539 (N_10539,N_8965,N_9500);
nand U10540 (N_10540,N_8867,N_9339);
or U10541 (N_10541,N_9487,N_9056);
and U10542 (N_10542,N_9592,N_9147);
nand U10543 (N_10543,N_9817,N_9119);
xnor U10544 (N_10544,N_9151,N_9773);
xnor U10545 (N_10545,N_9126,N_9008);
xor U10546 (N_10546,N_9814,N_9211);
and U10547 (N_10547,N_9022,N_9798);
or U10548 (N_10548,N_9667,N_9480);
or U10549 (N_10549,N_9681,N_9729);
xnor U10550 (N_10550,N_8750,N_9479);
or U10551 (N_10551,N_9519,N_9658);
nor U10552 (N_10552,N_8988,N_9043);
and U10553 (N_10553,N_9220,N_9092);
xor U10554 (N_10554,N_9107,N_9446);
nor U10555 (N_10555,N_8766,N_9352);
or U10556 (N_10556,N_9002,N_9348);
nor U10557 (N_10557,N_9342,N_9240);
and U10558 (N_10558,N_9445,N_8896);
xnor U10559 (N_10559,N_9250,N_9190);
or U10560 (N_10560,N_9042,N_9765);
xor U10561 (N_10561,N_9637,N_9704);
and U10562 (N_10562,N_9432,N_8968);
nor U10563 (N_10563,N_9412,N_9737);
xor U10564 (N_10564,N_9558,N_8943);
nor U10565 (N_10565,N_9966,N_9433);
xor U10566 (N_10566,N_8930,N_9629);
nand U10567 (N_10567,N_9529,N_8907);
and U10568 (N_10568,N_9655,N_9524);
nor U10569 (N_10569,N_9819,N_8991);
or U10570 (N_10570,N_9605,N_9595);
xnor U10571 (N_10571,N_8933,N_9158);
or U10572 (N_10572,N_8768,N_9187);
xor U10573 (N_10573,N_9090,N_8882);
nor U10574 (N_10574,N_9064,N_9085);
nand U10575 (N_10575,N_8954,N_9228);
or U10576 (N_10576,N_9712,N_9646);
xnor U10577 (N_10577,N_9615,N_9890);
nor U10578 (N_10578,N_9384,N_9784);
nor U10579 (N_10579,N_9464,N_8934);
nand U10580 (N_10580,N_9071,N_9238);
and U10581 (N_10581,N_8751,N_9657);
nand U10582 (N_10582,N_9839,N_9053);
xor U10583 (N_10583,N_9627,N_8833);
nand U10584 (N_10584,N_9744,N_9202);
or U10585 (N_10585,N_9337,N_9347);
xor U10586 (N_10586,N_8873,N_9925);
nor U10587 (N_10587,N_9427,N_8763);
and U10588 (N_10588,N_9103,N_8893);
and U10589 (N_10589,N_9442,N_9400);
nand U10590 (N_10590,N_9929,N_8784);
nor U10591 (N_10591,N_8793,N_9379);
xnor U10592 (N_10592,N_9951,N_9735);
nor U10593 (N_10593,N_9739,N_8939);
nor U10594 (N_10594,N_8796,N_9451);
or U10595 (N_10595,N_9736,N_9954);
or U10596 (N_10596,N_9547,N_8757);
and U10597 (N_10597,N_8913,N_8839);
nand U10598 (N_10598,N_9923,N_9388);
nand U10599 (N_10599,N_9259,N_9860);
and U10600 (N_10600,N_9094,N_9717);
and U10601 (N_10601,N_8998,N_9411);
and U10602 (N_10602,N_9594,N_9163);
nand U10603 (N_10603,N_9902,N_9831);
or U10604 (N_10604,N_8953,N_9269);
and U10605 (N_10605,N_9178,N_9093);
nor U10606 (N_10606,N_9413,N_9145);
nand U10607 (N_10607,N_9492,N_9052);
xor U10608 (N_10608,N_8935,N_9992);
or U10609 (N_10609,N_9800,N_9874);
nor U10610 (N_10610,N_9549,N_8816);
or U10611 (N_10611,N_9591,N_8985);
nor U10612 (N_10612,N_9628,N_8920);
nand U10613 (N_10613,N_9033,N_9974);
or U10614 (N_10614,N_9535,N_9134);
nor U10615 (N_10615,N_9606,N_9271);
nor U10616 (N_10616,N_9153,N_8788);
or U10617 (N_10617,N_8835,N_9012);
nand U10618 (N_10618,N_9887,N_8884);
nor U10619 (N_10619,N_9562,N_8869);
nor U10620 (N_10620,N_9358,N_9898);
nand U10621 (N_10621,N_9715,N_9567);
or U10622 (N_10622,N_8853,N_9846);
nor U10623 (N_10623,N_9356,N_9563);
and U10624 (N_10624,N_8756,N_9941);
xnor U10625 (N_10625,N_9646,N_9896);
xor U10626 (N_10626,N_9541,N_8995);
xnor U10627 (N_10627,N_9765,N_9702);
nor U10628 (N_10628,N_9932,N_8783);
nor U10629 (N_10629,N_8860,N_9227);
xor U10630 (N_10630,N_8981,N_9711);
nor U10631 (N_10631,N_9607,N_9315);
and U10632 (N_10632,N_9185,N_9757);
or U10633 (N_10633,N_9410,N_9898);
nor U10634 (N_10634,N_8903,N_9937);
xor U10635 (N_10635,N_9147,N_9119);
nand U10636 (N_10636,N_8803,N_9523);
xor U10637 (N_10637,N_9568,N_9061);
or U10638 (N_10638,N_9631,N_8837);
or U10639 (N_10639,N_9737,N_9108);
nor U10640 (N_10640,N_9872,N_9807);
xnor U10641 (N_10641,N_9066,N_9400);
and U10642 (N_10642,N_8775,N_9143);
nor U10643 (N_10643,N_9577,N_9208);
nand U10644 (N_10644,N_9065,N_9349);
and U10645 (N_10645,N_9475,N_8894);
or U10646 (N_10646,N_8907,N_9158);
or U10647 (N_10647,N_9021,N_9723);
xor U10648 (N_10648,N_9990,N_9096);
xnor U10649 (N_10649,N_9832,N_9295);
and U10650 (N_10650,N_8996,N_8770);
xnor U10651 (N_10651,N_9723,N_9897);
and U10652 (N_10652,N_9243,N_9872);
and U10653 (N_10653,N_8987,N_9536);
nand U10654 (N_10654,N_9972,N_9768);
nor U10655 (N_10655,N_9742,N_9418);
or U10656 (N_10656,N_9953,N_9830);
nor U10657 (N_10657,N_9268,N_9223);
xnor U10658 (N_10658,N_8756,N_9489);
nand U10659 (N_10659,N_9246,N_9096);
xnor U10660 (N_10660,N_8843,N_9242);
nor U10661 (N_10661,N_8999,N_9484);
and U10662 (N_10662,N_9341,N_9889);
nor U10663 (N_10663,N_8836,N_9043);
or U10664 (N_10664,N_9914,N_8903);
or U10665 (N_10665,N_8875,N_9973);
nor U10666 (N_10666,N_9470,N_9313);
or U10667 (N_10667,N_9952,N_9459);
or U10668 (N_10668,N_9267,N_9805);
xnor U10669 (N_10669,N_9237,N_9330);
nand U10670 (N_10670,N_9686,N_9370);
or U10671 (N_10671,N_9411,N_9919);
or U10672 (N_10672,N_8764,N_9398);
xor U10673 (N_10673,N_9043,N_9221);
or U10674 (N_10674,N_9300,N_9400);
or U10675 (N_10675,N_9526,N_9609);
nor U10676 (N_10676,N_9793,N_9650);
and U10677 (N_10677,N_9832,N_9640);
nor U10678 (N_10678,N_9457,N_9950);
or U10679 (N_10679,N_9076,N_9274);
nand U10680 (N_10680,N_8898,N_8959);
nand U10681 (N_10681,N_9182,N_9750);
and U10682 (N_10682,N_9585,N_9266);
and U10683 (N_10683,N_9265,N_9631);
nand U10684 (N_10684,N_9036,N_9516);
xnor U10685 (N_10685,N_9341,N_9060);
nand U10686 (N_10686,N_8956,N_9426);
nor U10687 (N_10687,N_9248,N_9526);
nor U10688 (N_10688,N_9466,N_9796);
and U10689 (N_10689,N_9389,N_8897);
or U10690 (N_10690,N_9427,N_9740);
nor U10691 (N_10691,N_9839,N_9749);
xnor U10692 (N_10692,N_9854,N_8759);
and U10693 (N_10693,N_9515,N_9415);
xor U10694 (N_10694,N_9167,N_8772);
xor U10695 (N_10695,N_9054,N_9332);
and U10696 (N_10696,N_9745,N_9601);
xor U10697 (N_10697,N_9606,N_9249);
nor U10698 (N_10698,N_9803,N_9175);
or U10699 (N_10699,N_9316,N_9162);
nor U10700 (N_10700,N_9670,N_9111);
and U10701 (N_10701,N_8775,N_9533);
or U10702 (N_10702,N_9963,N_9417);
nor U10703 (N_10703,N_9639,N_9279);
nor U10704 (N_10704,N_9426,N_8922);
nand U10705 (N_10705,N_9589,N_8977);
xnor U10706 (N_10706,N_9915,N_9739);
nand U10707 (N_10707,N_9831,N_9381);
and U10708 (N_10708,N_9190,N_9792);
nor U10709 (N_10709,N_9937,N_9664);
xnor U10710 (N_10710,N_9569,N_9563);
nor U10711 (N_10711,N_9951,N_9416);
or U10712 (N_10712,N_9493,N_8860);
nand U10713 (N_10713,N_9203,N_9010);
nor U10714 (N_10714,N_9724,N_9911);
nand U10715 (N_10715,N_9497,N_8861);
nor U10716 (N_10716,N_9934,N_9769);
nand U10717 (N_10717,N_9078,N_8766);
or U10718 (N_10718,N_9956,N_9388);
and U10719 (N_10719,N_9156,N_9734);
or U10720 (N_10720,N_9452,N_9861);
or U10721 (N_10721,N_9978,N_8841);
or U10722 (N_10722,N_9320,N_9588);
nand U10723 (N_10723,N_9705,N_9011);
nand U10724 (N_10724,N_8761,N_9929);
nor U10725 (N_10725,N_9597,N_8981);
and U10726 (N_10726,N_9523,N_9405);
or U10727 (N_10727,N_9814,N_9285);
or U10728 (N_10728,N_9348,N_9305);
nand U10729 (N_10729,N_9347,N_9117);
nor U10730 (N_10730,N_8951,N_8965);
nand U10731 (N_10731,N_9195,N_9889);
nor U10732 (N_10732,N_9395,N_9341);
or U10733 (N_10733,N_9270,N_9770);
nand U10734 (N_10734,N_9650,N_9773);
xnor U10735 (N_10735,N_9122,N_9820);
or U10736 (N_10736,N_9407,N_9576);
nand U10737 (N_10737,N_9183,N_8948);
xnor U10738 (N_10738,N_9944,N_9988);
nand U10739 (N_10739,N_9436,N_9717);
nand U10740 (N_10740,N_9348,N_9296);
and U10741 (N_10741,N_9708,N_9206);
nand U10742 (N_10742,N_8873,N_9452);
xnor U10743 (N_10743,N_9257,N_9317);
xnor U10744 (N_10744,N_9965,N_9140);
or U10745 (N_10745,N_9057,N_9481);
xnor U10746 (N_10746,N_9935,N_9276);
and U10747 (N_10747,N_9314,N_9114);
and U10748 (N_10748,N_8879,N_9909);
nand U10749 (N_10749,N_9085,N_8989);
and U10750 (N_10750,N_9272,N_8933);
xnor U10751 (N_10751,N_9913,N_8812);
nand U10752 (N_10752,N_9539,N_9971);
and U10753 (N_10753,N_9664,N_9534);
or U10754 (N_10754,N_9430,N_8935);
nand U10755 (N_10755,N_9243,N_8772);
or U10756 (N_10756,N_9048,N_8834);
nand U10757 (N_10757,N_9402,N_8812);
or U10758 (N_10758,N_9819,N_9434);
nor U10759 (N_10759,N_8888,N_9673);
and U10760 (N_10760,N_9338,N_9850);
nand U10761 (N_10761,N_9751,N_9814);
and U10762 (N_10762,N_9040,N_8939);
and U10763 (N_10763,N_9587,N_8897);
or U10764 (N_10764,N_9742,N_9781);
or U10765 (N_10765,N_9931,N_9895);
nor U10766 (N_10766,N_9112,N_9914);
nand U10767 (N_10767,N_9488,N_8773);
xor U10768 (N_10768,N_9202,N_9428);
xnor U10769 (N_10769,N_9543,N_9711);
nor U10770 (N_10770,N_9560,N_8804);
and U10771 (N_10771,N_9118,N_9256);
nand U10772 (N_10772,N_9571,N_9244);
or U10773 (N_10773,N_9357,N_9349);
nand U10774 (N_10774,N_8962,N_9541);
nor U10775 (N_10775,N_9032,N_9615);
and U10776 (N_10776,N_9003,N_9439);
nor U10777 (N_10777,N_9896,N_9107);
nand U10778 (N_10778,N_8975,N_9731);
nand U10779 (N_10779,N_9630,N_9563);
nand U10780 (N_10780,N_9722,N_8823);
nor U10781 (N_10781,N_9444,N_8767);
or U10782 (N_10782,N_9181,N_9652);
xor U10783 (N_10783,N_9140,N_9327);
nand U10784 (N_10784,N_8811,N_9208);
nor U10785 (N_10785,N_9910,N_9752);
xor U10786 (N_10786,N_9824,N_9457);
and U10787 (N_10787,N_9093,N_9794);
xor U10788 (N_10788,N_9761,N_9111);
nand U10789 (N_10789,N_9942,N_8794);
and U10790 (N_10790,N_9422,N_9608);
or U10791 (N_10791,N_9697,N_9328);
xor U10792 (N_10792,N_9247,N_9120);
and U10793 (N_10793,N_9653,N_8765);
xor U10794 (N_10794,N_9223,N_9179);
nand U10795 (N_10795,N_9668,N_9827);
nand U10796 (N_10796,N_9810,N_9593);
xor U10797 (N_10797,N_9436,N_9026);
xor U10798 (N_10798,N_9578,N_9744);
nand U10799 (N_10799,N_9135,N_8912);
and U10800 (N_10800,N_8863,N_9532);
xor U10801 (N_10801,N_9058,N_9744);
or U10802 (N_10802,N_9466,N_9747);
nand U10803 (N_10803,N_9260,N_9813);
nand U10804 (N_10804,N_8962,N_9054);
and U10805 (N_10805,N_9041,N_8807);
nand U10806 (N_10806,N_9668,N_9867);
and U10807 (N_10807,N_9080,N_9904);
and U10808 (N_10808,N_9721,N_9726);
nor U10809 (N_10809,N_8954,N_9621);
and U10810 (N_10810,N_9586,N_8969);
nand U10811 (N_10811,N_8924,N_9441);
nand U10812 (N_10812,N_8773,N_9800);
or U10813 (N_10813,N_9197,N_8898);
and U10814 (N_10814,N_9328,N_9669);
nand U10815 (N_10815,N_9630,N_8838);
nand U10816 (N_10816,N_9768,N_9367);
nor U10817 (N_10817,N_9240,N_8994);
nor U10818 (N_10818,N_9914,N_9751);
nand U10819 (N_10819,N_9928,N_9503);
or U10820 (N_10820,N_9271,N_9779);
nand U10821 (N_10821,N_9369,N_9186);
nand U10822 (N_10822,N_9776,N_9780);
nor U10823 (N_10823,N_9923,N_9951);
or U10824 (N_10824,N_9882,N_9079);
or U10825 (N_10825,N_9739,N_9107);
nand U10826 (N_10826,N_8774,N_9698);
and U10827 (N_10827,N_9723,N_9416);
nand U10828 (N_10828,N_9193,N_9548);
nand U10829 (N_10829,N_9789,N_9781);
or U10830 (N_10830,N_9887,N_9443);
and U10831 (N_10831,N_8836,N_9498);
or U10832 (N_10832,N_8981,N_9884);
or U10833 (N_10833,N_9600,N_9896);
nor U10834 (N_10834,N_9027,N_9041);
or U10835 (N_10835,N_9108,N_8939);
nor U10836 (N_10836,N_9474,N_8987);
xnor U10837 (N_10837,N_9346,N_8920);
nor U10838 (N_10838,N_8934,N_9833);
and U10839 (N_10839,N_9456,N_9429);
nand U10840 (N_10840,N_9958,N_8923);
nand U10841 (N_10841,N_9918,N_9282);
nand U10842 (N_10842,N_9468,N_9003);
xor U10843 (N_10843,N_8847,N_8817);
nor U10844 (N_10844,N_9822,N_9165);
and U10845 (N_10845,N_8961,N_9973);
nand U10846 (N_10846,N_9136,N_9423);
or U10847 (N_10847,N_8854,N_9076);
xor U10848 (N_10848,N_9220,N_9309);
and U10849 (N_10849,N_9999,N_8919);
xor U10850 (N_10850,N_8924,N_9973);
and U10851 (N_10851,N_8911,N_8765);
nor U10852 (N_10852,N_9948,N_9688);
and U10853 (N_10853,N_9494,N_9038);
and U10854 (N_10854,N_9016,N_9688);
nand U10855 (N_10855,N_9472,N_9547);
and U10856 (N_10856,N_9571,N_9781);
and U10857 (N_10857,N_9808,N_9391);
nand U10858 (N_10858,N_9080,N_9317);
nand U10859 (N_10859,N_9199,N_9045);
xor U10860 (N_10860,N_9570,N_9514);
or U10861 (N_10861,N_9776,N_9748);
xor U10862 (N_10862,N_9614,N_8846);
nand U10863 (N_10863,N_9491,N_8766);
and U10864 (N_10864,N_9875,N_8807);
nor U10865 (N_10865,N_9025,N_9623);
and U10866 (N_10866,N_9392,N_8946);
and U10867 (N_10867,N_9153,N_9618);
nor U10868 (N_10868,N_9337,N_9731);
and U10869 (N_10869,N_9797,N_8792);
xnor U10870 (N_10870,N_9481,N_9039);
xor U10871 (N_10871,N_9270,N_8780);
nor U10872 (N_10872,N_9950,N_8785);
nand U10873 (N_10873,N_9547,N_9336);
nand U10874 (N_10874,N_9712,N_9713);
nor U10875 (N_10875,N_9205,N_9614);
and U10876 (N_10876,N_9520,N_9158);
xnor U10877 (N_10877,N_9088,N_9166);
and U10878 (N_10878,N_9464,N_9767);
or U10879 (N_10879,N_8863,N_8939);
or U10880 (N_10880,N_9297,N_8939);
xnor U10881 (N_10881,N_9895,N_9317);
nor U10882 (N_10882,N_8879,N_8904);
and U10883 (N_10883,N_8856,N_9119);
nor U10884 (N_10884,N_9100,N_8883);
or U10885 (N_10885,N_9133,N_8947);
nand U10886 (N_10886,N_9834,N_8911);
or U10887 (N_10887,N_9707,N_8924);
nor U10888 (N_10888,N_9091,N_9380);
and U10889 (N_10889,N_9778,N_8758);
xor U10890 (N_10890,N_8910,N_9150);
xor U10891 (N_10891,N_9153,N_8976);
xnor U10892 (N_10892,N_9888,N_9809);
or U10893 (N_10893,N_9195,N_9181);
or U10894 (N_10894,N_9957,N_9394);
and U10895 (N_10895,N_9076,N_8887);
xnor U10896 (N_10896,N_8815,N_9797);
nor U10897 (N_10897,N_9737,N_9359);
or U10898 (N_10898,N_9253,N_8783);
or U10899 (N_10899,N_8773,N_9867);
xor U10900 (N_10900,N_9564,N_8844);
and U10901 (N_10901,N_9637,N_9787);
and U10902 (N_10902,N_9821,N_9658);
nand U10903 (N_10903,N_9688,N_9794);
xnor U10904 (N_10904,N_9114,N_8952);
nor U10905 (N_10905,N_9284,N_9187);
or U10906 (N_10906,N_8822,N_9725);
nand U10907 (N_10907,N_8818,N_9720);
or U10908 (N_10908,N_9862,N_8754);
xor U10909 (N_10909,N_9656,N_9431);
nor U10910 (N_10910,N_9914,N_8764);
nor U10911 (N_10911,N_9323,N_9012);
xnor U10912 (N_10912,N_9692,N_9658);
nand U10913 (N_10913,N_9399,N_8993);
nor U10914 (N_10914,N_9485,N_9375);
nand U10915 (N_10915,N_9393,N_9206);
nor U10916 (N_10916,N_9679,N_9203);
or U10917 (N_10917,N_9779,N_8928);
nor U10918 (N_10918,N_8777,N_9877);
xor U10919 (N_10919,N_9731,N_9176);
or U10920 (N_10920,N_9490,N_9004);
or U10921 (N_10921,N_9492,N_9290);
xor U10922 (N_10922,N_9920,N_9494);
nor U10923 (N_10923,N_9248,N_9785);
or U10924 (N_10924,N_9848,N_8841);
and U10925 (N_10925,N_9249,N_9323);
nor U10926 (N_10926,N_9607,N_9858);
and U10927 (N_10927,N_9949,N_9088);
nand U10928 (N_10928,N_9815,N_9869);
nand U10929 (N_10929,N_9065,N_9073);
xnor U10930 (N_10930,N_9632,N_8894);
and U10931 (N_10931,N_9111,N_9790);
nand U10932 (N_10932,N_9067,N_9622);
nand U10933 (N_10933,N_9099,N_9169);
and U10934 (N_10934,N_9748,N_9978);
and U10935 (N_10935,N_9454,N_9976);
nand U10936 (N_10936,N_9017,N_9195);
or U10937 (N_10937,N_9509,N_9199);
nand U10938 (N_10938,N_8880,N_9010);
xnor U10939 (N_10939,N_9772,N_9941);
nand U10940 (N_10940,N_9403,N_9318);
and U10941 (N_10941,N_9229,N_8940);
nand U10942 (N_10942,N_9551,N_9489);
or U10943 (N_10943,N_9349,N_9464);
nor U10944 (N_10944,N_9268,N_9740);
nand U10945 (N_10945,N_9575,N_9840);
nor U10946 (N_10946,N_9052,N_8931);
nor U10947 (N_10947,N_9080,N_9465);
xnor U10948 (N_10948,N_9749,N_9842);
nand U10949 (N_10949,N_9461,N_8826);
nor U10950 (N_10950,N_9867,N_9610);
xnor U10951 (N_10951,N_8962,N_9382);
xnor U10952 (N_10952,N_9294,N_9048);
or U10953 (N_10953,N_9979,N_9429);
or U10954 (N_10954,N_9771,N_9274);
or U10955 (N_10955,N_9397,N_8816);
and U10956 (N_10956,N_9697,N_9963);
and U10957 (N_10957,N_8945,N_9754);
nand U10958 (N_10958,N_9502,N_9240);
xor U10959 (N_10959,N_8881,N_8903);
nor U10960 (N_10960,N_9718,N_9571);
or U10961 (N_10961,N_9359,N_9823);
xnor U10962 (N_10962,N_9037,N_8949);
or U10963 (N_10963,N_9650,N_8954);
nand U10964 (N_10964,N_9420,N_9144);
or U10965 (N_10965,N_8947,N_9717);
or U10966 (N_10966,N_9647,N_9466);
and U10967 (N_10967,N_9591,N_8844);
nor U10968 (N_10968,N_9056,N_9339);
or U10969 (N_10969,N_8958,N_9672);
and U10970 (N_10970,N_9614,N_9430);
nand U10971 (N_10971,N_9689,N_8820);
nor U10972 (N_10972,N_9063,N_9809);
and U10973 (N_10973,N_9003,N_9001);
nand U10974 (N_10974,N_8753,N_8847);
or U10975 (N_10975,N_9522,N_9559);
nand U10976 (N_10976,N_9264,N_9062);
and U10977 (N_10977,N_9845,N_9697);
xnor U10978 (N_10978,N_8998,N_9448);
xor U10979 (N_10979,N_9039,N_8890);
and U10980 (N_10980,N_8910,N_9478);
and U10981 (N_10981,N_9770,N_9108);
and U10982 (N_10982,N_9357,N_9616);
and U10983 (N_10983,N_9696,N_8869);
nand U10984 (N_10984,N_9554,N_9492);
nand U10985 (N_10985,N_9361,N_9079);
and U10986 (N_10986,N_9427,N_9408);
and U10987 (N_10987,N_9501,N_9526);
and U10988 (N_10988,N_9530,N_9263);
and U10989 (N_10989,N_9532,N_9377);
xnor U10990 (N_10990,N_9740,N_9859);
nor U10991 (N_10991,N_9896,N_9775);
xnor U10992 (N_10992,N_9822,N_9913);
or U10993 (N_10993,N_9145,N_9878);
xnor U10994 (N_10994,N_9305,N_9611);
xnor U10995 (N_10995,N_9725,N_9438);
nor U10996 (N_10996,N_9816,N_9765);
or U10997 (N_10997,N_9861,N_9533);
nand U10998 (N_10998,N_8839,N_9518);
and U10999 (N_10999,N_9368,N_8803);
and U11000 (N_11000,N_9011,N_9201);
xnor U11001 (N_11001,N_8957,N_8799);
and U11002 (N_11002,N_9280,N_9906);
nand U11003 (N_11003,N_9303,N_9636);
nor U11004 (N_11004,N_9187,N_9103);
nor U11005 (N_11005,N_9293,N_9497);
and U11006 (N_11006,N_9356,N_9930);
and U11007 (N_11007,N_9558,N_8966);
and U11008 (N_11008,N_9780,N_8911);
nand U11009 (N_11009,N_9230,N_9996);
xor U11010 (N_11010,N_9209,N_9107);
nand U11011 (N_11011,N_8973,N_9881);
nor U11012 (N_11012,N_9978,N_9634);
nor U11013 (N_11013,N_9972,N_9999);
nor U11014 (N_11014,N_9928,N_9230);
nor U11015 (N_11015,N_9098,N_9976);
nor U11016 (N_11016,N_9447,N_8994);
nand U11017 (N_11017,N_9425,N_9746);
xor U11018 (N_11018,N_9636,N_8983);
or U11019 (N_11019,N_9185,N_9452);
and U11020 (N_11020,N_9170,N_8815);
and U11021 (N_11021,N_9003,N_9353);
and U11022 (N_11022,N_9088,N_9563);
nand U11023 (N_11023,N_9138,N_9223);
or U11024 (N_11024,N_9085,N_8779);
xnor U11025 (N_11025,N_9066,N_8970);
nand U11026 (N_11026,N_9197,N_9443);
nand U11027 (N_11027,N_9496,N_9658);
or U11028 (N_11028,N_9920,N_9043);
or U11029 (N_11029,N_9870,N_9986);
and U11030 (N_11030,N_9503,N_9843);
xnor U11031 (N_11031,N_9836,N_8754);
nand U11032 (N_11032,N_8755,N_8988);
nand U11033 (N_11033,N_9437,N_9826);
nand U11034 (N_11034,N_8889,N_9205);
and U11035 (N_11035,N_9428,N_9236);
and U11036 (N_11036,N_9831,N_8887);
or U11037 (N_11037,N_9033,N_9016);
xnor U11038 (N_11038,N_8870,N_9221);
xnor U11039 (N_11039,N_9880,N_9910);
or U11040 (N_11040,N_9206,N_8786);
nor U11041 (N_11041,N_9470,N_8813);
nor U11042 (N_11042,N_9482,N_9397);
nor U11043 (N_11043,N_9239,N_9743);
and U11044 (N_11044,N_9151,N_9256);
and U11045 (N_11045,N_9456,N_9514);
nand U11046 (N_11046,N_9889,N_9096);
nand U11047 (N_11047,N_9138,N_8887);
xor U11048 (N_11048,N_9236,N_9272);
xnor U11049 (N_11049,N_8996,N_8756);
xnor U11050 (N_11050,N_9458,N_9310);
nor U11051 (N_11051,N_9463,N_9342);
nand U11052 (N_11052,N_8966,N_9315);
and U11053 (N_11053,N_9243,N_8841);
nand U11054 (N_11054,N_9198,N_9577);
and U11055 (N_11055,N_9624,N_8993);
nor U11056 (N_11056,N_9440,N_9157);
and U11057 (N_11057,N_9653,N_9008);
or U11058 (N_11058,N_9338,N_9846);
or U11059 (N_11059,N_9058,N_9700);
or U11060 (N_11060,N_9516,N_9922);
xor U11061 (N_11061,N_9821,N_9310);
xor U11062 (N_11062,N_9196,N_9971);
nand U11063 (N_11063,N_9424,N_8819);
nand U11064 (N_11064,N_8834,N_9145);
nor U11065 (N_11065,N_9367,N_9962);
xor U11066 (N_11066,N_9069,N_8880);
nor U11067 (N_11067,N_9223,N_9604);
and U11068 (N_11068,N_9660,N_8890);
xor U11069 (N_11069,N_9241,N_9470);
xor U11070 (N_11070,N_9039,N_9210);
nand U11071 (N_11071,N_8891,N_9608);
and U11072 (N_11072,N_9712,N_9636);
nand U11073 (N_11073,N_8965,N_9111);
nor U11074 (N_11074,N_8780,N_9557);
and U11075 (N_11075,N_8757,N_9664);
nand U11076 (N_11076,N_9040,N_9474);
nor U11077 (N_11077,N_9682,N_9033);
nor U11078 (N_11078,N_9758,N_9189);
nand U11079 (N_11079,N_9665,N_9769);
nor U11080 (N_11080,N_8840,N_8886);
nor U11081 (N_11081,N_9804,N_9709);
nand U11082 (N_11082,N_9497,N_9532);
nand U11083 (N_11083,N_9222,N_9267);
nand U11084 (N_11084,N_8962,N_9621);
xor U11085 (N_11085,N_9872,N_9230);
nand U11086 (N_11086,N_9539,N_9849);
nand U11087 (N_11087,N_9965,N_8916);
nor U11088 (N_11088,N_9400,N_8855);
nand U11089 (N_11089,N_9271,N_9013);
and U11090 (N_11090,N_9839,N_8991);
nor U11091 (N_11091,N_8826,N_9878);
nand U11092 (N_11092,N_8816,N_9170);
nor U11093 (N_11093,N_9948,N_9073);
xnor U11094 (N_11094,N_9910,N_9625);
xnor U11095 (N_11095,N_9260,N_9405);
nand U11096 (N_11096,N_9915,N_9338);
and U11097 (N_11097,N_9300,N_8769);
or U11098 (N_11098,N_9960,N_9293);
xor U11099 (N_11099,N_9794,N_8762);
nor U11100 (N_11100,N_8927,N_9366);
or U11101 (N_11101,N_9200,N_9878);
nor U11102 (N_11102,N_8887,N_9250);
xnor U11103 (N_11103,N_9957,N_8994);
xor U11104 (N_11104,N_9902,N_8759);
and U11105 (N_11105,N_8786,N_9168);
nor U11106 (N_11106,N_9003,N_9303);
nor U11107 (N_11107,N_9267,N_9489);
and U11108 (N_11108,N_9571,N_8771);
xnor U11109 (N_11109,N_9994,N_9464);
and U11110 (N_11110,N_9158,N_9537);
or U11111 (N_11111,N_9889,N_9430);
or U11112 (N_11112,N_9625,N_9084);
and U11113 (N_11113,N_9380,N_9243);
xor U11114 (N_11114,N_8934,N_9858);
and U11115 (N_11115,N_9066,N_9245);
nor U11116 (N_11116,N_9911,N_9657);
nand U11117 (N_11117,N_9680,N_9675);
nand U11118 (N_11118,N_9098,N_9315);
nor U11119 (N_11119,N_9669,N_8921);
nor U11120 (N_11120,N_9398,N_9931);
nor U11121 (N_11121,N_9079,N_9037);
or U11122 (N_11122,N_9133,N_9335);
nor U11123 (N_11123,N_9194,N_8874);
or U11124 (N_11124,N_8888,N_9459);
nand U11125 (N_11125,N_9909,N_9819);
xor U11126 (N_11126,N_9924,N_8911);
nand U11127 (N_11127,N_9751,N_9200);
or U11128 (N_11128,N_9015,N_9938);
xnor U11129 (N_11129,N_9096,N_9981);
or U11130 (N_11130,N_9898,N_9175);
xnor U11131 (N_11131,N_9378,N_9435);
or U11132 (N_11132,N_9513,N_9506);
nor U11133 (N_11133,N_9001,N_8925);
or U11134 (N_11134,N_9528,N_9899);
nor U11135 (N_11135,N_9234,N_8811);
xor U11136 (N_11136,N_9819,N_8757);
or U11137 (N_11137,N_9889,N_9371);
xor U11138 (N_11138,N_9170,N_9318);
nor U11139 (N_11139,N_9031,N_9408);
nand U11140 (N_11140,N_9214,N_9226);
or U11141 (N_11141,N_9369,N_9115);
nor U11142 (N_11142,N_8878,N_9987);
and U11143 (N_11143,N_9667,N_9739);
and U11144 (N_11144,N_9330,N_9689);
nor U11145 (N_11145,N_9915,N_9881);
nand U11146 (N_11146,N_9130,N_9673);
nand U11147 (N_11147,N_8861,N_9144);
nor U11148 (N_11148,N_9476,N_9347);
or U11149 (N_11149,N_9360,N_9777);
xor U11150 (N_11150,N_9989,N_9710);
xnor U11151 (N_11151,N_8906,N_9430);
nand U11152 (N_11152,N_9622,N_8817);
nand U11153 (N_11153,N_9637,N_9507);
or U11154 (N_11154,N_9135,N_9366);
xnor U11155 (N_11155,N_9501,N_8771);
nand U11156 (N_11156,N_9314,N_8844);
nor U11157 (N_11157,N_9571,N_9567);
nand U11158 (N_11158,N_9496,N_9193);
xnor U11159 (N_11159,N_8838,N_9677);
and U11160 (N_11160,N_9089,N_9857);
nor U11161 (N_11161,N_8930,N_8936);
xnor U11162 (N_11162,N_8894,N_9317);
nor U11163 (N_11163,N_8909,N_9457);
xor U11164 (N_11164,N_9737,N_9762);
nor U11165 (N_11165,N_9612,N_9986);
and U11166 (N_11166,N_8992,N_9356);
and U11167 (N_11167,N_9294,N_9425);
xor U11168 (N_11168,N_9926,N_9292);
xnor U11169 (N_11169,N_9759,N_9619);
nand U11170 (N_11170,N_8862,N_9782);
and U11171 (N_11171,N_9955,N_9250);
or U11172 (N_11172,N_9135,N_9978);
nor U11173 (N_11173,N_9458,N_9993);
xnor U11174 (N_11174,N_9008,N_9400);
or U11175 (N_11175,N_9504,N_9016);
and U11176 (N_11176,N_9729,N_9898);
nor U11177 (N_11177,N_9916,N_9467);
or U11178 (N_11178,N_9613,N_9470);
xor U11179 (N_11179,N_8934,N_9090);
and U11180 (N_11180,N_9516,N_9749);
and U11181 (N_11181,N_9523,N_9943);
nor U11182 (N_11182,N_9120,N_9098);
nor U11183 (N_11183,N_9640,N_9339);
xor U11184 (N_11184,N_9243,N_8851);
nor U11185 (N_11185,N_8985,N_9438);
and U11186 (N_11186,N_9596,N_9931);
or U11187 (N_11187,N_9787,N_9662);
and U11188 (N_11188,N_8956,N_9150);
and U11189 (N_11189,N_9564,N_9538);
nor U11190 (N_11190,N_9234,N_8883);
xnor U11191 (N_11191,N_9625,N_9801);
and U11192 (N_11192,N_8830,N_9978);
or U11193 (N_11193,N_8941,N_9255);
and U11194 (N_11194,N_9710,N_9623);
nor U11195 (N_11195,N_9544,N_8824);
nand U11196 (N_11196,N_9985,N_9455);
nand U11197 (N_11197,N_9364,N_9650);
nand U11198 (N_11198,N_9010,N_9160);
nor U11199 (N_11199,N_9472,N_9790);
nand U11200 (N_11200,N_9855,N_9216);
xor U11201 (N_11201,N_9765,N_9734);
xnor U11202 (N_11202,N_9745,N_9059);
nand U11203 (N_11203,N_9507,N_9734);
xnor U11204 (N_11204,N_9474,N_9760);
nand U11205 (N_11205,N_8879,N_9929);
nor U11206 (N_11206,N_9559,N_9994);
or U11207 (N_11207,N_9773,N_9997);
nor U11208 (N_11208,N_9377,N_9395);
xnor U11209 (N_11209,N_9606,N_9405);
nand U11210 (N_11210,N_9515,N_9654);
nand U11211 (N_11211,N_8990,N_9769);
nor U11212 (N_11212,N_9789,N_9967);
nor U11213 (N_11213,N_8927,N_9678);
nor U11214 (N_11214,N_9167,N_9273);
nor U11215 (N_11215,N_9277,N_9092);
nor U11216 (N_11216,N_8757,N_9477);
or U11217 (N_11217,N_9395,N_9088);
or U11218 (N_11218,N_9600,N_9227);
nand U11219 (N_11219,N_9461,N_9279);
nor U11220 (N_11220,N_8830,N_9192);
and U11221 (N_11221,N_9581,N_9175);
xor U11222 (N_11222,N_9206,N_9689);
xor U11223 (N_11223,N_8916,N_9307);
or U11224 (N_11224,N_8809,N_9396);
nand U11225 (N_11225,N_9692,N_9024);
nand U11226 (N_11226,N_9081,N_9196);
and U11227 (N_11227,N_9957,N_9708);
xnor U11228 (N_11228,N_9389,N_9738);
nand U11229 (N_11229,N_9246,N_8925);
and U11230 (N_11230,N_8952,N_8892);
xor U11231 (N_11231,N_9354,N_9617);
nor U11232 (N_11232,N_9589,N_9141);
nor U11233 (N_11233,N_9581,N_9343);
nand U11234 (N_11234,N_9945,N_9566);
or U11235 (N_11235,N_8921,N_8798);
and U11236 (N_11236,N_9143,N_9114);
or U11237 (N_11237,N_9799,N_9173);
xnor U11238 (N_11238,N_9382,N_9421);
nand U11239 (N_11239,N_8809,N_9405);
xnor U11240 (N_11240,N_9473,N_8880);
nand U11241 (N_11241,N_9966,N_9906);
or U11242 (N_11242,N_9196,N_9591);
xor U11243 (N_11243,N_8758,N_9597);
nand U11244 (N_11244,N_8935,N_9796);
nor U11245 (N_11245,N_9059,N_9493);
and U11246 (N_11246,N_9898,N_9752);
or U11247 (N_11247,N_8964,N_9442);
and U11248 (N_11248,N_9917,N_8897);
and U11249 (N_11249,N_9796,N_9450);
or U11250 (N_11250,N_11115,N_10745);
nor U11251 (N_11251,N_10699,N_10439);
nor U11252 (N_11252,N_10487,N_10113);
nor U11253 (N_11253,N_11096,N_10001);
and U11254 (N_11254,N_10638,N_10491);
or U11255 (N_11255,N_11244,N_11010);
nand U11256 (N_11256,N_10870,N_10684);
nor U11257 (N_11257,N_11190,N_10226);
nand U11258 (N_11258,N_10622,N_10337);
xnor U11259 (N_11259,N_10136,N_10819);
nand U11260 (N_11260,N_11024,N_11229);
xor U11261 (N_11261,N_10237,N_10567);
nand U11262 (N_11262,N_11088,N_10164);
nand U11263 (N_11263,N_10719,N_10489);
xor U11264 (N_11264,N_10109,N_10677);
nand U11265 (N_11265,N_10633,N_10694);
and U11266 (N_11266,N_10325,N_10373);
nand U11267 (N_11267,N_10620,N_10752);
nand U11268 (N_11268,N_10347,N_10176);
nor U11269 (N_11269,N_11025,N_10030);
nor U11270 (N_11270,N_10857,N_10438);
and U11271 (N_11271,N_10406,N_10624);
nand U11272 (N_11272,N_10251,N_11112);
and U11273 (N_11273,N_10314,N_10845);
nand U11274 (N_11274,N_10805,N_10046);
or U11275 (N_11275,N_10957,N_10207);
nand U11276 (N_11276,N_10568,N_10602);
xnor U11277 (N_11277,N_10648,N_10312);
xnor U11278 (N_11278,N_11079,N_10322);
and U11279 (N_11279,N_10658,N_10381);
and U11280 (N_11280,N_10466,N_10728);
nor U11281 (N_11281,N_10405,N_10354);
nor U11282 (N_11282,N_10925,N_10274);
nand U11283 (N_11283,N_10261,N_10972);
xor U11284 (N_11284,N_10609,N_10588);
nand U11285 (N_11285,N_10475,N_10287);
nand U11286 (N_11286,N_10511,N_10838);
nand U11287 (N_11287,N_10157,N_10241);
xor U11288 (N_11288,N_11071,N_10024);
or U11289 (N_11289,N_10172,N_10636);
nor U11290 (N_11290,N_10121,N_10239);
or U11291 (N_11291,N_10167,N_10643);
nor U11292 (N_11292,N_10947,N_10931);
nand U11293 (N_11293,N_10402,N_11098);
and U11294 (N_11294,N_11133,N_10865);
nand U11295 (N_11295,N_11234,N_11018);
nor U11296 (N_11296,N_10666,N_10263);
xnor U11297 (N_11297,N_11152,N_10515);
nand U11298 (N_11298,N_10090,N_10125);
and U11299 (N_11299,N_10413,N_11198);
xnor U11300 (N_11300,N_11175,N_11162);
and U11301 (N_11301,N_10899,N_10985);
or U11302 (N_11302,N_10607,N_10232);
or U11303 (N_11303,N_10247,N_10929);
nor U11304 (N_11304,N_10321,N_10968);
nand U11305 (N_11305,N_10163,N_10344);
nand U11306 (N_11306,N_10143,N_10565);
and U11307 (N_11307,N_10131,N_11203);
or U11308 (N_11308,N_10371,N_10437);
xnor U11309 (N_11309,N_11072,N_10986);
xnor U11310 (N_11310,N_10970,N_10800);
nand U11311 (N_11311,N_10932,N_10123);
nand U11312 (N_11312,N_10988,N_10982);
xor U11313 (N_11313,N_11182,N_10890);
or U11314 (N_11314,N_10062,N_10478);
xnor U11315 (N_11315,N_10540,N_10732);
and U11316 (N_11316,N_10723,N_10353);
nor U11317 (N_11317,N_10161,N_10539);
nor U11318 (N_11318,N_10761,N_10180);
nor U11319 (N_11319,N_10403,N_10252);
and U11320 (N_11320,N_11180,N_11002);
xor U11321 (N_11321,N_10302,N_10014);
nor U11322 (N_11322,N_10702,N_10514);
or U11323 (N_11323,N_10996,N_10803);
xor U11324 (N_11324,N_11075,N_10502);
nor U11325 (N_11325,N_11150,N_10862);
and U11326 (N_11326,N_11011,N_10093);
or U11327 (N_11327,N_10115,N_11038);
and U11328 (N_11328,N_10335,N_10979);
or U11329 (N_11329,N_11099,N_11086);
nor U11330 (N_11330,N_10298,N_11247);
or U11331 (N_11331,N_10535,N_10114);
and U11332 (N_11332,N_10482,N_10356);
nand U11333 (N_11333,N_10903,N_10560);
nor U11334 (N_11334,N_10778,N_10612);
or U11335 (N_11335,N_11046,N_10610);
and U11336 (N_11336,N_10717,N_10348);
nand U11337 (N_11337,N_11087,N_10842);
and U11338 (N_11338,N_11246,N_11021);
nor U11339 (N_11339,N_10672,N_10757);
nor U11340 (N_11340,N_10811,N_11053);
xnor U11341 (N_11341,N_10944,N_10409);
nand U11342 (N_11342,N_11070,N_11212);
xnor U11343 (N_11343,N_10762,N_10202);
xor U11344 (N_11344,N_10149,N_10860);
nor U11345 (N_11345,N_10155,N_10372);
xnor U11346 (N_11346,N_10645,N_11248);
and U11347 (N_11347,N_10606,N_10965);
xnor U11348 (N_11348,N_10041,N_11055);
xor U11349 (N_11349,N_11197,N_10240);
and U11350 (N_11350,N_10179,N_11037);
nand U11351 (N_11351,N_10848,N_10178);
nand U11352 (N_11352,N_11137,N_10594);
or U11353 (N_11353,N_10910,N_11135);
xnor U11354 (N_11354,N_10993,N_10512);
or U11355 (N_11355,N_10122,N_10933);
nand U11356 (N_11356,N_10391,N_11184);
and U11357 (N_11357,N_10311,N_10559);
nor U11358 (N_11358,N_10912,N_10562);
or U11359 (N_11359,N_11176,N_10005);
or U11360 (N_11360,N_10962,N_11146);
nand U11361 (N_11361,N_10357,N_11149);
nor U11362 (N_11362,N_11016,N_10940);
nand U11363 (N_11363,N_11008,N_10906);
nand U11364 (N_11364,N_10147,N_10279);
or U11365 (N_11365,N_10936,N_10119);
nand U11366 (N_11366,N_10795,N_10966);
and U11367 (N_11367,N_10174,N_10215);
xnor U11368 (N_11368,N_10013,N_10448);
nor U11369 (N_11369,N_10937,N_10764);
nor U11370 (N_11370,N_10384,N_10952);
xor U11371 (N_11371,N_10880,N_10742);
nor U11372 (N_11372,N_10774,N_10023);
and U11373 (N_11373,N_10961,N_10255);
nand U11374 (N_11374,N_10159,N_11007);
nand U11375 (N_11375,N_11089,N_10632);
xor U11376 (N_11376,N_10958,N_10182);
nand U11377 (N_11377,N_10429,N_10729);
and U11378 (N_11378,N_10044,N_10854);
nor U11379 (N_11379,N_10470,N_10850);
xor U11380 (N_11380,N_10126,N_10901);
nor U11381 (N_11381,N_11210,N_10493);
or U11382 (N_11382,N_10999,N_10718);
xnor U11383 (N_11383,N_10110,N_10802);
and U11384 (N_11384,N_10206,N_10045);
and U11385 (N_11385,N_10118,N_11066);
nand U11386 (N_11386,N_10359,N_10276);
xnor U11387 (N_11387,N_10705,N_10821);
xor U11388 (N_11388,N_11104,N_10399);
xor U11389 (N_11389,N_10290,N_11056);
xor U11390 (N_11390,N_10080,N_10473);
xnor U11391 (N_11391,N_10809,N_11111);
nor U11392 (N_11392,N_11217,N_10676);
nor U11393 (N_11393,N_11042,N_10220);
xnor U11394 (N_11394,N_10871,N_10836);
nand U11395 (N_11395,N_10146,N_10522);
nor U11396 (N_11396,N_11123,N_10071);
nand U11397 (N_11397,N_10832,N_10716);
or U11398 (N_11398,N_10589,N_11033);
xor U11399 (N_11399,N_10479,N_10459);
nand U11400 (N_11400,N_11051,N_10526);
xnor U11401 (N_11401,N_10224,N_11142);
nor U11402 (N_11402,N_10410,N_11131);
and U11403 (N_11403,N_10389,N_11174);
nor U11404 (N_11404,N_10004,N_10012);
nor U11405 (N_11405,N_10987,N_10449);
xor U11406 (N_11406,N_10379,N_10316);
and U11407 (N_11407,N_11200,N_11035);
or U11408 (N_11408,N_11084,N_10219);
and U11409 (N_11409,N_10245,N_10746);
nor U11410 (N_11410,N_10758,N_10072);
nor U11411 (N_11411,N_10955,N_10657);
or U11412 (N_11412,N_10262,N_10997);
nor U11413 (N_11413,N_10704,N_10189);
and U11414 (N_11414,N_10160,N_10217);
and U11415 (N_11415,N_10555,N_10264);
or U11416 (N_11416,N_10564,N_10934);
xor U11417 (N_11417,N_10387,N_11122);
nor U11418 (N_11418,N_10888,N_10712);
or U11419 (N_11419,N_10443,N_10027);
and U11420 (N_11420,N_10376,N_10137);
xor U11421 (N_11421,N_11205,N_10198);
nand U11422 (N_11422,N_11110,N_10756);
nor U11423 (N_11423,N_10306,N_10411);
xor U11424 (N_11424,N_10840,N_10452);
nor U11425 (N_11425,N_10959,N_10297);
nor U11426 (N_11426,N_10843,N_10597);
or U11427 (N_11427,N_10599,N_10081);
nand U11428 (N_11428,N_10078,N_10875);
and U11429 (N_11429,N_10851,N_10886);
and U11430 (N_11430,N_10790,N_10408);
and U11431 (N_11431,N_10059,N_10395);
and U11432 (N_11432,N_10673,N_10289);
or U11433 (N_11433,N_10521,N_10652);
or U11434 (N_11434,N_10808,N_10055);
xor U11435 (N_11435,N_10796,N_10006);
and U11436 (N_11436,N_10726,N_11092);
nor U11437 (N_11437,N_10345,N_10601);
xnor U11438 (N_11438,N_10688,N_11219);
and U11439 (N_11439,N_10556,N_10751);
and U11440 (N_11440,N_10779,N_10770);
and U11441 (N_11441,N_10070,N_10169);
nor U11442 (N_11442,N_10407,N_10431);
nor U11443 (N_11443,N_10187,N_11103);
nand U11444 (N_11444,N_10709,N_10212);
and U11445 (N_11445,N_10692,N_10681);
and U11446 (N_11446,N_10120,N_10908);
nand U11447 (N_11447,N_10177,N_10374);
and U11448 (N_11448,N_10486,N_10532);
xor U11449 (N_11449,N_10530,N_10806);
and U11450 (N_11450,N_10739,N_10533);
xor U11451 (N_11451,N_10781,N_10483);
nand U11452 (N_11452,N_10000,N_10661);
or U11453 (N_11453,N_10035,N_10523);
nand U11454 (N_11454,N_10740,N_10361);
nor U11455 (N_11455,N_10741,N_10129);
or U11456 (N_11456,N_10858,N_11191);
nand U11457 (N_11457,N_10920,N_10960);
nor U11458 (N_11458,N_10388,N_10967);
xor U11459 (N_11459,N_11154,N_10102);
and U11460 (N_11460,N_11068,N_11134);
nand U11461 (N_11461,N_11178,N_10175);
and U11462 (N_11462,N_10363,N_10980);
and U11463 (N_11463,N_10789,N_10864);
xnor U11464 (N_11464,N_10984,N_10855);
nor U11465 (N_11465,N_10020,N_10266);
and U11466 (N_11466,N_10230,N_10735);
nand U11467 (N_11467,N_10707,N_10396);
nor U11468 (N_11468,N_11158,N_10504);
and U11469 (N_11469,N_10165,N_10827);
nor U11470 (N_11470,N_10668,N_10616);
xnor U11471 (N_11471,N_11169,N_10052);
or U11472 (N_11472,N_11000,N_10417);
and U11473 (N_11473,N_10272,N_10593);
nand U11474 (N_11474,N_11069,N_11231);
nand U11475 (N_11475,N_10519,N_11030);
nor U11476 (N_11476,N_10446,N_10185);
or U11477 (N_11477,N_10260,N_10008);
and U11478 (N_11478,N_10355,N_10797);
xnor U11479 (N_11479,N_10336,N_10744);
nand U11480 (N_11480,N_10693,N_10595);
xnor U11481 (N_11481,N_10339,N_10897);
nor U11482 (N_11482,N_11140,N_10398);
and U11483 (N_11483,N_10611,N_10981);
xor U11484 (N_11484,N_10553,N_11065);
nand U11485 (N_11485,N_10627,N_10507);
xnor U11486 (N_11486,N_11081,N_10566);
xor U11487 (N_11487,N_10846,N_10461);
xnor U11488 (N_11488,N_10977,N_10913);
xnor U11489 (N_11489,N_10303,N_11227);
and U11490 (N_11490,N_10916,N_10853);
nor U11491 (N_11491,N_11009,N_10725);
nor U11492 (N_11492,N_10280,N_10460);
and U11493 (N_11493,N_11116,N_10286);
and U11494 (N_11494,N_10656,N_10852);
nand U11495 (N_11495,N_11034,N_10085);
nand U11496 (N_11496,N_10308,N_10349);
xor U11497 (N_11497,N_10222,N_11097);
nor U11498 (N_11498,N_11173,N_10662);
or U11499 (N_11499,N_10878,N_10733);
xnor U11500 (N_11500,N_10768,N_10615);
and U11501 (N_11501,N_10623,N_10646);
nor U11502 (N_11502,N_10038,N_10294);
xor U11503 (N_11503,N_10524,N_10067);
and U11504 (N_11504,N_10151,N_10378);
xnor U11505 (N_11505,N_10089,N_10769);
and U11506 (N_11506,N_10456,N_10659);
or U11507 (N_11507,N_10414,N_10713);
xor U11508 (N_11508,N_10991,N_10863);
nor U11509 (N_11509,N_11126,N_10604);
or U11510 (N_11510,N_10690,N_10022);
or U11511 (N_11511,N_10869,N_10766);
nor U11512 (N_11512,N_10003,N_11003);
nor U11513 (N_11513,N_10678,N_10978);
nand U11514 (N_11514,N_10077,N_11241);
xor U11515 (N_11515,N_10651,N_10973);
nand U11516 (N_11516,N_10674,N_10928);
xor U11517 (N_11517,N_10053,N_10503);
nand U11518 (N_11518,N_10621,N_10112);
and U11519 (N_11519,N_10760,N_10773);
and U11520 (N_11520,N_10861,N_10647);
or U11521 (N_11521,N_10451,N_10467);
xor U11522 (N_11522,N_10107,N_10665);
or U11523 (N_11523,N_10103,N_10682);
nor U11524 (N_11524,N_10807,N_10191);
nor U11525 (N_11525,N_10710,N_10637);
xor U11526 (N_11526,N_10918,N_10605);
xor U11527 (N_11527,N_10743,N_11041);
or U11528 (N_11528,N_10313,N_11224);
and U11529 (N_11529,N_10700,N_11166);
nor U11530 (N_11530,N_10500,N_11063);
and U11531 (N_11531,N_10866,N_10847);
xor U11532 (N_11532,N_10584,N_10485);
and U11533 (N_11533,N_10590,N_10628);
nand U11534 (N_11534,N_10111,N_10557);
and U11535 (N_11535,N_10021,N_11236);
nand U11536 (N_11536,N_10088,N_10814);
nand U11537 (N_11537,N_10818,N_10675);
xnor U11538 (N_11538,N_10976,N_10318);
xnor U11539 (N_11539,N_10292,N_10749);
and U11540 (N_11540,N_10269,N_10755);
xor U11541 (N_11541,N_10450,N_11017);
xor U11542 (N_11542,N_10571,N_10882);
nand U11543 (N_11543,N_10481,N_10203);
nand U11544 (N_11544,N_10168,N_11028);
or U11545 (N_11545,N_10424,N_11032);
nor U11546 (N_11546,N_10104,N_11147);
nand U11547 (N_11547,N_10454,N_11101);
or U11548 (N_11548,N_10598,N_11006);
and U11549 (N_11549,N_10158,N_10299);
nor U11550 (N_11550,N_10951,N_10057);
nor U11551 (N_11551,N_10377,N_10351);
nor U11552 (N_11552,N_10066,N_10254);
or U11553 (N_11553,N_10236,N_10835);
and U11554 (N_11554,N_10772,N_11073);
and U11555 (N_11555,N_10892,N_10525);
nor U11556 (N_11556,N_10909,N_11083);
or U11557 (N_11557,N_10542,N_10550);
nor U11558 (N_11558,N_11232,N_11076);
nand U11559 (N_11559,N_10974,N_10826);
nand U11560 (N_11560,N_10065,N_10498);
xnor U11561 (N_11561,N_10792,N_10543);
and U11562 (N_11562,N_10798,N_10242);
or U11563 (N_11563,N_11179,N_11192);
xnor U11564 (N_11564,N_10380,N_10670);
nand U11565 (N_11565,N_11023,N_10170);
nand U11566 (N_11566,N_10270,N_10547);
and U11567 (N_11567,N_11168,N_10037);
and U11568 (N_11568,N_10285,N_10653);
and U11569 (N_11569,N_10150,N_10990);
or U11570 (N_11570,N_10581,N_11156);
or U11571 (N_11571,N_11213,N_10375);
and U11572 (N_11572,N_10091,N_10310);
nor U11573 (N_11573,N_10680,N_10697);
xor U11574 (N_11574,N_10196,N_10453);
nand U11575 (N_11575,N_10401,N_10634);
and U11576 (N_11576,N_10830,N_10333);
xor U11577 (N_11577,N_10572,N_11094);
xor U11578 (N_11578,N_10250,N_10816);
xor U11579 (N_11579,N_10534,N_10592);
or U11580 (N_11580,N_11136,N_11113);
nand U11581 (N_11581,N_11026,N_10246);
nand U11582 (N_11582,N_10209,N_11207);
xnor U11583 (N_11583,N_10092,N_10152);
nand U11584 (N_11584,N_10049,N_10786);
nor U11585 (N_11585,N_10135,N_11215);
and U11586 (N_11586,N_10753,N_10905);
nor U11587 (N_11587,N_11238,N_10018);
xnor U11588 (N_11588,N_10418,N_11242);
and U11589 (N_11589,N_11060,N_10667);
or U11590 (N_11590,N_10420,N_10267);
nor U11591 (N_11591,N_11188,N_10128);
nand U11592 (N_11592,N_10635,N_10428);
xor U11593 (N_11593,N_10334,N_10352);
or U11594 (N_11594,N_10708,N_10949);
nand U11595 (N_11595,N_11004,N_10914);
nor U11596 (N_11596,N_10366,N_10536);
and U11597 (N_11597,N_10223,N_10323);
nand U11598 (N_11598,N_10494,N_11049);
nor U11599 (N_11599,N_11061,N_10650);
nand U11600 (N_11600,N_10362,N_10441);
and U11601 (N_11601,N_10327,N_10501);
and U11602 (N_11602,N_10989,N_10703);
and U11603 (N_11603,N_11216,N_10162);
or U11604 (N_11604,N_10455,N_10569);
nor U11605 (N_11605,N_10492,N_10221);
and U11606 (N_11606,N_10698,N_10591);
or U11607 (N_11607,N_10421,N_10365);
xnor U11608 (N_11608,N_10679,N_10983);
xor U11609 (N_11609,N_10007,N_10586);
nor U11610 (N_11610,N_11189,N_11052);
nand U11611 (N_11611,N_10074,N_10412);
or U11612 (N_11612,N_11108,N_10884);
or U11613 (N_11613,N_10064,N_10608);
and U11614 (N_11614,N_10510,N_10810);
nand U11615 (N_11615,N_10484,N_10098);
xor U11616 (N_11616,N_10626,N_10923);
or U11617 (N_11617,N_11047,N_10499);
nor U11618 (N_11618,N_10048,N_11141);
nor U11619 (N_11619,N_10423,N_10876);
or U11620 (N_11620,N_10669,N_10338);
nor U11621 (N_11621,N_11208,N_10400);
xnor U11622 (N_11622,N_10060,N_11163);
or U11623 (N_11623,N_11161,N_10839);
or U11624 (N_11624,N_11214,N_11074);
and U11625 (N_11625,N_10243,N_10463);
and U11626 (N_11626,N_10714,N_10642);
nand U11627 (N_11627,N_10340,N_10887);
nor U11628 (N_11628,N_11039,N_10956);
nor U11629 (N_11629,N_10273,N_10942);
and U11630 (N_11630,N_11139,N_10537);
nand U11631 (N_11631,N_11019,N_10330);
nor U11632 (N_11632,N_10945,N_11233);
nand U11633 (N_11633,N_10794,N_10513);
nand U11634 (N_11634,N_10829,N_10033);
and U11635 (N_11635,N_10144,N_10529);
and U11636 (N_11636,N_10208,N_10051);
nand U11637 (N_11637,N_10181,N_10047);
or U11638 (N_11638,N_11230,N_11012);
nor U11639 (N_11639,N_10907,N_10265);
or U11640 (N_11640,N_10385,N_10383);
nor U11641 (N_11641,N_10153,N_10211);
xnor U11642 (N_11642,N_11165,N_10231);
nor U11643 (N_11643,N_10613,N_10393);
nor U11644 (N_11644,N_10791,N_10574);
and U11645 (N_11645,N_11057,N_10275);
and U11646 (N_11646,N_10040,N_10822);
nand U11647 (N_11647,N_10950,N_10036);
xor U11648 (N_11648,N_10192,N_11194);
nor U11649 (N_11649,N_11239,N_10497);
or U11650 (N_11650,N_10900,N_10281);
nor U11651 (N_11651,N_10577,N_10277);
and U11652 (N_11652,N_10364,N_10319);
nor U11653 (N_11653,N_10477,N_10083);
nor U11654 (N_11654,N_10392,N_10891);
xor U11655 (N_11655,N_10554,N_11064);
nand U11656 (N_11656,N_10516,N_10214);
or U11657 (N_11657,N_10465,N_10284);
nor U11658 (N_11658,N_10687,N_11050);
nand U11659 (N_11659,N_10031,N_10630);
xnor U11660 (N_11660,N_10367,N_10329);
xor U11661 (N_11661,N_10664,N_10930);
and U11662 (N_11662,N_10655,N_10938);
or U11663 (N_11663,N_10619,N_10141);
or U11664 (N_11664,N_10617,N_10343);
or U11665 (N_11665,N_11226,N_10992);
nand U11666 (N_11666,N_10307,N_10941);
nor U11667 (N_11667,N_11029,N_10813);
or U11668 (N_11668,N_10233,N_10856);
and U11669 (N_11669,N_10495,N_10032);
nand U11670 (N_11670,N_11202,N_11105);
and U11671 (N_11671,N_10326,N_10134);
or U11672 (N_11672,N_10278,N_10885);
and U11673 (N_11673,N_11067,N_10042);
xor U11674 (N_11674,N_10197,N_10082);
or U11675 (N_11675,N_10787,N_10506);
nor U11676 (N_11676,N_10283,N_10445);
nand U11677 (N_11677,N_10341,N_10654);
nor U11678 (N_11678,N_10904,N_10775);
xnor U11679 (N_11679,N_10259,N_10315);
and U11680 (N_11680,N_10317,N_11127);
or U11681 (N_11681,N_10127,N_11091);
nand U11682 (N_11682,N_11171,N_10010);
xor U11683 (N_11683,N_11221,N_10780);
nor U11684 (N_11684,N_10895,N_10063);
nor U11685 (N_11685,N_10935,N_10582);
or U11686 (N_11686,N_10184,N_10765);
and U11687 (N_11687,N_10011,N_11031);
nor U11688 (N_11688,N_11077,N_10520);
nor U11689 (N_11689,N_10881,N_10867);
nor U11690 (N_11690,N_11170,N_11225);
and U11691 (N_11691,N_10471,N_10799);
or U11692 (N_11692,N_10419,N_10328);
nand U11693 (N_11693,N_10953,N_10291);
xnor U11694 (N_11694,N_10695,N_10763);
nor U11695 (N_11695,N_10580,N_10924);
or U11696 (N_11696,N_10701,N_11043);
nor U11697 (N_11697,N_10545,N_11120);
or U11698 (N_11698,N_10138,N_10369);
and U11699 (N_11699,N_10029,N_11059);
xor U11700 (N_11700,N_10017,N_10225);
nor U11701 (N_11701,N_10076,N_11181);
and U11702 (N_11702,N_10815,N_10106);
nand U11703 (N_11703,N_10394,N_11144);
nand U11704 (N_11704,N_10879,N_11093);
nor U11705 (N_11705,N_11167,N_10841);
xnor U11706 (N_11706,N_10754,N_10844);
nand U11707 (N_11707,N_10995,N_10084);
xnor U11708 (N_11708,N_11164,N_10579);
nand U11709 (N_11709,N_10488,N_11249);
nor U11710 (N_11710,N_10148,N_11095);
nor U11711 (N_11711,N_10736,N_11125);
nand U11712 (N_11712,N_10346,N_10583);
or U11713 (N_11713,N_10404,N_10472);
xnor U11714 (N_11714,N_10300,N_10320);
xor U11715 (N_11715,N_10350,N_10722);
nand U11716 (N_11716,N_10186,N_10603);
nor U11717 (N_11717,N_10738,N_10309);
nand U11718 (N_11718,N_10447,N_10585);
nor U11719 (N_11719,N_10548,N_11100);
xnor U11720 (N_11720,N_10849,N_10573);
or U11721 (N_11721,N_11078,N_10894);
or U11722 (N_11722,N_10331,N_10531);
or U11723 (N_11723,N_11022,N_11090);
and U11724 (N_11724,N_11129,N_11045);
xnor U11725 (N_11725,N_10563,N_10649);
nor U11726 (N_11726,N_10025,N_10199);
or U11727 (N_11727,N_10238,N_10963);
or U11728 (N_11728,N_10464,N_10831);
and U11729 (N_11729,N_10288,N_10902);
and U11730 (N_11730,N_10828,N_10193);
or U11731 (N_11731,N_10720,N_10859);
nand U11732 (N_11732,N_10587,N_10073);
nand U11733 (N_11733,N_11121,N_11044);
nor U11734 (N_11734,N_10099,N_10939);
nor U11735 (N_11735,N_10544,N_11143);
nand U11736 (N_11736,N_10927,N_10561);
nor U11737 (N_11737,N_10730,N_11027);
and U11738 (N_11738,N_10382,N_10785);
and U11739 (N_11739,N_10079,N_11058);
nor U11740 (N_11740,N_11223,N_11220);
and U11741 (N_11741,N_10101,N_11211);
and U11742 (N_11742,N_10734,N_10508);
and U11743 (N_11743,N_10324,N_10724);
and U11744 (N_11744,N_11185,N_11132);
nor U11745 (N_11745,N_10696,N_10596);
nand U11746 (N_11746,N_10229,N_10527);
xor U11747 (N_11747,N_10009,N_10133);
xor U11748 (N_11748,N_11106,N_10457);
or U11749 (N_11749,N_10268,N_10139);
nor U11750 (N_11750,N_11048,N_10898);
nor U11751 (N_11751,N_10496,N_10683);
nand U11752 (N_11752,N_10825,N_10552);
nor U11753 (N_11753,N_10105,N_11036);
xor U11754 (N_11754,N_10788,N_10301);
nand U11755 (N_11755,N_10748,N_10360);
or U11756 (N_11756,N_10216,N_11082);
or U11757 (N_11757,N_10200,N_10889);
nor U11758 (N_11758,N_10784,N_10295);
or U11759 (N_11759,N_10948,N_11109);
nand U11760 (N_11760,N_11177,N_10368);
nand U11761 (N_11761,N_10706,N_10771);
or U11762 (N_11762,N_10426,N_11195);
or U11763 (N_11763,N_10204,N_10893);
or U11764 (N_11764,N_10776,N_10210);
xor U11765 (N_11765,N_10166,N_10711);
nand U11766 (N_11766,N_10922,N_10140);
or U11767 (N_11767,N_10994,N_10244);
or U11768 (N_11768,N_10332,N_10834);
or U11769 (N_11769,N_10868,N_10919);
or U11770 (N_11770,N_10715,N_10253);
nand U11771 (N_11771,N_10390,N_10782);
xor U11772 (N_11772,N_10094,N_11199);
xor U11773 (N_11773,N_10397,N_10296);
xor U11774 (N_11774,N_10458,N_10227);
and U11775 (N_11775,N_11128,N_10234);
and U11776 (N_11776,N_10190,N_10183);
nand U11777 (N_11777,N_10194,N_10969);
xnor U11778 (N_11778,N_11196,N_10257);
nor U11779 (N_11779,N_10416,N_10205);
nand U11780 (N_11780,N_10625,N_11013);
nor U11781 (N_11781,N_10921,N_11187);
nor U11782 (N_11782,N_10685,N_10069);
nor U11783 (N_11783,N_10946,N_10817);
xor U11784 (N_11784,N_10618,N_10019);
xnor U11785 (N_11785,N_10549,N_10824);
nor U11786 (N_11786,N_11206,N_10086);
nor U11787 (N_11787,N_10386,N_11153);
nand U11788 (N_11788,N_11186,N_10087);
nand U11789 (N_11789,N_11118,N_11209);
xnor U11790 (N_11790,N_11014,N_10474);
nor U11791 (N_11791,N_10570,N_11040);
nor U11792 (N_11792,N_10258,N_11119);
and U11793 (N_11793,N_11114,N_11157);
nand U11794 (N_11794,N_10436,N_10116);
xor U11795 (N_11795,N_10877,N_11015);
and U11796 (N_11796,N_10528,N_10444);
or U11797 (N_11797,N_10171,N_10468);
or U11798 (N_11798,N_10546,N_10015);
nand U11799 (N_11799,N_10068,N_11117);
nand U11800 (N_11800,N_10640,N_10462);
or U11801 (N_11801,N_10061,N_11204);
nand U11802 (N_11802,N_11183,N_10435);
nand U11803 (N_11803,N_10837,N_11243);
nor U11804 (N_11804,N_10342,N_10213);
and U11805 (N_11805,N_10293,N_11228);
xnor U11806 (N_11806,N_10639,N_10370);
and U11807 (N_11807,N_10541,N_10026);
nand U11808 (N_11808,N_10911,N_10433);
and U11809 (N_11809,N_10130,N_10002);
nand U11810 (N_11810,N_10915,N_10820);
nand U11811 (N_11811,N_10097,N_10777);
nand U11812 (N_11812,N_10823,N_11237);
or U11813 (N_11813,N_10551,N_10476);
nand U11814 (N_11814,N_11235,N_10964);
or U11815 (N_11815,N_10271,N_10721);
nor U11816 (N_11816,N_10663,N_10201);
and U11817 (N_11817,N_10480,N_10434);
and U11818 (N_11818,N_10108,N_10256);
nand U11819 (N_11819,N_11222,N_10578);
or U11820 (N_11820,N_10998,N_11085);
or U11821 (N_11821,N_10034,N_10644);
nor U11822 (N_11822,N_10538,N_10427);
nand U11823 (N_11823,N_10173,N_10727);
nor U11824 (N_11824,N_10425,N_10358);
and U11825 (N_11825,N_10783,N_10750);
and U11826 (N_11826,N_10142,N_11001);
nor U11827 (N_11827,N_10747,N_10188);
nor U11828 (N_11828,N_10558,N_11005);
nor U11829 (N_11829,N_10641,N_10629);
and U11830 (N_11830,N_10793,N_10469);
xor U11831 (N_11831,N_10660,N_10804);
nor U11832 (N_11832,N_10145,N_11062);
or U11833 (N_11833,N_10975,N_10249);
and U11834 (N_11834,N_10801,N_11240);
or U11835 (N_11835,N_11159,N_10971);
nand U11836 (N_11836,N_11130,N_11107);
nor U11837 (N_11837,N_10874,N_10039);
nor U11838 (N_11838,N_10432,N_10100);
and U11839 (N_11839,N_10731,N_11145);
nor U11840 (N_11840,N_10304,N_10833);
or U11841 (N_11841,N_10631,N_10415);
xnor U11842 (N_11842,N_10248,N_10505);
xnor U11843 (N_11843,N_10767,N_10896);
and U11844 (N_11844,N_10576,N_10873);
nor U11845 (N_11845,N_10305,N_10759);
nor U11846 (N_11846,N_10872,N_10056);
or U11847 (N_11847,N_11020,N_11138);
nand U11848 (N_11848,N_11080,N_10917);
nor U11849 (N_11849,N_10737,N_11218);
nor U11850 (N_11850,N_10689,N_11245);
nor U11851 (N_11851,N_11160,N_10156);
nand U11852 (N_11852,N_10686,N_11102);
xor U11853 (N_11853,N_10235,N_10132);
nor U11854 (N_11854,N_10195,N_11148);
nand U11855 (N_11855,N_11193,N_10671);
or U11856 (N_11856,N_11124,N_10075);
and U11857 (N_11857,N_10095,N_10218);
and U11858 (N_11858,N_10430,N_11155);
or U11859 (N_11859,N_10124,N_10043);
nor U11860 (N_11860,N_11151,N_10028);
and U11861 (N_11861,N_10600,N_10691);
xor U11862 (N_11862,N_10575,N_10490);
or U11863 (N_11863,N_10509,N_10812);
and U11864 (N_11864,N_10054,N_11172);
nand U11865 (N_11865,N_10614,N_10440);
xnor U11866 (N_11866,N_10050,N_10016);
nor U11867 (N_11867,N_10883,N_10954);
nand U11868 (N_11868,N_10926,N_10517);
or U11869 (N_11869,N_10422,N_11054);
xor U11870 (N_11870,N_10058,N_10282);
or U11871 (N_11871,N_10096,N_10442);
or U11872 (N_11872,N_10228,N_10943);
or U11873 (N_11873,N_10117,N_10518);
and U11874 (N_11874,N_11201,N_10154);
nor U11875 (N_11875,N_11031,N_10919);
and U11876 (N_11876,N_11112,N_10295);
nand U11877 (N_11877,N_10201,N_10980);
nand U11878 (N_11878,N_10958,N_10530);
or U11879 (N_11879,N_11224,N_10119);
or U11880 (N_11880,N_10990,N_11136);
or U11881 (N_11881,N_10609,N_10519);
or U11882 (N_11882,N_10315,N_10399);
nor U11883 (N_11883,N_10634,N_10166);
nor U11884 (N_11884,N_10495,N_11103);
nand U11885 (N_11885,N_10396,N_10299);
and U11886 (N_11886,N_10769,N_11016);
nor U11887 (N_11887,N_11087,N_10838);
or U11888 (N_11888,N_10132,N_10518);
xnor U11889 (N_11889,N_10712,N_10379);
nand U11890 (N_11890,N_10764,N_10342);
nand U11891 (N_11891,N_10815,N_10530);
nor U11892 (N_11892,N_10375,N_10765);
xor U11893 (N_11893,N_10264,N_11147);
nand U11894 (N_11894,N_11112,N_10754);
nor U11895 (N_11895,N_10667,N_10019);
nor U11896 (N_11896,N_10083,N_11134);
and U11897 (N_11897,N_10698,N_11081);
xnor U11898 (N_11898,N_11199,N_10526);
or U11899 (N_11899,N_10549,N_10490);
or U11900 (N_11900,N_10703,N_10248);
nor U11901 (N_11901,N_10540,N_10630);
or U11902 (N_11902,N_10967,N_11131);
nand U11903 (N_11903,N_11132,N_10547);
nand U11904 (N_11904,N_10356,N_10559);
nand U11905 (N_11905,N_10809,N_10430);
nand U11906 (N_11906,N_11020,N_10336);
nand U11907 (N_11907,N_10391,N_10107);
xnor U11908 (N_11908,N_10669,N_10152);
or U11909 (N_11909,N_10013,N_10185);
and U11910 (N_11910,N_10956,N_10633);
nand U11911 (N_11911,N_10200,N_11124);
xnor U11912 (N_11912,N_10660,N_11099);
nor U11913 (N_11913,N_10655,N_11017);
or U11914 (N_11914,N_10126,N_10639);
xor U11915 (N_11915,N_10968,N_11249);
nand U11916 (N_11916,N_10650,N_10223);
or U11917 (N_11917,N_10712,N_11062);
and U11918 (N_11918,N_10911,N_10587);
or U11919 (N_11919,N_10773,N_11081);
nand U11920 (N_11920,N_10777,N_10955);
nor U11921 (N_11921,N_10096,N_10422);
nand U11922 (N_11922,N_10552,N_10056);
or U11923 (N_11923,N_10068,N_11144);
nand U11924 (N_11924,N_10611,N_10578);
and U11925 (N_11925,N_10244,N_10888);
xnor U11926 (N_11926,N_10527,N_10969);
nand U11927 (N_11927,N_10810,N_11016);
and U11928 (N_11928,N_10301,N_10911);
and U11929 (N_11929,N_10206,N_11195);
and U11930 (N_11930,N_10602,N_11085);
nor U11931 (N_11931,N_10560,N_10378);
and U11932 (N_11932,N_11234,N_11154);
nand U11933 (N_11933,N_10157,N_10140);
and U11934 (N_11934,N_10119,N_10832);
and U11935 (N_11935,N_10261,N_10075);
xor U11936 (N_11936,N_10799,N_11225);
nor U11937 (N_11937,N_10883,N_10536);
and U11938 (N_11938,N_11139,N_10100);
xnor U11939 (N_11939,N_10336,N_10212);
and U11940 (N_11940,N_11222,N_10690);
and U11941 (N_11941,N_10419,N_11095);
or U11942 (N_11942,N_10382,N_10304);
xor U11943 (N_11943,N_11234,N_11212);
xor U11944 (N_11944,N_10280,N_10143);
nor U11945 (N_11945,N_10363,N_11128);
or U11946 (N_11946,N_10578,N_10547);
and U11947 (N_11947,N_10210,N_10174);
xnor U11948 (N_11948,N_10463,N_10598);
nor U11949 (N_11949,N_11068,N_11217);
xnor U11950 (N_11950,N_10032,N_10566);
and U11951 (N_11951,N_10558,N_10857);
and U11952 (N_11952,N_10810,N_11160);
xnor U11953 (N_11953,N_10674,N_10469);
xnor U11954 (N_11954,N_10233,N_11155);
or U11955 (N_11955,N_10487,N_10416);
or U11956 (N_11956,N_11057,N_10656);
nor U11957 (N_11957,N_10917,N_10676);
and U11958 (N_11958,N_10315,N_10988);
or U11959 (N_11959,N_10274,N_10870);
or U11960 (N_11960,N_10790,N_10592);
or U11961 (N_11961,N_10145,N_10993);
nor U11962 (N_11962,N_10512,N_10955);
nor U11963 (N_11963,N_10635,N_10446);
or U11964 (N_11964,N_11218,N_11165);
or U11965 (N_11965,N_10180,N_10791);
nand U11966 (N_11966,N_10462,N_10220);
xor U11967 (N_11967,N_10602,N_10026);
nand U11968 (N_11968,N_11121,N_11230);
xor U11969 (N_11969,N_10750,N_10463);
or U11970 (N_11970,N_10974,N_10135);
xor U11971 (N_11971,N_10603,N_10657);
nor U11972 (N_11972,N_10175,N_10599);
or U11973 (N_11973,N_10677,N_10840);
nor U11974 (N_11974,N_10918,N_10513);
or U11975 (N_11975,N_10840,N_10790);
nand U11976 (N_11976,N_10899,N_10961);
xor U11977 (N_11977,N_10086,N_11209);
nor U11978 (N_11978,N_10095,N_10421);
or U11979 (N_11979,N_10072,N_11242);
nor U11980 (N_11980,N_10639,N_11093);
and U11981 (N_11981,N_10747,N_11048);
and U11982 (N_11982,N_10723,N_11244);
nand U11983 (N_11983,N_11245,N_10575);
xnor U11984 (N_11984,N_10166,N_10545);
xor U11985 (N_11985,N_10401,N_10879);
or U11986 (N_11986,N_10311,N_10836);
or U11987 (N_11987,N_10858,N_10848);
nor U11988 (N_11988,N_11028,N_11119);
and U11989 (N_11989,N_10747,N_10221);
or U11990 (N_11990,N_11083,N_10098);
nand U11991 (N_11991,N_10172,N_10215);
nor U11992 (N_11992,N_11107,N_10784);
nor U11993 (N_11993,N_10035,N_11077);
and U11994 (N_11994,N_10377,N_10639);
nand U11995 (N_11995,N_10004,N_10069);
or U11996 (N_11996,N_10187,N_10878);
nor U11997 (N_11997,N_10736,N_11206);
nor U11998 (N_11998,N_10462,N_11219);
nand U11999 (N_11999,N_11153,N_10544);
nor U12000 (N_12000,N_10265,N_10262);
nor U12001 (N_12001,N_10614,N_11007);
nand U12002 (N_12002,N_10933,N_11101);
xnor U12003 (N_12003,N_10588,N_10600);
and U12004 (N_12004,N_10520,N_10240);
xor U12005 (N_12005,N_10398,N_10285);
or U12006 (N_12006,N_10732,N_10677);
or U12007 (N_12007,N_10399,N_11086);
nand U12008 (N_12008,N_10747,N_10362);
or U12009 (N_12009,N_10996,N_11088);
xnor U12010 (N_12010,N_10347,N_10381);
nor U12011 (N_12011,N_11198,N_11189);
and U12012 (N_12012,N_10323,N_11122);
xnor U12013 (N_12013,N_11212,N_11142);
nor U12014 (N_12014,N_10522,N_10396);
xnor U12015 (N_12015,N_10263,N_10001);
or U12016 (N_12016,N_10060,N_10064);
nor U12017 (N_12017,N_10596,N_11216);
nor U12018 (N_12018,N_10680,N_10595);
xor U12019 (N_12019,N_10819,N_10027);
xnor U12020 (N_12020,N_10005,N_10014);
nand U12021 (N_12021,N_10361,N_10928);
xnor U12022 (N_12022,N_11217,N_10340);
or U12023 (N_12023,N_10405,N_10408);
xor U12024 (N_12024,N_11043,N_10181);
and U12025 (N_12025,N_11025,N_10032);
nor U12026 (N_12026,N_10377,N_11135);
xor U12027 (N_12027,N_10197,N_11152);
or U12028 (N_12028,N_10493,N_10078);
or U12029 (N_12029,N_11210,N_10367);
nor U12030 (N_12030,N_10683,N_10582);
or U12031 (N_12031,N_10998,N_10440);
and U12032 (N_12032,N_11056,N_10617);
xor U12033 (N_12033,N_11082,N_10096);
and U12034 (N_12034,N_10996,N_11100);
and U12035 (N_12035,N_10779,N_10698);
nor U12036 (N_12036,N_11198,N_10215);
or U12037 (N_12037,N_10937,N_10541);
xor U12038 (N_12038,N_10146,N_11157);
and U12039 (N_12039,N_10949,N_10463);
or U12040 (N_12040,N_10301,N_10971);
xnor U12041 (N_12041,N_10467,N_10684);
and U12042 (N_12042,N_10401,N_11183);
and U12043 (N_12043,N_11058,N_11120);
xor U12044 (N_12044,N_10525,N_10294);
nor U12045 (N_12045,N_10094,N_10334);
nand U12046 (N_12046,N_10502,N_11102);
xor U12047 (N_12047,N_10889,N_10699);
nor U12048 (N_12048,N_11073,N_10380);
nand U12049 (N_12049,N_10980,N_10173);
xnor U12050 (N_12050,N_10901,N_10836);
or U12051 (N_12051,N_10908,N_10720);
or U12052 (N_12052,N_10840,N_10612);
or U12053 (N_12053,N_10215,N_10529);
or U12054 (N_12054,N_10808,N_10643);
and U12055 (N_12055,N_10014,N_11025);
nand U12056 (N_12056,N_10026,N_11101);
xnor U12057 (N_12057,N_10701,N_11071);
nor U12058 (N_12058,N_10336,N_10136);
nand U12059 (N_12059,N_10641,N_10154);
nor U12060 (N_12060,N_10166,N_10371);
nor U12061 (N_12061,N_10390,N_10548);
and U12062 (N_12062,N_10283,N_11248);
or U12063 (N_12063,N_11219,N_10584);
nor U12064 (N_12064,N_10062,N_10443);
nand U12065 (N_12065,N_11226,N_10430);
xor U12066 (N_12066,N_10092,N_10056);
xnor U12067 (N_12067,N_10903,N_10587);
nor U12068 (N_12068,N_11103,N_10909);
and U12069 (N_12069,N_10022,N_10441);
xnor U12070 (N_12070,N_10296,N_10630);
and U12071 (N_12071,N_11207,N_10219);
xor U12072 (N_12072,N_10114,N_11184);
xor U12073 (N_12073,N_10974,N_10079);
nand U12074 (N_12074,N_10466,N_10126);
nor U12075 (N_12075,N_10834,N_10206);
nand U12076 (N_12076,N_10304,N_10256);
xor U12077 (N_12077,N_10794,N_10408);
xor U12078 (N_12078,N_10674,N_10611);
nand U12079 (N_12079,N_10878,N_10969);
nand U12080 (N_12080,N_10436,N_10795);
or U12081 (N_12081,N_10094,N_10474);
and U12082 (N_12082,N_10453,N_10525);
nand U12083 (N_12083,N_11240,N_10901);
nor U12084 (N_12084,N_11079,N_10011);
xnor U12085 (N_12085,N_10564,N_10029);
xor U12086 (N_12086,N_10339,N_10595);
or U12087 (N_12087,N_10658,N_11236);
and U12088 (N_12088,N_10123,N_10782);
nor U12089 (N_12089,N_10839,N_11129);
or U12090 (N_12090,N_10672,N_10955);
nand U12091 (N_12091,N_10896,N_10477);
or U12092 (N_12092,N_10088,N_10395);
xor U12093 (N_12093,N_10175,N_11081);
and U12094 (N_12094,N_10635,N_10376);
nor U12095 (N_12095,N_10459,N_10910);
nor U12096 (N_12096,N_10694,N_10375);
or U12097 (N_12097,N_10553,N_10653);
nand U12098 (N_12098,N_10140,N_10960);
nand U12099 (N_12099,N_10706,N_10638);
nand U12100 (N_12100,N_10631,N_10715);
or U12101 (N_12101,N_10472,N_10478);
xor U12102 (N_12102,N_10958,N_10344);
xor U12103 (N_12103,N_11120,N_11104);
and U12104 (N_12104,N_10512,N_10338);
nor U12105 (N_12105,N_10927,N_11222);
and U12106 (N_12106,N_11070,N_11078);
nor U12107 (N_12107,N_10606,N_10510);
xor U12108 (N_12108,N_10296,N_11064);
and U12109 (N_12109,N_10555,N_10463);
and U12110 (N_12110,N_10432,N_10083);
nand U12111 (N_12111,N_11095,N_10754);
or U12112 (N_12112,N_10410,N_10276);
and U12113 (N_12113,N_11166,N_10986);
or U12114 (N_12114,N_10657,N_11055);
nor U12115 (N_12115,N_10552,N_10982);
and U12116 (N_12116,N_10765,N_10426);
xor U12117 (N_12117,N_10568,N_10591);
nor U12118 (N_12118,N_10055,N_11077);
or U12119 (N_12119,N_10293,N_10377);
nor U12120 (N_12120,N_10532,N_10469);
nor U12121 (N_12121,N_10752,N_10424);
nand U12122 (N_12122,N_10965,N_10686);
nor U12123 (N_12123,N_11174,N_10758);
xor U12124 (N_12124,N_11150,N_10948);
xor U12125 (N_12125,N_10353,N_10957);
nand U12126 (N_12126,N_10054,N_10011);
xnor U12127 (N_12127,N_11125,N_10068);
or U12128 (N_12128,N_10448,N_11047);
or U12129 (N_12129,N_10100,N_11176);
xnor U12130 (N_12130,N_11113,N_10788);
nand U12131 (N_12131,N_10471,N_10086);
and U12132 (N_12132,N_10066,N_10164);
xor U12133 (N_12133,N_10298,N_11095);
xnor U12134 (N_12134,N_10894,N_10979);
nand U12135 (N_12135,N_11048,N_10949);
xor U12136 (N_12136,N_10922,N_11140);
nor U12137 (N_12137,N_10383,N_10441);
and U12138 (N_12138,N_10157,N_10829);
and U12139 (N_12139,N_10967,N_10809);
and U12140 (N_12140,N_11188,N_10570);
or U12141 (N_12141,N_11083,N_10744);
or U12142 (N_12142,N_10573,N_10098);
or U12143 (N_12143,N_10332,N_11225);
nor U12144 (N_12144,N_10067,N_10422);
or U12145 (N_12145,N_10712,N_10382);
xnor U12146 (N_12146,N_10087,N_10798);
nor U12147 (N_12147,N_10221,N_10119);
or U12148 (N_12148,N_10140,N_10475);
nor U12149 (N_12149,N_10648,N_10589);
or U12150 (N_12150,N_10171,N_10910);
nor U12151 (N_12151,N_10080,N_10018);
nor U12152 (N_12152,N_10521,N_10316);
and U12153 (N_12153,N_10234,N_10649);
nor U12154 (N_12154,N_10513,N_10429);
and U12155 (N_12155,N_10575,N_10058);
xor U12156 (N_12156,N_10689,N_10705);
nand U12157 (N_12157,N_10770,N_10541);
nor U12158 (N_12158,N_11216,N_10913);
nor U12159 (N_12159,N_10676,N_10323);
and U12160 (N_12160,N_11121,N_10192);
and U12161 (N_12161,N_10535,N_10422);
nand U12162 (N_12162,N_10471,N_10006);
nor U12163 (N_12163,N_11045,N_10325);
nand U12164 (N_12164,N_10881,N_10183);
nor U12165 (N_12165,N_10946,N_10801);
or U12166 (N_12166,N_11155,N_10874);
xor U12167 (N_12167,N_10171,N_10690);
or U12168 (N_12168,N_10397,N_10590);
nor U12169 (N_12169,N_10955,N_10487);
xor U12170 (N_12170,N_10974,N_10735);
nand U12171 (N_12171,N_10105,N_10936);
xor U12172 (N_12172,N_11216,N_10829);
xnor U12173 (N_12173,N_10700,N_10332);
nand U12174 (N_12174,N_10555,N_10093);
nor U12175 (N_12175,N_11057,N_10231);
and U12176 (N_12176,N_10862,N_10157);
nor U12177 (N_12177,N_10727,N_10776);
nand U12178 (N_12178,N_11210,N_10964);
nor U12179 (N_12179,N_10996,N_11120);
nand U12180 (N_12180,N_11035,N_10696);
xnor U12181 (N_12181,N_11008,N_10659);
nor U12182 (N_12182,N_10134,N_10296);
nor U12183 (N_12183,N_10425,N_10521);
and U12184 (N_12184,N_10898,N_10551);
or U12185 (N_12185,N_11096,N_10724);
or U12186 (N_12186,N_10808,N_10908);
and U12187 (N_12187,N_10129,N_10737);
nand U12188 (N_12188,N_10873,N_10563);
or U12189 (N_12189,N_10150,N_10298);
or U12190 (N_12190,N_10450,N_10278);
nand U12191 (N_12191,N_10862,N_10119);
and U12192 (N_12192,N_10361,N_11111);
xor U12193 (N_12193,N_10472,N_10723);
or U12194 (N_12194,N_10620,N_10898);
or U12195 (N_12195,N_10322,N_10572);
nand U12196 (N_12196,N_10531,N_11035);
nor U12197 (N_12197,N_10611,N_11038);
nor U12198 (N_12198,N_10538,N_11060);
nor U12199 (N_12199,N_11058,N_10476);
and U12200 (N_12200,N_10621,N_10492);
and U12201 (N_12201,N_10939,N_10639);
xor U12202 (N_12202,N_10481,N_10037);
xor U12203 (N_12203,N_10148,N_11040);
nor U12204 (N_12204,N_10353,N_10453);
or U12205 (N_12205,N_11155,N_11054);
nor U12206 (N_12206,N_11033,N_10818);
or U12207 (N_12207,N_11196,N_11044);
nand U12208 (N_12208,N_10588,N_10456);
xor U12209 (N_12209,N_10037,N_10812);
or U12210 (N_12210,N_10489,N_10254);
or U12211 (N_12211,N_10384,N_10532);
xnor U12212 (N_12212,N_10624,N_10047);
or U12213 (N_12213,N_10683,N_10877);
or U12214 (N_12214,N_10458,N_11238);
nand U12215 (N_12215,N_10387,N_10389);
nand U12216 (N_12216,N_10420,N_10408);
and U12217 (N_12217,N_10243,N_10339);
or U12218 (N_12218,N_10859,N_10010);
nand U12219 (N_12219,N_10720,N_10922);
and U12220 (N_12220,N_11244,N_10633);
nand U12221 (N_12221,N_10266,N_10512);
nand U12222 (N_12222,N_10604,N_10915);
or U12223 (N_12223,N_10571,N_10765);
or U12224 (N_12224,N_11174,N_10173);
or U12225 (N_12225,N_10611,N_11131);
nor U12226 (N_12226,N_10125,N_10597);
or U12227 (N_12227,N_10962,N_11056);
or U12228 (N_12228,N_10205,N_11102);
xnor U12229 (N_12229,N_11234,N_10726);
or U12230 (N_12230,N_10459,N_10570);
and U12231 (N_12231,N_10431,N_10556);
nor U12232 (N_12232,N_10965,N_11142);
xnor U12233 (N_12233,N_10255,N_10501);
nand U12234 (N_12234,N_10941,N_11174);
and U12235 (N_12235,N_10028,N_10823);
nor U12236 (N_12236,N_11022,N_10239);
nor U12237 (N_12237,N_10955,N_10028);
xor U12238 (N_12238,N_10347,N_10368);
nor U12239 (N_12239,N_10502,N_10853);
and U12240 (N_12240,N_10874,N_10037);
nand U12241 (N_12241,N_11183,N_10700);
xor U12242 (N_12242,N_10785,N_10320);
and U12243 (N_12243,N_11219,N_10964);
xor U12244 (N_12244,N_10159,N_11195);
or U12245 (N_12245,N_10595,N_10721);
nor U12246 (N_12246,N_11159,N_11204);
or U12247 (N_12247,N_10040,N_10697);
and U12248 (N_12248,N_10463,N_10884);
and U12249 (N_12249,N_10665,N_10361);
and U12250 (N_12250,N_10481,N_10876);
xnor U12251 (N_12251,N_10461,N_11081);
nand U12252 (N_12252,N_10953,N_11195);
xor U12253 (N_12253,N_10243,N_10716);
nor U12254 (N_12254,N_10387,N_10278);
or U12255 (N_12255,N_10622,N_11023);
and U12256 (N_12256,N_10960,N_10948);
nand U12257 (N_12257,N_10464,N_10776);
and U12258 (N_12258,N_10999,N_10367);
xnor U12259 (N_12259,N_10330,N_10077);
nand U12260 (N_12260,N_11103,N_11122);
xnor U12261 (N_12261,N_10767,N_11216);
or U12262 (N_12262,N_10160,N_10877);
xor U12263 (N_12263,N_10982,N_11079);
and U12264 (N_12264,N_10026,N_10444);
nand U12265 (N_12265,N_11214,N_10130);
or U12266 (N_12266,N_11188,N_10744);
or U12267 (N_12267,N_10265,N_11143);
and U12268 (N_12268,N_10918,N_11160);
xnor U12269 (N_12269,N_10140,N_10980);
xor U12270 (N_12270,N_10378,N_10691);
and U12271 (N_12271,N_10247,N_10579);
and U12272 (N_12272,N_11235,N_10472);
nor U12273 (N_12273,N_10586,N_10172);
xor U12274 (N_12274,N_10841,N_10477);
nand U12275 (N_12275,N_10714,N_11078);
or U12276 (N_12276,N_10580,N_10843);
nand U12277 (N_12277,N_10143,N_10302);
xnor U12278 (N_12278,N_10562,N_11121);
nor U12279 (N_12279,N_10533,N_10144);
or U12280 (N_12280,N_11214,N_10303);
and U12281 (N_12281,N_10053,N_10462);
and U12282 (N_12282,N_10774,N_10367);
nand U12283 (N_12283,N_10814,N_10650);
or U12284 (N_12284,N_10452,N_10516);
or U12285 (N_12285,N_10417,N_10080);
nor U12286 (N_12286,N_11184,N_10306);
nor U12287 (N_12287,N_10805,N_10100);
nor U12288 (N_12288,N_10361,N_10909);
or U12289 (N_12289,N_11101,N_10362);
or U12290 (N_12290,N_10841,N_10656);
nand U12291 (N_12291,N_10641,N_10177);
nor U12292 (N_12292,N_10466,N_10940);
nand U12293 (N_12293,N_10847,N_11055);
nand U12294 (N_12294,N_10538,N_10085);
and U12295 (N_12295,N_10741,N_10001);
and U12296 (N_12296,N_10119,N_10559);
nor U12297 (N_12297,N_11146,N_10972);
and U12298 (N_12298,N_10177,N_10376);
or U12299 (N_12299,N_10599,N_10320);
or U12300 (N_12300,N_10587,N_10773);
nor U12301 (N_12301,N_10854,N_10034);
or U12302 (N_12302,N_10246,N_10382);
xnor U12303 (N_12303,N_11159,N_10473);
and U12304 (N_12304,N_11077,N_10719);
nor U12305 (N_12305,N_11063,N_10938);
and U12306 (N_12306,N_11090,N_10161);
and U12307 (N_12307,N_10749,N_10333);
and U12308 (N_12308,N_11201,N_11139);
xnor U12309 (N_12309,N_10081,N_10640);
xnor U12310 (N_12310,N_10646,N_10996);
or U12311 (N_12311,N_10389,N_10760);
and U12312 (N_12312,N_10662,N_10405);
xnor U12313 (N_12313,N_11056,N_10223);
and U12314 (N_12314,N_10074,N_10320);
xnor U12315 (N_12315,N_10808,N_10775);
and U12316 (N_12316,N_11150,N_10530);
and U12317 (N_12317,N_10953,N_10476);
or U12318 (N_12318,N_10726,N_10675);
xor U12319 (N_12319,N_10175,N_10232);
and U12320 (N_12320,N_10858,N_10428);
and U12321 (N_12321,N_10803,N_11095);
or U12322 (N_12322,N_10538,N_10612);
and U12323 (N_12323,N_10152,N_10224);
or U12324 (N_12324,N_10890,N_10489);
xor U12325 (N_12325,N_10530,N_10325);
or U12326 (N_12326,N_10513,N_11003);
nand U12327 (N_12327,N_10607,N_11125);
nand U12328 (N_12328,N_10833,N_11163);
or U12329 (N_12329,N_10544,N_10083);
and U12330 (N_12330,N_10276,N_10528);
xor U12331 (N_12331,N_11125,N_11089);
and U12332 (N_12332,N_10537,N_10409);
xnor U12333 (N_12333,N_10619,N_10510);
nand U12334 (N_12334,N_10535,N_10384);
nor U12335 (N_12335,N_10913,N_10064);
nor U12336 (N_12336,N_10955,N_10749);
or U12337 (N_12337,N_11048,N_10628);
or U12338 (N_12338,N_11037,N_11038);
nor U12339 (N_12339,N_10112,N_10777);
or U12340 (N_12340,N_10481,N_10711);
or U12341 (N_12341,N_10505,N_10465);
nand U12342 (N_12342,N_10101,N_10278);
nor U12343 (N_12343,N_11034,N_10296);
and U12344 (N_12344,N_10556,N_10941);
or U12345 (N_12345,N_10607,N_10432);
nor U12346 (N_12346,N_10265,N_10888);
or U12347 (N_12347,N_11081,N_10569);
nor U12348 (N_12348,N_10686,N_10012);
nand U12349 (N_12349,N_11034,N_10199);
or U12350 (N_12350,N_10981,N_10014);
and U12351 (N_12351,N_10958,N_11064);
and U12352 (N_12352,N_10762,N_10365);
and U12353 (N_12353,N_10372,N_10685);
nand U12354 (N_12354,N_11181,N_10365);
nor U12355 (N_12355,N_10460,N_10988);
nor U12356 (N_12356,N_10870,N_10900);
and U12357 (N_12357,N_11065,N_10043);
and U12358 (N_12358,N_10795,N_10452);
xnor U12359 (N_12359,N_10226,N_10715);
xnor U12360 (N_12360,N_10173,N_10602);
nor U12361 (N_12361,N_11236,N_10521);
or U12362 (N_12362,N_11053,N_11049);
and U12363 (N_12363,N_10401,N_11231);
xor U12364 (N_12364,N_10589,N_11232);
xor U12365 (N_12365,N_10754,N_10587);
nor U12366 (N_12366,N_11096,N_10779);
xor U12367 (N_12367,N_10333,N_10150);
nand U12368 (N_12368,N_10546,N_10922);
nor U12369 (N_12369,N_10934,N_11107);
nor U12370 (N_12370,N_11156,N_10707);
xor U12371 (N_12371,N_11113,N_11014);
and U12372 (N_12372,N_10463,N_11136);
nand U12373 (N_12373,N_10558,N_10562);
or U12374 (N_12374,N_10615,N_10915);
xor U12375 (N_12375,N_10870,N_10455);
nand U12376 (N_12376,N_10714,N_10109);
or U12377 (N_12377,N_10469,N_10045);
or U12378 (N_12378,N_11095,N_10808);
xnor U12379 (N_12379,N_10022,N_10902);
and U12380 (N_12380,N_10510,N_10018);
xor U12381 (N_12381,N_10666,N_10055);
nand U12382 (N_12382,N_10570,N_10527);
nor U12383 (N_12383,N_10639,N_10987);
xnor U12384 (N_12384,N_10628,N_10231);
xnor U12385 (N_12385,N_10284,N_10967);
nand U12386 (N_12386,N_10606,N_10948);
xor U12387 (N_12387,N_11197,N_10328);
or U12388 (N_12388,N_10027,N_10413);
nor U12389 (N_12389,N_10110,N_10654);
xor U12390 (N_12390,N_10720,N_10049);
xor U12391 (N_12391,N_10467,N_10080);
and U12392 (N_12392,N_10480,N_10385);
and U12393 (N_12393,N_10124,N_10597);
or U12394 (N_12394,N_11225,N_11158);
and U12395 (N_12395,N_10085,N_10444);
or U12396 (N_12396,N_10998,N_11172);
nand U12397 (N_12397,N_10413,N_11240);
nand U12398 (N_12398,N_10382,N_10188);
nor U12399 (N_12399,N_10144,N_10493);
and U12400 (N_12400,N_11104,N_11024);
xor U12401 (N_12401,N_11080,N_10623);
nand U12402 (N_12402,N_10696,N_10822);
nor U12403 (N_12403,N_11067,N_11209);
nand U12404 (N_12404,N_10014,N_10452);
xor U12405 (N_12405,N_10152,N_11133);
or U12406 (N_12406,N_10229,N_10284);
or U12407 (N_12407,N_10573,N_10563);
nand U12408 (N_12408,N_10050,N_11110);
nand U12409 (N_12409,N_11180,N_11118);
and U12410 (N_12410,N_10099,N_10636);
nand U12411 (N_12411,N_10272,N_10607);
or U12412 (N_12412,N_10542,N_10663);
nand U12413 (N_12413,N_10840,N_10337);
xor U12414 (N_12414,N_10004,N_11149);
nand U12415 (N_12415,N_10316,N_10000);
nand U12416 (N_12416,N_10335,N_10630);
nor U12417 (N_12417,N_10783,N_10090);
nand U12418 (N_12418,N_10415,N_11035);
nor U12419 (N_12419,N_10986,N_10056);
and U12420 (N_12420,N_11084,N_10992);
or U12421 (N_12421,N_10069,N_10621);
or U12422 (N_12422,N_10287,N_10425);
nor U12423 (N_12423,N_10281,N_10456);
nor U12424 (N_12424,N_10184,N_10768);
or U12425 (N_12425,N_10516,N_10914);
and U12426 (N_12426,N_10765,N_10150);
xor U12427 (N_12427,N_10209,N_10345);
and U12428 (N_12428,N_10888,N_10299);
nor U12429 (N_12429,N_10678,N_10238);
or U12430 (N_12430,N_10747,N_10670);
or U12431 (N_12431,N_10822,N_10845);
xnor U12432 (N_12432,N_10064,N_10161);
nor U12433 (N_12433,N_10190,N_10191);
and U12434 (N_12434,N_10449,N_10599);
or U12435 (N_12435,N_10566,N_10722);
or U12436 (N_12436,N_10185,N_10049);
nand U12437 (N_12437,N_10878,N_10933);
nor U12438 (N_12438,N_10849,N_10138);
or U12439 (N_12439,N_10031,N_10835);
nand U12440 (N_12440,N_10901,N_10360);
and U12441 (N_12441,N_10305,N_10111);
or U12442 (N_12442,N_10330,N_10011);
xnor U12443 (N_12443,N_11102,N_10544);
nand U12444 (N_12444,N_10705,N_10803);
and U12445 (N_12445,N_11143,N_10203);
nand U12446 (N_12446,N_11237,N_10113);
and U12447 (N_12447,N_10050,N_10001);
and U12448 (N_12448,N_10590,N_10822);
or U12449 (N_12449,N_10389,N_10208);
or U12450 (N_12450,N_10071,N_10880);
nor U12451 (N_12451,N_11189,N_10171);
nand U12452 (N_12452,N_11204,N_10613);
or U12453 (N_12453,N_10850,N_10635);
nand U12454 (N_12454,N_10763,N_11016);
nand U12455 (N_12455,N_10999,N_10385);
nor U12456 (N_12456,N_10905,N_10233);
and U12457 (N_12457,N_10785,N_10837);
or U12458 (N_12458,N_10666,N_10129);
nand U12459 (N_12459,N_10781,N_10377);
nor U12460 (N_12460,N_10328,N_11192);
xor U12461 (N_12461,N_10875,N_10581);
or U12462 (N_12462,N_10662,N_11147);
or U12463 (N_12463,N_10620,N_10319);
nand U12464 (N_12464,N_10868,N_10594);
xnor U12465 (N_12465,N_10993,N_10043);
nand U12466 (N_12466,N_11056,N_10980);
nand U12467 (N_12467,N_11102,N_10464);
or U12468 (N_12468,N_10883,N_10540);
xnor U12469 (N_12469,N_11206,N_11190);
or U12470 (N_12470,N_10266,N_11108);
nor U12471 (N_12471,N_10539,N_11165);
or U12472 (N_12472,N_10399,N_10159);
nor U12473 (N_12473,N_10159,N_11153);
or U12474 (N_12474,N_11202,N_10420);
or U12475 (N_12475,N_10997,N_11012);
and U12476 (N_12476,N_10737,N_10422);
nor U12477 (N_12477,N_10048,N_10203);
or U12478 (N_12478,N_10359,N_10993);
nand U12479 (N_12479,N_10741,N_10776);
nand U12480 (N_12480,N_10606,N_10463);
or U12481 (N_12481,N_10192,N_10795);
nand U12482 (N_12482,N_11180,N_10956);
nor U12483 (N_12483,N_10215,N_10716);
and U12484 (N_12484,N_10270,N_11242);
and U12485 (N_12485,N_10586,N_10821);
xor U12486 (N_12486,N_10961,N_10651);
nor U12487 (N_12487,N_10380,N_10160);
nand U12488 (N_12488,N_10041,N_10653);
or U12489 (N_12489,N_10790,N_11114);
xnor U12490 (N_12490,N_11197,N_10883);
xnor U12491 (N_12491,N_10629,N_10276);
and U12492 (N_12492,N_10269,N_11180);
nor U12493 (N_12493,N_11239,N_10011);
nand U12494 (N_12494,N_10508,N_10914);
or U12495 (N_12495,N_10782,N_10694);
or U12496 (N_12496,N_10345,N_10103);
nor U12497 (N_12497,N_11147,N_10933);
or U12498 (N_12498,N_10128,N_10163);
nor U12499 (N_12499,N_10789,N_10951);
nand U12500 (N_12500,N_12496,N_11689);
nor U12501 (N_12501,N_12064,N_12292);
nor U12502 (N_12502,N_12422,N_11871);
or U12503 (N_12503,N_12188,N_12439);
or U12504 (N_12504,N_12408,N_12048);
and U12505 (N_12505,N_11629,N_12053);
or U12506 (N_12506,N_11777,N_12202);
nor U12507 (N_12507,N_11553,N_11607);
xor U12508 (N_12508,N_11672,N_12010);
or U12509 (N_12509,N_11875,N_12432);
or U12510 (N_12510,N_11536,N_11865);
nor U12511 (N_12511,N_12070,N_11785);
or U12512 (N_12512,N_11469,N_11726);
or U12513 (N_12513,N_11575,N_12199);
and U12514 (N_12514,N_12276,N_12478);
or U12515 (N_12515,N_11491,N_12335);
nand U12516 (N_12516,N_12300,N_12039);
nand U12517 (N_12517,N_11953,N_11964);
nand U12518 (N_12518,N_11855,N_11988);
xor U12519 (N_12519,N_12215,N_12475);
nand U12520 (N_12520,N_12066,N_11428);
or U12521 (N_12521,N_12111,N_12195);
and U12522 (N_12522,N_12116,N_12433);
nand U12523 (N_12523,N_11878,N_11899);
or U12524 (N_12524,N_12406,N_12026);
nor U12525 (N_12525,N_11530,N_11654);
nor U12526 (N_12526,N_12012,N_11690);
or U12527 (N_12527,N_11405,N_12434);
nor U12528 (N_12528,N_11615,N_12370);
xnor U12529 (N_12529,N_11567,N_11359);
nor U12530 (N_12530,N_12394,N_12045);
xor U12531 (N_12531,N_11418,N_12431);
or U12532 (N_12532,N_11922,N_11681);
or U12533 (N_12533,N_12391,N_11515);
and U12534 (N_12534,N_12031,N_12062);
xnor U12535 (N_12535,N_11926,N_11912);
xnor U12536 (N_12536,N_12281,N_12378);
nand U12537 (N_12537,N_11872,N_11368);
nand U12538 (N_12538,N_12258,N_11741);
nor U12539 (N_12539,N_11829,N_11714);
nand U12540 (N_12540,N_12207,N_11773);
xor U12541 (N_12541,N_12119,N_12118);
xor U12542 (N_12542,N_11464,N_11774);
or U12543 (N_12543,N_12458,N_11967);
nand U12544 (N_12544,N_12454,N_11683);
nand U12545 (N_12545,N_12229,N_11622);
nand U12546 (N_12546,N_11397,N_12241);
or U12547 (N_12547,N_11549,N_11998);
nor U12548 (N_12548,N_12392,N_11627);
or U12549 (N_12549,N_11770,N_12283);
nor U12550 (N_12550,N_12459,N_12102);
and U12551 (N_12551,N_11273,N_11430);
nand U12552 (N_12552,N_12327,N_12137);
or U12553 (N_12553,N_11942,N_11422);
nor U12554 (N_12554,N_11753,N_11966);
or U12555 (N_12555,N_11749,N_11617);
or U12556 (N_12556,N_12447,N_12257);
nand U12557 (N_12557,N_12307,N_11279);
xor U12558 (N_12558,N_11700,N_12234);
xor U12559 (N_12559,N_11995,N_11792);
or U12560 (N_12560,N_12375,N_12329);
nand U12561 (N_12561,N_11825,N_11885);
and U12562 (N_12562,N_11501,N_12443);
and U12563 (N_12563,N_12106,N_12467);
xnor U12564 (N_12564,N_11302,N_11786);
nand U12565 (N_12565,N_12468,N_11606);
or U12566 (N_12566,N_11573,N_11623);
nand U12567 (N_12567,N_12349,N_12009);
nand U12568 (N_12568,N_11703,N_11844);
nand U12569 (N_12569,N_11594,N_11579);
nand U12570 (N_12570,N_12011,N_11781);
xnor U12571 (N_12571,N_12237,N_11776);
and U12572 (N_12572,N_12168,N_12180);
xnor U12573 (N_12573,N_12423,N_11642);
and U12574 (N_12574,N_11746,N_11718);
and U12575 (N_12575,N_11492,N_12022);
or U12576 (N_12576,N_11584,N_11434);
or U12577 (N_12577,N_11616,N_11559);
nand U12578 (N_12578,N_12186,N_11643);
nand U12579 (N_12579,N_11637,N_11443);
xor U12580 (N_12580,N_11975,N_11858);
nand U12581 (N_12581,N_11495,N_12206);
or U12582 (N_12582,N_11480,N_12428);
xnor U12583 (N_12583,N_11512,N_11389);
xor U12584 (N_12584,N_12196,N_12448);
nand U12585 (N_12585,N_11602,N_12044);
nand U12586 (N_12586,N_12270,N_11934);
or U12587 (N_12587,N_11997,N_11488);
xor U12588 (N_12588,N_12152,N_11601);
nand U12589 (N_12589,N_12249,N_12465);
and U12590 (N_12590,N_12181,N_11710);
or U12591 (N_12591,N_12008,N_12182);
nor U12592 (N_12592,N_11653,N_11386);
nand U12593 (N_12593,N_11465,N_12101);
xor U12594 (N_12594,N_11380,N_11752);
and U12595 (N_12595,N_11661,N_11704);
nor U12596 (N_12596,N_12125,N_11338);
xor U12597 (N_12597,N_11887,N_12295);
xnor U12598 (N_12598,N_11842,N_12001);
and U12599 (N_12599,N_11324,N_11687);
nand U12600 (N_12600,N_11748,N_11897);
or U12601 (N_12601,N_11592,N_11668);
nor U12602 (N_12602,N_11295,N_11659);
nor U12603 (N_12603,N_11271,N_11709);
nand U12604 (N_12604,N_11522,N_11437);
nor U12605 (N_12605,N_12185,N_12219);
nand U12606 (N_12606,N_12273,N_11727);
xor U12607 (N_12607,N_12282,N_12301);
nor U12608 (N_12608,N_11647,N_12387);
and U12609 (N_12609,N_11630,N_11846);
or U12610 (N_12610,N_11587,N_11980);
xnor U12611 (N_12611,N_11640,N_12252);
or U12612 (N_12612,N_11340,N_12204);
xnor U12613 (N_12613,N_11821,N_12201);
nor U12614 (N_12614,N_11904,N_11564);
or U12615 (N_12615,N_12140,N_11632);
nand U12616 (N_12616,N_12145,N_12463);
or U12617 (N_12617,N_11981,N_12487);
and U12618 (N_12618,N_11698,N_12404);
and U12619 (N_12619,N_11414,N_11784);
nor U12620 (N_12620,N_11985,N_12455);
xnor U12621 (N_12621,N_11276,N_12484);
and U12622 (N_12622,N_11365,N_11736);
or U12623 (N_12623,N_11543,N_12225);
xor U12624 (N_12624,N_11528,N_11369);
and U12625 (N_12625,N_11288,N_12124);
xor U12626 (N_12626,N_11470,N_11444);
xnor U12627 (N_12627,N_11673,N_11944);
xnor U12628 (N_12628,N_12228,N_11987);
and U12629 (N_12629,N_12223,N_11508);
or U12630 (N_12630,N_12357,N_11693);
xor U12631 (N_12631,N_11487,N_11525);
nand U12632 (N_12632,N_11345,N_11660);
or U12633 (N_12633,N_12081,N_12187);
xnor U12634 (N_12634,N_12025,N_11253);
xnor U12635 (N_12635,N_11984,N_11486);
nand U12636 (N_12636,N_11963,N_11524);
or U12637 (N_12637,N_12379,N_11992);
or U12638 (N_12638,N_11520,N_12351);
nor U12639 (N_12639,N_12035,N_11309);
nand U12640 (N_12640,N_11863,N_11809);
xor U12641 (N_12641,N_11577,N_11699);
nand U12642 (N_12642,N_11945,N_12261);
nor U12643 (N_12643,N_12013,N_12397);
and U12644 (N_12644,N_11826,N_12172);
or U12645 (N_12645,N_12189,N_11558);
or U12646 (N_12646,N_11381,N_12007);
nor U12647 (N_12647,N_11481,N_11823);
nand U12648 (N_12648,N_11466,N_11645);
nor U12649 (N_12649,N_11828,N_12127);
or U12650 (N_12650,N_11278,N_12359);
nand U12651 (N_12651,N_12193,N_11494);
nand U12652 (N_12652,N_12103,N_12176);
or U12653 (N_12653,N_12197,N_11835);
nand U12654 (N_12654,N_11320,N_12299);
nor U12655 (N_12655,N_12385,N_12499);
nor U12656 (N_12656,N_11420,N_11250);
and U12657 (N_12657,N_11316,N_11820);
and U12658 (N_12658,N_11895,N_11256);
or U12659 (N_12659,N_11837,N_11462);
nand U12660 (N_12660,N_12060,N_11356);
nand U12661 (N_12661,N_11590,N_12346);
and U12662 (N_12662,N_11747,N_11541);
or U12663 (N_12663,N_11586,N_12494);
xnor U12664 (N_12664,N_11918,N_12020);
nand U12665 (N_12665,N_11384,N_12369);
and U12666 (N_12666,N_12112,N_12485);
and U12667 (N_12667,N_12438,N_12266);
xnor U12668 (N_12668,N_11688,N_11952);
or U12669 (N_12669,N_11301,N_12398);
xor U12670 (N_12670,N_11857,N_12479);
nor U12671 (N_12671,N_11652,N_11403);
nor U12672 (N_12672,N_11388,N_12452);
or U12673 (N_12673,N_12161,N_11983);
xor U12674 (N_12674,N_11676,N_11290);
nor U12675 (N_12675,N_12141,N_12098);
or U12676 (N_12676,N_11377,N_12184);
and U12677 (N_12677,N_11373,N_11789);
nand U12678 (N_12678,N_11949,N_11956);
nand U12679 (N_12679,N_12361,N_12272);
and U12680 (N_12680,N_11516,N_11691);
and U12681 (N_12681,N_11419,N_11999);
xnor U12682 (N_12682,N_12497,N_11513);
or U12683 (N_12683,N_11533,N_11880);
xor U12684 (N_12684,N_11805,N_12040);
nand U12685 (N_12685,N_12156,N_11730);
or U12686 (N_12686,N_11901,N_12381);
and U12687 (N_12687,N_11599,N_11424);
nand U12688 (N_12688,N_11941,N_11286);
nor U12689 (N_12689,N_11604,N_11498);
nand U12690 (N_12690,N_11864,N_12440);
or U12691 (N_12691,N_11796,N_11542);
and U12692 (N_12692,N_11772,N_12003);
nand U12693 (N_12693,N_11296,N_11252);
xor U12694 (N_12694,N_12298,N_11951);
xor U12695 (N_12695,N_12100,N_11426);
and U12696 (N_12696,N_11475,N_11649);
or U12697 (N_12697,N_11595,N_11923);
and U12698 (N_12698,N_11908,N_12049);
or U12699 (N_12699,N_12306,N_11634);
and U12700 (N_12700,N_12260,N_11408);
and U12701 (N_12701,N_12233,N_11518);
nand U12702 (N_12702,N_12399,N_11308);
and U12703 (N_12703,N_12280,N_12303);
xnor U12704 (N_12704,N_11264,N_11717);
and U12705 (N_12705,N_12166,N_11790);
xor U12706 (N_12706,N_11743,N_11813);
xnor U12707 (N_12707,N_12079,N_11605);
nor U12708 (N_12708,N_11490,N_12173);
nor U12709 (N_12709,N_11755,N_11358);
and U12710 (N_12710,N_12004,N_11439);
xnor U12711 (N_12711,N_12212,N_12412);
xnor U12712 (N_12712,N_11385,N_11531);
xor U12713 (N_12713,N_11836,N_11500);
xor U12714 (N_12714,N_11280,N_12211);
and U12715 (N_12715,N_11331,N_12149);
or U12716 (N_12716,N_12200,N_11474);
or U12717 (N_12717,N_11968,N_11955);
nor U12718 (N_12718,N_11609,N_11803);
or U12719 (N_12719,N_11272,N_11351);
nand U12720 (N_12720,N_11565,N_11502);
and U12721 (N_12721,N_12371,N_11884);
or U12722 (N_12722,N_11757,N_12435);
nand U12723 (N_12723,N_11775,N_12084);
nand U12724 (N_12724,N_12123,N_11969);
nor U12725 (N_12725,N_12076,N_12492);
xnor U12726 (N_12726,N_12236,N_12338);
nor U12727 (N_12727,N_11454,N_12164);
and U12728 (N_12728,N_11666,N_12221);
nand U12729 (N_12729,N_11493,N_12238);
nor U12730 (N_12730,N_11390,N_12174);
nor U12731 (N_12731,N_12402,N_11732);
xor U12732 (N_12732,N_12462,N_11504);
or U12733 (N_12733,N_11337,N_11357);
or U12734 (N_12734,N_11436,N_11399);
and U12735 (N_12735,N_11832,N_11333);
and U12736 (N_12736,N_11519,N_12109);
xnor U12737 (N_12737,N_11978,N_11299);
nor U12738 (N_12738,N_11603,N_12409);
nand U12739 (N_12739,N_12445,N_12038);
nor U12740 (N_12740,N_11762,N_11862);
xor U12741 (N_12741,N_12469,N_12115);
and U12742 (N_12742,N_11557,N_11274);
and U12743 (N_12743,N_11538,N_11819);
and U12744 (N_12744,N_12471,N_12477);
or U12745 (N_12745,N_12348,N_12362);
nand U12746 (N_12746,N_11550,N_11737);
or U12747 (N_12747,N_12466,N_12470);
or U12748 (N_12748,N_12473,N_11562);
or U12749 (N_12749,N_11947,N_12364);
nand U12750 (N_12750,N_11348,N_11719);
nand U12751 (N_12751,N_11641,N_11868);
and U12752 (N_12752,N_12029,N_11334);
xor U12753 (N_12753,N_11341,N_11795);
xnor U12754 (N_12754,N_11970,N_11860);
and U12755 (N_12755,N_11371,N_11639);
and U12756 (N_12756,N_11489,N_11793);
nand U12757 (N_12757,N_12293,N_12092);
and U12758 (N_12758,N_11914,N_12099);
or U12759 (N_12759,N_11900,N_11453);
or U12760 (N_12760,N_11758,N_11903);
nor U12761 (N_12761,N_12311,N_11319);
nand U12762 (N_12762,N_11910,N_11539);
nor U12763 (N_12763,N_11263,N_11415);
xnor U12764 (N_12764,N_11665,N_11410);
nand U12765 (N_12765,N_11429,N_11658);
nand U12766 (N_12766,N_11935,N_12113);
xor U12767 (N_12767,N_11958,N_12322);
xnor U12768 (N_12768,N_12318,N_11725);
or U12769 (N_12769,N_12136,N_12388);
nand U12770 (N_12770,N_11906,N_11636);
or U12771 (N_12771,N_11435,N_11313);
nor U12772 (N_12772,N_11650,N_12155);
and U12773 (N_12773,N_11877,N_12489);
nor U12774 (N_12774,N_11363,N_11677);
nor U12775 (N_12775,N_12222,N_11794);
and U12776 (N_12776,N_11382,N_12146);
nand U12777 (N_12777,N_11684,N_12372);
or U12778 (N_12778,N_11750,N_12262);
nor U12779 (N_12779,N_12414,N_11303);
nor U12780 (N_12780,N_12177,N_12345);
nand U12781 (N_12781,N_11318,N_12368);
and U12782 (N_12782,N_12151,N_12305);
nand U12783 (N_12783,N_12417,N_11411);
or U12784 (N_12784,N_12218,N_11893);
or U12785 (N_12785,N_11920,N_12358);
and U12786 (N_12786,N_11670,N_12246);
nand U12787 (N_12787,N_12091,N_12042);
nand U12788 (N_12788,N_12481,N_12396);
nor U12789 (N_12789,N_11268,N_11433);
nand U12790 (N_12790,N_11578,N_11413);
nand U12791 (N_12791,N_11610,N_11378);
or U12792 (N_12792,N_11300,N_12165);
nand U12793 (N_12793,N_11305,N_12050);
or U12794 (N_12794,N_11529,N_11555);
nand U12795 (N_12795,N_11458,N_11767);
or U12796 (N_12796,N_12328,N_11343);
or U12797 (N_12797,N_11812,N_12179);
xnor U12798 (N_12798,N_11284,N_12107);
or U12799 (N_12799,N_12014,N_11817);
or U12800 (N_12800,N_12024,N_11355);
xor U12801 (N_12801,N_11898,N_11255);
and U12802 (N_12802,N_11838,N_11731);
nor U12803 (N_12803,N_12134,N_12167);
nand U12804 (N_12804,N_11655,N_11421);
nor U12805 (N_12805,N_12005,N_11635);
nor U12806 (N_12806,N_11756,N_11662);
nor U12807 (N_12807,N_11383,N_11619);
and U12808 (N_12808,N_11497,N_11322);
nor U12809 (N_12809,N_11976,N_11948);
xor U12810 (N_12810,N_12019,N_12190);
xor U12811 (N_12811,N_11568,N_12426);
or U12812 (N_12812,N_11409,N_11327);
xor U12813 (N_12813,N_11694,N_12080);
and U12814 (N_12814,N_11585,N_11769);
and U12815 (N_12815,N_11526,N_11505);
nor U12816 (N_12816,N_12336,N_12243);
nand U12817 (N_12817,N_12421,N_11972);
or U12818 (N_12818,N_12367,N_11251);
nor U12819 (N_12819,N_11275,N_12418);
nor U12820 (N_12820,N_11800,N_12491);
nor U12821 (N_12821,N_11993,N_12352);
nor U12822 (N_12822,N_11833,N_12095);
or U12823 (N_12823,N_11834,N_12425);
xor U12824 (N_12824,N_11818,N_11406);
nor U12825 (N_12825,N_12110,N_12446);
nand U12826 (N_12826,N_11851,N_12265);
nor U12827 (N_12827,N_12480,N_11569);
nor U12828 (N_12828,N_12169,N_11448);
xor U12829 (N_12829,N_11721,N_11315);
xnor U12830 (N_12830,N_12263,N_12380);
nand U12831 (N_12831,N_12383,N_11929);
and U12832 (N_12832,N_11994,N_11979);
nand U12833 (N_12833,N_12317,N_12316);
xor U12834 (N_12834,N_12490,N_12309);
and U12835 (N_12835,N_11452,N_12377);
xnor U12836 (N_12836,N_11277,N_11478);
or U12837 (N_12837,N_11574,N_11854);
xor U12838 (N_12838,N_11407,N_11745);
and U12839 (N_12839,N_11788,N_11467);
or U12840 (N_12840,N_11937,N_11631);
and U12841 (N_12841,N_12224,N_12302);
xnor U12842 (N_12842,N_11472,N_12374);
and U12843 (N_12843,N_12068,N_12386);
nand U12844 (N_12844,N_12245,N_11808);
and U12845 (N_12845,N_11423,N_11678);
nand U12846 (N_12846,N_11265,N_12122);
xor U12847 (N_12847,N_11674,N_12131);
xor U12848 (N_12848,N_11282,N_12356);
and U12849 (N_12849,N_11644,N_11664);
nand U12850 (N_12850,N_11722,N_12393);
xnor U12851 (N_12851,N_11551,N_11460);
nand U12852 (N_12852,N_11445,N_11896);
xor U12853 (N_12853,N_11950,N_12493);
or U12854 (N_12854,N_11881,N_11325);
xnor U12855 (N_12855,N_12271,N_12006);
nand U12856 (N_12856,N_11471,N_12442);
and U12857 (N_12857,N_11742,N_12077);
nor U12858 (N_12858,N_12023,N_12208);
nor U12859 (N_12859,N_11911,N_11889);
or U12860 (N_12860,N_12056,N_12373);
xnor U12861 (N_12861,N_12158,N_12139);
nand U12862 (N_12862,N_12148,N_12400);
nor U12863 (N_12863,N_11394,N_11392);
and U12864 (N_12864,N_11771,N_12153);
xnor U12865 (N_12865,N_11335,N_12451);
nor U12866 (N_12866,N_12170,N_12033);
xor U12867 (N_12867,N_12191,N_11600);
and U12868 (N_12868,N_11425,N_11523);
and U12869 (N_12869,N_12350,N_12287);
and U12870 (N_12870,N_11576,N_11807);
nand U12871 (N_12871,N_11989,N_12021);
nor U12872 (N_12872,N_12483,N_11907);
and U12873 (N_12873,N_11924,N_11571);
and U12874 (N_12874,N_11892,N_12097);
nor U12875 (N_12875,N_11375,N_11822);
xor U12876 (N_12876,N_11563,N_12032);
nand U12877 (N_12877,N_11883,N_12157);
and U12878 (N_12878,N_12002,N_11686);
nor U12879 (N_12879,N_11572,N_11810);
xnor U12880 (N_12880,N_12147,N_12120);
and U12881 (N_12881,N_12135,N_12331);
nor U12882 (N_12882,N_12363,N_11285);
and U12883 (N_12883,N_11283,N_11259);
xnor U12884 (N_12884,N_12420,N_11463);
or U12885 (N_12885,N_12213,N_11352);
xor U12886 (N_12886,N_11485,N_11957);
and U12887 (N_12887,N_11977,N_11442);
nor U12888 (N_12888,N_11905,N_12086);
nand U12889 (N_12889,N_12476,N_11974);
nand U12890 (N_12890,N_12144,N_11540);
nand U12891 (N_12891,N_11330,N_11449);
nor U12892 (N_12892,N_12132,N_12275);
and U12893 (N_12893,N_11715,N_11257);
or U12894 (N_12894,N_12194,N_12405);
xor U12895 (N_12895,N_12083,N_11927);
or U12896 (N_12896,N_11729,N_12126);
or U12897 (N_12897,N_11882,N_11593);
and U12898 (N_12898,N_11734,N_12339);
nand U12899 (N_12899,N_11759,N_12360);
nand U12900 (N_12900,N_12251,N_12067);
nor U12901 (N_12901,N_11740,N_11780);
nand U12902 (N_12902,N_11266,N_11427);
and U12903 (N_12903,N_12365,N_11298);
xor U12904 (N_12904,N_11991,N_11815);
or U12905 (N_12905,N_11801,N_12296);
or U12906 (N_12906,N_11560,N_12482);
xnor U12907 (N_12907,N_11936,N_12209);
xor U12908 (N_12908,N_12340,N_11724);
or U12909 (N_12909,N_11669,N_12074);
nor U12910 (N_12910,N_11479,N_11909);
nor U12911 (N_12911,N_11930,N_11638);
nor U12912 (N_12912,N_12376,N_12244);
or U12913 (N_12913,N_12078,N_12250);
or U12914 (N_12914,N_11633,N_11367);
xnor U12915 (N_12915,N_11798,N_12036);
and U12916 (N_12916,N_11986,N_11496);
and U12917 (N_12917,N_12216,N_11412);
and U12918 (N_12918,N_11451,N_12178);
nor U12919 (N_12919,N_11913,N_11393);
or U12920 (N_12920,N_11827,N_12324);
nor U12921 (N_12921,N_11326,N_11917);
or U12922 (N_12922,N_12389,N_12264);
nand U12923 (N_12923,N_11768,N_12429);
nor U12924 (N_12924,N_11267,N_12063);
nand U12925 (N_12925,N_11514,N_11570);
nor U12926 (N_12926,N_11431,N_12051);
or U12927 (N_12927,N_11919,N_11583);
or U12928 (N_12928,N_11712,N_12310);
nor U12929 (N_12929,N_12288,N_12474);
and U12930 (N_12930,N_11544,N_11806);
or U12931 (N_12931,N_11890,N_12284);
nor U12932 (N_12932,N_12332,N_11713);
nor U12933 (N_12933,N_11306,N_12093);
nor U12934 (N_12934,N_11360,N_12017);
xor U12935 (N_12935,N_12232,N_11545);
or U12936 (N_12936,N_11561,N_11840);
xnor U12937 (N_12937,N_11852,N_12312);
or U12938 (N_12938,N_12382,N_11395);
nand U12939 (N_12939,N_12415,N_12037);
or U12940 (N_12940,N_11962,N_11582);
nor U12941 (N_12941,N_12015,N_12088);
xor U12942 (N_12942,N_12105,N_11843);
and U12943 (N_12943,N_12150,N_11735);
xnor U12944 (N_12944,N_11446,N_12294);
xnor U12945 (N_12945,N_12138,N_12355);
xnor U12946 (N_12946,N_11738,N_12096);
or U12947 (N_12947,N_11656,N_12297);
xnor U12948 (N_12948,N_11613,N_11596);
xnor U12949 (N_12949,N_11350,N_11799);
or U12950 (N_12950,N_12085,N_11547);
nor U12951 (N_12951,N_11902,N_11961);
nand U12952 (N_12952,N_11971,N_11839);
nor U12953 (N_12953,N_11866,N_11733);
nand U12954 (N_12954,N_11310,N_11321);
xnor U12955 (N_12955,N_12046,N_11294);
and U12956 (N_12956,N_11754,N_12341);
xnor U12957 (N_12957,N_11402,N_11830);
nor U12958 (N_12958,N_11608,N_11261);
and U12959 (N_12959,N_12498,N_11626);
or U12960 (N_12960,N_12286,N_11816);
xnor U12961 (N_12961,N_11708,N_11482);
xnor U12962 (N_12962,N_11705,N_11939);
or U12963 (N_12963,N_11845,N_11891);
and U12964 (N_12964,N_12424,N_11778);
xnor U12965 (N_12965,N_12043,N_11332);
and U12966 (N_12966,N_11928,N_11940);
or U12967 (N_12967,N_12047,N_11802);
or U12968 (N_12968,N_11361,N_11447);
nand U12969 (N_12969,N_11459,N_12082);
nor U12970 (N_12970,N_11461,N_11695);
xnor U12971 (N_12971,N_11621,N_11269);
nand U12972 (N_12972,N_12220,N_11933);
nor U12973 (N_12973,N_11438,N_12242);
nand U12974 (N_12974,N_11618,N_12308);
and U12975 (N_12975,N_11648,N_12325);
and U12976 (N_12976,N_12071,N_11270);
nor U12977 (N_12977,N_11260,N_11346);
xor U12978 (N_12978,N_11293,N_11620);
nor U12979 (N_12979,N_11943,N_12163);
and U12980 (N_12980,N_11366,N_11954);
nand U12981 (N_12981,N_11362,N_12069);
and U12982 (N_12982,N_11783,N_11879);
or U12983 (N_12983,N_12256,N_11886);
and U12984 (N_12984,N_12291,N_12267);
or U12985 (N_12985,N_11938,N_12192);
and U12986 (N_12986,N_11646,N_11312);
nor U12987 (N_12987,N_11441,N_11292);
or U12988 (N_12988,N_11517,N_11317);
or U12989 (N_12989,N_12472,N_11307);
nor U12990 (N_12990,N_12027,N_12133);
xnor U12991 (N_12991,N_11849,N_11763);
and U12992 (N_12992,N_12090,N_11400);
xnor U12993 (N_12993,N_11888,N_12160);
nand U12994 (N_12994,N_11532,N_11537);
and U12995 (N_12995,N_12407,N_11473);
and U12996 (N_12996,N_12437,N_11336);
or U12997 (N_12997,N_12094,N_11728);
nand U12998 (N_12998,N_11682,N_11456);
and U12999 (N_12999,N_12253,N_11667);
nor U13000 (N_13000,N_12268,N_12436);
nand U13001 (N_13001,N_12230,N_11692);
and U13002 (N_13002,N_12128,N_11850);
nor U13003 (N_13003,N_12334,N_11262);
nand U13004 (N_13004,N_12354,N_11580);
nand U13005 (N_13005,N_12390,N_12108);
or U13006 (N_13006,N_11511,N_11787);
nor U13007 (N_13007,N_12488,N_12274);
or U13008 (N_13008,N_12205,N_11416);
nor U13009 (N_13009,N_11675,N_11965);
or U13010 (N_13010,N_11376,N_12330);
or U13011 (N_13011,N_11931,N_12052);
xor U13012 (N_13012,N_11372,N_11671);
nor U13013 (N_13013,N_11370,N_12456);
nor U13014 (N_13014,N_12259,N_11867);
xor U13015 (N_13015,N_11483,N_11848);
nand U13016 (N_13016,N_11814,N_12129);
nand U13017 (N_13017,N_11760,N_11339);
or U13018 (N_13018,N_12227,N_11476);
nand U13019 (N_13019,N_11401,N_12057);
nor U13020 (N_13020,N_11624,N_12104);
nor U13021 (N_13021,N_11347,N_11297);
and U13022 (N_13022,N_11873,N_11894);
nor U13023 (N_13023,N_12449,N_12059);
and U13024 (N_13024,N_12321,N_12411);
nand U13025 (N_13025,N_12117,N_12240);
nor U13026 (N_13026,N_12162,N_12313);
and U13027 (N_13027,N_12326,N_11831);
or U13028 (N_13028,N_11556,N_12034);
nand U13029 (N_13029,N_12217,N_12366);
xor U13030 (N_13030,N_11455,N_11797);
nand U13031 (N_13031,N_11663,N_11432);
nor U13032 (N_13032,N_12171,N_12114);
nor U13033 (N_13033,N_11811,N_11509);
nor U13034 (N_13034,N_11765,N_11611);
xnor U13035 (N_13035,N_11696,N_11353);
nand U13036 (N_13036,N_11499,N_11612);
or U13037 (N_13037,N_12000,N_11651);
or U13038 (N_13038,N_11761,N_11281);
nor U13039 (N_13039,N_12289,N_11304);
or U13040 (N_13040,N_12121,N_12028);
or U13041 (N_13041,N_11925,N_12278);
or U13042 (N_13042,N_12344,N_12065);
nor U13043 (N_13043,N_11982,N_12231);
and U13044 (N_13044,N_12430,N_11701);
and U13045 (N_13045,N_11342,N_11764);
nand U13046 (N_13046,N_12461,N_12154);
nand U13047 (N_13047,N_12315,N_11591);
nand U13048 (N_13048,N_12075,N_12235);
nor U13049 (N_13049,N_11861,N_12319);
nand U13050 (N_13050,N_11706,N_11680);
xor U13051 (N_13051,N_11468,N_12203);
nor U13052 (N_13052,N_11876,N_11396);
nand U13053 (N_13053,N_12143,N_12255);
xor U13054 (N_13054,N_11311,N_11374);
or U13055 (N_13055,N_11581,N_11506);
nand U13056 (N_13056,N_11685,N_11291);
nor U13057 (N_13057,N_11946,N_11554);
nand U13058 (N_13058,N_12495,N_12419);
xnor U13059 (N_13059,N_11697,N_12130);
or U13060 (N_13060,N_11507,N_12441);
nand U13061 (N_13061,N_12089,N_12304);
or U13062 (N_13062,N_12416,N_11588);
xnor U13063 (N_13063,N_12460,N_12486);
or U13064 (N_13064,N_12290,N_11625);
and U13065 (N_13065,N_12453,N_11398);
and U13066 (N_13066,N_11720,N_11870);
nor U13067 (N_13067,N_12087,N_12403);
nand U13068 (N_13068,N_12320,N_12450);
nand U13069 (N_13069,N_11959,N_12347);
and U13070 (N_13070,N_12333,N_11856);
nor U13071 (N_13071,N_11391,N_11440);
nand U13072 (N_13072,N_11841,N_11344);
or U13073 (N_13073,N_11782,N_11859);
nand U13074 (N_13074,N_12413,N_11552);
nor U13075 (N_13075,N_11589,N_11847);
nand U13076 (N_13076,N_11915,N_11853);
and U13077 (N_13077,N_12353,N_11990);
xor U13078 (N_13078,N_12279,N_11869);
or U13079 (N_13079,N_11597,N_11874);
or U13080 (N_13080,N_12342,N_11960);
or U13081 (N_13081,N_12041,N_12248);
or U13082 (N_13082,N_11707,N_11379);
xor U13083 (N_13083,N_11287,N_12285);
and U13084 (N_13084,N_11417,N_11566);
or U13085 (N_13085,N_11364,N_11527);
or U13086 (N_13086,N_12337,N_12457);
xor U13087 (N_13087,N_11779,N_11450);
or U13088 (N_13088,N_11503,N_12269);
xnor U13089 (N_13089,N_11329,N_11535);
xor U13090 (N_13090,N_11258,N_11548);
and U13091 (N_13091,N_12395,N_11323);
xnor U13092 (N_13092,N_12198,N_11387);
xor U13093 (N_13093,N_12214,N_12410);
nor U13094 (N_13094,N_12314,N_12073);
nor U13095 (N_13095,N_11521,N_11739);
nand U13096 (N_13096,N_11484,N_11744);
xnor U13097 (N_13097,N_12183,N_11996);
and U13098 (N_13098,N_11973,N_11916);
nand U13099 (N_13099,N_12343,N_11702);
or U13100 (N_13100,N_11510,N_12061);
and U13101 (N_13101,N_11534,N_12464);
xnor U13102 (N_13102,N_12072,N_11711);
or U13103 (N_13103,N_12401,N_11328);
nor U13104 (N_13104,N_11457,N_12054);
nor U13105 (N_13105,N_11804,N_12444);
or U13106 (N_13106,N_11628,N_11404);
or U13107 (N_13107,N_12018,N_12058);
xor U13108 (N_13108,N_12175,N_11791);
and U13109 (N_13109,N_11289,N_12254);
nor U13110 (N_13110,N_12239,N_11546);
nand U13111 (N_13111,N_12323,N_12247);
nand U13112 (N_13112,N_12210,N_11477);
and U13113 (N_13113,N_12384,N_12142);
nand U13114 (N_13114,N_11751,N_11932);
nor U13115 (N_13115,N_11354,N_11824);
xor U13116 (N_13116,N_11314,N_12277);
or U13117 (N_13117,N_11254,N_11614);
nor U13118 (N_13118,N_11598,N_11716);
and U13119 (N_13119,N_12016,N_11921);
or U13120 (N_13120,N_11679,N_11657);
nand U13121 (N_13121,N_11723,N_11349);
xor U13122 (N_13122,N_12055,N_12159);
and U13123 (N_13123,N_12226,N_12427);
xnor U13124 (N_13124,N_12030,N_11766);
xor U13125 (N_13125,N_11549,N_11641);
xor U13126 (N_13126,N_12248,N_11475);
nand U13127 (N_13127,N_12058,N_12043);
nor U13128 (N_13128,N_11730,N_12203);
or U13129 (N_13129,N_11621,N_11582);
xnor U13130 (N_13130,N_12424,N_11897);
xnor U13131 (N_13131,N_12016,N_11950);
xnor U13132 (N_13132,N_11289,N_12285);
or U13133 (N_13133,N_11342,N_11485);
nor U13134 (N_13134,N_12308,N_11947);
nor U13135 (N_13135,N_12403,N_11404);
nor U13136 (N_13136,N_12195,N_11318);
or U13137 (N_13137,N_12499,N_11926);
and U13138 (N_13138,N_12427,N_11984);
nand U13139 (N_13139,N_12210,N_12486);
and U13140 (N_13140,N_11676,N_12428);
nor U13141 (N_13141,N_12221,N_11252);
and U13142 (N_13142,N_11343,N_11734);
xnor U13143 (N_13143,N_11846,N_11926);
xnor U13144 (N_13144,N_12058,N_11982);
xor U13145 (N_13145,N_11836,N_11587);
nor U13146 (N_13146,N_11906,N_11489);
xnor U13147 (N_13147,N_11592,N_11968);
nor U13148 (N_13148,N_11344,N_12108);
nand U13149 (N_13149,N_12284,N_11324);
nand U13150 (N_13150,N_11822,N_11888);
nand U13151 (N_13151,N_11265,N_11478);
and U13152 (N_13152,N_11273,N_11801);
and U13153 (N_13153,N_11406,N_12467);
or U13154 (N_13154,N_12129,N_11860);
nor U13155 (N_13155,N_12324,N_11361);
xnor U13156 (N_13156,N_11502,N_11744);
nand U13157 (N_13157,N_11866,N_11703);
and U13158 (N_13158,N_11805,N_11490);
or U13159 (N_13159,N_11934,N_11489);
and U13160 (N_13160,N_11304,N_11371);
nor U13161 (N_13161,N_12395,N_12162);
nand U13162 (N_13162,N_11674,N_11928);
nor U13163 (N_13163,N_11750,N_11880);
xor U13164 (N_13164,N_11370,N_11471);
xnor U13165 (N_13165,N_11984,N_12315);
nor U13166 (N_13166,N_12028,N_11425);
nand U13167 (N_13167,N_11717,N_11639);
nor U13168 (N_13168,N_12486,N_12396);
and U13169 (N_13169,N_11829,N_12060);
or U13170 (N_13170,N_11412,N_11601);
and U13171 (N_13171,N_12024,N_12172);
xor U13172 (N_13172,N_11608,N_11930);
and U13173 (N_13173,N_11982,N_12083);
xor U13174 (N_13174,N_12270,N_12485);
and U13175 (N_13175,N_11579,N_12276);
nor U13176 (N_13176,N_12379,N_11616);
xor U13177 (N_13177,N_11659,N_11358);
nand U13178 (N_13178,N_11701,N_11439);
nand U13179 (N_13179,N_12332,N_12083);
nand U13180 (N_13180,N_11842,N_11314);
nand U13181 (N_13181,N_12437,N_11988);
xnor U13182 (N_13182,N_11594,N_11984);
xor U13183 (N_13183,N_11978,N_12429);
nor U13184 (N_13184,N_11745,N_11897);
and U13185 (N_13185,N_11631,N_11481);
nand U13186 (N_13186,N_11979,N_11839);
or U13187 (N_13187,N_12377,N_12265);
nand U13188 (N_13188,N_12406,N_11290);
and U13189 (N_13189,N_12109,N_11332);
nor U13190 (N_13190,N_12053,N_12160);
xnor U13191 (N_13191,N_11367,N_11338);
nor U13192 (N_13192,N_11532,N_11906);
xor U13193 (N_13193,N_11755,N_12359);
xnor U13194 (N_13194,N_11927,N_12218);
xor U13195 (N_13195,N_12144,N_12329);
xor U13196 (N_13196,N_11646,N_12277);
or U13197 (N_13197,N_11546,N_11584);
nor U13198 (N_13198,N_11686,N_12330);
nor U13199 (N_13199,N_12198,N_11508);
or U13200 (N_13200,N_11270,N_12315);
nand U13201 (N_13201,N_12475,N_12250);
or U13202 (N_13202,N_11756,N_12423);
xor U13203 (N_13203,N_12184,N_11849);
nand U13204 (N_13204,N_11564,N_12438);
or U13205 (N_13205,N_11774,N_11351);
or U13206 (N_13206,N_11861,N_12096);
and U13207 (N_13207,N_12063,N_11492);
and U13208 (N_13208,N_12395,N_11892);
nand U13209 (N_13209,N_12445,N_11366);
nand U13210 (N_13210,N_11605,N_12319);
nor U13211 (N_13211,N_12086,N_12008);
nor U13212 (N_13212,N_12171,N_11804);
and U13213 (N_13213,N_11282,N_11552);
or U13214 (N_13214,N_11636,N_11879);
or U13215 (N_13215,N_11983,N_11604);
nor U13216 (N_13216,N_11599,N_11340);
or U13217 (N_13217,N_12339,N_12413);
nand U13218 (N_13218,N_11821,N_11415);
or U13219 (N_13219,N_12040,N_11750);
or U13220 (N_13220,N_12483,N_11960);
nor U13221 (N_13221,N_12073,N_12333);
and U13222 (N_13222,N_11944,N_11955);
nand U13223 (N_13223,N_11324,N_11271);
nand U13224 (N_13224,N_11764,N_11265);
or U13225 (N_13225,N_11992,N_12343);
nand U13226 (N_13226,N_11740,N_11608);
and U13227 (N_13227,N_12434,N_11661);
or U13228 (N_13228,N_11897,N_11341);
xnor U13229 (N_13229,N_11564,N_11861);
nor U13230 (N_13230,N_12388,N_12172);
and U13231 (N_13231,N_12425,N_11385);
and U13232 (N_13232,N_11309,N_12397);
xnor U13233 (N_13233,N_12477,N_12401);
nand U13234 (N_13234,N_11783,N_11861);
nor U13235 (N_13235,N_11856,N_12430);
nor U13236 (N_13236,N_12367,N_12422);
xor U13237 (N_13237,N_11744,N_12348);
nand U13238 (N_13238,N_11843,N_11329);
nand U13239 (N_13239,N_11801,N_12014);
xnor U13240 (N_13240,N_11804,N_11908);
and U13241 (N_13241,N_11685,N_11470);
or U13242 (N_13242,N_12004,N_11779);
nor U13243 (N_13243,N_12451,N_11887);
and U13244 (N_13244,N_11659,N_12088);
and U13245 (N_13245,N_11418,N_11952);
and U13246 (N_13246,N_12349,N_11566);
nor U13247 (N_13247,N_12253,N_12133);
nor U13248 (N_13248,N_11485,N_11857);
nand U13249 (N_13249,N_11939,N_11995);
nor U13250 (N_13250,N_12015,N_12165);
nand U13251 (N_13251,N_11867,N_11442);
nor U13252 (N_13252,N_11884,N_11434);
xnor U13253 (N_13253,N_11823,N_11959);
or U13254 (N_13254,N_11996,N_11850);
nor U13255 (N_13255,N_11846,N_12380);
and U13256 (N_13256,N_11718,N_11874);
nor U13257 (N_13257,N_11419,N_11677);
nor U13258 (N_13258,N_11954,N_12317);
and U13259 (N_13259,N_12223,N_12108);
or U13260 (N_13260,N_12109,N_12309);
nand U13261 (N_13261,N_11606,N_11761);
nand U13262 (N_13262,N_12192,N_12491);
or U13263 (N_13263,N_11474,N_12375);
nor U13264 (N_13264,N_12367,N_11359);
or U13265 (N_13265,N_12196,N_12001);
nand U13266 (N_13266,N_12251,N_11782);
or U13267 (N_13267,N_11311,N_11317);
or U13268 (N_13268,N_11987,N_12435);
or U13269 (N_13269,N_11484,N_11930);
and U13270 (N_13270,N_12110,N_11948);
xor U13271 (N_13271,N_11315,N_11876);
xor U13272 (N_13272,N_12393,N_11649);
nand U13273 (N_13273,N_11908,N_11675);
and U13274 (N_13274,N_12185,N_11874);
xor U13275 (N_13275,N_11643,N_11650);
nor U13276 (N_13276,N_11868,N_12076);
or U13277 (N_13277,N_12260,N_11760);
and U13278 (N_13278,N_11508,N_11661);
xnor U13279 (N_13279,N_12490,N_11887);
nor U13280 (N_13280,N_12472,N_11456);
or U13281 (N_13281,N_11465,N_11413);
nor U13282 (N_13282,N_11378,N_11893);
xnor U13283 (N_13283,N_12365,N_11319);
nor U13284 (N_13284,N_11978,N_12265);
or U13285 (N_13285,N_12113,N_12293);
or U13286 (N_13286,N_11320,N_11992);
nor U13287 (N_13287,N_11764,N_12124);
nand U13288 (N_13288,N_12012,N_12169);
nand U13289 (N_13289,N_11351,N_12366);
or U13290 (N_13290,N_12367,N_11486);
or U13291 (N_13291,N_11627,N_12327);
nor U13292 (N_13292,N_11938,N_12450);
xor U13293 (N_13293,N_12140,N_12189);
or U13294 (N_13294,N_11259,N_12384);
nor U13295 (N_13295,N_12133,N_11922);
nand U13296 (N_13296,N_12390,N_12367);
or U13297 (N_13297,N_12206,N_11800);
xnor U13298 (N_13298,N_12390,N_11796);
xnor U13299 (N_13299,N_11494,N_11771);
nor U13300 (N_13300,N_12240,N_11631);
xor U13301 (N_13301,N_11988,N_12252);
or U13302 (N_13302,N_12325,N_12305);
nand U13303 (N_13303,N_11999,N_11778);
and U13304 (N_13304,N_11651,N_12324);
nor U13305 (N_13305,N_11406,N_11385);
nor U13306 (N_13306,N_12362,N_12203);
nand U13307 (N_13307,N_11689,N_11446);
or U13308 (N_13308,N_11778,N_11392);
or U13309 (N_13309,N_12493,N_11849);
and U13310 (N_13310,N_11262,N_11900);
nand U13311 (N_13311,N_11311,N_12203);
nand U13312 (N_13312,N_11657,N_12494);
or U13313 (N_13313,N_12235,N_12244);
xor U13314 (N_13314,N_11451,N_12129);
xor U13315 (N_13315,N_11377,N_11339);
xor U13316 (N_13316,N_12427,N_12280);
and U13317 (N_13317,N_11939,N_11297);
xor U13318 (N_13318,N_11806,N_12339);
xor U13319 (N_13319,N_12497,N_12391);
nand U13320 (N_13320,N_12462,N_12093);
xor U13321 (N_13321,N_11654,N_11651);
or U13322 (N_13322,N_11612,N_12230);
and U13323 (N_13323,N_11608,N_11875);
or U13324 (N_13324,N_11917,N_11971);
xor U13325 (N_13325,N_11835,N_11745);
nand U13326 (N_13326,N_12270,N_11993);
nand U13327 (N_13327,N_12096,N_12413);
nor U13328 (N_13328,N_12059,N_12078);
xnor U13329 (N_13329,N_12494,N_12078);
nor U13330 (N_13330,N_12359,N_11855);
nor U13331 (N_13331,N_11951,N_11881);
xnor U13332 (N_13332,N_11689,N_12337);
and U13333 (N_13333,N_12462,N_11832);
or U13334 (N_13334,N_12050,N_11275);
xnor U13335 (N_13335,N_12039,N_12270);
nand U13336 (N_13336,N_11574,N_12059);
xor U13337 (N_13337,N_12290,N_12215);
nor U13338 (N_13338,N_12401,N_11826);
xnor U13339 (N_13339,N_11853,N_11687);
nand U13340 (N_13340,N_11362,N_11985);
xor U13341 (N_13341,N_11925,N_11439);
xor U13342 (N_13342,N_11857,N_11440);
or U13343 (N_13343,N_11722,N_11746);
or U13344 (N_13344,N_11724,N_11771);
xnor U13345 (N_13345,N_11739,N_12052);
or U13346 (N_13346,N_12136,N_12152);
xor U13347 (N_13347,N_12035,N_12045);
or U13348 (N_13348,N_12104,N_11931);
nor U13349 (N_13349,N_12471,N_11714);
and U13350 (N_13350,N_12425,N_12006);
xnor U13351 (N_13351,N_11605,N_11284);
and U13352 (N_13352,N_12481,N_11436);
nand U13353 (N_13353,N_12204,N_11665);
nand U13354 (N_13354,N_12223,N_12449);
xor U13355 (N_13355,N_11639,N_11560);
xor U13356 (N_13356,N_11966,N_12474);
nor U13357 (N_13357,N_12198,N_11859);
nand U13358 (N_13358,N_11684,N_11709);
nand U13359 (N_13359,N_12146,N_11964);
or U13360 (N_13360,N_11770,N_11929);
and U13361 (N_13361,N_11424,N_11472);
or U13362 (N_13362,N_11914,N_11723);
and U13363 (N_13363,N_11883,N_12366);
and U13364 (N_13364,N_12276,N_11403);
and U13365 (N_13365,N_11945,N_11881);
and U13366 (N_13366,N_12440,N_11938);
and U13367 (N_13367,N_11714,N_11378);
nor U13368 (N_13368,N_12302,N_12058);
xor U13369 (N_13369,N_11878,N_11263);
nand U13370 (N_13370,N_11686,N_12112);
and U13371 (N_13371,N_11265,N_12232);
nand U13372 (N_13372,N_11642,N_12354);
or U13373 (N_13373,N_11441,N_11658);
and U13374 (N_13374,N_12421,N_11980);
nor U13375 (N_13375,N_11767,N_11759);
or U13376 (N_13376,N_11610,N_11784);
nor U13377 (N_13377,N_11444,N_12480);
or U13378 (N_13378,N_11783,N_11335);
and U13379 (N_13379,N_11340,N_12446);
or U13380 (N_13380,N_11696,N_11610);
and U13381 (N_13381,N_11420,N_12126);
and U13382 (N_13382,N_11412,N_11914);
nand U13383 (N_13383,N_11766,N_11385);
nand U13384 (N_13384,N_11818,N_11627);
nand U13385 (N_13385,N_11749,N_12310);
nor U13386 (N_13386,N_11890,N_11394);
nand U13387 (N_13387,N_11838,N_12135);
nand U13388 (N_13388,N_11872,N_11783);
or U13389 (N_13389,N_11818,N_12055);
xnor U13390 (N_13390,N_11686,N_11888);
nand U13391 (N_13391,N_12068,N_12100);
nand U13392 (N_13392,N_11904,N_11294);
nand U13393 (N_13393,N_11720,N_12144);
or U13394 (N_13394,N_11635,N_12069);
nor U13395 (N_13395,N_11422,N_12451);
xor U13396 (N_13396,N_11666,N_12351);
nor U13397 (N_13397,N_11821,N_11880);
xor U13398 (N_13398,N_11346,N_11484);
xnor U13399 (N_13399,N_11722,N_11379);
nand U13400 (N_13400,N_11369,N_11349);
nand U13401 (N_13401,N_11717,N_11524);
nand U13402 (N_13402,N_11483,N_12035);
xnor U13403 (N_13403,N_11493,N_11905);
xnor U13404 (N_13404,N_12206,N_12221);
xnor U13405 (N_13405,N_11831,N_12002);
nand U13406 (N_13406,N_12052,N_12232);
or U13407 (N_13407,N_11725,N_11862);
and U13408 (N_13408,N_11760,N_12450);
or U13409 (N_13409,N_11835,N_11468);
nand U13410 (N_13410,N_12220,N_12324);
nand U13411 (N_13411,N_11504,N_11569);
xnor U13412 (N_13412,N_12467,N_11583);
xor U13413 (N_13413,N_11473,N_12301);
nor U13414 (N_13414,N_11669,N_12447);
nand U13415 (N_13415,N_11293,N_11535);
or U13416 (N_13416,N_11611,N_11785);
nand U13417 (N_13417,N_12472,N_11790);
nor U13418 (N_13418,N_11258,N_11283);
xnor U13419 (N_13419,N_11699,N_11716);
or U13420 (N_13420,N_11385,N_11895);
or U13421 (N_13421,N_11270,N_12230);
nand U13422 (N_13422,N_12076,N_11459);
nand U13423 (N_13423,N_12297,N_12281);
nor U13424 (N_13424,N_12452,N_12114);
nand U13425 (N_13425,N_12263,N_11681);
nand U13426 (N_13426,N_12002,N_12360);
nor U13427 (N_13427,N_11905,N_11900);
and U13428 (N_13428,N_12378,N_11731);
or U13429 (N_13429,N_12472,N_12440);
xnor U13430 (N_13430,N_11723,N_11870);
xor U13431 (N_13431,N_12201,N_12249);
nor U13432 (N_13432,N_12390,N_11795);
or U13433 (N_13433,N_11516,N_11426);
nor U13434 (N_13434,N_11788,N_11843);
nor U13435 (N_13435,N_11567,N_11324);
or U13436 (N_13436,N_11317,N_12409);
and U13437 (N_13437,N_11952,N_12455);
nor U13438 (N_13438,N_11305,N_11912);
xor U13439 (N_13439,N_11942,N_11340);
and U13440 (N_13440,N_11970,N_12347);
or U13441 (N_13441,N_11826,N_11587);
or U13442 (N_13442,N_11945,N_11805);
xnor U13443 (N_13443,N_12161,N_11583);
nor U13444 (N_13444,N_11927,N_11322);
nor U13445 (N_13445,N_12014,N_11518);
and U13446 (N_13446,N_12064,N_12428);
or U13447 (N_13447,N_12333,N_12497);
and U13448 (N_13448,N_12087,N_12213);
nand U13449 (N_13449,N_11642,N_12182);
xor U13450 (N_13450,N_11463,N_12066);
or U13451 (N_13451,N_11785,N_11844);
xor U13452 (N_13452,N_12487,N_12069);
and U13453 (N_13453,N_11652,N_11893);
and U13454 (N_13454,N_11477,N_11786);
nor U13455 (N_13455,N_11565,N_11264);
nor U13456 (N_13456,N_11455,N_11716);
nor U13457 (N_13457,N_11752,N_11888);
nand U13458 (N_13458,N_12466,N_12385);
or U13459 (N_13459,N_11524,N_11676);
xor U13460 (N_13460,N_11555,N_11363);
nor U13461 (N_13461,N_11970,N_11993);
nor U13462 (N_13462,N_12006,N_11420);
xor U13463 (N_13463,N_11837,N_11932);
or U13464 (N_13464,N_11797,N_11390);
nand U13465 (N_13465,N_11912,N_11485);
nor U13466 (N_13466,N_12364,N_12192);
and U13467 (N_13467,N_12148,N_11926);
nand U13468 (N_13468,N_11966,N_12114);
and U13469 (N_13469,N_12486,N_11785);
or U13470 (N_13470,N_12219,N_11988);
nand U13471 (N_13471,N_12100,N_11259);
xnor U13472 (N_13472,N_12476,N_11376);
nand U13473 (N_13473,N_12161,N_11596);
nand U13474 (N_13474,N_11364,N_12281);
xor U13475 (N_13475,N_11961,N_12472);
and U13476 (N_13476,N_11980,N_11532);
xor U13477 (N_13477,N_11628,N_11860);
nor U13478 (N_13478,N_11272,N_11801);
nand U13479 (N_13479,N_12001,N_11519);
xnor U13480 (N_13480,N_12432,N_11854);
and U13481 (N_13481,N_11811,N_12388);
and U13482 (N_13482,N_11811,N_11943);
or U13483 (N_13483,N_11777,N_11813);
and U13484 (N_13484,N_11257,N_12066);
nor U13485 (N_13485,N_11602,N_11954);
and U13486 (N_13486,N_12069,N_12371);
and U13487 (N_13487,N_11553,N_12184);
nor U13488 (N_13488,N_11403,N_12169);
nand U13489 (N_13489,N_12252,N_11450);
nand U13490 (N_13490,N_11841,N_11297);
xor U13491 (N_13491,N_11930,N_11850);
nand U13492 (N_13492,N_12468,N_12191);
xor U13493 (N_13493,N_11448,N_11968);
nand U13494 (N_13494,N_12216,N_12442);
xnor U13495 (N_13495,N_12345,N_11543);
xnor U13496 (N_13496,N_11259,N_11276);
xor U13497 (N_13497,N_11751,N_11404);
nand U13498 (N_13498,N_11658,N_12149);
xnor U13499 (N_13499,N_11681,N_11614);
xor U13500 (N_13500,N_11652,N_12268);
xor U13501 (N_13501,N_12404,N_11621);
and U13502 (N_13502,N_11702,N_11902);
xnor U13503 (N_13503,N_11940,N_11826);
and U13504 (N_13504,N_11395,N_11845);
xnor U13505 (N_13505,N_12132,N_11739);
nand U13506 (N_13506,N_11298,N_11627);
and U13507 (N_13507,N_11272,N_11975);
or U13508 (N_13508,N_11580,N_12009);
xor U13509 (N_13509,N_11559,N_11785);
or U13510 (N_13510,N_12374,N_11854);
nor U13511 (N_13511,N_11575,N_12275);
or U13512 (N_13512,N_11697,N_12154);
and U13513 (N_13513,N_12272,N_11521);
xnor U13514 (N_13514,N_11808,N_11798);
or U13515 (N_13515,N_12277,N_12324);
nand U13516 (N_13516,N_11605,N_11804);
and U13517 (N_13517,N_11431,N_12036);
nand U13518 (N_13518,N_11561,N_12138);
nand U13519 (N_13519,N_12212,N_12159);
and U13520 (N_13520,N_11619,N_12263);
or U13521 (N_13521,N_12020,N_12053);
nand U13522 (N_13522,N_12353,N_11337);
nor U13523 (N_13523,N_12242,N_11791);
nor U13524 (N_13524,N_12438,N_12416);
or U13525 (N_13525,N_11900,N_11471);
xnor U13526 (N_13526,N_11445,N_11841);
nor U13527 (N_13527,N_11310,N_12021);
xor U13528 (N_13528,N_11983,N_11941);
and U13529 (N_13529,N_11338,N_11427);
or U13530 (N_13530,N_11466,N_11601);
and U13531 (N_13531,N_12203,N_12092);
or U13532 (N_13532,N_12248,N_12393);
xnor U13533 (N_13533,N_11318,N_12167);
and U13534 (N_13534,N_11727,N_11975);
and U13535 (N_13535,N_12310,N_11532);
nand U13536 (N_13536,N_12210,N_12320);
and U13537 (N_13537,N_12066,N_11775);
xnor U13538 (N_13538,N_12089,N_11409);
and U13539 (N_13539,N_11274,N_11463);
and U13540 (N_13540,N_11457,N_12322);
xor U13541 (N_13541,N_11311,N_12436);
nand U13542 (N_13542,N_12129,N_12294);
or U13543 (N_13543,N_11749,N_12003);
xor U13544 (N_13544,N_11541,N_11991);
xnor U13545 (N_13545,N_11278,N_12070);
nand U13546 (N_13546,N_11377,N_12209);
nand U13547 (N_13547,N_11463,N_11742);
nor U13548 (N_13548,N_11593,N_11671);
xor U13549 (N_13549,N_12315,N_11921);
nand U13550 (N_13550,N_11551,N_11673);
nor U13551 (N_13551,N_12189,N_12499);
or U13552 (N_13552,N_12196,N_12086);
xnor U13553 (N_13553,N_11787,N_11415);
nor U13554 (N_13554,N_11920,N_11256);
or U13555 (N_13555,N_11359,N_11651);
nand U13556 (N_13556,N_11418,N_12193);
nor U13557 (N_13557,N_12197,N_11517);
xnor U13558 (N_13558,N_11929,N_12371);
xor U13559 (N_13559,N_12079,N_11891);
xnor U13560 (N_13560,N_12052,N_11827);
or U13561 (N_13561,N_11340,N_11959);
nand U13562 (N_13562,N_12480,N_11711);
and U13563 (N_13563,N_12332,N_12286);
nand U13564 (N_13564,N_12387,N_11633);
or U13565 (N_13565,N_11436,N_11838);
and U13566 (N_13566,N_12397,N_11795);
xor U13567 (N_13567,N_11968,N_12087);
xnor U13568 (N_13568,N_11294,N_11292);
xnor U13569 (N_13569,N_12322,N_12402);
nor U13570 (N_13570,N_11468,N_11679);
nor U13571 (N_13571,N_11560,N_11601);
nand U13572 (N_13572,N_12070,N_12442);
and U13573 (N_13573,N_11612,N_11919);
or U13574 (N_13574,N_11354,N_11489);
nor U13575 (N_13575,N_12261,N_12413);
xnor U13576 (N_13576,N_11489,N_11683);
nand U13577 (N_13577,N_12102,N_11802);
nor U13578 (N_13578,N_11814,N_12347);
or U13579 (N_13579,N_11308,N_11427);
nor U13580 (N_13580,N_11402,N_11821);
nand U13581 (N_13581,N_11886,N_11787);
nor U13582 (N_13582,N_12484,N_12317);
and U13583 (N_13583,N_12080,N_11476);
nand U13584 (N_13584,N_11613,N_11770);
nor U13585 (N_13585,N_11893,N_11488);
or U13586 (N_13586,N_11680,N_12306);
xor U13587 (N_13587,N_11954,N_11355);
nand U13588 (N_13588,N_11436,N_11464);
nand U13589 (N_13589,N_11711,N_12207);
and U13590 (N_13590,N_11823,N_11520);
nor U13591 (N_13591,N_11509,N_12330);
xor U13592 (N_13592,N_11634,N_12311);
nand U13593 (N_13593,N_11356,N_11627);
nor U13594 (N_13594,N_12214,N_12220);
nand U13595 (N_13595,N_11511,N_12139);
nor U13596 (N_13596,N_11394,N_12236);
or U13597 (N_13597,N_12252,N_12341);
and U13598 (N_13598,N_12280,N_11969);
and U13599 (N_13599,N_12460,N_11789);
xnor U13600 (N_13600,N_12176,N_11939);
nand U13601 (N_13601,N_12358,N_11715);
or U13602 (N_13602,N_12048,N_11385);
nor U13603 (N_13603,N_11617,N_11378);
xor U13604 (N_13604,N_11626,N_12349);
nor U13605 (N_13605,N_11873,N_12330);
and U13606 (N_13606,N_11955,N_11656);
nand U13607 (N_13607,N_12332,N_12058);
nand U13608 (N_13608,N_12036,N_11520);
and U13609 (N_13609,N_11829,N_11601);
xnor U13610 (N_13610,N_11785,N_12333);
or U13611 (N_13611,N_12063,N_11993);
or U13612 (N_13612,N_12225,N_11354);
or U13613 (N_13613,N_12350,N_11572);
xnor U13614 (N_13614,N_11380,N_12062);
xnor U13615 (N_13615,N_12008,N_12244);
and U13616 (N_13616,N_11913,N_11298);
and U13617 (N_13617,N_11708,N_12232);
or U13618 (N_13618,N_12039,N_12127);
nor U13619 (N_13619,N_11702,N_12102);
xnor U13620 (N_13620,N_11721,N_11788);
nand U13621 (N_13621,N_12451,N_11314);
nand U13622 (N_13622,N_12268,N_11524);
nor U13623 (N_13623,N_11890,N_11813);
or U13624 (N_13624,N_11765,N_11529);
and U13625 (N_13625,N_12472,N_11593);
nand U13626 (N_13626,N_11877,N_11808);
nand U13627 (N_13627,N_11772,N_12244);
nand U13628 (N_13628,N_12196,N_12464);
xnor U13629 (N_13629,N_12112,N_11294);
and U13630 (N_13630,N_12348,N_12408);
xor U13631 (N_13631,N_12092,N_11932);
nor U13632 (N_13632,N_12065,N_11342);
nor U13633 (N_13633,N_11640,N_12423);
nand U13634 (N_13634,N_11527,N_11899);
xnor U13635 (N_13635,N_12238,N_12463);
nand U13636 (N_13636,N_12322,N_12206);
nand U13637 (N_13637,N_11281,N_11905);
nand U13638 (N_13638,N_11991,N_11966);
or U13639 (N_13639,N_12051,N_12369);
nand U13640 (N_13640,N_11475,N_12120);
nor U13641 (N_13641,N_11613,N_12404);
or U13642 (N_13642,N_11821,N_12303);
xnor U13643 (N_13643,N_12094,N_11731);
nand U13644 (N_13644,N_11515,N_11877);
and U13645 (N_13645,N_11922,N_12482);
nor U13646 (N_13646,N_12067,N_12369);
nand U13647 (N_13647,N_11371,N_11830);
and U13648 (N_13648,N_12277,N_11922);
or U13649 (N_13649,N_11502,N_11782);
and U13650 (N_13650,N_11605,N_12091);
or U13651 (N_13651,N_11609,N_11419);
nand U13652 (N_13652,N_12128,N_11920);
or U13653 (N_13653,N_12338,N_11805);
xor U13654 (N_13654,N_11446,N_11814);
nand U13655 (N_13655,N_11899,N_12405);
and U13656 (N_13656,N_11858,N_11894);
nand U13657 (N_13657,N_11766,N_11719);
and U13658 (N_13658,N_12097,N_11958);
xnor U13659 (N_13659,N_12260,N_11330);
or U13660 (N_13660,N_12489,N_11318);
xor U13661 (N_13661,N_11894,N_12243);
nand U13662 (N_13662,N_11771,N_12110);
or U13663 (N_13663,N_12231,N_12389);
or U13664 (N_13664,N_12085,N_11784);
nor U13665 (N_13665,N_11389,N_12049);
and U13666 (N_13666,N_12244,N_11522);
xnor U13667 (N_13667,N_11256,N_11339);
xnor U13668 (N_13668,N_11912,N_12183);
xnor U13669 (N_13669,N_12423,N_12024);
and U13670 (N_13670,N_12237,N_11511);
nor U13671 (N_13671,N_11831,N_12238);
or U13672 (N_13672,N_12228,N_12447);
and U13673 (N_13673,N_12412,N_12037);
xor U13674 (N_13674,N_12061,N_12177);
or U13675 (N_13675,N_11449,N_12353);
or U13676 (N_13676,N_11893,N_11908);
and U13677 (N_13677,N_11423,N_11654);
nand U13678 (N_13678,N_11890,N_11883);
or U13679 (N_13679,N_12084,N_11917);
xor U13680 (N_13680,N_12476,N_11574);
nand U13681 (N_13681,N_11384,N_12258);
or U13682 (N_13682,N_11505,N_11374);
nand U13683 (N_13683,N_12464,N_12254);
xnor U13684 (N_13684,N_11833,N_11596);
xor U13685 (N_13685,N_11674,N_12446);
or U13686 (N_13686,N_11707,N_11268);
xor U13687 (N_13687,N_11810,N_12031);
and U13688 (N_13688,N_12411,N_12163);
or U13689 (N_13689,N_12427,N_11272);
and U13690 (N_13690,N_12455,N_11999);
nor U13691 (N_13691,N_11995,N_11305);
or U13692 (N_13692,N_12352,N_12396);
nor U13693 (N_13693,N_12163,N_11973);
nor U13694 (N_13694,N_12019,N_11777);
nand U13695 (N_13695,N_11411,N_11568);
nand U13696 (N_13696,N_11513,N_11622);
xor U13697 (N_13697,N_11911,N_12003);
and U13698 (N_13698,N_11471,N_11522);
nand U13699 (N_13699,N_12270,N_11641);
nand U13700 (N_13700,N_11392,N_12094);
and U13701 (N_13701,N_12102,N_12050);
or U13702 (N_13702,N_12371,N_11268);
and U13703 (N_13703,N_12173,N_11730);
nor U13704 (N_13704,N_11432,N_11581);
or U13705 (N_13705,N_12476,N_12311);
or U13706 (N_13706,N_12042,N_12207);
xnor U13707 (N_13707,N_12138,N_11933);
nor U13708 (N_13708,N_11994,N_12170);
and U13709 (N_13709,N_11598,N_11892);
or U13710 (N_13710,N_11368,N_11281);
and U13711 (N_13711,N_12383,N_12392);
nand U13712 (N_13712,N_12403,N_11751);
nor U13713 (N_13713,N_11271,N_11907);
nand U13714 (N_13714,N_11687,N_11795);
or U13715 (N_13715,N_12123,N_11495);
nand U13716 (N_13716,N_11546,N_11938);
or U13717 (N_13717,N_11599,N_12317);
nor U13718 (N_13718,N_11803,N_11665);
and U13719 (N_13719,N_11546,N_11741);
nor U13720 (N_13720,N_11577,N_12059);
xnor U13721 (N_13721,N_11812,N_11719);
xnor U13722 (N_13722,N_11677,N_11695);
or U13723 (N_13723,N_12269,N_11694);
or U13724 (N_13724,N_11608,N_12365);
xor U13725 (N_13725,N_11297,N_11680);
or U13726 (N_13726,N_11733,N_11815);
nand U13727 (N_13727,N_12427,N_11691);
nor U13728 (N_13728,N_11355,N_11416);
nor U13729 (N_13729,N_12413,N_12265);
nand U13730 (N_13730,N_11375,N_11746);
and U13731 (N_13731,N_11738,N_12437);
and U13732 (N_13732,N_11720,N_11688);
xor U13733 (N_13733,N_11272,N_11619);
nor U13734 (N_13734,N_12364,N_12419);
and U13735 (N_13735,N_12018,N_11835);
and U13736 (N_13736,N_11723,N_11755);
and U13737 (N_13737,N_12133,N_11632);
nor U13738 (N_13738,N_11321,N_11676);
and U13739 (N_13739,N_12341,N_11307);
and U13740 (N_13740,N_11485,N_11418);
xnor U13741 (N_13741,N_11350,N_11874);
xor U13742 (N_13742,N_11734,N_11991);
nor U13743 (N_13743,N_11434,N_11999);
or U13744 (N_13744,N_12102,N_11682);
xor U13745 (N_13745,N_12461,N_12153);
or U13746 (N_13746,N_11966,N_11370);
xor U13747 (N_13747,N_11868,N_11349);
or U13748 (N_13748,N_11849,N_11700);
xnor U13749 (N_13749,N_12320,N_12100);
or U13750 (N_13750,N_12744,N_13626);
nor U13751 (N_13751,N_13159,N_13725);
nand U13752 (N_13752,N_12601,N_13132);
xnor U13753 (N_13753,N_13104,N_12922);
xnor U13754 (N_13754,N_12812,N_12931);
nor U13755 (N_13755,N_13405,N_12898);
nor U13756 (N_13756,N_13459,N_12533);
nor U13757 (N_13757,N_13627,N_13361);
nand U13758 (N_13758,N_12924,N_12659);
nor U13759 (N_13759,N_13697,N_12614);
nor U13760 (N_13760,N_12865,N_13449);
nand U13761 (N_13761,N_13732,N_13658);
nand U13762 (N_13762,N_13582,N_13069);
nor U13763 (N_13763,N_13356,N_13407);
xor U13764 (N_13764,N_12799,N_12937);
nand U13765 (N_13765,N_13207,N_13044);
or U13766 (N_13766,N_12768,N_12581);
nor U13767 (N_13767,N_13527,N_13063);
xnor U13768 (N_13768,N_12873,N_13475);
xor U13769 (N_13769,N_12693,N_12883);
and U13770 (N_13770,N_13078,N_12523);
and U13771 (N_13771,N_13244,N_12594);
or U13772 (N_13772,N_13483,N_12616);
or U13773 (N_13773,N_12964,N_12961);
or U13774 (N_13774,N_13480,N_13260);
and U13775 (N_13775,N_13030,N_12675);
and U13776 (N_13776,N_13665,N_12847);
and U13777 (N_13777,N_12682,N_12950);
and U13778 (N_13778,N_13437,N_12608);
nand U13779 (N_13779,N_12963,N_13341);
or U13780 (N_13780,N_12633,N_13070);
nand U13781 (N_13781,N_12947,N_13301);
xor U13782 (N_13782,N_12597,N_12997);
or U13783 (N_13783,N_12665,N_12926);
xnor U13784 (N_13784,N_13233,N_13007);
and U13785 (N_13785,N_13579,N_12936);
xor U13786 (N_13786,N_13742,N_13517);
and U13787 (N_13787,N_13254,N_12554);
nand U13788 (N_13788,N_13488,N_13531);
or U13789 (N_13789,N_13592,N_12881);
nor U13790 (N_13790,N_12838,N_12876);
xnor U13791 (N_13791,N_12986,N_13614);
xor U13792 (N_13792,N_12816,N_13027);
and U13793 (N_13793,N_13525,N_13662);
or U13794 (N_13794,N_12823,N_13102);
nand U13795 (N_13795,N_13564,N_13438);
nor U13796 (N_13796,N_13738,N_13261);
nand U13797 (N_13797,N_13304,N_13682);
and U13798 (N_13798,N_12643,N_12697);
nor U13799 (N_13799,N_13045,N_13546);
nor U13800 (N_13800,N_13289,N_13644);
nor U13801 (N_13801,N_12804,N_12655);
nand U13802 (N_13802,N_12989,N_13451);
xor U13803 (N_13803,N_13000,N_13171);
nor U13804 (N_13804,N_12730,N_13013);
or U13805 (N_13805,N_13043,N_13089);
and U13806 (N_13806,N_12741,N_13436);
xnor U13807 (N_13807,N_13079,N_12746);
or U13808 (N_13808,N_13467,N_13619);
xnor U13809 (N_13809,N_12854,N_13705);
and U13810 (N_13810,N_12801,N_13332);
or U13811 (N_13811,N_13290,N_12543);
and U13812 (N_13812,N_12946,N_13291);
or U13813 (N_13813,N_13190,N_12637);
or U13814 (N_13814,N_12545,N_12830);
nor U13815 (N_13815,N_13319,N_13298);
or U13816 (N_13816,N_12651,N_13688);
or U13817 (N_13817,N_13059,N_13121);
and U13818 (N_13818,N_12559,N_13417);
nor U13819 (N_13819,N_13421,N_13106);
or U13820 (N_13820,N_13635,N_12953);
nand U13821 (N_13821,N_12681,N_13181);
nand U13822 (N_13822,N_12713,N_12716);
or U13823 (N_13823,N_12930,N_13153);
nand U13824 (N_13824,N_13501,N_13601);
or U13825 (N_13825,N_12751,N_13607);
or U13826 (N_13826,N_12564,N_13033);
or U13827 (N_13827,N_13606,N_12829);
nand U13828 (N_13828,N_12699,N_13350);
and U13829 (N_13829,N_12837,N_12618);
or U13830 (N_13830,N_13378,N_13279);
xnor U13831 (N_13831,N_13504,N_12894);
xor U13832 (N_13832,N_13015,N_12563);
nor U13833 (N_13833,N_12982,N_13684);
xor U13834 (N_13834,N_13236,N_12561);
and U13835 (N_13835,N_13162,N_12504);
xor U13836 (N_13836,N_12756,N_13408);
or U13837 (N_13837,N_13391,N_12776);
nand U13838 (N_13838,N_13225,N_12864);
nand U13839 (N_13839,N_13492,N_12539);
nor U13840 (N_13840,N_13482,N_13180);
or U13841 (N_13841,N_13074,N_13404);
and U13842 (N_13842,N_13274,N_12737);
or U13843 (N_13843,N_12785,N_12720);
and U13844 (N_13844,N_12732,N_13556);
nand U13845 (N_13845,N_12705,N_13557);
nor U13846 (N_13846,N_12727,N_13383);
xnor U13847 (N_13847,N_13381,N_13183);
xor U13848 (N_13848,N_12506,N_13499);
or U13849 (N_13849,N_13166,N_13511);
nand U13850 (N_13850,N_12870,N_13072);
or U13851 (N_13851,N_12646,N_13731);
xor U13852 (N_13852,N_12770,N_13710);
nand U13853 (N_13853,N_13285,N_12587);
nand U13854 (N_13854,N_13338,N_12755);
nand U13855 (N_13855,N_13217,N_12516);
or U13856 (N_13856,N_13318,N_13232);
xnor U13857 (N_13857,N_13354,N_13562);
nor U13858 (N_13858,N_13555,N_12688);
or U13859 (N_13859,N_13567,N_12548);
or U13860 (N_13860,N_13672,N_12576);
xor U13861 (N_13861,N_13359,N_12684);
or U13862 (N_13862,N_13680,N_12769);
nor U13863 (N_13863,N_13143,N_13222);
nor U13864 (N_13864,N_12531,N_12942);
or U13865 (N_13865,N_13196,N_12957);
xnor U13866 (N_13866,N_13311,N_13523);
and U13867 (N_13867,N_13263,N_13170);
and U13868 (N_13868,N_13726,N_13513);
nor U13869 (N_13869,N_12851,N_13657);
nand U13870 (N_13870,N_13435,N_13390);
nand U13871 (N_13871,N_13655,N_13639);
nand U13872 (N_13872,N_12540,N_13453);
and U13873 (N_13873,N_13594,N_13495);
nand U13874 (N_13874,N_13653,N_13117);
or U13875 (N_13875,N_13073,N_12690);
or U13876 (N_13876,N_13179,N_13270);
xnor U13877 (N_13877,N_12856,N_12983);
nor U13878 (N_13878,N_13317,N_13518);
or U13879 (N_13879,N_13266,N_12871);
xor U13880 (N_13880,N_13092,N_13347);
and U13881 (N_13881,N_13194,N_12609);
nor U13882 (N_13882,N_12954,N_12800);
nor U13883 (N_13883,N_13123,N_12869);
xnor U13884 (N_13884,N_13004,N_12825);
nand U13885 (N_13885,N_13508,N_13049);
and U13886 (N_13886,N_12968,N_12604);
nand U13887 (N_13887,N_13510,N_13091);
nor U13888 (N_13888,N_12918,N_12939);
xnor U13889 (N_13889,N_12753,N_12839);
and U13890 (N_13890,N_12951,N_13188);
nor U13891 (N_13891,N_12912,N_12915);
and U13892 (N_13892,N_12975,N_12831);
and U13893 (N_13893,N_13571,N_13110);
xor U13894 (N_13894,N_12658,N_13704);
xnor U13895 (N_13895,N_13160,N_13479);
xnor U13896 (N_13896,N_13745,N_13551);
nand U13897 (N_13897,N_12927,N_13723);
or U13898 (N_13898,N_12923,N_13315);
nand U13899 (N_13899,N_13258,N_13071);
or U13900 (N_13900,N_13292,N_12731);
and U13901 (N_13901,N_12575,N_13740);
xnor U13902 (N_13902,N_13568,N_13549);
or U13903 (N_13903,N_13450,N_13014);
nand U13904 (N_13904,N_13692,N_12878);
and U13905 (N_13905,N_13215,N_13563);
nor U13906 (N_13906,N_13409,N_13721);
or U13907 (N_13907,N_12844,N_12525);
nand U13908 (N_13908,N_12696,N_13604);
and U13909 (N_13909,N_12882,N_12537);
xor U13910 (N_13910,N_13623,N_13161);
or U13911 (N_13911,N_13415,N_12771);
or U13912 (N_13912,N_12893,N_13313);
nor U13913 (N_13913,N_13191,N_12635);
and U13914 (N_13914,N_12965,N_12528);
nand U13915 (N_13915,N_13135,N_12875);
and U13916 (N_13916,N_13701,N_13558);
nor U13917 (N_13917,N_12952,N_13309);
xor U13918 (N_13918,N_13681,N_12657);
and U13919 (N_13919,N_13220,N_13545);
and U13920 (N_13920,N_12821,N_13139);
and U13921 (N_13921,N_13445,N_13703);
xnor U13922 (N_13922,N_13661,N_13651);
or U13923 (N_13923,N_12556,N_13142);
xnor U13924 (N_13924,N_13533,N_13320);
and U13925 (N_13925,N_13476,N_13018);
xor U13926 (N_13926,N_13020,N_13214);
nand U13927 (N_13927,N_13137,N_13282);
nor U13928 (N_13928,N_12920,N_12670);
or U13929 (N_13929,N_13719,N_13148);
nor U13930 (N_13930,N_12943,N_12652);
or U13931 (N_13931,N_13595,N_13589);
nor U13932 (N_13932,N_13230,N_13609);
or U13933 (N_13933,N_13528,N_12623);
and U13934 (N_13934,N_13094,N_13691);
nor U13935 (N_13935,N_12663,N_13387);
and U13936 (N_13936,N_13029,N_12555);
or U13937 (N_13937,N_13683,N_12591);
or U13938 (N_13938,N_12599,N_12760);
or U13939 (N_13939,N_13543,N_13638);
or U13940 (N_13940,N_13418,N_13218);
and U13941 (N_13941,N_12656,N_12858);
nor U13942 (N_13942,N_13597,N_13255);
and U13943 (N_13943,N_12861,N_13668);
nor U13944 (N_13944,N_13444,N_12779);
or U13945 (N_13945,N_12536,N_12546);
or U13946 (N_13946,N_13693,N_12967);
nand U13947 (N_13947,N_13096,N_13376);
nor U13948 (N_13948,N_13101,N_12562);
xnor U13949 (N_13949,N_13466,N_13534);
nand U13950 (N_13950,N_13734,N_12627);
xor U13951 (N_13951,N_12860,N_12932);
nand U13952 (N_13952,N_12761,N_13257);
or U13953 (N_13953,N_13477,N_13133);
or U13954 (N_13954,N_13461,N_12557);
nand U13955 (N_13955,N_12919,N_13038);
nand U13956 (N_13956,N_12520,N_12680);
nor U13957 (N_13957,N_13288,N_12569);
nor U13958 (N_13958,N_13677,N_13530);
nor U13959 (N_13959,N_13468,N_13722);
xor U13960 (N_13960,N_13471,N_13709);
nand U13961 (N_13961,N_13120,N_13088);
xor U13962 (N_13962,N_13443,N_12789);
or U13963 (N_13963,N_13717,N_13219);
nor U13964 (N_13964,N_13294,N_13025);
and U13965 (N_13965,N_12902,N_13400);
and U13966 (N_13966,N_13521,N_12999);
or U13967 (N_13967,N_13583,N_12909);
xor U13968 (N_13968,N_12895,N_13082);
nor U13969 (N_13969,N_12791,N_13446);
or U13970 (N_13970,N_13613,N_12676);
nor U13971 (N_13971,N_13130,N_13398);
nor U13972 (N_13972,N_13307,N_12827);
nor U13973 (N_13973,N_13654,N_13576);
or U13974 (N_13974,N_13377,N_12767);
xnor U13975 (N_13975,N_13645,N_13195);
xnor U13976 (N_13976,N_13086,N_13365);
or U13977 (N_13977,N_12905,N_12817);
nor U13978 (N_13978,N_13464,N_12503);
and U13979 (N_13979,N_13362,N_12565);
nand U13980 (N_13980,N_12622,N_12984);
nand U13981 (N_13981,N_13259,N_12662);
or U13982 (N_13982,N_13593,N_12798);
or U13983 (N_13983,N_12974,N_12736);
nand U13984 (N_13984,N_13569,N_13348);
nor U13985 (N_13985,N_12510,N_13502);
and U13986 (N_13986,N_13629,N_12530);
nor U13987 (N_13987,N_13224,N_13529);
or U13988 (N_13988,N_13720,N_12891);
nand U13989 (N_13989,N_13189,N_13034);
or U13990 (N_13990,N_12749,N_13695);
xor U13991 (N_13991,N_13023,N_12813);
nor U13992 (N_13992,N_13620,N_13429);
nand U13993 (N_13993,N_12972,N_12505);
or U13994 (N_13994,N_13055,N_12866);
nand U13995 (N_13995,N_12850,N_13542);
or U13996 (N_13996,N_13384,N_13131);
and U13997 (N_13997,N_13032,N_12691);
or U13998 (N_13998,N_13519,N_13548);
nand U13999 (N_13999,N_12880,N_12745);
or U14000 (N_14000,N_13305,N_13009);
and U14001 (N_14001,N_13630,N_12824);
nor U14002 (N_14002,N_12848,N_13602);
nand U14003 (N_14003,N_13500,N_12976);
nand U14004 (N_14004,N_13646,N_13212);
or U14005 (N_14005,N_12867,N_13741);
xnor U14006 (N_14006,N_12994,N_12872);
xor U14007 (N_14007,N_13177,N_12724);
nor U14008 (N_14008,N_12512,N_12790);
xnor U14009 (N_14009,N_13022,N_13382);
or U14010 (N_14010,N_13107,N_13412);
and U14011 (N_14011,N_12683,N_12797);
nor U14012 (N_14012,N_13577,N_12707);
nand U14013 (N_14013,N_13269,N_13441);
and U14014 (N_14014,N_13458,N_13119);
nor U14015 (N_14015,N_12846,N_13243);
nand U14016 (N_14016,N_13397,N_12721);
xnor U14017 (N_14017,N_12887,N_13690);
or U14018 (N_14018,N_13634,N_13184);
or U14019 (N_14019,N_13590,N_13659);
nand U14020 (N_14020,N_12885,N_12507);
xnor U14021 (N_14021,N_12611,N_13514);
nand U14022 (N_14022,N_12811,N_12842);
or U14023 (N_14023,N_12709,N_13118);
nor U14024 (N_14024,N_13208,N_12593);
nor U14025 (N_14025,N_13448,N_13204);
nand U14026 (N_14026,N_13156,N_13414);
and U14027 (N_14027,N_13707,N_13216);
or U14028 (N_14028,N_13008,N_13050);
and U14029 (N_14029,N_13748,N_12687);
or U14030 (N_14030,N_12552,N_13363);
and U14031 (N_14031,N_12748,N_12668);
xor U14032 (N_14032,N_13011,N_12762);
xor U14033 (N_14033,N_13447,N_13141);
nor U14034 (N_14034,N_12759,N_13241);
xor U14035 (N_14035,N_13735,N_12549);
nand U14036 (N_14036,N_12532,N_12678);
nand U14037 (N_14037,N_13494,N_13077);
nor U14038 (N_14038,N_13474,N_12819);
or U14039 (N_14039,N_12765,N_12522);
nand U14040 (N_14040,N_13612,N_13371);
xor U14041 (N_14041,N_12541,N_13581);
nand U14042 (N_14042,N_13083,N_13368);
and U14043 (N_14043,N_13031,N_13718);
nand U14044 (N_14044,N_13713,N_12782);
and U14045 (N_14045,N_13395,N_13633);
or U14046 (N_14046,N_13578,N_12916);
nand U14047 (N_14047,N_13503,N_12711);
nand U14048 (N_14048,N_13048,N_13134);
nor U14049 (N_14049,N_12845,N_13221);
or U14050 (N_14050,N_12928,N_12589);
xor U14051 (N_14051,N_13481,N_13231);
xor U14052 (N_14052,N_12729,N_13664);
or U14053 (N_14053,N_13084,N_12940);
nand U14054 (N_14054,N_12757,N_13273);
nor U14055 (N_14055,N_13287,N_13267);
nor U14056 (N_14056,N_13739,N_12710);
nor U14057 (N_14057,N_13312,N_12901);
nor U14058 (N_14058,N_13253,N_13105);
nor U14059 (N_14059,N_13642,N_13650);
and U14060 (N_14060,N_13251,N_13355);
or U14061 (N_14061,N_13686,N_13042);
xnor U14062 (N_14062,N_13358,N_13201);
or U14063 (N_14063,N_12701,N_12996);
nand U14064 (N_14064,N_12805,N_13636);
nand U14065 (N_14065,N_13125,N_13168);
and U14066 (N_14066,N_13246,N_12585);
and U14067 (N_14067,N_12877,N_12859);
or U14068 (N_14068,N_12679,N_13694);
and U14069 (N_14069,N_12733,N_13392);
and U14070 (N_14070,N_13052,N_12517);
xnor U14071 (N_14071,N_13399,N_12632);
xor U14072 (N_14072,N_13584,N_12832);
nor U14073 (N_14073,N_13316,N_13747);
or U14074 (N_14074,N_13711,N_12807);
and U14075 (N_14075,N_13605,N_13154);
nand U14076 (N_14076,N_12995,N_12903);
xor U14077 (N_14077,N_13652,N_13128);
and U14078 (N_14078,N_13496,N_12971);
xnor U14079 (N_14079,N_13454,N_12578);
or U14080 (N_14080,N_12990,N_12834);
and U14081 (N_14081,N_13616,N_13506);
nand U14082 (N_14082,N_12592,N_13565);
nor U14083 (N_14083,N_13423,N_12913);
nand U14084 (N_14084,N_13226,N_13340);
nand U14085 (N_14085,N_13553,N_13323);
or U14086 (N_14086,N_12695,N_13432);
and U14087 (N_14087,N_13389,N_13268);
xor U14088 (N_14088,N_12900,N_13374);
and U14089 (N_14089,N_13028,N_12630);
nand U14090 (N_14090,N_13300,N_12518);
or U14091 (N_14091,N_12583,N_13164);
nor U14092 (N_14092,N_13696,N_12666);
nor U14093 (N_14093,N_13056,N_13345);
nand U14094 (N_14094,N_13357,N_12501);
nand U14095 (N_14095,N_12948,N_13112);
nand U14096 (N_14096,N_12644,N_12542);
xor U14097 (N_14097,N_12934,N_13169);
nand U14098 (N_14098,N_13081,N_12615);
or U14099 (N_14099,N_13010,N_12787);
xnor U14100 (N_14100,N_13588,N_13364);
nor U14101 (N_14101,N_12777,N_13598);
nor U14102 (N_14102,N_13284,N_12500);
or U14103 (N_14103,N_13192,N_12544);
nand U14104 (N_14104,N_12796,N_12925);
xnor U14105 (N_14105,N_13676,N_13001);
and U14106 (N_14106,N_12973,N_12723);
nand U14107 (N_14107,N_13698,N_13098);
xnor U14108 (N_14108,N_13322,N_13271);
or U14109 (N_14109,N_13671,N_13003);
nor U14110 (N_14110,N_13062,N_13144);
nor U14111 (N_14111,N_12841,N_12788);
xnor U14112 (N_14112,N_13205,N_13237);
or U14113 (N_14113,N_12734,N_13625);
or U14114 (N_14114,N_13729,N_13026);
xnor U14115 (N_14115,N_12582,N_12689);
and U14116 (N_14116,N_13047,N_13152);
or U14117 (N_14117,N_12669,N_12588);
xor U14118 (N_14118,N_12778,N_12508);
xor U14119 (N_14119,N_12890,N_13505);
xor U14120 (N_14120,N_12764,N_12677);
and U14121 (N_14121,N_12560,N_12810);
nand U14122 (N_14122,N_13064,N_12649);
nand U14123 (N_14123,N_12843,N_12911);
nand U14124 (N_14124,N_12641,N_13336);
and U14125 (N_14125,N_13380,N_13497);
or U14126 (N_14126,N_12978,N_13736);
nand U14127 (N_14127,N_13329,N_12621);
xor U14128 (N_14128,N_12814,N_12624);
nor U14129 (N_14129,N_13297,N_12551);
and U14130 (N_14130,N_13249,N_13352);
xnor U14131 (N_14131,N_13465,N_13113);
nand U14132 (N_14132,N_13238,N_12857);
nor U14133 (N_14133,N_13280,N_12613);
nand U14134 (N_14134,N_12714,N_12580);
nor U14135 (N_14135,N_12667,N_13085);
or U14136 (N_14136,N_12853,N_13182);
nand U14137 (N_14137,N_12653,N_13596);
and U14138 (N_14138,N_13649,N_13452);
xnor U14139 (N_14139,N_12566,N_13520);
or U14140 (N_14140,N_13334,N_13175);
or U14141 (N_14141,N_12598,N_12849);
and U14142 (N_14142,N_13325,N_12577);
or U14143 (N_14143,N_13040,N_13470);
nand U14144 (N_14144,N_12979,N_13245);
nor U14145 (N_14145,N_12879,N_13544);
or U14146 (N_14146,N_13127,N_12639);
nand U14147 (N_14147,N_13442,N_13116);
xor U14148 (N_14148,N_13559,N_13002);
nor U14149 (N_14149,N_13673,N_13158);
xor U14150 (N_14150,N_13574,N_12944);
nand U14151 (N_14151,N_13587,N_12553);
and U14152 (N_14152,N_12970,N_13328);
and U14153 (N_14153,N_12620,N_12855);
nand U14154 (N_14154,N_13335,N_13617);
or U14155 (N_14155,N_12783,N_13498);
and U14156 (N_14156,N_13174,N_13603);
nor U14157 (N_14157,N_13054,N_12573);
xor U14158 (N_14158,N_13223,N_12803);
and U14159 (N_14159,N_12567,N_12524);
or U14160 (N_14160,N_12572,N_13099);
and U14161 (N_14161,N_13663,N_13431);
xor U14162 (N_14162,N_13669,N_13211);
nor U14163 (N_14163,N_13433,N_13367);
xnor U14164 (N_14164,N_13037,N_12625);
and U14165 (N_14165,N_12579,N_12766);
xor U14166 (N_14166,N_12672,N_12595);
and U14167 (N_14167,N_12642,N_12535);
nor U14168 (N_14168,N_12692,N_13068);
and U14169 (N_14169,N_13469,N_13679);
nor U14170 (N_14170,N_13303,N_13067);
nor U14171 (N_14171,N_13608,N_13314);
nand U14172 (N_14172,N_13039,N_13343);
or U14173 (N_14173,N_13666,N_12527);
and U14174 (N_14174,N_13293,N_13599);
nand U14175 (N_14175,N_13331,N_12862);
nand U14176 (N_14176,N_13535,N_12929);
nor U14177 (N_14177,N_13388,N_13570);
xnor U14178 (N_14178,N_12584,N_13393);
nor U14179 (N_14179,N_13532,N_13321);
xor U14180 (N_14180,N_13250,N_12664);
nand U14181 (N_14181,N_12758,N_12673);
or U14182 (N_14182,N_13647,N_13685);
nor U14183 (N_14183,N_12935,N_13440);
nor U14184 (N_14184,N_12889,N_13122);
or U14185 (N_14185,N_13353,N_13427);
or U14186 (N_14186,N_12590,N_12750);
nand U14187 (N_14187,N_13737,N_12795);
nand U14188 (N_14188,N_13410,N_13715);
or U14189 (N_14189,N_13485,N_13610);
xor U14190 (N_14190,N_12600,N_12596);
nor U14191 (N_14191,N_13540,N_13541);
xnor U14192 (N_14192,N_13641,N_13193);
xnor U14193 (N_14193,N_12607,N_13566);
or U14194 (N_14194,N_13058,N_13228);
nand U14195 (N_14195,N_13455,N_12908);
nand U14196 (N_14196,N_13276,N_13370);
and U14197 (N_14197,N_12897,N_13296);
nor U14198 (N_14198,N_13147,N_12826);
and U14199 (N_14199,N_13227,N_13699);
or U14200 (N_14200,N_12784,N_13360);
nor U14201 (N_14201,N_13744,N_12886);
xor U14202 (N_14202,N_12603,N_12809);
nor U14203 (N_14203,N_12617,N_13507);
nand U14204 (N_14204,N_13283,N_12509);
xnor U14205 (N_14205,N_13552,N_13235);
nor U14206 (N_14206,N_13024,N_13333);
xor U14207 (N_14207,N_12945,N_12513);
xor U14208 (N_14208,N_13247,N_12981);
nor U14209 (N_14209,N_12706,N_12956);
nand U14210 (N_14210,N_12547,N_13486);
nand U14211 (N_14211,N_12586,N_12700);
and U14212 (N_14212,N_13344,N_13585);
and U14213 (N_14213,N_13150,N_12619);
or U14214 (N_14214,N_12671,N_13006);
xor U14215 (N_14215,N_12661,N_13108);
xor U14216 (N_14216,N_13173,N_12980);
and U14217 (N_14217,N_13016,N_13572);
or U14218 (N_14218,N_13615,N_13674);
or U14219 (N_14219,N_13229,N_13021);
nand U14220 (N_14220,N_13200,N_12896);
or U14221 (N_14221,N_12571,N_13339);
and U14222 (N_14222,N_13491,N_13202);
nor U14223 (N_14223,N_13386,N_13252);
xnor U14224 (N_14224,N_13157,N_12907);
nand U14225 (N_14225,N_13522,N_12726);
and U14226 (N_14226,N_12781,N_13310);
nor U14227 (N_14227,N_12949,N_12868);
xor U14228 (N_14228,N_12794,N_13369);
or U14229 (N_14229,N_13413,N_12960);
or U14230 (N_14230,N_13733,N_13155);
or U14231 (N_14231,N_12650,N_13342);
nor U14232 (N_14232,N_12574,N_12793);
nand U14233 (N_14233,N_13727,N_13203);
nor U14234 (N_14234,N_12708,N_13430);
or U14235 (N_14235,N_13493,N_13337);
or U14236 (N_14236,N_13197,N_13728);
or U14237 (N_14237,N_13743,N_12992);
or U14238 (N_14238,N_13176,N_12874);
nor U14239 (N_14239,N_13422,N_13373);
or U14240 (N_14240,N_12993,N_13547);
xnor U14241 (N_14241,N_13667,N_13420);
nor U14242 (N_14242,N_13349,N_12534);
or U14243 (N_14243,N_12969,N_12835);
nor U14244 (N_14244,N_12966,N_13439);
and U14245 (N_14245,N_13242,N_13586);
nand U14246 (N_14246,N_12735,N_13209);
and U14247 (N_14247,N_13366,N_13621);
or U14248 (N_14248,N_12704,N_13095);
nor U14249 (N_14249,N_13411,N_13640);
and U14250 (N_14250,N_13111,N_12786);
nand U14251 (N_14251,N_12775,N_13080);
or U14252 (N_14252,N_12634,N_12998);
and U14253 (N_14253,N_13185,N_12852);
and U14254 (N_14254,N_12742,N_13165);
or U14255 (N_14255,N_13061,N_13554);
nor U14256 (N_14256,N_13005,N_13706);
or U14257 (N_14257,N_13524,N_12550);
xnor U14258 (N_14258,N_12806,N_13066);
nor U14259 (N_14259,N_13489,N_13473);
or U14260 (N_14260,N_13631,N_13234);
xor U14261 (N_14261,N_12754,N_13379);
and U14262 (N_14262,N_13017,N_13622);
nor U14263 (N_14263,N_13656,N_13478);
or U14264 (N_14264,N_12955,N_12962);
nor U14265 (N_14265,N_13140,N_13053);
or U14266 (N_14266,N_12828,N_12660);
or U14267 (N_14267,N_13490,N_12674);
or U14268 (N_14268,N_13306,N_12772);
nor U14269 (N_14269,N_13256,N_12636);
nor U14270 (N_14270,N_13714,N_13538);
nand U14271 (N_14271,N_13515,N_13199);
nor U14272 (N_14272,N_12612,N_12833);
or U14273 (N_14273,N_13426,N_13167);
nand U14274 (N_14274,N_13264,N_12987);
nand U14275 (N_14275,N_12977,N_13660);
and U14276 (N_14276,N_13600,N_12892);
xor U14277 (N_14277,N_13402,N_12938);
nor U14278 (N_14278,N_13041,N_13178);
or U14279 (N_14279,N_13324,N_12502);
xnor U14280 (N_14280,N_13115,N_12933);
and U14281 (N_14281,N_13716,N_13428);
xor U14282 (N_14282,N_13643,N_13580);
nand U14283 (N_14283,N_13299,N_13035);
and U14284 (N_14284,N_12802,N_13406);
nor U14285 (N_14285,N_13460,N_12910);
nor U14286 (N_14286,N_12991,N_12904);
or U14287 (N_14287,N_13145,N_13187);
nand U14288 (N_14288,N_12628,N_13172);
xor U14289 (N_14289,N_12921,N_13611);
or U14290 (N_14290,N_12685,N_13512);
nand U14291 (N_14291,N_13724,N_12725);
xor U14292 (N_14292,N_12959,N_13146);
xnor U14293 (N_14293,N_13248,N_12519);
or U14294 (N_14294,N_12941,N_12648);
or U14295 (N_14295,N_13425,N_13097);
xor U14296 (N_14296,N_13550,N_12820);
or U14297 (N_14297,N_13457,N_13375);
nand U14298 (N_14298,N_12694,N_13281);
nor U14299 (N_14299,N_13286,N_13372);
xnor U14300 (N_14300,N_12773,N_12686);
nand U14301 (N_14301,N_13687,N_12605);
xnor U14302 (N_14302,N_12774,N_13240);
or U14303 (N_14303,N_13065,N_12743);
nor U14304 (N_14304,N_12822,N_13302);
nor U14305 (N_14305,N_13206,N_13618);
xor U14306 (N_14306,N_13702,N_13126);
nor U14307 (N_14307,N_12747,N_12640);
and U14308 (N_14308,N_12645,N_12836);
nand U14309 (N_14309,N_12728,N_13019);
nand U14310 (N_14310,N_13689,N_12863);
nor U14311 (N_14311,N_13124,N_13278);
or U14312 (N_14312,N_13419,N_13624);
nor U14313 (N_14313,N_13060,N_13539);
nand U14314 (N_14314,N_12717,N_13100);
and U14315 (N_14315,N_12638,N_12988);
xor U14316 (N_14316,N_12602,N_12703);
or U14317 (N_14317,N_12631,N_13103);
or U14318 (N_14318,N_13138,N_13708);
and U14319 (N_14319,N_13136,N_12780);
xor U14320 (N_14320,N_13272,N_13632);
nand U14321 (N_14321,N_13330,N_12752);
or U14322 (N_14322,N_12568,N_12715);
nand U14323 (N_14323,N_13036,N_13509);
nor U14324 (N_14324,N_12647,N_12884);
nand U14325 (N_14325,N_12529,N_13093);
or U14326 (N_14326,N_13087,N_13057);
xnor U14327 (N_14327,N_12718,N_12610);
nor U14328 (N_14328,N_12526,N_12740);
nand U14329 (N_14329,N_13012,N_12958);
and U14330 (N_14330,N_13076,N_13424);
or U14331 (N_14331,N_13648,N_13591);
xor U14332 (N_14332,N_12914,N_13401);
and U14333 (N_14333,N_13295,N_13456);
nand U14334 (N_14334,N_13712,N_12719);
nor U14335 (N_14335,N_12888,N_12985);
and U14336 (N_14336,N_13628,N_13675);
or U14337 (N_14337,N_13308,N_13463);
xnor U14338 (N_14338,N_12570,N_12906);
nand U14339 (N_14339,N_13526,N_13090);
xnor U14340 (N_14340,N_12515,N_13536);
or U14341 (N_14341,N_13472,N_13484);
and U14342 (N_14342,N_13462,N_13573);
or U14343 (N_14343,N_13198,N_13746);
xor U14344 (N_14344,N_13678,N_13385);
or U14345 (N_14345,N_12626,N_13075);
and U14346 (N_14346,N_12558,N_13560);
nor U14347 (N_14347,N_12739,N_13210);
and U14348 (N_14348,N_12917,N_13109);
xnor U14349 (N_14349,N_13149,N_13265);
xor U14350 (N_14350,N_12698,N_12818);
xor U14351 (N_14351,N_12521,N_12629);
xor U14352 (N_14352,N_13326,N_12722);
or U14353 (N_14353,N_12808,N_13670);
or U14354 (N_14354,N_13700,N_12606);
xor U14355 (N_14355,N_12815,N_13277);
xnor U14356 (N_14356,N_13046,N_12514);
xor U14357 (N_14357,N_12538,N_12712);
xor U14358 (N_14358,N_13351,N_13434);
and U14359 (N_14359,N_13151,N_13114);
nor U14360 (N_14360,N_13239,N_12763);
nand U14361 (N_14361,N_13394,N_13487);
or U14362 (N_14362,N_13730,N_13213);
and U14363 (N_14363,N_12702,N_13327);
and U14364 (N_14364,N_13186,N_13051);
or U14365 (N_14365,N_12899,N_13416);
and U14366 (N_14366,N_13637,N_13262);
or U14367 (N_14367,N_13275,N_12738);
nor U14368 (N_14368,N_13163,N_12840);
nand U14369 (N_14369,N_13129,N_13575);
nand U14370 (N_14370,N_12792,N_13749);
and U14371 (N_14371,N_12511,N_13396);
xor U14372 (N_14372,N_13346,N_13403);
xnor U14373 (N_14373,N_13561,N_12654);
xnor U14374 (N_14374,N_13537,N_13516);
nor U14375 (N_14375,N_12569,N_13035);
or U14376 (N_14376,N_12536,N_13275);
nand U14377 (N_14377,N_13731,N_13653);
xnor U14378 (N_14378,N_13677,N_13207);
or U14379 (N_14379,N_13706,N_13424);
xnor U14380 (N_14380,N_12814,N_12848);
or U14381 (N_14381,N_13638,N_13433);
xor U14382 (N_14382,N_12923,N_13648);
or U14383 (N_14383,N_13689,N_12892);
nor U14384 (N_14384,N_13214,N_13182);
xor U14385 (N_14385,N_13046,N_13023);
xor U14386 (N_14386,N_12841,N_12720);
or U14387 (N_14387,N_12684,N_12925);
or U14388 (N_14388,N_12646,N_13129);
nor U14389 (N_14389,N_13072,N_12824);
or U14390 (N_14390,N_13375,N_13664);
or U14391 (N_14391,N_13214,N_13281);
nand U14392 (N_14392,N_13031,N_13179);
xor U14393 (N_14393,N_12785,N_13443);
or U14394 (N_14394,N_13358,N_12632);
xor U14395 (N_14395,N_13596,N_12521);
xnor U14396 (N_14396,N_13286,N_12633);
and U14397 (N_14397,N_12973,N_13183);
nor U14398 (N_14398,N_12831,N_13189);
xor U14399 (N_14399,N_13132,N_13133);
xnor U14400 (N_14400,N_12500,N_13732);
xor U14401 (N_14401,N_13636,N_13632);
xnor U14402 (N_14402,N_13269,N_12964);
nor U14403 (N_14403,N_12967,N_12667);
nor U14404 (N_14404,N_13299,N_13346);
and U14405 (N_14405,N_12515,N_13715);
and U14406 (N_14406,N_12854,N_13172);
or U14407 (N_14407,N_13421,N_13562);
and U14408 (N_14408,N_13152,N_12917);
and U14409 (N_14409,N_13042,N_13408);
nand U14410 (N_14410,N_12810,N_13170);
xnor U14411 (N_14411,N_13662,N_13648);
xor U14412 (N_14412,N_12656,N_12933);
nor U14413 (N_14413,N_13146,N_13583);
and U14414 (N_14414,N_12623,N_12613);
nand U14415 (N_14415,N_13012,N_13002);
and U14416 (N_14416,N_13134,N_12612);
xor U14417 (N_14417,N_13123,N_12701);
and U14418 (N_14418,N_13726,N_13168);
xnor U14419 (N_14419,N_13715,N_12757);
or U14420 (N_14420,N_13748,N_12670);
or U14421 (N_14421,N_13004,N_13141);
nor U14422 (N_14422,N_13527,N_13247);
and U14423 (N_14423,N_13013,N_13747);
or U14424 (N_14424,N_12884,N_12889);
and U14425 (N_14425,N_13592,N_13497);
xor U14426 (N_14426,N_12939,N_13745);
and U14427 (N_14427,N_12577,N_12894);
nor U14428 (N_14428,N_13551,N_12786);
nor U14429 (N_14429,N_12798,N_12783);
nor U14430 (N_14430,N_13262,N_12898);
or U14431 (N_14431,N_12633,N_13204);
nor U14432 (N_14432,N_12554,N_13591);
xnor U14433 (N_14433,N_12558,N_12919);
nor U14434 (N_14434,N_13238,N_12612);
or U14435 (N_14435,N_13238,N_13067);
nand U14436 (N_14436,N_13172,N_13292);
and U14437 (N_14437,N_13553,N_13359);
and U14438 (N_14438,N_13279,N_13098);
nor U14439 (N_14439,N_13093,N_13017);
xnor U14440 (N_14440,N_13236,N_12649);
xnor U14441 (N_14441,N_13049,N_12932);
nand U14442 (N_14442,N_13689,N_13456);
and U14443 (N_14443,N_12613,N_13635);
nor U14444 (N_14444,N_13284,N_13454);
nor U14445 (N_14445,N_13599,N_13606);
and U14446 (N_14446,N_12964,N_13272);
and U14447 (N_14447,N_13245,N_13542);
xor U14448 (N_14448,N_12604,N_13007);
and U14449 (N_14449,N_13599,N_12555);
and U14450 (N_14450,N_12719,N_13099);
xor U14451 (N_14451,N_13577,N_12995);
nand U14452 (N_14452,N_13671,N_13270);
and U14453 (N_14453,N_13512,N_13187);
nand U14454 (N_14454,N_12678,N_12628);
nand U14455 (N_14455,N_12650,N_13171);
nor U14456 (N_14456,N_13351,N_13265);
nor U14457 (N_14457,N_13070,N_13702);
or U14458 (N_14458,N_13350,N_13141);
nor U14459 (N_14459,N_13695,N_13305);
xor U14460 (N_14460,N_12707,N_12703);
xor U14461 (N_14461,N_12708,N_12563);
xor U14462 (N_14462,N_13126,N_12820);
or U14463 (N_14463,N_13165,N_13220);
xnor U14464 (N_14464,N_13002,N_13250);
xor U14465 (N_14465,N_13208,N_13067);
nor U14466 (N_14466,N_13566,N_13241);
nand U14467 (N_14467,N_13367,N_13514);
or U14468 (N_14468,N_13573,N_13278);
xnor U14469 (N_14469,N_13350,N_13505);
and U14470 (N_14470,N_13461,N_12924);
or U14471 (N_14471,N_13641,N_13725);
or U14472 (N_14472,N_12889,N_13218);
and U14473 (N_14473,N_13582,N_13192);
nand U14474 (N_14474,N_13616,N_13455);
and U14475 (N_14475,N_12988,N_13141);
nor U14476 (N_14476,N_12603,N_13293);
and U14477 (N_14477,N_13618,N_12932);
nor U14478 (N_14478,N_13429,N_13092);
nand U14479 (N_14479,N_13530,N_13432);
xnor U14480 (N_14480,N_12836,N_13156);
nor U14481 (N_14481,N_13254,N_12668);
xor U14482 (N_14482,N_13097,N_13202);
nor U14483 (N_14483,N_12571,N_12921);
and U14484 (N_14484,N_13276,N_13450);
or U14485 (N_14485,N_13206,N_13559);
xor U14486 (N_14486,N_13163,N_13216);
and U14487 (N_14487,N_13629,N_12864);
xor U14488 (N_14488,N_13565,N_13088);
xnor U14489 (N_14489,N_13619,N_13278);
nor U14490 (N_14490,N_13269,N_12841);
nor U14491 (N_14491,N_12555,N_12742);
nand U14492 (N_14492,N_13547,N_13063);
xnor U14493 (N_14493,N_12670,N_13291);
and U14494 (N_14494,N_12749,N_12822);
xor U14495 (N_14495,N_12582,N_13642);
nand U14496 (N_14496,N_13675,N_13651);
nand U14497 (N_14497,N_12665,N_13168);
xor U14498 (N_14498,N_13342,N_13109);
or U14499 (N_14499,N_13402,N_12692);
nor U14500 (N_14500,N_13088,N_12508);
nor U14501 (N_14501,N_12676,N_13697);
or U14502 (N_14502,N_13239,N_12874);
and U14503 (N_14503,N_12889,N_13117);
nand U14504 (N_14504,N_13580,N_13015);
xnor U14505 (N_14505,N_12652,N_12786);
and U14506 (N_14506,N_13703,N_13690);
and U14507 (N_14507,N_13225,N_12683);
and U14508 (N_14508,N_13634,N_13176);
xor U14509 (N_14509,N_13517,N_12652);
nand U14510 (N_14510,N_13123,N_12718);
nand U14511 (N_14511,N_13005,N_13074);
xnor U14512 (N_14512,N_13238,N_12685);
nand U14513 (N_14513,N_12829,N_13729);
and U14514 (N_14514,N_13055,N_12711);
and U14515 (N_14515,N_12909,N_13316);
or U14516 (N_14516,N_13322,N_13304);
and U14517 (N_14517,N_13168,N_13227);
xnor U14518 (N_14518,N_12648,N_12748);
nor U14519 (N_14519,N_13387,N_12671);
or U14520 (N_14520,N_13500,N_13657);
nor U14521 (N_14521,N_12938,N_12898);
nand U14522 (N_14522,N_12586,N_12642);
nor U14523 (N_14523,N_13224,N_12830);
nor U14524 (N_14524,N_12518,N_12633);
nand U14525 (N_14525,N_13413,N_12678);
xor U14526 (N_14526,N_12503,N_13676);
or U14527 (N_14527,N_13545,N_13151);
xnor U14528 (N_14528,N_12524,N_12509);
nor U14529 (N_14529,N_12659,N_13701);
nor U14530 (N_14530,N_13007,N_12690);
and U14531 (N_14531,N_13252,N_12693);
and U14532 (N_14532,N_12567,N_13598);
and U14533 (N_14533,N_13210,N_13326);
or U14534 (N_14534,N_13451,N_12547);
and U14535 (N_14535,N_12527,N_13406);
xnor U14536 (N_14536,N_13033,N_13472);
or U14537 (N_14537,N_12594,N_12932);
nand U14538 (N_14538,N_13402,N_12735);
and U14539 (N_14539,N_13427,N_13365);
nand U14540 (N_14540,N_13606,N_13161);
nand U14541 (N_14541,N_13629,N_13607);
or U14542 (N_14542,N_13349,N_13235);
nor U14543 (N_14543,N_13191,N_12678);
xor U14544 (N_14544,N_12801,N_13687);
nor U14545 (N_14545,N_13354,N_12507);
or U14546 (N_14546,N_12845,N_12734);
nor U14547 (N_14547,N_13446,N_12572);
xnor U14548 (N_14548,N_12546,N_13739);
or U14549 (N_14549,N_12640,N_12657);
or U14550 (N_14550,N_13041,N_12907);
or U14551 (N_14551,N_13377,N_12600);
xnor U14552 (N_14552,N_13324,N_13078);
xnor U14553 (N_14553,N_12861,N_13231);
nor U14554 (N_14554,N_13426,N_12725);
or U14555 (N_14555,N_12695,N_13131);
nand U14556 (N_14556,N_12724,N_13641);
or U14557 (N_14557,N_13346,N_13515);
or U14558 (N_14558,N_12518,N_13080);
nand U14559 (N_14559,N_12575,N_13136);
xor U14560 (N_14560,N_13353,N_12807);
xor U14561 (N_14561,N_13538,N_13635);
nand U14562 (N_14562,N_12646,N_12864);
or U14563 (N_14563,N_12864,N_13591);
and U14564 (N_14564,N_12837,N_12642);
nand U14565 (N_14565,N_13050,N_12653);
nor U14566 (N_14566,N_13029,N_13044);
nand U14567 (N_14567,N_13179,N_12984);
nand U14568 (N_14568,N_13653,N_13123);
and U14569 (N_14569,N_13205,N_12573);
nand U14570 (N_14570,N_13711,N_12854);
and U14571 (N_14571,N_13106,N_12665);
xor U14572 (N_14572,N_13425,N_13070);
nand U14573 (N_14573,N_12640,N_13630);
nand U14574 (N_14574,N_12912,N_12539);
nand U14575 (N_14575,N_13389,N_13718);
or U14576 (N_14576,N_12729,N_12740);
or U14577 (N_14577,N_13062,N_13174);
or U14578 (N_14578,N_13378,N_13656);
xor U14579 (N_14579,N_12510,N_12984);
and U14580 (N_14580,N_12929,N_13572);
nand U14581 (N_14581,N_13464,N_13409);
and U14582 (N_14582,N_13002,N_13310);
nand U14583 (N_14583,N_13480,N_13270);
and U14584 (N_14584,N_13001,N_12942);
and U14585 (N_14585,N_13322,N_13664);
or U14586 (N_14586,N_13728,N_13168);
nand U14587 (N_14587,N_13304,N_13748);
nand U14588 (N_14588,N_13606,N_12879);
and U14589 (N_14589,N_13720,N_12630);
and U14590 (N_14590,N_12861,N_12582);
nand U14591 (N_14591,N_13276,N_13664);
and U14592 (N_14592,N_13735,N_13338);
nor U14593 (N_14593,N_13744,N_12660);
and U14594 (N_14594,N_13224,N_12809);
and U14595 (N_14595,N_12600,N_13227);
and U14596 (N_14596,N_12530,N_12582);
or U14597 (N_14597,N_13545,N_13113);
or U14598 (N_14598,N_13587,N_12749);
and U14599 (N_14599,N_13059,N_13105);
and U14600 (N_14600,N_13568,N_13382);
nor U14601 (N_14601,N_13244,N_13481);
nand U14602 (N_14602,N_13735,N_13666);
xor U14603 (N_14603,N_12655,N_12843);
nor U14604 (N_14604,N_12885,N_13468);
xor U14605 (N_14605,N_13328,N_13401);
nand U14606 (N_14606,N_12781,N_12623);
nand U14607 (N_14607,N_13493,N_13089);
nor U14608 (N_14608,N_12556,N_13173);
nor U14609 (N_14609,N_13134,N_12854);
xnor U14610 (N_14610,N_13107,N_12719);
nand U14611 (N_14611,N_13046,N_12561);
or U14612 (N_14612,N_13627,N_13413);
and U14613 (N_14613,N_12611,N_13282);
and U14614 (N_14614,N_13013,N_13201);
nor U14615 (N_14615,N_13287,N_13491);
and U14616 (N_14616,N_12866,N_13288);
and U14617 (N_14617,N_12644,N_13094);
or U14618 (N_14618,N_13016,N_12936);
xnor U14619 (N_14619,N_13239,N_13483);
and U14620 (N_14620,N_12645,N_12531);
or U14621 (N_14621,N_13456,N_12800);
xor U14622 (N_14622,N_12878,N_13548);
or U14623 (N_14623,N_12838,N_13591);
or U14624 (N_14624,N_12691,N_12683);
nor U14625 (N_14625,N_12774,N_12674);
or U14626 (N_14626,N_12948,N_12867);
nand U14627 (N_14627,N_12825,N_12726);
xor U14628 (N_14628,N_13735,N_12582);
or U14629 (N_14629,N_12795,N_13602);
nor U14630 (N_14630,N_12607,N_12939);
and U14631 (N_14631,N_12710,N_12666);
xnor U14632 (N_14632,N_12891,N_12759);
xor U14633 (N_14633,N_13032,N_12614);
nor U14634 (N_14634,N_13687,N_13649);
or U14635 (N_14635,N_12581,N_12752);
or U14636 (N_14636,N_12977,N_12625);
and U14637 (N_14637,N_13481,N_13745);
and U14638 (N_14638,N_13359,N_12746);
nand U14639 (N_14639,N_12795,N_12818);
or U14640 (N_14640,N_13613,N_13119);
and U14641 (N_14641,N_13234,N_13149);
and U14642 (N_14642,N_13490,N_13114);
nand U14643 (N_14643,N_12537,N_13266);
nand U14644 (N_14644,N_12526,N_13598);
nor U14645 (N_14645,N_12747,N_12563);
nor U14646 (N_14646,N_13052,N_12714);
and U14647 (N_14647,N_13169,N_13237);
or U14648 (N_14648,N_12761,N_13511);
or U14649 (N_14649,N_12984,N_13313);
and U14650 (N_14650,N_12534,N_12512);
nand U14651 (N_14651,N_13380,N_13290);
or U14652 (N_14652,N_13124,N_13181);
or U14653 (N_14653,N_13747,N_13049);
xor U14654 (N_14654,N_13497,N_12787);
nor U14655 (N_14655,N_13553,N_13504);
xor U14656 (N_14656,N_13727,N_12578);
or U14657 (N_14657,N_13411,N_13354);
and U14658 (N_14658,N_13350,N_13675);
and U14659 (N_14659,N_12579,N_13159);
and U14660 (N_14660,N_13203,N_13346);
nand U14661 (N_14661,N_13573,N_12972);
nor U14662 (N_14662,N_13177,N_13537);
xnor U14663 (N_14663,N_13274,N_12639);
nand U14664 (N_14664,N_12905,N_13215);
xor U14665 (N_14665,N_13276,N_12527);
nor U14666 (N_14666,N_13113,N_12857);
and U14667 (N_14667,N_12675,N_13523);
nand U14668 (N_14668,N_13240,N_13167);
nor U14669 (N_14669,N_12652,N_12797);
nand U14670 (N_14670,N_13599,N_13634);
or U14671 (N_14671,N_12776,N_13498);
xnor U14672 (N_14672,N_12577,N_12703);
nand U14673 (N_14673,N_12511,N_13283);
xnor U14674 (N_14674,N_12511,N_13549);
nand U14675 (N_14675,N_12976,N_12802);
or U14676 (N_14676,N_13603,N_13676);
nand U14677 (N_14677,N_13040,N_12516);
nor U14678 (N_14678,N_13519,N_13179);
or U14679 (N_14679,N_13625,N_13261);
xor U14680 (N_14680,N_13352,N_12894);
nor U14681 (N_14681,N_13592,N_12980);
xnor U14682 (N_14682,N_13178,N_12818);
nand U14683 (N_14683,N_12763,N_13012);
nand U14684 (N_14684,N_13466,N_13585);
or U14685 (N_14685,N_13457,N_13158);
xnor U14686 (N_14686,N_13712,N_13423);
nand U14687 (N_14687,N_12975,N_12776);
or U14688 (N_14688,N_12627,N_12513);
and U14689 (N_14689,N_13500,N_12975);
nor U14690 (N_14690,N_13301,N_12909);
xnor U14691 (N_14691,N_12604,N_12939);
nor U14692 (N_14692,N_12845,N_13145);
and U14693 (N_14693,N_13601,N_13737);
and U14694 (N_14694,N_13335,N_13463);
nand U14695 (N_14695,N_12628,N_13299);
nor U14696 (N_14696,N_12774,N_13161);
nand U14697 (N_14697,N_12779,N_13078);
nor U14698 (N_14698,N_13465,N_12581);
nor U14699 (N_14699,N_13676,N_13250);
and U14700 (N_14700,N_13088,N_12916);
nor U14701 (N_14701,N_13534,N_13705);
xnor U14702 (N_14702,N_13374,N_13331);
xnor U14703 (N_14703,N_13025,N_13733);
xor U14704 (N_14704,N_13022,N_13597);
nand U14705 (N_14705,N_13269,N_13287);
xor U14706 (N_14706,N_13428,N_13021);
or U14707 (N_14707,N_12808,N_12574);
and U14708 (N_14708,N_12853,N_13661);
xnor U14709 (N_14709,N_13632,N_12574);
or U14710 (N_14710,N_13361,N_13564);
nor U14711 (N_14711,N_12542,N_13115);
or U14712 (N_14712,N_12980,N_13321);
and U14713 (N_14713,N_13027,N_13590);
nand U14714 (N_14714,N_13087,N_12561);
and U14715 (N_14715,N_12730,N_13714);
and U14716 (N_14716,N_12857,N_13593);
or U14717 (N_14717,N_12524,N_12645);
and U14718 (N_14718,N_12686,N_12522);
or U14719 (N_14719,N_13530,N_13126);
nor U14720 (N_14720,N_12994,N_13303);
xor U14721 (N_14721,N_13446,N_13530);
nand U14722 (N_14722,N_13712,N_12921);
nand U14723 (N_14723,N_12886,N_12992);
or U14724 (N_14724,N_12907,N_13143);
xnor U14725 (N_14725,N_13703,N_13249);
and U14726 (N_14726,N_13664,N_12515);
nor U14727 (N_14727,N_12789,N_13210);
or U14728 (N_14728,N_13118,N_13658);
nand U14729 (N_14729,N_13664,N_13133);
xor U14730 (N_14730,N_12582,N_13719);
and U14731 (N_14731,N_13664,N_13359);
nand U14732 (N_14732,N_13443,N_12620);
nand U14733 (N_14733,N_12847,N_13339);
or U14734 (N_14734,N_12722,N_12958);
nor U14735 (N_14735,N_13677,N_12857);
nand U14736 (N_14736,N_13309,N_13747);
nor U14737 (N_14737,N_12737,N_12527);
or U14738 (N_14738,N_12764,N_12610);
xnor U14739 (N_14739,N_12533,N_12890);
nor U14740 (N_14740,N_12921,N_13231);
or U14741 (N_14741,N_13550,N_12916);
or U14742 (N_14742,N_13457,N_13580);
xor U14743 (N_14743,N_12965,N_12636);
nor U14744 (N_14744,N_13543,N_12855);
nand U14745 (N_14745,N_12956,N_13572);
and U14746 (N_14746,N_12872,N_13383);
nor U14747 (N_14747,N_12920,N_13081);
nand U14748 (N_14748,N_13041,N_13010);
xor U14749 (N_14749,N_13707,N_13548);
and U14750 (N_14750,N_13645,N_13739);
and U14751 (N_14751,N_13595,N_13576);
xor U14752 (N_14752,N_13129,N_12853);
nor U14753 (N_14753,N_13005,N_12643);
or U14754 (N_14754,N_12583,N_13240);
xor U14755 (N_14755,N_13288,N_12671);
nand U14756 (N_14756,N_13644,N_13174);
xor U14757 (N_14757,N_13254,N_13466);
nand U14758 (N_14758,N_12848,N_12653);
nand U14759 (N_14759,N_12601,N_12573);
nor U14760 (N_14760,N_13385,N_12642);
nand U14761 (N_14761,N_13605,N_12567);
nor U14762 (N_14762,N_13693,N_12912);
nand U14763 (N_14763,N_13644,N_12682);
and U14764 (N_14764,N_13569,N_12761);
and U14765 (N_14765,N_13628,N_13064);
xor U14766 (N_14766,N_13713,N_13072);
nand U14767 (N_14767,N_12953,N_13054);
nor U14768 (N_14768,N_13225,N_12762);
and U14769 (N_14769,N_13097,N_13465);
or U14770 (N_14770,N_13181,N_12766);
nand U14771 (N_14771,N_13075,N_13236);
xor U14772 (N_14772,N_13137,N_13197);
or U14773 (N_14773,N_12709,N_13458);
nand U14774 (N_14774,N_13370,N_13414);
xor U14775 (N_14775,N_13342,N_12553);
xnor U14776 (N_14776,N_12572,N_12854);
nor U14777 (N_14777,N_12895,N_12773);
or U14778 (N_14778,N_12927,N_13005);
nand U14779 (N_14779,N_13451,N_13739);
xor U14780 (N_14780,N_13187,N_12915);
xnor U14781 (N_14781,N_13062,N_13695);
or U14782 (N_14782,N_13645,N_13581);
and U14783 (N_14783,N_12989,N_13043);
or U14784 (N_14784,N_12745,N_13020);
nand U14785 (N_14785,N_12854,N_12639);
nor U14786 (N_14786,N_13291,N_13423);
nand U14787 (N_14787,N_12849,N_13275);
and U14788 (N_14788,N_12871,N_12893);
nand U14789 (N_14789,N_13618,N_13739);
and U14790 (N_14790,N_12666,N_13333);
and U14791 (N_14791,N_13488,N_12885);
and U14792 (N_14792,N_13281,N_13671);
nor U14793 (N_14793,N_13442,N_12785);
or U14794 (N_14794,N_12835,N_12616);
nor U14795 (N_14795,N_13289,N_12891);
and U14796 (N_14796,N_12927,N_13707);
xor U14797 (N_14797,N_12557,N_12937);
nand U14798 (N_14798,N_12625,N_13372);
and U14799 (N_14799,N_12810,N_13287);
and U14800 (N_14800,N_13051,N_13321);
nor U14801 (N_14801,N_12710,N_13289);
xor U14802 (N_14802,N_12998,N_12603);
or U14803 (N_14803,N_13340,N_12935);
xnor U14804 (N_14804,N_13229,N_13174);
and U14805 (N_14805,N_13020,N_13357);
or U14806 (N_14806,N_13270,N_12645);
xor U14807 (N_14807,N_13004,N_12829);
nand U14808 (N_14808,N_13527,N_13717);
or U14809 (N_14809,N_12612,N_12729);
nor U14810 (N_14810,N_13484,N_12859);
or U14811 (N_14811,N_13065,N_12710);
xor U14812 (N_14812,N_12973,N_13050);
or U14813 (N_14813,N_12530,N_12794);
nand U14814 (N_14814,N_13394,N_12965);
nand U14815 (N_14815,N_12764,N_12525);
xor U14816 (N_14816,N_13235,N_12643);
xor U14817 (N_14817,N_12805,N_12904);
xor U14818 (N_14818,N_12766,N_12744);
nand U14819 (N_14819,N_13447,N_12958);
xnor U14820 (N_14820,N_13171,N_12622);
and U14821 (N_14821,N_13627,N_13541);
or U14822 (N_14822,N_12806,N_13032);
and U14823 (N_14823,N_12631,N_12860);
or U14824 (N_14824,N_12641,N_13506);
xnor U14825 (N_14825,N_12586,N_13283);
nor U14826 (N_14826,N_13280,N_12611);
and U14827 (N_14827,N_12754,N_12577);
xor U14828 (N_14828,N_12689,N_12589);
nor U14829 (N_14829,N_12994,N_12926);
and U14830 (N_14830,N_13481,N_12690);
nor U14831 (N_14831,N_13599,N_12989);
nand U14832 (N_14832,N_12594,N_12549);
nand U14833 (N_14833,N_12674,N_13284);
nor U14834 (N_14834,N_13215,N_13749);
xor U14835 (N_14835,N_12700,N_12982);
xnor U14836 (N_14836,N_13022,N_12890);
and U14837 (N_14837,N_13661,N_13051);
nor U14838 (N_14838,N_13242,N_12878);
and U14839 (N_14839,N_13367,N_13487);
and U14840 (N_14840,N_13098,N_12584);
xnor U14841 (N_14841,N_13637,N_13058);
xnor U14842 (N_14842,N_13330,N_13155);
nand U14843 (N_14843,N_13490,N_13483);
nor U14844 (N_14844,N_13622,N_12924);
and U14845 (N_14845,N_12885,N_12850);
xnor U14846 (N_14846,N_13095,N_13156);
nand U14847 (N_14847,N_13152,N_13608);
nor U14848 (N_14848,N_13336,N_12723);
xor U14849 (N_14849,N_12920,N_13142);
or U14850 (N_14850,N_12699,N_12867);
or U14851 (N_14851,N_12965,N_13041);
and U14852 (N_14852,N_12606,N_12747);
xor U14853 (N_14853,N_13088,N_12969);
nand U14854 (N_14854,N_13716,N_13044);
xor U14855 (N_14855,N_13663,N_13351);
nand U14856 (N_14856,N_13583,N_12943);
nand U14857 (N_14857,N_12955,N_12633);
and U14858 (N_14858,N_12879,N_13384);
and U14859 (N_14859,N_12525,N_13004);
xor U14860 (N_14860,N_12546,N_12939);
and U14861 (N_14861,N_13133,N_13735);
or U14862 (N_14862,N_12871,N_13318);
xnor U14863 (N_14863,N_13303,N_13086);
or U14864 (N_14864,N_12579,N_13120);
or U14865 (N_14865,N_13548,N_12922);
nor U14866 (N_14866,N_13469,N_12524);
nand U14867 (N_14867,N_13533,N_13088);
nor U14868 (N_14868,N_12895,N_12647);
nor U14869 (N_14869,N_13486,N_12875);
nor U14870 (N_14870,N_12576,N_13090);
xor U14871 (N_14871,N_13438,N_13705);
or U14872 (N_14872,N_12943,N_13667);
or U14873 (N_14873,N_13135,N_12773);
xnor U14874 (N_14874,N_13574,N_13650);
nor U14875 (N_14875,N_12800,N_13635);
or U14876 (N_14876,N_13223,N_13528);
nor U14877 (N_14877,N_13200,N_13227);
or U14878 (N_14878,N_13632,N_13239);
xor U14879 (N_14879,N_13572,N_13369);
and U14880 (N_14880,N_12984,N_13390);
nand U14881 (N_14881,N_13642,N_12935);
xnor U14882 (N_14882,N_12623,N_13579);
xor U14883 (N_14883,N_13568,N_13209);
and U14884 (N_14884,N_13454,N_13401);
or U14885 (N_14885,N_13486,N_13627);
and U14886 (N_14886,N_12655,N_13253);
xor U14887 (N_14887,N_12845,N_12720);
nor U14888 (N_14888,N_13743,N_13725);
nand U14889 (N_14889,N_13639,N_13285);
xor U14890 (N_14890,N_13045,N_13099);
nand U14891 (N_14891,N_12988,N_13058);
nor U14892 (N_14892,N_12944,N_12629);
xnor U14893 (N_14893,N_13639,N_13413);
nor U14894 (N_14894,N_12678,N_13315);
or U14895 (N_14895,N_12750,N_13593);
or U14896 (N_14896,N_13671,N_13249);
xnor U14897 (N_14897,N_13139,N_12997);
nand U14898 (N_14898,N_13576,N_13196);
nor U14899 (N_14899,N_12716,N_13719);
nand U14900 (N_14900,N_12709,N_13734);
xor U14901 (N_14901,N_13564,N_13203);
xnor U14902 (N_14902,N_13692,N_13107);
nand U14903 (N_14903,N_12688,N_13502);
and U14904 (N_14904,N_13737,N_12962);
or U14905 (N_14905,N_13370,N_13472);
nand U14906 (N_14906,N_12568,N_12954);
and U14907 (N_14907,N_13232,N_13026);
nand U14908 (N_14908,N_13444,N_12830);
nor U14909 (N_14909,N_12557,N_13334);
nor U14910 (N_14910,N_12908,N_13511);
or U14911 (N_14911,N_12699,N_13356);
or U14912 (N_14912,N_12621,N_12783);
and U14913 (N_14913,N_13507,N_13396);
and U14914 (N_14914,N_12980,N_12733);
or U14915 (N_14915,N_12796,N_13253);
nor U14916 (N_14916,N_12808,N_12536);
or U14917 (N_14917,N_13382,N_12573);
or U14918 (N_14918,N_12915,N_12655);
or U14919 (N_14919,N_12513,N_12788);
and U14920 (N_14920,N_13411,N_12950);
nand U14921 (N_14921,N_12987,N_13727);
nor U14922 (N_14922,N_12988,N_13504);
nand U14923 (N_14923,N_12844,N_12860);
nor U14924 (N_14924,N_13355,N_12784);
or U14925 (N_14925,N_13498,N_13328);
xor U14926 (N_14926,N_13607,N_13088);
xnor U14927 (N_14927,N_12747,N_12961);
nand U14928 (N_14928,N_13295,N_13591);
nand U14929 (N_14929,N_13235,N_12595);
or U14930 (N_14930,N_12652,N_12712);
nor U14931 (N_14931,N_13736,N_12508);
and U14932 (N_14932,N_12534,N_13025);
or U14933 (N_14933,N_12527,N_13315);
nand U14934 (N_14934,N_13033,N_13022);
and U14935 (N_14935,N_13706,N_13102);
xnor U14936 (N_14936,N_13497,N_12728);
nand U14937 (N_14937,N_12564,N_13511);
and U14938 (N_14938,N_12771,N_12896);
nand U14939 (N_14939,N_13716,N_12942);
nor U14940 (N_14940,N_12943,N_13575);
nor U14941 (N_14941,N_13420,N_13074);
xor U14942 (N_14942,N_12641,N_13307);
and U14943 (N_14943,N_13040,N_13735);
nand U14944 (N_14944,N_12629,N_13184);
nand U14945 (N_14945,N_12714,N_13430);
or U14946 (N_14946,N_12651,N_12747);
xor U14947 (N_14947,N_13185,N_13614);
nor U14948 (N_14948,N_12920,N_12851);
nand U14949 (N_14949,N_13710,N_13560);
nor U14950 (N_14950,N_13198,N_13559);
xnor U14951 (N_14951,N_12603,N_13419);
nand U14952 (N_14952,N_13678,N_13606);
nand U14953 (N_14953,N_13282,N_12985);
nand U14954 (N_14954,N_12942,N_13739);
xor U14955 (N_14955,N_12529,N_12850);
nor U14956 (N_14956,N_13168,N_13121);
nand U14957 (N_14957,N_13544,N_12575);
or U14958 (N_14958,N_13504,N_12875);
nand U14959 (N_14959,N_13530,N_13280);
xnor U14960 (N_14960,N_13144,N_13553);
nand U14961 (N_14961,N_13510,N_12609);
and U14962 (N_14962,N_13047,N_13061);
nand U14963 (N_14963,N_13161,N_13413);
nor U14964 (N_14964,N_13292,N_13282);
or U14965 (N_14965,N_13138,N_12591);
xnor U14966 (N_14966,N_13535,N_13045);
or U14967 (N_14967,N_12655,N_13377);
nand U14968 (N_14968,N_12652,N_13645);
nand U14969 (N_14969,N_12942,N_12650);
nor U14970 (N_14970,N_12611,N_12663);
nor U14971 (N_14971,N_13126,N_12903);
xor U14972 (N_14972,N_12598,N_13572);
nand U14973 (N_14973,N_13732,N_13195);
and U14974 (N_14974,N_13564,N_12604);
and U14975 (N_14975,N_13685,N_13346);
and U14976 (N_14976,N_12818,N_13355);
nand U14977 (N_14977,N_13470,N_13255);
nand U14978 (N_14978,N_13524,N_12515);
and U14979 (N_14979,N_12925,N_13546);
nor U14980 (N_14980,N_12904,N_13114);
nor U14981 (N_14981,N_12775,N_13520);
and U14982 (N_14982,N_13536,N_13718);
nor U14983 (N_14983,N_12503,N_12804);
nor U14984 (N_14984,N_12914,N_13167);
xor U14985 (N_14985,N_12695,N_13039);
nor U14986 (N_14986,N_12655,N_12997);
xnor U14987 (N_14987,N_12860,N_13636);
or U14988 (N_14988,N_13044,N_12981);
nor U14989 (N_14989,N_13144,N_13157);
nor U14990 (N_14990,N_13668,N_12689);
xnor U14991 (N_14991,N_13716,N_12515);
xnor U14992 (N_14992,N_13715,N_12907);
and U14993 (N_14993,N_13145,N_12758);
nor U14994 (N_14994,N_12680,N_13115);
nand U14995 (N_14995,N_13047,N_12831);
nand U14996 (N_14996,N_13525,N_12992);
nand U14997 (N_14997,N_12974,N_13546);
and U14998 (N_14998,N_13528,N_13340);
nor U14999 (N_14999,N_12725,N_12976);
xor U15000 (N_15000,N_13804,N_14276);
or U15001 (N_15001,N_14574,N_14132);
and U15002 (N_15002,N_13767,N_14859);
nand U15003 (N_15003,N_14399,N_14945);
or U15004 (N_15004,N_14179,N_14134);
or U15005 (N_15005,N_14192,N_14886);
and U15006 (N_15006,N_13797,N_14553);
or U15007 (N_15007,N_14170,N_14277);
nor U15008 (N_15008,N_14707,N_14249);
xor U15009 (N_15009,N_14567,N_14382);
nand U15010 (N_15010,N_14002,N_14877);
nand U15011 (N_15011,N_13918,N_14594);
nand U15012 (N_15012,N_13807,N_14472);
xor U15013 (N_15013,N_14576,N_14280);
and U15014 (N_15014,N_13853,N_14298);
xor U15015 (N_15015,N_14048,N_14517);
nor U15016 (N_15016,N_14366,N_14747);
nand U15017 (N_15017,N_14824,N_14414);
and U15018 (N_15018,N_14214,N_14614);
nor U15019 (N_15019,N_14496,N_14869);
xor U15020 (N_15020,N_14921,N_14938);
nand U15021 (N_15021,N_14865,N_14846);
and U15022 (N_15022,N_14081,N_14626);
nor U15023 (N_15023,N_14584,N_14686);
or U15024 (N_15024,N_14705,N_13985);
xnor U15025 (N_15025,N_14473,N_14805);
or U15026 (N_15026,N_14789,N_14979);
nand U15027 (N_15027,N_14844,N_14702);
or U15028 (N_15028,N_14813,N_14448);
and U15029 (N_15029,N_14142,N_14578);
or U15030 (N_15030,N_14294,N_14841);
or U15031 (N_15031,N_13915,N_13983);
and U15032 (N_15032,N_14332,N_14203);
and U15033 (N_15033,N_14773,N_14286);
or U15034 (N_15034,N_14531,N_14794);
xor U15035 (N_15035,N_14776,N_14477);
or U15036 (N_15036,N_14720,N_14289);
nand U15037 (N_15037,N_14333,N_14852);
nor U15038 (N_15038,N_14459,N_14281);
or U15039 (N_15039,N_14334,N_13887);
or U15040 (N_15040,N_14356,N_14968);
or U15041 (N_15041,N_14949,N_14906);
nor U15042 (N_15042,N_14548,N_14954);
nand U15043 (N_15043,N_13798,N_14245);
and U15044 (N_15044,N_14084,N_14480);
nand U15045 (N_15045,N_14244,N_14648);
xnor U15046 (N_15046,N_14812,N_14840);
nor U15047 (N_15047,N_13870,N_14788);
nor U15048 (N_15048,N_14185,N_14427);
nand U15049 (N_15049,N_14308,N_13862);
and U15050 (N_15050,N_14215,N_14947);
xor U15051 (N_15051,N_14030,N_14229);
and U15052 (N_15052,N_14232,N_14903);
xnor U15053 (N_15053,N_14407,N_14975);
and U15054 (N_15054,N_14020,N_14741);
xor U15055 (N_15055,N_14549,N_13879);
or U15056 (N_15056,N_14823,N_14733);
or U15057 (N_15057,N_14853,N_13991);
xnor U15058 (N_15058,N_14934,N_14128);
or U15059 (N_15059,N_14994,N_14821);
nor U15060 (N_15060,N_14072,N_13987);
xnor U15061 (N_15061,N_14113,N_14038);
nand U15062 (N_15062,N_13855,N_14816);
nand U15063 (N_15063,N_14898,N_14624);
nand U15064 (N_15064,N_14362,N_14351);
xor U15065 (N_15065,N_13792,N_13871);
xor U15066 (N_15066,N_14312,N_14438);
or U15067 (N_15067,N_14115,N_14653);
xor U15068 (N_15068,N_13825,N_14564);
xor U15069 (N_15069,N_14116,N_13913);
nand U15070 (N_15070,N_14739,N_14725);
nand U15071 (N_15071,N_14470,N_14166);
nand U15072 (N_15072,N_14011,N_14354);
nand U15073 (N_15073,N_14835,N_14446);
nand U15074 (N_15074,N_14176,N_14951);
and U15075 (N_15075,N_14090,N_14087);
xnor U15076 (N_15076,N_14264,N_14041);
or U15077 (N_15077,N_14242,N_14655);
xor U15078 (N_15078,N_14696,N_14323);
nand U15079 (N_15079,N_14629,N_14717);
xor U15080 (N_15080,N_13924,N_14457);
or U15081 (N_15081,N_14905,N_13828);
nor U15082 (N_15082,N_13838,N_14631);
xnor U15083 (N_15083,N_14093,N_13884);
or U15084 (N_15084,N_14487,N_14984);
nor U15085 (N_15085,N_13858,N_14443);
and U15086 (N_15086,N_14123,N_13824);
xnor U15087 (N_15087,N_13908,N_14524);
nor U15088 (N_15088,N_14490,N_14909);
xor U15089 (N_15089,N_14914,N_14940);
or U15090 (N_15090,N_14783,N_14522);
or U15091 (N_15091,N_14714,N_14328);
nor U15092 (N_15092,N_14617,N_14027);
or U15093 (N_15093,N_14770,N_14317);
xnor U15094 (N_15094,N_14408,N_14801);
nand U15095 (N_15095,N_14143,N_14378);
or U15096 (N_15096,N_14642,N_14661);
nor U15097 (N_15097,N_14300,N_14601);
nor U15098 (N_15098,N_14296,N_13809);
xor U15099 (N_15099,N_14061,N_14969);
or U15100 (N_15100,N_13770,N_14726);
xnor U15101 (N_15101,N_14431,N_14077);
or U15102 (N_15102,N_14603,N_14119);
or U15103 (N_15103,N_14887,N_13823);
xor U15104 (N_15104,N_13889,N_14533);
and U15105 (N_15105,N_14899,N_14868);
nor U15106 (N_15106,N_14201,N_14510);
nand U15107 (N_15107,N_13947,N_14257);
nand U15108 (N_15108,N_14191,N_14110);
xnor U15109 (N_15109,N_14095,N_14656);
and U15110 (N_15110,N_14013,N_14799);
nor U15111 (N_15111,N_14337,N_13953);
or U15112 (N_15112,N_14863,N_14521);
nand U15113 (N_15113,N_14715,N_14340);
and U15114 (N_15114,N_14809,N_14238);
xor U15115 (N_15115,N_14645,N_14543);
nand U15116 (N_15116,N_14220,N_14461);
nand U15117 (N_15117,N_13826,N_14034);
or U15118 (N_15118,N_13859,N_13920);
nor U15119 (N_15119,N_14297,N_14929);
nor U15120 (N_15120,N_14953,N_13793);
or U15121 (N_15121,N_14358,N_14508);
or U15122 (N_15122,N_14664,N_14767);
and U15123 (N_15123,N_14625,N_14729);
nor U15124 (N_15124,N_14073,N_14600);
nor U15125 (N_15125,N_13805,N_14772);
nor U15126 (N_15126,N_14153,N_14983);
or U15127 (N_15127,N_14186,N_14850);
xor U15128 (N_15128,N_14096,N_14247);
xor U15129 (N_15129,N_14708,N_14442);
or U15130 (N_15130,N_14152,N_14724);
and U15131 (N_15131,N_14550,N_13764);
and U15132 (N_15132,N_14336,N_13754);
nand U15133 (N_15133,N_14019,N_14195);
or U15134 (N_15134,N_14076,N_14120);
nor U15135 (N_15135,N_14795,N_14671);
and U15136 (N_15136,N_13976,N_14313);
or U15137 (N_15137,N_14124,N_13989);
nor U15138 (N_15138,N_14912,N_14223);
or U15139 (N_15139,N_14409,N_14764);
and U15140 (N_15140,N_14043,N_14558);
nand U15141 (N_15141,N_14107,N_14917);
xor U15142 (N_15142,N_13979,N_13949);
or U15143 (N_15143,N_14608,N_14923);
xor U15144 (N_15144,N_14540,N_14069);
and U15145 (N_15145,N_14270,N_14634);
or U15146 (N_15146,N_14737,N_14891);
xor U15147 (N_15147,N_14430,N_14727);
or U15148 (N_15148,N_14613,N_13932);
and U15149 (N_15149,N_13863,N_13821);
and U15150 (N_15150,N_14632,N_13790);
and U15151 (N_15151,N_13750,N_14721);
or U15152 (N_15152,N_14620,N_14818);
nand U15153 (N_15153,N_13752,N_14098);
nand U15154 (N_15154,N_14800,N_14454);
nor U15155 (N_15155,N_14883,N_14165);
nand U15156 (N_15156,N_14941,N_14897);
or U15157 (N_15157,N_14082,N_14663);
nor U15158 (N_15158,N_14782,N_14911);
nand U15159 (N_15159,N_14598,N_13917);
xnor U15160 (N_15160,N_14527,N_14676);
nand U15161 (N_15161,N_14820,N_14506);
xnor U15162 (N_15162,N_14562,N_14746);
nor U15163 (N_15163,N_13951,N_14713);
or U15164 (N_15164,N_14042,N_14856);
xor U15165 (N_15165,N_13929,N_14144);
and U15166 (N_15166,N_14927,N_14207);
or U15167 (N_15167,N_14920,N_13990);
nor U15168 (N_15168,N_14039,N_13995);
nand U15169 (N_15169,N_14516,N_14761);
or U15170 (N_15170,N_14150,N_14682);
xor U15171 (N_15171,N_14698,N_14651);
nor U15172 (N_15172,N_14749,N_14109);
and U15173 (N_15173,N_14557,N_14924);
nand U15174 (N_15174,N_14592,N_14140);
or U15175 (N_15175,N_14224,N_14748);
or U15176 (N_15176,N_14063,N_14248);
nand U15177 (N_15177,N_14704,N_13851);
nor U15178 (N_15178,N_14751,N_14138);
xnor U15179 (N_15179,N_14610,N_13844);
nor U15180 (N_15180,N_13931,N_14993);
and U15181 (N_15181,N_14503,N_14709);
xnor U15182 (N_15182,N_14094,N_14167);
xnor U15183 (N_15183,N_14383,N_14274);
xor U15184 (N_15184,N_14568,N_14998);
nand U15185 (N_15185,N_14847,N_14037);
or U15186 (N_15186,N_14985,N_14484);
nor U15187 (N_15187,N_14440,N_14211);
nand U15188 (N_15188,N_14602,N_14010);
nor U15189 (N_15189,N_14106,N_14070);
and U15190 (N_15190,N_14593,N_13776);
nand U15191 (N_15191,N_14606,N_14875);
or U15192 (N_15192,N_14139,N_14449);
nand U15193 (N_15193,N_14363,N_14114);
nor U15194 (N_15194,N_14990,N_13897);
and U15195 (N_15195,N_13799,N_13774);
xor U15196 (N_15196,N_14768,N_13854);
and U15197 (N_15197,N_14206,N_14599);
nor U15198 (N_15198,N_14973,N_14701);
nand U15199 (N_15199,N_14980,N_14502);
nor U15200 (N_15200,N_14666,N_14250);
xor U15201 (N_15201,N_14423,N_14827);
xnor U15202 (N_15202,N_14633,N_14193);
xor U15203 (N_15203,N_14759,N_14828);
or U15204 (N_15204,N_14960,N_14986);
and U15205 (N_15205,N_13775,N_14851);
xnor U15206 (N_15206,N_14403,N_14916);
nand U15207 (N_15207,N_14971,N_14319);
nor U15208 (N_15208,N_14901,N_14755);
nand U15209 (N_15209,N_14209,N_14667);
xor U15210 (N_15210,N_14722,N_14894);
xor U15211 (N_15211,N_14341,N_14504);
nor U15212 (N_15212,N_14965,N_14650);
nand U15213 (N_15213,N_14062,N_13998);
xnor U15214 (N_15214,N_14157,N_14494);
and U15215 (N_15215,N_14529,N_14586);
or U15216 (N_15216,N_14588,N_13941);
or U15217 (N_15217,N_14475,N_13848);
nand U15218 (N_15218,N_14672,N_13843);
nor U15219 (N_15219,N_14266,N_14829);
nor U15220 (N_15220,N_14311,N_14133);
nand U15221 (N_15221,N_14252,N_13846);
nand U15222 (N_15222,N_14329,N_13937);
nor U15223 (N_15223,N_14199,N_14267);
nor U15224 (N_15224,N_13883,N_14398);
and U15225 (N_15225,N_14743,N_14194);
xor U15226 (N_15226,N_14051,N_14479);
nand U15227 (N_15227,N_14417,N_14159);
or U15228 (N_15228,N_14180,N_14777);
nor U15229 (N_15229,N_13972,N_14752);
nand U15230 (N_15230,N_14053,N_14371);
and U15231 (N_15231,N_14639,N_14991);
or U15232 (N_15232,N_14925,N_14200);
nor U15233 (N_15233,N_13768,N_14445);
nor U15234 (N_15234,N_14866,N_14488);
xor U15235 (N_15235,N_14754,N_13811);
nand U15236 (N_15236,N_14943,N_13999);
xnor U15237 (N_15237,N_14305,N_14129);
or U15238 (N_15238,N_14318,N_14992);
nor U15239 (N_15239,N_14067,N_13751);
nor U15240 (N_15240,N_14511,N_14429);
or U15241 (N_15241,N_13778,N_14885);
and U15242 (N_15242,N_14630,N_14055);
nand U15243 (N_15243,N_14158,N_13784);
or U15244 (N_15244,N_14627,N_13833);
xnor U15245 (N_15245,N_14178,N_14774);
xnor U15246 (N_15246,N_14697,N_13868);
or U15247 (N_15247,N_14616,N_14118);
and U15248 (N_15248,N_14239,N_14187);
and U15249 (N_15249,N_14691,N_14033);
xor U15250 (N_15250,N_14003,N_13815);
and U15251 (N_15251,N_14240,N_14740);
or U15252 (N_15252,N_14915,N_14719);
and U15253 (N_15253,N_14939,N_13818);
xor U15254 (N_15254,N_14552,N_14551);
nor U15255 (N_15255,N_13902,N_14190);
xor U15256 (N_15256,N_14685,N_14532);
nand U15257 (N_15257,N_13922,N_14926);
nor U15258 (N_15258,N_13956,N_14836);
or U15259 (N_15259,N_14862,N_14175);
nand U15260 (N_15260,N_14227,N_14830);
or U15261 (N_15261,N_13861,N_14338);
nor U15262 (N_15262,N_14324,N_13831);
or U15263 (N_15263,N_14291,N_14744);
and U15264 (N_15264,N_13885,N_14460);
or U15265 (N_15265,N_14391,N_13935);
nor U15266 (N_15266,N_14416,N_13869);
or U15267 (N_15267,N_14365,N_14972);
nand U15268 (N_15268,N_14386,N_14309);
nand U15269 (N_15269,N_14346,N_14254);
xnor U15270 (N_15270,N_13975,N_13779);
or U15271 (N_15271,N_14556,N_14775);
xnor U15272 (N_15272,N_13923,N_14879);
and U15273 (N_15273,N_13945,N_14561);
nand U15274 (N_15274,N_14703,N_14355);
xnor U15275 (N_15275,N_14299,N_14463);
nor U15276 (N_15276,N_14060,N_14834);
and U15277 (N_15277,N_13970,N_14679);
nand U15278 (N_15278,N_13919,N_14732);
and U15279 (N_15279,N_13903,N_14628);
nand U15280 (N_15280,N_14888,N_14900);
and U15281 (N_15281,N_14058,N_13934);
xnor U15282 (N_15282,N_14258,N_14837);
and U15283 (N_15283,N_14218,N_14904);
and U15284 (N_15284,N_14253,N_14565);
and U15285 (N_15285,N_14233,N_13977);
nand U15286 (N_15286,N_14230,N_14001);
and U15287 (N_15287,N_14327,N_13755);
nand U15288 (N_15288,N_14471,N_14579);
xor U15289 (N_15289,N_14146,N_14216);
nand U15290 (N_15290,N_14873,N_13968);
or U15291 (N_15291,N_14083,N_14962);
nand U15292 (N_15292,N_13780,N_14155);
and U15293 (N_15293,N_14147,N_13771);
and U15294 (N_15294,N_14347,N_14262);
or U15295 (N_15295,N_14434,N_14519);
or U15296 (N_15296,N_14874,N_14950);
nand U15297 (N_15297,N_14512,N_14538);
xor U15298 (N_15298,N_14590,N_14314);
nand U15299 (N_15299,N_13842,N_14674);
nand U15300 (N_15300,N_14316,N_13969);
nand U15301 (N_15301,N_14287,N_14681);
xnor U15302 (N_15302,N_14374,N_14320);
nor U15303 (N_15303,N_14982,N_14996);
nand U15304 (N_15304,N_14235,N_13974);
nand U15305 (N_15305,N_13994,N_14117);
nor U15306 (N_15306,N_14474,N_14079);
xnor U15307 (N_15307,N_14815,N_14591);
or U15308 (N_15308,N_14217,N_14112);
xnor U15309 (N_15309,N_14988,N_14014);
or U15310 (N_15310,N_13830,N_14738);
or U15311 (N_15311,N_14647,N_14177);
and U15312 (N_15312,N_14970,N_14910);
and U15313 (N_15313,N_14541,N_14793);
and U15314 (N_15314,N_13819,N_13791);
xnor U15315 (N_15315,N_14222,N_14458);
nand U15316 (N_15316,N_14831,N_14451);
and U15317 (N_15317,N_14455,N_14271);
nor U15318 (N_15318,N_13874,N_14078);
or U15319 (N_15319,N_14573,N_14210);
xor U15320 (N_15320,N_13850,N_13827);
and U15321 (N_15321,N_14306,N_14342);
or U15322 (N_15322,N_14394,N_14164);
nor U15323 (N_15323,N_14000,N_14161);
xor U15324 (N_15324,N_14699,N_14101);
nor U15325 (N_15325,N_14961,N_14622);
nor U15326 (N_15326,N_14044,N_14638);
nand U15327 (N_15327,N_14498,N_14208);
nand U15328 (N_15328,N_14880,N_14845);
nand U15329 (N_15329,N_14884,N_14678);
nand U15330 (N_15330,N_14481,N_14221);
nor U15331 (N_15331,N_14958,N_14860);
xor U15332 (N_15332,N_14495,N_13982);
nand U15333 (N_15333,N_14745,N_13898);
nand U15334 (N_15334,N_13986,N_14535);
nand U15335 (N_15335,N_14189,N_14413);
or U15336 (N_15336,N_14263,N_13783);
nor U15337 (N_15337,N_13939,N_14295);
and U15338 (N_15338,N_14765,N_13813);
nor U15339 (N_15339,N_14560,N_14169);
and U15340 (N_15340,N_14184,N_13758);
xnor U15341 (N_15341,N_14520,N_14855);
nor U15342 (N_15342,N_14537,N_14005);
and U15343 (N_15343,N_14811,N_14711);
xnor U15344 (N_15344,N_14290,N_14097);
xnor U15345 (N_15345,N_14467,N_14435);
or U15346 (N_15346,N_14424,N_14325);
xnor U15347 (N_15347,N_14546,N_14056);
or U15348 (N_15348,N_14544,N_14085);
nand U15349 (N_15349,N_14539,N_14361);
and U15350 (N_15350,N_14604,N_14932);
and U15351 (N_15351,N_14605,N_14367);
nor U15352 (N_15352,N_14902,N_14256);
xor U15353 (N_15353,N_14870,N_13930);
and U15354 (N_15354,N_14397,N_13925);
and U15355 (N_15355,N_13927,N_14976);
xor U15356 (N_15356,N_14370,N_14483);
or U15357 (N_15357,N_14452,N_14350);
and U15358 (N_15358,N_14690,N_14896);
nor U15359 (N_15359,N_14231,N_14188);
nand U15360 (N_15360,N_13808,N_14406);
nor U15361 (N_15361,N_13928,N_14563);
nor U15362 (N_15362,N_14395,N_14833);
nor U15363 (N_15363,N_14804,N_14068);
or U15364 (N_15364,N_14771,N_14769);
or U15365 (N_15365,N_14282,N_14518);
nor U15366 (N_15366,N_14074,N_14890);
or U15367 (N_15367,N_14279,N_13960);
and U15368 (N_15368,N_14021,N_14680);
xnor U15369 (N_15369,N_14581,N_13954);
or U15370 (N_15370,N_14065,N_14352);
and U15371 (N_15371,N_14421,N_14571);
nand U15372 (N_15372,N_13880,N_14525);
xnor U15373 (N_15373,N_14753,N_14023);
nand U15374 (N_15374,N_14612,N_13849);
nand U15375 (N_15375,N_14802,N_14967);
xor U15376 (N_15376,N_14436,N_14963);
xor U15377 (N_15377,N_14344,N_14689);
nand U15378 (N_15378,N_14331,N_13964);
xnor U15379 (N_15379,N_14575,N_14787);
or U15380 (N_15380,N_14384,N_14842);
nand U15381 (N_15381,N_14712,N_14955);
nand U15382 (N_15382,N_14644,N_14587);
xnor U15383 (N_15383,N_14349,N_14237);
or U15384 (N_15384,N_14577,N_13943);
nor U15385 (N_15385,N_14047,N_14780);
and U15386 (N_15386,N_14930,N_14657);
or U15387 (N_15387,N_14497,N_14779);
nor U15388 (N_15388,N_13832,N_14760);
nand U15389 (N_15389,N_14677,N_14659);
nand U15390 (N_15390,N_13906,N_14125);
xnor U15391 (N_15391,N_14103,N_14654);
nor U15392 (N_15392,N_14570,N_14688);
or U15393 (N_15393,N_14456,N_13800);
or U15394 (N_15394,N_14031,N_14007);
nand U15395 (N_15395,N_14173,N_13980);
nor U15396 (N_15396,N_13801,N_13763);
and U15397 (N_15397,N_14377,N_13864);
and U15398 (N_15398,N_14046,N_14465);
xnor U15399 (N_15399,N_14500,N_14127);
and U15400 (N_15400,N_14838,N_14045);
xnor U15401 (N_15401,N_14609,N_13944);
xor U15402 (N_15402,N_14236,N_14507);
nor U15403 (N_15403,N_13782,N_14260);
and U15404 (N_15404,N_14392,N_14372);
xor U15405 (N_15405,N_13786,N_14411);
nor U15406 (N_15406,N_14611,N_13904);
xor U15407 (N_15407,N_14432,N_14872);
or U15408 (N_15408,N_14088,N_14861);
xnor U15409 (N_15409,N_13777,N_13914);
or U15410 (N_15410,N_14381,N_13837);
and U15411 (N_15411,N_13963,N_13860);
nor U15412 (N_15412,N_14693,N_14931);
nor U15413 (N_15413,N_14808,N_13973);
xor U15414 (N_15414,N_14018,N_13895);
nand U15415 (N_15415,N_14401,N_14205);
or U15416 (N_15416,N_13952,N_14105);
xnor U15417 (N_15417,N_13788,N_14566);
xnor U15418 (N_15418,N_14024,N_14700);
or U15419 (N_15419,N_13959,N_14649);
nand U15420 (N_15420,N_14389,N_14100);
xor U15421 (N_15421,N_14995,N_14637);
nor U15422 (N_15422,N_14987,N_13841);
nor U15423 (N_15423,N_13961,N_14437);
xnor U15424 (N_15424,N_14212,N_14036);
and U15425 (N_15425,N_13891,N_13796);
nand U15426 (N_15426,N_14049,N_14302);
nand U15427 (N_15427,N_14615,N_13873);
or U15428 (N_15428,N_13822,N_13948);
and U15429 (N_15429,N_13877,N_14148);
nand U15430 (N_15430,N_14476,N_13955);
or U15431 (N_15431,N_13896,N_13942);
or U15432 (N_15432,N_14269,N_14806);
and U15433 (N_15433,N_14756,N_13946);
nand U15434 (N_15434,N_14989,N_13856);
and U15435 (N_15435,N_14154,N_14854);
xor U15436 (N_15436,N_14066,N_14526);
xnor U15437 (N_15437,N_14670,N_14304);
xor U15438 (N_15438,N_14272,N_14464);
nor U15439 (N_15439,N_14373,N_14402);
or U15440 (N_15440,N_13894,N_13761);
or U15441 (N_15441,N_14784,N_14405);
or U15442 (N_15442,N_14814,N_14687);
and U15443 (N_15443,N_14420,N_14636);
nand U15444 (N_15444,N_14798,N_14335);
and U15445 (N_15445,N_14360,N_14035);
xnor U15446 (N_15446,N_14695,N_13769);
nand U15447 (N_15447,N_13881,N_14321);
and U15448 (N_15448,N_13866,N_13760);
or U15449 (N_15449,N_13907,N_14822);
xor U15450 (N_15450,N_13795,N_14439);
nor U15451 (N_15451,N_14052,N_14284);
or U15452 (N_15452,N_13814,N_13966);
and U15453 (N_15453,N_13981,N_13996);
nor U15454 (N_15454,N_14493,N_14559);
or U15455 (N_15455,N_14999,N_13835);
and U15456 (N_15456,N_14307,N_14919);
nand U15457 (N_15457,N_14742,N_14182);
or U15458 (N_15458,N_14646,N_14137);
nand U15459 (N_15459,N_14956,N_14889);
or U15460 (N_15460,N_14623,N_14933);
or U15461 (N_15461,N_13890,N_14937);
or U15462 (N_15462,N_13802,N_14265);
nor U15463 (N_15463,N_14668,N_14278);
xnor U15464 (N_15464,N_14966,N_14162);
nand U15465 (N_15465,N_14936,N_14015);
or U15466 (N_15466,N_14959,N_14283);
and U15467 (N_15467,N_14736,N_14136);
nor U15468 (N_15468,N_13756,N_14466);
or U15469 (N_15469,N_14683,N_14364);
xnor U15470 (N_15470,N_14099,N_14425);
nand U15471 (N_15471,N_14268,N_14913);
nand U15472 (N_15472,N_14583,N_14660);
nand U15473 (N_15473,N_13816,N_14343);
and U15474 (N_15474,N_14022,N_13984);
nor U15475 (N_15475,N_14542,N_14259);
nor U15476 (N_15476,N_14326,N_14054);
nand U15477 (N_15477,N_14426,N_14219);
nand U15478 (N_15478,N_14895,N_14807);
nand U15479 (N_15479,N_14135,N_14198);
and U15480 (N_15480,N_14641,N_14981);
xor U15481 (N_15481,N_13967,N_14528);
or U15482 (N_15482,N_14785,N_14908);
xor U15483 (N_15483,N_14016,N_14163);
and U15484 (N_15484,N_14893,N_14428);
nor U15485 (N_15485,N_14368,N_13971);
and U15486 (N_15486,N_14716,N_14330);
or U15487 (N_15487,N_14580,N_13812);
and U15488 (N_15488,N_14582,N_14597);
xnor U15489 (N_15489,N_13794,N_14607);
nand U15490 (N_15490,N_14515,N_14353);
nor U15491 (N_15491,N_14523,N_14075);
nor U15492 (N_15492,N_14817,N_14126);
nor U15493 (N_15493,N_14204,N_14554);
and U15494 (N_15494,N_14345,N_14735);
or U15495 (N_15495,N_14684,N_14181);
nor U15496 (N_15496,N_13803,N_14501);
xor U15497 (N_15497,N_14675,N_14730);
and U15498 (N_15498,N_13787,N_14149);
or U15499 (N_15499,N_14357,N_14555);
and U15500 (N_15500,N_13845,N_14412);
nand U15501 (N_15501,N_13900,N_13892);
nor U15502 (N_15502,N_14652,N_14944);
nand U15503 (N_15503,N_14462,N_14791);
nand U15504 (N_15504,N_13950,N_14183);
or U15505 (N_15505,N_14922,N_13997);
xor U15506 (N_15506,N_14393,N_13865);
nand U15507 (N_15507,N_14102,N_13785);
or U15508 (N_15508,N_14225,N_13852);
xor U15509 (N_15509,N_14757,N_14665);
xor U15510 (N_15510,N_13766,N_13888);
or U15511 (N_15511,N_13936,N_13836);
or U15512 (N_15512,N_14781,N_14882);
nor U15513 (N_15513,N_14585,N_14410);
nand U15514 (N_15514,N_14728,N_13829);
or U15515 (N_15515,N_14064,N_14168);
xor U15516 (N_15516,N_14226,N_14151);
and U15517 (N_15517,N_13957,N_14275);
nor U15518 (N_15518,N_14876,N_14071);
nor U15519 (N_15519,N_14339,N_14878);
and U15520 (N_15520,N_14589,N_13781);
and U15521 (N_15521,N_14032,N_14243);
nor U15522 (N_15522,N_14017,N_14723);
and U15523 (N_15523,N_14796,N_13905);
or U15524 (N_15524,N_14505,N_14978);
nand U15525 (N_15525,N_13762,N_13857);
xor U15526 (N_15526,N_14658,N_14499);
xor U15527 (N_15527,N_14864,N_14288);
xnor U15528 (N_15528,N_14758,N_14694);
and U15529 (N_15529,N_14643,N_13933);
nand U15530 (N_15530,N_14080,N_14881);
or U15531 (N_15531,N_14619,N_14692);
nand U15532 (N_15532,N_14731,N_14662);
nand U15533 (N_15533,N_14482,N_14572);
and U15534 (N_15534,N_14977,N_14935);
and U15535 (N_15535,N_13810,N_13773);
nand U15536 (N_15536,N_13899,N_14418);
or U15537 (N_15537,N_14145,N_14108);
nor U15538 (N_15538,N_14385,N_14948);
xnor U15539 (N_15539,N_13912,N_14131);
nand U15540 (N_15540,N_14618,N_14025);
or U15541 (N_15541,N_14545,N_14121);
nand U15542 (N_15542,N_14197,N_13938);
or U15543 (N_15543,N_14478,N_14858);
xnor U15544 (N_15544,N_14763,N_13988);
nand U15545 (N_15545,N_14379,N_14012);
nand U15546 (N_15546,N_14778,N_14040);
xnor U15547 (N_15547,N_14415,N_14396);
nor U15548 (N_15548,N_14050,N_14848);
xor U15549 (N_15549,N_14322,N_14028);
nor U15550 (N_15550,N_14441,N_14008);
or U15551 (N_15551,N_13840,N_14857);
and U15552 (N_15552,N_14928,N_14485);
xnor U15553 (N_15553,N_14292,N_13882);
and U15554 (N_15554,N_14673,N_14825);
and U15555 (N_15555,N_14130,N_14710);
nand U15556 (N_15556,N_14530,N_14285);
or U15557 (N_15557,N_13867,N_14228);
nand U15558 (N_15558,N_14255,N_14009);
xnor U15559 (N_15559,N_13753,N_14453);
nand U15560 (N_15560,N_14004,N_14400);
and U15561 (N_15561,N_14839,N_14536);
or U15562 (N_15562,N_13876,N_14315);
or U15563 (N_15563,N_14974,N_14826);
and U15564 (N_15564,N_14918,N_14790);
and U15565 (N_15565,N_13958,N_14762);
nand U15566 (N_15566,N_13911,N_14964);
nand U15567 (N_15567,N_14867,N_14734);
and U15568 (N_15568,N_14892,N_14375);
nand U15569 (N_15569,N_14513,N_14390);
or U15570 (N_15570,N_14202,N_14444);
or U15571 (N_15571,N_14086,N_14026);
or U15572 (N_15572,N_14669,N_14750);
or U15573 (N_15573,N_13978,N_14489);
and U15574 (N_15574,N_14261,N_13993);
nand U15575 (N_15575,N_14387,N_14380);
xnor U15576 (N_15576,N_14348,N_14635);
nand U15577 (N_15577,N_14509,N_14156);
and U15578 (N_15578,N_14786,N_14213);
nor U15579 (N_15579,N_14832,N_14621);
nand U15580 (N_15580,N_13789,N_14310);
nor U15581 (N_15581,N_14369,N_14942);
nand U15582 (N_15582,N_14871,N_14172);
nor U15583 (N_15583,N_14640,N_14006);
nand U15584 (N_15584,N_14486,N_13965);
nor U15585 (N_15585,N_14596,N_14419);
and U15586 (N_15586,N_13901,N_14388);
or U15587 (N_15587,N_14957,N_13757);
xnor U15588 (N_15588,N_14196,N_14122);
or U15589 (N_15589,N_14447,N_13962);
or U15590 (N_15590,N_13940,N_14234);
and U15591 (N_15591,N_13893,N_14468);
or U15592 (N_15592,N_14171,N_14797);
and U15593 (N_15593,N_14246,N_14706);
or U15594 (N_15594,N_14595,N_14273);
nor U15595 (N_15595,N_14141,N_14491);
xor U15596 (N_15596,N_14293,N_13817);
or U15597 (N_15597,N_14160,N_14174);
nor U15598 (N_15598,N_14469,N_14492);
xnor U15599 (N_15599,N_14514,N_14907);
nor U15600 (N_15600,N_14997,N_14718);
or U15601 (N_15601,N_13765,N_14547);
or U15602 (N_15602,N_14422,N_13909);
nand U15603 (N_15603,N_14092,N_14810);
and U15604 (N_15604,N_14359,N_13926);
nor U15605 (N_15605,N_14111,N_14952);
nor U15606 (N_15606,N_14303,N_14241);
nor U15607 (N_15607,N_14057,N_14569);
xnor U15608 (N_15608,N_13992,N_13910);
xor U15609 (N_15609,N_14433,N_14450);
nor U15610 (N_15610,N_14792,N_14849);
or U15611 (N_15611,N_14946,N_14766);
or U15612 (N_15612,N_14534,N_13916);
nor U15613 (N_15613,N_13847,N_13886);
or U15614 (N_15614,N_14251,N_14089);
nor U15615 (N_15615,N_13759,N_14843);
nor U15616 (N_15616,N_14091,N_14819);
nor U15617 (N_15617,N_14059,N_13872);
or U15618 (N_15618,N_14404,N_14376);
nor U15619 (N_15619,N_13772,N_13839);
or U15620 (N_15620,N_14803,N_14029);
nand U15621 (N_15621,N_13878,N_13875);
or U15622 (N_15622,N_13806,N_13921);
and U15623 (N_15623,N_13820,N_14301);
nand U15624 (N_15624,N_14104,N_13834);
and U15625 (N_15625,N_14936,N_14741);
nor U15626 (N_15626,N_14995,N_14307);
xor U15627 (N_15627,N_14427,N_14288);
nand U15628 (N_15628,N_14431,N_14670);
xnor U15629 (N_15629,N_14915,N_13932);
nand U15630 (N_15630,N_14441,N_14596);
xnor U15631 (N_15631,N_14684,N_14426);
xnor U15632 (N_15632,N_14784,N_14950);
nand U15633 (N_15633,N_13877,N_13869);
nor U15634 (N_15634,N_14526,N_14162);
and U15635 (N_15635,N_14029,N_14427);
nand U15636 (N_15636,N_14667,N_14840);
nor U15637 (N_15637,N_14295,N_14040);
xnor U15638 (N_15638,N_14662,N_14744);
nand U15639 (N_15639,N_14863,N_14684);
nor U15640 (N_15640,N_14562,N_14971);
or U15641 (N_15641,N_14319,N_13876);
and U15642 (N_15642,N_14227,N_14897);
nor U15643 (N_15643,N_14810,N_14596);
nor U15644 (N_15644,N_14770,N_13983);
or U15645 (N_15645,N_14826,N_14430);
and U15646 (N_15646,N_14126,N_13893);
and U15647 (N_15647,N_14229,N_14590);
xor U15648 (N_15648,N_14918,N_13865);
nor U15649 (N_15649,N_14547,N_14529);
or U15650 (N_15650,N_14376,N_14768);
nand U15651 (N_15651,N_14626,N_14638);
xnor U15652 (N_15652,N_13990,N_14954);
xnor U15653 (N_15653,N_13966,N_14087);
xor U15654 (N_15654,N_14573,N_14122);
or U15655 (N_15655,N_14014,N_14724);
nor U15656 (N_15656,N_13751,N_14787);
xor U15657 (N_15657,N_14854,N_13857);
nor U15658 (N_15658,N_13755,N_14409);
or U15659 (N_15659,N_13953,N_14729);
nor U15660 (N_15660,N_13908,N_14658);
or U15661 (N_15661,N_14603,N_14490);
and U15662 (N_15662,N_14012,N_14433);
and U15663 (N_15663,N_14354,N_13893);
nor U15664 (N_15664,N_14524,N_14766);
or U15665 (N_15665,N_14622,N_14272);
xnor U15666 (N_15666,N_14924,N_14244);
nand U15667 (N_15667,N_14151,N_14166);
or U15668 (N_15668,N_14241,N_14769);
xor U15669 (N_15669,N_13983,N_14906);
and U15670 (N_15670,N_13820,N_14954);
nand U15671 (N_15671,N_14548,N_13947);
or U15672 (N_15672,N_14426,N_14000);
xnor U15673 (N_15673,N_14977,N_14296);
xor U15674 (N_15674,N_14540,N_14182);
nand U15675 (N_15675,N_13922,N_14297);
and U15676 (N_15676,N_14538,N_13940);
and U15677 (N_15677,N_14281,N_13786);
and U15678 (N_15678,N_13948,N_14739);
xnor U15679 (N_15679,N_14044,N_14951);
nor U15680 (N_15680,N_13840,N_14333);
or U15681 (N_15681,N_13755,N_14603);
nand U15682 (N_15682,N_14264,N_14470);
nor U15683 (N_15683,N_14700,N_14802);
and U15684 (N_15684,N_14179,N_14534);
xnor U15685 (N_15685,N_14322,N_14209);
or U15686 (N_15686,N_14677,N_14812);
or U15687 (N_15687,N_14967,N_14502);
nand U15688 (N_15688,N_14432,N_14017);
nor U15689 (N_15689,N_13918,N_14013);
nor U15690 (N_15690,N_13814,N_13750);
or U15691 (N_15691,N_14697,N_14048);
nand U15692 (N_15692,N_13947,N_14615);
or U15693 (N_15693,N_14149,N_14932);
nor U15694 (N_15694,N_14236,N_13847);
or U15695 (N_15695,N_14968,N_14913);
and U15696 (N_15696,N_14563,N_14072);
nand U15697 (N_15697,N_13908,N_14834);
or U15698 (N_15698,N_14865,N_14590);
nor U15699 (N_15699,N_14303,N_13984);
or U15700 (N_15700,N_14809,N_14588);
and U15701 (N_15701,N_14341,N_14545);
and U15702 (N_15702,N_14795,N_14116);
xor U15703 (N_15703,N_14360,N_13809);
nand U15704 (N_15704,N_14891,N_14241);
and U15705 (N_15705,N_14277,N_13788);
nand U15706 (N_15706,N_14659,N_14109);
or U15707 (N_15707,N_14106,N_14188);
xor U15708 (N_15708,N_14385,N_13952);
nand U15709 (N_15709,N_13971,N_13833);
and U15710 (N_15710,N_14838,N_13926);
and U15711 (N_15711,N_13996,N_13991);
xnor U15712 (N_15712,N_14607,N_13952);
xnor U15713 (N_15713,N_14563,N_14077);
nand U15714 (N_15714,N_14985,N_13886);
and U15715 (N_15715,N_14502,N_14588);
or U15716 (N_15716,N_14359,N_14488);
and U15717 (N_15717,N_13867,N_14500);
nor U15718 (N_15718,N_14166,N_13903);
xor U15719 (N_15719,N_13799,N_13795);
or U15720 (N_15720,N_14537,N_14607);
nand U15721 (N_15721,N_14117,N_14743);
nor U15722 (N_15722,N_14053,N_14211);
nand U15723 (N_15723,N_14233,N_14789);
or U15724 (N_15724,N_14541,N_14005);
and U15725 (N_15725,N_14154,N_14709);
nor U15726 (N_15726,N_14152,N_14144);
xnor U15727 (N_15727,N_14400,N_14532);
and U15728 (N_15728,N_13874,N_13879);
or U15729 (N_15729,N_14120,N_14923);
nand U15730 (N_15730,N_14980,N_14216);
xnor U15731 (N_15731,N_14458,N_14817);
or U15732 (N_15732,N_14407,N_14713);
nand U15733 (N_15733,N_14772,N_13800);
and U15734 (N_15734,N_14666,N_14654);
nor U15735 (N_15735,N_14927,N_14910);
nand U15736 (N_15736,N_14627,N_14708);
nand U15737 (N_15737,N_13936,N_14146);
nand U15738 (N_15738,N_14072,N_14674);
xor U15739 (N_15739,N_13925,N_14793);
and U15740 (N_15740,N_14435,N_14449);
nand U15741 (N_15741,N_14852,N_14646);
nand U15742 (N_15742,N_14892,N_14331);
nor U15743 (N_15743,N_13870,N_14970);
nand U15744 (N_15744,N_13936,N_14467);
nand U15745 (N_15745,N_13927,N_14373);
or U15746 (N_15746,N_14788,N_14173);
nand U15747 (N_15747,N_14864,N_14711);
xor U15748 (N_15748,N_14093,N_14799);
or U15749 (N_15749,N_14601,N_14852);
nand U15750 (N_15750,N_14488,N_14594);
and U15751 (N_15751,N_14557,N_13831);
nand U15752 (N_15752,N_14193,N_14925);
nand U15753 (N_15753,N_14310,N_14332);
nand U15754 (N_15754,N_14995,N_13928);
nand U15755 (N_15755,N_13761,N_14551);
xor U15756 (N_15756,N_13875,N_14241);
or U15757 (N_15757,N_14754,N_14540);
xnor U15758 (N_15758,N_14382,N_14283);
nand U15759 (N_15759,N_14284,N_14119);
xnor U15760 (N_15760,N_14650,N_13996);
xor U15761 (N_15761,N_14181,N_14937);
xor U15762 (N_15762,N_14363,N_14324);
xor U15763 (N_15763,N_13911,N_14344);
or U15764 (N_15764,N_14817,N_13859);
and U15765 (N_15765,N_14655,N_13924);
and U15766 (N_15766,N_14002,N_14623);
and U15767 (N_15767,N_14974,N_14953);
and U15768 (N_15768,N_14116,N_14004);
or U15769 (N_15769,N_13766,N_14221);
xnor U15770 (N_15770,N_14123,N_14698);
nand U15771 (N_15771,N_13850,N_13824);
and U15772 (N_15772,N_14661,N_13977);
or U15773 (N_15773,N_14466,N_14187);
and U15774 (N_15774,N_14897,N_14157);
nand U15775 (N_15775,N_13798,N_14898);
nor U15776 (N_15776,N_14652,N_14323);
and U15777 (N_15777,N_14518,N_14079);
nor U15778 (N_15778,N_14485,N_13862);
or U15779 (N_15779,N_14011,N_14426);
xnor U15780 (N_15780,N_14904,N_14337);
xnor U15781 (N_15781,N_14407,N_13910);
nor U15782 (N_15782,N_14027,N_14940);
or U15783 (N_15783,N_14587,N_14627);
and U15784 (N_15784,N_14483,N_14722);
nor U15785 (N_15785,N_13947,N_14041);
nor U15786 (N_15786,N_14406,N_14012);
and U15787 (N_15787,N_14767,N_13995);
or U15788 (N_15788,N_14208,N_14016);
and U15789 (N_15789,N_14970,N_13943);
or U15790 (N_15790,N_14211,N_14371);
nor U15791 (N_15791,N_14812,N_13813);
xor U15792 (N_15792,N_14583,N_13904);
and U15793 (N_15793,N_14298,N_13936);
and U15794 (N_15794,N_14472,N_13922);
and U15795 (N_15795,N_14194,N_13815);
nand U15796 (N_15796,N_14094,N_13935);
nor U15797 (N_15797,N_14060,N_14660);
and U15798 (N_15798,N_14393,N_14828);
nor U15799 (N_15799,N_14506,N_14275);
nand U15800 (N_15800,N_14029,N_14102);
and U15801 (N_15801,N_13860,N_14329);
nand U15802 (N_15802,N_14533,N_13752);
xnor U15803 (N_15803,N_13829,N_14252);
xor U15804 (N_15804,N_14892,N_14201);
nand U15805 (N_15805,N_14366,N_14735);
xnor U15806 (N_15806,N_14458,N_14510);
nor U15807 (N_15807,N_14275,N_14898);
nand U15808 (N_15808,N_14416,N_14307);
xor U15809 (N_15809,N_14598,N_14554);
xor U15810 (N_15810,N_13840,N_14441);
nor U15811 (N_15811,N_14701,N_14343);
and U15812 (N_15812,N_14056,N_14747);
nor U15813 (N_15813,N_14279,N_14052);
nor U15814 (N_15814,N_14763,N_14654);
xnor U15815 (N_15815,N_14974,N_14184);
nand U15816 (N_15816,N_14655,N_13997);
xor U15817 (N_15817,N_14274,N_13974);
xnor U15818 (N_15818,N_13791,N_14859);
or U15819 (N_15819,N_14367,N_14429);
xor U15820 (N_15820,N_13995,N_14273);
xor U15821 (N_15821,N_14716,N_14491);
and U15822 (N_15822,N_14156,N_14148);
and U15823 (N_15823,N_14306,N_14480);
nand U15824 (N_15824,N_14773,N_14027);
and U15825 (N_15825,N_14108,N_13793);
and U15826 (N_15826,N_14425,N_14496);
nor U15827 (N_15827,N_14741,N_14979);
or U15828 (N_15828,N_14890,N_14947);
nand U15829 (N_15829,N_14761,N_14916);
and U15830 (N_15830,N_14582,N_14444);
xnor U15831 (N_15831,N_14089,N_13866);
nand U15832 (N_15832,N_13984,N_13895);
xnor U15833 (N_15833,N_14943,N_14782);
xor U15834 (N_15834,N_14223,N_14068);
nand U15835 (N_15835,N_14978,N_14919);
xor U15836 (N_15836,N_14446,N_14638);
and U15837 (N_15837,N_14165,N_14010);
or U15838 (N_15838,N_14093,N_14087);
nor U15839 (N_15839,N_13786,N_14534);
nor U15840 (N_15840,N_14492,N_14746);
or U15841 (N_15841,N_13833,N_14737);
nor U15842 (N_15842,N_14269,N_14458);
xnor U15843 (N_15843,N_14881,N_14648);
nor U15844 (N_15844,N_14552,N_14470);
and U15845 (N_15845,N_14695,N_13902);
and U15846 (N_15846,N_14693,N_14365);
xnor U15847 (N_15847,N_14537,N_14083);
and U15848 (N_15848,N_14636,N_13796);
nand U15849 (N_15849,N_14484,N_14047);
and U15850 (N_15850,N_13869,N_14093);
xor U15851 (N_15851,N_13765,N_14208);
nor U15852 (N_15852,N_13950,N_14386);
xnor U15853 (N_15853,N_14756,N_14351);
or U15854 (N_15854,N_14313,N_14165);
nor U15855 (N_15855,N_13923,N_14513);
and U15856 (N_15856,N_13961,N_14058);
nand U15857 (N_15857,N_13942,N_13954);
or U15858 (N_15858,N_14447,N_14537);
xor U15859 (N_15859,N_13950,N_14940);
xnor U15860 (N_15860,N_14540,N_14231);
nor U15861 (N_15861,N_14748,N_14010);
xnor U15862 (N_15862,N_14119,N_14962);
nand U15863 (N_15863,N_13804,N_14521);
xor U15864 (N_15864,N_14079,N_14629);
and U15865 (N_15865,N_14674,N_14661);
and U15866 (N_15866,N_14660,N_13949);
nand U15867 (N_15867,N_14843,N_14907);
nand U15868 (N_15868,N_14892,N_14797);
or U15869 (N_15869,N_14155,N_13948);
xor U15870 (N_15870,N_14793,N_14196);
and U15871 (N_15871,N_14680,N_14845);
nand U15872 (N_15872,N_14392,N_14018);
nand U15873 (N_15873,N_14283,N_14466);
nand U15874 (N_15874,N_14265,N_14210);
xor U15875 (N_15875,N_13954,N_13939);
and U15876 (N_15876,N_14219,N_14120);
nor U15877 (N_15877,N_13943,N_14183);
xor U15878 (N_15878,N_14208,N_14089);
xnor U15879 (N_15879,N_14156,N_13938);
nor U15880 (N_15880,N_14500,N_14426);
or U15881 (N_15881,N_14806,N_14999);
xor U15882 (N_15882,N_14957,N_13878);
and U15883 (N_15883,N_14845,N_13875);
xnor U15884 (N_15884,N_13973,N_14279);
xor U15885 (N_15885,N_14878,N_14737);
nor U15886 (N_15886,N_14635,N_14191);
or U15887 (N_15887,N_14606,N_14514);
nand U15888 (N_15888,N_14347,N_14990);
or U15889 (N_15889,N_14447,N_14929);
xnor U15890 (N_15890,N_14712,N_14487);
nand U15891 (N_15891,N_14571,N_14925);
nor U15892 (N_15892,N_14580,N_13996);
nor U15893 (N_15893,N_13951,N_14558);
xnor U15894 (N_15894,N_14809,N_14574);
xnor U15895 (N_15895,N_14287,N_14897);
nand U15896 (N_15896,N_14979,N_13768);
nand U15897 (N_15897,N_13853,N_14195);
or U15898 (N_15898,N_13952,N_14997);
nand U15899 (N_15899,N_13815,N_14282);
xor U15900 (N_15900,N_14848,N_14371);
xor U15901 (N_15901,N_14878,N_14320);
nor U15902 (N_15902,N_14330,N_13794);
and U15903 (N_15903,N_14634,N_14190);
nand U15904 (N_15904,N_14270,N_14098);
nor U15905 (N_15905,N_13967,N_14505);
and U15906 (N_15906,N_14269,N_14895);
nor U15907 (N_15907,N_14129,N_14784);
and U15908 (N_15908,N_13934,N_14603);
nand U15909 (N_15909,N_14519,N_14437);
xnor U15910 (N_15910,N_14394,N_14780);
and U15911 (N_15911,N_14774,N_14396);
and U15912 (N_15912,N_14332,N_14491);
xor U15913 (N_15913,N_14795,N_14613);
or U15914 (N_15914,N_14187,N_13782);
nor U15915 (N_15915,N_14938,N_14129);
nand U15916 (N_15916,N_14280,N_14607);
and U15917 (N_15917,N_14798,N_14533);
nand U15918 (N_15918,N_14871,N_14296);
nand U15919 (N_15919,N_14458,N_14842);
nand U15920 (N_15920,N_14547,N_14896);
nor U15921 (N_15921,N_14534,N_13750);
nor U15922 (N_15922,N_13955,N_14930);
and U15923 (N_15923,N_14049,N_14853);
nand U15924 (N_15924,N_14475,N_14108);
and U15925 (N_15925,N_13963,N_14281);
nand U15926 (N_15926,N_14713,N_14486);
or U15927 (N_15927,N_14450,N_14201);
nand U15928 (N_15928,N_14879,N_14484);
nor U15929 (N_15929,N_14461,N_13792);
or U15930 (N_15930,N_14964,N_14437);
or U15931 (N_15931,N_14730,N_14487);
or U15932 (N_15932,N_14662,N_14502);
xor U15933 (N_15933,N_14453,N_14575);
nor U15934 (N_15934,N_14026,N_14481);
and U15935 (N_15935,N_14313,N_14470);
or U15936 (N_15936,N_14828,N_13886);
and U15937 (N_15937,N_14341,N_14017);
or U15938 (N_15938,N_14418,N_14751);
nand U15939 (N_15939,N_14427,N_14334);
or U15940 (N_15940,N_14075,N_14057);
and U15941 (N_15941,N_14799,N_14583);
nor U15942 (N_15942,N_14465,N_14533);
xor U15943 (N_15943,N_14303,N_14704);
nor U15944 (N_15944,N_14223,N_13985);
or U15945 (N_15945,N_14839,N_14978);
xor U15946 (N_15946,N_14444,N_14973);
nor U15947 (N_15947,N_14657,N_14512);
and U15948 (N_15948,N_14182,N_13941);
nor U15949 (N_15949,N_14014,N_13934);
nand U15950 (N_15950,N_13790,N_13889);
nand U15951 (N_15951,N_14530,N_14304);
and U15952 (N_15952,N_14488,N_14556);
nand U15953 (N_15953,N_14511,N_13961);
xor U15954 (N_15954,N_14219,N_14492);
nand U15955 (N_15955,N_14078,N_14355);
xnor U15956 (N_15956,N_13838,N_14594);
nand U15957 (N_15957,N_14258,N_14340);
xnor U15958 (N_15958,N_14297,N_14188);
and U15959 (N_15959,N_14280,N_13900);
nand U15960 (N_15960,N_14934,N_14390);
xnor U15961 (N_15961,N_14635,N_14875);
and U15962 (N_15962,N_14350,N_14630);
and U15963 (N_15963,N_14173,N_14879);
nor U15964 (N_15964,N_14747,N_14912);
nor U15965 (N_15965,N_13776,N_13863);
and U15966 (N_15966,N_14673,N_14283);
xnor U15967 (N_15967,N_14340,N_14947);
or U15968 (N_15968,N_14499,N_14677);
and U15969 (N_15969,N_14555,N_14939);
nand U15970 (N_15970,N_13751,N_14972);
and U15971 (N_15971,N_13841,N_14735);
and U15972 (N_15972,N_14182,N_13823);
xnor U15973 (N_15973,N_14999,N_14299);
and U15974 (N_15974,N_13998,N_14894);
xnor U15975 (N_15975,N_13861,N_14056);
and U15976 (N_15976,N_14967,N_13840);
and U15977 (N_15977,N_14317,N_14641);
xnor U15978 (N_15978,N_14737,N_14243);
nor U15979 (N_15979,N_13823,N_14439);
nor U15980 (N_15980,N_14914,N_14279);
and U15981 (N_15981,N_14741,N_14527);
nand U15982 (N_15982,N_13838,N_14542);
or U15983 (N_15983,N_14095,N_14963);
nand U15984 (N_15984,N_14879,N_14509);
nor U15985 (N_15985,N_14613,N_14783);
nor U15986 (N_15986,N_14826,N_14029);
nand U15987 (N_15987,N_14751,N_14943);
nand U15988 (N_15988,N_14776,N_14914);
and U15989 (N_15989,N_14983,N_14372);
nor U15990 (N_15990,N_14457,N_14557);
nor U15991 (N_15991,N_14985,N_14941);
and U15992 (N_15992,N_13905,N_14529);
xnor U15993 (N_15993,N_14238,N_14956);
xor U15994 (N_15994,N_14343,N_13870);
xnor U15995 (N_15995,N_14880,N_14138);
and U15996 (N_15996,N_13807,N_14027);
nand U15997 (N_15997,N_13952,N_14829);
and U15998 (N_15998,N_14059,N_13761);
and U15999 (N_15999,N_14653,N_14267);
or U16000 (N_16000,N_13794,N_13846);
xnor U16001 (N_16001,N_14228,N_13763);
and U16002 (N_16002,N_13828,N_14396);
nor U16003 (N_16003,N_13756,N_13753);
xor U16004 (N_16004,N_14859,N_13882);
or U16005 (N_16005,N_14257,N_14592);
nand U16006 (N_16006,N_14536,N_14414);
nand U16007 (N_16007,N_14576,N_14603);
xnor U16008 (N_16008,N_14185,N_14666);
xnor U16009 (N_16009,N_14428,N_14061);
nor U16010 (N_16010,N_14368,N_14980);
nor U16011 (N_16011,N_14535,N_14294);
and U16012 (N_16012,N_14922,N_14852);
nand U16013 (N_16013,N_13779,N_14833);
or U16014 (N_16014,N_14778,N_14666);
xor U16015 (N_16015,N_14534,N_14248);
nor U16016 (N_16016,N_13822,N_14506);
nor U16017 (N_16017,N_14313,N_13993);
and U16018 (N_16018,N_14256,N_14162);
or U16019 (N_16019,N_14308,N_14820);
and U16020 (N_16020,N_14763,N_14087);
nor U16021 (N_16021,N_14162,N_14096);
nand U16022 (N_16022,N_14669,N_14388);
or U16023 (N_16023,N_14313,N_13966);
and U16024 (N_16024,N_14030,N_14333);
xnor U16025 (N_16025,N_14285,N_14508);
nor U16026 (N_16026,N_14649,N_13876);
or U16027 (N_16027,N_14461,N_14542);
or U16028 (N_16028,N_13934,N_14992);
nand U16029 (N_16029,N_14074,N_13864);
and U16030 (N_16030,N_14485,N_14517);
or U16031 (N_16031,N_13880,N_14766);
xnor U16032 (N_16032,N_13806,N_14474);
nor U16033 (N_16033,N_14756,N_14606);
nor U16034 (N_16034,N_14679,N_14272);
nand U16035 (N_16035,N_14413,N_13831);
xor U16036 (N_16036,N_14125,N_14977);
and U16037 (N_16037,N_13851,N_14620);
nor U16038 (N_16038,N_14149,N_14633);
or U16039 (N_16039,N_14697,N_14955);
nand U16040 (N_16040,N_14712,N_13842);
nor U16041 (N_16041,N_14323,N_14543);
and U16042 (N_16042,N_13844,N_13764);
xnor U16043 (N_16043,N_14442,N_14600);
and U16044 (N_16044,N_14936,N_14704);
and U16045 (N_16045,N_14531,N_13943);
nor U16046 (N_16046,N_14719,N_14523);
nand U16047 (N_16047,N_14782,N_14852);
xor U16048 (N_16048,N_14999,N_14183);
nand U16049 (N_16049,N_14689,N_14954);
xnor U16050 (N_16050,N_14657,N_14419);
nand U16051 (N_16051,N_14495,N_14306);
xnor U16052 (N_16052,N_14498,N_14295);
nand U16053 (N_16053,N_14101,N_13948);
xnor U16054 (N_16054,N_14424,N_14154);
xnor U16055 (N_16055,N_14649,N_14519);
xnor U16056 (N_16056,N_14261,N_14023);
nor U16057 (N_16057,N_14574,N_14492);
and U16058 (N_16058,N_14633,N_14604);
or U16059 (N_16059,N_14769,N_13845);
nand U16060 (N_16060,N_13750,N_13837);
nand U16061 (N_16061,N_14039,N_14873);
nand U16062 (N_16062,N_13935,N_14930);
or U16063 (N_16063,N_13799,N_14227);
nand U16064 (N_16064,N_14544,N_14606);
nand U16065 (N_16065,N_14366,N_13981);
and U16066 (N_16066,N_14136,N_14036);
nor U16067 (N_16067,N_14799,N_14660);
xor U16068 (N_16068,N_13827,N_14000);
nor U16069 (N_16069,N_14911,N_13931);
nor U16070 (N_16070,N_13862,N_14409);
nor U16071 (N_16071,N_14823,N_14970);
or U16072 (N_16072,N_14659,N_14887);
nor U16073 (N_16073,N_14189,N_14556);
nand U16074 (N_16074,N_14347,N_14499);
xnor U16075 (N_16075,N_14323,N_13766);
xor U16076 (N_16076,N_14027,N_14823);
and U16077 (N_16077,N_14825,N_14731);
and U16078 (N_16078,N_14354,N_14016);
xor U16079 (N_16079,N_14915,N_14447);
and U16080 (N_16080,N_14431,N_14889);
nand U16081 (N_16081,N_14580,N_14337);
nand U16082 (N_16082,N_14507,N_14202);
and U16083 (N_16083,N_13928,N_14089);
nor U16084 (N_16084,N_14586,N_13957);
nand U16085 (N_16085,N_14863,N_14912);
nor U16086 (N_16086,N_14957,N_14371);
and U16087 (N_16087,N_14741,N_14836);
or U16088 (N_16088,N_14386,N_14897);
nand U16089 (N_16089,N_14457,N_14957);
and U16090 (N_16090,N_14851,N_14286);
and U16091 (N_16091,N_14019,N_14547);
or U16092 (N_16092,N_14176,N_14364);
and U16093 (N_16093,N_14612,N_14719);
nand U16094 (N_16094,N_14828,N_14508);
nand U16095 (N_16095,N_13757,N_14889);
xnor U16096 (N_16096,N_14452,N_14911);
nor U16097 (N_16097,N_14267,N_14058);
and U16098 (N_16098,N_14581,N_14614);
and U16099 (N_16099,N_14981,N_14264);
and U16100 (N_16100,N_14815,N_14665);
nand U16101 (N_16101,N_14773,N_14406);
nor U16102 (N_16102,N_14084,N_14422);
nand U16103 (N_16103,N_14697,N_14296);
nor U16104 (N_16104,N_14419,N_14923);
and U16105 (N_16105,N_14889,N_14579);
nor U16106 (N_16106,N_14663,N_14592);
xor U16107 (N_16107,N_14075,N_14755);
or U16108 (N_16108,N_14363,N_14639);
and U16109 (N_16109,N_14835,N_14787);
nor U16110 (N_16110,N_14555,N_14826);
nor U16111 (N_16111,N_14131,N_14738);
xor U16112 (N_16112,N_14873,N_14897);
or U16113 (N_16113,N_13874,N_14218);
or U16114 (N_16114,N_14310,N_14888);
and U16115 (N_16115,N_14364,N_14789);
or U16116 (N_16116,N_14395,N_13912);
nand U16117 (N_16117,N_14916,N_14119);
or U16118 (N_16118,N_14152,N_13822);
and U16119 (N_16119,N_13974,N_14392);
xnor U16120 (N_16120,N_14581,N_14009);
nor U16121 (N_16121,N_14614,N_13764);
xor U16122 (N_16122,N_14748,N_14626);
nor U16123 (N_16123,N_14252,N_14804);
or U16124 (N_16124,N_14088,N_14294);
nor U16125 (N_16125,N_14848,N_14864);
nor U16126 (N_16126,N_14036,N_14062);
xnor U16127 (N_16127,N_13879,N_14368);
nor U16128 (N_16128,N_13910,N_14967);
nor U16129 (N_16129,N_14940,N_14749);
nand U16130 (N_16130,N_13877,N_13902);
nor U16131 (N_16131,N_14285,N_14873);
xor U16132 (N_16132,N_13859,N_13907);
nand U16133 (N_16133,N_14723,N_14041);
nand U16134 (N_16134,N_13834,N_14325);
and U16135 (N_16135,N_14207,N_13972);
or U16136 (N_16136,N_14181,N_14404);
or U16137 (N_16137,N_14641,N_14625);
xnor U16138 (N_16138,N_13954,N_14052);
or U16139 (N_16139,N_13989,N_13773);
or U16140 (N_16140,N_14818,N_14354);
nand U16141 (N_16141,N_14374,N_14107);
and U16142 (N_16142,N_14350,N_14661);
xnor U16143 (N_16143,N_14210,N_14521);
xor U16144 (N_16144,N_14379,N_14005);
nor U16145 (N_16145,N_13931,N_14148);
xor U16146 (N_16146,N_14130,N_14031);
xnor U16147 (N_16147,N_14172,N_14225);
or U16148 (N_16148,N_13897,N_13814);
nand U16149 (N_16149,N_14976,N_13988);
nand U16150 (N_16150,N_14059,N_14344);
nand U16151 (N_16151,N_14183,N_14361);
or U16152 (N_16152,N_14926,N_14732);
or U16153 (N_16153,N_14604,N_14819);
nand U16154 (N_16154,N_14525,N_13918);
nand U16155 (N_16155,N_14801,N_14759);
and U16156 (N_16156,N_14308,N_14026);
or U16157 (N_16157,N_14562,N_14121);
and U16158 (N_16158,N_14917,N_14772);
nand U16159 (N_16159,N_14856,N_14244);
or U16160 (N_16160,N_14935,N_13842);
and U16161 (N_16161,N_14602,N_14345);
or U16162 (N_16162,N_14173,N_14348);
nor U16163 (N_16163,N_14419,N_14457);
and U16164 (N_16164,N_14052,N_14709);
xor U16165 (N_16165,N_13874,N_13814);
or U16166 (N_16166,N_14366,N_14363);
xnor U16167 (N_16167,N_13952,N_13860);
xnor U16168 (N_16168,N_14574,N_14171);
nand U16169 (N_16169,N_13904,N_14033);
xnor U16170 (N_16170,N_14997,N_14343);
nor U16171 (N_16171,N_14574,N_13940);
and U16172 (N_16172,N_14306,N_14737);
nor U16173 (N_16173,N_14554,N_14801);
and U16174 (N_16174,N_13775,N_14311);
or U16175 (N_16175,N_14144,N_14695);
and U16176 (N_16176,N_14895,N_14322);
xnor U16177 (N_16177,N_14030,N_14405);
and U16178 (N_16178,N_14419,N_13986);
nand U16179 (N_16179,N_13773,N_13789);
nor U16180 (N_16180,N_14816,N_14195);
or U16181 (N_16181,N_14696,N_14494);
nand U16182 (N_16182,N_14835,N_13759);
nor U16183 (N_16183,N_14722,N_13915);
nand U16184 (N_16184,N_14497,N_14706);
and U16185 (N_16185,N_14155,N_14088);
and U16186 (N_16186,N_14772,N_14172);
or U16187 (N_16187,N_13996,N_14714);
or U16188 (N_16188,N_14032,N_14519);
xor U16189 (N_16189,N_14451,N_14556);
nand U16190 (N_16190,N_14189,N_14810);
and U16191 (N_16191,N_14502,N_13840);
or U16192 (N_16192,N_14691,N_14940);
and U16193 (N_16193,N_14789,N_13787);
xor U16194 (N_16194,N_13857,N_14076);
or U16195 (N_16195,N_14433,N_13889);
xor U16196 (N_16196,N_14179,N_13866);
and U16197 (N_16197,N_14915,N_13835);
xnor U16198 (N_16198,N_13990,N_14566);
nand U16199 (N_16199,N_13924,N_14241);
and U16200 (N_16200,N_14674,N_14949);
xnor U16201 (N_16201,N_13840,N_14130);
and U16202 (N_16202,N_14451,N_13971);
xnor U16203 (N_16203,N_14324,N_14990);
and U16204 (N_16204,N_14647,N_13851);
or U16205 (N_16205,N_14852,N_14417);
or U16206 (N_16206,N_14394,N_13953);
nor U16207 (N_16207,N_14933,N_14309);
nor U16208 (N_16208,N_14986,N_13922);
or U16209 (N_16209,N_14903,N_13940);
or U16210 (N_16210,N_14656,N_14232);
or U16211 (N_16211,N_14114,N_13985);
nor U16212 (N_16212,N_13894,N_14920);
and U16213 (N_16213,N_14635,N_14322);
xnor U16214 (N_16214,N_14779,N_14417);
xnor U16215 (N_16215,N_14271,N_14416);
and U16216 (N_16216,N_14142,N_14624);
and U16217 (N_16217,N_14855,N_14540);
nand U16218 (N_16218,N_14869,N_13956);
nor U16219 (N_16219,N_14350,N_14242);
or U16220 (N_16220,N_13882,N_14965);
nand U16221 (N_16221,N_13891,N_14627);
or U16222 (N_16222,N_14550,N_14098);
xnor U16223 (N_16223,N_14711,N_14948);
nand U16224 (N_16224,N_14120,N_14165);
nand U16225 (N_16225,N_14827,N_14523);
or U16226 (N_16226,N_13921,N_13763);
and U16227 (N_16227,N_14595,N_14657);
nand U16228 (N_16228,N_14031,N_14289);
or U16229 (N_16229,N_14644,N_14866);
and U16230 (N_16230,N_14145,N_14916);
nand U16231 (N_16231,N_14757,N_14074);
nor U16232 (N_16232,N_13932,N_14710);
nand U16233 (N_16233,N_13781,N_14916);
and U16234 (N_16234,N_14006,N_14023);
nand U16235 (N_16235,N_13780,N_14511);
or U16236 (N_16236,N_14822,N_14636);
nand U16237 (N_16237,N_14135,N_14662);
xnor U16238 (N_16238,N_14796,N_14215);
or U16239 (N_16239,N_14692,N_14094);
and U16240 (N_16240,N_13757,N_13989);
and U16241 (N_16241,N_14265,N_14204);
nand U16242 (N_16242,N_14578,N_14467);
nor U16243 (N_16243,N_14642,N_14715);
nand U16244 (N_16244,N_14788,N_14104);
and U16245 (N_16245,N_13912,N_14492);
or U16246 (N_16246,N_14440,N_14207);
nor U16247 (N_16247,N_13808,N_14603);
or U16248 (N_16248,N_14661,N_14700);
or U16249 (N_16249,N_13929,N_14872);
or U16250 (N_16250,N_15743,N_16069);
xnor U16251 (N_16251,N_15477,N_15409);
and U16252 (N_16252,N_16056,N_15322);
nand U16253 (N_16253,N_15786,N_15985);
and U16254 (N_16254,N_15083,N_15902);
nand U16255 (N_16255,N_15053,N_16162);
nor U16256 (N_16256,N_16124,N_15724);
nand U16257 (N_16257,N_15520,N_15126);
and U16258 (N_16258,N_15741,N_15887);
nor U16259 (N_16259,N_15058,N_15880);
nor U16260 (N_16260,N_15577,N_16220);
nor U16261 (N_16261,N_15745,N_15769);
nor U16262 (N_16262,N_16008,N_15450);
nor U16263 (N_16263,N_16027,N_15653);
or U16264 (N_16264,N_15181,N_15529);
xnor U16265 (N_16265,N_15495,N_16138);
nor U16266 (N_16266,N_16089,N_15262);
or U16267 (N_16267,N_16244,N_15390);
nor U16268 (N_16268,N_15562,N_15919);
nand U16269 (N_16269,N_15997,N_16209);
xor U16270 (N_16270,N_15899,N_15537);
or U16271 (N_16271,N_16018,N_15216);
nor U16272 (N_16272,N_15344,N_15736);
nand U16273 (N_16273,N_15479,N_15356);
nor U16274 (N_16274,N_15306,N_16107);
nor U16275 (N_16275,N_16043,N_15867);
and U16276 (N_16276,N_15145,N_15052);
xor U16277 (N_16277,N_15774,N_15313);
and U16278 (N_16278,N_16063,N_15473);
xnor U16279 (N_16279,N_15609,N_15418);
and U16280 (N_16280,N_15565,N_15631);
xnor U16281 (N_16281,N_15217,N_16144);
nand U16282 (N_16282,N_15290,N_15925);
and U16283 (N_16283,N_15698,N_15550);
xor U16284 (N_16284,N_15160,N_15253);
nor U16285 (N_16285,N_15267,N_15593);
nor U16286 (N_16286,N_15980,N_15664);
nand U16287 (N_16287,N_15911,N_15872);
nand U16288 (N_16288,N_16172,N_15699);
nand U16289 (N_16289,N_15048,N_15019);
nand U16290 (N_16290,N_15784,N_15326);
nor U16291 (N_16291,N_15033,N_15864);
nand U16292 (N_16292,N_16136,N_15352);
xor U16293 (N_16293,N_15511,N_15116);
and U16294 (N_16294,N_15594,N_15968);
or U16295 (N_16295,N_15431,N_16077);
or U16296 (N_16296,N_15333,N_16216);
xor U16297 (N_16297,N_15556,N_16071);
nand U16298 (N_16298,N_15121,N_15112);
nand U16299 (N_16299,N_15044,N_15242);
xor U16300 (N_16300,N_15885,N_16115);
nor U16301 (N_16301,N_15994,N_15739);
and U16302 (N_16302,N_15255,N_15122);
or U16303 (N_16303,N_15688,N_15028);
nor U16304 (N_16304,N_15041,N_16178);
or U16305 (N_16305,N_15336,N_15378);
and U16306 (N_16306,N_15965,N_15626);
nor U16307 (N_16307,N_15991,N_16053);
xor U16308 (N_16308,N_15377,N_16085);
and U16309 (N_16309,N_16134,N_15798);
xnor U16310 (N_16310,N_15568,N_15192);
nor U16311 (N_16311,N_15797,N_15913);
nand U16312 (N_16312,N_15815,N_16076);
nand U16313 (N_16313,N_15440,N_15690);
and U16314 (N_16314,N_15389,N_15092);
xor U16315 (N_16315,N_15627,N_15817);
or U16316 (N_16316,N_15951,N_15767);
nor U16317 (N_16317,N_15008,N_15304);
xor U16318 (N_16318,N_15931,N_15437);
or U16319 (N_16319,N_16098,N_15247);
and U16320 (N_16320,N_15413,N_15071);
nand U16321 (N_16321,N_15350,N_15227);
nand U16322 (N_16322,N_15410,N_15995);
xnor U16323 (N_16323,N_15775,N_16101);
and U16324 (N_16324,N_15927,N_15283);
nand U16325 (N_16325,N_15254,N_15307);
xor U16326 (N_16326,N_15882,N_15605);
or U16327 (N_16327,N_15497,N_15771);
or U16328 (N_16328,N_15792,N_15689);
xnor U16329 (N_16329,N_16030,N_16205);
nor U16330 (N_16330,N_15823,N_15737);
nor U16331 (N_16331,N_16066,N_15194);
nor U16332 (N_16332,N_15155,N_15671);
or U16333 (N_16333,N_16061,N_16102);
xnor U16334 (N_16334,N_15448,N_15579);
and U16335 (N_16335,N_15584,N_15123);
nand U16336 (N_16336,N_16149,N_15422);
nand U16337 (N_16337,N_15308,N_15848);
nor U16338 (N_16338,N_15235,N_15148);
or U16339 (N_16339,N_15607,N_16128);
nand U16340 (N_16340,N_15695,N_15660);
nor U16341 (N_16341,N_15528,N_15417);
nand U16342 (N_16342,N_15635,N_16150);
nand U16343 (N_16343,N_16094,N_15563);
and U16344 (N_16344,N_15040,N_15632);
nor U16345 (N_16345,N_15030,N_16086);
or U16346 (N_16346,N_15187,N_15655);
xnor U16347 (N_16347,N_15038,N_15500);
or U16348 (N_16348,N_15018,N_15481);
nor U16349 (N_16349,N_16013,N_16116);
nand U16350 (N_16350,N_15001,N_15049);
xor U16351 (N_16351,N_16233,N_15982);
and U16352 (N_16352,N_15270,N_15424);
and U16353 (N_16353,N_15000,N_15429);
nand U16354 (N_16354,N_15282,N_15299);
xnor U16355 (N_16355,N_16111,N_15938);
nand U16356 (N_16356,N_15130,N_15031);
nand U16357 (N_16357,N_15067,N_16169);
and U16358 (N_16358,N_15375,N_15933);
or U16359 (N_16359,N_16127,N_15170);
or U16360 (N_16360,N_15742,N_15293);
nor U16361 (N_16361,N_16230,N_15648);
nand U16362 (N_16362,N_15491,N_15929);
xor U16363 (N_16363,N_15989,N_15447);
nand U16364 (N_16364,N_15177,N_15022);
nor U16365 (N_16365,N_15858,N_15060);
or U16366 (N_16366,N_15171,N_15531);
or U16367 (N_16367,N_15534,N_16006);
or U16368 (N_16368,N_15677,N_15955);
xor U16369 (N_16369,N_15103,N_15538);
nand U16370 (N_16370,N_15638,N_15351);
and U16371 (N_16371,N_16218,N_15438);
and U16372 (N_16372,N_15611,N_15725);
nor U16373 (N_16373,N_15199,N_15761);
nand U16374 (N_16374,N_15156,N_15098);
or U16375 (N_16375,N_15603,N_15970);
nor U16376 (N_16376,N_15641,N_16040);
nand U16377 (N_16377,N_15824,N_15713);
nor U16378 (N_16378,N_15166,N_15813);
and U16379 (N_16379,N_15251,N_16106);
and U16380 (N_16380,N_15070,N_15339);
or U16381 (N_16381,N_16087,N_15361);
and U16382 (N_16382,N_15539,N_15596);
xnor U16383 (N_16383,N_16015,N_15915);
nand U16384 (N_16384,N_15812,N_15464);
or U16385 (N_16385,N_15893,N_15347);
and U16386 (N_16386,N_15907,N_16159);
and U16387 (N_16387,N_15667,N_16185);
or U16388 (N_16388,N_16122,N_15768);
and U16389 (N_16389,N_16227,N_15973);
or U16390 (N_16390,N_15753,N_15937);
or U16391 (N_16391,N_15394,N_15856);
nand U16392 (N_16392,N_16221,N_16133);
xnor U16393 (N_16393,N_15825,N_15958);
nand U16394 (N_16394,N_15622,N_15621);
nor U16395 (N_16395,N_16195,N_15346);
nand U16396 (N_16396,N_15969,N_15211);
and U16397 (N_16397,N_15708,N_15240);
and U16398 (N_16398,N_15328,N_15035);
and U16399 (N_16399,N_15583,N_15458);
nor U16400 (N_16400,N_15934,N_15633);
or U16401 (N_16401,N_16023,N_15486);
nand U16402 (N_16402,N_15248,N_15710);
xor U16403 (N_16403,N_15150,N_15644);
xor U16404 (N_16404,N_16206,N_15032);
nand U16405 (N_16405,N_15613,N_16219);
nand U16406 (N_16406,N_15136,N_15021);
or U16407 (N_16407,N_15666,N_15532);
xnor U16408 (N_16408,N_15023,N_15452);
nor U16409 (N_16409,N_15244,N_16224);
nand U16410 (N_16410,N_16100,N_15757);
or U16411 (N_16411,N_15966,N_15256);
nor U16412 (N_16412,N_16114,N_15017);
xnor U16413 (N_16413,N_15470,N_15780);
or U16414 (N_16414,N_15526,N_15209);
xnor U16415 (N_16415,N_15421,N_15920);
nand U16416 (N_16416,N_15056,N_15879);
nor U16417 (N_16417,N_15201,N_15066);
and U16418 (N_16418,N_16109,N_15206);
xnor U16419 (N_16419,N_15517,N_15950);
nand U16420 (N_16420,N_15158,N_15694);
nand U16421 (N_16421,N_15278,N_15914);
or U16422 (N_16422,N_15682,N_16225);
nor U16423 (N_16423,N_15546,N_15800);
and U16424 (N_16424,N_15237,N_15860);
nor U16425 (N_16425,N_15947,N_16062);
nand U16426 (N_16426,N_15013,N_16110);
and U16427 (N_16427,N_16075,N_15901);
nor U16428 (N_16428,N_15324,N_16155);
and U16429 (N_16429,N_15159,N_16131);
xor U16430 (N_16430,N_15898,N_15912);
and U16431 (N_16431,N_15161,N_16078);
nor U16432 (N_16432,N_15337,N_15803);
nand U16433 (N_16433,N_15547,N_15752);
nand U16434 (N_16434,N_15986,N_15503);
and U16435 (N_16435,N_15645,N_16234);
and U16436 (N_16436,N_15615,N_15099);
nand U16437 (N_16437,N_16037,N_15176);
or U16438 (N_16438,N_16117,N_15718);
nand U16439 (N_16439,N_15788,N_16044);
nor U16440 (N_16440,N_16207,N_15770);
or U16441 (N_16441,N_15175,N_15439);
nor U16442 (N_16442,N_15338,N_15600);
xnor U16443 (N_16443,N_16045,N_15364);
nand U16444 (N_16444,N_15445,N_15303);
nor U16445 (N_16445,N_15599,N_15818);
nor U16446 (N_16446,N_16092,N_15320);
nor U16447 (N_16447,N_15987,N_15670);
xor U16448 (N_16448,N_16095,N_15005);
nor U16449 (N_16449,N_16041,N_15095);
xor U16450 (N_16450,N_16164,N_16154);
nor U16451 (N_16451,N_15681,N_15238);
and U16452 (N_16452,N_15851,N_16072);
or U16453 (N_16453,N_15466,N_15129);
xor U16454 (N_16454,N_15407,N_16208);
and U16455 (N_16455,N_15395,N_15425);
nand U16456 (N_16456,N_15492,N_15379);
or U16457 (N_16457,N_15811,N_15212);
xor U16458 (N_16458,N_15077,N_15250);
nor U16459 (N_16459,N_15174,N_16046);
and U16460 (N_16460,N_15312,N_15488);
nand U16461 (N_16461,N_16187,N_15702);
nor U16462 (N_16462,N_15790,N_15229);
xor U16463 (N_16463,N_15459,N_16157);
or U16464 (N_16464,N_15665,N_16239);
xor U16465 (N_16465,N_15654,N_15524);
and U16466 (N_16466,N_16229,N_15456);
xnor U16467 (N_16467,N_15471,N_15513);
nor U16468 (N_16468,N_15266,N_15944);
or U16469 (N_16469,N_15432,N_15084);
nand U16470 (N_16470,N_15779,N_15243);
nor U16471 (N_16471,N_16033,N_16082);
xnor U16472 (N_16472,N_15016,N_15522);
or U16473 (N_16473,N_15288,N_15762);
nor U16474 (N_16474,N_15793,N_15311);
nor U16475 (N_16475,N_15285,N_15329);
nor U16476 (N_16476,N_15572,N_15449);
xnor U16477 (N_16477,N_15264,N_15372);
and U16478 (N_16478,N_15423,N_15142);
and U16479 (N_16479,N_15691,N_16147);
and U16480 (N_16480,N_16145,N_16104);
nand U16481 (N_16481,N_15334,N_15110);
xnor U16482 (N_16482,N_15383,N_15590);
nor U16483 (N_16483,N_15196,N_15153);
nand U16484 (N_16484,N_15214,N_16012);
xor U16485 (N_16485,N_15419,N_16212);
xnor U16486 (N_16486,N_15616,N_16241);
or U16487 (N_16487,N_15367,N_15263);
nand U16488 (N_16488,N_15575,N_15834);
and U16489 (N_16489,N_15086,N_15113);
nor U16490 (N_16490,N_15292,N_15623);
or U16491 (N_16491,N_16180,N_16024);
or U16492 (N_16492,N_15434,N_15003);
and U16493 (N_16493,N_15415,N_15839);
or U16494 (N_16494,N_15629,N_15904);
nor U16495 (N_16495,N_16140,N_15265);
nor U16496 (N_16496,N_15012,N_16158);
nand U16497 (N_16497,N_15140,N_15186);
xor U16498 (N_16498,N_15932,N_16148);
or U16499 (N_16499,N_16194,N_15853);
xor U16500 (N_16500,N_15705,N_16079);
xor U16501 (N_16501,N_16146,N_16065);
nor U16502 (N_16502,N_15223,N_16051);
nor U16503 (N_16503,N_15883,N_15543);
nor U16504 (N_16504,N_15802,N_15637);
xnor U16505 (N_16505,N_15772,N_15183);
xor U16506 (N_16506,N_16031,N_15791);
or U16507 (N_16507,N_15144,N_16074);
or U16508 (N_16508,N_15598,N_15412);
nand U16509 (N_16509,N_16231,N_15551);
nand U16510 (N_16510,N_16246,N_15921);
xor U16511 (N_16511,N_15972,N_15318);
nor U16512 (N_16512,N_15941,N_15465);
xor U16513 (N_16513,N_15198,N_15863);
or U16514 (N_16514,N_15760,N_15039);
xnor U16515 (N_16515,N_15386,N_16025);
xnor U16516 (N_16516,N_16123,N_15618);
xor U16517 (N_16517,N_15561,N_16168);
nand U16518 (N_16518,N_15544,N_15340);
and U16519 (N_16519,N_16237,N_15601);
or U16520 (N_16520,N_15435,N_15732);
nor U16521 (N_16521,N_15715,N_15795);
or U16522 (N_16522,N_15845,N_15549);
nor U16523 (N_16523,N_15809,N_15219);
nor U16524 (N_16524,N_15474,N_15273);
and U16525 (N_16525,N_15533,N_15178);
and U16526 (N_16526,N_15910,N_15894);
or U16527 (N_16527,N_15037,N_15696);
xor U16528 (N_16528,N_15147,N_15096);
nand U16529 (N_16529,N_15442,N_15873);
xnor U16530 (N_16530,N_15519,N_15085);
or U16531 (N_16531,N_15990,N_16038);
nand U16532 (N_16532,N_16059,N_15015);
or U16533 (N_16533,N_15309,N_15202);
nor U16534 (N_16534,N_15707,N_15081);
nor U16535 (N_16535,N_15119,N_15400);
and U16536 (N_16536,N_15487,N_15485);
nand U16537 (N_16537,N_16113,N_15193);
nor U16538 (N_16538,N_15010,N_15781);
or U16539 (N_16539,N_15570,N_16047);
nand U16540 (N_16540,N_15874,N_15200);
or U16541 (N_16541,N_16055,N_15636);
xor U16542 (N_16542,N_15298,N_15639);
nor U16543 (N_16543,N_15179,N_16105);
and U16544 (N_16544,N_15428,N_15744);
nor U16545 (N_16545,N_15173,N_15408);
xnor U16546 (N_16546,N_15974,N_15230);
and U16547 (N_16547,N_16236,N_15763);
or U16548 (N_16548,N_16068,N_15109);
or U16549 (N_16549,N_15135,N_15020);
or U16550 (N_16550,N_15054,N_16151);
xor U16551 (N_16551,N_15079,N_15108);
xnor U16552 (N_16552,N_15963,N_15068);
xnor U16553 (N_16553,N_16139,N_15335);
nor U16554 (N_16554,N_16039,N_15755);
nor U16555 (N_16555,N_16248,N_16120);
xnor U16556 (N_16556,N_15365,N_15133);
nand U16557 (N_16557,N_15062,N_16193);
nor U16558 (N_16558,N_15317,N_15844);
or U16559 (N_16559,N_15234,N_15512);
or U16560 (N_16560,N_15646,N_15801);
nor U16561 (N_16561,N_16058,N_16016);
and U16562 (N_16562,N_16067,N_15029);
and U16563 (N_16563,N_15567,N_15891);
or U16564 (N_16564,N_15816,N_15617);
or U16565 (N_16565,N_15806,N_15560);
nor U16566 (N_16566,N_15711,N_16081);
nand U16567 (N_16567,N_15906,N_16213);
xor U16568 (N_16568,N_15499,N_16001);
nor U16569 (N_16569,N_16232,N_15405);
or U16570 (N_16570,N_15097,N_15960);
nor U16571 (N_16571,N_16245,N_15945);
nand U16572 (N_16572,N_15117,N_15859);
or U16573 (N_16573,N_15002,N_15131);
nand U16574 (N_16574,N_15731,N_15369);
and U16575 (N_16575,N_16064,N_16184);
nor U16576 (N_16576,N_15063,N_15162);
xor U16577 (N_16577,N_15011,N_16215);
nand U16578 (N_16578,N_15861,N_15354);
xnor U16579 (N_16579,N_15443,N_15475);
or U16580 (N_16580,N_15895,N_15709);
and U16581 (N_16581,N_16093,N_15125);
and U16582 (N_16582,N_15535,N_15905);
or U16583 (N_16583,N_15703,N_15586);
nand U16584 (N_16584,N_16009,N_15956);
and U16585 (N_16585,N_15362,N_16021);
and U16586 (N_16586,N_15436,N_15257);
and U16587 (N_16587,N_16247,N_16090);
nand U16588 (N_16588,N_15685,N_15576);
and U16589 (N_16589,N_15404,N_15735);
nor U16590 (N_16590,N_15983,N_15239);
xor U16591 (N_16591,N_15280,N_16235);
or U16592 (N_16592,N_15870,N_15589);
and U16593 (N_16593,N_15523,N_16129);
nand U16594 (N_16594,N_15558,N_15924);
and U16595 (N_16595,N_15074,N_15917);
and U16596 (N_16596,N_15889,N_15357);
and U16597 (N_16597,N_15608,N_15420);
and U16598 (N_16598,N_15542,N_15050);
and U16599 (N_16599,N_16143,N_15676);
and U16600 (N_16600,N_15909,N_16174);
nand U16601 (N_16601,N_16202,N_16189);
nor U16602 (N_16602,N_16142,N_16108);
or U16603 (N_16603,N_15402,N_15167);
nand U16604 (N_16604,N_15678,N_15953);
nand U16605 (N_16605,N_16011,N_15215);
nor U16606 (N_16606,N_16125,N_15294);
xnor U16607 (N_16607,N_15722,N_16049);
or U16608 (N_16608,N_15082,N_15051);
nor U16609 (N_16609,N_16060,N_15114);
xor U16610 (N_16610,N_15004,N_15876);
xnor U16611 (N_16611,N_15172,N_15669);
or U16612 (N_16612,N_15249,N_15540);
nand U16613 (N_16613,N_16183,N_15507);
or U16614 (N_16614,N_15843,N_15988);
nor U16615 (N_16615,N_15047,N_15451);
nor U16616 (N_16616,N_15191,N_15684);
nor U16617 (N_16617,N_15325,N_15961);
or U16618 (N_16618,N_15620,N_15319);
nand U16619 (N_16619,N_15749,N_15930);
or U16620 (N_16620,N_15730,N_15647);
and U16621 (N_16621,N_15782,N_16176);
or U16622 (N_16622,N_15076,N_15559);
nand U16623 (N_16623,N_15700,N_15602);
or U16624 (N_16624,N_15808,N_15675);
xor U16625 (N_16625,N_15805,N_16050);
or U16626 (N_16626,N_15628,N_15832);
xor U16627 (N_16627,N_16014,N_16199);
nor U16628 (N_16628,N_15042,N_15430);
and U16629 (N_16629,N_15461,N_15182);
and U16630 (N_16630,N_15279,N_15733);
nor U16631 (N_16631,N_15588,N_15124);
nor U16632 (N_16632,N_15276,N_15469);
and U16633 (N_16633,N_15692,N_15157);
or U16634 (N_16634,N_16200,N_15830);
nor U16635 (N_16635,N_15726,N_15064);
or U16636 (N_16636,N_15224,N_15127);
and U16637 (N_16637,N_15866,N_15025);
and U16638 (N_16638,N_15332,N_15530);
or U16639 (N_16639,N_15472,N_15587);
xor U16640 (N_16640,N_15065,N_15414);
nand U16641 (N_16641,N_16137,N_15154);
nor U16642 (N_16642,N_16119,N_15948);
nand U16643 (N_16643,N_15766,N_15446);
nand U16644 (N_16644,N_15979,N_16249);
nand U16645 (N_16645,N_15258,N_15785);
nand U16646 (N_16646,N_15069,N_15120);
or U16647 (N_16647,N_15773,N_15463);
and U16648 (N_16648,N_15087,N_15923);
and U16649 (N_16649,N_15518,N_16073);
nor U16650 (N_16650,N_15261,N_15978);
nor U16651 (N_16651,N_16026,N_15850);
nand U16652 (N_16652,N_16022,N_15075);
xnor U16653 (N_16653,N_15807,N_15833);
nand U16654 (N_16654,N_15504,N_15197);
nor U16655 (N_16655,N_15959,N_15716);
and U16656 (N_16656,N_16019,N_15441);
xnor U16657 (N_16657,N_15819,N_15205);
xor U16658 (N_16658,N_15467,N_15935);
nand U16659 (N_16659,N_15869,N_15776);
nand U16660 (N_16660,N_15847,N_15396);
nand U16661 (N_16661,N_15926,N_15536);
nand U16662 (N_16662,N_16135,N_15521);
xnor U16663 (N_16663,N_15759,N_16161);
xnor U16664 (N_16664,N_15661,N_15454);
xor U16665 (N_16665,N_15525,N_15720);
and U16666 (N_16666,N_15218,N_15604);
or U16667 (N_16667,N_16198,N_16211);
nand U16668 (N_16668,N_15846,N_16173);
nor U16669 (N_16669,N_16091,N_15168);
nand U16670 (N_16670,N_15836,N_15094);
or U16671 (N_16671,N_15679,N_15835);
xor U16672 (N_16672,N_15165,N_15489);
xnor U16673 (N_16673,N_15026,N_15107);
and U16674 (N_16674,N_15650,N_15295);
xor U16675 (N_16675,N_15360,N_16191);
and U16676 (N_16676,N_15105,N_15634);
nor U16677 (N_16677,N_15756,N_15277);
nor U16678 (N_16678,N_15697,N_15043);
nor U16679 (N_16679,N_15574,N_15624);
and U16680 (N_16680,N_16080,N_15406);
and U16681 (N_16681,N_15349,N_15680);
nand U16682 (N_16682,N_15509,N_15385);
xor U16683 (N_16683,N_15208,N_15592);
nor U16684 (N_16684,N_15185,N_15829);
nor U16685 (N_16685,N_15892,N_15490);
xor U16686 (N_16686,N_15009,N_15348);
nand U16687 (N_16687,N_15401,N_15100);
nand U16688 (N_16688,N_15640,N_15453);
and U16689 (N_16689,N_15188,N_15241);
xnor U16690 (N_16690,N_16166,N_15663);
or U16691 (N_16691,N_15721,N_16217);
nor U16692 (N_16692,N_15291,N_15221);
and U16693 (N_16693,N_15706,N_15842);
xor U16694 (N_16694,N_15180,N_15139);
nor U16695 (N_16695,N_15838,N_15992);
nand U16696 (N_16696,N_15034,N_15297);
nor U16697 (N_16697,N_16242,N_15566);
nor U16698 (N_16698,N_15246,N_15210);
and U16699 (N_16699,N_15723,N_15233);
xor U16700 (N_16700,N_15686,N_16160);
and U16701 (N_16701,N_16054,N_15552);
and U16702 (N_16702,N_15046,N_15928);
nand U16703 (N_16703,N_15169,N_15651);
nand U16704 (N_16704,N_16048,N_16036);
or U16705 (N_16705,N_15496,N_15286);
xor U16706 (N_16706,N_15061,N_15841);
nor U16707 (N_16707,N_16029,N_15922);
nand U16708 (N_16708,N_15976,N_16070);
nor U16709 (N_16709,N_15750,N_15310);
xnor U16710 (N_16710,N_15143,N_15896);
nand U16711 (N_16711,N_16096,N_15810);
nor U16712 (N_16712,N_15939,N_15137);
xor U16713 (N_16713,N_16228,N_15527);
or U16714 (N_16714,N_15388,N_16171);
nand U16715 (N_16715,N_16099,N_15738);
or U16716 (N_16716,N_15977,N_15088);
nand U16717 (N_16717,N_15146,N_15510);
nand U16718 (N_16718,N_15036,N_15787);
nand U16719 (N_16719,N_16084,N_15203);
and U16720 (N_16720,N_16175,N_16188);
nor U16721 (N_16721,N_15506,N_15149);
xor U16722 (N_16722,N_15998,N_15478);
xnor U16723 (N_16723,N_15382,N_15614);
nand U16724 (N_16724,N_15220,N_15564);
or U16725 (N_16725,N_15658,N_15498);
nand U16726 (N_16726,N_15881,N_15865);
and U16727 (N_16727,N_15837,N_16156);
xnor U16728 (N_16728,N_15748,N_15952);
or U16729 (N_16729,N_15946,N_16177);
nor U16730 (N_16730,N_15740,N_15118);
xnor U16731 (N_16731,N_15368,N_15854);
nor U16732 (N_16732,N_16003,N_15444);
xnor U16733 (N_16733,N_16057,N_15072);
xor U16734 (N_16734,N_16152,N_15101);
xor U16735 (N_16735,N_15821,N_16197);
or U16736 (N_16736,N_15804,N_16052);
nor U16737 (N_16737,N_15555,N_15245);
nor U16738 (N_16738,N_16112,N_15305);
nor U16739 (N_16739,N_15943,N_15515);
nand U16740 (N_16740,N_15416,N_15252);
nor U16741 (N_16741,N_15975,N_16132);
xnor U16742 (N_16742,N_16222,N_15073);
nand U16743 (N_16743,N_16126,N_15799);
xor U16744 (N_16744,N_15849,N_16165);
nor U16745 (N_16745,N_15996,N_15852);
nand U16746 (N_16746,N_15457,N_15502);
xor U16747 (N_16747,N_15656,N_15758);
nor U16748 (N_16748,N_15964,N_15272);
nand U16749 (N_16749,N_16226,N_15163);
nor U16750 (N_16750,N_15057,N_15548);
nor U16751 (N_16751,N_15897,N_15232);
nor U16752 (N_16752,N_15330,N_15314);
and U16753 (N_16753,N_15501,N_15204);
and U16754 (N_16754,N_15342,N_15657);
xnor U16755 (N_16755,N_15289,N_16163);
nor U16756 (N_16756,N_15619,N_15376);
xnor U16757 (N_16757,N_16192,N_15747);
nor U16758 (N_16758,N_15358,N_15236);
nor U16759 (N_16759,N_15794,N_16201);
nor U16760 (N_16760,N_15455,N_15719);
xor U16761 (N_16761,N_16004,N_15152);
nor U16762 (N_16762,N_15207,N_15693);
nand U16763 (N_16763,N_16017,N_15302);
nor U16764 (N_16764,N_15886,N_15585);
nand U16765 (N_16765,N_15226,N_16010);
xnor U16766 (N_16766,N_15541,N_15301);
and U16767 (N_16767,N_15765,N_15091);
xor U16768 (N_16768,N_15345,N_15397);
nand U16769 (N_16769,N_16000,N_15778);
nor U16770 (N_16770,N_15476,N_15132);
nor U16771 (N_16771,N_15260,N_15268);
or U16772 (N_16772,N_16181,N_15373);
and U16773 (N_16773,N_15916,N_15391);
nor U16774 (N_16774,N_15999,N_15093);
or U16775 (N_16775,N_15796,N_15433);
nand U16776 (N_16776,N_15878,N_15918);
nand U16777 (N_16777,N_15908,N_15746);
xor U16778 (N_16778,N_15981,N_15826);
and U16779 (N_16779,N_15890,N_15840);
nor U16780 (N_16780,N_16121,N_16210);
nand U16781 (N_16781,N_15371,N_15427);
nand U16782 (N_16782,N_15936,N_15967);
nor U16783 (N_16783,N_15275,N_15827);
nor U16784 (N_16784,N_15014,N_15597);
nand U16785 (N_16785,N_15580,N_16141);
xor U16786 (N_16786,N_15828,N_15630);
or U16787 (N_16787,N_15734,N_15764);
nand U16788 (N_16788,N_15387,N_15341);
nand U16789 (N_16789,N_15553,N_15059);
or U16790 (N_16790,N_16243,N_15228);
nand U16791 (N_16791,N_15259,N_16118);
and U16792 (N_16792,N_15399,N_15353);
nor U16793 (N_16793,N_15321,N_15189);
or U16794 (N_16794,N_16182,N_16196);
xor U16795 (N_16795,N_16007,N_15006);
or U16796 (N_16796,N_15355,N_16032);
and U16797 (N_16797,N_15729,N_15777);
nor U16798 (N_16798,N_15460,N_15184);
nor U16799 (N_16799,N_15190,N_15557);
and U16800 (N_16800,N_15868,N_15662);
xor U16801 (N_16801,N_15717,N_15569);
nor U16802 (N_16802,N_15673,N_16002);
nor U16803 (N_16803,N_15871,N_15483);
nor U16804 (N_16804,N_16153,N_16179);
and U16805 (N_16805,N_15393,N_15111);
nor U16806 (N_16806,N_15751,N_15296);
nand U16807 (N_16807,N_15582,N_15089);
and U16808 (N_16808,N_15683,N_16204);
and U16809 (N_16809,N_15606,N_15134);
or U16810 (N_16810,N_15141,N_15649);
and U16811 (N_16811,N_15494,N_15855);
or U16812 (N_16812,N_15225,N_15573);
nand U16813 (N_16813,N_15115,N_15954);
nor U16814 (N_16814,N_15480,N_16190);
and U16815 (N_16815,N_15045,N_15151);
or U16816 (N_16816,N_16028,N_15957);
nand U16817 (N_16817,N_15701,N_15659);
and U16818 (N_16818,N_15610,N_15381);
and U16819 (N_16819,N_15578,N_15195);
or U16820 (N_16820,N_15754,N_15090);
xor U16821 (N_16821,N_15468,N_16223);
nor U16822 (N_16822,N_15940,N_15643);
xor U16823 (N_16823,N_15392,N_16167);
xor U16824 (N_16824,N_15222,N_15591);
or U16825 (N_16825,N_15595,N_15728);
or U16826 (N_16826,N_15359,N_16042);
xnor U16827 (N_16827,N_15323,N_16238);
and U16828 (N_16828,N_15514,N_16005);
and U16829 (N_16829,N_16214,N_15138);
or U16830 (N_16830,N_15984,N_15687);
and U16831 (N_16831,N_15363,N_16020);
nor U16832 (N_16832,N_15287,N_15789);
xnor U16833 (N_16833,N_15080,N_15213);
or U16834 (N_16834,N_15398,N_15505);
and U16835 (N_16835,N_15426,N_15374);
nand U16836 (N_16836,N_16097,N_15949);
and U16837 (N_16837,N_15104,N_15102);
nor U16838 (N_16838,N_15857,N_16034);
nand U16839 (N_16839,N_15888,N_15462);
nor U16840 (N_16840,N_15484,N_15712);
xnor U16841 (N_16841,N_15411,N_16103);
or U16842 (N_16842,N_15900,N_15642);
and U16843 (N_16843,N_15316,N_16240);
xor U16844 (N_16844,N_15581,N_16130);
nand U16845 (N_16845,N_15674,N_15814);
and U16846 (N_16846,N_15993,N_15820);
nand U16847 (N_16847,N_15831,N_15274);
or U16848 (N_16848,N_15007,N_15055);
nand U16849 (N_16849,N_15612,N_15884);
and U16850 (N_16850,N_15271,N_16203);
or U16851 (N_16851,N_15625,N_15281);
nand U16852 (N_16852,N_15327,N_15024);
or U16853 (N_16853,N_15384,N_15942);
or U16854 (N_16854,N_15231,N_16088);
nand U16855 (N_16855,N_15078,N_15668);
xor U16856 (N_16856,N_15516,N_15128);
or U16857 (N_16857,N_15903,N_15284);
nor U16858 (N_16858,N_15366,N_16083);
xor U16859 (N_16859,N_15380,N_15877);
nand U16860 (N_16860,N_15164,N_15822);
or U16861 (N_16861,N_15652,N_15554);
nor U16862 (N_16862,N_15672,N_15106);
and U16863 (N_16863,N_15545,N_16170);
nor U16864 (N_16864,N_15971,N_15862);
xnor U16865 (N_16865,N_15343,N_15962);
nand U16866 (N_16866,N_16035,N_15704);
or U16867 (N_16867,N_15315,N_15875);
and U16868 (N_16868,N_15493,N_15727);
or U16869 (N_16869,N_15482,N_15300);
nand U16870 (N_16870,N_15714,N_15508);
or U16871 (N_16871,N_15783,N_15331);
and U16872 (N_16872,N_16186,N_15269);
and U16873 (N_16873,N_15027,N_15370);
nor U16874 (N_16874,N_15403,N_15571);
or U16875 (N_16875,N_15183,N_15263);
nand U16876 (N_16876,N_16119,N_16166);
xnor U16877 (N_16877,N_15027,N_15476);
nor U16878 (N_16878,N_15745,N_15248);
xor U16879 (N_16879,N_15627,N_15591);
xnor U16880 (N_16880,N_15730,N_16020);
or U16881 (N_16881,N_15965,N_15240);
or U16882 (N_16882,N_15299,N_15683);
nor U16883 (N_16883,N_15956,N_15636);
nor U16884 (N_16884,N_15826,N_15699);
and U16885 (N_16885,N_15465,N_15030);
nand U16886 (N_16886,N_15705,N_15901);
xnor U16887 (N_16887,N_15717,N_15558);
or U16888 (N_16888,N_15647,N_16217);
nor U16889 (N_16889,N_15583,N_15432);
xor U16890 (N_16890,N_15789,N_15715);
or U16891 (N_16891,N_15437,N_15432);
xnor U16892 (N_16892,N_15277,N_16007);
or U16893 (N_16893,N_15245,N_15242);
nand U16894 (N_16894,N_16054,N_16053);
nor U16895 (N_16895,N_15907,N_15644);
and U16896 (N_16896,N_15219,N_15877);
xor U16897 (N_16897,N_16145,N_16178);
and U16898 (N_16898,N_16039,N_16199);
xnor U16899 (N_16899,N_15542,N_16102);
nand U16900 (N_16900,N_15207,N_15009);
or U16901 (N_16901,N_15711,N_15467);
xnor U16902 (N_16902,N_15982,N_15915);
nor U16903 (N_16903,N_15305,N_15016);
or U16904 (N_16904,N_15531,N_16135);
nand U16905 (N_16905,N_15014,N_15213);
xor U16906 (N_16906,N_16074,N_15883);
xor U16907 (N_16907,N_15591,N_16045);
xnor U16908 (N_16908,N_15816,N_15564);
or U16909 (N_16909,N_15972,N_15745);
nand U16910 (N_16910,N_15590,N_15247);
and U16911 (N_16911,N_15366,N_15564);
or U16912 (N_16912,N_15280,N_15173);
or U16913 (N_16913,N_16216,N_15296);
or U16914 (N_16914,N_15557,N_15756);
or U16915 (N_16915,N_15941,N_16101);
nand U16916 (N_16916,N_16040,N_15147);
xor U16917 (N_16917,N_15900,N_15200);
xor U16918 (N_16918,N_16065,N_15658);
or U16919 (N_16919,N_15603,N_15210);
or U16920 (N_16920,N_15126,N_15844);
nand U16921 (N_16921,N_15580,N_15445);
nand U16922 (N_16922,N_15490,N_15296);
nor U16923 (N_16923,N_15231,N_15567);
nor U16924 (N_16924,N_15234,N_15317);
and U16925 (N_16925,N_15576,N_15074);
nor U16926 (N_16926,N_15723,N_15621);
or U16927 (N_16927,N_16145,N_15778);
and U16928 (N_16928,N_15241,N_15011);
nand U16929 (N_16929,N_15033,N_16096);
nand U16930 (N_16930,N_15647,N_15855);
and U16931 (N_16931,N_15499,N_15694);
nand U16932 (N_16932,N_15117,N_15005);
xnor U16933 (N_16933,N_15773,N_16122);
or U16934 (N_16934,N_15959,N_15211);
or U16935 (N_16935,N_16187,N_16030);
xnor U16936 (N_16936,N_15178,N_15041);
nor U16937 (N_16937,N_15153,N_15015);
nand U16938 (N_16938,N_15041,N_16106);
xnor U16939 (N_16939,N_15317,N_15544);
and U16940 (N_16940,N_15155,N_15367);
xnor U16941 (N_16941,N_15153,N_15125);
and U16942 (N_16942,N_15482,N_15179);
nand U16943 (N_16943,N_16210,N_15782);
and U16944 (N_16944,N_16234,N_15570);
and U16945 (N_16945,N_15102,N_16183);
xor U16946 (N_16946,N_15015,N_15903);
nor U16947 (N_16947,N_16164,N_15117);
and U16948 (N_16948,N_16186,N_16224);
nand U16949 (N_16949,N_15383,N_15191);
nand U16950 (N_16950,N_15058,N_15885);
nor U16951 (N_16951,N_15943,N_15067);
or U16952 (N_16952,N_15199,N_16203);
xor U16953 (N_16953,N_15015,N_15228);
and U16954 (N_16954,N_15557,N_15160);
nand U16955 (N_16955,N_15169,N_15678);
or U16956 (N_16956,N_16233,N_15593);
and U16957 (N_16957,N_15493,N_15061);
xnor U16958 (N_16958,N_15258,N_15010);
or U16959 (N_16959,N_15215,N_15607);
and U16960 (N_16960,N_15720,N_15954);
xor U16961 (N_16961,N_15943,N_15707);
and U16962 (N_16962,N_15605,N_15812);
nand U16963 (N_16963,N_15029,N_15847);
and U16964 (N_16964,N_15395,N_15151);
nor U16965 (N_16965,N_15807,N_15547);
and U16966 (N_16966,N_15933,N_15147);
nor U16967 (N_16967,N_16000,N_15390);
nor U16968 (N_16968,N_15539,N_15766);
nand U16969 (N_16969,N_15699,N_15338);
or U16970 (N_16970,N_15888,N_15313);
nand U16971 (N_16971,N_15100,N_15835);
xor U16972 (N_16972,N_15564,N_16121);
or U16973 (N_16973,N_15405,N_15765);
or U16974 (N_16974,N_15227,N_16085);
or U16975 (N_16975,N_16232,N_15855);
nor U16976 (N_16976,N_15272,N_15878);
nand U16977 (N_16977,N_15965,N_15367);
and U16978 (N_16978,N_15456,N_15292);
nor U16979 (N_16979,N_15878,N_15928);
or U16980 (N_16980,N_15052,N_15866);
nand U16981 (N_16981,N_15215,N_15016);
or U16982 (N_16982,N_15690,N_15255);
and U16983 (N_16983,N_15742,N_15727);
nand U16984 (N_16984,N_15576,N_15784);
nand U16985 (N_16985,N_16173,N_15950);
nand U16986 (N_16986,N_15891,N_15853);
nor U16987 (N_16987,N_15245,N_15842);
xnor U16988 (N_16988,N_15791,N_15211);
xnor U16989 (N_16989,N_15215,N_16221);
nor U16990 (N_16990,N_15347,N_15867);
and U16991 (N_16991,N_16246,N_16004);
and U16992 (N_16992,N_16178,N_15524);
or U16993 (N_16993,N_16144,N_15805);
nand U16994 (N_16994,N_15945,N_16056);
or U16995 (N_16995,N_15066,N_15873);
xnor U16996 (N_16996,N_15117,N_16192);
or U16997 (N_16997,N_15307,N_15501);
nand U16998 (N_16998,N_15908,N_15130);
nand U16999 (N_16999,N_15708,N_15274);
xor U17000 (N_17000,N_15791,N_15444);
xnor U17001 (N_17001,N_15575,N_16063);
xnor U17002 (N_17002,N_15571,N_15164);
or U17003 (N_17003,N_16065,N_15366);
nor U17004 (N_17004,N_15393,N_15250);
nor U17005 (N_17005,N_15408,N_15421);
nand U17006 (N_17006,N_15592,N_15540);
and U17007 (N_17007,N_15454,N_16082);
nand U17008 (N_17008,N_15884,N_15887);
or U17009 (N_17009,N_15233,N_15460);
and U17010 (N_17010,N_16187,N_15119);
nand U17011 (N_17011,N_15561,N_15566);
nand U17012 (N_17012,N_15882,N_15572);
nand U17013 (N_17013,N_15540,N_15490);
nor U17014 (N_17014,N_15322,N_15517);
nand U17015 (N_17015,N_15502,N_15709);
or U17016 (N_17016,N_15804,N_15250);
and U17017 (N_17017,N_15630,N_15331);
nand U17018 (N_17018,N_15125,N_15994);
nand U17019 (N_17019,N_15228,N_15531);
xor U17020 (N_17020,N_15376,N_15239);
or U17021 (N_17021,N_15670,N_16151);
nand U17022 (N_17022,N_15951,N_15005);
or U17023 (N_17023,N_15963,N_15238);
and U17024 (N_17024,N_15680,N_15311);
and U17025 (N_17025,N_15401,N_15080);
or U17026 (N_17026,N_15100,N_15301);
nor U17027 (N_17027,N_15916,N_15425);
or U17028 (N_17028,N_15523,N_15884);
nor U17029 (N_17029,N_15223,N_15197);
nand U17030 (N_17030,N_15276,N_15255);
nand U17031 (N_17031,N_15273,N_16242);
nor U17032 (N_17032,N_15342,N_16130);
xor U17033 (N_17033,N_15073,N_15593);
or U17034 (N_17034,N_15495,N_15935);
nor U17035 (N_17035,N_15393,N_15666);
or U17036 (N_17036,N_15875,N_16097);
nor U17037 (N_17037,N_15483,N_15106);
or U17038 (N_17038,N_15344,N_15109);
and U17039 (N_17039,N_15664,N_15572);
nand U17040 (N_17040,N_15509,N_15882);
nand U17041 (N_17041,N_16034,N_15237);
and U17042 (N_17042,N_15033,N_15598);
nor U17043 (N_17043,N_15702,N_15064);
or U17044 (N_17044,N_15561,N_15503);
nand U17045 (N_17045,N_15297,N_15861);
nor U17046 (N_17046,N_15139,N_15157);
nor U17047 (N_17047,N_15589,N_15771);
xor U17048 (N_17048,N_15803,N_15868);
nand U17049 (N_17049,N_16204,N_16048);
nand U17050 (N_17050,N_15116,N_16168);
xor U17051 (N_17051,N_15070,N_15543);
or U17052 (N_17052,N_15744,N_16171);
or U17053 (N_17053,N_15253,N_15004);
and U17054 (N_17054,N_15581,N_15628);
xor U17055 (N_17055,N_15146,N_15390);
or U17056 (N_17056,N_16097,N_16118);
nor U17057 (N_17057,N_15485,N_15840);
or U17058 (N_17058,N_16138,N_15790);
nor U17059 (N_17059,N_15172,N_15662);
nand U17060 (N_17060,N_15053,N_16103);
nand U17061 (N_17061,N_15422,N_15721);
nand U17062 (N_17062,N_15638,N_16173);
nor U17063 (N_17063,N_15899,N_15536);
or U17064 (N_17064,N_15545,N_15869);
nand U17065 (N_17065,N_15740,N_15389);
nor U17066 (N_17066,N_15547,N_15660);
and U17067 (N_17067,N_15817,N_16122);
nand U17068 (N_17068,N_15762,N_15111);
xnor U17069 (N_17069,N_15850,N_16174);
nor U17070 (N_17070,N_15396,N_15177);
and U17071 (N_17071,N_15629,N_16138);
nor U17072 (N_17072,N_15520,N_15378);
xnor U17073 (N_17073,N_15812,N_15909);
xor U17074 (N_17074,N_16112,N_15651);
and U17075 (N_17075,N_16212,N_15268);
nor U17076 (N_17076,N_15604,N_16028);
nor U17077 (N_17077,N_15397,N_16247);
nor U17078 (N_17078,N_15483,N_15273);
nand U17079 (N_17079,N_15457,N_15908);
or U17080 (N_17080,N_15621,N_15581);
nor U17081 (N_17081,N_15873,N_16190);
and U17082 (N_17082,N_16178,N_15956);
xor U17083 (N_17083,N_15493,N_15507);
or U17084 (N_17084,N_15063,N_15314);
or U17085 (N_17085,N_15488,N_15593);
xor U17086 (N_17086,N_15803,N_15077);
xor U17087 (N_17087,N_15864,N_16075);
or U17088 (N_17088,N_15473,N_15666);
nor U17089 (N_17089,N_15781,N_15602);
nand U17090 (N_17090,N_15229,N_15051);
nor U17091 (N_17091,N_15934,N_15413);
xnor U17092 (N_17092,N_15375,N_15817);
nor U17093 (N_17093,N_15005,N_16104);
or U17094 (N_17094,N_15778,N_15560);
xor U17095 (N_17095,N_15615,N_15178);
or U17096 (N_17096,N_15831,N_15380);
and U17097 (N_17097,N_15663,N_15842);
or U17098 (N_17098,N_15385,N_15340);
or U17099 (N_17099,N_15423,N_16099);
or U17100 (N_17100,N_15581,N_15016);
xor U17101 (N_17101,N_15405,N_15631);
or U17102 (N_17102,N_15253,N_16079);
xnor U17103 (N_17103,N_15790,N_16084);
nor U17104 (N_17104,N_15367,N_16156);
and U17105 (N_17105,N_15571,N_15070);
nand U17106 (N_17106,N_15019,N_15230);
and U17107 (N_17107,N_15950,N_16077);
or U17108 (N_17108,N_15333,N_15037);
xor U17109 (N_17109,N_16234,N_15972);
xnor U17110 (N_17110,N_15722,N_16105);
nand U17111 (N_17111,N_16202,N_15045);
nor U17112 (N_17112,N_15861,N_15908);
nand U17113 (N_17113,N_15216,N_16185);
or U17114 (N_17114,N_15980,N_15738);
and U17115 (N_17115,N_15812,N_15152);
nand U17116 (N_17116,N_15421,N_15541);
nor U17117 (N_17117,N_15050,N_15780);
xor U17118 (N_17118,N_15280,N_15858);
nor U17119 (N_17119,N_15085,N_15183);
nor U17120 (N_17120,N_15055,N_16208);
nor U17121 (N_17121,N_15252,N_15892);
nand U17122 (N_17122,N_15806,N_15448);
and U17123 (N_17123,N_15533,N_15600);
nor U17124 (N_17124,N_15906,N_16084);
and U17125 (N_17125,N_15934,N_15528);
or U17126 (N_17126,N_15906,N_15789);
nand U17127 (N_17127,N_15211,N_15212);
xor U17128 (N_17128,N_15721,N_16116);
and U17129 (N_17129,N_16141,N_16134);
and U17130 (N_17130,N_16223,N_16237);
or U17131 (N_17131,N_16070,N_15099);
nand U17132 (N_17132,N_15104,N_15512);
xor U17133 (N_17133,N_15874,N_15843);
nand U17134 (N_17134,N_16138,N_15599);
or U17135 (N_17135,N_16178,N_15434);
and U17136 (N_17136,N_16156,N_15864);
and U17137 (N_17137,N_15418,N_15851);
nand U17138 (N_17138,N_15419,N_15756);
nor U17139 (N_17139,N_15053,N_15448);
nor U17140 (N_17140,N_16045,N_15851);
or U17141 (N_17141,N_15392,N_15866);
xnor U17142 (N_17142,N_16143,N_15130);
xnor U17143 (N_17143,N_15145,N_15482);
nand U17144 (N_17144,N_15937,N_15311);
nand U17145 (N_17145,N_15394,N_15429);
or U17146 (N_17146,N_15159,N_15218);
nand U17147 (N_17147,N_15470,N_15022);
nor U17148 (N_17148,N_15220,N_16203);
or U17149 (N_17149,N_15198,N_15094);
and U17150 (N_17150,N_15824,N_15520);
or U17151 (N_17151,N_15255,N_15607);
and U17152 (N_17152,N_15331,N_16230);
xor U17153 (N_17153,N_16042,N_16009);
or U17154 (N_17154,N_15435,N_16216);
or U17155 (N_17155,N_15955,N_15185);
nand U17156 (N_17156,N_15807,N_15498);
or U17157 (N_17157,N_15379,N_16230);
nor U17158 (N_17158,N_15964,N_15234);
nand U17159 (N_17159,N_15494,N_16113);
and U17160 (N_17160,N_15512,N_15708);
xor U17161 (N_17161,N_15236,N_15023);
xnor U17162 (N_17162,N_16164,N_15725);
nor U17163 (N_17163,N_15892,N_16164);
and U17164 (N_17164,N_15065,N_15102);
nor U17165 (N_17165,N_15027,N_15991);
xnor U17166 (N_17166,N_15068,N_15541);
nor U17167 (N_17167,N_15770,N_15114);
and U17168 (N_17168,N_15087,N_15352);
and U17169 (N_17169,N_15575,N_15810);
and U17170 (N_17170,N_15711,N_15132);
nor U17171 (N_17171,N_15448,N_15691);
or U17172 (N_17172,N_15925,N_15274);
and U17173 (N_17173,N_15231,N_15781);
nand U17174 (N_17174,N_16018,N_15782);
nor U17175 (N_17175,N_15805,N_15506);
or U17176 (N_17176,N_16091,N_15444);
or U17177 (N_17177,N_15696,N_15048);
xnor U17178 (N_17178,N_16182,N_16108);
or U17179 (N_17179,N_15034,N_15863);
xnor U17180 (N_17180,N_15767,N_16230);
and U17181 (N_17181,N_16226,N_16212);
nor U17182 (N_17182,N_15355,N_15285);
nor U17183 (N_17183,N_15057,N_16243);
nand U17184 (N_17184,N_15005,N_15494);
nor U17185 (N_17185,N_15278,N_15857);
xor U17186 (N_17186,N_15991,N_15023);
and U17187 (N_17187,N_15338,N_15175);
xnor U17188 (N_17188,N_15532,N_15291);
or U17189 (N_17189,N_15923,N_16215);
nor U17190 (N_17190,N_15600,N_15112);
and U17191 (N_17191,N_15144,N_16097);
nand U17192 (N_17192,N_15661,N_15522);
or U17193 (N_17193,N_15399,N_15801);
xnor U17194 (N_17194,N_15252,N_15865);
nor U17195 (N_17195,N_15255,N_15182);
xor U17196 (N_17196,N_15346,N_16165);
nand U17197 (N_17197,N_15029,N_16129);
nand U17198 (N_17198,N_15848,N_15335);
nor U17199 (N_17199,N_15814,N_15216);
nand U17200 (N_17200,N_16225,N_15482);
and U17201 (N_17201,N_16120,N_15385);
nand U17202 (N_17202,N_15664,N_15084);
or U17203 (N_17203,N_15713,N_15886);
nor U17204 (N_17204,N_15071,N_15087);
or U17205 (N_17205,N_15493,N_15604);
or U17206 (N_17206,N_15122,N_15466);
xor U17207 (N_17207,N_15977,N_15476);
or U17208 (N_17208,N_15464,N_15187);
nand U17209 (N_17209,N_16173,N_16142);
and U17210 (N_17210,N_15615,N_15508);
xor U17211 (N_17211,N_16200,N_15190);
nand U17212 (N_17212,N_15496,N_15944);
nor U17213 (N_17213,N_15539,N_15091);
xor U17214 (N_17214,N_16096,N_15537);
xor U17215 (N_17215,N_15928,N_16172);
nor U17216 (N_17216,N_15722,N_15297);
xnor U17217 (N_17217,N_15705,N_16049);
xnor U17218 (N_17218,N_15765,N_15088);
nand U17219 (N_17219,N_15531,N_15324);
nand U17220 (N_17220,N_15750,N_15535);
nor U17221 (N_17221,N_16196,N_16145);
and U17222 (N_17222,N_15480,N_15440);
nor U17223 (N_17223,N_15335,N_15584);
nand U17224 (N_17224,N_15450,N_15355);
nor U17225 (N_17225,N_15195,N_15757);
nor U17226 (N_17226,N_15357,N_16174);
or U17227 (N_17227,N_15175,N_15598);
or U17228 (N_17228,N_15999,N_15957);
or U17229 (N_17229,N_15486,N_15636);
nand U17230 (N_17230,N_15890,N_15346);
xor U17231 (N_17231,N_15679,N_15291);
or U17232 (N_17232,N_15111,N_15508);
nand U17233 (N_17233,N_15475,N_15400);
or U17234 (N_17234,N_16025,N_15780);
xnor U17235 (N_17235,N_15223,N_15348);
or U17236 (N_17236,N_16230,N_15360);
nor U17237 (N_17237,N_15364,N_16150);
nor U17238 (N_17238,N_15656,N_15310);
nor U17239 (N_17239,N_16074,N_15592);
or U17240 (N_17240,N_15599,N_15162);
nand U17241 (N_17241,N_15245,N_16210);
nor U17242 (N_17242,N_15591,N_15327);
and U17243 (N_17243,N_15431,N_15153);
nand U17244 (N_17244,N_15499,N_15570);
or U17245 (N_17245,N_15303,N_15662);
nor U17246 (N_17246,N_15447,N_16087);
xnor U17247 (N_17247,N_15908,N_15538);
nand U17248 (N_17248,N_15327,N_15158);
nor U17249 (N_17249,N_15627,N_15075);
nor U17250 (N_17250,N_15416,N_15299);
and U17251 (N_17251,N_15231,N_15538);
xnor U17252 (N_17252,N_15179,N_15863);
and U17253 (N_17253,N_15574,N_15893);
nand U17254 (N_17254,N_15799,N_15455);
xnor U17255 (N_17255,N_15983,N_15245);
or U17256 (N_17256,N_15869,N_15004);
or U17257 (N_17257,N_16156,N_15309);
and U17258 (N_17258,N_15192,N_15254);
or U17259 (N_17259,N_15080,N_15119);
nand U17260 (N_17260,N_15935,N_15153);
xnor U17261 (N_17261,N_15245,N_15742);
nand U17262 (N_17262,N_15037,N_15516);
nand U17263 (N_17263,N_15835,N_15902);
or U17264 (N_17264,N_16019,N_15903);
and U17265 (N_17265,N_15814,N_15829);
and U17266 (N_17266,N_15085,N_15091);
xnor U17267 (N_17267,N_15539,N_15353);
nand U17268 (N_17268,N_15175,N_15467);
nor U17269 (N_17269,N_15098,N_15552);
and U17270 (N_17270,N_15435,N_15479);
nand U17271 (N_17271,N_16107,N_15026);
or U17272 (N_17272,N_15431,N_15126);
and U17273 (N_17273,N_16022,N_16076);
or U17274 (N_17274,N_16132,N_15972);
nor U17275 (N_17275,N_16218,N_15126);
xor U17276 (N_17276,N_16246,N_15376);
and U17277 (N_17277,N_15046,N_15688);
or U17278 (N_17278,N_15698,N_15731);
nand U17279 (N_17279,N_15623,N_16061);
and U17280 (N_17280,N_15343,N_15573);
nand U17281 (N_17281,N_15226,N_16244);
and U17282 (N_17282,N_15950,N_16200);
xnor U17283 (N_17283,N_15673,N_15601);
nand U17284 (N_17284,N_15437,N_15604);
nor U17285 (N_17285,N_15896,N_15550);
nand U17286 (N_17286,N_15009,N_15295);
or U17287 (N_17287,N_15320,N_15193);
xor U17288 (N_17288,N_15631,N_15104);
or U17289 (N_17289,N_16063,N_15615);
or U17290 (N_17290,N_15611,N_15148);
xor U17291 (N_17291,N_15542,N_15084);
or U17292 (N_17292,N_15060,N_16232);
nand U17293 (N_17293,N_15446,N_16010);
or U17294 (N_17294,N_15348,N_15834);
nand U17295 (N_17295,N_16007,N_15644);
or U17296 (N_17296,N_15843,N_15710);
and U17297 (N_17297,N_15799,N_15256);
nor U17298 (N_17298,N_15313,N_15191);
or U17299 (N_17299,N_16015,N_15411);
xor U17300 (N_17300,N_15181,N_16190);
nor U17301 (N_17301,N_15809,N_15799);
nand U17302 (N_17302,N_15818,N_15438);
and U17303 (N_17303,N_15094,N_15068);
nor U17304 (N_17304,N_15791,N_15829);
and U17305 (N_17305,N_15741,N_15389);
xor U17306 (N_17306,N_15226,N_15837);
xor U17307 (N_17307,N_16078,N_15873);
nand U17308 (N_17308,N_15707,N_15332);
and U17309 (N_17309,N_15741,N_15792);
or U17310 (N_17310,N_16051,N_15452);
and U17311 (N_17311,N_16193,N_15696);
and U17312 (N_17312,N_15486,N_15731);
nand U17313 (N_17313,N_15809,N_15080);
nand U17314 (N_17314,N_15385,N_15232);
or U17315 (N_17315,N_15998,N_15177);
and U17316 (N_17316,N_15490,N_15426);
xnor U17317 (N_17317,N_15859,N_15966);
and U17318 (N_17318,N_15028,N_15031);
and U17319 (N_17319,N_15262,N_15563);
nand U17320 (N_17320,N_15794,N_15925);
nand U17321 (N_17321,N_15197,N_16058);
nor U17322 (N_17322,N_15641,N_15502);
nor U17323 (N_17323,N_15599,N_15001);
nor U17324 (N_17324,N_15642,N_15183);
and U17325 (N_17325,N_15135,N_15862);
or U17326 (N_17326,N_15119,N_15513);
nand U17327 (N_17327,N_15153,N_15785);
nor U17328 (N_17328,N_15089,N_15691);
nand U17329 (N_17329,N_15182,N_15787);
or U17330 (N_17330,N_15380,N_15133);
nor U17331 (N_17331,N_16033,N_16153);
xnor U17332 (N_17332,N_15738,N_15175);
or U17333 (N_17333,N_16159,N_15672);
or U17334 (N_17334,N_15849,N_15514);
nor U17335 (N_17335,N_15864,N_15683);
nand U17336 (N_17336,N_15405,N_15490);
and U17337 (N_17337,N_15607,N_15023);
xnor U17338 (N_17338,N_15564,N_15737);
or U17339 (N_17339,N_16076,N_16016);
nand U17340 (N_17340,N_15963,N_15580);
and U17341 (N_17341,N_15897,N_15940);
and U17342 (N_17342,N_15133,N_15630);
xor U17343 (N_17343,N_15629,N_15190);
nand U17344 (N_17344,N_15980,N_16243);
or U17345 (N_17345,N_16038,N_15499);
nor U17346 (N_17346,N_16018,N_15476);
and U17347 (N_17347,N_15504,N_15360);
xor U17348 (N_17348,N_15737,N_16158);
nand U17349 (N_17349,N_15159,N_16017);
and U17350 (N_17350,N_15765,N_15582);
nand U17351 (N_17351,N_15298,N_15024);
or U17352 (N_17352,N_16204,N_15585);
or U17353 (N_17353,N_16083,N_15610);
and U17354 (N_17354,N_15917,N_15559);
or U17355 (N_17355,N_15808,N_15487);
nand U17356 (N_17356,N_16086,N_15914);
or U17357 (N_17357,N_15908,N_15655);
and U17358 (N_17358,N_15413,N_15058);
xnor U17359 (N_17359,N_16030,N_15653);
xnor U17360 (N_17360,N_15001,N_15288);
nand U17361 (N_17361,N_15276,N_15805);
nand U17362 (N_17362,N_16002,N_16046);
nor U17363 (N_17363,N_15935,N_15374);
xnor U17364 (N_17364,N_15431,N_15566);
or U17365 (N_17365,N_15018,N_15488);
nand U17366 (N_17366,N_15308,N_16222);
xnor U17367 (N_17367,N_15873,N_16079);
nand U17368 (N_17368,N_15814,N_15495);
nor U17369 (N_17369,N_15041,N_15599);
xnor U17370 (N_17370,N_15706,N_15965);
nand U17371 (N_17371,N_15941,N_16159);
nand U17372 (N_17372,N_15100,N_15595);
nand U17373 (N_17373,N_15227,N_15231);
nor U17374 (N_17374,N_15138,N_15267);
or U17375 (N_17375,N_15023,N_15744);
nor U17376 (N_17376,N_15518,N_15095);
nand U17377 (N_17377,N_15203,N_15773);
nand U17378 (N_17378,N_15698,N_15792);
and U17379 (N_17379,N_15694,N_15474);
or U17380 (N_17380,N_15171,N_16222);
xor U17381 (N_17381,N_15233,N_15819);
nand U17382 (N_17382,N_16021,N_15699);
or U17383 (N_17383,N_16113,N_15608);
or U17384 (N_17384,N_15621,N_16244);
nand U17385 (N_17385,N_15083,N_15599);
and U17386 (N_17386,N_15216,N_16031);
nor U17387 (N_17387,N_15306,N_15971);
nor U17388 (N_17388,N_15961,N_15820);
or U17389 (N_17389,N_16140,N_15532);
xnor U17390 (N_17390,N_15490,N_15144);
nand U17391 (N_17391,N_16052,N_15889);
xnor U17392 (N_17392,N_15479,N_16025);
nor U17393 (N_17393,N_15702,N_16051);
nand U17394 (N_17394,N_15385,N_15782);
or U17395 (N_17395,N_16085,N_15644);
and U17396 (N_17396,N_15372,N_15476);
or U17397 (N_17397,N_15519,N_16046);
xnor U17398 (N_17398,N_15781,N_15493);
xnor U17399 (N_17399,N_15186,N_15264);
nor U17400 (N_17400,N_16000,N_15096);
xor U17401 (N_17401,N_15324,N_15000);
xnor U17402 (N_17402,N_15201,N_15766);
nor U17403 (N_17403,N_16247,N_15170);
or U17404 (N_17404,N_15456,N_15285);
or U17405 (N_17405,N_16136,N_15180);
and U17406 (N_17406,N_15025,N_15455);
and U17407 (N_17407,N_16203,N_16010);
nor U17408 (N_17408,N_16009,N_16165);
nor U17409 (N_17409,N_15193,N_16076);
and U17410 (N_17410,N_15384,N_15717);
nor U17411 (N_17411,N_15880,N_15627);
nand U17412 (N_17412,N_16248,N_15051);
nand U17413 (N_17413,N_15028,N_15511);
and U17414 (N_17414,N_15814,N_16000);
and U17415 (N_17415,N_16122,N_15110);
or U17416 (N_17416,N_15776,N_16155);
nor U17417 (N_17417,N_15973,N_16138);
nand U17418 (N_17418,N_15105,N_16235);
and U17419 (N_17419,N_16020,N_15173);
nand U17420 (N_17420,N_15756,N_15384);
nand U17421 (N_17421,N_15574,N_15459);
nor U17422 (N_17422,N_15377,N_15991);
or U17423 (N_17423,N_15845,N_15419);
nor U17424 (N_17424,N_15941,N_15473);
or U17425 (N_17425,N_16205,N_15308);
and U17426 (N_17426,N_15182,N_16184);
xor U17427 (N_17427,N_15306,N_15127);
nand U17428 (N_17428,N_15387,N_15754);
xnor U17429 (N_17429,N_15831,N_15738);
nor U17430 (N_17430,N_15802,N_15348);
nand U17431 (N_17431,N_16200,N_15794);
and U17432 (N_17432,N_15107,N_15418);
or U17433 (N_17433,N_15246,N_15616);
and U17434 (N_17434,N_15027,N_15255);
nor U17435 (N_17435,N_16209,N_15114);
and U17436 (N_17436,N_16122,N_15415);
xnor U17437 (N_17437,N_16215,N_15550);
or U17438 (N_17438,N_15627,N_15703);
nand U17439 (N_17439,N_16184,N_15037);
and U17440 (N_17440,N_15237,N_15597);
nand U17441 (N_17441,N_15460,N_15485);
nor U17442 (N_17442,N_15827,N_16123);
xnor U17443 (N_17443,N_16064,N_15317);
xnor U17444 (N_17444,N_15787,N_15465);
nand U17445 (N_17445,N_15667,N_15399);
nand U17446 (N_17446,N_16249,N_15082);
and U17447 (N_17447,N_15735,N_15256);
or U17448 (N_17448,N_15874,N_15388);
xor U17449 (N_17449,N_15346,N_15272);
and U17450 (N_17450,N_15978,N_15352);
xor U17451 (N_17451,N_15900,N_15045);
nor U17452 (N_17452,N_15525,N_15372);
and U17453 (N_17453,N_15892,N_15864);
nand U17454 (N_17454,N_16121,N_15960);
and U17455 (N_17455,N_16017,N_15115);
nor U17456 (N_17456,N_15035,N_15669);
and U17457 (N_17457,N_15330,N_15015);
and U17458 (N_17458,N_15369,N_16108);
xnor U17459 (N_17459,N_15064,N_15935);
nand U17460 (N_17460,N_15213,N_15875);
and U17461 (N_17461,N_15604,N_15878);
nor U17462 (N_17462,N_15122,N_15492);
xor U17463 (N_17463,N_15726,N_15145);
and U17464 (N_17464,N_15942,N_15604);
xnor U17465 (N_17465,N_15741,N_15689);
and U17466 (N_17466,N_16063,N_15897);
nand U17467 (N_17467,N_15357,N_15728);
nand U17468 (N_17468,N_15038,N_15798);
and U17469 (N_17469,N_15041,N_15764);
or U17470 (N_17470,N_15017,N_16061);
and U17471 (N_17471,N_15539,N_15527);
nor U17472 (N_17472,N_16175,N_15447);
and U17473 (N_17473,N_16203,N_15538);
nor U17474 (N_17474,N_15360,N_15076);
nand U17475 (N_17475,N_16072,N_16083);
xnor U17476 (N_17476,N_15001,N_15545);
nor U17477 (N_17477,N_15532,N_15998);
or U17478 (N_17478,N_16210,N_15837);
nor U17479 (N_17479,N_15436,N_15663);
nor U17480 (N_17480,N_15572,N_15875);
xor U17481 (N_17481,N_15233,N_16191);
nor U17482 (N_17482,N_15458,N_16100);
and U17483 (N_17483,N_15861,N_16016);
xor U17484 (N_17484,N_15228,N_15920);
nand U17485 (N_17485,N_15877,N_16234);
or U17486 (N_17486,N_15373,N_15149);
nand U17487 (N_17487,N_15761,N_16140);
or U17488 (N_17488,N_15265,N_15306);
and U17489 (N_17489,N_15286,N_16195);
nand U17490 (N_17490,N_15873,N_15378);
nor U17491 (N_17491,N_15406,N_15588);
and U17492 (N_17492,N_15030,N_15393);
or U17493 (N_17493,N_15129,N_15319);
nand U17494 (N_17494,N_15364,N_15081);
xnor U17495 (N_17495,N_16165,N_16174);
or U17496 (N_17496,N_15959,N_15752);
and U17497 (N_17497,N_16092,N_15281);
nand U17498 (N_17498,N_15829,N_15772);
and U17499 (N_17499,N_15879,N_15540);
xnor U17500 (N_17500,N_17381,N_16748);
or U17501 (N_17501,N_17090,N_16798);
and U17502 (N_17502,N_16419,N_17086);
nor U17503 (N_17503,N_16953,N_17398);
nor U17504 (N_17504,N_17261,N_17068);
or U17505 (N_17505,N_16653,N_16918);
and U17506 (N_17506,N_16837,N_16478);
nor U17507 (N_17507,N_17229,N_16860);
xnor U17508 (N_17508,N_16904,N_17298);
xnor U17509 (N_17509,N_17383,N_16335);
or U17510 (N_17510,N_16611,N_16888);
or U17511 (N_17511,N_16381,N_16267);
and U17512 (N_17512,N_16483,N_17001);
nor U17513 (N_17513,N_16965,N_16972);
and U17514 (N_17514,N_17319,N_17313);
nand U17515 (N_17515,N_17131,N_16537);
nand U17516 (N_17516,N_16818,N_16557);
or U17517 (N_17517,N_16664,N_16411);
xnor U17518 (N_17518,N_17278,N_16944);
nand U17519 (N_17519,N_16598,N_16574);
or U17520 (N_17520,N_16449,N_16722);
nand U17521 (N_17521,N_16539,N_16415);
nor U17522 (N_17522,N_17253,N_16609);
nor U17523 (N_17523,N_16811,N_17394);
nor U17524 (N_17524,N_17129,N_16887);
xnor U17525 (N_17525,N_17374,N_16641);
nand U17526 (N_17526,N_17152,N_17225);
nand U17527 (N_17527,N_16399,N_17162);
nor U17528 (N_17528,N_16690,N_17296);
nor U17529 (N_17529,N_16289,N_17244);
or U17530 (N_17530,N_16558,N_17339);
xnor U17531 (N_17531,N_16422,N_17489);
xor U17532 (N_17532,N_16864,N_16951);
or U17533 (N_17533,N_16568,N_16750);
or U17534 (N_17534,N_16548,N_17186);
and U17535 (N_17535,N_17156,N_17017);
or U17536 (N_17536,N_16746,N_16317);
and U17537 (N_17537,N_16886,N_16346);
nor U17538 (N_17538,N_16662,N_16266);
or U17539 (N_17539,N_16355,N_16742);
and U17540 (N_17540,N_17228,N_16783);
nand U17541 (N_17541,N_16785,N_16708);
or U17542 (N_17542,N_17290,N_16626);
nor U17543 (N_17543,N_17214,N_16545);
or U17544 (N_17544,N_16424,N_16627);
xor U17545 (N_17545,N_16356,N_16554);
nand U17546 (N_17546,N_17392,N_16648);
and U17547 (N_17547,N_16352,N_16853);
and U17548 (N_17548,N_17440,N_16529);
nand U17549 (N_17549,N_16561,N_17443);
xnor U17550 (N_17550,N_16398,N_17027);
nor U17551 (N_17551,N_16271,N_16949);
or U17552 (N_17552,N_16337,N_17144);
nand U17553 (N_17553,N_16591,N_17200);
and U17554 (N_17554,N_17456,N_16890);
xor U17555 (N_17555,N_17273,N_16931);
and U17556 (N_17556,N_16897,N_17187);
nor U17557 (N_17557,N_17277,N_16547);
and U17558 (N_17558,N_17410,N_16300);
nor U17559 (N_17559,N_16929,N_16276);
and U17560 (N_17560,N_16606,N_16534);
nand U17561 (N_17561,N_16987,N_16768);
and U17562 (N_17562,N_17437,N_17060);
nand U17563 (N_17563,N_16787,N_16391);
nor U17564 (N_17564,N_16971,N_17424);
nand U17565 (N_17565,N_16582,N_16821);
or U17566 (N_17566,N_16333,N_16520);
xnor U17567 (N_17567,N_17262,N_17176);
and U17568 (N_17568,N_17400,N_17128);
nand U17569 (N_17569,N_16556,N_16644);
and U17570 (N_17570,N_16601,N_16717);
or U17571 (N_17571,N_17105,N_16402);
nand U17572 (N_17572,N_17478,N_16714);
xnor U17573 (N_17573,N_17356,N_16417);
xnor U17574 (N_17574,N_17430,N_16675);
and U17575 (N_17575,N_16859,N_16621);
nand U17576 (N_17576,N_17472,N_16268);
nor U17577 (N_17577,N_16567,N_17243);
xnor U17578 (N_17578,N_17488,N_16366);
xor U17579 (N_17579,N_17093,N_16321);
or U17580 (N_17580,N_16993,N_16470);
nor U17581 (N_17581,N_17352,N_16677);
or U17582 (N_17582,N_16286,N_17391);
xnor U17583 (N_17583,N_16964,N_16631);
xor U17584 (N_17584,N_16939,N_17486);
nor U17585 (N_17585,N_17153,N_16790);
or U17586 (N_17586,N_16998,N_16867);
or U17587 (N_17587,N_17107,N_17238);
nand U17588 (N_17588,N_16585,N_16728);
nor U17589 (N_17589,N_17476,N_17155);
nand U17590 (N_17590,N_17405,N_17401);
nor U17591 (N_17591,N_17118,N_16516);
nand U17592 (N_17592,N_17124,N_16438);
nand U17593 (N_17593,N_16476,N_16928);
and U17594 (N_17594,N_16846,N_17444);
nand U17595 (N_17595,N_17188,N_16819);
xor U17596 (N_17596,N_17497,N_16880);
nand U17597 (N_17597,N_16423,N_16786);
xor U17598 (N_17598,N_16498,N_17442);
or U17599 (N_17599,N_17191,N_17211);
nor U17600 (N_17600,N_16313,N_16553);
or U17601 (N_17601,N_16581,N_16418);
or U17602 (N_17602,N_17378,N_16699);
nor U17603 (N_17603,N_16408,N_17032);
nor U17604 (N_17604,N_16795,N_17487);
xor U17605 (N_17605,N_16353,N_17414);
and U17606 (N_17606,N_17283,N_17431);
nand U17607 (N_17607,N_16633,N_16979);
and U17608 (N_17608,N_16632,N_16397);
and U17609 (N_17609,N_16265,N_16459);
or U17610 (N_17610,N_17425,N_16608);
and U17611 (N_17611,N_16405,N_17030);
or U17612 (N_17612,N_17172,N_17037);
and U17613 (N_17613,N_17012,N_17451);
or U17614 (N_17614,N_16685,N_16958);
nand U17615 (N_17615,N_17455,N_16761);
or U17616 (N_17616,N_16946,N_16889);
or U17617 (N_17617,N_17077,N_16385);
and U17618 (N_17618,N_16436,N_16839);
nor U17619 (N_17619,N_17227,N_16511);
xnor U17620 (N_17620,N_16920,N_16715);
nor U17621 (N_17621,N_16977,N_17035);
xnor U17622 (N_17622,N_17458,N_17138);
and U17623 (N_17623,N_16395,N_16320);
xor U17624 (N_17624,N_17098,N_16776);
or U17625 (N_17625,N_16260,N_16610);
xnor U17626 (N_17626,N_17119,N_17370);
nand U17627 (N_17627,N_16517,N_17023);
nor U17628 (N_17628,N_17239,N_16940);
xnor U17629 (N_17629,N_17483,N_17242);
nor U17630 (N_17630,N_16603,N_17372);
nor U17631 (N_17631,N_16713,N_16532);
nand U17632 (N_17632,N_16272,N_16309);
nor U17633 (N_17633,N_17047,N_16596);
or U17634 (N_17634,N_17469,N_17323);
nand U17635 (N_17635,N_17146,N_16661);
nor U17636 (N_17636,N_17452,N_16844);
or U17637 (N_17637,N_17226,N_17484);
or U17638 (N_17638,N_16341,N_17168);
nand U17639 (N_17639,N_16723,N_16737);
nand U17640 (N_17640,N_17259,N_16872);
xnor U17641 (N_17641,N_16310,N_16325);
xor U17642 (N_17642,N_16925,N_17382);
nor U17643 (N_17643,N_16629,N_16826);
nor U17644 (N_17644,N_16825,N_17385);
nand U17645 (N_17645,N_17390,N_16968);
nor U17646 (N_17646,N_16809,N_17065);
xnor U17647 (N_17647,N_17288,N_16784);
nor U17648 (N_17648,N_17429,N_16814);
or U17649 (N_17649,N_16584,N_17071);
or U17650 (N_17650,N_17005,N_17348);
or U17651 (N_17651,N_16756,N_17457);
nand U17652 (N_17652,N_16796,N_17018);
or U17653 (N_17653,N_16383,N_16995);
and U17654 (N_17654,N_17280,N_17088);
or U17655 (N_17655,N_17208,N_16451);
and U17656 (N_17656,N_16669,N_16643);
or U17657 (N_17657,N_17494,N_17240);
nand U17658 (N_17658,N_16635,N_17263);
nor U17659 (N_17659,N_16707,N_17059);
and U17660 (N_17660,N_16503,N_16425);
nor U17661 (N_17661,N_16850,N_17013);
nor U17662 (N_17662,N_16515,N_16698);
or U17663 (N_17663,N_17206,N_16463);
nor U17664 (N_17664,N_16565,N_16280);
nor U17665 (N_17665,N_17022,N_16299);
or U17666 (N_17666,N_16740,N_17083);
and U17667 (N_17667,N_16816,N_17493);
or U17668 (N_17668,N_16474,N_17117);
and U17669 (N_17669,N_16358,N_16579);
xnor U17670 (N_17670,N_17380,N_16736);
nand U17671 (N_17671,N_16878,N_16832);
or U17672 (N_17672,N_16681,N_16588);
or U17673 (N_17673,N_17351,N_16453);
nand U17674 (N_17674,N_16739,N_16583);
nand U17675 (N_17675,N_16440,N_16540);
nor U17676 (N_17676,N_16646,N_16657);
or U17677 (N_17677,N_17078,N_16901);
nand U17678 (N_17678,N_16854,N_17407);
or U17679 (N_17679,N_17250,N_16763);
nor U17680 (N_17680,N_16650,N_16710);
nor U17681 (N_17681,N_16492,N_16573);
nor U17682 (N_17682,N_17435,N_16360);
and U17683 (N_17683,N_17041,N_16834);
nor U17684 (N_17684,N_16465,N_16663);
xnor U17685 (N_17685,N_17171,N_16909);
nor U17686 (N_17686,N_17289,N_17066);
xnor U17687 (N_17687,N_16917,N_16343);
nor U17688 (N_17688,N_17123,N_16523);
xor U17689 (N_17689,N_16820,N_16807);
or U17690 (N_17690,N_17219,N_16559);
xor U17691 (N_17691,N_17441,N_16528);
xnor U17692 (N_17692,N_16347,N_17257);
or U17693 (N_17693,N_17415,N_16509);
and U17694 (N_17694,N_16817,N_16803);
or U17695 (N_17695,N_17194,N_17293);
and U17696 (N_17696,N_16308,N_16883);
xor U17697 (N_17697,N_16702,N_17079);
and U17698 (N_17698,N_17040,N_16334);
and U17699 (N_17699,N_16665,N_16893);
xor U17700 (N_17700,N_17073,N_17492);
xnor U17701 (N_17701,N_16259,N_16873);
nand U17702 (N_17702,N_16607,N_17334);
or U17703 (N_17703,N_16857,N_16255);
xor U17704 (N_17704,N_17204,N_17048);
and U17705 (N_17705,N_16913,N_16412);
or U17706 (N_17706,N_16871,N_17076);
or U17707 (N_17707,N_16876,N_16769);
xor U17708 (N_17708,N_16638,N_16342);
and U17709 (N_17709,N_17338,N_17254);
xnor U17710 (N_17710,N_17341,N_17470);
or U17711 (N_17711,N_17311,N_17161);
nor U17712 (N_17712,N_17221,N_17366);
or U17713 (N_17713,N_17106,N_16594);
and U17714 (N_17714,N_17006,N_17142);
or U17715 (N_17715,N_17173,N_17315);
nor U17716 (N_17716,N_16730,N_17258);
xor U17717 (N_17717,N_16328,N_16421);
nand U17718 (N_17718,N_16563,N_16812);
nand U17719 (N_17719,N_16709,N_17375);
and U17720 (N_17720,N_16442,N_16733);
nand U17721 (N_17721,N_17306,N_17222);
and U17722 (N_17722,N_16618,N_16911);
and U17723 (N_17723,N_17074,N_17149);
nor U17724 (N_17724,N_16759,N_17089);
and U17725 (N_17725,N_16486,N_16256);
and U17726 (N_17726,N_17011,N_17433);
and U17727 (N_17727,N_17485,N_17096);
xor U17728 (N_17728,N_17423,N_16612);
and U17729 (N_17729,N_17099,N_16304);
nor U17730 (N_17730,N_16894,N_16764);
and U17731 (N_17731,N_16693,N_16620);
and U17732 (N_17732,N_17318,N_16930);
xor U17733 (N_17733,N_17406,N_16264);
nor U17734 (N_17734,N_16326,N_16674);
nor U17735 (N_17735,N_16943,N_17103);
nand U17736 (N_17736,N_17220,N_16354);
or U17737 (N_17737,N_16912,N_16916);
nor U17738 (N_17738,N_16393,N_16379);
nor U17739 (N_17739,N_17114,N_17084);
and U17740 (N_17740,N_17413,N_17184);
xnor U17741 (N_17741,N_16487,N_16284);
nor U17742 (N_17742,N_16937,N_16287);
xnor U17743 (N_17743,N_16863,N_16948);
xnor U17744 (N_17744,N_16396,N_16504);
or U17745 (N_17745,N_17365,N_16477);
or U17746 (N_17746,N_17051,N_16472);
nor U17747 (N_17747,N_16311,N_17180);
xnor U17748 (N_17748,N_16514,N_17126);
and U17749 (N_17749,N_17421,N_16975);
or U17750 (N_17750,N_17046,N_16962);
xnor U17751 (N_17751,N_16312,N_17213);
xor U17752 (N_17752,N_17448,N_16732);
xnor U17753 (N_17753,N_17237,N_17317);
xnor U17754 (N_17754,N_17196,N_16969);
xor U17755 (N_17755,N_16485,N_16941);
and U17756 (N_17756,N_16285,N_17094);
nor U17757 (N_17757,N_17309,N_17368);
nand U17758 (N_17758,N_17234,N_17342);
or U17759 (N_17759,N_16570,N_16303);
xnor U17760 (N_17760,N_16772,N_17045);
xnor U17761 (N_17761,N_16444,N_17233);
xnor U17762 (N_17762,N_17357,N_17463);
or U17763 (N_17763,N_16697,N_16505);
and U17764 (N_17764,N_16506,N_16954);
and U17765 (N_17765,N_16404,N_16720);
nor U17766 (N_17766,N_16986,N_16981);
and U17767 (N_17767,N_17294,N_17052);
nand U17768 (N_17768,N_17361,N_16336);
nor U17769 (N_17769,N_16329,N_16592);
xor U17770 (N_17770,N_16858,N_16555);
or U17771 (N_17771,N_17354,N_16651);
and U17772 (N_17772,N_17295,N_17034);
xor U17773 (N_17773,N_16518,N_17270);
nor U17774 (N_17774,N_16744,N_17217);
and U17775 (N_17775,N_17111,N_16647);
nand U17776 (N_17776,N_16458,N_16655);
nand U17777 (N_17777,N_16959,N_16645);
or U17778 (N_17778,N_16757,N_17154);
nor U17779 (N_17779,N_16874,N_17266);
xnor U17780 (N_17780,N_16782,N_16367);
and U17781 (N_17781,N_17169,N_16359);
xor U17782 (N_17782,N_17031,N_16315);
or U17783 (N_17783,N_17439,N_17092);
nand U17784 (N_17784,N_17008,N_17490);
or U17785 (N_17785,N_17460,N_16755);
xnor U17786 (N_17786,N_16414,N_16640);
or U17787 (N_17787,N_16741,N_17300);
nand U17788 (N_17788,N_16552,N_17019);
nand U17789 (N_17789,N_17082,N_16673);
and U17790 (N_17790,N_16323,N_16544);
or U17791 (N_17791,N_17466,N_17459);
xnor U17792 (N_17792,N_17087,N_16703);
and U17793 (N_17793,N_17189,N_17025);
xnor U17794 (N_17794,N_17028,N_16957);
xor U17795 (N_17795,N_17434,N_16519);
xor U17796 (N_17796,N_17163,N_16881);
and U17797 (N_17797,N_17054,N_17202);
xor U17798 (N_17798,N_17133,N_16891);
nor U17799 (N_17799,N_16569,N_17397);
nor U17800 (N_17800,N_17132,N_16351);
or U17801 (N_17801,N_16777,N_17411);
xnor U17802 (N_17802,N_16683,N_16745);
xor U17803 (N_17803,N_17067,N_16512);
and U17804 (N_17804,N_17369,N_16489);
nor U17805 (N_17805,N_16617,N_16447);
xnor U17806 (N_17806,N_16926,N_16749);
nand U17807 (N_17807,N_17481,N_16274);
or U17808 (N_17808,N_16293,N_17377);
nand U17809 (N_17809,N_16992,N_16595);
xnor U17810 (N_17810,N_16794,N_17064);
nand U17811 (N_17811,N_16428,N_17388);
and U17812 (N_17812,N_17148,N_16900);
or U17813 (N_17813,N_16377,N_16670);
nor U17814 (N_17814,N_17281,N_17321);
and U17815 (N_17815,N_16340,N_17358);
xor U17816 (N_17816,N_16919,N_16374);
or U17817 (N_17817,N_17480,N_17327);
or U17818 (N_17818,N_16802,N_16448);
or U17819 (N_17819,N_17312,N_16441);
nand U17820 (N_17820,N_17418,N_16842);
or U17821 (N_17821,N_16615,N_16991);
or U17822 (N_17822,N_17303,N_16823);
nand U17823 (N_17823,N_16950,N_16510);
xor U17824 (N_17824,N_17260,N_17215);
or U17825 (N_17825,N_16822,N_17495);
nand U17826 (N_17826,N_16985,N_17322);
and U17827 (N_17827,N_16590,N_16797);
or U17828 (N_17828,N_16905,N_17347);
and U17829 (N_17829,N_16597,N_16614);
nand U17830 (N_17830,N_16371,N_17276);
nor U17831 (N_17831,N_16613,N_16536);
nor U17832 (N_17832,N_16394,N_16933);
and U17833 (N_17833,N_16257,N_17235);
xnor U17834 (N_17834,N_16619,N_17265);
nand U17835 (N_17835,N_16956,N_17272);
nor U17836 (N_17836,N_17137,N_16862);
and U17837 (N_17837,N_16624,N_16416);
xnor U17838 (N_17838,N_16679,N_17038);
nand U17839 (N_17839,N_16400,N_17095);
or U17840 (N_17840,N_16497,N_17461);
or U17841 (N_17841,N_16792,N_17335);
or U17842 (N_17842,N_16751,N_16292);
nand U17843 (N_17843,N_16835,N_16378);
xor U17844 (N_17844,N_16530,N_16362);
nand U17845 (N_17845,N_16845,N_17373);
and U17846 (N_17846,N_17284,N_16357);
or U17847 (N_17847,N_16468,N_16773);
nor U17848 (N_17848,N_16339,N_16830);
xnor U17849 (N_17849,N_16847,N_17002);
nor U17850 (N_17850,N_17159,N_17473);
nor U17851 (N_17851,N_17299,N_16808);
nor U17852 (N_17852,N_17336,N_16302);
nor U17853 (N_17853,N_16580,N_17232);
or U17854 (N_17854,N_17120,N_16380);
nor U17855 (N_17855,N_17043,N_17345);
or U17856 (N_17856,N_16869,N_16471);
xor U17857 (N_17857,N_17097,N_16947);
nand U17858 (N_17858,N_16560,N_16427);
nand U17859 (N_17859,N_16499,N_16735);
and U17860 (N_17860,N_17015,N_17201);
nand U17861 (N_17861,N_16250,N_16283);
xnor U17862 (N_17862,N_16966,N_16671);
and U17863 (N_17863,N_16521,N_16432);
or U17864 (N_17864,N_17231,N_16914);
xor U17865 (N_17865,N_16479,N_17412);
nand U17866 (N_17866,N_16908,N_17241);
xor U17867 (N_17867,N_16533,N_17285);
xnor U17868 (N_17868,N_16988,N_16649);
and U17869 (N_17869,N_16298,N_17376);
xnor U17870 (N_17870,N_17248,N_16884);
nand U17871 (N_17871,N_17399,N_17216);
nor U17872 (N_17872,N_16306,N_16875);
and U17873 (N_17873,N_16467,N_16711);
and U17874 (N_17874,N_17224,N_17247);
nor U17875 (N_17875,N_16628,N_17209);
or U17876 (N_17876,N_16892,N_16718);
and U17877 (N_17877,N_16488,N_16437);
and U17878 (N_17878,N_17499,N_16789);
xnor U17879 (N_17879,N_16942,N_16989);
or U17880 (N_17880,N_17183,N_16294);
nand U17881 (N_17881,N_16462,N_16433);
nand U17882 (N_17882,N_17475,N_17102);
nor U17883 (N_17883,N_16843,N_17326);
nor U17884 (N_17884,N_16524,N_16967);
nand U17885 (N_17885,N_16704,N_17333);
nand U17886 (N_17886,N_16338,N_16729);
and U17887 (N_17887,N_16550,N_16253);
xnor U17888 (N_17888,N_17212,N_17127);
xnor U17889 (N_17889,N_17282,N_17121);
nand U17890 (N_17890,N_17292,N_16369);
xnor U17891 (N_17891,N_17199,N_16278);
and U17892 (N_17892,N_16725,N_17113);
and U17893 (N_17893,N_16652,N_16426);
nand U17894 (N_17894,N_16660,N_16252);
nor U17895 (N_17895,N_16602,N_16762);
nor U17896 (N_17896,N_16571,N_16774);
nand U17897 (N_17897,N_17016,N_17274);
or U17898 (N_17898,N_17160,N_16861);
nor U17899 (N_17899,N_17350,N_17449);
or U17900 (N_17900,N_16599,N_17371);
xnor U17901 (N_17901,N_16849,N_17190);
nor U17902 (N_17902,N_17359,N_16262);
and U17903 (N_17903,N_17471,N_16882);
or U17904 (N_17904,N_16452,N_17166);
and U17905 (N_17905,N_16758,N_17178);
nand U17906 (N_17906,N_17426,N_17454);
or U17907 (N_17907,N_16577,N_16734);
nand U17908 (N_17908,N_17020,N_16330);
xor U17909 (N_17909,N_16983,N_16678);
or U17910 (N_17910,N_16927,N_17355);
xor U17911 (N_17911,N_16616,N_17151);
or U17912 (N_17912,N_17462,N_16324);
or U17913 (N_17913,N_16295,N_16996);
xor U17914 (N_17914,N_17181,N_17134);
nor U17915 (N_17915,N_16586,N_16800);
or U17916 (N_17916,N_17174,N_16507);
and U17917 (N_17917,N_17205,N_17337);
or U17918 (N_17918,N_16716,N_17387);
and U17919 (N_17919,N_16277,N_17344);
nor U17920 (N_17920,N_16799,N_16576);
and U17921 (N_17921,N_16502,N_16403);
nand U17922 (N_17922,N_16407,N_17069);
nor U17923 (N_17923,N_16923,N_16903);
or U17924 (N_17924,N_16982,N_16401);
nand U17925 (N_17925,N_16686,N_16778);
xnor U17926 (N_17926,N_16508,N_17310);
nor U17927 (N_17927,N_17343,N_17384);
or U17928 (N_17928,N_17245,N_17496);
or U17929 (N_17929,N_17367,N_17389);
nand U17930 (N_17930,N_17039,N_16727);
nor U17931 (N_17931,N_17268,N_16482);
xor U17932 (N_17932,N_16368,N_16829);
nand U17933 (N_17933,N_16770,N_16752);
or U17934 (N_17934,N_16910,N_16793);
nand U17935 (N_17935,N_17026,N_17236);
xor U17936 (N_17936,N_16543,N_16319);
xnor U17937 (N_17937,N_17147,N_16984);
nand U17938 (N_17938,N_16434,N_17230);
nor U17939 (N_17939,N_16654,N_17197);
or U17940 (N_17940,N_16288,N_16254);
or U17941 (N_17941,N_17177,N_16373);
nand U17942 (N_17942,N_17207,N_16696);
nand U17943 (N_17943,N_16695,N_16258);
nand U17944 (N_17944,N_16322,N_17193);
nand U17945 (N_17945,N_16445,N_16915);
nand U17946 (N_17946,N_17122,N_17104);
nand U17947 (N_17947,N_17464,N_17275);
nand U17948 (N_17948,N_17479,N_16251);
nand U17949 (N_17949,N_16868,N_17145);
or U17950 (N_17950,N_17150,N_17416);
nand U17951 (N_17951,N_16997,N_16921);
nor U17952 (N_17952,N_16435,N_17010);
xnor U17953 (N_17953,N_16466,N_17498);
and U17954 (N_17954,N_16721,N_17198);
nand U17955 (N_17955,N_17297,N_17396);
or U17956 (N_17956,N_16980,N_16961);
and U17957 (N_17957,N_16687,N_16767);
nand U17958 (N_17958,N_17110,N_16705);
or U17959 (N_17959,N_16481,N_17324);
or U17960 (N_17960,N_16974,N_16281);
xor U17961 (N_17961,N_16484,N_16999);
nand U17962 (N_17962,N_16455,N_17465);
nand U17963 (N_17963,N_17125,N_17320);
nor U17964 (N_17964,N_16726,N_16513);
and U17965 (N_17965,N_17252,N_16813);
nand U17966 (N_17966,N_16305,N_16775);
and U17967 (N_17967,N_16578,N_17246);
nor U17968 (N_17968,N_17332,N_17393);
xnor U17969 (N_17969,N_17286,N_16604);
nor U17970 (N_17970,N_16406,N_16430);
xor U17971 (N_17971,N_17447,N_17139);
or U17972 (N_17972,N_16376,N_17185);
or U17973 (N_17973,N_16766,N_16546);
xnor U17974 (N_17974,N_16637,N_16945);
nand U17975 (N_17975,N_17049,N_17438);
or U17976 (N_17976,N_16364,N_16297);
and U17977 (N_17977,N_16439,N_16781);
nor U17978 (N_17978,N_16450,N_16390);
nand U17979 (N_17979,N_17130,N_17436);
and U17980 (N_17980,N_16370,N_16700);
nor U17981 (N_17981,N_16840,N_17085);
or U17982 (N_17982,N_16331,N_16496);
nor U17983 (N_17983,N_16639,N_17033);
or U17984 (N_17984,N_16724,N_17063);
or U17985 (N_17985,N_16384,N_16389);
nand U17986 (N_17986,N_17362,N_16658);
nor U17987 (N_17987,N_17353,N_16898);
xnor U17988 (N_17988,N_17328,N_17432);
xnor U17989 (N_17989,N_17170,N_16572);
nor U17990 (N_17990,N_17477,N_16771);
nor U17991 (N_17991,N_16656,N_17003);
or U17992 (N_17992,N_16273,N_17075);
nor U17993 (N_17993,N_16747,N_16851);
and U17994 (N_17994,N_16738,N_17340);
nand U17995 (N_17995,N_16848,N_17044);
and U17996 (N_17996,N_16841,N_17256);
nand U17997 (N_17997,N_17360,N_16994);
nand U17998 (N_17998,N_17467,N_17055);
nand U17999 (N_17999,N_16446,N_17325);
xnor U18000 (N_18000,N_17062,N_17307);
xnor U18001 (N_18001,N_17182,N_16856);
nand U18002 (N_18002,N_16831,N_16263);
xnor U18003 (N_18003,N_17000,N_16623);
nor U18004 (N_18004,N_16801,N_17331);
xnor U18005 (N_18005,N_16866,N_16935);
or U18006 (N_18006,N_16970,N_16952);
and U18007 (N_18007,N_16575,N_16634);
and U18008 (N_18008,N_16535,N_17363);
xor U18009 (N_18009,N_16743,N_16345);
or U18010 (N_18010,N_17158,N_16318);
xor U18011 (N_18011,N_17057,N_16531);
and U18012 (N_18012,N_17072,N_16865);
or U18013 (N_18013,N_16712,N_16314);
nand U18014 (N_18014,N_16827,N_16805);
and U18015 (N_18015,N_17379,N_17136);
nor U18016 (N_18016,N_16551,N_16765);
and U18017 (N_18017,N_16429,N_17179);
nand U18018 (N_18018,N_16493,N_17302);
nor U18019 (N_18019,N_16261,N_16824);
and U18020 (N_18020,N_16990,N_17314);
nor U18021 (N_18021,N_16895,N_16932);
or U18022 (N_18022,N_16382,N_17422);
nor U18023 (N_18023,N_16372,N_16754);
nand U18024 (N_18024,N_16978,N_16833);
and U18025 (N_18025,N_17364,N_17061);
or U18026 (N_18026,N_16541,N_17036);
and U18027 (N_18027,N_16269,N_16788);
or U18028 (N_18028,N_16779,N_16538);
nand U18029 (N_18029,N_17279,N_16636);
nand U18030 (N_18030,N_16279,N_16667);
nor U18031 (N_18031,N_17450,N_16549);
or U18032 (N_18032,N_16410,N_16828);
and U18033 (N_18033,N_17140,N_17210);
nor U18034 (N_18034,N_16902,N_16922);
nand U18035 (N_18035,N_16938,N_16495);
nor U18036 (N_18036,N_16413,N_16332);
xnor U18037 (N_18037,N_17417,N_16885);
xnor U18038 (N_18038,N_16388,N_16852);
or U18039 (N_18039,N_16870,N_17349);
or U18040 (N_18040,N_17267,N_17255);
or U18041 (N_18041,N_16684,N_16672);
nor U18042 (N_18042,N_17308,N_17081);
and U18043 (N_18043,N_17157,N_16527);
or U18044 (N_18044,N_17403,N_17004);
nand U18045 (N_18045,N_16855,N_16838);
or U18046 (N_18046,N_16836,N_16456);
nor U18047 (N_18047,N_16804,N_16291);
nor U18048 (N_18048,N_17007,N_17264);
nand U18049 (N_18049,N_17404,N_16500);
and U18050 (N_18050,N_17100,N_17402);
or U18051 (N_18051,N_16349,N_16692);
or U18052 (N_18052,N_17386,N_17428);
xor U18053 (N_18053,N_16680,N_16361);
and U18054 (N_18054,N_16316,N_17453);
xnor U18055 (N_18055,N_16457,N_16936);
and U18056 (N_18056,N_16526,N_16363);
nand U18057 (N_18057,N_16791,N_17445);
or U18058 (N_18058,N_16386,N_17029);
xnor U18059 (N_18059,N_16562,N_16806);
nand U18060 (N_18060,N_16409,N_16475);
and U18061 (N_18061,N_16375,N_16963);
or U18062 (N_18062,N_17291,N_16960);
or U18063 (N_18063,N_17053,N_16666);
xnor U18064 (N_18064,N_16810,N_16630);
xnor U18065 (N_18065,N_16815,N_16701);
nor U18066 (N_18066,N_17108,N_16625);
or U18067 (N_18067,N_16600,N_17316);
and U18068 (N_18068,N_16392,N_17024);
xor U18069 (N_18069,N_16642,N_16461);
or U18070 (N_18070,N_17112,N_16542);
nor U18071 (N_18071,N_16491,N_16564);
nor U18072 (N_18072,N_17491,N_16348);
xnor U18073 (N_18073,N_16689,N_17021);
nand U18074 (N_18074,N_17419,N_17091);
nor U18075 (N_18075,N_17305,N_17192);
xor U18076 (N_18076,N_16593,N_17141);
or U18077 (N_18077,N_16494,N_16955);
or U18078 (N_18078,N_17330,N_16907);
xnor U18079 (N_18079,N_17167,N_16906);
nor U18080 (N_18080,N_16924,N_17203);
nand U18081 (N_18081,N_17301,N_17409);
xnor U18082 (N_18082,N_17143,N_17164);
or U18083 (N_18083,N_17420,N_17304);
nor U18084 (N_18084,N_16896,N_16387);
or U18085 (N_18085,N_16566,N_16307);
xor U18086 (N_18086,N_16431,N_17395);
and U18087 (N_18087,N_16879,N_17115);
or U18088 (N_18088,N_16694,N_17101);
or U18089 (N_18089,N_16454,N_16899);
and U18090 (N_18090,N_16659,N_17468);
nand U18091 (N_18091,N_17329,N_16490);
nand U18092 (N_18092,N_16522,N_16691);
xor U18093 (N_18093,N_17195,N_16282);
nor U18094 (N_18094,N_17014,N_17223);
or U18095 (N_18095,N_16469,N_17218);
nor U18096 (N_18096,N_16420,N_16350);
and U18097 (N_18097,N_17346,N_16525);
and U18098 (N_18098,N_17056,N_16605);
nor U18099 (N_18099,N_16301,N_16587);
nor U18100 (N_18100,N_16973,N_16668);
or U18101 (N_18101,N_16622,N_16877);
nand U18102 (N_18102,N_16296,N_17287);
and U18103 (N_18103,N_16290,N_17042);
xnor U18104 (N_18104,N_16934,N_16706);
nor U18105 (N_18105,N_17175,N_17271);
nand U18106 (N_18106,N_17080,N_17482);
nor U18107 (N_18107,N_16731,N_16688);
and U18108 (N_18108,N_16464,N_17165);
or U18109 (N_18109,N_16473,N_16365);
nand U18110 (N_18110,N_17050,N_16676);
xnor U18111 (N_18111,N_16682,N_17251);
nor U18112 (N_18112,N_17474,N_17070);
xor U18113 (N_18113,N_17427,N_17009);
nand U18114 (N_18114,N_16344,N_16443);
and U18115 (N_18115,N_17408,N_16275);
xnor U18116 (N_18116,N_16270,N_16753);
and U18117 (N_18117,N_17249,N_16589);
nand U18118 (N_18118,N_16780,N_16501);
nor U18119 (N_18119,N_17109,N_16480);
and U18120 (N_18120,N_16760,N_16460);
nand U18121 (N_18121,N_17269,N_16719);
nand U18122 (N_18122,N_17058,N_16327);
xor U18123 (N_18123,N_17116,N_17446);
or U18124 (N_18124,N_16976,N_17135);
xor U18125 (N_18125,N_17282,N_17302);
xor U18126 (N_18126,N_16682,N_17350);
or U18127 (N_18127,N_16681,N_17298);
xor U18128 (N_18128,N_16306,N_16937);
xor U18129 (N_18129,N_16904,N_16828);
xnor U18130 (N_18130,N_16971,N_16600);
xor U18131 (N_18131,N_16687,N_16519);
xnor U18132 (N_18132,N_16771,N_17174);
and U18133 (N_18133,N_17291,N_17416);
xnor U18134 (N_18134,N_16415,N_16803);
xnor U18135 (N_18135,N_16524,N_17143);
nor U18136 (N_18136,N_16505,N_17041);
nand U18137 (N_18137,N_16492,N_16600);
and U18138 (N_18138,N_16847,N_16501);
or U18139 (N_18139,N_16700,N_16374);
nor U18140 (N_18140,N_16704,N_17123);
xor U18141 (N_18141,N_16853,N_17443);
nand U18142 (N_18142,N_17253,N_16836);
nor U18143 (N_18143,N_16522,N_16312);
nand U18144 (N_18144,N_17101,N_16290);
nand U18145 (N_18145,N_17405,N_16844);
nand U18146 (N_18146,N_17076,N_16251);
or U18147 (N_18147,N_16389,N_17474);
or U18148 (N_18148,N_16842,N_17298);
or U18149 (N_18149,N_17061,N_16640);
nor U18150 (N_18150,N_16316,N_17489);
xor U18151 (N_18151,N_16615,N_17181);
nor U18152 (N_18152,N_16477,N_16575);
nor U18153 (N_18153,N_17491,N_16501);
nor U18154 (N_18154,N_16905,N_16968);
xnor U18155 (N_18155,N_17476,N_16370);
nor U18156 (N_18156,N_16675,N_16946);
xor U18157 (N_18157,N_16979,N_17442);
nand U18158 (N_18158,N_16717,N_16833);
and U18159 (N_18159,N_16360,N_16675);
and U18160 (N_18160,N_17329,N_16373);
or U18161 (N_18161,N_16349,N_16778);
nor U18162 (N_18162,N_16298,N_17257);
or U18163 (N_18163,N_17311,N_16876);
nand U18164 (N_18164,N_16302,N_17370);
and U18165 (N_18165,N_17034,N_17074);
nor U18166 (N_18166,N_16252,N_16656);
and U18167 (N_18167,N_16442,N_16251);
nand U18168 (N_18168,N_16707,N_16877);
or U18169 (N_18169,N_17398,N_17323);
nor U18170 (N_18170,N_17243,N_16983);
nand U18171 (N_18171,N_17438,N_16921);
nand U18172 (N_18172,N_16404,N_17229);
nor U18173 (N_18173,N_16312,N_16859);
and U18174 (N_18174,N_17022,N_17192);
and U18175 (N_18175,N_17287,N_16284);
and U18176 (N_18176,N_17087,N_17069);
and U18177 (N_18177,N_16358,N_16931);
or U18178 (N_18178,N_16718,N_17199);
or U18179 (N_18179,N_17132,N_16292);
and U18180 (N_18180,N_17408,N_17134);
or U18181 (N_18181,N_16986,N_16669);
xnor U18182 (N_18182,N_16553,N_16801);
or U18183 (N_18183,N_16579,N_16573);
and U18184 (N_18184,N_17210,N_16735);
xnor U18185 (N_18185,N_17402,N_16619);
nor U18186 (N_18186,N_16408,N_16326);
nand U18187 (N_18187,N_16397,N_17346);
nor U18188 (N_18188,N_16799,N_16512);
or U18189 (N_18189,N_16965,N_16919);
nor U18190 (N_18190,N_16932,N_17069);
or U18191 (N_18191,N_17387,N_16579);
xor U18192 (N_18192,N_17376,N_17461);
nand U18193 (N_18193,N_17251,N_16656);
xor U18194 (N_18194,N_17334,N_16866);
and U18195 (N_18195,N_16622,N_17252);
and U18196 (N_18196,N_16335,N_16577);
nor U18197 (N_18197,N_17469,N_16749);
nand U18198 (N_18198,N_16536,N_16889);
nand U18199 (N_18199,N_16466,N_16305);
xnor U18200 (N_18200,N_16492,N_17345);
and U18201 (N_18201,N_16450,N_16265);
nor U18202 (N_18202,N_17485,N_17208);
xor U18203 (N_18203,N_16422,N_16809);
xor U18204 (N_18204,N_16386,N_17397);
xnor U18205 (N_18205,N_16617,N_16339);
or U18206 (N_18206,N_16300,N_16559);
nand U18207 (N_18207,N_16321,N_17348);
and U18208 (N_18208,N_16531,N_16837);
nor U18209 (N_18209,N_16274,N_17100);
or U18210 (N_18210,N_17317,N_16644);
and U18211 (N_18211,N_17243,N_16991);
nand U18212 (N_18212,N_17322,N_16717);
and U18213 (N_18213,N_17025,N_16756);
nand U18214 (N_18214,N_16635,N_16926);
and U18215 (N_18215,N_17409,N_16803);
xor U18216 (N_18216,N_17438,N_16624);
nand U18217 (N_18217,N_16583,N_16340);
nor U18218 (N_18218,N_17005,N_16343);
or U18219 (N_18219,N_17157,N_17273);
xnor U18220 (N_18220,N_17463,N_16794);
and U18221 (N_18221,N_16669,N_17497);
xnor U18222 (N_18222,N_16448,N_17068);
nand U18223 (N_18223,N_16438,N_16734);
and U18224 (N_18224,N_17493,N_16756);
nor U18225 (N_18225,N_16538,N_16294);
nor U18226 (N_18226,N_17180,N_16716);
or U18227 (N_18227,N_17116,N_17338);
or U18228 (N_18228,N_17068,N_16921);
nor U18229 (N_18229,N_17310,N_17175);
nand U18230 (N_18230,N_16959,N_17277);
and U18231 (N_18231,N_17074,N_17413);
xor U18232 (N_18232,N_17323,N_16503);
nor U18233 (N_18233,N_16612,N_16843);
or U18234 (N_18234,N_16686,N_16717);
xnor U18235 (N_18235,N_16361,N_17261);
and U18236 (N_18236,N_17084,N_17258);
or U18237 (N_18237,N_16703,N_17347);
nand U18238 (N_18238,N_17295,N_16938);
and U18239 (N_18239,N_16792,N_16882);
nand U18240 (N_18240,N_16800,N_16655);
nand U18241 (N_18241,N_17410,N_16451);
nand U18242 (N_18242,N_17107,N_16528);
xnor U18243 (N_18243,N_17178,N_16727);
or U18244 (N_18244,N_16635,N_16954);
nand U18245 (N_18245,N_16380,N_16838);
nand U18246 (N_18246,N_17212,N_16722);
or U18247 (N_18247,N_17157,N_16682);
nand U18248 (N_18248,N_17211,N_17429);
and U18249 (N_18249,N_17172,N_17459);
nand U18250 (N_18250,N_17307,N_16408);
nor U18251 (N_18251,N_16563,N_17295);
or U18252 (N_18252,N_17345,N_16512);
nor U18253 (N_18253,N_17125,N_16362);
xor U18254 (N_18254,N_16900,N_17023);
and U18255 (N_18255,N_17141,N_17112);
xor U18256 (N_18256,N_17302,N_16414);
nand U18257 (N_18257,N_16784,N_16701);
nor U18258 (N_18258,N_16298,N_16335);
xor U18259 (N_18259,N_17236,N_17105);
and U18260 (N_18260,N_16993,N_17033);
nand U18261 (N_18261,N_17250,N_17056);
xnor U18262 (N_18262,N_16274,N_17430);
nand U18263 (N_18263,N_17259,N_17158);
nand U18264 (N_18264,N_17058,N_17014);
or U18265 (N_18265,N_16780,N_16554);
xor U18266 (N_18266,N_16298,N_16591);
xnor U18267 (N_18267,N_17344,N_16265);
nor U18268 (N_18268,N_16295,N_16697);
nor U18269 (N_18269,N_16395,N_17161);
nand U18270 (N_18270,N_16481,N_17266);
xnor U18271 (N_18271,N_16452,N_17090);
or U18272 (N_18272,N_16441,N_16868);
xor U18273 (N_18273,N_17092,N_17355);
nor U18274 (N_18274,N_16653,N_16806);
nor U18275 (N_18275,N_16519,N_16965);
nor U18276 (N_18276,N_16810,N_16628);
xor U18277 (N_18277,N_16270,N_16566);
xor U18278 (N_18278,N_17074,N_17371);
nor U18279 (N_18279,N_16592,N_16927);
or U18280 (N_18280,N_16387,N_16371);
or U18281 (N_18281,N_16994,N_16534);
xnor U18282 (N_18282,N_16999,N_16523);
nor U18283 (N_18283,N_17074,N_17405);
and U18284 (N_18284,N_16606,N_17464);
nor U18285 (N_18285,N_16708,N_16510);
nor U18286 (N_18286,N_16811,N_16590);
or U18287 (N_18287,N_16786,N_16869);
or U18288 (N_18288,N_16650,N_17253);
or U18289 (N_18289,N_17318,N_17341);
xnor U18290 (N_18290,N_16323,N_16801);
xor U18291 (N_18291,N_16711,N_16682);
nor U18292 (N_18292,N_17344,N_16773);
or U18293 (N_18293,N_17403,N_16629);
and U18294 (N_18294,N_16631,N_17016);
nand U18295 (N_18295,N_17297,N_16611);
xnor U18296 (N_18296,N_16817,N_16809);
xnor U18297 (N_18297,N_17324,N_17459);
or U18298 (N_18298,N_17402,N_16769);
xnor U18299 (N_18299,N_16580,N_17259);
xor U18300 (N_18300,N_16406,N_16397);
nand U18301 (N_18301,N_16663,N_16476);
and U18302 (N_18302,N_17154,N_16924);
or U18303 (N_18303,N_16746,N_16307);
and U18304 (N_18304,N_16318,N_17078);
xnor U18305 (N_18305,N_17157,N_16747);
nand U18306 (N_18306,N_16982,N_17290);
and U18307 (N_18307,N_16476,N_16296);
and U18308 (N_18308,N_16466,N_17376);
and U18309 (N_18309,N_17455,N_17167);
and U18310 (N_18310,N_16544,N_16701);
xnor U18311 (N_18311,N_17123,N_17340);
or U18312 (N_18312,N_17069,N_17393);
nand U18313 (N_18313,N_16806,N_16472);
or U18314 (N_18314,N_17153,N_16610);
nand U18315 (N_18315,N_16678,N_17320);
nand U18316 (N_18316,N_16532,N_16631);
and U18317 (N_18317,N_16366,N_17205);
xor U18318 (N_18318,N_17330,N_16704);
or U18319 (N_18319,N_16893,N_16309);
or U18320 (N_18320,N_16969,N_16647);
nor U18321 (N_18321,N_16693,N_16344);
xnor U18322 (N_18322,N_16255,N_17397);
xnor U18323 (N_18323,N_17052,N_16592);
nor U18324 (N_18324,N_16737,N_16741);
nor U18325 (N_18325,N_16777,N_17187);
xnor U18326 (N_18326,N_17412,N_16810);
and U18327 (N_18327,N_16539,N_17050);
and U18328 (N_18328,N_16490,N_17414);
and U18329 (N_18329,N_16522,N_17200);
and U18330 (N_18330,N_17323,N_16747);
or U18331 (N_18331,N_16578,N_16559);
nand U18332 (N_18332,N_17494,N_17171);
or U18333 (N_18333,N_17266,N_17042);
nor U18334 (N_18334,N_16674,N_17439);
and U18335 (N_18335,N_16921,N_16485);
and U18336 (N_18336,N_16484,N_16963);
xnor U18337 (N_18337,N_17401,N_16615);
nand U18338 (N_18338,N_16284,N_16358);
nand U18339 (N_18339,N_16381,N_16635);
nor U18340 (N_18340,N_17156,N_17398);
nand U18341 (N_18341,N_16335,N_16800);
and U18342 (N_18342,N_17406,N_17439);
nand U18343 (N_18343,N_16380,N_16561);
or U18344 (N_18344,N_16388,N_17036);
xnor U18345 (N_18345,N_16322,N_16998);
xor U18346 (N_18346,N_17153,N_16612);
nor U18347 (N_18347,N_16760,N_17148);
nand U18348 (N_18348,N_16862,N_17191);
nor U18349 (N_18349,N_17194,N_16509);
and U18350 (N_18350,N_16909,N_16903);
xor U18351 (N_18351,N_16254,N_16733);
or U18352 (N_18352,N_16827,N_16803);
nor U18353 (N_18353,N_16933,N_16646);
and U18354 (N_18354,N_17167,N_17081);
nand U18355 (N_18355,N_17022,N_16673);
or U18356 (N_18356,N_17472,N_16641);
or U18357 (N_18357,N_17385,N_16601);
nand U18358 (N_18358,N_17158,N_16516);
or U18359 (N_18359,N_16704,N_17226);
nor U18360 (N_18360,N_17372,N_16813);
and U18361 (N_18361,N_17108,N_16968);
xor U18362 (N_18362,N_17173,N_16856);
and U18363 (N_18363,N_16457,N_16531);
and U18364 (N_18364,N_16652,N_16717);
nor U18365 (N_18365,N_16703,N_17301);
xor U18366 (N_18366,N_16933,N_16431);
nand U18367 (N_18367,N_17410,N_16433);
nand U18368 (N_18368,N_17227,N_16733);
xnor U18369 (N_18369,N_16782,N_16252);
nand U18370 (N_18370,N_16777,N_17257);
and U18371 (N_18371,N_16401,N_16860);
nor U18372 (N_18372,N_17109,N_17296);
or U18373 (N_18373,N_16859,N_17486);
xnor U18374 (N_18374,N_16747,N_16813);
or U18375 (N_18375,N_17368,N_17011);
and U18376 (N_18376,N_16953,N_17102);
nor U18377 (N_18377,N_16887,N_16337);
xnor U18378 (N_18378,N_16761,N_17441);
or U18379 (N_18379,N_17307,N_16823);
nand U18380 (N_18380,N_16368,N_16672);
or U18381 (N_18381,N_17180,N_16401);
nand U18382 (N_18382,N_17095,N_17352);
and U18383 (N_18383,N_16564,N_17336);
or U18384 (N_18384,N_17349,N_16693);
xnor U18385 (N_18385,N_16987,N_16723);
or U18386 (N_18386,N_17184,N_16521);
or U18387 (N_18387,N_16541,N_16413);
or U18388 (N_18388,N_17248,N_17251);
nor U18389 (N_18389,N_16464,N_16528);
nand U18390 (N_18390,N_17418,N_16536);
nand U18391 (N_18391,N_17349,N_16581);
nand U18392 (N_18392,N_16491,N_17377);
nand U18393 (N_18393,N_16387,N_17326);
and U18394 (N_18394,N_17356,N_16406);
and U18395 (N_18395,N_16970,N_16323);
xor U18396 (N_18396,N_17497,N_17083);
or U18397 (N_18397,N_16906,N_17125);
nor U18398 (N_18398,N_17479,N_16629);
nor U18399 (N_18399,N_17333,N_17000);
and U18400 (N_18400,N_16333,N_17306);
nor U18401 (N_18401,N_16304,N_17145);
xnor U18402 (N_18402,N_17333,N_16282);
nand U18403 (N_18403,N_16959,N_16969);
nor U18404 (N_18404,N_17188,N_16402);
nand U18405 (N_18405,N_17366,N_16523);
nand U18406 (N_18406,N_17296,N_17006);
xor U18407 (N_18407,N_16833,N_16461);
or U18408 (N_18408,N_17463,N_16398);
xor U18409 (N_18409,N_16288,N_17143);
nor U18410 (N_18410,N_16686,N_16750);
and U18411 (N_18411,N_17081,N_16505);
xor U18412 (N_18412,N_16549,N_17400);
xor U18413 (N_18413,N_16653,N_16336);
and U18414 (N_18414,N_17375,N_17155);
and U18415 (N_18415,N_16414,N_16872);
and U18416 (N_18416,N_16997,N_16961);
nor U18417 (N_18417,N_17230,N_16607);
nand U18418 (N_18418,N_16559,N_16680);
xor U18419 (N_18419,N_16347,N_16565);
xor U18420 (N_18420,N_17139,N_17401);
xor U18421 (N_18421,N_17008,N_16879);
xor U18422 (N_18422,N_16562,N_17056);
or U18423 (N_18423,N_17259,N_16852);
or U18424 (N_18424,N_16633,N_17090);
and U18425 (N_18425,N_17460,N_16779);
nor U18426 (N_18426,N_16796,N_16445);
nand U18427 (N_18427,N_16692,N_16924);
and U18428 (N_18428,N_16539,N_17258);
nand U18429 (N_18429,N_17355,N_16510);
xor U18430 (N_18430,N_17352,N_16366);
or U18431 (N_18431,N_17113,N_17384);
and U18432 (N_18432,N_17425,N_16837);
nor U18433 (N_18433,N_17493,N_17138);
xor U18434 (N_18434,N_17413,N_17258);
nand U18435 (N_18435,N_16794,N_16301);
or U18436 (N_18436,N_17350,N_16794);
or U18437 (N_18437,N_16337,N_17422);
nand U18438 (N_18438,N_17166,N_16841);
nor U18439 (N_18439,N_17150,N_17303);
nand U18440 (N_18440,N_16325,N_16785);
nand U18441 (N_18441,N_17221,N_17468);
nand U18442 (N_18442,N_17305,N_17140);
and U18443 (N_18443,N_17181,N_17493);
or U18444 (N_18444,N_17398,N_17406);
or U18445 (N_18445,N_17273,N_16743);
or U18446 (N_18446,N_17250,N_16405);
and U18447 (N_18447,N_17099,N_16283);
nand U18448 (N_18448,N_16561,N_16500);
nor U18449 (N_18449,N_16956,N_16978);
xnor U18450 (N_18450,N_16717,N_17251);
or U18451 (N_18451,N_17346,N_17019);
or U18452 (N_18452,N_17277,N_16847);
nor U18453 (N_18453,N_17458,N_16787);
nand U18454 (N_18454,N_17482,N_17274);
nor U18455 (N_18455,N_17266,N_17260);
xnor U18456 (N_18456,N_16736,N_16457);
and U18457 (N_18457,N_16406,N_16276);
and U18458 (N_18458,N_16348,N_16854);
and U18459 (N_18459,N_16926,N_16446);
and U18460 (N_18460,N_16669,N_16292);
xnor U18461 (N_18461,N_16432,N_16671);
or U18462 (N_18462,N_16317,N_17433);
nor U18463 (N_18463,N_16475,N_16470);
or U18464 (N_18464,N_16551,N_17121);
nand U18465 (N_18465,N_16322,N_17047);
xor U18466 (N_18466,N_17016,N_16665);
and U18467 (N_18467,N_17408,N_17186);
xnor U18468 (N_18468,N_17267,N_17230);
nand U18469 (N_18469,N_16597,N_16367);
nand U18470 (N_18470,N_16605,N_17467);
nand U18471 (N_18471,N_17017,N_17416);
xor U18472 (N_18472,N_17161,N_17028);
xor U18473 (N_18473,N_17029,N_16390);
nor U18474 (N_18474,N_17198,N_17374);
or U18475 (N_18475,N_16806,N_16599);
and U18476 (N_18476,N_16566,N_16756);
nand U18477 (N_18477,N_16442,N_16271);
and U18478 (N_18478,N_16488,N_16357);
and U18479 (N_18479,N_16688,N_16886);
nor U18480 (N_18480,N_16617,N_16279);
nand U18481 (N_18481,N_16499,N_16918);
nor U18482 (N_18482,N_16649,N_16896);
nor U18483 (N_18483,N_16523,N_17287);
and U18484 (N_18484,N_17127,N_17458);
nor U18485 (N_18485,N_17449,N_17056);
nand U18486 (N_18486,N_17366,N_16450);
or U18487 (N_18487,N_17075,N_16356);
nor U18488 (N_18488,N_16469,N_16674);
xor U18489 (N_18489,N_17446,N_16781);
or U18490 (N_18490,N_16529,N_16258);
or U18491 (N_18491,N_16471,N_17167);
nor U18492 (N_18492,N_17004,N_16617);
xor U18493 (N_18493,N_17165,N_17376);
and U18494 (N_18494,N_16423,N_16998);
nand U18495 (N_18495,N_17156,N_16715);
nor U18496 (N_18496,N_16495,N_17380);
and U18497 (N_18497,N_16923,N_16695);
and U18498 (N_18498,N_16759,N_16442);
xnor U18499 (N_18499,N_16867,N_17005);
and U18500 (N_18500,N_17249,N_16967);
nor U18501 (N_18501,N_16703,N_17008);
and U18502 (N_18502,N_16877,N_17284);
and U18503 (N_18503,N_17085,N_16257);
xnor U18504 (N_18504,N_16473,N_16533);
and U18505 (N_18505,N_16634,N_17199);
and U18506 (N_18506,N_16780,N_17414);
xor U18507 (N_18507,N_16647,N_17425);
and U18508 (N_18508,N_17370,N_16607);
nor U18509 (N_18509,N_16705,N_17466);
or U18510 (N_18510,N_16748,N_16752);
nand U18511 (N_18511,N_16867,N_17218);
xnor U18512 (N_18512,N_16304,N_17038);
nor U18513 (N_18513,N_17403,N_17141);
nand U18514 (N_18514,N_17055,N_16571);
nand U18515 (N_18515,N_17201,N_17309);
nor U18516 (N_18516,N_17368,N_16929);
and U18517 (N_18517,N_17239,N_16507);
xor U18518 (N_18518,N_17446,N_16624);
nor U18519 (N_18519,N_16679,N_16728);
or U18520 (N_18520,N_16591,N_17418);
and U18521 (N_18521,N_17311,N_17355);
nand U18522 (N_18522,N_17038,N_16755);
nor U18523 (N_18523,N_16999,N_16656);
or U18524 (N_18524,N_16452,N_17434);
nor U18525 (N_18525,N_16787,N_16753);
and U18526 (N_18526,N_16886,N_16560);
or U18527 (N_18527,N_17131,N_17431);
and U18528 (N_18528,N_16285,N_16576);
and U18529 (N_18529,N_16901,N_16956);
xnor U18530 (N_18530,N_17403,N_16747);
and U18531 (N_18531,N_16487,N_17273);
nor U18532 (N_18532,N_17379,N_17130);
or U18533 (N_18533,N_17491,N_17133);
and U18534 (N_18534,N_16483,N_16828);
xor U18535 (N_18535,N_16485,N_17324);
and U18536 (N_18536,N_16940,N_16881);
and U18537 (N_18537,N_17324,N_17192);
or U18538 (N_18538,N_17387,N_16928);
or U18539 (N_18539,N_17216,N_16571);
xor U18540 (N_18540,N_16313,N_16642);
xor U18541 (N_18541,N_17048,N_16817);
nor U18542 (N_18542,N_16871,N_17304);
nand U18543 (N_18543,N_16933,N_17258);
nand U18544 (N_18544,N_16306,N_16589);
or U18545 (N_18545,N_16655,N_17257);
nor U18546 (N_18546,N_16550,N_16493);
and U18547 (N_18547,N_16717,N_16907);
nand U18548 (N_18548,N_16943,N_16962);
and U18549 (N_18549,N_16271,N_17203);
nand U18550 (N_18550,N_16930,N_16252);
nand U18551 (N_18551,N_16584,N_17342);
nand U18552 (N_18552,N_17165,N_16315);
nor U18553 (N_18553,N_17140,N_17161);
and U18554 (N_18554,N_16886,N_17232);
nand U18555 (N_18555,N_16672,N_17155);
nand U18556 (N_18556,N_16694,N_16556);
or U18557 (N_18557,N_17129,N_17321);
or U18558 (N_18558,N_17415,N_16826);
nor U18559 (N_18559,N_17403,N_16267);
nor U18560 (N_18560,N_17162,N_16730);
and U18561 (N_18561,N_17134,N_16395);
or U18562 (N_18562,N_16622,N_16853);
xnor U18563 (N_18563,N_16735,N_16968);
or U18564 (N_18564,N_17414,N_16641);
xnor U18565 (N_18565,N_16847,N_16303);
nor U18566 (N_18566,N_16805,N_16682);
and U18567 (N_18567,N_17376,N_16890);
nor U18568 (N_18568,N_17230,N_17358);
xnor U18569 (N_18569,N_16835,N_17316);
xnor U18570 (N_18570,N_16833,N_16877);
nor U18571 (N_18571,N_16515,N_16263);
nor U18572 (N_18572,N_16486,N_16880);
and U18573 (N_18573,N_17007,N_17010);
xor U18574 (N_18574,N_17039,N_17331);
nor U18575 (N_18575,N_16536,N_16999);
nor U18576 (N_18576,N_17026,N_17349);
or U18577 (N_18577,N_16998,N_16776);
and U18578 (N_18578,N_16853,N_17298);
and U18579 (N_18579,N_17045,N_17056);
nor U18580 (N_18580,N_16415,N_17231);
or U18581 (N_18581,N_17245,N_16964);
nor U18582 (N_18582,N_17166,N_17288);
xnor U18583 (N_18583,N_17297,N_16564);
and U18584 (N_18584,N_16533,N_16393);
nand U18585 (N_18585,N_16323,N_17445);
xor U18586 (N_18586,N_16819,N_17232);
nand U18587 (N_18587,N_16618,N_17196);
xor U18588 (N_18588,N_16453,N_16910);
or U18589 (N_18589,N_16281,N_16538);
nand U18590 (N_18590,N_16955,N_16852);
or U18591 (N_18591,N_16533,N_17164);
nand U18592 (N_18592,N_16572,N_17226);
and U18593 (N_18593,N_16557,N_16399);
nor U18594 (N_18594,N_16452,N_16475);
nor U18595 (N_18595,N_16697,N_16691);
or U18596 (N_18596,N_16891,N_16885);
xnor U18597 (N_18597,N_16867,N_16693);
xnor U18598 (N_18598,N_16644,N_17318);
and U18599 (N_18599,N_17190,N_17443);
or U18600 (N_18600,N_16983,N_17286);
xnor U18601 (N_18601,N_16307,N_16972);
and U18602 (N_18602,N_16662,N_17302);
and U18603 (N_18603,N_16994,N_16969);
and U18604 (N_18604,N_17134,N_17040);
xor U18605 (N_18605,N_16626,N_16569);
and U18606 (N_18606,N_17481,N_17145);
xnor U18607 (N_18607,N_17042,N_17104);
or U18608 (N_18608,N_17429,N_16901);
or U18609 (N_18609,N_17098,N_17489);
nor U18610 (N_18610,N_17346,N_16511);
and U18611 (N_18611,N_17100,N_17254);
nor U18612 (N_18612,N_17396,N_17263);
nor U18613 (N_18613,N_17214,N_16313);
nor U18614 (N_18614,N_17224,N_17256);
nor U18615 (N_18615,N_17285,N_16461);
nor U18616 (N_18616,N_17378,N_16936);
nor U18617 (N_18617,N_17022,N_17056);
and U18618 (N_18618,N_17120,N_17151);
or U18619 (N_18619,N_16885,N_17397);
or U18620 (N_18620,N_17478,N_16735);
nand U18621 (N_18621,N_16409,N_16811);
or U18622 (N_18622,N_16449,N_16903);
or U18623 (N_18623,N_17430,N_17432);
nor U18624 (N_18624,N_16330,N_17424);
and U18625 (N_18625,N_16449,N_16777);
or U18626 (N_18626,N_16287,N_17057);
nand U18627 (N_18627,N_16630,N_16440);
or U18628 (N_18628,N_17352,N_16305);
or U18629 (N_18629,N_16401,N_16633);
xnor U18630 (N_18630,N_16892,N_16444);
nor U18631 (N_18631,N_16625,N_16965);
nor U18632 (N_18632,N_16725,N_16958);
or U18633 (N_18633,N_16949,N_17194);
xor U18634 (N_18634,N_16975,N_16565);
nand U18635 (N_18635,N_17245,N_16813);
or U18636 (N_18636,N_16619,N_17125);
xnor U18637 (N_18637,N_17286,N_16926);
and U18638 (N_18638,N_16361,N_16544);
and U18639 (N_18639,N_16310,N_16822);
xnor U18640 (N_18640,N_16329,N_16257);
nand U18641 (N_18641,N_16688,N_17071);
xnor U18642 (N_18642,N_16951,N_17334);
or U18643 (N_18643,N_17498,N_16435);
xor U18644 (N_18644,N_16300,N_17458);
nor U18645 (N_18645,N_16763,N_16491);
nand U18646 (N_18646,N_17309,N_16294);
and U18647 (N_18647,N_17418,N_17108);
or U18648 (N_18648,N_16510,N_16684);
or U18649 (N_18649,N_16803,N_16720);
and U18650 (N_18650,N_17322,N_16557);
and U18651 (N_18651,N_16952,N_17199);
xor U18652 (N_18652,N_16523,N_16726);
and U18653 (N_18653,N_17149,N_16400);
xor U18654 (N_18654,N_17177,N_16372);
nand U18655 (N_18655,N_17229,N_17352);
xor U18656 (N_18656,N_16451,N_16874);
nor U18657 (N_18657,N_17296,N_17267);
nor U18658 (N_18658,N_16284,N_17100);
xor U18659 (N_18659,N_16683,N_16949);
nor U18660 (N_18660,N_17498,N_16501);
and U18661 (N_18661,N_16871,N_17346);
nor U18662 (N_18662,N_17391,N_16753);
xnor U18663 (N_18663,N_17092,N_17304);
and U18664 (N_18664,N_17104,N_16772);
xor U18665 (N_18665,N_16308,N_17400);
and U18666 (N_18666,N_16380,N_17373);
nand U18667 (N_18667,N_16551,N_17077);
and U18668 (N_18668,N_16634,N_17482);
or U18669 (N_18669,N_16306,N_17358);
or U18670 (N_18670,N_16282,N_17211);
xnor U18671 (N_18671,N_16310,N_16888);
and U18672 (N_18672,N_16760,N_16471);
or U18673 (N_18673,N_17471,N_17074);
nor U18674 (N_18674,N_16353,N_16858);
and U18675 (N_18675,N_17261,N_16336);
nor U18676 (N_18676,N_16738,N_16900);
xnor U18677 (N_18677,N_16467,N_16276);
nand U18678 (N_18678,N_16931,N_16334);
or U18679 (N_18679,N_17453,N_17487);
nand U18680 (N_18680,N_16715,N_17199);
nor U18681 (N_18681,N_16840,N_16375);
or U18682 (N_18682,N_16281,N_17034);
and U18683 (N_18683,N_16834,N_17360);
nor U18684 (N_18684,N_16417,N_16451);
nand U18685 (N_18685,N_17065,N_17474);
or U18686 (N_18686,N_17393,N_16899);
nor U18687 (N_18687,N_17045,N_16931);
and U18688 (N_18688,N_16718,N_17185);
or U18689 (N_18689,N_16268,N_16536);
nor U18690 (N_18690,N_17195,N_16976);
and U18691 (N_18691,N_17442,N_16255);
and U18692 (N_18692,N_17203,N_17409);
xnor U18693 (N_18693,N_16299,N_16678);
nand U18694 (N_18694,N_16970,N_17446);
nand U18695 (N_18695,N_16437,N_17352);
and U18696 (N_18696,N_17248,N_16710);
nand U18697 (N_18697,N_17206,N_17276);
or U18698 (N_18698,N_17032,N_17217);
or U18699 (N_18699,N_16918,N_16643);
xor U18700 (N_18700,N_16899,N_16481);
and U18701 (N_18701,N_17083,N_16645);
nand U18702 (N_18702,N_17033,N_16983);
nand U18703 (N_18703,N_17481,N_16520);
nand U18704 (N_18704,N_17389,N_17409);
nand U18705 (N_18705,N_16254,N_17260);
and U18706 (N_18706,N_17341,N_16346);
nand U18707 (N_18707,N_17061,N_16728);
nor U18708 (N_18708,N_16689,N_16625);
nand U18709 (N_18709,N_16828,N_16311);
xnor U18710 (N_18710,N_16569,N_17386);
nand U18711 (N_18711,N_17202,N_17280);
nor U18712 (N_18712,N_17198,N_16644);
and U18713 (N_18713,N_16957,N_16643);
and U18714 (N_18714,N_17232,N_17186);
nand U18715 (N_18715,N_16887,N_16390);
nand U18716 (N_18716,N_16353,N_16692);
nor U18717 (N_18717,N_16569,N_16519);
or U18718 (N_18718,N_17018,N_16580);
and U18719 (N_18719,N_17381,N_17485);
nand U18720 (N_18720,N_17037,N_16420);
or U18721 (N_18721,N_16904,N_16318);
nor U18722 (N_18722,N_16312,N_17005);
nand U18723 (N_18723,N_16489,N_16983);
nor U18724 (N_18724,N_17080,N_16281);
and U18725 (N_18725,N_16795,N_17141);
nor U18726 (N_18726,N_16716,N_17013);
xnor U18727 (N_18727,N_16868,N_17491);
xor U18728 (N_18728,N_16979,N_16981);
nor U18729 (N_18729,N_16809,N_16870);
nand U18730 (N_18730,N_17105,N_17220);
or U18731 (N_18731,N_16675,N_17036);
xor U18732 (N_18732,N_16597,N_16315);
or U18733 (N_18733,N_17374,N_17071);
or U18734 (N_18734,N_16376,N_17274);
nand U18735 (N_18735,N_16525,N_16948);
or U18736 (N_18736,N_17129,N_17216);
xnor U18737 (N_18737,N_17491,N_16998);
or U18738 (N_18738,N_16954,N_16251);
and U18739 (N_18739,N_16566,N_16410);
or U18740 (N_18740,N_17141,N_16818);
nand U18741 (N_18741,N_16370,N_16592);
xor U18742 (N_18742,N_17087,N_16662);
and U18743 (N_18743,N_16835,N_16832);
nor U18744 (N_18744,N_17005,N_17203);
xor U18745 (N_18745,N_16418,N_17039);
nand U18746 (N_18746,N_16476,N_16852);
and U18747 (N_18747,N_17473,N_17305);
xor U18748 (N_18748,N_17483,N_16294);
or U18749 (N_18749,N_16665,N_17496);
and U18750 (N_18750,N_18264,N_18287);
xnor U18751 (N_18751,N_18472,N_17931);
nand U18752 (N_18752,N_18466,N_18276);
and U18753 (N_18753,N_17663,N_18705);
nand U18754 (N_18754,N_18307,N_18223);
or U18755 (N_18755,N_18163,N_17774);
nor U18756 (N_18756,N_18405,N_18365);
or U18757 (N_18757,N_18039,N_18314);
and U18758 (N_18758,N_17706,N_17802);
or U18759 (N_18759,N_18310,N_18278);
and U18760 (N_18760,N_18660,N_17721);
nor U18761 (N_18761,N_17744,N_17712);
or U18762 (N_18762,N_17860,N_18052);
and U18763 (N_18763,N_17707,N_18411);
nand U18764 (N_18764,N_18316,N_18524);
nor U18765 (N_18765,N_18739,N_17697);
or U18766 (N_18766,N_17694,N_18549);
or U18767 (N_18767,N_17616,N_17560);
and U18768 (N_18768,N_18017,N_17859);
nor U18769 (N_18769,N_17577,N_18266);
xnor U18770 (N_18770,N_17564,N_18084);
nand U18771 (N_18771,N_18185,N_18409);
and U18772 (N_18772,N_18481,N_17785);
xnor U18773 (N_18773,N_17894,N_18697);
or U18774 (N_18774,N_18722,N_17834);
nand U18775 (N_18775,N_17809,N_18116);
nand U18776 (N_18776,N_18193,N_17923);
and U18777 (N_18777,N_18150,N_17557);
nand U18778 (N_18778,N_18249,N_17562);
and U18779 (N_18779,N_18237,N_18628);
or U18780 (N_18780,N_18572,N_18174);
and U18781 (N_18781,N_18347,N_18020);
or U18782 (N_18782,N_18568,N_17844);
nor U18783 (N_18783,N_18215,N_17905);
and U18784 (N_18784,N_17570,N_18669);
and U18785 (N_18785,N_18344,N_17530);
nor U18786 (N_18786,N_17730,N_18312);
and U18787 (N_18787,N_18746,N_17546);
and U18788 (N_18788,N_18086,N_18681);
or U18789 (N_18789,N_18128,N_17673);
or U18790 (N_18790,N_18233,N_18734);
nor U18791 (N_18791,N_18257,N_18170);
nand U18792 (N_18792,N_17637,N_17880);
and U18793 (N_18793,N_18304,N_18471);
nand U18794 (N_18794,N_17734,N_17680);
or U18795 (N_18795,N_18637,N_17563);
or U18796 (N_18796,N_18186,N_18557);
and U18797 (N_18797,N_17765,N_18033);
xor U18798 (N_18798,N_18200,N_18323);
nand U18799 (N_18799,N_17580,N_17764);
or U18800 (N_18800,N_18248,N_18535);
xor U18801 (N_18801,N_17925,N_17622);
nand U18802 (N_18802,N_18674,N_17756);
and U18803 (N_18803,N_17757,N_17709);
and U18804 (N_18804,N_18723,N_17607);
nand U18805 (N_18805,N_18588,N_18007);
xor U18806 (N_18806,N_17889,N_17606);
nand U18807 (N_18807,N_18213,N_17733);
and U18808 (N_18808,N_17893,N_18520);
xor U18809 (N_18809,N_17897,N_18635);
or U18810 (N_18810,N_18726,N_18353);
nor U18811 (N_18811,N_17977,N_17961);
and U18812 (N_18812,N_18602,N_17542);
or U18813 (N_18813,N_18636,N_17520);
nand U18814 (N_18814,N_18601,N_18041);
xor U18815 (N_18815,N_18640,N_18350);
and U18816 (N_18816,N_18443,N_18262);
nor U18817 (N_18817,N_18491,N_18715);
and U18818 (N_18818,N_17821,N_17715);
nor U18819 (N_18819,N_18500,N_18013);
nor U18820 (N_18820,N_18188,N_17535);
or U18821 (N_18821,N_18127,N_18707);
or U18822 (N_18822,N_18258,N_17836);
and U18823 (N_18823,N_18085,N_18267);
and U18824 (N_18824,N_17888,N_18517);
nor U18825 (N_18825,N_18137,N_17918);
nor U18826 (N_18826,N_17526,N_18046);
nor U18827 (N_18827,N_17583,N_18704);
nor U18828 (N_18828,N_17735,N_18179);
nand U18829 (N_18829,N_18684,N_17674);
and U18830 (N_18830,N_17999,N_18748);
nor U18831 (N_18831,N_18232,N_18245);
or U18832 (N_18832,N_17725,N_17780);
and U18833 (N_18833,N_18690,N_18198);
nand U18834 (N_18834,N_18428,N_17509);
or U18835 (N_18835,N_17512,N_17521);
nand U18836 (N_18836,N_17758,N_17511);
and U18837 (N_18837,N_18358,N_17829);
or U18838 (N_18838,N_18173,N_18357);
and U18839 (N_18839,N_17991,N_18387);
nand U18840 (N_18840,N_17672,N_17784);
nor U18841 (N_18841,N_18247,N_18696);
xnor U18842 (N_18842,N_18082,N_17769);
xor U18843 (N_18843,N_18454,N_17936);
nor U18844 (N_18844,N_18093,N_18414);
and U18845 (N_18845,N_18489,N_18110);
xor U18846 (N_18846,N_18378,N_18080);
nand U18847 (N_18847,N_18418,N_18225);
xnor U18848 (N_18848,N_17996,N_17574);
or U18849 (N_18849,N_18587,N_17551);
xor U18850 (N_18850,N_18555,N_17742);
and U18851 (N_18851,N_18712,N_18625);
xor U18852 (N_18852,N_17679,N_18565);
nand U18853 (N_18853,N_18023,N_18590);
nor U18854 (N_18854,N_18457,N_18577);
nand U18855 (N_18855,N_17972,N_18112);
xor U18856 (N_18856,N_18009,N_18620);
nor U18857 (N_18857,N_17523,N_17945);
xor U18858 (N_18858,N_18528,N_17950);
xnor U18859 (N_18859,N_18716,N_17753);
and U18860 (N_18860,N_17561,N_18176);
and U18861 (N_18861,N_17656,N_18586);
nor U18862 (N_18862,N_18079,N_17746);
and U18863 (N_18863,N_17837,N_17921);
nor U18864 (N_18864,N_18741,N_17934);
or U18865 (N_18865,N_18283,N_18239);
nor U18866 (N_18866,N_17608,N_17932);
xnor U18867 (N_18867,N_17963,N_18400);
xnor U18868 (N_18868,N_17614,N_18594);
nor U18869 (N_18869,N_18146,N_18274);
xnor U18870 (N_18870,N_17502,N_17586);
nand U18871 (N_18871,N_17832,N_18218);
nand U18872 (N_18872,N_18497,N_18114);
and U18873 (N_18873,N_17724,N_18177);
or U18874 (N_18874,N_18412,N_18165);
or U18875 (N_18875,N_17857,N_18596);
nand U18876 (N_18876,N_18117,N_18332);
and U18877 (N_18877,N_18228,N_18180);
nand U18878 (N_18878,N_17875,N_18144);
nand U18879 (N_18879,N_18706,N_18210);
and U18880 (N_18880,N_17776,N_18534);
xor U18881 (N_18881,N_17675,N_18195);
nand U18882 (N_18882,N_18680,N_17532);
and U18883 (N_18883,N_18570,N_18003);
xnor U18884 (N_18884,N_18359,N_18703);
nand U18885 (N_18885,N_18465,N_18214);
and U18886 (N_18886,N_18121,N_18191);
nand U18887 (N_18887,N_18463,N_17545);
nor U18888 (N_18888,N_17669,N_18012);
and U18889 (N_18889,N_17567,N_18038);
nand U18890 (N_18890,N_17610,N_18429);
xor U18891 (N_18891,N_17942,N_18607);
nor U18892 (N_18892,N_17920,N_18404);
nor U18893 (N_18893,N_18611,N_18394);
nand U18894 (N_18894,N_18324,N_18675);
xor U18895 (N_18895,N_18139,N_17693);
xor U18896 (N_18896,N_18401,N_17946);
and U18897 (N_18897,N_17993,N_17529);
or U18898 (N_18898,N_17895,N_18686);
nand U18899 (N_18899,N_17591,N_18492);
xor U18900 (N_18900,N_18553,N_18682);
xor U18901 (N_18901,N_17791,N_18051);
or U18902 (N_18902,N_18000,N_18632);
and U18903 (N_18903,N_18496,N_18338);
nor U18904 (N_18904,N_17814,N_18091);
or U18905 (N_18905,N_17690,N_18380);
nand U18906 (N_18906,N_17685,N_17768);
and U18907 (N_18907,N_18280,N_18192);
xor U18908 (N_18908,N_17646,N_18385);
nand U18909 (N_18909,N_18364,N_18181);
or U18910 (N_18910,N_18279,N_18651);
or U18911 (N_18911,N_18419,N_18229);
nand U18912 (N_18912,N_18189,N_17850);
or U18913 (N_18913,N_17882,N_17877);
xor U18914 (N_18914,N_17617,N_18367);
nand U18915 (N_18915,N_18661,N_17536);
nor U18916 (N_18916,N_18202,N_18199);
xnor U18917 (N_18917,N_18689,N_17812);
xor U18918 (N_18918,N_18598,N_17909);
or U18919 (N_18919,N_18074,N_18356);
or U18920 (N_18920,N_18105,N_17632);
or U18921 (N_18921,N_17643,N_18360);
and U18922 (N_18922,N_17652,N_17726);
or U18923 (N_18923,N_17914,N_18135);
nand U18924 (N_18924,N_18349,N_18563);
nor U18925 (N_18925,N_17751,N_18479);
xor U18926 (N_18926,N_18334,N_18317);
or U18927 (N_18927,N_17667,N_18374);
and U18928 (N_18928,N_18488,N_17813);
xor U18929 (N_18929,N_17695,N_18442);
nor U18930 (N_18930,N_17896,N_18145);
or U18931 (N_18931,N_18536,N_18030);
and U18932 (N_18932,N_17696,N_17626);
and U18933 (N_18933,N_18355,N_17899);
and U18934 (N_18934,N_18194,N_18423);
nor U18935 (N_18935,N_18060,N_18544);
xor U18936 (N_18936,N_18441,N_17964);
nor U18937 (N_18937,N_18081,N_17736);
or U18938 (N_18938,N_18643,N_18325);
or U18939 (N_18939,N_17668,N_18475);
nor U18940 (N_18940,N_18345,N_17618);
nand U18941 (N_18941,N_18700,N_17929);
nor U18942 (N_18942,N_17940,N_17782);
nand U18943 (N_18943,N_18333,N_18119);
and U18944 (N_18944,N_18502,N_17910);
or U18945 (N_18945,N_17716,N_17600);
xnor U18946 (N_18946,N_18095,N_17830);
and U18947 (N_18947,N_18608,N_17554);
nand U18948 (N_18948,N_18271,N_17869);
nor U18949 (N_18949,N_18609,N_18432);
nor U18950 (N_18950,N_17794,N_17750);
nor U18951 (N_18951,N_17884,N_18453);
nor U18952 (N_18952,N_18425,N_18614);
nor U18953 (N_18953,N_18670,N_17901);
and U18954 (N_18954,N_18103,N_18571);
xnor U18955 (N_18955,N_18666,N_18040);
nand U18956 (N_18956,N_18284,N_18190);
nor U18957 (N_18957,N_17661,N_18075);
or U18958 (N_18958,N_18717,N_17777);
xor U18959 (N_18959,N_17689,N_18389);
xnor U18960 (N_18960,N_17933,N_18612);
nand U18961 (N_18961,N_18290,N_18542);
or U18962 (N_18962,N_18653,N_18123);
nand U18963 (N_18963,N_17941,N_18747);
nand U18964 (N_18964,N_17913,N_18499);
nor U18965 (N_18965,N_17788,N_18275);
nor U18966 (N_18966,N_17770,N_18527);
or U18967 (N_18967,N_18254,N_17579);
nor U18968 (N_18968,N_17633,N_17662);
nand U18969 (N_18969,N_17612,N_17822);
and U18970 (N_18970,N_18037,N_17846);
nor U18971 (N_18971,N_18659,N_18049);
xnor U18972 (N_18972,N_18291,N_18372);
and U18973 (N_18973,N_18390,N_18582);
and U18974 (N_18974,N_18595,N_18495);
and U18975 (N_18975,N_17639,N_17701);
and U18976 (N_18976,N_17902,N_17898);
and U18977 (N_18977,N_18483,N_17973);
or U18978 (N_18978,N_17823,N_18336);
nor U18979 (N_18979,N_17795,N_18448);
and U18980 (N_18980,N_18131,N_17852);
and U18981 (N_18981,N_17810,N_17702);
xnor U18982 (N_18982,N_17740,N_17870);
and U18983 (N_18983,N_18072,N_17981);
nor U18984 (N_18984,N_17534,N_18381);
or U18985 (N_18985,N_18560,N_18159);
nor U18986 (N_18986,N_18631,N_18731);
nor U18987 (N_18987,N_17767,N_17620);
nand U18988 (N_18988,N_18541,N_17856);
or U18989 (N_18989,N_18227,N_18226);
nand U18990 (N_18990,N_17628,N_18519);
or U18991 (N_18991,N_18071,N_18327);
or U18992 (N_18992,N_18109,N_17853);
xnor U18993 (N_18993,N_17518,N_17904);
or U18994 (N_18994,N_17660,N_18025);
or U18995 (N_18995,N_17503,N_17807);
nand U18996 (N_18996,N_17651,N_18664);
and U18997 (N_18997,N_17980,N_17760);
xnor U18998 (N_18998,N_17678,N_18222);
or U18999 (N_18999,N_18141,N_18521);
nand U19000 (N_19000,N_18298,N_18749);
nor U19001 (N_19001,N_17590,N_17816);
xor U19002 (N_19002,N_18610,N_17828);
xnor U19003 (N_19003,N_17500,N_18066);
nand U19004 (N_19004,N_17754,N_17833);
nor U19005 (N_19005,N_18580,N_17783);
and U19006 (N_19006,N_18050,N_17817);
xnor U19007 (N_19007,N_18576,N_18744);
nand U19008 (N_19008,N_18259,N_17581);
nor U19009 (N_19009,N_18140,N_18720);
nand U19010 (N_19010,N_18297,N_17949);
and U19011 (N_19011,N_18308,N_18263);
xor U19012 (N_19012,N_17826,N_17842);
nand U19013 (N_19013,N_17992,N_18016);
nor U19014 (N_19014,N_17858,N_17513);
xor U19015 (N_19015,N_18493,N_18008);
or U19016 (N_19016,N_18171,N_18398);
xnor U19017 (N_19017,N_17594,N_18099);
nand U19018 (N_19018,N_18311,N_17881);
or U19019 (N_19019,N_17625,N_18599);
or U19020 (N_19020,N_17719,N_18511);
nor U19021 (N_19021,N_18626,N_18231);
xor U19022 (N_19022,N_18124,N_18652);
nand U19023 (N_19023,N_18638,N_17623);
and U19024 (N_19024,N_18246,N_18092);
nor U19025 (N_19025,N_17575,N_18339);
or U19026 (N_19026,N_17762,N_18070);
or U19027 (N_19027,N_18467,N_18476);
and U19028 (N_19028,N_18004,N_17845);
nand U19029 (N_19029,N_17874,N_17516);
xnor U19030 (N_19030,N_17599,N_18474);
or U19031 (N_19031,N_17671,N_18444);
xor U19032 (N_19032,N_18745,N_18348);
and U19033 (N_19033,N_17863,N_17605);
and U19034 (N_19034,N_17939,N_17861);
xnor U19035 (N_19035,N_17501,N_18045);
or U19036 (N_19036,N_18002,N_18566);
and U19037 (N_19037,N_18581,N_17907);
nor U19038 (N_19038,N_18437,N_17772);
xor U19039 (N_19039,N_17843,N_18480);
and U19040 (N_19040,N_18106,N_17630);
and U19041 (N_19041,N_17631,N_17815);
nand U19042 (N_19042,N_18113,N_17995);
xnor U19043 (N_19043,N_17713,N_18593);
or U19044 (N_19044,N_17743,N_18011);
nand U19045 (N_19045,N_18629,N_18219);
xnor U19046 (N_19046,N_17952,N_18455);
xor U19047 (N_19047,N_18242,N_17808);
nor U19048 (N_19048,N_18592,N_18294);
xnor U19049 (N_19049,N_18209,N_18439);
nand U19050 (N_19050,N_18721,N_18505);
or U19051 (N_19051,N_18343,N_18416);
nor U19052 (N_19052,N_18073,N_17990);
or U19053 (N_19053,N_17647,N_18313);
nand U19054 (N_19054,N_17926,N_17958);
nor U19055 (N_19055,N_17773,N_18067);
nand U19056 (N_19056,N_18083,N_18162);
or U19057 (N_19057,N_17699,N_18477);
and U19058 (N_19058,N_17947,N_18440);
nor U19059 (N_19059,N_18044,N_18687);
and U19060 (N_19060,N_18167,N_17988);
xnor U19061 (N_19061,N_17510,N_17611);
or U19062 (N_19062,N_18515,N_17967);
nor U19063 (N_19063,N_18667,N_18464);
or U19064 (N_19064,N_17944,N_18406);
xor U19065 (N_19065,N_18305,N_18341);
nand U19066 (N_19066,N_17571,N_17885);
nand U19067 (N_19067,N_17872,N_17820);
or U19068 (N_19068,N_18513,N_18714);
xor U19069 (N_19069,N_18244,N_18402);
and U19070 (N_19070,N_17835,N_18584);
nor U19071 (N_19071,N_17759,N_18111);
and U19072 (N_19072,N_17714,N_17705);
or U19073 (N_19073,N_18330,N_18693);
or U19074 (N_19074,N_18329,N_18583);
and U19075 (N_19075,N_17969,N_18371);
or U19076 (N_19076,N_18328,N_18470);
nand U19077 (N_19077,N_17555,N_18024);
xnor U19078 (N_19078,N_17670,N_17737);
nand U19079 (N_19079,N_18393,N_18654);
nor U19080 (N_19080,N_18270,N_17576);
or U19081 (N_19081,N_18035,N_18063);
nand U19082 (N_19082,N_18695,N_18136);
and U19083 (N_19083,N_18379,N_17819);
nand U19084 (N_19084,N_18561,N_18574);
or U19085 (N_19085,N_17708,N_18685);
nand U19086 (N_19086,N_17650,N_17866);
nand U19087 (N_19087,N_17641,N_18624);
nor U19088 (N_19088,N_18567,N_17922);
nand U19089 (N_19089,N_18164,N_17627);
nand U19090 (N_19090,N_18613,N_17524);
nor U19091 (N_19091,N_18363,N_17798);
and U19092 (N_19092,N_18203,N_18711);
xor U19093 (N_19093,N_18537,N_18713);
and U19094 (N_19094,N_17505,N_18143);
and U19095 (N_19095,N_18473,N_17644);
xor U19096 (N_19096,N_18427,N_18320);
xor U19097 (N_19097,N_18318,N_17558);
nand U19098 (N_19098,N_18391,N_18322);
xnor U19099 (N_19099,N_17738,N_18207);
xor U19100 (N_19100,N_18692,N_17873);
nor U19101 (N_19101,N_18054,N_17722);
or U19102 (N_19102,N_17635,N_18420);
nand U19103 (N_19103,N_18399,N_17710);
or U19104 (N_19104,N_18028,N_18742);
nor U19105 (N_19105,N_18518,N_17659);
nor U19106 (N_19106,N_18042,N_17589);
xor U19107 (N_19107,N_18384,N_17839);
or U19108 (N_19108,N_18450,N_18281);
and U19109 (N_19109,N_18445,N_18047);
and U19110 (N_19110,N_18386,N_17803);
nor U19111 (N_19111,N_17615,N_17504);
or U19112 (N_19112,N_18240,N_18014);
or U19113 (N_19113,N_17766,N_18005);
or U19114 (N_19114,N_17911,N_18677);
or U19115 (N_19115,N_17919,N_18148);
and U19116 (N_19116,N_18646,N_17649);
nand U19117 (N_19117,N_18478,N_17723);
nand U19118 (N_19118,N_17732,N_17704);
nor U19119 (N_19119,N_17686,N_17968);
or U19120 (N_19120,N_18168,N_17666);
nor U19121 (N_19121,N_18433,N_17544);
nor U19122 (N_19122,N_18649,N_17786);
xor U19123 (N_19123,N_18321,N_17636);
or U19124 (N_19124,N_17824,N_18289);
nor U19125 (N_19125,N_18510,N_17597);
nand U19126 (N_19126,N_18027,N_17789);
nor U19127 (N_19127,N_18260,N_18241);
nand U19128 (N_19128,N_18550,N_17556);
nor U19129 (N_19129,N_18370,N_18265);
xor U19130 (N_19130,N_18702,N_17588);
or U19131 (N_19131,N_18115,N_18134);
and U19132 (N_19132,N_18062,N_17531);
and U19133 (N_19133,N_18490,N_18569);
xnor U19134 (N_19134,N_18617,N_18648);
or U19135 (N_19135,N_17976,N_18373);
xor U19136 (N_19136,N_18514,N_18250);
and U19137 (N_19137,N_17975,N_18485);
nand U19138 (N_19138,N_17848,N_18238);
nor U19139 (N_19139,N_18383,N_17539);
and U19140 (N_19140,N_18430,N_18740);
nor U19141 (N_19141,N_17655,N_18337);
nand U19142 (N_19142,N_18034,N_18120);
and U19143 (N_19143,N_18048,N_18157);
xnor U19144 (N_19144,N_18104,N_18089);
nor U19145 (N_19145,N_18354,N_18306);
nor U19146 (N_19146,N_17868,N_18288);
or U19147 (N_19147,N_17514,N_18451);
and U19148 (N_19148,N_17886,N_18556);
nand U19149 (N_19149,N_18001,N_18619);
nand U19150 (N_19150,N_18107,N_18547);
and U19151 (N_19151,N_18392,N_18616);
nor U19152 (N_19152,N_18655,N_18299);
and U19153 (N_19153,N_18529,N_17878);
nand U19154 (N_19154,N_18057,N_18591);
nand U19155 (N_19155,N_17974,N_18484);
nor U19156 (N_19156,N_18633,N_18701);
nand U19157 (N_19157,N_17890,N_18340);
or U19158 (N_19158,N_17847,N_18126);
or U19159 (N_19159,N_18600,N_18447);
nand U19160 (N_19160,N_18197,N_18589);
xor U19161 (N_19161,N_17645,N_18078);
nor U19162 (N_19162,N_18132,N_18277);
nand U19163 (N_19163,N_18158,N_17887);
nor U19164 (N_19164,N_17747,N_17593);
and U19165 (N_19165,N_17519,N_17957);
and U19166 (N_19166,N_17982,N_17506);
xnor U19167 (N_19167,N_17998,N_18606);
and U19168 (N_19168,N_18382,N_18216);
xnor U19169 (N_19169,N_18413,N_17664);
xnor U19170 (N_19170,N_17688,N_17854);
nand U19171 (N_19171,N_18462,N_17965);
nand U19172 (N_19172,N_17609,N_17879);
xnor U19173 (N_19173,N_17537,N_17924);
nor U19174 (N_19174,N_18662,N_17749);
and U19175 (N_19175,N_18710,N_18417);
and U19176 (N_19176,N_18019,N_18508);
or U19177 (N_19177,N_17778,N_17515);
nor U19178 (N_19178,N_17797,N_18724);
and U19179 (N_19179,N_18644,N_18501);
nor U19180 (N_19180,N_17900,N_18368);
or U19181 (N_19181,N_18055,N_18282);
or U19182 (N_19182,N_17684,N_18388);
nor U19183 (N_19183,N_17796,N_18361);
or U19184 (N_19184,N_17790,N_18426);
xor U19185 (N_19185,N_17849,N_17891);
nor U19186 (N_19186,N_18183,N_17818);
or U19187 (N_19187,N_18639,N_18196);
nor U19188 (N_19188,N_18676,N_17987);
nor U19189 (N_19189,N_18053,N_17543);
nor U19190 (N_19190,N_18494,N_18509);
or U19191 (N_19191,N_18504,N_18579);
nand U19192 (N_19192,N_18506,N_18699);
and U19193 (N_19193,N_18261,N_18302);
or U19194 (N_19194,N_18331,N_18184);
nor U19195 (N_19195,N_18255,N_18498);
or U19196 (N_19196,N_18029,N_18152);
nand U19197 (N_19197,N_18187,N_18679);
nor U19198 (N_19198,N_17892,N_18458);
or U19199 (N_19199,N_18205,N_18395);
nand U19200 (N_19200,N_17805,N_17676);
nand U19201 (N_19201,N_18424,N_17569);
xor U19202 (N_19202,N_18036,N_18603);
nor U19203 (N_19203,N_18272,N_18551);
and U19204 (N_19204,N_18285,N_18068);
nand U19205 (N_19205,N_17739,N_18059);
xnor U19206 (N_19206,N_17522,N_17657);
nor U19207 (N_19207,N_17938,N_17989);
or U19208 (N_19208,N_18727,N_17642);
nor U19209 (N_19209,N_18621,N_18683);
nor U19210 (N_19210,N_17935,N_17917);
xnor U19211 (N_19211,N_17978,N_18461);
nand U19212 (N_19212,N_18220,N_18102);
nor U19213 (N_19213,N_17984,N_17953);
nor U19214 (N_19214,N_18096,N_18630);
nand U19215 (N_19215,N_17728,N_18545);
or U19216 (N_19216,N_18558,N_18147);
nor U19217 (N_19217,N_17775,N_17781);
nor U19218 (N_19218,N_18326,N_17827);
nand U19219 (N_19219,N_18018,N_17598);
or U19220 (N_19220,N_18292,N_17720);
nand U19221 (N_19221,N_17687,N_18303);
nand U19222 (N_19222,N_18065,N_18407);
xor U19223 (N_19223,N_18351,N_17584);
nand U19224 (N_19224,N_18069,N_17596);
xnor U19225 (N_19225,N_18236,N_17956);
nand U19226 (N_19226,N_18234,N_18154);
or U19227 (N_19227,N_17508,N_17578);
nor U19228 (N_19228,N_17937,N_18641);
and U19229 (N_19229,N_17871,N_18100);
nor U19230 (N_19230,N_18156,N_17613);
xnor U19231 (N_19231,N_18403,N_18268);
xor U19232 (N_19232,N_18342,N_18088);
nand U19233 (N_19233,N_17629,N_18032);
xnor U19234 (N_19234,N_17951,N_18108);
or U19235 (N_19235,N_17592,N_18431);
nor U19236 (N_19236,N_18737,N_18718);
nand U19237 (N_19237,N_18438,N_17800);
and U19238 (N_19238,N_18142,N_18155);
xor U19239 (N_19239,N_17717,N_18459);
nand U19240 (N_19240,N_17799,N_17986);
nand U19241 (N_19241,N_18087,N_18161);
nand U19242 (N_19242,N_18533,N_17533);
nor U19243 (N_19243,N_18252,N_17568);
xor U19244 (N_19244,N_18315,N_18396);
and U19245 (N_19245,N_17883,N_18286);
and U19246 (N_19246,N_18530,N_17634);
xor U19247 (N_19247,N_18204,N_17549);
nor U19248 (N_19248,N_18729,N_17654);
xor U19249 (N_19249,N_17729,N_18206);
nor U19250 (N_19250,N_17831,N_18452);
nor U19251 (N_19251,N_17550,N_18605);
or U19252 (N_19252,N_17681,N_17587);
xnor U19253 (N_19253,N_18169,N_17763);
and U19254 (N_19254,N_18369,N_17994);
and U19255 (N_19255,N_18319,N_17865);
xor U19256 (N_19256,N_17548,N_18296);
nand U19257 (N_19257,N_18709,N_18562);
nand U19258 (N_19258,N_18575,N_18251);
and U19259 (N_19259,N_17517,N_18456);
or U19260 (N_19260,N_17682,N_18658);
or U19261 (N_19261,N_18212,N_18634);
nand U19262 (N_19262,N_18436,N_17985);
nand U19263 (N_19263,N_18585,N_17638);
or U19264 (N_19264,N_18397,N_18077);
nand U19265 (N_19265,N_17553,N_18362);
and U19266 (N_19266,N_18094,N_18221);
and U19267 (N_19267,N_17698,N_18552);
nor U19268 (N_19268,N_18058,N_18573);
and U19269 (N_19269,N_17876,N_18482);
nand U19270 (N_19270,N_18522,N_17566);
and U19271 (N_19271,N_18149,N_18719);
and U19272 (N_19272,N_18293,N_18656);
xnor U19273 (N_19273,N_17841,N_17983);
and U19274 (N_19274,N_18523,N_18597);
xor U19275 (N_19275,N_17711,N_18129);
xor U19276 (N_19276,N_17801,N_17761);
and U19277 (N_19277,N_17811,N_17624);
and U19278 (N_19278,N_17538,N_18578);
nand U19279 (N_19279,N_17838,N_17601);
or U19280 (N_19280,N_17540,N_18446);
nand U19281 (N_19281,N_17912,N_17928);
and U19282 (N_19282,N_18732,N_17525);
xor U19283 (N_19283,N_17867,N_18738);
xnor U19284 (N_19284,N_18604,N_17507);
and U19285 (N_19285,N_17943,N_17915);
nor U19286 (N_19286,N_18623,N_18300);
nor U19287 (N_19287,N_17748,N_18671);
and U19288 (N_19288,N_17573,N_18516);
or U19289 (N_19289,N_18178,N_17962);
nor U19290 (N_19290,N_17752,N_18064);
and U19291 (N_19291,N_18422,N_17948);
or U19292 (N_19292,N_18688,N_17851);
or U19293 (N_19293,N_18531,N_18301);
and U19294 (N_19294,N_18434,N_18026);
nand U19295 (N_19295,N_18243,N_17572);
or U19296 (N_19296,N_18098,N_17960);
or U19297 (N_19297,N_17665,N_18201);
nand U19298 (N_19298,N_17619,N_17604);
and U19299 (N_19299,N_18366,N_18101);
and U19300 (N_19300,N_17527,N_18021);
and U19301 (N_19301,N_17677,N_17692);
and U19302 (N_19302,N_18235,N_18468);
xnor U19303 (N_19303,N_18672,N_18090);
or U19304 (N_19304,N_18130,N_17966);
or U19305 (N_19305,N_18122,N_18554);
xnor U19306 (N_19306,N_17792,N_18487);
nand U19307 (N_19307,N_18151,N_18061);
and U19308 (N_19308,N_17603,N_17979);
xnor U19309 (N_19309,N_18253,N_17585);
nand U19310 (N_19310,N_18335,N_18532);
and U19311 (N_19311,N_18097,N_18076);
or U19312 (N_19312,N_18512,N_17653);
nand U19313 (N_19313,N_17541,N_17547);
or U19314 (N_19314,N_17930,N_18410);
nor U19315 (N_19315,N_18056,N_18460);
and U19316 (N_19316,N_18172,N_18736);
or U19317 (N_19317,N_17840,N_17582);
and U19318 (N_19318,N_18182,N_17779);
nor U19319 (N_19319,N_18153,N_17771);
nor U19320 (N_19320,N_17565,N_18622);
or U19321 (N_19321,N_18352,N_17903);
nor U19322 (N_19322,N_18118,N_18160);
and U19323 (N_19323,N_17691,N_18309);
xnor U19324 (N_19324,N_18469,N_17954);
nand U19325 (N_19325,N_18415,N_18376);
and U19326 (N_19326,N_17559,N_18125);
xnor U19327 (N_19327,N_18211,N_18377);
nand U19328 (N_19328,N_18691,N_17727);
and U19329 (N_19329,N_17658,N_18618);
and U19330 (N_19330,N_18022,N_18503);
nor U19331 (N_19331,N_18138,N_18698);
nand U19332 (N_19332,N_17552,N_18708);
and U19333 (N_19333,N_18694,N_18735);
nor U19334 (N_19334,N_18526,N_18408);
and U19335 (N_19335,N_18486,N_18548);
or U19336 (N_19336,N_17906,N_17793);
and U19337 (N_19337,N_18539,N_17804);
or U19338 (N_19338,N_18295,N_17927);
and U19339 (N_19339,N_17595,N_17640);
or U19340 (N_19340,N_18043,N_17703);
or U19341 (N_19341,N_17806,N_18175);
xnor U19342 (N_19342,N_18725,N_18449);
and U19343 (N_19343,N_17855,N_18543);
nor U19344 (N_19344,N_18743,N_18647);
and U19345 (N_19345,N_18540,N_18421);
or U19346 (N_19346,N_18730,N_17862);
or U19347 (N_19347,N_18230,N_18546);
nor U19348 (N_19348,N_17908,N_18375);
nand U19349 (N_19349,N_17755,N_18208);
nor U19350 (N_19350,N_17731,N_17916);
or U19351 (N_19351,N_17997,N_18668);
nor U19352 (N_19352,N_18166,N_18678);
nor U19353 (N_19353,N_17602,N_17970);
or U19354 (N_19354,N_18435,N_17683);
nand U19355 (N_19355,N_18006,N_18538);
nor U19356 (N_19356,N_18133,N_18657);
or U19357 (N_19357,N_18645,N_18273);
or U19358 (N_19358,N_17825,N_18665);
or U19359 (N_19359,N_18031,N_18733);
nand U19360 (N_19360,N_17700,N_18650);
nand U19361 (N_19361,N_18010,N_18256);
and U19362 (N_19362,N_17787,N_18217);
xor U19363 (N_19363,N_18673,N_18663);
nand U19364 (N_19364,N_18346,N_17955);
nor U19365 (N_19365,N_17621,N_18507);
nor U19366 (N_19366,N_18627,N_17648);
or U19367 (N_19367,N_18564,N_17864);
and U19368 (N_19368,N_18728,N_18525);
xnor U19369 (N_19369,N_18224,N_18269);
xor U19370 (N_19370,N_18615,N_17745);
nor U19371 (N_19371,N_18559,N_17741);
and U19372 (N_19372,N_17528,N_17971);
xnor U19373 (N_19373,N_18642,N_18015);
xor U19374 (N_19374,N_17959,N_17718);
and U19375 (N_19375,N_17846,N_18383);
nor U19376 (N_19376,N_17620,N_18682);
xnor U19377 (N_19377,N_17728,N_17732);
nor U19378 (N_19378,N_18531,N_17624);
nand U19379 (N_19379,N_17929,N_18299);
and U19380 (N_19380,N_18358,N_18300);
xor U19381 (N_19381,N_18290,N_17797);
or U19382 (N_19382,N_18411,N_17541);
and U19383 (N_19383,N_18221,N_17746);
nor U19384 (N_19384,N_18676,N_18555);
xnor U19385 (N_19385,N_17912,N_17945);
nor U19386 (N_19386,N_18156,N_17985);
nor U19387 (N_19387,N_17986,N_17911);
xnor U19388 (N_19388,N_18027,N_18686);
xnor U19389 (N_19389,N_18724,N_18296);
nand U19390 (N_19390,N_17635,N_18193);
nor U19391 (N_19391,N_18311,N_17597);
nand U19392 (N_19392,N_18630,N_18708);
and U19393 (N_19393,N_17849,N_17630);
nor U19394 (N_19394,N_18728,N_18595);
nor U19395 (N_19395,N_18101,N_18417);
xnor U19396 (N_19396,N_17610,N_17706);
and U19397 (N_19397,N_18389,N_18341);
or U19398 (N_19398,N_17798,N_17695);
nor U19399 (N_19399,N_18560,N_17721);
nor U19400 (N_19400,N_17987,N_17642);
nand U19401 (N_19401,N_17892,N_17861);
or U19402 (N_19402,N_17776,N_18343);
xnor U19403 (N_19403,N_18266,N_17587);
nor U19404 (N_19404,N_18463,N_18471);
nor U19405 (N_19405,N_18280,N_17962);
or U19406 (N_19406,N_18576,N_18585);
and U19407 (N_19407,N_18288,N_17794);
nor U19408 (N_19408,N_18212,N_17683);
nand U19409 (N_19409,N_18064,N_17820);
or U19410 (N_19410,N_18246,N_18489);
nand U19411 (N_19411,N_18398,N_18698);
or U19412 (N_19412,N_17514,N_17802);
or U19413 (N_19413,N_18394,N_18391);
nand U19414 (N_19414,N_17944,N_18520);
nand U19415 (N_19415,N_17959,N_18553);
xnor U19416 (N_19416,N_18486,N_18718);
nor U19417 (N_19417,N_17658,N_17517);
nand U19418 (N_19418,N_18015,N_17853);
nor U19419 (N_19419,N_18210,N_18347);
nand U19420 (N_19420,N_18051,N_17532);
xor U19421 (N_19421,N_17732,N_18512);
nand U19422 (N_19422,N_17561,N_17742);
or U19423 (N_19423,N_18447,N_17749);
nand U19424 (N_19424,N_18280,N_18028);
and U19425 (N_19425,N_18124,N_18021);
xnor U19426 (N_19426,N_18739,N_17559);
xor U19427 (N_19427,N_17953,N_18355);
or U19428 (N_19428,N_17632,N_17983);
nand U19429 (N_19429,N_17691,N_17773);
and U19430 (N_19430,N_18531,N_17796);
xnor U19431 (N_19431,N_17736,N_17690);
xnor U19432 (N_19432,N_18018,N_17636);
nor U19433 (N_19433,N_18521,N_17599);
xor U19434 (N_19434,N_18171,N_18167);
xnor U19435 (N_19435,N_17581,N_18267);
xor U19436 (N_19436,N_18630,N_18053);
nand U19437 (N_19437,N_18211,N_18600);
xnor U19438 (N_19438,N_17754,N_18223);
xnor U19439 (N_19439,N_18203,N_17626);
nor U19440 (N_19440,N_18477,N_17997);
xor U19441 (N_19441,N_18435,N_18411);
nor U19442 (N_19442,N_17770,N_18613);
nand U19443 (N_19443,N_18063,N_18651);
and U19444 (N_19444,N_17815,N_18203);
or U19445 (N_19445,N_18308,N_17938);
and U19446 (N_19446,N_18392,N_18571);
and U19447 (N_19447,N_17538,N_18589);
and U19448 (N_19448,N_17663,N_18498);
xor U19449 (N_19449,N_18093,N_18057);
or U19450 (N_19450,N_17795,N_17805);
nand U19451 (N_19451,N_18092,N_17748);
xor U19452 (N_19452,N_17736,N_18652);
nor U19453 (N_19453,N_17669,N_18571);
nand U19454 (N_19454,N_18165,N_18301);
xnor U19455 (N_19455,N_18294,N_17602);
xnor U19456 (N_19456,N_18599,N_17883);
xnor U19457 (N_19457,N_17612,N_18368);
xnor U19458 (N_19458,N_17850,N_18017);
or U19459 (N_19459,N_18267,N_18596);
nor U19460 (N_19460,N_17986,N_17716);
or U19461 (N_19461,N_17791,N_18090);
nor U19462 (N_19462,N_18658,N_18091);
nor U19463 (N_19463,N_18145,N_18030);
nand U19464 (N_19464,N_18324,N_17949);
nand U19465 (N_19465,N_17715,N_18325);
xnor U19466 (N_19466,N_18078,N_17557);
and U19467 (N_19467,N_17823,N_17528);
nor U19468 (N_19468,N_18633,N_18576);
nand U19469 (N_19469,N_17580,N_17775);
nand U19470 (N_19470,N_18615,N_17679);
or U19471 (N_19471,N_18123,N_18269);
nand U19472 (N_19472,N_18579,N_18210);
xor U19473 (N_19473,N_18423,N_18074);
xor U19474 (N_19474,N_18489,N_17758);
nand U19475 (N_19475,N_18136,N_18655);
xnor U19476 (N_19476,N_18461,N_17793);
and U19477 (N_19477,N_17841,N_18115);
nand U19478 (N_19478,N_18342,N_18281);
or U19479 (N_19479,N_18594,N_17847);
nand U19480 (N_19480,N_18305,N_18626);
nand U19481 (N_19481,N_17621,N_17623);
and U19482 (N_19482,N_18449,N_18532);
nand U19483 (N_19483,N_18279,N_18107);
nor U19484 (N_19484,N_18056,N_18139);
nand U19485 (N_19485,N_18535,N_17814);
nor U19486 (N_19486,N_18703,N_18461);
or U19487 (N_19487,N_17827,N_18455);
nor U19488 (N_19488,N_17946,N_18697);
or U19489 (N_19489,N_18681,N_18304);
xor U19490 (N_19490,N_18726,N_17816);
and U19491 (N_19491,N_18498,N_17965);
nor U19492 (N_19492,N_17799,N_18265);
nand U19493 (N_19493,N_17505,N_18116);
nand U19494 (N_19494,N_18125,N_18069);
nor U19495 (N_19495,N_18619,N_17937);
nor U19496 (N_19496,N_18313,N_18285);
nor U19497 (N_19497,N_17854,N_18463);
or U19498 (N_19498,N_18268,N_17620);
xor U19499 (N_19499,N_18317,N_18296);
or U19500 (N_19500,N_18463,N_17989);
xnor U19501 (N_19501,N_18371,N_17965);
xnor U19502 (N_19502,N_17719,N_18337);
xnor U19503 (N_19503,N_18474,N_18109);
nor U19504 (N_19504,N_18415,N_18040);
nand U19505 (N_19505,N_17770,N_18117);
xnor U19506 (N_19506,N_18301,N_18362);
and U19507 (N_19507,N_18455,N_18124);
and U19508 (N_19508,N_18460,N_17616);
or U19509 (N_19509,N_17523,N_17765);
and U19510 (N_19510,N_18463,N_17876);
nor U19511 (N_19511,N_17581,N_17692);
xor U19512 (N_19512,N_18527,N_17525);
nor U19513 (N_19513,N_17502,N_18524);
nand U19514 (N_19514,N_17883,N_18154);
and U19515 (N_19515,N_17811,N_18549);
nand U19516 (N_19516,N_17904,N_18180);
nand U19517 (N_19517,N_18359,N_17606);
nor U19518 (N_19518,N_18291,N_18466);
and U19519 (N_19519,N_17667,N_18240);
nand U19520 (N_19520,N_18029,N_18012);
or U19521 (N_19521,N_18095,N_18072);
nand U19522 (N_19522,N_17552,N_17643);
or U19523 (N_19523,N_17695,N_18443);
nand U19524 (N_19524,N_18449,N_18055);
nor U19525 (N_19525,N_18046,N_17608);
nand U19526 (N_19526,N_18590,N_18300);
nor U19527 (N_19527,N_17779,N_18074);
nand U19528 (N_19528,N_18062,N_18301);
nor U19529 (N_19529,N_18684,N_18187);
nand U19530 (N_19530,N_18231,N_18550);
xnor U19531 (N_19531,N_17637,N_18217);
nor U19532 (N_19532,N_18545,N_17709);
nand U19533 (N_19533,N_18148,N_18368);
nor U19534 (N_19534,N_17982,N_17871);
or U19535 (N_19535,N_18501,N_17772);
nor U19536 (N_19536,N_18369,N_18674);
and U19537 (N_19537,N_17999,N_18060);
nand U19538 (N_19538,N_18159,N_18276);
and U19539 (N_19539,N_17928,N_18662);
or U19540 (N_19540,N_17919,N_17573);
or U19541 (N_19541,N_18003,N_18327);
xor U19542 (N_19542,N_18046,N_18423);
xnor U19543 (N_19543,N_18150,N_17902);
nand U19544 (N_19544,N_18508,N_17582);
and U19545 (N_19545,N_18607,N_17702);
xor U19546 (N_19546,N_18711,N_18487);
xnor U19547 (N_19547,N_18622,N_18399);
or U19548 (N_19548,N_17529,N_18206);
xnor U19549 (N_19549,N_17501,N_17614);
nor U19550 (N_19550,N_17810,N_18729);
or U19551 (N_19551,N_18285,N_18551);
xor U19552 (N_19552,N_18594,N_18051);
nor U19553 (N_19553,N_18320,N_18596);
nor U19554 (N_19554,N_18479,N_18235);
nand U19555 (N_19555,N_18516,N_18394);
xor U19556 (N_19556,N_18320,N_18382);
nor U19557 (N_19557,N_18417,N_18137);
or U19558 (N_19558,N_18710,N_18059);
nor U19559 (N_19559,N_17633,N_18149);
xor U19560 (N_19560,N_18248,N_18073);
and U19561 (N_19561,N_18402,N_18556);
and U19562 (N_19562,N_17500,N_18530);
nand U19563 (N_19563,N_18261,N_17587);
and U19564 (N_19564,N_17785,N_17828);
or U19565 (N_19565,N_18452,N_17791);
or U19566 (N_19566,N_18038,N_17927);
xor U19567 (N_19567,N_18672,N_17862);
xnor U19568 (N_19568,N_18088,N_18295);
and U19569 (N_19569,N_18634,N_17538);
or U19570 (N_19570,N_17770,N_18329);
and U19571 (N_19571,N_18474,N_18068);
nor U19572 (N_19572,N_17588,N_17514);
or U19573 (N_19573,N_18499,N_17806);
xor U19574 (N_19574,N_18445,N_17838);
or U19575 (N_19575,N_17879,N_18314);
and U19576 (N_19576,N_18067,N_18594);
nor U19577 (N_19577,N_17792,N_18144);
nand U19578 (N_19578,N_18261,N_18382);
nor U19579 (N_19579,N_18333,N_17954);
nand U19580 (N_19580,N_17648,N_18377);
nor U19581 (N_19581,N_17755,N_18717);
and U19582 (N_19582,N_17643,N_18040);
nand U19583 (N_19583,N_17722,N_17666);
and U19584 (N_19584,N_17677,N_17905);
xnor U19585 (N_19585,N_18691,N_18471);
nand U19586 (N_19586,N_18628,N_18300);
nand U19587 (N_19587,N_18506,N_17623);
nand U19588 (N_19588,N_18741,N_18161);
or U19589 (N_19589,N_17976,N_18035);
nand U19590 (N_19590,N_17590,N_17607);
nand U19591 (N_19591,N_18534,N_18412);
nand U19592 (N_19592,N_18529,N_17537);
xnor U19593 (N_19593,N_17753,N_18040);
nor U19594 (N_19594,N_18231,N_18660);
nor U19595 (N_19595,N_18082,N_18363);
nor U19596 (N_19596,N_18711,N_17659);
xnor U19597 (N_19597,N_17668,N_18218);
or U19598 (N_19598,N_18637,N_17914);
or U19599 (N_19599,N_18485,N_18066);
nand U19600 (N_19600,N_18581,N_18292);
xnor U19601 (N_19601,N_18041,N_17778);
nand U19602 (N_19602,N_17709,N_17664);
xor U19603 (N_19603,N_18028,N_18069);
xor U19604 (N_19604,N_18506,N_17543);
nand U19605 (N_19605,N_18624,N_18026);
nor U19606 (N_19606,N_17937,N_18448);
nor U19607 (N_19607,N_18377,N_18318);
and U19608 (N_19608,N_18296,N_18089);
nor U19609 (N_19609,N_17632,N_18316);
or U19610 (N_19610,N_18368,N_17832);
or U19611 (N_19611,N_18569,N_18336);
nor U19612 (N_19612,N_18460,N_18450);
nand U19613 (N_19613,N_17675,N_17616);
nor U19614 (N_19614,N_18616,N_18378);
nor U19615 (N_19615,N_17589,N_18295);
and U19616 (N_19616,N_18464,N_17933);
and U19617 (N_19617,N_18296,N_18580);
and U19618 (N_19618,N_18289,N_18672);
nand U19619 (N_19619,N_18601,N_17536);
xnor U19620 (N_19620,N_18394,N_17624);
nor U19621 (N_19621,N_18738,N_17808);
nor U19622 (N_19622,N_18489,N_18293);
nor U19623 (N_19623,N_18460,N_17951);
or U19624 (N_19624,N_18371,N_18578);
nor U19625 (N_19625,N_17965,N_17628);
nand U19626 (N_19626,N_17727,N_18202);
or U19627 (N_19627,N_18282,N_18498);
and U19628 (N_19628,N_18465,N_17747);
nand U19629 (N_19629,N_18087,N_17813);
nand U19630 (N_19630,N_18430,N_18534);
nand U19631 (N_19631,N_18473,N_17720);
and U19632 (N_19632,N_17966,N_18579);
or U19633 (N_19633,N_18113,N_18018);
or U19634 (N_19634,N_18440,N_18100);
xor U19635 (N_19635,N_18430,N_18404);
nand U19636 (N_19636,N_18126,N_17638);
nand U19637 (N_19637,N_18331,N_18110);
nor U19638 (N_19638,N_17828,N_18440);
and U19639 (N_19639,N_18604,N_18298);
nor U19640 (N_19640,N_18144,N_18243);
nand U19641 (N_19641,N_18114,N_17814);
xor U19642 (N_19642,N_17819,N_18148);
and U19643 (N_19643,N_18328,N_18232);
and U19644 (N_19644,N_18002,N_17529);
nor U19645 (N_19645,N_17803,N_17509);
xnor U19646 (N_19646,N_18471,N_18267);
or U19647 (N_19647,N_17656,N_18733);
xnor U19648 (N_19648,N_18183,N_18206);
nand U19649 (N_19649,N_18489,N_17661);
nand U19650 (N_19650,N_18609,N_17744);
xor U19651 (N_19651,N_18729,N_18695);
nor U19652 (N_19652,N_18446,N_17655);
xor U19653 (N_19653,N_18358,N_17538);
nor U19654 (N_19654,N_17881,N_18202);
nor U19655 (N_19655,N_18299,N_18108);
nand U19656 (N_19656,N_18619,N_18630);
and U19657 (N_19657,N_17763,N_17995);
nor U19658 (N_19658,N_17882,N_18333);
or U19659 (N_19659,N_18040,N_17624);
nor U19660 (N_19660,N_18255,N_18128);
and U19661 (N_19661,N_18260,N_17752);
and U19662 (N_19662,N_18463,N_17513);
nand U19663 (N_19663,N_18151,N_18305);
and U19664 (N_19664,N_17676,N_18341);
or U19665 (N_19665,N_17677,N_18551);
or U19666 (N_19666,N_18697,N_18025);
and U19667 (N_19667,N_17524,N_17942);
and U19668 (N_19668,N_17705,N_18738);
or U19669 (N_19669,N_18680,N_18291);
nor U19670 (N_19670,N_18212,N_18599);
nor U19671 (N_19671,N_18642,N_17865);
nor U19672 (N_19672,N_18642,N_18382);
and U19673 (N_19673,N_18664,N_18625);
xnor U19674 (N_19674,N_18339,N_18283);
or U19675 (N_19675,N_17854,N_18684);
xor U19676 (N_19676,N_18453,N_18735);
nor U19677 (N_19677,N_18117,N_17802);
xnor U19678 (N_19678,N_18065,N_18580);
or U19679 (N_19679,N_18433,N_17729);
or U19680 (N_19680,N_18435,N_17906);
xor U19681 (N_19681,N_18268,N_18346);
nand U19682 (N_19682,N_18679,N_17719);
and U19683 (N_19683,N_18611,N_17720);
nor U19684 (N_19684,N_17501,N_17780);
xor U19685 (N_19685,N_17533,N_18265);
or U19686 (N_19686,N_18223,N_18266);
and U19687 (N_19687,N_17671,N_18652);
nor U19688 (N_19688,N_18662,N_18075);
or U19689 (N_19689,N_18264,N_18647);
nor U19690 (N_19690,N_17528,N_18520);
xnor U19691 (N_19691,N_18563,N_17920);
or U19692 (N_19692,N_18309,N_17953);
nand U19693 (N_19693,N_17613,N_18196);
nor U19694 (N_19694,N_18380,N_18289);
and U19695 (N_19695,N_17726,N_17504);
xnor U19696 (N_19696,N_17696,N_18466);
and U19697 (N_19697,N_18108,N_18161);
or U19698 (N_19698,N_17935,N_18338);
and U19699 (N_19699,N_17931,N_18337);
nor U19700 (N_19700,N_17559,N_18000);
xnor U19701 (N_19701,N_18301,N_18478);
nand U19702 (N_19702,N_18120,N_18186);
xor U19703 (N_19703,N_18655,N_18747);
xor U19704 (N_19704,N_17863,N_18425);
and U19705 (N_19705,N_17853,N_17919);
or U19706 (N_19706,N_17538,N_17566);
nand U19707 (N_19707,N_18180,N_17906);
and U19708 (N_19708,N_18103,N_17688);
or U19709 (N_19709,N_17564,N_17718);
and U19710 (N_19710,N_17959,N_17727);
nand U19711 (N_19711,N_18058,N_18381);
nand U19712 (N_19712,N_17511,N_17726);
xnor U19713 (N_19713,N_18649,N_17582);
nor U19714 (N_19714,N_17899,N_17952);
nor U19715 (N_19715,N_18647,N_18170);
or U19716 (N_19716,N_18101,N_17943);
or U19717 (N_19717,N_18679,N_17628);
and U19718 (N_19718,N_17915,N_18184);
xnor U19719 (N_19719,N_18298,N_17984);
and U19720 (N_19720,N_17589,N_18279);
or U19721 (N_19721,N_18199,N_17696);
nor U19722 (N_19722,N_17928,N_18057);
or U19723 (N_19723,N_18056,N_17842);
nor U19724 (N_19724,N_18077,N_17990);
nor U19725 (N_19725,N_18067,N_17998);
nand U19726 (N_19726,N_18648,N_17732);
nand U19727 (N_19727,N_18074,N_18419);
nor U19728 (N_19728,N_18216,N_18427);
nand U19729 (N_19729,N_17894,N_17672);
xor U19730 (N_19730,N_17771,N_18713);
and U19731 (N_19731,N_18438,N_18742);
nor U19732 (N_19732,N_17983,N_18692);
and U19733 (N_19733,N_18695,N_17919);
or U19734 (N_19734,N_17999,N_18074);
nor U19735 (N_19735,N_18062,N_18475);
nor U19736 (N_19736,N_18368,N_18113);
or U19737 (N_19737,N_17670,N_18052);
or U19738 (N_19738,N_18699,N_18268);
xor U19739 (N_19739,N_18134,N_18582);
nand U19740 (N_19740,N_17656,N_18170);
nor U19741 (N_19741,N_18289,N_17708);
nand U19742 (N_19742,N_17841,N_18017);
or U19743 (N_19743,N_18398,N_18443);
and U19744 (N_19744,N_17891,N_18554);
xor U19745 (N_19745,N_18279,N_18703);
or U19746 (N_19746,N_17683,N_18310);
nand U19747 (N_19747,N_17984,N_17588);
nor U19748 (N_19748,N_18110,N_17619);
and U19749 (N_19749,N_17584,N_18231);
nor U19750 (N_19750,N_17675,N_18110);
and U19751 (N_19751,N_18317,N_17949);
nand U19752 (N_19752,N_18373,N_18091);
and U19753 (N_19753,N_18435,N_17594);
xnor U19754 (N_19754,N_18138,N_18355);
xor U19755 (N_19755,N_18419,N_17615);
and U19756 (N_19756,N_18676,N_18559);
and U19757 (N_19757,N_18582,N_18192);
nand U19758 (N_19758,N_18075,N_18678);
nand U19759 (N_19759,N_18494,N_18055);
nand U19760 (N_19760,N_18137,N_18632);
xnor U19761 (N_19761,N_18273,N_18153);
xor U19762 (N_19762,N_17639,N_17516);
nor U19763 (N_19763,N_18459,N_18719);
and U19764 (N_19764,N_17696,N_18688);
or U19765 (N_19765,N_18234,N_17508);
and U19766 (N_19766,N_18556,N_17812);
or U19767 (N_19767,N_17727,N_18086);
and U19768 (N_19768,N_17504,N_18575);
or U19769 (N_19769,N_18281,N_18155);
nand U19770 (N_19770,N_17640,N_17910);
and U19771 (N_19771,N_18164,N_17586);
and U19772 (N_19772,N_18694,N_17923);
nor U19773 (N_19773,N_18282,N_17952);
and U19774 (N_19774,N_18366,N_18712);
and U19775 (N_19775,N_17606,N_17894);
nor U19776 (N_19776,N_18308,N_18374);
nand U19777 (N_19777,N_18387,N_17840);
or U19778 (N_19778,N_18620,N_17634);
xnor U19779 (N_19779,N_17570,N_18486);
or U19780 (N_19780,N_17519,N_17919);
xnor U19781 (N_19781,N_18004,N_18657);
nand U19782 (N_19782,N_18540,N_17906);
xnor U19783 (N_19783,N_17594,N_18361);
or U19784 (N_19784,N_18195,N_17638);
nor U19785 (N_19785,N_17804,N_18255);
or U19786 (N_19786,N_18729,N_18589);
nor U19787 (N_19787,N_17702,N_17910);
nor U19788 (N_19788,N_18475,N_18458);
nor U19789 (N_19789,N_18530,N_18250);
nor U19790 (N_19790,N_18358,N_17918);
or U19791 (N_19791,N_18294,N_17756);
nand U19792 (N_19792,N_18040,N_17771);
xnor U19793 (N_19793,N_18544,N_18155);
nor U19794 (N_19794,N_18410,N_17893);
nor U19795 (N_19795,N_18745,N_18609);
nor U19796 (N_19796,N_18489,N_17818);
nand U19797 (N_19797,N_18344,N_17552);
and U19798 (N_19798,N_18478,N_18444);
nor U19799 (N_19799,N_17951,N_17554);
xor U19800 (N_19800,N_17864,N_17700);
xor U19801 (N_19801,N_18002,N_18557);
nand U19802 (N_19802,N_18520,N_18151);
xnor U19803 (N_19803,N_17967,N_18411);
xor U19804 (N_19804,N_18388,N_17699);
xor U19805 (N_19805,N_18088,N_18271);
nor U19806 (N_19806,N_18333,N_18150);
and U19807 (N_19807,N_18151,N_17501);
or U19808 (N_19808,N_18521,N_17725);
or U19809 (N_19809,N_17517,N_18356);
or U19810 (N_19810,N_18358,N_17505);
nand U19811 (N_19811,N_18253,N_18489);
nor U19812 (N_19812,N_18350,N_18042);
nor U19813 (N_19813,N_18065,N_17672);
and U19814 (N_19814,N_17732,N_18596);
or U19815 (N_19815,N_17671,N_18463);
or U19816 (N_19816,N_17728,N_17512);
xnor U19817 (N_19817,N_18347,N_18315);
and U19818 (N_19818,N_17815,N_18340);
nand U19819 (N_19819,N_18364,N_17653);
xor U19820 (N_19820,N_18216,N_18456);
xor U19821 (N_19821,N_18749,N_18365);
or U19822 (N_19822,N_17514,N_18244);
xor U19823 (N_19823,N_18423,N_17764);
nor U19824 (N_19824,N_18679,N_18216);
nor U19825 (N_19825,N_17909,N_17643);
nor U19826 (N_19826,N_18655,N_17602);
or U19827 (N_19827,N_18498,N_18189);
nor U19828 (N_19828,N_18139,N_18215);
or U19829 (N_19829,N_17970,N_17615);
nor U19830 (N_19830,N_18110,N_17701);
xnor U19831 (N_19831,N_17563,N_18108);
nor U19832 (N_19832,N_18501,N_18531);
xor U19833 (N_19833,N_18354,N_18233);
nand U19834 (N_19834,N_18526,N_18167);
or U19835 (N_19835,N_18520,N_17670);
or U19836 (N_19836,N_18458,N_18602);
xnor U19837 (N_19837,N_17820,N_17804);
nand U19838 (N_19838,N_18096,N_17775);
nand U19839 (N_19839,N_17510,N_17926);
nor U19840 (N_19840,N_18010,N_18201);
xor U19841 (N_19841,N_17864,N_17523);
xnor U19842 (N_19842,N_18007,N_17697);
xnor U19843 (N_19843,N_17793,N_18668);
and U19844 (N_19844,N_18700,N_17910);
xnor U19845 (N_19845,N_17743,N_18469);
nand U19846 (N_19846,N_17714,N_18022);
and U19847 (N_19847,N_17735,N_18502);
or U19848 (N_19848,N_18557,N_18301);
xnor U19849 (N_19849,N_17505,N_18499);
and U19850 (N_19850,N_18548,N_17733);
and U19851 (N_19851,N_17745,N_17884);
nand U19852 (N_19852,N_18185,N_18149);
nand U19853 (N_19853,N_18495,N_18290);
nor U19854 (N_19854,N_18205,N_18671);
or U19855 (N_19855,N_17998,N_18026);
and U19856 (N_19856,N_18684,N_17989);
nand U19857 (N_19857,N_17894,N_18743);
nand U19858 (N_19858,N_18067,N_17524);
or U19859 (N_19859,N_17647,N_17919);
xor U19860 (N_19860,N_18657,N_18711);
or U19861 (N_19861,N_17762,N_18240);
and U19862 (N_19862,N_18498,N_18577);
nand U19863 (N_19863,N_18008,N_18047);
nor U19864 (N_19864,N_17875,N_18694);
nand U19865 (N_19865,N_17711,N_17744);
and U19866 (N_19866,N_18697,N_18047);
and U19867 (N_19867,N_17699,N_18270);
nand U19868 (N_19868,N_17595,N_18440);
or U19869 (N_19869,N_18670,N_17624);
nand U19870 (N_19870,N_18545,N_18662);
nand U19871 (N_19871,N_18713,N_18698);
or U19872 (N_19872,N_18288,N_17708);
xor U19873 (N_19873,N_17792,N_17691);
and U19874 (N_19874,N_17758,N_18220);
nand U19875 (N_19875,N_18283,N_17563);
and U19876 (N_19876,N_18126,N_17854);
or U19877 (N_19877,N_18108,N_18107);
or U19878 (N_19878,N_18693,N_18104);
nand U19879 (N_19879,N_18356,N_17988);
or U19880 (N_19880,N_17835,N_18065);
xnor U19881 (N_19881,N_18016,N_17550);
and U19882 (N_19882,N_17721,N_18470);
nor U19883 (N_19883,N_18722,N_18149);
or U19884 (N_19884,N_17580,N_18602);
nand U19885 (N_19885,N_18575,N_18667);
xnor U19886 (N_19886,N_18734,N_18074);
or U19887 (N_19887,N_18533,N_18450);
or U19888 (N_19888,N_17943,N_17574);
nand U19889 (N_19889,N_17719,N_17654);
xor U19890 (N_19890,N_17719,N_18205);
nand U19891 (N_19891,N_18265,N_17885);
nor U19892 (N_19892,N_17872,N_17536);
nand U19893 (N_19893,N_18693,N_18585);
xnor U19894 (N_19894,N_18582,N_17829);
xor U19895 (N_19895,N_17693,N_18339);
or U19896 (N_19896,N_17923,N_17554);
nor U19897 (N_19897,N_18313,N_17819);
or U19898 (N_19898,N_18479,N_18307);
nand U19899 (N_19899,N_18116,N_18699);
xor U19900 (N_19900,N_17985,N_18725);
and U19901 (N_19901,N_18135,N_18472);
or U19902 (N_19902,N_18484,N_18550);
nand U19903 (N_19903,N_18183,N_17507);
nand U19904 (N_19904,N_18532,N_18359);
and U19905 (N_19905,N_17658,N_17948);
nor U19906 (N_19906,N_18252,N_18710);
or U19907 (N_19907,N_17504,N_17593);
or U19908 (N_19908,N_18006,N_18490);
nor U19909 (N_19909,N_18213,N_17877);
and U19910 (N_19910,N_18210,N_18341);
xnor U19911 (N_19911,N_18092,N_18090);
nand U19912 (N_19912,N_18069,N_18643);
or U19913 (N_19913,N_17527,N_18686);
nor U19914 (N_19914,N_18001,N_17821);
xnor U19915 (N_19915,N_17848,N_18605);
nand U19916 (N_19916,N_17930,N_17855);
xor U19917 (N_19917,N_18503,N_17903);
xor U19918 (N_19918,N_18646,N_18063);
nor U19919 (N_19919,N_18599,N_18272);
nor U19920 (N_19920,N_17860,N_18557);
nor U19921 (N_19921,N_18667,N_18229);
and U19922 (N_19922,N_18564,N_17888);
and U19923 (N_19923,N_18507,N_17505);
nand U19924 (N_19924,N_18360,N_17694);
and U19925 (N_19925,N_17878,N_17590);
and U19926 (N_19926,N_18346,N_17880);
and U19927 (N_19927,N_17756,N_17982);
xor U19928 (N_19928,N_18112,N_18358);
xor U19929 (N_19929,N_18074,N_17563);
xnor U19930 (N_19930,N_18225,N_18555);
and U19931 (N_19931,N_18413,N_18608);
or U19932 (N_19932,N_17816,N_18436);
nand U19933 (N_19933,N_18541,N_18177);
nor U19934 (N_19934,N_18084,N_18092);
nand U19935 (N_19935,N_18436,N_17980);
and U19936 (N_19936,N_17918,N_18649);
xnor U19937 (N_19937,N_17950,N_18551);
or U19938 (N_19938,N_17961,N_17755);
and U19939 (N_19939,N_18612,N_18715);
and U19940 (N_19940,N_18312,N_17727);
nand U19941 (N_19941,N_18716,N_18165);
or U19942 (N_19942,N_17812,N_18041);
xor U19943 (N_19943,N_18016,N_18473);
nand U19944 (N_19944,N_18364,N_18552);
or U19945 (N_19945,N_18463,N_17878);
and U19946 (N_19946,N_18588,N_17669);
xnor U19947 (N_19947,N_18624,N_18434);
or U19948 (N_19948,N_18270,N_18402);
xor U19949 (N_19949,N_17822,N_18315);
nor U19950 (N_19950,N_18411,N_18283);
nor U19951 (N_19951,N_18003,N_17760);
and U19952 (N_19952,N_18344,N_18079);
nand U19953 (N_19953,N_18089,N_18489);
or U19954 (N_19954,N_18727,N_17794);
or U19955 (N_19955,N_18116,N_18202);
nor U19956 (N_19956,N_18415,N_18066);
and U19957 (N_19957,N_17762,N_17588);
and U19958 (N_19958,N_18241,N_17958);
xor U19959 (N_19959,N_17878,N_17772);
xnor U19960 (N_19960,N_18379,N_18098);
xor U19961 (N_19961,N_17513,N_18661);
nor U19962 (N_19962,N_18638,N_18687);
or U19963 (N_19963,N_18091,N_18186);
and U19964 (N_19964,N_18539,N_18572);
and U19965 (N_19965,N_17957,N_17580);
and U19966 (N_19966,N_18468,N_17703);
nand U19967 (N_19967,N_17741,N_18705);
nand U19968 (N_19968,N_17615,N_17529);
nand U19969 (N_19969,N_18738,N_17873);
or U19970 (N_19970,N_18255,N_18448);
or U19971 (N_19971,N_18561,N_17661);
and U19972 (N_19972,N_18084,N_18030);
nor U19973 (N_19973,N_18255,N_18652);
and U19974 (N_19974,N_18369,N_18668);
or U19975 (N_19975,N_17806,N_17719);
and U19976 (N_19976,N_18444,N_18228);
nor U19977 (N_19977,N_17997,N_18222);
and U19978 (N_19978,N_18651,N_17609);
xor U19979 (N_19979,N_18092,N_18679);
nor U19980 (N_19980,N_17581,N_18023);
and U19981 (N_19981,N_18700,N_17974);
and U19982 (N_19982,N_17932,N_18368);
nand U19983 (N_19983,N_18240,N_17810);
nand U19984 (N_19984,N_18510,N_17937);
and U19985 (N_19985,N_18435,N_17900);
nor U19986 (N_19986,N_17658,N_17779);
or U19987 (N_19987,N_18056,N_18737);
nand U19988 (N_19988,N_18359,N_18099);
and U19989 (N_19989,N_18594,N_18439);
xnor U19990 (N_19990,N_17857,N_18132);
and U19991 (N_19991,N_17910,N_17786);
nand U19992 (N_19992,N_18553,N_18486);
xor U19993 (N_19993,N_17818,N_18051);
or U19994 (N_19994,N_18067,N_17569);
xnor U19995 (N_19995,N_18099,N_17956);
and U19996 (N_19996,N_17694,N_18692);
nor U19997 (N_19997,N_18553,N_17808);
or U19998 (N_19998,N_17545,N_18365);
nor U19999 (N_19999,N_17688,N_18658);
or U20000 (N_20000,N_19733,N_19551);
nor U20001 (N_20001,N_19252,N_19529);
nor U20002 (N_20002,N_19774,N_19548);
nor U20003 (N_20003,N_19656,N_19520);
nor U20004 (N_20004,N_19176,N_19228);
nor U20005 (N_20005,N_19293,N_19157);
nor U20006 (N_20006,N_18989,N_19368);
xnor U20007 (N_20007,N_19862,N_19486);
nor U20008 (N_20008,N_18941,N_19756);
and U20009 (N_20009,N_19268,N_19650);
nor U20010 (N_20010,N_19623,N_19246);
nand U20011 (N_20011,N_19519,N_19029);
xnor U20012 (N_20012,N_19309,N_19041);
nor U20013 (N_20013,N_19023,N_19513);
or U20014 (N_20014,N_19026,N_18971);
nand U20015 (N_20015,N_19682,N_19393);
nor U20016 (N_20016,N_18902,N_18822);
nand U20017 (N_20017,N_19641,N_19159);
or U20018 (N_20018,N_19104,N_19578);
nor U20019 (N_20019,N_19540,N_19069);
xor U20020 (N_20020,N_18806,N_19407);
nand U20021 (N_20021,N_19345,N_19531);
nor U20022 (N_20022,N_19165,N_18825);
or U20023 (N_20023,N_19585,N_19688);
xor U20024 (N_20024,N_18947,N_19201);
xor U20025 (N_20025,N_19598,N_18762);
xor U20026 (N_20026,N_19828,N_18828);
nor U20027 (N_20027,N_19395,N_19544);
nand U20028 (N_20028,N_19036,N_19621);
and U20029 (N_20029,N_19112,N_19214);
nand U20030 (N_20030,N_19587,N_19824);
and U20031 (N_20031,N_19062,N_19166);
xnor U20032 (N_20032,N_19975,N_19329);
xnor U20033 (N_20033,N_19132,N_19213);
nand U20034 (N_20034,N_19199,N_19851);
or U20035 (N_20035,N_18854,N_19521);
or U20036 (N_20036,N_19010,N_19786);
nand U20037 (N_20037,N_19586,N_19194);
or U20038 (N_20038,N_18830,N_19234);
or U20039 (N_20039,N_18942,N_19045);
or U20040 (N_20040,N_19924,N_19633);
and U20041 (N_20041,N_19775,N_19326);
xor U20042 (N_20042,N_19319,N_19356);
nand U20043 (N_20043,N_18761,N_19505);
nand U20044 (N_20044,N_19861,N_19180);
or U20045 (N_20045,N_19766,N_19831);
xor U20046 (N_20046,N_19111,N_19574);
or U20047 (N_20047,N_19514,N_19547);
xor U20048 (N_20048,N_19316,N_19328);
nor U20049 (N_20049,N_19880,N_18995);
xnor U20050 (N_20050,N_19868,N_18945);
or U20051 (N_20051,N_19225,N_19966);
nand U20052 (N_20052,N_18931,N_19860);
nor U20053 (N_20053,N_18804,N_19624);
or U20054 (N_20054,N_19318,N_18798);
and U20055 (N_20055,N_19003,N_19264);
and U20056 (N_20056,N_19764,N_19058);
or U20057 (N_20057,N_18789,N_19818);
nor U20058 (N_20058,N_19147,N_19219);
nor U20059 (N_20059,N_19464,N_19954);
xor U20060 (N_20060,N_19651,N_19631);
nand U20061 (N_20061,N_19281,N_19289);
or U20062 (N_20062,N_19363,N_18969);
nand U20063 (N_20063,N_18927,N_18937);
nand U20064 (N_20064,N_19899,N_19353);
nor U20065 (N_20065,N_19497,N_19394);
xnor U20066 (N_20066,N_19116,N_18778);
and U20067 (N_20067,N_19526,N_19592);
and U20068 (N_20068,N_19992,N_19681);
or U20069 (N_20069,N_19857,N_19156);
and U20070 (N_20070,N_19061,N_19875);
nand U20071 (N_20071,N_19536,N_19099);
or U20072 (N_20072,N_19122,N_19427);
and U20073 (N_20073,N_19605,N_19424);
nor U20074 (N_20074,N_19702,N_19898);
xor U20075 (N_20075,N_19034,N_19739);
or U20076 (N_20076,N_19064,N_19606);
nand U20077 (N_20077,N_19794,N_19988);
and U20078 (N_20078,N_19654,N_19782);
or U20079 (N_20079,N_19414,N_19662);
or U20080 (N_20080,N_19713,N_19488);
or U20081 (N_20081,N_18881,N_18901);
nor U20082 (N_20082,N_19802,N_18752);
nand U20083 (N_20083,N_19995,N_19622);
or U20084 (N_20084,N_19974,N_19172);
and U20085 (N_20085,N_19640,N_19461);
xor U20086 (N_20086,N_19173,N_18932);
xor U20087 (N_20087,N_18985,N_18811);
nand U20088 (N_20088,N_19181,N_19660);
nor U20089 (N_20089,N_19618,N_19434);
xor U20090 (N_20090,N_19355,N_19302);
and U20091 (N_20091,N_18990,N_19404);
or U20092 (N_20092,N_19803,N_19384);
xor U20093 (N_20093,N_19002,N_19576);
nor U20094 (N_20094,N_18832,N_18867);
nor U20095 (N_20095,N_19174,N_19085);
and U20096 (N_20096,N_19680,N_19674);
and U20097 (N_20097,N_19842,N_19426);
nand U20098 (N_20098,N_19479,N_19960);
xor U20099 (N_20099,N_19443,N_19380);
nor U20100 (N_20100,N_18781,N_19789);
xor U20101 (N_20101,N_19007,N_19179);
nor U20102 (N_20102,N_19557,N_19757);
xnor U20103 (N_20103,N_19823,N_19770);
xnor U20104 (N_20104,N_18754,N_18810);
or U20105 (N_20105,N_19241,N_19535);
or U20106 (N_20106,N_19858,N_19288);
nand U20107 (N_20107,N_19878,N_19236);
nand U20108 (N_20108,N_18772,N_19202);
and U20109 (N_20109,N_18793,N_19152);
and U20110 (N_20110,N_19925,N_18908);
xnor U20111 (N_20111,N_19990,N_19311);
and U20112 (N_20112,N_19447,N_19616);
xnor U20113 (N_20113,N_19939,N_19611);
nand U20114 (N_20114,N_19726,N_18835);
or U20115 (N_20115,N_19245,N_19170);
xnor U20116 (N_20116,N_18952,N_19080);
nor U20117 (N_20117,N_19283,N_18776);
or U20118 (N_20118,N_19324,N_19107);
xor U20119 (N_20119,N_18999,N_19977);
and U20120 (N_20120,N_19303,N_18758);
nand U20121 (N_20121,N_18957,N_19599);
xor U20122 (N_20122,N_19204,N_19678);
xor U20123 (N_20123,N_19383,N_19541);
xor U20124 (N_20124,N_19836,N_18919);
nand U20125 (N_20125,N_19435,N_19337);
nor U20126 (N_20126,N_19564,N_19422);
xnor U20127 (N_20127,N_18784,N_19504);
xor U20128 (N_20128,N_19182,N_19719);
or U20129 (N_20129,N_19523,N_19837);
nor U20130 (N_20130,N_19418,N_19556);
nand U20131 (N_20131,N_19666,N_19187);
or U20132 (N_20132,N_19809,N_19402);
nor U20133 (N_20133,N_18975,N_19387);
nand U20134 (N_20134,N_18950,N_19591);
and U20135 (N_20135,N_19723,N_18777);
and U20136 (N_20136,N_19516,N_19015);
and U20137 (N_20137,N_19922,N_19121);
or U20138 (N_20138,N_19391,N_19762);
nor U20139 (N_20139,N_19101,N_19820);
xor U20140 (N_20140,N_19866,N_19817);
or U20141 (N_20141,N_18893,N_19243);
or U20142 (N_20142,N_19889,N_19330);
nand U20143 (N_20143,N_18792,N_19450);
and U20144 (N_20144,N_19462,N_19495);
xnor U20145 (N_20145,N_18805,N_18800);
nand U20146 (N_20146,N_19184,N_19158);
or U20147 (N_20147,N_19411,N_19758);
nor U20148 (N_20148,N_19962,N_19049);
xnor U20149 (N_20149,N_19949,N_19232);
and U20150 (N_20150,N_19271,N_18954);
xor U20151 (N_20151,N_19507,N_19763);
nand U20152 (N_20152,N_19509,N_19783);
nor U20153 (N_20153,N_19886,N_19242);
or U20154 (N_20154,N_18883,N_19291);
or U20155 (N_20155,N_19115,N_19050);
or U20156 (N_20156,N_19732,N_19684);
and U20157 (N_20157,N_19095,N_18868);
nor U20158 (N_20158,N_18786,N_19437);
xnor U20159 (N_20159,N_19927,N_19475);
and U20160 (N_20160,N_19200,N_18944);
nand U20161 (N_20161,N_19872,N_18885);
xor U20162 (N_20162,N_19139,N_19942);
or U20163 (N_20163,N_18785,N_18986);
xnor U20164 (N_20164,N_19257,N_19738);
or U20165 (N_20165,N_19814,N_18850);
or U20166 (N_20166,N_18926,N_19700);
and U20167 (N_20167,N_19221,N_18824);
xor U20168 (N_20168,N_19140,N_19338);
or U20169 (N_20169,N_18795,N_19073);
xnor U20170 (N_20170,N_19423,N_18879);
or U20171 (N_20171,N_19558,N_18962);
nand U20172 (N_20172,N_19928,N_19039);
xor U20173 (N_20173,N_19077,N_19038);
nor U20174 (N_20174,N_19968,N_19908);
nand U20175 (N_20175,N_19150,N_19492);
xor U20176 (N_20176,N_19776,N_19994);
nor U20177 (N_20177,N_19750,N_19575);
or U20178 (N_20178,N_19580,N_18951);
and U20179 (N_20179,N_19594,N_19349);
nand U20180 (N_20180,N_19206,N_18787);
nand U20181 (N_20181,N_19525,N_18922);
xnor U20182 (N_20182,N_18924,N_19390);
nor U20183 (N_20183,N_19619,N_19458);
xnor U20184 (N_20184,N_18973,N_19562);
or U20185 (N_20185,N_19494,N_18848);
nor U20186 (N_20186,N_19067,N_19795);
and U20187 (N_20187,N_19377,N_19445);
xnor U20188 (N_20188,N_19696,N_19694);
and U20189 (N_20189,N_19300,N_19113);
or U20190 (N_20190,N_19256,N_19884);
and U20191 (N_20191,N_19093,N_19471);
or U20192 (N_20192,N_19685,N_19322);
nand U20193 (N_20193,N_19192,N_19630);
nor U20194 (N_20194,N_18856,N_19855);
nor U20195 (N_20195,N_19028,N_18773);
xnor U20196 (N_20196,N_19873,N_19483);
and U20197 (N_20197,N_19946,N_18880);
or U20198 (N_20198,N_19568,N_19597);
nor U20199 (N_20199,N_19210,N_19369);
nor U20200 (N_20200,N_19907,N_19561);
nor U20201 (N_20201,N_18866,N_19129);
and U20202 (N_20202,N_19911,N_19930);
and U20203 (N_20203,N_19603,N_19935);
and U20204 (N_20204,N_18812,N_19790);
or U20205 (N_20205,N_19500,N_19084);
or U20206 (N_20206,N_18750,N_19255);
nand U20207 (N_20207,N_18788,N_19545);
nand U20208 (N_20208,N_19822,N_19405);
nor U20209 (N_20209,N_19844,N_19323);
or U20210 (N_20210,N_19304,N_18888);
or U20211 (N_20211,N_18871,N_18935);
or U20212 (N_20212,N_18807,N_18863);
xnor U20213 (N_20213,N_19358,N_19767);
xnor U20214 (N_20214,N_19686,N_18840);
or U20215 (N_20215,N_18940,N_19070);
nor U20216 (N_20216,N_19542,N_19496);
nor U20217 (N_20217,N_19499,N_18790);
or U20218 (N_20218,N_19183,N_19826);
or U20219 (N_20219,N_18974,N_19971);
and U20220 (N_20220,N_19819,N_19013);
nand U20221 (N_20221,N_18909,N_19801);
xor U20222 (N_20222,N_19493,N_19989);
or U20223 (N_20223,N_19382,N_19560);
nand U20224 (N_20224,N_18889,N_19452);
xor U20225 (N_20225,N_19498,N_19639);
or U20226 (N_20226,N_19903,N_19792);
and U20227 (N_20227,N_19117,N_18803);
xnor U20228 (N_20228,N_19885,N_19065);
or U20229 (N_20229,N_19951,N_19731);
nand U20230 (N_20230,N_19251,N_18873);
nand U20231 (N_20231,N_19127,N_18977);
nor U20232 (N_20232,N_19563,N_18799);
nand U20233 (N_20233,N_19196,N_19325);
and U20234 (N_20234,N_19695,N_19279);
or U20235 (N_20235,N_19403,N_19066);
nand U20236 (N_20236,N_19307,N_19583);
xnor U20237 (N_20237,N_19584,N_19871);
or U20238 (N_20238,N_19835,N_19511);
or U20239 (N_20239,N_19613,N_18833);
xnor U20240 (N_20240,N_19808,N_19354);
and U20241 (N_20241,N_19569,N_19800);
nand U20242 (N_20242,N_19490,N_19918);
xnor U20243 (N_20243,N_18972,N_19295);
xnor U20244 (N_20244,N_18915,N_19033);
nor U20245 (N_20245,N_19420,N_19047);
or U20246 (N_20246,N_18916,N_19915);
and U20247 (N_20247,N_19301,N_18782);
nor U20248 (N_20248,N_19779,N_18899);
and U20249 (N_20249,N_19687,N_19463);
and U20250 (N_20250,N_19429,N_19299);
and U20251 (N_20251,N_19009,N_18917);
or U20252 (N_20252,N_19321,N_19430);
and U20253 (N_20253,N_19408,N_18763);
and U20254 (N_20254,N_19691,N_19102);
nand U20255 (N_20255,N_19059,N_19667);
and U20256 (N_20256,N_19195,N_19566);
nor U20257 (N_20257,N_19890,N_19484);
or U20258 (N_20258,N_19290,N_19254);
and U20259 (N_20259,N_19863,N_19530);
nor U20260 (N_20260,N_19491,N_19538);
and U20261 (N_20261,N_19969,N_19190);
and U20262 (N_20262,N_19707,N_19317);
and U20263 (N_20263,N_19796,N_19852);
nand U20264 (N_20264,N_19850,N_18780);
nand U20265 (N_20265,N_19142,N_19673);
or U20266 (N_20266,N_19669,N_19769);
nor U20267 (N_20267,N_19216,N_18929);
nand U20268 (N_20268,N_18898,N_19001);
and U20269 (N_20269,N_19999,N_19386);
nor U20270 (N_20270,N_19442,N_19751);
xor U20271 (N_20271,N_19063,N_19957);
nand U20272 (N_20272,N_19344,N_19357);
nand U20273 (N_20273,N_19436,N_18823);
or U20274 (N_20274,N_19433,N_19428);
xnor U20275 (N_20275,N_18934,N_18755);
xor U20276 (N_20276,N_18914,N_19864);
or U20277 (N_20277,N_19169,N_19269);
nor U20278 (N_20278,N_19672,N_19222);
xnor U20279 (N_20279,N_19698,N_19054);
nor U20280 (N_20280,N_19474,N_19397);
nand U20281 (N_20281,N_19658,N_18783);
xor U20282 (N_20282,N_19848,N_19665);
or U20283 (N_20283,N_18984,N_19993);
and U20284 (N_20284,N_18872,N_18837);
xnor U20285 (N_20285,N_19090,N_19853);
xnor U20286 (N_20286,N_19017,N_19760);
and U20287 (N_20287,N_18939,N_18894);
and U20288 (N_20288,N_19781,N_19748);
nand U20289 (N_20289,N_19217,N_19743);
xnor U20290 (N_20290,N_19805,N_19634);
or U20291 (N_20291,N_18831,N_19921);
or U20292 (N_20292,N_19668,N_19735);
or U20293 (N_20293,N_19936,N_19198);
and U20294 (N_20294,N_19472,N_19653);
and U20295 (N_20295,N_19040,N_19730);
nor U20296 (N_20296,N_19503,N_19056);
and U20297 (N_20297,N_19203,N_19788);
or U20298 (N_20298,N_19032,N_19043);
and U20299 (N_20299,N_18933,N_18904);
nor U20300 (N_20300,N_19105,N_19454);
nand U20301 (N_20301,N_19375,N_19266);
nor U20302 (N_20302,N_19137,N_19938);
nor U20303 (N_20303,N_19806,N_18991);
nor U20304 (N_20304,N_19725,N_19421);
nor U20305 (N_20305,N_19340,N_19609);
nand U20306 (N_20306,N_18895,N_18882);
xor U20307 (N_20307,N_19883,N_19759);
xor U20308 (N_20308,N_18928,N_18876);
and U20309 (N_20309,N_18820,N_19487);
nand U20310 (N_20310,N_19876,N_19468);
nor U20311 (N_20311,N_19125,N_19027);
nor U20312 (N_20312,N_19670,N_19867);
or U20313 (N_20313,N_19339,N_19554);
xnor U20314 (N_20314,N_19991,N_19088);
and U20315 (N_20315,N_19952,N_19648);
nand U20316 (N_20316,N_19742,N_19896);
and U20317 (N_20317,N_19292,N_19131);
xor U20318 (N_20318,N_18896,N_19089);
or U20319 (N_20319,N_19708,N_19714);
xor U20320 (N_20320,N_19917,N_18836);
nand U20321 (N_20321,N_19679,N_18816);
xnor U20322 (N_20322,N_18955,N_19467);
nor U20323 (N_20323,N_19919,N_19331);
nand U20324 (N_20324,N_19997,N_19155);
and U20325 (N_20325,N_19970,N_18918);
or U20326 (N_20326,N_19025,N_19508);
and U20327 (N_20327,N_19197,N_18925);
and U20328 (N_20328,N_19109,N_19825);
or U20329 (N_20329,N_19754,N_19133);
nor U20330 (N_20330,N_19297,N_19715);
or U20331 (N_20331,N_18870,N_18855);
nor U20332 (N_20332,N_18923,N_19956);
nand U20333 (N_20333,N_19235,N_19167);
or U20334 (N_20334,N_18801,N_18981);
or U20335 (N_20335,N_19753,N_19106);
nand U20336 (N_20336,N_19626,N_19947);
xor U20337 (N_20337,N_19144,N_19108);
and U20338 (N_20338,N_19787,N_19914);
nand U20339 (N_20339,N_18886,N_19539);
nor U20340 (N_20340,N_19410,N_19171);
xor U20341 (N_20341,N_19079,N_19466);
or U20342 (N_20342,N_19231,N_18980);
xor U20343 (N_20343,N_19186,N_19632);
and U20344 (N_20344,N_19449,N_19870);
and U20345 (N_20345,N_19877,N_19312);
nand U20346 (N_20346,N_18966,N_19193);
xnor U20347 (N_20347,N_19798,N_19335);
and U20348 (N_20348,N_19777,N_19706);
xnor U20349 (N_20349,N_19388,N_19126);
or U20350 (N_20350,N_19734,N_19572);
nor U20351 (N_20351,N_19986,N_19900);
nor U20352 (N_20352,N_19559,N_19920);
and U20353 (N_20353,N_19829,N_19267);
nor U20354 (N_20354,N_19145,N_19072);
nand U20355 (N_20355,N_19978,N_19985);
xor U20356 (N_20356,N_19270,N_19346);
or U20357 (N_20357,N_18938,N_19350);
nor U20358 (N_20358,N_18967,N_19772);
or U20359 (N_20359,N_18757,N_19711);
and U20360 (N_20360,N_19655,N_19854);
nand U20361 (N_20361,N_19097,N_19249);
nor U20362 (N_20362,N_19676,N_19315);
nor U20363 (N_20363,N_19083,N_19506);
xnor U20364 (N_20364,N_19976,N_19982);
nor U20365 (N_20365,N_19151,N_19019);
nor U20366 (N_20366,N_19298,N_18844);
and U20367 (N_20367,N_19261,N_19160);
xnor U20368 (N_20368,N_19811,N_19549);
nor U20369 (N_20369,N_19348,N_18797);
xor U20370 (N_20370,N_19501,N_18992);
nand U20371 (N_20371,N_19469,N_18849);
xor U20372 (N_20372,N_19933,N_19894);
nand U20373 (N_20373,N_19524,N_19987);
xnor U20374 (N_20374,N_19590,N_19943);
xor U20375 (N_20375,N_19087,N_19478);
nor U20376 (N_20376,N_19163,N_19413);
nor U20377 (N_20377,N_19909,N_18808);
and U20378 (N_20378,N_19815,N_19887);
or U20379 (N_20379,N_19205,N_19177);
nand U20380 (N_20380,N_19916,N_19663);
nand U20381 (N_20381,N_19923,N_18948);
xor U20382 (N_20382,N_19709,N_18875);
or U20383 (N_20383,N_19000,N_18907);
nand U20384 (N_20384,N_19593,N_19849);
nand U20385 (N_20385,N_18892,N_18826);
and U20386 (N_20386,N_19114,N_19262);
or U20387 (N_20387,N_19148,N_18983);
or U20388 (N_20388,N_19717,N_19627);
nand U20389 (N_20389,N_19533,N_19233);
xnor U20390 (N_20390,N_19373,N_19517);
xor U20391 (N_20391,N_19720,N_19929);
or U20392 (N_20392,N_19865,N_19342);
or U20393 (N_20393,N_19162,N_19642);
xor U20394 (N_20394,N_19961,N_19212);
xnor U20395 (N_20395,N_19124,N_19489);
nor U20396 (N_20396,N_19588,N_19444);
or U20397 (N_20397,N_18769,N_19473);
or U20398 (N_20398,N_19021,N_19341);
and U20399 (N_20399,N_19671,N_19308);
and U20400 (N_20400,N_19459,N_19998);
nor U20401 (N_20401,N_19367,N_19372);
xor U20402 (N_20402,N_19737,N_19074);
nor U20403 (N_20403,N_19768,N_19168);
or U20404 (N_20404,N_19438,N_19522);
nand U20405 (N_20405,N_19343,N_18943);
nand U20406 (N_20406,N_18903,N_19608);
or U20407 (N_20407,N_19582,N_18900);
nor U20408 (N_20408,N_18920,N_19629);
xor U20409 (N_20409,N_19661,N_19869);
or U20410 (N_20410,N_19830,N_19191);
nand U20411 (N_20411,N_19275,N_18994);
and U20412 (N_20412,N_19272,N_19096);
nand U20413 (N_20413,N_19973,N_18987);
and U20414 (N_20414,N_19965,N_19237);
and U20415 (N_20415,N_19161,N_19773);
nor U20416 (N_20416,N_19981,N_19637);
and U20417 (N_20417,N_19881,N_18965);
xor U20418 (N_20418,N_18764,N_18959);
or U20419 (N_20419,N_19123,N_19718);
nand U20420 (N_20420,N_19224,N_19534);
and U20421 (N_20421,N_19018,N_19244);
xor U20422 (N_20422,N_19510,N_19389);
or U20423 (N_20423,N_18964,N_19780);
or U20424 (N_20424,N_19024,N_19385);
and U20425 (N_20425,N_18869,N_19457);
and U20426 (N_20426,N_19797,N_19845);
nor U20427 (N_20427,N_19327,N_19274);
xor U20428 (N_20428,N_18897,N_19625);
or U20429 (N_20429,N_19657,N_19265);
and U20430 (N_20430,N_18963,N_18768);
nor U20431 (N_20431,N_19604,N_19595);
and U20432 (N_20432,N_19379,N_18794);
and U20433 (N_20433,N_19940,N_19071);
or U20434 (N_20434,N_19476,N_18775);
or U20435 (N_20435,N_19832,N_19644);
nand U20436 (N_20436,N_19567,N_19736);
and U20437 (N_20437,N_19953,N_18821);
or U20438 (N_20438,N_19360,N_19481);
and U20439 (N_20439,N_19636,N_19602);
nor U20440 (N_20440,N_19659,N_19398);
xnor U20441 (N_20441,N_18843,N_19004);
or U20442 (N_20442,N_19164,N_19596);
and U20443 (N_20443,N_19897,N_19258);
nand U20444 (N_20444,N_19314,N_19370);
nor U20445 (N_20445,N_18953,N_19189);
or U20446 (N_20446,N_18911,N_19838);
nand U20447 (N_20447,N_18771,N_19502);
xor U20448 (N_20448,N_19276,N_19705);
xnor U20449 (N_20449,N_19581,N_19784);
xnor U20450 (N_20450,N_19532,N_19745);
nor U20451 (N_20451,N_19752,N_19810);
and U20452 (N_20452,N_19416,N_19693);
nand U20453 (N_20453,N_19146,N_19904);
and U20454 (N_20454,N_19692,N_19550);
and U20455 (N_20455,N_19901,N_18910);
nand U20456 (N_20456,N_18842,N_19816);
xnor U20457 (N_20457,N_19950,N_19841);
and U20458 (N_20458,N_19888,N_19135);
or U20459 (N_20459,N_19218,N_19984);
nor U20460 (N_20460,N_19701,N_19294);
xor U20461 (N_20461,N_19729,N_18988);
and U20462 (N_20462,N_18853,N_19926);
or U20463 (N_20463,N_18766,N_19359);
nand U20464 (N_20464,N_18814,N_19892);
and U20465 (N_20465,N_19675,N_19856);
nor U20466 (N_20466,N_18813,N_18958);
xor U20467 (N_20467,N_19432,N_18834);
or U20468 (N_20468,N_19130,N_19746);
nor U20469 (N_20469,N_19963,N_19724);
xnor U20470 (N_20470,N_19075,N_19906);
xnor U20471 (N_20471,N_19376,N_19647);
and U20472 (N_20472,N_19515,N_19215);
nor U20473 (N_20473,N_19552,N_18852);
nor U20474 (N_20474,N_18860,N_19366);
nand U20475 (N_20475,N_19138,N_18993);
xor U20476 (N_20476,N_19728,N_18845);
nand U20477 (N_20477,N_18819,N_19485);
or U20478 (N_20478,N_19527,N_19250);
nor U20479 (N_20479,N_19282,N_19804);
nand U20480 (N_20480,N_18751,N_19082);
and U20481 (N_20481,N_19570,N_18912);
nor U20482 (N_20482,N_19807,N_19118);
and U20483 (N_20483,N_18979,N_19477);
and U20484 (N_20484,N_19638,N_19967);
nor U20485 (N_20485,N_18818,N_19110);
or U20486 (N_20486,N_18851,N_19843);
xnor U20487 (N_20487,N_19690,N_19260);
nor U20488 (N_20488,N_19296,N_18846);
and U20489 (N_20489,N_19931,N_19401);
xor U20490 (N_20490,N_18815,N_19347);
and U20491 (N_20491,N_19100,N_18857);
and U20492 (N_20492,N_19902,N_19365);
nor U20493 (N_20493,N_19175,N_19239);
nor U20494 (N_20494,N_19827,N_19601);
xor U20495 (N_20495,N_19284,N_19646);
and U20496 (N_20496,N_19577,N_19078);
nor U20497 (N_20497,N_19381,N_19400);
xor U20498 (N_20498,N_18779,N_18791);
or U20499 (N_20499,N_19081,N_19912);
and U20500 (N_20500,N_19419,N_19703);
xor U20501 (N_20501,N_19141,N_19006);
nor U20502 (N_20502,N_19277,N_19617);
nand U20503 (N_20503,N_19154,N_19937);
and U20504 (N_20504,N_18829,N_19362);
nor U20505 (N_20505,N_19310,N_19910);
or U20506 (N_20506,N_18817,N_19482);
nand U20507 (N_20507,N_19229,N_19451);
nand U20508 (N_20508,N_19313,N_19697);
and U20509 (N_20509,N_19406,N_19364);
xor U20510 (N_20510,N_19710,N_19247);
nand U20511 (N_20511,N_19415,N_18753);
xnor U20512 (N_20512,N_19834,N_19378);
xor U20513 (N_20513,N_19227,N_19614);
nor U20514 (N_20514,N_19399,N_19334);
and U20515 (N_20515,N_18838,N_19944);
xnor U20516 (N_20516,N_18774,N_19374);
and U20517 (N_20517,N_19188,N_18968);
nor U20518 (N_20518,N_19749,N_19068);
or U20519 (N_20519,N_19840,N_19208);
xor U20520 (N_20520,N_19812,N_19448);
nor U20521 (N_20521,N_19882,N_19470);
or U20522 (N_20522,N_19980,N_19716);
and U20523 (N_20523,N_19280,N_19051);
nand U20524 (N_20524,N_19833,N_19076);
nor U20525 (N_20525,N_18839,N_19689);
nor U20526 (N_20526,N_18890,N_19417);
nand U20527 (N_20527,N_19913,N_19799);
nor U20528 (N_20528,N_19546,N_19821);
nor U20529 (N_20529,N_19439,N_19628);
and U20530 (N_20530,N_19286,N_19453);
and U20531 (N_20531,N_19057,N_19553);
and U20532 (N_20532,N_19958,N_19371);
nor U20533 (N_20533,N_18865,N_19425);
xnor U20534 (N_20534,N_19053,N_19959);
or U20535 (N_20535,N_19465,N_19253);
or U20536 (N_20536,N_19149,N_18976);
nand U20537 (N_20537,N_19945,N_19761);
or U20538 (N_20538,N_19652,N_19305);
nand U20539 (N_20539,N_19456,N_19008);
xor U20540 (N_20540,N_18891,N_18913);
xnor U20541 (N_20541,N_19320,N_19412);
or U20542 (N_20542,N_19683,N_19979);
nand U20543 (N_20543,N_19747,N_18946);
xnor U20544 (N_20544,N_18997,N_19278);
or U20545 (N_20545,N_19446,N_18767);
and U20546 (N_20546,N_18921,N_19612);
and U20547 (N_20547,N_19791,N_19589);
nor U20548 (N_20548,N_18996,N_18756);
xnor U20549 (N_20549,N_18827,N_19934);
nand U20550 (N_20550,N_19263,N_19094);
and U20551 (N_20551,N_19226,N_19248);
and U20552 (N_20552,N_18859,N_19120);
and U20553 (N_20553,N_19932,N_18878);
and U20554 (N_20554,N_18858,N_19664);
and U20555 (N_20555,N_19610,N_18861);
xnor U20556 (N_20556,N_19528,N_19891);
nor U20557 (N_20557,N_19793,N_19895);
and U20558 (N_20558,N_19238,N_19441);
or U20559 (N_20559,N_19431,N_19012);
nor U20560 (N_20560,N_18862,N_19143);
or U20561 (N_20561,N_19352,N_18877);
or U20562 (N_20562,N_19643,N_19119);
nor U20563 (N_20563,N_19955,N_19392);
xnor U20564 (N_20564,N_19153,N_18956);
nand U20565 (N_20565,N_19874,N_19207);
xnor U20566 (N_20566,N_19512,N_19092);
and U20567 (N_20567,N_19351,N_19361);
nor U20568 (N_20568,N_19839,N_18847);
nor U20569 (N_20569,N_19211,N_18949);
nor U20570 (N_20570,N_19016,N_19048);
nor U20571 (N_20571,N_19741,N_18802);
and U20572 (N_20572,N_18930,N_19042);
or U20573 (N_20573,N_19046,N_18905);
xor U20574 (N_20574,N_19103,N_19571);
or U20575 (N_20575,N_19785,N_18884);
nor U20576 (N_20576,N_19230,N_19455);
and U20577 (N_20577,N_19722,N_18936);
or U20578 (N_20578,N_19905,N_19771);
xor U20579 (N_20579,N_19091,N_18961);
nand U20580 (N_20580,N_19964,N_19543);
nor U20581 (N_20581,N_19677,N_18887);
and U20582 (N_20582,N_19755,N_19098);
nor U20583 (N_20583,N_18765,N_19055);
or U20584 (N_20584,N_19060,N_19333);
xnor U20585 (N_20585,N_19336,N_19178);
and U20586 (N_20586,N_19712,N_18759);
or U20587 (N_20587,N_18982,N_19699);
or U20588 (N_20588,N_19273,N_18906);
and U20589 (N_20589,N_18809,N_19136);
nor U20590 (N_20590,N_18960,N_19537);
xnor U20591 (N_20591,N_19555,N_18841);
or U20592 (N_20592,N_19014,N_19020);
nand U20593 (N_20593,N_19600,N_18998);
nor U20594 (N_20594,N_19579,N_19704);
or U20595 (N_20595,N_19765,N_19740);
nor U20596 (N_20596,N_19332,N_19030);
nor U20597 (N_20597,N_19607,N_19134);
and U20598 (N_20598,N_19223,N_19086);
and U20599 (N_20599,N_19052,N_18864);
or U20600 (N_20600,N_19209,N_19721);
and U20601 (N_20601,N_19037,N_18770);
nand U20602 (N_20602,N_19259,N_19480);
and U20603 (N_20603,N_19306,N_19778);
and U20604 (N_20604,N_19240,N_19285);
xor U20605 (N_20605,N_19813,N_19035);
nand U20606 (N_20606,N_19948,N_19518);
and U20607 (N_20607,N_19287,N_19460);
nor U20608 (N_20608,N_19893,N_19972);
and U20609 (N_20609,N_19649,N_19996);
nand U20610 (N_20610,N_19573,N_18796);
or U20611 (N_20611,N_19635,N_18978);
or U20612 (N_20612,N_19440,N_19011);
and U20613 (N_20613,N_19396,N_19615);
nand U20614 (N_20614,N_19983,N_19022);
and U20615 (N_20615,N_19565,N_19220);
or U20616 (N_20616,N_19128,N_19185);
nor U20617 (N_20617,N_19846,N_19031);
xor U20618 (N_20618,N_18760,N_19005);
nand U20619 (N_20619,N_19620,N_19879);
and U20620 (N_20620,N_19859,N_19409);
nand U20621 (N_20621,N_19727,N_19044);
xnor U20622 (N_20622,N_19645,N_18970);
and U20623 (N_20623,N_19941,N_18874);
xor U20624 (N_20624,N_19847,N_19744);
nand U20625 (N_20625,N_18822,N_19436);
or U20626 (N_20626,N_19254,N_18800);
nand U20627 (N_20627,N_19317,N_19023);
xor U20628 (N_20628,N_18869,N_19899);
and U20629 (N_20629,N_19577,N_19801);
nor U20630 (N_20630,N_19689,N_19130);
xnor U20631 (N_20631,N_19338,N_19193);
and U20632 (N_20632,N_19737,N_19484);
nor U20633 (N_20633,N_19547,N_19190);
or U20634 (N_20634,N_19783,N_19179);
nor U20635 (N_20635,N_19967,N_19142);
xnor U20636 (N_20636,N_18781,N_19067);
or U20637 (N_20637,N_18976,N_18997);
and U20638 (N_20638,N_18793,N_19394);
or U20639 (N_20639,N_19374,N_19025);
xor U20640 (N_20640,N_19986,N_19154);
or U20641 (N_20641,N_18974,N_19524);
nor U20642 (N_20642,N_19068,N_18954);
xor U20643 (N_20643,N_19387,N_19604);
xor U20644 (N_20644,N_19492,N_18819);
or U20645 (N_20645,N_18830,N_19990);
and U20646 (N_20646,N_19970,N_19984);
nand U20647 (N_20647,N_19179,N_19115);
or U20648 (N_20648,N_19880,N_19907);
or U20649 (N_20649,N_19820,N_19094);
nor U20650 (N_20650,N_18953,N_19458);
and U20651 (N_20651,N_19006,N_19674);
xnor U20652 (N_20652,N_19441,N_18916);
or U20653 (N_20653,N_19713,N_19042);
or U20654 (N_20654,N_19639,N_19643);
nand U20655 (N_20655,N_19480,N_19331);
nor U20656 (N_20656,N_19854,N_18806);
nor U20657 (N_20657,N_19250,N_19437);
or U20658 (N_20658,N_19485,N_18784);
nor U20659 (N_20659,N_19191,N_19410);
nor U20660 (N_20660,N_19409,N_18782);
nor U20661 (N_20661,N_19235,N_18753);
nor U20662 (N_20662,N_18805,N_18831);
or U20663 (N_20663,N_18975,N_19738);
xor U20664 (N_20664,N_19387,N_19602);
or U20665 (N_20665,N_18876,N_19420);
nand U20666 (N_20666,N_19281,N_19041);
nor U20667 (N_20667,N_19692,N_19405);
or U20668 (N_20668,N_18804,N_19733);
xor U20669 (N_20669,N_19921,N_19254);
nor U20670 (N_20670,N_19435,N_19588);
xor U20671 (N_20671,N_18878,N_19784);
and U20672 (N_20672,N_19410,N_19335);
or U20673 (N_20673,N_19065,N_19211);
xor U20674 (N_20674,N_19000,N_19576);
xor U20675 (N_20675,N_19753,N_19792);
xor U20676 (N_20676,N_19146,N_19135);
xnor U20677 (N_20677,N_19289,N_19579);
xnor U20678 (N_20678,N_18806,N_19926);
nand U20679 (N_20679,N_19467,N_18773);
xor U20680 (N_20680,N_18969,N_19029);
nor U20681 (N_20681,N_19989,N_19942);
nor U20682 (N_20682,N_19981,N_19551);
nand U20683 (N_20683,N_19734,N_18911);
nor U20684 (N_20684,N_19327,N_19218);
and U20685 (N_20685,N_19832,N_19330);
or U20686 (N_20686,N_19929,N_19482);
nand U20687 (N_20687,N_19478,N_19764);
or U20688 (N_20688,N_19495,N_19025);
and U20689 (N_20689,N_19144,N_19423);
and U20690 (N_20690,N_19052,N_19063);
or U20691 (N_20691,N_19888,N_18860);
or U20692 (N_20692,N_19011,N_19033);
or U20693 (N_20693,N_18912,N_19680);
or U20694 (N_20694,N_19106,N_19737);
nor U20695 (N_20695,N_19636,N_19135);
xor U20696 (N_20696,N_19185,N_19281);
nand U20697 (N_20697,N_19430,N_18909);
xnor U20698 (N_20698,N_19053,N_19150);
nor U20699 (N_20699,N_19458,N_19491);
or U20700 (N_20700,N_19636,N_19248);
nand U20701 (N_20701,N_19880,N_19494);
or U20702 (N_20702,N_19235,N_19549);
and U20703 (N_20703,N_18953,N_19093);
and U20704 (N_20704,N_19670,N_19039);
xor U20705 (N_20705,N_19108,N_19327);
and U20706 (N_20706,N_19465,N_18950);
nand U20707 (N_20707,N_18852,N_19201);
or U20708 (N_20708,N_19370,N_19167);
xnor U20709 (N_20709,N_19042,N_19838);
and U20710 (N_20710,N_19744,N_19800);
and U20711 (N_20711,N_19275,N_19195);
nor U20712 (N_20712,N_18984,N_19676);
and U20713 (N_20713,N_19285,N_19545);
nor U20714 (N_20714,N_19361,N_19804);
nand U20715 (N_20715,N_19270,N_18869);
xor U20716 (N_20716,N_19320,N_19027);
nor U20717 (N_20717,N_19983,N_19440);
nand U20718 (N_20718,N_19793,N_19075);
xnor U20719 (N_20719,N_19937,N_18864);
nor U20720 (N_20720,N_19649,N_18871);
or U20721 (N_20721,N_19455,N_19772);
or U20722 (N_20722,N_19919,N_19545);
and U20723 (N_20723,N_19864,N_19965);
nand U20724 (N_20724,N_19292,N_19145);
nor U20725 (N_20725,N_19518,N_18888);
and U20726 (N_20726,N_19034,N_19741);
or U20727 (N_20727,N_19444,N_19719);
or U20728 (N_20728,N_19401,N_19832);
nand U20729 (N_20729,N_19045,N_19709);
and U20730 (N_20730,N_18770,N_19417);
or U20731 (N_20731,N_18768,N_19772);
xor U20732 (N_20732,N_19839,N_19343);
or U20733 (N_20733,N_19520,N_19612);
and U20734 (N_20734,N_19697,N_19056);
nor U20735 (N_20735,N_19479,N_19813);
xor U20736 (N_20736,N_19387,N_19912);
nand U20737 (N_20737,N_19548,N_19412);
nand U20738 (N_20738,N_19437,N_19422);
nand U20739 (N_20739,N_19407,N_19191);
and U20740 (N_20740,N_19591,N_19246);
xnor U20741 (N_20741,N_19795,N_18866);
xnor U20742 (N_20742,N_19479,N_19001);
nand U20743 (N_20743,N_19473,N_19359);
or U20744 (N_20744,N_19371,N_18844);
nor U20745 (N_20745,N_19689,N_19027);
xor U20746 (N_20746,N_19293,N_18783);
nand U20747 (N_20747,N_18799,N_19511);
and U20748 (N_20748,N_19338,N_19171);
xnor U20749 (N_20749,N_19610,N_19758);
nor U20750 (N_20750,N_19222,N_19303);
nor U20751 (N_20751,N_18755,N_19537);
and U20752 (N_20752,N_19497,N_18784);
nor U20753 (N_20753,N_19372,N_19720);
or U20754 (N_20754,N_19358,N_19067);
xnor U20755 (N_20755,N_19101,N_19292);
nand U20756 (N_20756,N_19384,N_19131);
nor U20757 (N_20757,N_19153,N_18991);
or U20758 (N_20758,N_18805,N_19901);
nor U20759 (N_20759,N_19972,N_19284);
and U20760 (N_20760,N_19635,N_18945);
nand U20761 (N_20761,N_19029,N_19951);
nand U20762 (N_20762,N_18967,N_19348);
and U20763 (N_20763,N_19335,N_19726);
nor U20764 (N_20764,N_18816,N_19899);
nand U20765 (N_20765,N_18966,N_18826);
or U20766 (N_20766,N_19312,N_19198);
xnor U20767 (N_20767,N_18930,N_19436);
nor U20768 (N_20768,N_18835,N_19520);
or U20769 (N_20769,N_19259,N_18940);
xnor U20770 (N_20770,N_19636,N_19691);
nor U20771 (N_20771,N_19574,N_19883);
or U20772 (N_20772,N_19063,N_19715);
nand U20773 (N_20773,N_19419,N_19473);
and U20774 (N_20774,N_18868,N_18966);
xnor U20775 (N_20775,N_19208,N_19432);
nand U20776 (N_20776,N_19198,N_19055);
nand U20777 (N_20777,N_19982,N_18860);
nor U20778 (N_20778,N_18975,N_18881);
and U20779 (N_20779,N_19977,N_19443);
nand U20780 (N_20780,N_18946,N_19694);
or U20781 (N_20781,N_18860,N_19722);
nor U20782 (N_20782,N_19661,N_19118);
and U20783 (N_20783,N_19267,N_19755);
nand U20784 (N_20784,N_19984,N_19736);
xor U20785 (N_20785,N_19974,N_18793);
nand U20786 (N_20786,N_19908,N_19660);
nand U20787 (N_20787,N_19974,N_19214);
nand U20788 (N_20788,N_18806,N_19240);
nor U20789 (N_20789,N_19419,N_19175);
or U20790 (N_20790,N_19360,N_19249);
and U20791 (N_20791,N_19271,N_19031);
nand U20792 (N_20792,N_19603,N_19434);
and U20793 (N_20793,N_19727,N_19683);
and U20794 (N_20794,N_19345,N_19169);
xnor U20795 (N_20795,N_19477,N_19660);
nor U20796 (N_20796,N_18810,N_18822);
xor U20797 (N_20797,N_18903,N_19106);
nor U20798 (N_20798,N_19545,N_19840);
and U20799 (N_20799,N_19259,N_19665);
xor U20800 (N_20800,N_18951,N_19121);
nand U20801 (N_20801,N_19541,N_19246);
xor U20802 (N_20802,N_19510,N_19082);
and U20803 (N_20803,N_19463,N_19298);
nand U20804 (N_20804,N_19015,N_19352);
and U20805 (N_20805,N_18767,N_19023);
nand U20806 (N_20806,N_18932,N_19688);
nand U20807 (N_20807,N_19623,N_19344);
xnor U20808 (N_20808,N_19862,N_19765);
or U20809 (N_20809,N_19899,N_19434);
or U20810 (N_20810,N_19958,N_19075);
nand U20811 (N_20811,N_19149,N_19512);
and U20812 (N_20812,N_19262,N_19601);
or U20813 (N_20813,N_19846,N_19560);
or U20814 (N_20814,N_19374,N_19774);
and U20815 (N_20815,N_19843,N_19248);
or U20816 (N_20816,N_19380,N_19225);
xnor U20817 (N_20817,N_19617,N_19859);
and U20818 (N_20818,N_19756,N_19084);
xnor U20819 (N_20819,N_18839,N_18766);
and U20820 (N_20820,N_18821,N_19321);
and U20821 (N_20821,N_19260,N_19926);
nor U20822 (N_20822,N_18951,N_19877);
xnor U20823 (N_20823,N_19587,N_19891);
nand U20824 (N_20824,N_19565,N_19083);
nor U20825 (N_20825,N_18887,N_19619);
and U20826 (N_20826,N_19780,N_18797);
and U20827 (N_20827,N_19636,N_19640);
xnor U20828 (N_20828,N_19806,N_19586);
and U20829 (N_20829,N_19198,N_19669);
nand U20830 (N_20830,N_19895,N_19858);
nand U20831 (N_20831,N_19363,N_19143);
nor U20832 (N_20832,N_19705,N_19537);
xnor U20833 (N_20833,N_19589,N_19214);
xor U20834 (N_20834,N_19703,N_19115);
nor U20835 (N_20835,N_19265,N_19237);
nor U20836 (N_20836,N_19283,N_19368);
and U20837 (N_20837,N_19771,N_19821);
or U20838 (N_20838,N_18867,N_19379);
or U20839 (N_20839,N_19077,N_19567);
and U20840 (N_20840,N_19296,N_19679);
nand U20841 (N_20841,N_19099,N_19400);
nor U20842 (N_20842,N_19074,N_19744);
nor U20843 (N_20843,N_19567,N_19032);
nand U20844 (N_20844,N_19888,N_19194);
or U20845 (N_20845,N_19307,N_19969);
xor U20846 (N_20846,N_19566,N_19601);
nor U20847 (N_20847,N_18876,N_19056);
xnor U20848 (N_20848,N_19395,N_19413);
or U20849 (N_20849,N_19517,N_19833);
or U20850 (N_20850,N_19735,N_18770);
and U20851 (N_20851,N_18758,N_18805);
and U20852 (N_20852,N_19792,N_19698);
xnor U20853 (N_20853,N_19921,N_18881);
nor U20854 (N_20854,N_19410,N_19441);
xnor U20855 (N_20855,N_18851,N_19352);
nand U20856 (N_20856,N_19736,N_19743);
nand U20857 (N_20857,N_19977,N_19254);
xnor U20858 (N_20858,N_19905,N_19866);
xnor U20859 (N_20859,N_19352,N_19213);
nor U20860 (N_20860,N_18965,N_19064);
nand U20861 (N_20861,N_19042,N_19074);
xnor U20862 (N_20862,N_19418,N_19016);
or U20863 (N_20863,N_19419,N_19898);
or U20864 (N_20864,N_19409,N_19505);
and U20865 (N_20865,N_19807,N_19090);
and U20866 (N_20866,N_19444,N_18939);
nand U20867 (N_20867,N_19426,N_19132);
or U20868 (N_20868,N_18891,N_19405);
xor U20869 (N_20869,N_19123,N_19788);
xor U20870 (N_20870,N_18901,N_19986);
and U20871 (N_20871,N_18934,N_19215);
nor U20872 (N_20872,N_19342,N_19112);
or U20873 (N_20873,N_19531,N_19412);
nor U20874 (N_20874,N_19415,N_19910);
and U20875 (N_20875,N_19080,N_18950);
nand U20876 (N_20876,N_18967,N_19089);
xor U20877 (N_20877,N_19962,N_19526);
xor U20878 (N_20878,N_19606,N_19174);
xnor U20879 (N_20879,N_19242,N_18755);
nand U20880 (N_20880,N_18768,N_19777);
or U20881 (N_20881,N_19845,N_19950);
nand U20882 (N_20882,N_19931,N_19409);
xnor U20883 (N_20883,N_19444,N_19615);
or U20884 (N_20884,N_19123,N_19106);
nand U20885 (N_20885,N_18979,N_19079);
and U20886 (N_20886,N_19835,N_19210);
xor U20887 (N_20887,N_19981,N_19979);
xor U20888 (N_20888,N_19611,N_18898);
nand U20889 (N_20889,N_19140,N_19918);
nand U20890 (N_20890,N_19215,N_19627);
nor U20891 (N_20891,N_19137,N_18883);
or U20892 (N_20892,N_19874,N_18851);
or U20893 (N_20893,N_19869,N_19578);
nand U20894 (N_20894,N_18952,N_19647);
xor U20895 (N_20895,N_19977,N_18927);
nor U20896 (N_20896,N_19263,N_18813);
and U20897 (N_20897,N_18769,N_18937);
and U20898 (N_20898,N_19868,N_19552);
nor U20899 (N_20899,N_19935,N_19334);
and U20900 (N_20900,N_19071,N_19351);
nor U20901 (N_20901,N_19764,N_18883);
xor U20902 (N_20902,N_18874,N_19266);
xor U20903 (N_20903,N_19572,N_19813);
nor U20904 (N_20904,N_19740,N_19131);
and U20905 (N_20905,N_19793,N_18924);
and U20906 (N_20906,N_18855,N_19981);
xnor U20907 (N_20907,N_19869,N_19456);
or U20908 (N_20908,N_19294,N_18876);
nand U20909 (N_20909,N_19561,N_19255);
nand U20910 (N_20910,N_18983,N_19505);
nor U20911 (N_20911,N_19917,N_18779);
or U20912 (N_20912,N_19862,N_19048);
nand U20913 (N_20913,N_18811,N_19967);
nand U20914 (N_20914,N_18815,N_19107);
or U20915 (N_20915,N_19800,N_19872);
nor U20916 (N_20916,N_19845,N_19881);
nand U20917 (N_20917,N_19122,N_19714);
nor U20918 (N_20918,N_19180,N_19589);
and U20919 (N_20919,N_19832,N_19885);
and U20920 (N_20920,N_19865,N_19114);
xnor U20921 (N_20921,N_19367,N_19244);
and U20922 (N_20922,N_19468,N_19802);
nand U20923 (N_20923,N_19509,N_18883);
or U20924 (N_20924,N_19022,N_18912);
and U20925 (N_20925,N_19692,N_19526);
xor U20926 (N_20926,N_19704,N_19478);
nor U20927 (N_20927,N_19215,N_19664);
and U20928 (N_20928,N_18871,N_19772);
nor U20929 (N_20929,N_19280,N_19900);
or U20930 (N_20930,N_19143,N_19869);
nor U20931 (N_20931,N_19414,N_19975);
and U20932 (N_20932,N_19643,N_19996);
nand U20933 (N_20933,N_19687,N_19417);
nor U20934 (N_20934,N_18762,N_18942);
xor U20935 (N_20935,N_19676,N_18928);
nor U20936 (N_20936,N_19554,N_19674);
nor U20937 (N_20937,N_18859,N_19674);
nor U20938 (N_20938,N_19044,N_19989);
or U20939 (N_20939,N_18910,N_18791);
nor U20940 (N_20940,N_19178,N_19712);
and U20941 (N_20941,N_19785,N_19470);
nand U20942 (N_20942,N_19257,N_18759);
and U20943 (N_20943,N_19529,N_19343);
and U20944 (N_20944,N_19227,N_19302);
xnor U20945 (N_20945,N_18783,N_18822);
xor U20946 (N_20946,N_19697,N_19170);
nor U20947 (N_20947,N_19492,N_19525);
and U20948 (N_20948,N_19463,N_18885);
xnor U20949 (N_20949,N_18951,N_18839);
xor U20950 (N_20950,N_19527,N_18834);
xnor U20951 (N_20951,N_19363,N_19698);
and U20952 (N_20952,N_19032,N_19574);
xor U20953 (N_20953,N_18778,N_19598);
xor U20954 (N_20954,N_18912,N_19333);
nor U20955 (N_20955,N_18947,N_19574);
nand U20956 (N_20956,N_19043,N_19606);
nand U20957 (N_20957,N_18860,N_19423);
nand U20958 (N_20958,N_19041,N_19858);
xor U20959 (N_20959,N_19736,N_19128);
nor U20960 (N_20960,N_19693,N_19976);
and U20961 (N_20961,N_19220,N_19626);
or U20962 (N_20962,N_19096,N_19603);
and U20963 (N_20963,N_19652,N_19950);
nand U20964 (N_20964,N_19628,N_19399);
xor U20965 (N_20965,N_19880,N_19257);
nand U20966 (N_20966,N_19052,N_19993);
nor U20967 (N_20967,N_18872,N_19403);
nor U20968 (N_20968,N_18914,N_19506);
nor U20969 (N_20969,N_19354,N_19811);
and U20970 (N_20970,N_19280,N_19797);
xor U20971 (N_20971,N_18992,N_19093);
xor U20972 (N_20972,N_19614,N_19914);
nor U20973 (N_20973,N_19256,N_19125);
xnor U20974 (N_20974,N_19550,N_19037);
and U20975 (N_20975,N_19412,N_19356);
nand U20976 (N_20976,N_19723,N_19840);
nor U20977 (N_20977,N_18791,N_19822);
nand U20978 (N_20978,N_19288,N_18890);
and U20979 (N_20979,N_19619,N_19071);
nor U20980 (N_20980,N_19563,N_19371);
and U20981 (N_20981,N_19963,N_19019);
xor U20982 (N_20982,N_19866,N_18931);
or U20983 (N_20983,N_19446,N_19855);
xor U20984 (N_20984,N_19202,N_19988);
nor U20985 (N_20985,N_19095,N_19534);
and U20986 (N_20986,N_19343,N_19257);
xor U20987 (N_20987,N_19802,N_19226);
or U20988 (N_20988,N_19087,N_18817);
nand U20989 (N_20989,N_19344,N_19049);
nand U20990 (N_20990,N_19929,N_18754);
nand U20991 (N_20991,N_18762,N_19391);
or U20992 (N_20992,N_18909,N_18993);
xnor U20993 (N_20993,N_19767,N_19830);
or U20994 (N_20994,N_19061,N_19451);
and U20995 (N_20995,N_19344,N_18955);
and U20996 (N_20996,N_18881,N_19947);
and U20997 (N_20997,N_19817,N_19989);
nand U20998 (N_20998,N_19531,N_18819);
xor U20999 (N_20999,N_19022,N_19769);
nand U21000 (N_21000,N_19172,N_19821);
nand U21001 (N_21001,N_19272,N_19116);
nand U21002 (N_21002,N_19863,N_19103);
xor U21003 (N_21003,N_19449,N_19962);
or U21004 (N_21004,N_19531,N_18901);
or U21005 (N_21005,N_19096,N_18791);
and U21006 (N_21006,N_19579,N_19583);
nand U21007 (N_21007,N_19530,N_19807);
xnor U21008 (N_21008,N_18894,N_19568);
and U21009 (N_21009,N_19509,N_19775);
or U21010 (N_21010,N_19378,N_19563);
nor U21011 (N_21011,N_18874,N_18812);
or U21012 (N_21012,N_19491,N_19477);
nand U21013 (N_21013,N_19139,N_19560);
xor U21014 (N_21014,N_19393,N_19780);
nor U21015 (N_21015,N_19772,N_19161);
nand U21016 (N_21016,N_18886,N_18815);
nand U21017 (N_21017,N_19658,N_19346);
and U21018 (N_21018,N_19921,N_19552);
or U21019 (N_21019,N_18774,N_19467);
nand U21020 (N_21020,N_19549,N_19353);
xor U21021 (N_21021,N_18982,N_19138);
or U21022 (N_21022,N_18928,N_18856);
or U21023 (N_21023,N_19126,N_19445);
and U21024 (N_21024,N_19544,N_19307);
nand U21025 (N_21025,N_19420,N_19168);
nor U21026 (N_21026,N_18866,N_19261);
and U21027 (N_21027,N_19417,N_19427);
or U21028 (N_21028,N_19708,N_18777);
and U21029 (N_21029,N_19051,N_18760);
nand U21030 (N_21030,N_19504,N_18899);
and U21031 (N_21031,N_19243,N_19149);
nor U21032 (N_21032,N_19874,N_19863);
or U21033 (N_21033,N_19573,N_19762);
or U21034 (N_21034,N_19064,N_19297);
and U21035 (N_21035,N_18845,N_19688);
nor U21036 (N_21036,N_19354,N_19305);
xor U21037 (N_21037,N_19461,N_19685);
nand U21038 (N_21038,N_19100,N_19910);
and U21039 (N_21039,N_19348,N_18895);
nor U21040 (N_21040,N_19690,N_19804);
and U21041 (N_21041,N_19613,N_19158);
xor U21042 (N_21042,N_18767,N_18985);
xnor U21043 (N_21043,N_19925,N_19723);
and U21044 (N_21044,N_19778,N_18956);
and U21045 (N_21045,N_19548,N_18804);
nand U21046 (N_21046,N_19127,N_19363);
nand U21047 (N_21047,N_18890,N_19122);
nor U21048 (N_21048,N_19377,N_19790);
or U21049 (N_21049,N_19523,N_19099);
nand U21050 (N_21050,N_19824,N_19206);
nor U21051 (N_21051,N_19295,N_19829);
nand U21052 (N_21052,N_18970,N_19962);
and U21053 (N_21053,N_18987,N_18840);
xnor U21054 (N_21054,N_19808,N_18868);
or U21055 (N_21055,N_19612,N_19460);
or U21056 (N_21056,N_19183,N_19521);
xor U21057 (N_21057,N_19253,N_18756);
xnor U21058 (N_21058,N_19883,N_19222);
nor U21059 (N_21059,N_18978,N_19055);
nor U21060 (N_21060,N_19584,N_19180);
nand U21061 (N_21061,N_19613,N_19600);
or U21062 (N_21062,N_19069,N_19314);
nor U21063 (N_21063,N_19299,N_19241);
or U21064 (N_21064,N_19681,N_19685);
xnor U21065 (N_21065,N_19551,N_19700);
nor U21066 (N_21066,N_19513,N_19168);
nor U21067 (N_21067,N_19149,N_19348);
or U21068 (N_21068,N_19996,N_18851);
xor U21069 (N_21069,N_18992,N_19042);
nand U21070 (N_21070,N_19277,N_19637);
xor U21071 (N_21071,N_19666,N_19853);
and U21072 (N_21072,N_19072,N_19505);
nor U21073 (N_21073,N_19236,N_19615);
nand U21074 (N_21074,N_19762,N_19318);
xnor U21075 (N_21075,N_19575,N_19244);
xnor U21076 (N_21076,N_19523,N_19626);
nor U21077 (N_21077,N_19724,N_19766);
or U21078 (N_21078,N_19352,N_18790);
nor U21079 (N_21079,N_19861,N_19201);
and U21080 (N_21080,N_19092,N_19681);
or U21081 (N_21081,N_19738,N_19795);
nor U21082 (N_21082,N_18858,N_19366);
or U21083 (N_21083,N_18825,N_19544);
xnor U21084 (N_21084,N_19418,N_19931);
and U21085 (N_21085,N_19377,N_19243);
or U21086 (N_21086,N_19933,N_19062);
nor U21087 (N_21087,N_19741,N_19905);
xnor U21088 (N_21088,N_19676,N_19005);
and U21089 (N_21089,N_18883,N_19932);
or U21090 (N_21090,N_19203,N_18898);
xor U21091 (N_21091,N_18906,N_18948);
xor U21092 (N_21092,N_19590,N_19770);
xor U21093 (N_21093,N_19552,N_19762);
xor U21094 (N_21094,N_19282,N_19629);
nor U21095 (N_21095,N_19541,N_19060);
xor U21096 (N_21096,N_18797,N_19065);
and U21097 (N_21097,N_19102,N_19510);
nand U21098 (N_21098,N_19480,N_19902);
nand U21099 (N_21099,N_19524,N_18820);
nand U21100 (N_21100,N_18757,N_19069);
or U21101 (N_21101,N_19040,N_19215);
xnor U21102 (N_21102,N_18817,N_19275);
nand U21103 (N_21103,N_19030,N_19826);
nand U21104 (N_21104,N_19571,N_19921);
xnor U21105 (N_21105,N_18910,N_18988);
and U21106 (N_21106,N_19686,N_19320);
and U21107 (N_21107,N_19496,N_19699);
or U21108 (N_21108,N_18810,N_19803);
nor U21109 (N_21109,N_19206,N_19425);
or U21110 (N_21110,N_18998,N_19818);
or U21111 (N_21111,N_18997,N_18795);
nand U21112 (N_21112,N_18752,N_18860);
or U21113 (N_21113,N_19455,N_19956);
nor U21114 (N_21114,N_19751,N_19499);
nand U21115 (N_21115,N_18911,N_19879);
or U21116 (N_21116,N_19216,N_19137);
xor U21117 (N_21117,N_19314,N_19959);
xnor U21118 (N_21118,N_19173,N_19750);
nand U21119 (N_21119,N_18915,N_19184);
and U21120 (N_21120,N_19835,N_18792);
nor U21121 (N_21121,N_19612,N_19105);
nor U21122 (N_21122,N_18999,N_18756);
xor U21123 (N_21123,N_19530,N_19557);
nand U21124 (N_21124,N_19986,N_19880);
xnor U21125 (N_21125,N_19806,N_19673);
nand U21126 (N_21126,N_19383,N_19620);
nor U21127 (N_21127,N_19924,N_19339);
and U21128 (N_21128,N_19442,N_19451);
or U21129 (N_21129,N_19037,N_19461);
nand U21130 (N_21130,N_19991,N_19275);
xor U21131 (N_21131,N_18835,N_19840);
nand U21132 (N_21132,N_19713,N_19470);
or U21133 (N_21133,N_19158,N_18759);
and U21134 (N_21134,N_18993,N_18866);
and U21135 (N_21135,N_18931,N_19554);
or U21136 (N_21136,N_19926,N_19547);
xor U21137 (N_21137,N_19413,N_19353);
xor U21138 (N_21138,N_19285,N_19841);
nor U21139 (N_21139,N_18894,N_18897);
xnor U21140 (N_21140,N_19404,N_19286);
nor U21141 (N_21141,N_19541,N_19740);
nor U21142 (N_21142,N_19839,N_19066);
and U21143 (N_21143,N_18960,N_19587);
and U21144 (N_21144,N_19796,N_19786);
nor U21145 (N_21145,N_19737,N_18875);
and U21146 (N_21146,N_19570,N_19439);
or U21147 (N_21147,N_19879,N_19580);
and U21148 (N_21148,N_18997,N_19948);
or U21149 (N_21149,N_19206,N_19341);
nor U21150 (N_21150,N_19202,N_19401);
and U21151 (N_21151,N_19463,N_19377);
nor U21152 (N_21152,N_19672,N_18858);
xor U21153 (N_21153,N_19049,N_19369);
or U21154 (N_21154,N_19690,N_19106);
nand U21155 (N_21155,N_19215,N_19639);
nor U21156 (N_21156,N_19490,N_19699);
xnor U21157 (N_21157,N_19481,N_19938);
and U21158 (N_21158,N_19325,N_19343);
and U21159 (N_21159,N_19811,N_18842);
and U21160 (N_21160,N_19140,N_19706);
or U21161 (N_21161,N_19728,N_19916);
nand U21162 (N_21162,N_19462,N_19542);
and U21163 (N_21163,N_19780,N_19042);
nand U21164 (N_21164,N_19998,N_18907);
nand U21165 (N_21165,N_19560,N_19555);
nor U21166 (N_21166,N_19755,N_19463);
or U21167 (N_21167,N_18959,N_19461);
or U21168 (N_21168,N_19586,N_18840);
and U21169 (N_21169,N_19754,N_19741);
nor U21170 (N_21170,N_19069,N_19278);
nor U21171 (N_21171,N_19633,N_19598);
and U21172 (N_21172,N_19275,N_19759);
nand U21173 (N_21173,N_19673,N_19913);
xor U21174 (N_21174,N_19882,N_19284);
or U21175 (N_21175,N_19417,N_19819);
or U21176 (N_21176,N_19736,N_19486);
and U21177 (N_21177,N_19969,N_19648);
xor U21178 (N_21178,N_19308,N_18853);
nor U21179 (N_21179,N_18912,N_19903);
xor U21180 (N_21180,N_19540,N_19119);
xnor U21181 (N_21181,N_18847,N_19406);
nand U21182 (N_21182,N_19372,N_19342);
nor U21183 (N_21183,N_19938,N_19092);
nand U21184 (N_21184,N_18808,N_18806);
and U21185 (N_21185,N_19587,N_19833);
nor U21186 (N_21186,N_19097,N_19316);
nor U21187 (N_21187,N_19504,N_19065);
or U21188 (N_21188,N_19016,N_19961);
nor U21189 (N_21189,N_18935,N_18855);
xnor U21190 (N_21190,N_19321,N_19480);
or U21191 (N_21191,N_19659,N_19970);
or U21192 (N_21192,N_19573,N_19370);
nand U21193 (N_21193,N_19218,N_19555);
or U21194 (N_21194,N_19297,N_19956);
or U21195 (N_21195,N_18769,N_19014);
nand U21196 (N_21196,N_19888,N_18759);
xor U21197 (N_21197,N_19306,N_19347);
nand U21198 (N_21198,N_19186,N_19260);
and U21199 (N_21199,N_19462,N_19376);
nor U21200 (N_21200,N_18870,N_19442);
and U21201 (N_21201,N_18873,N_18867);
and U21202 (N_21202,N_18973,N_18844);
xnor U21203 (N_21203,N_18930,N_19993);
and U21204 (N_21204,N_19263,N_19709);
or U21205 (N_21205,N_18805,N_19587);
xnor U21206 (N_21206,N_19703,N_19934);
nand U21207 (N_21207,N_19191,N_19471);
xnor U21208 (N_21208,N_19038,N_19799);
nand U21209 (N_21209,N_18983,N_19788);
and U21210 (N_21210,N_18776,N_19054);
or U21211 (N_21211,N_19686,N_18907);
nor U21212 (N_21212,N_19942,N_19567);
or U21213 (N_21213,N_19275,N_19220);
and U21214 (N_21214,N_19371,N_19079);
xor U21215 (N_21215,N_18941,N_19064);
nand U21216 (N_21216,N_19439,N_19687);
nand U21217 (N_21217,N_18944,N_19760);
nor U21218 (N_21218,N_18862,N_19475);
or U21219 (N_21219,N_19917,N_19725);
and U21220 (N_21220,N_19732,N_19634);
or U21221 (N_21221,N_18968,N_19334);
nand U21222 (N_21222,N_19174,N_19471);
nor U21223 (N_21223,N_19381,N_19636);
and U21224 (N_21224,N_19731,N_18897);
or U21225 (N_21225,N_19762,N_19222);
nand U21226 (N_21226,N_19412,N_19732);
nand U21227 (N_21227,N_18860,N_18804);
and U21228 (N_21228,N_18907,N_19488);
xor U21229 (N_21229,N_19090,N_19881);
nand U21230 (N_21230,N_19435,N_19510);
nor U21231 (N_21231,N_19354,N_18915);
and U21232 (N_21232,N_19961,N_19316);
nand U21233 (N_21233,N_19986,N_18866);
nor U21234 (N_21234,N_18813,N_18799);
or U21235 (N_21235,N_18963,N_18810);
and U21236 (N_21236,N_19714,N_19377);
or U21237 (N_21237,N_19554,N_19075);
nor U21238 (N_21238,N_19513,N_19435);
and U21239 (N_21239,N_19143,N_19093);
and U21240 (N_21240,N_19237,N_19978);
xor U21241 (N_21241,N_18935,N_19819);
xnor U21242 (N_21242,N_19127,N_19661);
nor U21243 (N_21243,N_19321,N_19109);
or U21244 (N_21244,N_18760,N_19707);
xnor U21245 (N_21245,N_19973,N_19831);
nand U21246 (N_21246,N_19128,N_19391);
nor U21247 (N_21247,N_19207,N_19193);
nand U21248 (N_21248,N_18996,N_19559);
xnor U21249 (N_21249,N_18979,N_18766);
nand U21250 (N_21250,N_21131,N_21105);
or U21251 (N_21251,N_21058,N_21101);
or U21252 (N_21252,N_20011,N_20669);
and U21253 (N_21253,N_20149,N_20302);
xor U21254 (N_21254,N_21174,N_20244);
nor U21255 (N_21255,N_20278,N_20092);
and U21256 (N_21256,N_20164,N_20965);
nor U21257 (N_21257,N_20635,N_20785);
and U21258 (N_21258,N_20286,N_21113);
or U21259 (N_21259,N_20409,N_20346);
nor U21260 (N_21260,N_20437,N_20502);
nor U21261 (N_21261,N_21138,N_20827);
xor U21262 (N_21262,N_20717,N_20883);
nand U21263 (N_21263,N_21239,N_20249);
xnor U21264 (N_21264,N_20866,N_20279);
xor U21265 (N_21265,N_20751,N_20536);
nor U21266 (N_21266,N_20850,N_21163);
nand U21267 (N_21267,N_20903,N_20018);
nor U21268 (N_21268,N_20436,N_20742);
nor U21269 (N_21269,N_20255,N_20939);
or U21270 (N_21270,N_20985,N_20837);
and U21271 (N_21271,N_20446,N_20445);
nand U21272 (N_21272,N_21097,N_20479);
nand U21273 (N_21273,N_20563,N_20604);
nor U21274 (N_21274,N_21036,N_20429);
nand U21275 (N_21275,N_21205,N_20661);
nor U21276 (N_21276,N_21184,N_20841);
and U21277 (N_21277,N_20304,N_21209);
or U21278 (N_21278,N_20095,N_20687);
nand U21279 (N_21279,N_20540,N_20703);
or U21280 (N_21280,N_20838,N_21090);
nor U21281 (N_21281,N_20747,N_20078);
and U21282 (N_21282,N_20498,N_21094);
or U21283 (N_21283,N_21236,N_20013);
nor U21284 (N_21284,N_20217,N_20443);
xor U21285 (N_21285,N_20642,N_20031);
or U21286 (N_21286,N_20594,N_20280);
nand U21287 (N_21287,N_20268,N_20801);
nor U21288 (N_21288,N_20177,N_21040);
xor U21289 (N_21289,N_20601,N_20514);
nand U21290 (N_21290,N_20069,N_20824);
xnor U21291 (N_21291,N_20607,N_20526);
or U21292 (N_21292,N_20836,N_21162);
nand U21293 (N_21293,N_21079,N_21132);
xnor U21294 (N_21294,N_20958,N_20968);
nand U21295 (N_21295,N_21054,N_20954);
nand U21296 (N_21296,N_20943,N_20105);
nor U21297 (N_21297,N_20351,N_20768);
and U21298 (N_21298,N_20267,N_20758);
nor U21299 (N_21299,N_20276,N_20401);
or U21300 (N_21300,N_20405,N_20690);
xnor U21301 (N_21301,N_21008,N_20251);
nand U21302 (N_21302,N_20885,N_20061);
or U21303 (N_21303,N_20593,N_20929);
nand U21304 (N_21304,N_20561,N_20241);
and U21305 (N_21305,N_20822,N_20422);
or U21306 (N_21306,N_20362,N_20353);
and U21307 (N_21307,N_21213,N_20997);
and U21308 (N_21308,N_20226,N_20157);
xor U21309 (N_21309,N_20951,N_20388);
xor U21310 (N_21310,N_20865,N_21196);
or U21311 (N_21311,N_21023,N_21150);
nor U21312 (N_21312,N_20392,N_20355);
nor U21313 (N_21313,N_20343,N_21042);
xor U21314 (N_21314,N_20963,N_21026);
xor U21315 (N_21315,N_20732,N_20860);
or U21316 (N_21316,N_20432,N_20010);
and U21317 (N_21317,N_20222,N_20789);
nand U21318 (N_21318,N_20535,N_20356);
and U21319 (N_21319,N_20052,N_20724);
or U21320 (N_21320,N_20495,N_20833);
nor U21321 (N_21321,N_20935,N_20472);
nand U21322 (N_21322,N_20532,N_21207);
or U21323 (N_21323,N_21043,N_20391);
or U21324 (N_21324,N_20757,N_20266);
xor U21325 (N_21325,N_20488,N_20839);
or U21326 (N_21326,N_20112,N_21165);
or U21327 (N_21327,N_20066,N_21035);
and U21328 (N_21328,N_20274,N_20447);
nor U21329 (N_21329,N_20589,N_20761);
and U21330 (N_21330,N_20901,N_20908);
nor U21331 (N_21331,N_20085,N_20250);
nor U21332 (N_21332,N_21219,N_20277);
nor U21333 (N_21333,N_20017,N_21224);
nor U21334 (N_21334,N_20229,N_20987);
nand U21335 (N_21335,N_20133,N_20897);
and U21336 (N_21336,N_20281,N_21048);
and U21337 (N_21337,N_20097,N_20870);
or U21338 (N_21338,N_20109,N_21084);
nor U21339 (N_21339,N_20537,N_20120);
and U21340 (N_21340,N_21197,N_21228);
or U21341 (N_21341,N_20547,N_20867);
and U21342 (N_21342,N_20888,N_21231);
nor U21343 (N_21343,N_20397,N_20370);
and U21344 (N_21344,N_20764,N_21067);
xnor U21345 (N_21345,N_21160,N_20887);
xnor U21346 (N_21346,N_20981,N_20360);
xnor U21347 (N_21347,N_21137,N_20350);
nor U21348 (N_21348,N_21088,N_20273);
nand U21349 (N_21349,N_20609,N_20787);
nor U21350 (N_21350,N_21147,N_21248);
nand U21351 (N_21351,N_20671,N_20380);
xor U21352 (N_21352,N_20725,N_20913);
xor U21353 (N_21353,N_20199,N_21214);
or U21354 (N_21354,N_20975,N_20426);
xnor U21355 (N_21355,N_20541,N_20420);
xnor U21356 (N_21356,N_20332,N_20922);
xnor U21357 (N_21357,N_20745,N_21059);
nor U21358 (N_21358,N_20524,N_20419);
xor U21359 (N_21359,N_20826,N_20947);
nand U21360 (N_21360,N_20167,N_20904);
or U21361 (N_21361,N_20932,N_20723);
and U21362 (N_21362,N_20428,N_21051);
and U21363 (N_21363,N_20361,N_20118);
nor U21364 (N_21364,N_20040,N_20709);
nand U21365 (N_21365,N_21225,N_20666);
nor U21366 (N_21366,N_20802,N_20618);
xor U21367 (N_21367,N_20091,N_20608);
xor U21368 (N_21368,N_20243,N_20086);
xnor U21369 (N_21369,N_21047,N_21107);
nor U21370 (N_21370,N_20170,N_20633);
or U21371 (N_21371,N_20211,N_20795);
and U21372 (N_21372,N_20966,N_20704);
or U21373 (N_21373,N_20510,N_20894);
xor U21374 (N_21374,N_20363,N_20813);
nor U21375 (N_21375,N_20191,N_20053);
nor U21376 (N_21376,N_20708,N_21186);
xnor U21377 (N_21377,N_20235,N_20832);
nand U21378 (N_21378,N_21151,N_20319);
nand U21379 (N_21379,N_20744,N_21216);
or U21380 (N_21380,N_20676,N_20743);
and U21381 (N_21381,N_20679,N_20693);
xnor U21382 (N_21382,N_20046,N_21055);
and U21383 (N_21383,N_20068,N_20777);
xnor U21384 (N_21384,N_20588,N_20686);
xor U21385 (N_21385,N_20408,N_20478);
and U21386 (N_21386,N_20734,N_20512);
nor U21387 (N_21387,N_20634,N_21111);
xor U21388 (N_21388,N_20342,N_21100);
and U21389 (N_21389,N_20174,N_21112);
nor U21390 (N_21390,N_20299,N_20560);
nand U21391 (N_21391,N_21108,N_20135);
nand U21392 (N_21392,N_20315,N_20600);
and U21393 (N_21393,N_20579,N_20469);
or U21394 (N_21394,N_21103,N_20859);
nand U21395 (N_21395,N_20400,N_21077);
nor U21396 (N_21396,N_21096,N_20624);
and U21397 (N_21397,N_21235,N_20379);
nor U21398 (N_21398,N_20658,N_20944);
and U21399 (N_21399,N_21156,N_20729);
nor U21400 (N_21400,N_21030,N_21007);
or U21401 (N_21401,N_20493,N_20584);
and U21402 (N_21402,N_20875,N_20372);
or U21403 (N_21403,N_20741,N_21016);
nor U21404 (N_21404,N_21172,N_20387);
nor U21405 (N_21405,N_20182,N_20863);
nor U21406 (N_21406,N_20873,N_20145);
and U21407 (N_21407,N_20337,N_20270);
nor U21408 (N_21408,N_20035,N_20938);
or U21409 (N_21409,N_21117,N_20127);
and U21410 (N_21410,N_21130,N_21063);
and U21411 (N_21411,N_20236,N_20992);
nor U21412 (N_21412,N_20962,N_20995);
and U21413 (N_21413,N_21179,N_20204);
nor U21414 (N_21414,N_20808,N_20489);
and U21415 (N_21415,N_20978,N_21182);
nor U21416 (N_21416,N_20759,N_20440);
or U21417 (N_21417,N_20779,N_20680);
nand U21418 (N_21418,N_20988,N_20718);
or U21419 (N_21419,N_20189,N_20862);
or U21420 (N_21420,N_21126,N_20716);
nor U21421 (N_21421,N_20208,N_20007);
nand U21422 (N_21422,N_21073,N_20934);
nor U21423 (N_21423,N_20989,N_20188);
xnor U21424 (N_21424,N_20874,N_20821);
nor U21425 (N_21425,N_20016,N_20272);
nor U21426 (N_21426,N_20702,N_20119);
nand U21427 (N_21427,N_21052,N_20444);
xnor U21428 (N_21428,N_20684,N_20321);
or U21429 (N_21429,N_20413,N_20014);
or U21430 (N_21430,N_20258,N_20575);
or U21431 (N_21431,N_20653,N_21173);
and U21432 (N_21432,N_20074,N_21245);
nand U21433 (N_21433,N_20287,N_20663);
xnor U21434 (N_21434,N_20364,N_20650);
and U21435 (N_21435,N_21099,N_20291);
nor U21436 (N_21436,N_20316,N_20647);
nand U21437 (N_21437,N_20848,N_20621);
nand U21438 (N_21438,N_20238,N_20158);
xor U21439 (N_21439,N_20622,N_20282);
xnor U21440 (N_21440,N_20871,N_20187);
or U21441 (N_21441,N_20660,N_20615);
or U21442 (N_21442,N_20854,N_20314);
xnor U21443 (N_21443,N_20701,N_20322);
nand U21444 (N_21444,N_21218,N_20142);
or U21445 (N_21445,N_20856,N_20890);
nor U21446 (N_21446,N_20610,N_20386);
nor U21447 (N_21447,N_20089,N_21102);
or U21448 (N_21448,N_20843,N_20937);
nor U21449 (N_21449,N_20060,N_20691);
or U21450 (N_21450,N_20739,N_20946);
nor U21451 (N_21451,N_21064,N_20193);
nand U21452 (N_21452,N_20215,N_20721);
xor U21453 (N_21453,N_20090,N_20398);
nand U21454 (N_21454,N_20899,N_20218);
nand U21455 (N_21455,N_20829,N_20039);
xor U21456 (N_21456,N_21001,N_20156);
nor U21457 (N_21457,N_21208,N_21068);
nor U21458 (N_21458,N_20318,N_21085);
nor U21459 (N_21459,N_20054,N_20203);
or U21460 (N_21460,N_20959,N_20245);
nor U21461 (N_21461,N_21009,N_20763);
nand U21462 (N_21462,N_20034,N_21164);
nand U21463 (N_21463,N_20043,N_20956);
and U21464 (N_21464,N_20809,N_20945);
xnor U21465 (N_21465,N_20186,N_20375);
or U21466 (N_21466,N_20916,N_20309);
and U21467 (N_21467,N_20571,N_20819);
nor U21468 (N_21468,N_21161,N_20210);
or U21469 (N_21469,N_20325,N_20688);
or U21470 (N_21470,N_20807,N_21221);
nor U21471 (N_21471,N_21154,N_20804);
nor U21472 (N_21472,N_20008,N_21081);
or U21473 (N_21473,N_20465,N_21038);
nand U21474 (N_21474,N_20448,N_20825);
and U21475 (N_21475,N_20626,N_21191);
xor U21476 (N_21476,N_20000,N_20855);
nand U21477 (N_21477,N_20404,N_20207);
or U21478 (N_21478,N_20760,N_20161);
xnor U21479 (N_21479,N_20698,N_20065);
xnor U21480 (N_21480,N_20221,N_20651);
and U21481 (N_21481,N_20116,N_21033);
xor U21482 (N_21482,N_20129,N_20410);
nor U21483 (N_21483,N_20376,N_20652);
or U21484 (N_21484,N_21168,N_20383);
nand U21485 (N_21485,N_20574,N_21141);
xnor U21486 (N_21486,N_20898,N_20662);
nand U21487 (N_21487,N_20788,N_20290);
nand U21488 (N_21488,N_20835,N_21241);
xor U21489 (N_21489,N_21198,N_20632);
nor U21490 (N_21490,N_20190,N_20692);
nand U21491 (N_21491,N_20394,N_20339);
xor U21492 (N_21492,N_20590,N_20817);
nor U21493 (N_21493,N_21069,N_20872);
xnor U21494 (N_21494,N_20303,N_20998);
and U21495 (N_21495,N_20476,N_20949);
nor U21496 (N_21496,N_20453,N_20513);
xnor U21497 (N_21497,N_20449,N_20631);
nand U21498 (N_21498,N_21065,N_20461);
or U21499 (N_21499,N_20033,N_21127);
nand U21500 (N_21500,N_20056,N_20301);
nand U21501 (N_21501,N_20131,N_20638);
xnor U21502 (N_21502,N_20330,N_20504);
nor U21503 (N_21503,N_20545,N_20727);
nand U21504 (N_21504,N_21183,N_21187);
and U21505 (N_21505,N_20749,N_21136);
and U21506 (N_21506,N_20275,N_20549);
and U21507 (N_21507,N_20672,N_20578);
and U21508 (N_21508,N_20715,N_21249);
xor U21509 (N_21509,N_20424,N_20689);
nor U21510 (N_21510,N_20214,N_20490);
nand U21511 (N_21511,N_20811,N_21017);
or U21512 (N_21512,N_20644,N_20002);
nor U21513 (N_21513,N_20463,N_20613);
and U21514 (N_21514,N_20227,N_21233);
nand U21515 (N_21515,N_20736,N_20507);
xnor U21516 (N_21516,N_20543,N_20096);
nand U21517 (N_21517,N_20623,N_20531);
and U21518 (N_21518,N_20783,N_20990);
xnor U21519 (N_21519,N_20076,N_21206);
nor U21520 (N_21520,N_20983,N_20231);
and U21521 (N_21521,N_20637,N_20773);
and U21522 (N_21522,N_20884,N_20844);
xnor U21523 (N_21523,N_20402,N_20442);
nand U21524 (N_21524,N_20026,N_20766);
or U21525 (N_21525,N_20906,N_20880);
xor U21526 (N_21526,N_21222,N_20641);
nand U21527 (N_21527,N_20412,N_20212);
nor U21528 (N_21528,N_20617,N_20123);
nor U21529 (N_21529,N_20840,N_20542);
or U21530 (N_21530,N_20924,N_20602);
xnor U21531 (N_21531,N_21075,N_20786);
nor U21532 (N_21532,N_20497,N_20746);
xor U21533 (N_21533,N_20972,N_20247);
and U21534 (N_21534,N_20357,N_20639);
nand U21535 (N_21535,N_21135,N_21010);
or U21536 (N_21536,N_20657,N_20707);
or U21537 (N_21537,N_21142,N_20735);
or U21538 (N_21538,N_20328,N_20996);
xnor U21539 (N_21539,N_20029,N_20414);
nand U21540 (N_21540,N_20668,N_21159);
or U21541 (N_21541,N_20919,N_20103);
or U21542 (N_21542,N_20506,N_20460);
or U21543 (N_21543,N_20101,N_20242);
and U21544 (N_21544,N_20847,N_20952);
and U21545 (N_21545,N_20077,N_20100);
nor U21546 (N_21546,N_21238,N_21133);
nor U21547 (N_21547,N_21177,N_21110);
xnor U21548 (N_21548,N_21181,N_21109);
nor U21549 (N_21549,N_20473,N_20964);
and U21550 (N_21550,N_20341,N_20114);
or U21551 (N_21551,N_20697,N_20931);
nor U21552 (N_21552,N_20682,N_20955);
nand U21553 (N_21553,N_20921,N_20640);
nor U21554 (N_21554,N_20816,N_20382);
nor U21555 (N_21555,N_20781,N_20685);
nor U21556 (N_21556,N_20780,N_20544);
or U21557 (N_21557,N_20019,N_20696);
xnor U21558 (N_21558,N_20784,N_20327);
nor U21559 (N_21559,N_20475,N_20812);
nor U21560 (N_21560,N_20079,N_21202);
nor U21561 (N_21561,N_20232,N_20705);
xor U21562 (N_21562,N_20451,N_20891);
or U21563 (N_21563,N_20102,N_20366);
nand U21564 (N_21564,N_20620,N_20160);
and U21565 (N_21565,N_20948,N_20522);
nand U21566 (N_21566,N_20311,N_20527);
nor U21567 (N_21567,N_20137,N_20798);
or U21568 (N_21568,N_20907,N_20467);
xor U21569 (N_21569,N_20455,N_21018);
nor U21570 (N_21570,N_20771,N_21074);
nand U21571 (N_21571,N_20458,N_20775);
nand U21572 (N_21572,N_20909,N_20726);
nand U21573 (N_21573,N_20028,N_21003);
or U21574 (N_21574,N_20940,N_20511);
nor U21575 (N_21575,N_20411,N_20846);
nor U21576 (N_21576,N_20861,N_20345);
xor U21577 (N_21577,N_20059,N_20122);
and U21578 (N_21578,N_21095,N_20038);
and U21579 (N_21579,N_20005,N_20099);
or U21580 (N_21580,N_20960,N_21149);
xor U21581 (N_21581,N_20139,N_20348);
xnor U21582 (N_21582,N_21106,N_20587);
nor U21583 (N_21583,N_20283,N_21024);
nor U21584 (N_21584,N_20765,N_20853);
nand U21585 (N_21585,N_21050,N_21145);
and U21586 (N_21586,N_20331,N_21015);
xnor U21587 (N_21587,N_21140,N_20581);
nand U21588 (N_21588,N_20979,N_20298);
xnor U21589 (N_21589,N_20113,N_20292);
or U21590 (N_21590,N_20313,N_20597);
xnor U21591 (N_21591,N_21226,N_20168);
nand U21592 (N_21592,N_20200,N_20499);
and U21593 (N_21593,N_20810,N_20566);
and U21594 (N_21594,N_20317,N_20665);
nor U21595 (N_21595,N_20159,N_20224);
nor U21596 (N_21596,N_20044,N_20599);
nand U21597 (N_21597,N_20596,N_20456);
and U21598 (N_21598,N_20125,N_20580);
and U21599 (N_21599,N_21201,N_20487);
nor U21600 (N_21600,N_21004,N_20198);
or U21601 (N_21601,N_20239,N_20171);
nor U21602 (N_21602,N_20605,N_20431);
xor U21603 (N_21603,N_21062,N_20967);
and U21604 (N_21604,N_20072,N_20154);
or U21605 (N_21605,N_20295,N_20664);
or U21606 (N_21606,N_20329,N_21028);
nand U21607 (N_21607,N_20518,N_20416);
or U21608 (N_21608,N_20659,N_20627);
or U21609 (N_21609,N_20138,N_20823);
nor U21610 (N_21610,N_20982,N_20121);
nor U21611 (N_21611,N_20418,N_20740);
and U21612 (N_21612,N_20369,N_20003);
or U21613 (N_21613,N_20755,N_20213);
and U21614 (N_21614,N_21148,N_21114);
nor U21615 (N_21615,N_20141,N_20928);
xor U21616 (N_21616,N_21022,N_20306);
xor U21617 (N_21617,N_20774,N_21217);
or U21618 (N_21618,N_20485,N_20434);
xnor U21619 (N_21619,N_20307,N_20737);
nand U21620 (N_21620,N_20554,N_20023);
nor U21621 (N_21621,N_20869,N_20770);
and U21622 (N_21622,N_20886,N_20305);
or U21623 (N_21623,N_20895,N_20851);
and U21624 (N_21624,N_20257,N_20673);
nand U21625 (N_21625,N_20654,N_20675);
nand U21626 (N_21626,N_20248,N_20427);
nand U21627 (N_21627,N_21002,N_20374);
xnor U21628 (N_21628,N_20548,N_20094);
xor U21629 (N_21629,N_21123,N_20108);
nand U21630 (N_21630,N_20083,N_20564);
or U21631 (N_21631,N_20373,N_20009);
nand U21632 (N_21632,N_20491,N_20389);
or U21633 (N_21633,N_20803,N_20438);
nand U21634 (N_21634,N_20797,N_21053);
or U21635 (N_21635,N_20132,N_20585);
xnor U21636 (N_21636,N_21080,N_20629);
nor U21637 (N_21637,N_20269,N_20284);
nand U21638 (N_21638,N_20515,N_21246);
xnor U21639 (N_21639,N_20616,N_20324);
or U21640 (N_21640,N_20681,N_21082);
nand U21641 (N_21641,N_20530,N_20896);
nor U21642 (N_21642,N_20147,N_20184);
and U21643 (N_21643,N_20857,N_20523);
xnor U21644 (N_21644,N_20902,N_20165);
nand U21645 (N_21645,N_20205,N_20572);
and U21646 (N_21646,N_20344,N_20365);
nor U21647 (N_21647,N_21083,N_20253);
nor U21648 (N_21648,N_20457,N_21061);
or U21649 (N_21649,N_20220,N_21029);
xor U21650 (N_21650,N_20030,N_21121);
xor U21651 (N_21651,N_20842,N_20927);
xnor U21652 (N_21652,N_20569,N_20501);
or U21653 (N_21653,N_20155,N_20503);
or U21654 (N_21654,N_20918,N_20057);
and U21655 (N_21655,N_20070,N_21171);
nor U21656 (N_21656,N_20219,N_20583);
nand U21657 (N_21657,N_20876,N_21020);
nor U21658 (N_21658,N_20553,N_20381);
or U21659 (N_21659,N_20984,N_20175);
xor U21660 (N_21660,N_20892,N_20022);
nor U21661 (N_21661,N_20466,N_21034);
nor U21662 (N_21662,N_20953,N_20603);
and U21663 (N_21663,N_20970,N_20399);
or U21664 (N_21664,N_20630,N_20012);
or U21665 (N_21665,N_20265,N_20176);
or U21666 (N_21666,N_21158,N_20063);
xnor U21667 (N_21667,N_20058,N_21193);
xnor U21668 (N_21668,N_20694,N_20971);
or U21669 (N_21669,N_20024,N_20223);
nor U21670 (N_21670,N_20371,N_21066);
nand U21671 (N_21671,N_20738,N_20293);
and U21672 (N_21672,N_20452,N_20648);
and U21673 (N_21673,N_20338,N_20925);
or U21674 (N_21674,N_20912,N_20556);
nor U21675 (N_21675,N_20252,N_20969);
nor U21676 (N_21676,N_21115,N_20259);
nor U21677 (N_21677,N_20368,N_21119);
nand U21678 (N_21678,N_20733,N_20312);
or U21679 (N_21679,N_21232,N_20577);
or U21680 (N_21680,N_20152,N_20550);
xor U21681 (N_21681,N_20300,N_20976);
and U21682 (N_21682,N_20481,N_21215);
nand U21683 (N_21683,N_20468,N_21178);
nand U21684 (N_21684,N_20144,N_21078);
or U21685 (N_21685,N_20706,N_20195);
nor U21686 (N_21686,N_21046,N_21089);
and U21687 (N_21687,N_20271,N_20815);
nand U21688 (N_21688,N_21210,N_20710);
nor U21689 (N_21689,N_20288,N_20881);
nand U21690 (N_21690,N_20649,N_20980);
nor U21691 (N_21691,N_20950,N_20516);
and U21692 (N_21692,N_20772,N_20877);
and U21693 (N_21693,N_20525,N_20534);
xor U21694 (N_21694,N_21072,N_20471);
and U21695 (N_21695,N_20519,N_20800);
xnor U21696 (N_21696,N_20233,N_20591);
nand U21697 (N_21697,N_21176,N_21189);
or U21698 (N_21698,N_21153,N_20678);
xnor U21699 (N_21699,N_20730,N_21025);
xnor U21700 (N_21700,N_21146,N_21044);
nor U21701 (N_21701,N_20169,N_20423);
and U21702 (N_21702,N_20683,N_20335);
nand U21703 (N_21703,N_20462,N_20562);
or U21704 (N_21704,N_20042,N_20163);
nor U21705 (N_21705,N_21060,N_20047);
or U21706 (N_21706,N_20197,N_20778);
nor U21707 (N_21707,N_20320,N_20477);
nand U21708 (N_21708,N_21143,N_20831);
nand U21709 (N_21709,N_21155,N_20748);
nand U21710 (N_21710,N_21139,N_20674);
nor U21711 (N_21711,N_21247,N_20474);
xor U21712 (N_21712,N_20695,N_20606);
xor U21713 (N_21713,N_20500,N_21021);
nand U21714 (N_21714,N_20036,N_20923);
and U21715 (N_21715,N_21125,N_21005);
nor U21716 (N_21716,N_21212,N_20570);
xnor U21717 (N_21717,N_20576,N_20050);
nand U21718 (N_21718,N_21031,N_20878);
and U21719 (N_21719,N_20041,N_20528);
or U21720 (N_21720,N_21128,N_21124);
xnor U21721 (N_21721,N_20879,N_20776);
or U21722 (N_21722,N_20075,N_20538);
or U21723 (N_21723,N_20670,N_20196);
xnor U21724 (N_21724,N_20558,N_21116);
nand U21725 (N_21725,N_20614,N_20403);
xnor U21726 (N_21726,N_20087,N_21188);
or U21727 (N_21727,N_20308,N_20517);
nor U21728 (N_21728,N_20889,N_20194);
or U21729 (N_21729,N_20910,N_21234);
nor U21730 (N_21730,N_20568,N_21190);
nand U21731 (N_21731,N_21057,N_20920);
nor U21732 (N_21732,N_21071,N_20020);
nand U21733 (N_21733,N_20181,N_21170);
nand U21734 (N_21734,N_20323,N_20917);
nand U21735 (N_21735,N_20565,N_21144);
and U21736 (N_21736,N_20991,N_20310);
xnor U21737 (N_21737,N_21169,N_20237);
nor U21738 (N_21738,N_20082,N_20459);
and U21739 (N_21739,N_20110,N_20941);
xnor U21740 (N_21740,N_20722,N_20793);
and U21741 (N_21741,N_20062,N_20820);
xor U21742 (N_21742,N_20858,N_20260);
nand U21743 (N_21743,N_21230,N_21152);
and U21744 (N_21744,N_20354,N_20520);
xor U21745 (N_21745,N_20792,N_20464);
xnor U21746 (N_21746,N_20025,N_20150);
xor U21747 (N_21747,N_21227,N_20994);
xnor U21748 (N_21748,N_20173,N_20667);
nand U21749 (N_21749,N_21200,N_20711);
nand U21750 (N_21750,N_20297,N_20914);
xnor U21751 (N_21751,N_20492,N_21122);
nand U21752 (N_21752,N_20004,N_20806);
nand U21753 (N_21753,N_20555,N_20107);
nor U21754 (N_21754,N_20055,N_20961);
nand U21755 (N_21755,N_20973,N_20926);
nor U21756 (N_21756,N_20240,N_21242);
or U21757 (N_21757,N_20111,N_20435);
nand U21758 (N_21758,N_21204,N_21192);
and U21759 (N_21759,N_20830,N_20071);
and U21760 (N_21760,N_21180,N_20454);
or U21761 (N_21761,N_20128,N_20868);
nand U21762 (N_21762,N_20336,N_20552);
or U21763 (N_21763,N_20713,N_20201);
and U21764 (N_21764,N_20643,N_20999);
nor U21765 (N_21765,N_20900,N_21157);
xnor U21766 (N_21766,N_20148,N_20415);
or U21767 (N_21767,N_20700,N_20080);
xor U21768 (N_21768,N_21041,N_21049);
nand U21769 (N_21769,N_21006,N_20093);
nor U21770 (N_21770,N_21087,N_20104);
nor U21771 (N_21771,N_21039,N_20533);
nor U21772 (N_21772,N_20592,N_20334);
xor U21773 (N_21773,N_20551,N_20180);
and U21774 (N_21774,N_20645,N_21012);
nor U21775 (N_21775,N_20699,N_20067);
nor U21776 (N_21776,N_20384,N_20098);
and U21777 (N_21777,N_20172,N_20814);
nor U21778 (N_21778,N_21019,N_20450);
and U21779 (N_21779,N_21076,N_20508);
nand U21780 (N_21780,N_20559,N_21244);
nand U21781 (N_21781,N_20421,N_21129);
xnor U21782 (N_21782,N_20216,N_20529);
or U21783 (N_21783,N_20720,N_20598);
nor U21784 (N_21784,N_21011,N_20767);
nor U21785 (N_21785,N_20993,N_21086);
nand U21786 (N_21786,N_20791,N_20263);
and U21787 (N_21787,N_21243,N_20378);
nand U21788 (N_21788,N_21032,N_21037);
or U21789 (N_21789,N_21220,N_20646);
xnor U21790 (N_21790,N_20754,N_21175);
or U21791 (N_21791,N_21056,N_20539);
xnor U21792 (N_21792,N_20796,N_20192);
nand U21793 (N_21793,N_20957,N_20496);
nor U21794 (N_21794,N_20206,N_21013);
nor U21795 (N_21795,N_20852,N_20393);
xor U21796 (N_21796,N_20655,N_20794);
or U21797 (N_21797,N_20179,N_20073);
xnor U21798 (N_21798,N_20162,N_20385);
and U21799 (N_21799,N_20864,N_20045);
xor U21800 (N_21800,N_20509,N_20143);
or U21801 (N_21801,N_20977,N_20048);
or U21802 (N_21802,N_20126,N_20470);
or U21803 (N_21803,N_20390,N_20911);
xnor U21804 (N_21804,N_21118,N_20352);
nor U21805 (N_21805,N_20088,N_20377);
nor U21806 (N_21806,N_20049,N_20882);
nand U21807 (N_21807,N_20234,N_20818);
nor U21808 (N_21808,N_20505,N_20262);
xor U21809 (N_21809,N_20051,N_20612);
or U21810 (N_21810,N_21211,N_20230);
or U21811 (N_21811,N_20942,N_20762);
or U21812 (N_21812,N_20081,N_20084);
nand U21813 (N_21813,N_20586,N_20358);
and U21814 (N_21814,N_20769,N_20611);
and U21815 (N_21815,N_20015,N_20930);
nand U21816 (N_21816,N_20677,N_20254);
nand U21817 (N_21817,N_20482,N_20359);
xnor U21818 (N_21818,N_21167,N_20752);
nor U21819 (N_21819,N_21014,N_20936);
nor U21820 (N_21820,N_20021,N_20595);
and U21821 (N_21821,N_21098,N_21229);
nand U21822 (N_21822,N_20294,N_20396);
xnor U21823 (N_21823,N_20441,N_20712);
nor U21824 (N_21824,N_20246,N_20185);
nor U21825 (N_21825,N_20347,N_20106);
nand U21826 (N_21826,N_21237,N_20285);
nor U21827 (N_21827,N_20625,N_20828);
nand U21828 (N_21828,N_20202,N_20480);
or U21829 (N_21829,N_20407,N_20484);
nand U21830 (N_21830,N_20140,N_21203);
or U21831 (N_21831,N_20750,N_20834);
nand U21832 (N_21832,N_20166,N_20915);
xnor U21833 (N_21833,N_20134,N_21104);
xor U21834 (N_21834,N_20636,N_20546);
xor U21835 (N_21835,N_20582,N_21045);
nor U21836 (N_21836,N_20731,N_20439);
nor U21837 (N_21837,N_20494,N_20296);
or U21838 (N_21838,N_21092,N_20425);
or U21839 (N_21839,N_20486,N_20289);
xnor U21840 (N_21840,N_20130,N_20183);
and U21841 (N_21841,N_20986,N_20845);
nor U21842 (N_21842,N_20905,N_20782);
and U21843 (N_21843,N_20264,N_21185);
and U21844 (N_21844,N_21091,N_20153);
and U21845 (N_21845,N_20656,N_20151);
xor U21846 (N_21846,N_20006,N_20124);
xor U21847 (N_21847,N_20333,N_20430);
nand U21848 (N_21848,N_21166,N_20557);
or U21849 (N_21849,N_20849,N_20037);
nand U21850 (N_21850,N_20032,N_20753);
nand U21851 (N_21851,N_20573,N_20256);
nor U21852 (N_21852,N_20395,N_20714);
nand U21853 (N_21853,N_20001,N_20756);
xnor U21854 (N_21854,N_20326,N_20349);
nand U21855 (N_21855,N_20115,N_20790);
nor U21856 (N_21856,N_21093,N_21194);
or U21857 (N_21857,N_20340,N_21134);
or U21858 (N_21858,N_20027,N_20567);
or U21859 (N_21859,N_20974,N_20178);
and U21860 (N_21860,N_20228,N_20117);
or U21861 (N_21861,N_20805,N_20367);
nand U21862 (N_21862,N_21240,N_20483);
xor U21863 (N_21863,N_20799,N_20146);
nand U21864 (N_21864,N_21000,N_21027);
nand U21865 (N_21865,N_20619,N_21070);
or U21866 (N_21866,N_21223,N_20628);
and U21867 (N_21867,N_20728,N_20136);
xnor U21868 (N_21868,N_21120,N_20521);
nor U21869 (N_21869,N_20893,N_20261);
xnor U21870 (N_21870,N_20417,N_20719);
xnor U21871 (N_21871,N_20406,N_20933);
and U21872 (N_21872,N_20225,N_20209);
and U21873 (N_21873,N_21195,N_20433);
or U21874 (N_21874,N_20064,N_21199);
nand U21875 (N_21875,N_20298,N_20972);
nor U21876 (N_21876,N_20088,N_20265);
nor U21877 (N_21877,N_20216,N_21011);
xor U21878 (N_21878,N_21019,N_20435);
and U21879 (N_21879,N_20523,N_20491);
nand U21880 (N_21880,N_20547,N_20962);
or U21881 (N_21881,N_21113,N_20519);
nand U21882 (N_21882,N_21245,N_20143);
and U21883 (N_21883,N_20714,N_20520);
and U21884 (N_21884,N_21019,N_20771);
and U21885 (N_21885,N_20518,N_20880);
or U21886 (N_21886,N_21247,N_20706);
and U21887 (N_21887,N_20524,N_20347);
or U21888 (N_21888,N_20721,N_21113);
nor U21889 (N_21889,N_21046,N_20861);
and U21890 (N_21890,N_20067,N_20960);
xnor U21891 (N_21891,N_21057,N_20265);
nand U21892 (N_21892,N_20119,N_20253);
nand U21893 (N_21893,N_20694,N_20623);
xor U21894 (N_21894,N_21202,N_20045);
nand U21895 (N_21895,N_20714,N_21040);
xor U21896 (N_21896,N_20719,N_20234);
and U21897 (N_21897,N_20160,N_20302);
nand U21898 (N_21898,N_20732,N_20049);
nand U21899 (N_21899,N_20408,N_20250);
xor U21900 (N_21900,N_20863,N_20658);
and U21901 (N_21901,N_21240,N_20777);
nor U21902 (N_21902,N_20079,N_20179);
xnor U21903 (N_21903,N_20810,N_20273);
xor U21904 (N_21904,N_20779,N_20487);
nor U21905 (N_21905,N_20660,N_21152);
nand U21906 (N_21906,N_20221,N_20448);
or U21907 (N_21907,N_20287,N_21199);
and U21908 (N_21908,N_20566,N_21214);
xor U21909 (N_21909,N_20030,N_20693);
nor U21910 (N_21910,N_20069,N_21130);
nor U21911 (N_21911,N_21207,N_20117);
nand U21912 (N_21912,N_20378,N_20148);
and U21913 (N_21913,N_20457,N_20131);
or U21914 (N_21914,N_20760,N_20615);
and U21915 (N_21915,N_21207,N_20181);
nor U21916 (N_21916,N_21069,N_21013);
or U21917 (N_21917,N_20773,N_20482);
and U21918 (N_21918,N_21134,N_20634);
and U21919 (N_21919,N_21069,N_20071);
nand U21920 (N_21920,N_20378,N_20542);
or U21921 (N_21921,N_20862,N_20898);
nand U21922 (N_21922,N_21231,N_20021);
nand U21923 (N_21923,N_20969,N_21069);
or U21924 (N_21924,N_20275,N_20805);
or U21925 (N_21925,N_20229,N_20077);
or U21926 (N_21926,N_20636,N_20226);
or U21927 (N_21927,N_21164,N_20119);
xor U21928 (N_21928,N_20209,N_20547);
and U21929 (N_21929,N_20598,N_20276);
and U21930 (N_21930,N_20594,N_20060);
and U21931 (N_21931,N_20050,N_20199);
nor U21932 (N_21932,N_20731,N_20706);
nand U21933 (N_21933,N_21157,N_20912);
and U21934 (N_21934,N_20069,N_20541);
nand U21935 (N_21935,N_21144,N_21028);
xnor U21936 (N_21936,N_20137,N_20311);
or U21937 (N_21937,N_21240,N_20708);
nand U21938 (N_21938,N_20346,N_20247);
and U21939 (N_21939,N_20477,N_20403);
xnor U21940 (N_21940,N_21107,N_21236);
or U21941 (N_21941,N_20853,N_21025);
and U21942 (N_21942,N_21193,N_20639);
and U21943 (N_21943,N_20293,N_20812);
nand U21944 (N_21944,N_20664,N_21213);
xor U21945 (N_21945,N_21013,N_20945);
and U21946 (N_21946,N_20425,N_20052);
nor U21947 (N_21947,N_20188,N_20610);
or U21948 (N_21948,N_20036,N_20429);
and U21949 (N_21949,N_20555,N_20539);
nand U21950 (N_21950,N_20420,N_20861);
nor U21951 (N_21951,N_20753,N_20891);
nand U21952 (N_21952,N_20846,N_20378);
xor U21953 (N_21953,N_21180,N_20241);
or U21954 (N_21954,N_21233,N_20908);
nor U21955 (N_21955,N_20594,N_21172);
and U21956 (N_21956,N_20155,N_20169);
nor U21957 (N_21957,N_20235,N_20603);
xor U21958 (N_21958,N_20289,N_21231);
and U21959 (N_21959,N_20302,N_21243);
and U21960 (N_21960,N_20965,N_20062);
xnor U21961 (N_21961,N_20713,N_20042);
nand U21962 (N_21962,N_20470,N_21131);
xor U21963 (N_21963,N_20356,N_20739);
or U21964 (N_21964,N_20275,N_20009);
or U21965 (N_21965,N_20882,N_20607);
xnor U21966 (N_21966,N_20806,N_20849);
nor U21967 (N_21967,N_20564,N_20609);
nor U21968 (N_21968,N_20459,N_21241);
nor U21969 (N_21969,N_20636,N_20980);
or U21970 (N_21970,N_21151,N_20728);
or U21971 (N_21971,N_20415,N_20629);
nand U21972 (N_21972,N_20838,N_20287);
xnor U21973 (N_21973,N_21141,N_20190);
nor U21974 (N_21974,N_21239,N_20981);
xor U21975 (N_21975,N_20052,N_21222);
and U21976 (N_21976,N_21119,N_20770);
nor U21977 (N_21977,N_20029,N_20737);
or U21978 (N_21978,N_20708,N_21156);
xor U21979 (N_21979,N_20658,N_20840);
nand U21980 (N_21980,N_20485,N_21085);
nand U21981 (N_21981,N_21231,N_20570);
and U21982 (N_21982,N_20348,N_21086);
nand U21983 (N_21983,N_20671,N_20897);
and U21984 (N_21984,N_20739,N_20246);
or U21985 (N_21985,N_20290,N_21147);
nor U21986 (N_21986,N_21156,N_20131);
nand U21987 (N_21987,N_20710,N_21131);
nand U21988 (N_21988,N_20618,N_20508);
nand U21989 (N_21989,N_20310,N_20534);
nand U21990 (N_21990,N_20276,N_20887);
xnor U21991 (N_21991,N_20070,N_20518);
or U21992 (N_21992,N_20661,N_20428);
and U21993 (N_21993,N_20277,N_20795);
and U21994 (N_21994,N_20595,N_21015);
or U21995 (N_21995,N_20363,N_20725);
and U21996 (N_21996,N_20601,N_20989);
and U21997 (N_21997,N_20735,N_20138);
and U21998 (N_21998,N_20422,N_20746);
nand U21999 (N_21999,N_20106,N_20586);
or U22000 (N_22000,N_20038,N_21056);
or U22001 (N_22001,N_20319,N_20984);
nand U22002 (N_22002,N_20617,N_20479);
or U22003 (N_22003,N_20964,N_20922);
or U22004 (N_22004,N_20676,N_20271);
xnor U22005 (N_22005,N_20720,N_20345);
nand U22006 (N_22006,N_20325,N_20843);
nor U22007 (N_22007,N_20048,N_20841);
xnor U22008 (N_22008,N_20421,N_20528);
xor U22009 (N_22009,N_21182,N_20687);
or U22010 (N_22010,N_20009,N_20861);
nor U22011 (N_22011,N_20040,N_20564);
and U22012 (N_22012,N_20046,N_20948);
nand U22013 (N_22013,N_20612,N_20163);
xnor U22014 (N_22014,N_20539,N_20241);
or U22015 (N_22015,N_20153,N_20746);
xnor U22016 (N_22016,N_21038,N_20967);
and U22017 (N_22017,N_20447,N_20032);
nand U22018 (N_22018,N_20305,N_20401);
xnor U22019 (N_22019,N_20637,N_20821);
and U22020 (N_22020,N_20831,N_20187);
and U22021 (N_22021,N_21134,N_21142);
or U22022 (N_22022,N_21092,N_20061);
and U22023 (N_22023,N_20773,N_20422);
nor U22024 (N_22024,N_20733,N_21041);
and U22025 (N_22025,N_20200,N_20273);
nand U22026 (N_22026,N_20549,N_20880);
or U22027 (N_22027,N_20861,N_21028);
and U22028 (N_22028,N_20025,N_20037);
and U22029 (N_22029,N_20324,N_21013);
and U22030 (N_22030,N_20624,N_20481);
or U22031 (N_22031,N_20302,N_20802);
nor U22032 (N_22032,N_21211,N_20473);
xnor U22033 (N_22033,N_20262,N_21122);
nor U22034 (N_22034,N_20674,N_20305);
nor U22035 (N_22035,N_21102,N_20671);
xnor U22036 (N_22036,N_20883,N_20389);
nor U22037 (N_22037,N_20175,N_20822);
nor U22038 (N_22038,N_20674,N_20777);
nor U22039 (N_22039,N_20550,N_20336);
xor U22040 (N_22040,N_21109,N_20422);
or U22041 (N_22041,N_21087,N_20475);
or U22042 (N_22042,N_20298,N_20389);
and U22043 (N_22043,N_20819,N_20082);
xnor U22044 (N_22044,N_20584,N_20324);
nand U22045 (N_22045,N_21199,N_20114);
xnor U22046 (N_22046,N_20644,N_21163);
xor U22047 (N_22047,N_20097,N_20107);
or U22048 (N_22048,N_20843,N_20758);
nand U22049 (N_22049,N_20694,N_21155);
and U22050 (N_22050,N_20173,N_21104);
nand U22051 (N_22051,N_20930,N_20438);
nor U22052 (N_22052,N_20775,N_20590);
and U22053 (N_22053,N_20664,N_21201);
nor U22054 (N_22054,N_21169,N_20555);
nor U22055 (N_22055,N_20041,N_20004);
nand U22056 (N_22056,N_20683,N_20344);
nand U22057 (N_22057,N_21246,N_20828);
xor U22058 (N_22058,N_20959,N_20564);
or U22059 (N_22059,N_20485,N_21045);
and U22060 (N_22060,N_20703,N_21026);
nand U22061 (N_22061,N_20994,N_21048);
xnor U22062 (N_22062,N_20250,N_20935);
or U22063 (N_22063,N_20098,N_21169);
nand U22064 (N_22064,N_20854,N_20176);
nor U22065 (N_22065,N_20352,N_20318);
nand U22066 (N_22066,N_20943,N_20950);
xnor U22067 (N_22067,N_20810,N_20463);
nand U22068 (N_22068,N_20857,N_21060);
nand U22069 (N_22069,N_20208,N_20413);
xor U22070 (N_22070,N_20465,N_20295);
and U22071 (N_22071,N_20761,N_20668);
nand U22072 (N_22072,N_20289,N_21097);
and U22073 (N_22073,N_20557,N_20778);
nor U22074 (N_22074,N_20212,N_20219);
and U22075 (N_22075,N_20085,N_21107);
and U22076 (N_22076,N_20662,N_20944);
xnor U22077 (N_22077,N_21025,N_20412);
nand U22078 (N_22078,N_20610,N_20042);
xor U22079 (N_22079,N_20866,N_20481);
xor U22080 (N_22080,N_21102,N_20158);
or U22081 (N_22081,N_20229,N_21177);
and U22082 (N_22082,N_20395,N_21109);
nor U22083 (N_22083,N_20105,N_21242);
or U22084 (N_22084,N_20881,N_21125);
or U22085 (N_22085,N_21021,N_20419);
nor U22086 (N_22086,N_20683,N_20557);
or U22087 (N_22087,N_20889,N_20187);
and U22088 (N_22088,N_21192,N_20126);
and U22089 (N_22089,N_20334,N_20891);
xor U22090 (N_22090,N_21129,N_20670);
and U22091 (N_22091,N_20634,N_21183);
xnor U22092 (N_22092,N_20117,N_21008);
or U22093 (N_22093,N_20940,N_20011);
nand U22094 (N_22094,N_20781,N_21048);
and U22095 (N_22095,N_20179,N_20676);
and U22096 (N_22096,N_20583,N_21004);
and U22097 (N_22097,N_20793,N_20648);
or U22098 (N_22098,N_21224,N_20047);
or U22099 (N_22099,N_20228,N_20313);
nor U22100 (N_22100,N_20330,N_20471);
nand U22101 (N_22101,N_20395,N_20000);
nand U22102 (N_22102,N_20567,N_21163);
nand U22103 (N_22103,N_21001,N_21247);
nand U22104 (N_22104,N_21009,N_20910);
nand U22105 (N_22105,N_20892,N_20176);
or U22106 (N_22106,N_20338,N_21116);
xnor U22107 (N_22107,N_20366,N_20589);
nand U22108 (N_22108,N_20786,N_20471);
xor U22109 (N_22109,N_20814,N_20893);
or U22110 (N_22110,N_20534,N_20921);
nor U22111 (N_22111,N_20254,N_20044);
and U22112 (N_22112,N_20698,N_20266);
nor U22113 (N_22113,N_20964,N_20655);
xor U22114 (N_22114,N_20232,N_21243);
and U22115 (N_22115,N_20889,N_20887);
nor U22116 (N_22116,N_20993,N_20011);
and U22117 (N_22117,N_20759,N_20704);
xor U22118 (N_22118,N_20964,N_20861);
nand U22119 (N_22119,N_20220,N_20975);
and U22120 (N_22120,N_20287,N_21014);
nor U22121 (N_22121,N_20052,N_20614);
nor U22122 (N_22122,N_20052,N_20302);
nor U22123 (N_22123,N_20695,N_20297);
or U22124 (N_22124,N_20567,N_20261);
xor U22125 (N_22125,N_20489,N_20417);
or U22126 (N_22126,N_21145,N_20969);
xnor U22127 (N_22127,N_21025,N_20519);
xnor U22128 (N_22128,N_20605,N_21069);
xnor U22129 (N_22129,N_21227,N_20156);
and U22130 (N_22130,N_20122,N_20931);
nand U22131 (N_22131,N_20692,N_20846);
and U22132 (N_22132,N_20192,N_21114);
or U22133 (N_22133,N_20665,N_20867);
and U22134 (N_22134,N_20896,N_21045);
or U22135 (N_22135,N_21157,N_20757);
nor U22136 (N_22136,N_20483,N_20264);
and U22137 (N_22137,N_20758,N_20483);
xor U22138 (N_22138,N_20165,N_20390);
xnor U22139 (N_22139,N_20981,N_20890);
or U22140 (N_22140,N_20940,N_21060);
and U22141 (N_22141,N_20459,N_20817);
nor U22142 (N_22142,N_21124,N_20324);
nand U22143 (N_22143,N_20013,N_20952);
xnor U22144 (N_22144,N_20919,N_20979);
and U22145 (N_22145,N_20392,N_20929);
nand U22146 (N_22146,N_21055,N_20030);
nor U22147 (N_22147,N_20473,N_20458);
nand U22148 (N_22148,N_20523,N_20020);
nor U22149 (N_22149,N_20527,N_21068);
xnor U22150 (N_22150,N_20602,N_20247);
xor U22151 (N_22151,N_20369,N_20995);
xnor U22152 (N_22152,N_20319,N_20522);
and U22153 (N_22153,N_20937,N_20635);
or U22154 (N_22154,N_21232,N_20162);
and U22155 (N_22155,N_20991,N_20553);
nor U22156 (N_22156,N_20468,N_20319);
or U22157 (N_22157,N_20021,N_20213);
xnor U22158 (N_22158,N_20432,N_20561);
nand U22159 (N_22159,N_20761,N_21196);
and U22160 (N_22160,N_21073,N_20868);
and U22161 (N_22161,N_20019,N_20618);
and U22162 (N_22162,N_20533,N_20557);
or U22163 (N_22163,N_20476,N_21010);
nor U22164 (N_22164,N_20374,N_20813);
and U22165 (N_22165,N_20950,N_20169);
xor U22166 (N_22166,N_21075,N_20245);
xor U22167 (N_22167,N_20008,N_20530);
nand U22168 (N_22168,N_20525,N_20376);
xor U22169 (N_22169,N_20264,N_20110);
and U22170 (N_22170,N_20642,N_21185);
and U22171 (N_22171,N_20344,N_20425);
nor U22172 (N_22172,N_20051,N_20814);
nor U22173 (N_22173,N_20107,N_20931);
nor U22174 (N_22174,N_20832,N_20982);
xnor U22175 (N_22175,N_20634,N_20476);
or U22176 (N_22176,N_20994,N_21037);
nor U22177 (N_22177,N_20979,N_21081);
nor U22178 (N_22178,N_20979,N_20923);
nand U22179 (N_22179,N_20717,N_20451);
nand U22180 (N_22180,N_20139,N_20820);
and U22181 (N_22181,N_20459,N_20535);
or U22182 (N_22182,N_21154,N_20047);
and U22183 (N_22183,N_20519,N_20103);
nor U22184 (N_22184,N_20879,N_20545);
or U22185 (N_22185,N_20250,N_21067);
or U22186 (N_22186,N_20390,N_20371);
xor U22187 (N_22187,N_20644,N_21091);
nand U22188 (N_22188,N_20396,N_21231);
or U22189 (N_22189,N_20511,N_20734);
nor U22190 (N_22190,N_20776,N_20241);
or U22191 (N_22191,N_20843,N_20237);
and U22192 (N_22192,N_20881,N_21169);
or U22193 (N_22193,N_21225,N_20808);
xnor U22194 (N_22194,N_20500,N_20145);
or U22195 (N_22195,N_20473,N_21177);
nand U22196 (N_22196,N_21004,N_20842);
and U22197 (N_22197,N_20400,N_20441);
and U22198 (N_22198,N_20879,N_20257);
nor U22199 (N_22199,N_20114,N_20535);
nor U22200 (N_22200,N_20899,N_21173);
and U22201 (N_22201,N_20893,N_21068);
nand U22202 (N_22202,N_20722,N_20201);
and U22203 (N_22203,N_20688,N_21039);
xor U22204 (N_22204,N_20743,N_20128);
or U22205 (N_22205,N_20384,N_20673);
or U22206 (N_22206,N_20832,N_20105);
xnor U22207 (N_22207,N_20750,N_20956);
or U22208 (N_22208,N_20477,N_20641);
xor U22209 (N_22209,N_20472,N_20680);
nor U22210 (N_22210,N_20691,N_20177);
or U22211 (N_22211,N_20199,N_20891);
xnor U22212 (N_22212,N_20499,N_20371);
xor U22213 (N_22213,N_20944,N_20693);
and U22214 (N_22214,N_20943,N_20208);
nor U22215 (N_22215,N_21094,N_21158);
xnor U22216 (N_22216,N_21234,N_20280);
xnor U22217 (N_22217,N_20631,N_20689);
nand U22218 (N_22218,N_21085,N_21155);
xor U22219 (N_22219,N_20485,N_20914);
and U22220 (N_22220,N_20455,N_20145);
xnor U22221 (N_22221,N_20272,N_20350);
nand U22222 (N_22222,N_20342,N_21172);
or U22223 (N_22223,N_20268,N_20328);
and U22224 (N_22224,N_20989,N_21225);
xor U22225 (N_22225,N_20350,N_21077);
or U22226 (N_22226,N_20066,N_20165);
or U22227 (N_22227,N_21206,N_21161);
and U22228 (N_22228,N_20372,N_20401);
nand U22229 (N_22229,N_20523,N_20468);
and U22230 (N_22230,N_20651,N_20055);
and U22231 (N_22231,N_20183,N_21105);
nor U22232 (N_22232,N_20499,N_20344);
xnor U22233 (N_22233,N_20236,N_21124);
xnor U22234 (N_22234,N_20103,N_21094);
nand U22235 (N_22235,N_20445,N_21058);
and U22236 (N_22236,N_20136,N_20407);
nor U22237 (N_22237,N_21008,N_20535);
and U22238 (N_22238,N_20256,N_20232);
or U22239 (N_22239,N_20752,N_20136);
xnor U22240 (N_22240,N_20421,N_20346);
xnor U22241 (N_22241,N_21017,N_20208);
or U22242 (N_22242,N_21030,N_20221);
nor U22243 (N_22243,N_21160,N_21071);
nand U22244 (N_22244,N_20542,N_20289);
and U22245 (N_22245,N_20047,N_20399);
and U22246 (N_22246,N_20920,N_20530);
and U22247 (N_22247,N_20129,N_20968);
or U22248 (N_22248,N_20441,N_20904);
xor U22249 (N_22249,N_20842,N_20065);
and U22250 (N_22250,N_20469,N_21096);
and U22251 (N_22251,N_20742,N_20260);
and U22252 (N_22252,N_21169,N_20872);
or U22253 (N_22253,N_20932,N_20036);
xnor U22254 (N_22254,N_21141,N_20647);
and U22255 (N_22255,N_20831,N_20708);
or U22256 (N_22256,N_20543,N_21073);
or U22257 (N_22257,N_20209,N_20501);
or U22258 (N_22258,N_20556,N_20722);
nor U22259 (N_22259,N_20084,N_20835);
nand U22260 (N_22260,N_20013,N_20141);
or U22261 (N_22261,N_20383,N_20055);
nand U22262 (N_22262,N_20377,N_20271);
or U22263 (N_22263,N_20601,N_20546);
and U22264 (N_22264,N_21049,N_20966);
nand U22265 (N_22265,N_20930,N_20149);
xor U22266 (N_22266,N_20980,N_20240);
xnor U22267 (N_22267,N_20000,N_21114);
nand U22268 (N_22268,N_20543,N_20019);
nor U22269 (N_22269,N_20188,N_20687);
nor U22270 (N_22270,N_20967,N_20716);
nand U22271 (N_22271,N_21208,N_20485);
nor U22272 (N_22272,N_21152,N_20868);
nor U22273 (N_22273,N_20587,N_20426);
nand U22274 (N_22274,N_20276,N_20078);
xor U22275 (N_22275,N_20297,N_20404);
nand U22276 (N_22276,N_20741,N_20671);
nor U22277 (N_22277,N_20885,N_20477);
xnor U22278 (N_22278,N_20238,N_20574);
and U22279 (N_22279,N_20233,N_20603);
and U22280 (N_22280,N_20340,N_20846);
or U22281 (N_22281,N_20498,N_20802);
nor U22282 (N_22282,N_20022,N_20555);
xnor U22283 (N_22283,N_20529,N_20428);
or U22284 (N_22284,N_20050,N_20755);
and U22285 (N_22285,N_21230,N_20658);
xnor U22286 (N_22286,N_20179,N_20917);
nor U22287 (N_22287,N_21211,N_20643);
nor U22288 (N_22288,N_20351,N_21190);
or U22289 (N_22289,N_20202,N_20239);
nand U22290 (N_22290,N_20932,N_20438);
nand U22291 (N_22291,N_20662,N_20603);
nor U22292 (N_22292,N_20989,N_20869);
and U22293 (N_22293,N_20429,N_20515);
nand U22294 (N_22294,N_20192,N_20147);
nand U22295 (N_22295,N_20341,N_20134);
nor U22296 (N_22296,N_20952,N_20722);
or U22297 (N_22297,N_20613,N_20033);
and U22298 (N_22298,N_20139,N_20075);
or U22299 (N_22299,N_20883,N_21233);
xor U22300 (N_22300,N_20678,N_21119);
nor U22301 (N_22301,N_20099,N_21113);
xnor U22302 (N_22302,N_20276,N_20839);
xor U22303 (N_22303,N_21055,N_20330);
nand U22304 (N_22304,N_20282,N_20823);
nand U22305 (N_22305,N_20249,N_20257);
xor U22306 (N_22306,N_20590,N_20159);
nand U22307 (N_22307,N_20201,N_20508);
xnor U22308 (N_22308,N_20795,N_21142);
xor U22309 (N_22309,N_20159,N_20850);
or U22310 (N_22310,N_21200,N_20302);
or U22311 (N_22311,N_20731,N_20211);
or U22312 (N_22312,N_20106,N_20899);
nand U22313 (N_22313,N_20871,N_20186);
nor U22314 (N_22314,N_20520,N_20482);
xnor U22315 (N_22315,N_20698,N_20396);
xnor U22316 (N_22316,N_20704,N_20492);
nor U22317 (N_22317,N_21137,N_20077);
nand U22318 (N_22318,N_20178,N_21059);
xnor U22319 (N_22319,N_21150,N_20325);
and U22320 (N_22320,N_20435,N_21062);
and U22321 (N_22321,N_20784,N_20105);
nand U22322 (N_22322,N_21069,N_20213);
or U22323 (N_22323,N_20999,N_20655);
nand U22324 (N_22324,N_20194,N_20706);
nor U22325 (N_22325,N_21107,N_20700);
nor U22326 (N_22326,N_20650,N_20141);
nand U22327 (N_22327,N_20281,N_21154);
nand U22328 (N_22328,N_21049,N_20911);
and U22329 (N_22329,N_20641,N_20582);
nor U22330 (N_22330,N_20869,N_21078);
or U22331 (N_22331,N_20056,N_20486);
nor U22332 (N_22332,N_20594,N_20278);
or U22333 (N_22333,N_21055,N_20258);
nor U22334 (N_22334,N_20695,N_20895);
nand U22335 (N_22335,N_20174,N_20973);
nand U22336 (N_22336,N_20435,N_21204);
nand U22337 (N_22337,N_20546,N_20418);
nand U22338 (N_22338,N_20145,N_21001);
or U22339 (N_22339,N_20310,N_21202);
xor U22340 (N_22340,N_21180,N_20024);
nand U22341 (N_22341,N_20698,N_20338);
nor U22342 (N_22342,N_20411,N_20175);
nand U22343 (N_22343,N_21198,N_21210);
or U22344 (N_22344,N_20178,N_21080);
xor U22345 (N_22345,N_20537,N_20920);
and U22346 (N_22346,N_20934,N_20909);
xor U22347 (N_22347,N_20386,N_20126);
nand U22348 (N_22348,N_20351,N_20080);
and U22349 (N_22349,N_20468,N_20124);
nand U22350 (N_22350,N_21085,N_20131);
nor U22351 (N_22351,N_20271,N_21140);
xor U22352 (N_22352,N_20287,N_21021);
nor U22353 (N_22353,N_21046,N_20609);
xnor U22354 (N_22354,N_20700,N_21156);
or U22355 (N_22355,N_20264,N_20169);
xnor U22356 (N_22356,N_20276,N_20282);
xor U22357 (N_22357,N_20640,N_20444);
nand U22358 (N_22358,N_21161,N_21046);
and U22359 (N_22359,N_20617,N_21188);
or U22360 (N_22360,N_20707,N_20596);
nand U22361 (N_22361,N_20164,N_20201);
nor U22362 (N_22362,N_20939,N_20431);
or U22363 (N_22363,N_20801,N_20035);
nor U22364 (N_22364,N_21101,N_20426);
or U22365 (N_22365,N_21170,N_20526);
nor U22366 (N_22366,N_20056,N_20987);
xor U22367 (N_22367,N_20590,N_20567);
nand U22368 (N_22368,N_20391,N_20451);
xnor U22369 (N_22369,N_20831,N_20926);
or U22370 (N_22370,N_20731,N_21143);
xor U22371 (N_22371,N_20418,N_20108);
nand U22372 (N_22372,N_20647,N_20645);
or U22373 (N_22373,N_20183,N_21209);
or U22374 (N_22374,N_21070,N_20970);
nand U22375 (N_22375,N_20975,N_20310);
or U22376 (N_22376,N_20917,N_20060);
xor U22377 (N_22377,N_20420,N_20680);
or U22378 (N_22378,N_20246,N_21215);
xnor U22379 (N_22379,N_20872,N_20301);
or U22380 (N_22380,N_20459,N_20772);
or U22381 (N_22381,N_20749,N_21084);
nor U22382 (N_22382,N_21196,N_20755);
xor U22383 (N_22383,N_20135,N_20660);
or U22384 (N_22384,N_20801,N_20334);
nor U22385 (N_22385,N_20253,N_20878);
nand U22386 (N_22386,N_21025,N_20570);
nor U22387 (N_22387,N_21098,N_20453);
or U22388 (N_22388,N_20865,N_20825);
xnor U22389 (N_22389,N_20464,N_20123);
and U22390 (N_22390,N_20510,N_20676);
nand U22391 (N_22391,N_21038,N_20944);
xor U22392 (N_22392,N_20675,N_20818);
nor U22393 (N_22393,N_20064,N_20803);
and U22394 (N_22394,N_20199,N_20606);
nand U22395 (N_22395,N_20991,N_20168);
xor U22396 (N_22396,N_20803,N_20167);
nand U22397 (N_22397,N_20045,N_21087);
and U22398 (N_22398,N_20254,N_20433);
or U22399 (N_22399,N_20757,N_20422);
xor U22400 (N_22400,N_20507,N_20655);
or U22401 (N_22401,N_20667,N_20790);
xnor U22402 (N_22402,N_20222,N_20932);
xnor U22403 (N_22403,N_20123,N_20004);
or U22404 (N_22404,N_20482,N_20657);
or U22405 (N_22405,N_20982,N_20517);
and U22406 (N_22406,N_20747,N_20021);
nand U22407 (N_22407,N_20174,N_20316);
and U22408 (N_22408,N_20924,N_20574);
xor U22409 (N_22409,N_20668,N_20570);
and U22410 (N_22410,N_21175,N_20030);
nor U22411 (N_22411,N_20939,N_21179);
nand U22412 (N_22412,N_20788,N_20474);
nand U22413 (N_22413,N_20344,N_21229);
or U22414 (N_22414,N_20504,N_20840);
xnor U22415 (N_22415,N_20962,N_20412);
or U22416 (N_22416,N_20785,N_20517);
nor U22417 (N_22417,N_20225,N_21164);
or U22418 (N_22418,N_20504,N_20373);
xnor U22419 (N_22419,N_20660,N_20068);
and U22420 (N_22420,N_20555,N_20809);
nor U22421 (N_22421,N_20774,N_20975);
and U22422 (N_22422,N_20080,N_21129);
xor U22423 (N_22423,N_20257,N_20965);
or U22424 (N_22424,N_20475,N_20410);
nor U22425 (N_22425,N_20762,N_20008);
xor U22426 (N_22426,N_20562,N_20457);
or U22427 (N_22427,N_21120,N_20370);
xnor U22428 (N_22428,N_21214,N_20500);
nor U22429 (N_22429,N_20559,N_20011);
or U22430 (N_22430,N_20033,N_20369);
and U22431 (N_22431,N_20830,N_21093);
nand U22432 (N_22432,N_20467,N_20022);
and U22433 (N_22433,N_20851,N_20226);
and U22434 (N_22434,N_20844,N_20233);
or U22435 (N_22435,N_21015,N_20976);
xnor U22436 (N_22436,N_20298,N_20316);
or U22437 (N_22437,N_21059,N_21166);
or U22438 (N_22438,N_21109,N_20404);
nand U22439 (N_22439,N_20232,N_20978);
nor U22440 (N_22440,N_20960,N_20537);
and U22441 (N_22441,N_20467,N_20870);
xor U22442 (N_22442,N_20259,N_20684);
and U22443 (N_22443,N_20750,N_20661);
nand U22444 (N_22444,N_20550,N_20775);
nor U22445 (N_22445,N_20392,N_20087);
nand U22446 (N_22446,N_20244,N_20357);
xor U22447 (N_22447,N_20733,N_20154);
xnor U22448 (N_22448,N_20970,N_20178);
nand U22449 (N_22449,N_20979,N_20718);
nor U22450 (N_22450,N_21054,N_20102);
or U22451 (N_22451,N_20776,N_20075);
and U22452 (N_22452,N_21081,N_21196);
and U22453 (N_22453,N_20030,N_20595);
xor U22454 (N_22454,N_21073,N_20080);
xnor U22455 (N_22455,N_20221,N_21152);
nor U22456 (N_22456,N_20929,N_20919);
and U22457 (N_22457,N_20072,N_20018);
and U22458 (N_22458,N_20161,N_20169);
or U22459 (N_22459,N_20612,N_20746);
xnor U22460 (N_22460,N_20965,N_20220);
nand U22461 (N_22461,N_21173,N_20435);
xnor U22462 (N_22462,N_21086,N_20114);
xnor U22463 (N_22463,N_20023,N_20031);
nor U22464 (N_22464,N_20588,N_20412);
and U22465 (N_22465,N_20682,N_20099);
nor U22466 (N_22466,N_21172,N_21177);
and U22467 (N_22467,N_20193,N_20698);
nand U22468 (N_22468,N_21186,N_20973);
nand U22469 (N_22469,N_20319,N_20374);
nor U22470 (N_22470,N_20075,N_20991);
nand U22471 (N_22471,N_20274,N_20190);
xor U22472 (N_22472,N_20179,N_20844);
and U22473 (N_22473,N_21171,N_20312);
nor U22474 (N_22474,N_20707,N_20453);
or U22475 (N_22475,N_20997,N_21232);
or U22476 (N_22476,N_20883,N_20775);
and U22477 (N_22477,N_20606,N_20146);
and U22478 (N_22478,N_20289,N_20680);
and U22479 (N_22479,N_20762,N_21021);
and U22480 (N_22480,N_20131,N_21225);
nand U22481 (N_22481,N_20862,N_20766);
nor U22482 (N_22482,N_21066,N_20655);
xnor U22483 (N_22483,N_20374,N_20242);
nor U22484 (N_22484,N_20191,N_20682);
or U22485 (N_22485,N_20998,N_20847);
and U22486 (N_22486,N_20971,N_20859);
and U22487 (N_22487,N_20324,N_20759);
nor U22488 (N_22488,N_20746,N_20605);
nor U22489 (N_22489,N_20033,N_20845);
xor U22490 (N_22490,N_20503,N_21094);
nor U22491 (N_22491,N_21229,N_21245);
xor U22492 (N_22492,N_20084,N_20802);
xnor U22493 (N_22493,N_20991,N_20558);
xor U22494 (N_22494,N_20515,N_20258);
and U22495 (N_22495,N_20385,N_20187);
nand U22496 (N_22496,N_21111,N_20607);
nand U22497 (N_22497,N_20378,N_20917);
nand U22498 (N_22498,N_20599,N_20869);
and U22499 (N_22499,N_20425,N_20322);
nor U22500 (N_22500,N_21535,N_21667);
and U22501 (N_22501,N_22216,N_22222);
xnor U22502 (N_22502,N_22427,N_22358);
nor U22503 (N_22503,N_21605,N_22303);
xnor U22504 (N_22504,N_21959,N_21522);
or U22505 (N_22505,N_21969,N_21483);
nor U22506 (N_22506,N_22212,N_22025);
nor U22507 (N_22507,N_21830,N_21364);
and U22508 (N_22508,N_21986,N_21611);
nor U22509 (N_22509,N_21351,N_21271);
nor U22510 (N_22510,N_21337,N_21454);
nand U22511 (N_22511,N_21948,N_21903);
nand U22512 (N_22512,N_21938,N_21550);
nor U22513 (N_22513,N_22257,N_21593);
xor U22514 (N_22514,N_21877,N_21459);
and U22515 (N_22515,N_21477,N_21915);
nand U22516 (N_22516,N_21353,N_22041);
nor U22517 (N_22517,N_21523,N_21625);
xor U22518 (N_22518,N_21272,N_21510);
nand U22519 (N_22519,N_22274,N_21651);
nand U22520 (N_22520,N_21398,N_21416);
nand U22521 (N_22521,N_22142,N_21842);
nor U22522 (N_22522,N_21331,N_22400);
nor U22523 (N_22523,N_21414,N_21812);
and U22524 (N_22524,N_22035,N_22316);
nand U22525 (N_22525,N_21970,N_22136);
xor U22526 (N_22526,N_21860,N_21530);
and U22527 (N_22527,N_22218,N_22267);
nand U22528 (N_22528,N_22113,N_22098);
nor U22529 (N_22529,N_21995,N_22333);
nor U22530 (N_22530,N_21690,N_22000);
and U22531 (N_22531,N_21595,N_21793);
or U22532 (N_22532,N_22151,N_21551);
and U22533 (N_22533,N_21655,N_22414);
nand U22534 (N_22534,N_22309,N_21939);
and U22535 (N_22535,N_21971,N_21332);
or U22536 (N_22536,N_22210,N_22045);
xnor U22537 (N_22537,N_22217,N_21548);
nand U22538 (N_22538,N_22269,N_21834);
and U22539 (N_22539,N_22122,N_21964);
nand U22540 (N_22540,N_22287,N_22256);
or U22541 (N_22541,N_21998,N_22154);
nor U22542 (N_22542,N_22091,N_21304);
nor U22543 (N_22543,N_21253,N_21963);
nor U22544 (N_22544,N_21958,N_21475);
nor U22545 (N_22545,N_21580,N_22039);
nor U22546 (N_22546,N_22207,N_21904);
nand U22547 (N_22547,N_21572,N_22445);
xor U22548 (N_22548,N_21932,N_22378);
or U22549 (N_22549,N_22268,N_22312);
or U22550 (N_22550,N_22239,N_21965);
xnor U22551 (N_22551,N_21709,N_22370);
xor U22552 (N_22552,N_21960,N_21979);
nor U22553 (N_22553,N_21761,N_22024);
xnor U22554 (N_22554,N_21867,N_21916);
or U22555 (N_22555,N_21432,N_22363);
nor U22556 (N_22556,N_21309,N_22022);
nand U22557 (N_22557,N_21807,N_22473);
nand U22558 (N_22558,N_21363,N_22120);
and U22559 (N_22559,N_21492,N_21669);
nand U22560 (N_22560,N_21678,N_22069);
and U22561 (N_22561,N_21798,N_21512);
xnor U22562 (N_22562,N_22092,N_21565);
nand U22563 (N_22563,N_21924,N_21395);
nor U22564 (N_22564,N_21665,N_21562);
nor U22565 (N_22565,N_22483,N_21790);
and U22566 (N_22566,N_22481,N_21968);
xnor U22567 (N_22567,N_22096,N_21388);
and U22568 (N_22568,N_22332,N_21436);
or U22569 (N_22569,N_22127,N_22443);
or U22570 (N_22570,N_21858,N_22432);
nand U22571 (N_22571,N_22172,N_22408);
or U22572 (N_22572,N_22491,N_22146);
nor U22573 (N_22573,N_21883,N_22461);
or U22574 (N_22574,N_21452,N_21508);
nand U22575 (N_22575,N_21897,N_21317);
and U22576 (N_22576,N_21503,N_22319);
nand U22577 (N_22577,N_21973,N_22004);
xnor U22578 (N_22578,N_22040,N_21374);
nand U22579 (N_22579,N_22175,N_22464);
or U22580 (N_22580,N_21270,N_21300);
nand U22581 (N_22581,N_21460,N_21598);
nand U22582 (N_22582,N_21980,N_22047);
or U22583 (N_22583,N_21738,N_21458);
or U22584 (N_22584,N_21334,N_21673);
nor U22585 (N_22585,N_21603,N_21767);
xor U22586 (N_22586,N_22364,N_21461);
nor U22587 (N_22587,N_22074,N_22438);
or U22588 (N_22588,N_21828,N_22019);
and U22589 (N_22589,N_21526,N_21758);
nand U22590 (N_22590,N_21619,N_21365);
and U22591 (N_22591,N_22442,N_22359);
nor U22592 (N_22592,N_21996,N_21536);
nor U22593 (N_22593,N_21990,N_22411);
or U22594 (N_22594,N_22447,N_22140);
nand U22595 (N_22595,N_22030,N_22021);
nor U22596 (N_22596,N_21840,N_21355);
and U22597 (N_22597,N_21560,N_21833);
nor U22598 (N_22598,N_22452,N_21789);
and U22599 (N_22599,N_21473,N_22472);
nand U22600 (N_22600,N_22020,N_22211);
xnor U22601 (N_22601,N_21600,N_22345);
xor U22602 (N_22602,N_22357,N_21283);
or U22603 (N_22603,N_22093,N_21463);
nand U22604 (N_22604,N_21260,N_22228);
nor U22605 (N_22605,N_22141,N_22075);
nand U22606 (N_22606,N_21515,N_21746);
nand U22607 (N_22607,N_22453,N_21301);
nand U22608 (N_22608,N_22388,N_21601);
and U22609 (N_22609,N_21722,N_21715);
nand U22610 (N_22610,N_22107,N_22235);
nand U22611 (N_22611,N_21585,N_22318);
and U22612 (N_22612,N_22051,N_22492);
or U22613 (N_22613,N_21590,N_22067);
and U22614 (N_22614,N_22335,N_21975);
nand U22615 (N_22615,N_21294,N_21918);
xnor U22616 (N_22616,N_21400,N_21267);
and U22617 (N_22617,N_21443,N_21422);
or U22618 (N_22618,N_21437,N_21836);
nand U22619 (N_22619,N_22480,N_22458);
nand U22620 (N_22620,N_21684,N_22402);
nand U22621 (N_22621,N_21768,N_21544);
nand U22622 (N_22622,N_21701,N_21534);
xnor U22623 (N_22623,N_22306,N_21552);
or U22624 (N_22624,N_22204,N_21424);
nor U22625 (N_22625,N_22460,N_21756);
nor U22626 (N_22626,N_22374,N_21373);
or U22627 (N_22627,N_21794,N_21435);
or U22628 (N_22628,N_21806,N_21874);
nor U22629 (N_22629,N_21984,N_22339);
nand U22630 (N_22630,N_21345,N_21926);
and U22631 (N_22631,N_22409,N_21481);
or U22632 (N_22632,N_21307,N_22328);
and U22633 (N_22633,N_21274,N_21569);
nor U22634 (N_22634,N_22253,N_21962);
nor U22635 (N_22635,N_21917,N_21765);
nand U22636 (N_22636,N_22242,N_21561);
nand U22637 (N_22637,N_21788,N_22076);
and U22638 (N_22638,N_21541,N_22278);
nor U22639 (N_22639,N_21531,N_21547);
or U22640 (N_22640,N_21800,N_22490);
xor U22641 (N_22641,N_21375,N_22016);
or U22642 (N_22642,N_22455,N_21927);
xor U22643 (N_22643,N_21431,N_21446);
xor U22644 (N_22644,N_21647,N_21450);
and U22645 (N_22645,N_22214,N_22285);
nor U22646 (N_22646,N_21251,N_22023);
nor U22647 (N_22647,N_21567,N_22187);
xor U22648 (N_22648,N_22106,N_21940);
nand U22649 (N_22649,N_21699,N_22238);
xor U22650 (N_22650,N_21404,N_22246);
or U22651 (N_22651,N_21533,N_21896);
nor U22652 (N_22652,N_22273,N_22459);
and U22653 (N_22653,N_22231,N_22086);
nor U22654 (N_22654,N_21729,N_22186);
nor U22655 (N_22655,N_21258,N_22315);
nor U22656 (N_22656,N_22152,N_21724);
and U22657 (N_22657,N_21381,N_22038);
or U22658 (N_22658,N_21708,N_21869);
or U22659 (N_22659,N_21773,N_21397);
xor U22660 (N_22660,N_21685,N_22351);
or U22661 (N_22661,N_22227,N_21895);
xor U22662 (N_22662,N_21818,N_21406);
or U22663 (N_22663,N_21991,N_21875);
and U22664 (N_22664,N_22484,N_21344);
nor U22665 (N_22665,N_21848,N_21468);
or U22666 (N_22666,N_22262,N_21859);
xnor U22667 (N_22667,N_22065,N_22396);
nand U22668 (N_22668,N_22372,N_21941);
nor U22669 (N_22669,N_21616,N_22277);
xnor U22670 (N_22670,N_22084,N_22463);
or U22671 (N_22671,N_22013,N_21913);
nor U22672 (N_22672,N_21417,N_22355);
nor U22673 (N_22673,N_21324,N_21607);
xnor U22674 (N_22674,N_22422,N_21465);
nor U22675 (N_22675,N_21976,N_22115);
or U22676 (N_22676,N_21440,N_21378);
or U22677 (N_22677,N_21537,N_21866);
and U22678 (N_22678,N_21745,N_22353);
nor U22679 (N_22679,N_22245,N_21719);
or U22680 (N_22680,N_21546,N_21770);
nor U22681 (N_22681,N_22289,N_21442);
or U22682 (N_22682,N_22249,N_22184);
nand U22683 (N_22683,N_22469,N_21657);
xnor U22684 (N_22684,N_22385,N_21954);
nand U22685 (N_22685,N_21827,N_22340);
or U22686 (N_22686,N_22323,N_22382);
or U22687 (N_22687,N_21396,N_21319);
or U22688 (N_22688,N_21499,N_22145);
and U22689 (N_22689,N_22167,N_21441);
and U22690 (N_22690,N_22346,N_21327);
nor U22691 (N_22691,N_21371,N_21650);
and U22692 (N_22692,N_21584,N_22320);
xor U22693 (N_22693,N_21582,N_21920);
nor U22694 (N_22694,N_21372,N_21634);
nor U22695 (N_22695,N_21656,N_21814);
and U22696 (N_22696,N_22054,N_21674);
nand U22697 (N_22697,N_21636,N_21297);
and U22698 (N_22698,N_21529,N_22259);
and U22699 (N_22699,N_22173,N_22178);
nor U22700 (N_22700,N_21826,N_22125);
nor U22701 (N_22701,N_22170,N_21675);
nor U22702 (N_22702,N_21387,N_22104);
xnor U22703 (N_22703,N_21769,N_22121);
nand U22704 (N_22704,N_22250,N_21356);
and U22705 (N_22705,N_22362,N_22423);
and U22706 (N_22706,N_21449,N_22329);
or U22707 (N_22707,N_22478,N_21776);
or U22708 (N_22708,N_22042,N_21384);
or U22709 (N_22709,N_21726,N_21403);
nor U22710 (N_22710,N_22404,N_21772);
xor U22711 (N_22711,N_21322,N_21925);
xor U22712 (N_22712,N_21705,N_21539);
and U22713 (N_22713,N_21929,N_21802);
or U22714 (N_22714,N_22230,N_22037);
or U22715 (N_22715,N_21887,N_22102);
nand U22716 (N_22716,N_21997,N_22226);
or U22717 (N_22717,N_22361,N_21447);
nor U22718 (N_22718,N_21652,N_21741);
nand U22719 (N_22719,N_21841,N_21706);
nor U22720 (N_22720,N_21592,N_21779);
or U22721 (N_22721,N_21872,N_21594);
xnor U22722 (N_22722,N_22094,N_22163);
nor U22723 (N_22723,N_21318,N_21486);
or U22724 (N_22724,N_21306,N_21612);
nand U22725 (N_22725,N_21945,N_22079);
nor U22726 (N_22726,N_22196,N_22428);
nor U22727 (N_22727,N_21370,N_21415);
and U22728 (N_22728,N_22108,N_22430);
nand U22729 (N_22729,N_21907,N_21527);
nor U22730 (N_22730,N_21467,N_21434);
and U22731 (N_22731,N_21495,N_21727);
nand U22732 (N_22732,N_22044,N_22325);
or U22733 (N_22733,N_22405,N_22283);
xor U22734 (N_22734,N_22087,N_22377);
or U22735 (N_22735,N_21464,N_21262);
xnor U22736 (N_22736,N_22454,N_21393);
nor U22737 (N_22737,N_22334,N_22281);
and U22738 (N_22738,N_21981,N_21750);
xnor U22739 (N_22739,N_21734,N_21632);
or U22740 (N_22740,N_21554,N_21518);
and U22741 (N_22741,N_21766,N_21972);
nor U22742 (N_22742,N_22446,N_21586);
xor U22743 (N_22743,N_21884,N_21613);
or U22744 (N_22744,N_22134,N_21553);
and U22745 (N_22745,N_21640,N_22027);
or U22746 (N_22746,N_22387,N_21873);
nor U22747 (N_22747,N_21792,N_22095);
and U22748 (N_22748,N_21302,N_21937);
nand U22749 (N_22749,N_22341,N_22090);
nor U22750 (N_22750,N_22080,N_21289);
xnor U22751 (N_22751,N_22389,N_22159);
xnor U22752 (N_22752,N_21822,N_21256);
or U22753 (N_22753,N_21753,N_21579);
nor U22754 (N_22754,N_21942,N_21643);
xnor U22755 (N_22755,N_22229,N_22448);
nand U22756 (N_22756,N_21797,N_21296);
nor U22757 (N_22757,N_22467,N_21894);
xor U22758 (N_22758,N_22271,N_21608);
nor U22759 (N_22759,N_21936,N_22008);
xor U22760 (N_22760,N_21407,N_21854);
and U22761 (N_22761,N_21666,N_21795);
xor U22762 (N_22762,N_22034,N_21731);
nand U22763 (N_22763,N_21777,N_22489);
nand U22764 (N_22764,N_21341,N_21614);
xnor U22765 (N_22765,N_21287,N_22380);
and U22766 (N_22766,N_21457,N_22336);
nand U22767 (N_22767,N_21733,N_21755);
or U22768 (N_22768,N_21338,N_21316);
nor U22769 (N_22769,N_21293,N_22252);
or U22770 (N_22770,N_21852,N_22433);
nand U22771 (N_22771,N_21497,N_22055);
nand U22772 (N_22772,N_21782,N_22410);
xnor U22773 (N_22773,N_22183,N_22350);
xnor U22774 (N_22774,N_21754,N_22485);
or U22775 (N_22775,N_22118,N_21951);
or U22776 (N_22776,N_21538,N_21956);
or U22777 (N_22777,N_21379,N_21346);
or U22778 (N_22778,N_22138,N_22059);
xor U22779 (N_22779,N_22006,N_21849);
xor U22780 (N_22780,N_21308,N_22270);
xor U22781 (N_22781,N_21559,N_21557);
nand U22782 (N_22782,N_21695,N_22441);
and U22783 (N_22783,N_22191,N_21462);
and U22784 (N_22784,N_21688,N_21618);
nand U22785 (N_22785,N_21399,N_21480);
xnor U22786 (N_22786,N_22232,N_21892);
or U22787 (N_22787,N_21732,N_21933);
xor U22788 (N_22788,N_21484,N_21359);
and U22789 (N_22789,N_22308,N_21908);
and U22790 (N_22790,N_22487,N_21783);
xor U22791 (N_22791,N_21329,N_21350);
and U22792 (N_22792,N_21882,N_22036);
or U22793 (N_22793,N_21983,N_21456);
nand U22794 (N_22794,N_21914,N_21816);
nand U22795 (N_22795,N_21735,N_22028);
or U22796 (N_22796,N_21988,N_21491);
xor U22797 (N_22797,N_22243,N_21389);
or U22798 (N_22798,N_22203,N_21796);
xor U22799 (N_22799,N_21507,N_21587);
nand U22800 (N_22800,N_22457,N_22296);
nand U22801 (N_22801,N_22060,N_21881);
nand U22802 (N_22802,N_21330,N_22190);
and U22803 (N_22803,N_21644,N_21702);
xnor U22804 (N_22804,N_21771,N_21298);
nor U22805 (N_22805,N_21711,N_21739);
and U22806 (N_22806,N_21482,N_21747);
and U22807 (N_22807,N_21433,N_22294);
nor U22808 (N_22808,N_22444,N_22164);
and U22809 (N_22809,N_22407,N_21259);
and U22810 (N_22810,N_21950,N_22168);
nand U22811 (N_22811,N_21857,N_21946);
xnor U22812 (N_22812,N_21288,N_21851);
nand U22813 (N_22813,N_21799,N_21813);
nand U22814 (N_22814,N_22302,N_21472);
nand U22815 (N_22815,N_21455,N_21514);
xnor U22816 (N_22816,N_21845,N_22160);
and U22817 (N_22817,N_22321,N_22495);
xnor U22818 (N_22818,N_21509,N_21850);
and U22819 (N_22819,N_21323,N_22043);
xnor U22820 (N_22820,N_21697,N_21994);
or U22821 (N_22821,N_21519,N_21269);
and U22822 (N_22822,N_22426,N_22344);
and U22823 (N_22823,N_21430,N_22486);
xnor U22824 (N_22824,N_21532,N_22293);
xor U22825 (N_22825,N_21281,N_21376);
and U22826 (N_22826,N_22352,N_22149);
nand U22827 (N_22827,N_22147,N_21689);
and U22828 (N_22828,N_22496,N_21775);
nor U22829 (N_22829,N_21543,N_22169);
nor U22830 (N_22830,N_22068,N_21325);
xnor U22831 (N_22831,N_21668,N_21354);
or U22832 (N_22832,N_22384,N_21646);
and U22833 (N_22833,N_21934,N_22424);
xor U22834 (N_22834,N_21284,N_22071);
nor U22835 (N_22835,N_21380,N_22179);
xnor U22836 (N_22836,N_21413,N_22189);
or U22837 (N_22837,N_22010,N_21863);
or U22838 (N_22838,N_22116,N_21909);
or U22839 (N_22839,N_21808,N_22456);
and U22840 (N_22840,N_21252,N_22011);
nor U22841 (N_22841,N_21438,N_21588);
and U22842 (N_22842,N_22063,N_21681);
xnor U22843 (N_22843,N_22097,N_21728);
xnor U22844 (N_22844,N_21313,N_21409);
nor U22845 (N_22845,N_21266,N_21853);
and U22846 (N_22846,N_21639,N_22081);
and U22847 (N_22847,N_21340,N_21265);
or U22848 (N_22848,N_21279,N_22192);
or U22849 (N_22849,N_22394,N_21752);
or U22850 (N_22850,N_21791,N_22208);
or U22851 (N_22851,N_21989,N_22434);
nor U22852 (N_22852,N_22161,N_21693);
xor U22853 (N_22853,N_21649,N_21428);
and U22854 (N_22854,N_22462,N_21819);
or U22855 (N_22855,N_22265,N_22199);
nand U22856 (N_22856,N_21824,N_22261);
nand U22857 (N_22857,N_22009,N_21844);
and U22858 (N_22858,N_21425,N_21906);
xor U22859 (N_22859,N_21679,N_22347);
nor U22860 (N_22860,N_22126,N_21268);
nor U22861 (N_22861,N_21774,N_21928);
xnor U22862 (N_22862,N_22383,N_21419);
or U22863 (N_22863,N_21861,N_22412);
and U22864 (N_22864,N_21787,N_22139);
and U22865 (N_22865,N_21876,N_22322);
or U22866 (N_22866,N_22114,N_21856);
nor U22867 (N_22867,N_21922,N_22419);
nand U22868 (N_22868,N_21911,N_21847);
and U22869 (N_22869,N_22416,N_22395);
nor U22870 (N_22870,N_22015,N_21716);
and U22871 (N_22871,N_22465,N_21444);
or U22872 (N_22872,N_22052,N_22221);
nor U22873 (N_22873,N_21624,N_21427);
xor U22874 (N_22874,N_22012,N_21622);
xnor U22875 (N_22875,N_22479,N_21687);
nand U22876 (N_22876,N_22266,N_21286);
nand U22877 (N_22877,N_21751,N_21742);
or U22878 (N_22878,N_21961,N_21662);
and U22879 (N_22879,N_21520,N_22450);
and U22880 (N_22880,N_21846,N_21880);
or U22881 (N_22881,N_21292,N_21889);
and U22882 (N_22882,N_22148,N_21943);
xor U22883 (N_22883,N_21670,N_21478);
xnor U22884 (N_22884,N_21832,N_22180);
xnor U22885 (N_22885,N_21574,N_22155);
nor U22886 (N_22886,N_21659,N_21367);
nor U22887 (N_22887,N_22247,N_21571);
xor U22888 (N_22888,N_22066,N_22110);
xnor U22889 (N_22889,N_22048,N_22244);
xor U22890 (N_22890,N_21361,N_21500);
and U22891 (N_22891,N_22397,N_22390);
xor U22892 (N_22892,N_22371,N_21890);
nand U22893 (N_22893,N_21521,N_21336);
nand U22894 (N_22894,N_21597,N_21764);
or U22895 (N_22895,N_22156,N_22421);
or U22896 (N_22896,N_22365,N_22119);
nor U22897 (N_22897,N_22026,N_21978);
and U22898 (N_22898,N_21278,N_22470);
nand U22899 (N_22899,N_22174,N_21410);
and U22900 (N_22900,N_22219,N_21620);
or U22901 (N_22901,N_22153,N_22275);
nand U22902 (N_22902,N_21623,N_21310);
xnor U22903 (N_22903,N_21825,N_21506);
nand U22904 (N_22904,N_21947,N_21470);
or U22905 (N_22905,N_21982,N_22280);
nor U22906 (N_22906,N_21525,N_21352);
nor U22907 (N_22907,N_21581,N_21648);
nor U22908 (N_22908,N_21935,N_21899);
and U22909 (N_22909,N_22279,N_21910);
or U22910 (N_22910,N_21879,N_22135);
and U22911 (N_22911,N_22258,N_21564);
xnor U22912 (N_22912,N_21686,N_21555);
and U22913 (N_22913,N_21255,N_21348);
xnor U22914 (N_22914,N_22194,N_21606);
or U22915 (N_22915,N_22299,N_21312);
and U22916 (N_22916,N_21930,N_21575);
nor U22917 (N_22917,N_21691,N_22349);
xor U22918 (N_22918,N_21676,N_22165);
or U22919 (N_22919,N_21263,N_22050);
nor U22920 (N_22920,N_21609,N_21653);
nand U22921 (N_22921,N_22403,N_22018);
and U22922 (N_22922,N_21280,N_22284);
xor U22923 (N_22923,N_22085,N_22391);
or U22924 (N_22924,N_21762,N_21641);
or U22925 (N_22925,N_22089,N_21839);
nor U22926 (N_22926,N_22077,N_22356);
xnor U22927 (N_22927,N_22197,N_22143);
xor U22928 (N_22928,N_22200,N_22498);
xnor U22929 (N_22929,N_21394,N_21261);
xor U22930 (N_22930,N_22124,N_22062);
nor U22931 (N_22931,N_21589,N_22112);
or U22932 (N_22932,N_22157,N_21439);
and U22933 (N_22933,N_21487,N_21493);
and U22934 (N_22934,N_21577,N_21683);
or U22935 (N_22935,N_22215,N_22058);
nor U22936 (N_22936,N_22420,N_22171);
and U22937 (N_22937,N_21999,N_22436);
nand U22938 (N_22938,N_21627,N_22100);
or U22939 (N_22939,N_22331,N_21923);
or U22940 (N_22940,N_22220,N_21700);
nand U22941 (N_22941,N_22276,N_22413);
nand U22942 (N_22942,N_21540,N_21498);
nand U22943 (N_22943,N_21635,N_21821);
nor U22944 (N_22944,N_21974,N_21418);
or U22945 (N_22945,N_21474,N_21944);
xor U22946 (N_22946,N_22264,N_22327);
and U22947 (N_22947,N_21451,N_21599);
and U22948 (N_22948,N_22418,N_21664);
xor U22949 (N_22949,N_21843,N_22429);
nand U22950 (N_22950,N_22475,N_21391);
and U22951 (N_22951,N_21804,N_22311);
and U22952 (N_22952,N_21785,N_22466);
and U22953 (N_22953,N_22082,N_22307);
and U22954 (N_22954,N_22002,N_21368);
or U22955 (N_22955,N_21494,N_21328);
xor U22956 (N_22956,N_21919,N_21382);
nand U22957 (N_22957,N_21912,N_22476);
nand U22958 (N_22958,N_21902,N_22286);
nor U22959 (N_22959,N_21871,N_22255);
or U22960 (N_22960,N_21426,N_21893);
and U22961 (N_22961,N_21898,N_21390);
nand U22962 (N_22962,N_21596,N_22083);
or U22963 (N_22963,N_21282,N_22406);
or U22964 (N_22964,N_22301,N_21886);
xor U22965 (N_22965,N_22223,N_21273);
and U22966 (N_22966,N_22376,N_21250);
nor U22967 (N_22967,N_21621,N_21496);
nand U22968 (N_22968,N_22292,N_21992);
nand U22969 (N_22969,N_22282,N_22290);
nor U22970 (N_22970,N_22130,N_22078);
xnor U22971 (N_22971,N_21987,N_21831);
nor U22972 (N_22972,N_22003,N_22417);
xnor U22973 (N_22973,N_21703,N_21386);
nand U22974 (N_22974,N_22482,N_21704);
and U22975 (N_22975,N_21736,N_22375);
or U22976 (N_22976,N_21931,N_21862);
or U22977 (N_22977,N_21993,N_21710);
or U22978 (N_22978,N_22474,N_22237);
nor U22979 (N_22979,N_21967,N_21511);
nand U22980 (N_22980,N_21466,N_21421);
or U22981 (N_22981,N_21524,N_21411);
xor U22982 (N_22982,N_21542,N_22367);
or U22983 (N_22983,N_21748,N_21905);
nor U22984 (N_22984,N_22029,N_21629);
xnor U22985 (N_22985,N_22234,N_22305);
nand U22986 (N_22986,N_21744,N_21602);
and U22987 (N_22987,N_21335,N_21885);
or U22988 (N_22988,N_22326,N_22193);
nand U22989 (N_22989,N_22014,N_21275);
or U22990 (N_22990,N_21865,N_21402);
or U22991 (N_22991,N_21642,N_22132);
and U22992 (N_22992,N_22185,N_22123);
or U22993 (N_22993,N_21630,N_21901);
nor U22994 (N_22994,N_22338,N_21985);
xnor U22995 (N_22995,N_21966,N_21290);
nand U22996 (N_22996,N_21957,N_21809);
nand U22997 (N_22997,N_22437,N_21528);
xnor U22998 (N_22998,N_21504,N_22497);
or U22999 (N_22999,N_22348,N_22471);
nand U23000 (N_23000,N_21476,N_21778);
and U23001 (N_23001,N_22468,N_21479);
nand U23002 (N_23002,N_22342,N_21326);
and U23003 (N_23003,N_21725,N_22072);
and U23004 (N_23004,N_22401,N_22225);
or U23005 (N_23005,N_21358,N_21712);
nand U23006 (N_23006,N_22103,N_22392);
nor U23007 (N_23007,N_21786,N_22101);
nand U23008 (N_23008,N_21660,N_21763);
nor U23009 (N_23009,N_21573,N_22360);
xor U23010 (N_23010,N_21392,N_22451);
nor U23011 (N_23011,N_21658,N_22181);
and U23012 (N_23012,N_22260,N_21321);
nand U23013 (N_23013,N_21721,N_22206);
or U23014 (N_23014,N_21868,N_22001);
xnor U23015 (N_23015,N_21671,N_22129);
nand U23016 (N_23016,N_22297,N_22288);
and U23017 (N_23017,N_21254,N_21633);
or U23018 (N_23018,N_21717,N_21377);
nand U23019 (N_23019,N_22324,N_22298);
or U23020 (N_23020,N_21864,N_22176);
or U23021 (N_23021,N_21891,N_22314);
nand U23022 (N_23022,N_22477,N_22070);
or U23023 (N_23023,N_21820,N_22295);
nand U23024 (N_23024,N_21408,N_22053);
nor U23025 (N_23025,N_22368,N_22366);
xor U23026 (N_23026,N_21631,N_21610);
nor U23027 (N_23027,N_21837,N_22213);
nand U23028 (N_23028,N_21677,N_21714);
nor U23029 (N_23029,N_21342,N_22449);
nor U23030 (N_23030,N_21362,N_21617);
xor U23031 (N_23031,N_22205,N_22056);
xor U23032 (N_23032,N_21977,N_21952);
or U23033 (N_23033,N_21815,N_22201);
xor U23034 (N_23034,N_22166,N_22254);
nand U23035 (N_23035,N_22310,N_22088);
xnor U23036 (N_23036,N_21545,N_22032);
nor U23037 (N_23037,N_21568,N_21835);
or U23038 (N_23038,N_21591,N_21888);
nor U23039 (N_23039,N_21921,N_21488);
and U23040 (N_23040,N_21311,N_21360);
nand U23041 (N_23041,N_21578,N_21453);
nand U23042 (N_23042,N_22300,N_21383);
xnor U23043 (N_23043,N_21489,N_21502);
nand U23044 (N_23044,N_22188,N_22398);
or U23045 (N_23045,N_22005,N_21490);
nor U23046 (N_23046,N_21720,N_21445);
or U23047 (N_23047,N_21423,N_22177);
xor U23048 (N_23048,N_21781,N_22182);
or U23049 (N_23049,N_22209,N_21737);
xnor U23050 (N_23050,N_22233,N_21501);
xor U23051 (N_23051,N_22343,N_22488);
or U23052 (N_23052,N_22128,N_21730);
nand U23053 (N_23053,N_21412,N_21257);
and U23054 (N_23054,N_21661,N_21485);
nand U23055 (N_23055,N_21276,N_22198);
nor U23056 (N_23056,N_21672,N_22263);
nor U23057 (N_23057,N_22007,N_21900);
or U23058 (N_23058,N_21366,N_21801);
and U23059 (N_23059,N_21566,N_22241);
or U23060 (N_23060,N_21305,N_21749);
or U23061 (N_23061,N_21645,N_21870);
or U23062 (N_23062,N_21784,N_21654);
nor U23063 (N_23063,N_21694,N_22202);
nand U23064 (N_23064,N_21692,N_22248);
nor U23065 (N_23065,N_21855,N_22195);
and U23066 (N_23066,N_21405,N_21448);
or U23067 (N_23067,N_21385,N_21823);
or U23068 (N_23068,N_21838,N_22064);
nor U23069 (N_23069,N_21549,N_22105);
nor U23070 (N_23070,N_21401,N_22144);
nand U23071 (N_23071,N_21314,N_21743);
nor U23072 (N_23072,N_21563,N_22251);
nor U23073 (N_23073,N_21349,N_21955);
nor U23074 (N_23074,N_22330,N_22499);
xnor U23075 (N_23075,N_21277,N_21556);
xor U23076 (N_23076,N_21757,N_21469);
nand U23077 (N_23077,N_22399,N_22099);
and U23078 (N_23078,N_21740,N_21315);
and U23079 (N_23079,N_21347,N_21759);
and U23080 (N_23080,N_21558,N_21707);
nand U23081 (N_23081,N_21583,N_21878);
xor U23082 (N_23082,N_21803,N_22031);
and U23083 (N_23083,N_21505,N_21682);
xnor U23084 (N_23084,N_22224,N_21357);
nand U23085 (N_23085,N_22073,N_21320);
and U23086 (N_23086,N_21637,N_21626);
xor U23087 (N_23087,N_21663,N_21615);
nor U23088 (N_23088,N_21333,N_21817);
or U23089 (N_23089,N_22313,N_22033);
and U23090 (N_23090,N_22373,N_21680);
nand U23091 (N_23091,N_21516,N_22440);
xnor U23092 (N_23092,N_21471,N_21339);
and U23093 (N_23093,N_22435,N_21811);
and U23094 (N_23094,N_21299,N_22381);
or U23095 (N_23095,N_21696,N_22109);
xor U23096 (N_23096,N_22061,N_22162);
nand U23097 (N_23097,N_22304,N_21698);
or U23098 (N_23098,N_22150,N_21604);
and U23099 (N_23099,N_21264,N_21517);
and U23100 (N_23100,N_21810,N_21723);
nor U23101 (N_23101,N_22046,N_21829);
xnor U23102 (N_23102,N_21343,N_21949);
nand U23103 (N_23103,N_21628,N_22049);
or U23104 (N_23104,N_22158,N_22439);
xor U23105 (N_23105,N_22291,N_22111);
nor U23106 (N_23106,N_22133,N_21303);
or U23107 (N_23107,N_21576,N_21570);
xor U23108 (N_23108,N_22493,N_21285);
xor U23109 (N_23109,N_22272,N_22117);
nor U23110 (N_23110,N_21805,N_22137);
xnor U23111 (N_23111,N_21295,N_21369);
nor U23112 (N_23112,N_22393,N_21291);
xnor U23113 (N_23113,N_22425,N_22236);
nor U23114 (N_23114,N_22131,N_22494);
nand U23115 (N_23115,N_22057,N_22240);
xnor U23116 (N_23116,N_21513,N_21638);
or U23117 (N_23117,N_22337,N_21780);
and U23118 (N_23118,N_22354,N_22386);
nor U23119 (N_23119,N_22379,N_21420);
nand U23120 (N_23120,N_22317,N_21429);
nand U23121 (N_23121,N_21953,N_21760);
and U23122 (N_23122,N_22017,N_22369);
or U23123 (N_23123,N_22415,N_22431);
xor U23124 (N_23124,N_21718,N_21713);
xor U23125 (N_23125,N_22351,N_21372);
nor U23126 (N_23126,N_22103,N_21796);
or U23127 (N_23127,N_21402,N_21630);
nor U23128 (N_23128,N_22110,N_21684);
or U23129 (N_23129,N_21742,N_22293);
or U23130 (N_23130,N_21348,N_21415);
xnor U23131 (N_23131,N_22217,N_21530);
xnor U23132 (N_23132,N_21289,N_21800);
nor U23133 (N_23133,N_21456,N_21988);
nor U23134 (N_23134,N_22123,N_22229);
and U23135 (N_23135,N_21440,N_22345);
or U23136 (N_23136,N_21849,N_21782);
xor U23137 (N_23137,N_21798,N_21861);
and U23138 (N_23138,N_22399,N_21813);
and U23139 (N_23139,N_21906,N_21718);
nor U23140 (N_23140,N_21325,N_21429);
nand U23141 (N_23141,N_21587,N_22388);
xnor U23142 (N_23142,N_22068,N_21947);
nor U23143 (N_23143,N_21448,N_21784);
nor U23144 (N_23144,N_22150,N_22498);
xor U23145 (N_23145,N_22216,N_22118);
nor U23146 (N_23146,N_21671,N_21425);
xor U23147 (N_23147,N_22066,N_22341);
nor U23148 (N_23148,N_22411,N_22064);
nor U23149 (N_23149,N_21800,N_22499);
xor U23150 (N_23150,N_21778,N_21840);
nor U23151 (N_23151,N_21360,N_21971);
and U23152 (N_23152,N_22281,N_21272);
and U23153 (N_23153,N_22437,N_21902);
and U23154 (N_23154,N_21791,N_21586);
xnor U23155 (N_23155,N_22112,N_22208);
and U23156 (N_23156,N_21878,N_21454);
nand U23157 (N_23157,N_22033,N_21357);
or U23158 (N_23158,N_21365,N_21503);
xnor U23159 (N_23159,N_21658,N_21527);
xnor U23160 (N_23160,N_21462,N_22163);
xnor U23161 (N_23161,N_22365,N_21282);
or U23162 (N_23162,N_21552,N_21461);
nor U23163 (N_23163,N_21585,N_21326);
xnor U23164 (N_23164,N_22111,N_21945);
nor U23165 (N_23165,N_21582,N_22411);
or U23166 (N_23166,N_21953,N_21570);
and U23167 (N_23167,N_21620,N_22287);
nand U23168 (N_23168,N_21645,N_21934);
nand U23169 (N_23169,N_21810,N_21741);
nor U23170 (N_23170,N_21437,N_21560);
xnor U23171 (N_23171,N_21851,N_22161);
nor U23172 (N_23172,N_22068,N_22213);
and U23173 (N_23173,N_21849,N_21540);
nor U23174 (N_23174,N_21554,N_21704);
nand U23175 (N_23175,N_21666,N_21264);
nor U23176 (N_23176,N_21549,N_22124);
or U23177 (N_23177,N_22154,N_22471);
nor U23178 (N_23178,N_22313,N_22244);
xnor U23179 (N_23179,N_21459,N_22405);
nand U23180 (N_23180,N_21806,N_21461);
nor U23181 (N_23181,N_21417,N_21563);
nor U23182 (N_23182,N_22454,N_22037);
nand U23183 (N_23183,N_21575,N_21683);
or U23184 (N_23184,N_22236,N_22304);
and U23185 (N_23185,N_21759,N_21886);
and U23186 (N_23186,N_21880,N_21356);
or U23187 (N_23187,N_21748,N_21916);
nor U23188 (N_23188,N_21786,N_22001);
xor U23189 (N_23189,N_22184,N_21903);
or U23190 (N_23190,N_21336,N_21803);
and U23191 (N_23191,N_21252,N_21760);
xor U23192 (N_23192,N_21828,N_22313);
nand U23193 (N_23193,N_22189,N_21873);
nand U23194 (N_23194,N_21425,N_22361);
xor U23195 (N_23195,N_22157,N_21773);
xnor U23196 (N_23196,N_22079,N_22324);
xnor U23197 (N_23197,N_21657,N_22486);
nand U23198 (N_23198,N_21685,N_21578);
and U23199 (N_23199,N_22441,N_22251);
or U23200 (N_23200,N_22409,N_21332);
and U23201 (N_23201,N_22006,N_22352);
or U23202 (N_23202,N_22475,N_21993);
or U23203 (N_23203,N_22399,N_21892);
or U23204 (N_23204,N_21924,N_21620);
or U23205 (N_23205,N_22150,N_22111);
xnor U23206 (N_23206,N_21666,N_22070);
nand U23207 (N_23207,N_22102,N_22275);
and U23208 (N_23208,N_21948,N_22243);
nor U23209 (N_23209,N_21949,N_21784);
and U23210 (N_23210,N_22441,N_21254);
or U23211 (N_23211,N_21941,N_21825);
nand U23212 (N_23212,N_21349,N_21811);
or U23213 (N_23213,N_21915,N_21530);
xor U23214 (N_23214,N_22337,N_21428);
nor U23215 (N_23215,N_22315,N_22404);
nor U23216 (N_23216,N_21343,N_22168);
and U23217 (N_23217,N_21709,N_21635);
xnor U23218 (N_23218,N_22138,N_22442);
and U23219 (N_23219,N_22434,N_21592);
or U23220 (N_23220,N_22437,N_22361);
xor U23221 (N_23221,N_21355,N_21383);
and U23222 (N_23222,N_22347,N_22318);
nor U23223 (N_23223,N_22294,N_21743);
nand U23224 (N_23224,N_21925,N_22286);
nor U23225 (N_23225,N_22367,N_21684);
xnor U23226 (N_23226,N_21947,N_22207);
nand U23227 (N_23227,N_21970,N_21726);
xor U23228 (N_23228,N_21633,N_21877);
and U23229 (N_23229,N_22399,N_22353);
nor U23230 (N_23230,N_21316,N_22119);
nor U23231 (N_23231,N_21617,N_21977);
nor U23232 (N_23232,N_21953,N_21331);
and U23233 (N_23233,N_21598,N_21317);
nand U23234 (N_23234,N_21757,N_21354);
and U23235 (N_23235,N_22043,N_21704);
nand U23236 (N_23236,N_21622,N_21288);
nor U23237 (N_23237,N_21824,N_21886);
nor U23238 (N_23238,N_21852,N_21585);
xnor U23239 (N_23239,N_22138,N_21326);
and U23240 (N_23240,N_22166,N_21879);
and U23241 (N_23241,N_21529,N_22421);
nor U23242 (N_23242,N_22333,N_22492);
xnor U23243 (N_23243,N_22173,N_21741);
xnor U23244 (N_23244,N_22205,N_21747);
xnor U23245 (N_23245,N_21478,N_22091);
nor U23246 (N_23246,N_22097,N_22455);
nor U23247 (N_23247,N_21279,N_21526);
nand U23248 (N_23248,N_22438,N_21445);
nor U23249 (N_23249,N_22195,N_22087);
xor U23250 (N_23250,N_22133,N_21897);
and U23251 (N_23251,N_22116,N_21960);
or U23252 (N_23252,N_21460,N_21916);
or U23253 (N_23253,N_21490,N_21365);
and U23254 (N_23254,N_22399,N_21726);
and U23255 (N_23255,N_22430,N_21874);
or U23256 (N_23256,N_22030,N_21728);
or U23257 (N_23257,N_21899,N_21289);
and U23258 (N_23258,N_22427,N_21763);
or U23259 (N_23259,N_21926,N_22014);
nand U23260 (N_23260,N_21945,N_21295);
nand U23261 (N_23261,N_22265,N_21906);
and U23262 (N_23262,N_21292,N_21708);
or U23263 (N_23263,N_21436,N_21843);
or U23264 (N_23264,N_21547,N_22166);
nand U23265 (N_23265,N_21771,N_22377);
nor U23266 (N_23266,N_21489,N_22202);
and U23267 (N_23267,N_22106,N_22103);
and U23268 (N_23268,N_22337,N_22174);
and U23269 (N_23269,N_21520,N_22456);
and U23270 (N_23270,N_22295,N_21643);
nor U23271 (N_23271,N_22401,N_21926);
and U23272 (N_23272,N_21686,N_21457);
xor U23273 (N_23273,N_21421,N_21304);
xor U23274 (N_23274,N_22098,N_22316);
or U23275 (N_23275,N_21861,N_21871);
nand U23276 (N_23276,N_21338,N_21515);
nor U23277 (N_23277,N_22166,N_21896);
or U23278 (N_23278,N_22098,N_21776);
or U23279 (N_23279,N_21284,N_22053);
xor U23280 (N_23280,N_22313,N_21339);
nor U23281 (N_23281,N_22451,N_21417);
and U23282 (N_23282,N_21944,N_22035);
or U23283 (N_23283,N_22166,N_21796);
nand U23284 (N_23284,N_21361,N_21356);
nor U23285 (N_23285,N_21864,N_21665);
nor U23286 (N_23286,N_21583,N_21600);
and U23287 (N_23287,N_21883,N_21252);
nand U23288 (N_23288,N_21828,N_21914);
xor U23289 (N_23289,N_22478,N_22304);
or U23290 (N_23290,N_21709,N_21675);
xnor U23291 (N_23291,N_21365,N_21275);
or U23292 (N_23292,N_21284,N_22322);
or U23293 (N_23293,N_21656,N_22026);
xnor U23294 (N_23294,N_21425,N_21293);
and U23295 (N_23295,N_21862,N_21591);
xor U23296 (N_23296,N_22038,N_21457);
or U23297 (N_23297,N_22448,N_21777);
nand U23298 (N_23298,N_22041,N_21858);
and U23299 (N_23299,N_21805,N_21992);
nand U23300 (N_23300,N_22312,N_21666);
xor U23301 (N_23301,N_21737,N_22031);
nor U23302 (N_23302,N_22301,N_22197);
nor U23303 (N_23303,N_22155,N_21837);
nand U23304 (N_23304,N_22404,N_21933);
xor U23305 (N_23305,N_21736,N_22426);
nor U23306 (N_23306,N_22381,N_21785);
or U23307 (N_23307,N_22471,N_21799);
nand U23308 (N_23308,N_21430,N_22365);
nand U23309 (N_23309,N_21932,N_21740);
or U23310 (N_23310,N_22065,N_22315);
nand U23311 (N_23311,N_22043,N_21890);
xor U23312 (N_23312,N_22288,N_21773);
nor U23313 (N_23313,N_22449,N_22259);
nor U23314 (N_23314,N_21295,N_21378);
and U23315 (N_23315,N_22271,N_21583);
xnor U23316 (N_23316,N_21848,N_21743);
xor U23317 (N_23317,N_22495,N_22398);
or U23318 (N_23318,N_21763,N_22256);
and U23319 (N_23319,N_22333,N_21886);
nand U23320 (N_23320,N_22416,N_21771);
nand U23321 (N_23321,N_21549,N_21591);
nor U23322 (N_23322,N_22354,N_22099);
and U23323 (N_23323,N_21702,N_22472);
or U23324 (N_23324,N_22463,N_21437);
and U23325 (N_23325,N_21834,N_21267);
nand U23326 (N_23326,N_22433,N_21737);
and U23327 (N_23327,N_21437,N_21698);
nand U23328 (N_23328,N_21846,N_21529);
nor U23329 (N_23329,N_21295,N_21269);
and U23330 (N_23330,N_22438,N_22072);
nand U23331 (N_23331,N_21290,N_21957);
nor U23332 (N_23332,N_21593,N_22408);
xnor U23333 (N_23333,N_21739,N_21494);
and U23334 (N_23334,N_21536,N_21580);
nor U23335 (N_23335,N_21578,N_22043);
and U23336 (N_23336,N_22168,N_22100);
and U23337 (N_23337,N_21866,N_21742);
or U23338 (N_23338,N_21273,N_22052);
or U23339 (N_23339,N_21343,N_22267);
and U23340 (N_23340,N_21712,N_21536);
nor U23341 (N_23341,N_22151,N_22142);
xor U23342 (N_23342,N_22026,N_22356);
xor U23343 (N_23343,N_22346,N_21544);
and U23344 (N_23344,N_21476,N_22033);
nor U23345 (N_23345,N_22069,N_22422);
and U23346 (N_23346,N_22114,N_22278);
nor U23347 (N_23347,N_21736,N_22324);
nor U23348 (N_23348,N_22033,N_22431);
or U23349 (N_23349,N_22293,N_21334);
xnor U23350 (N_23350,N_21983,N_22031);
xor U23351 (N_23351,N_21251,N_22303);
nand U23352 (N_23352,N_22353,N_21252);
nor U23353 (N_23353,N_21822,N_22315);
and U23354 (N_23354,N_21293,N_21433);
or U23355 (N_23355,N_21740,N_21821);
xnor U23356 (N_23356,N_21364,N_21500);
nor U23357 (N_23357,N_21622,N_21818);
nand U23358 (N_23358,N_21504,N_21567);
nor U23359 (N_23359,N_22083,N_21310);
or U23360 (N_23360,N_21542,N_22180);
or U23361 (N_23361,N_21548,N_21479);
or U23362 (N_23362,N_21620,N_22275);
nor U23363 (N_23363,N_21806,N_21274);
nand U23364 (N_23364,N_21652,N_22419);
nor U23365 (N_23365,N_21948,N_21799);
nand U23366 (N_23366,N_21420,N_21462);
nor U23367 (N_23367,N_21710,N_22088);
xor U23368 (N_23368,N_21371,N_22135);
or U23369 (N_23369,N_21989,N_22288);
nor U23370 (N_23370,N_22355,N_22435);
and U23371 (N_23371,N_22373,N_21509);
and U23372 (N_23372,N_21363,N_22078);
and U23373 (N_23373,N_22094,N_22348);
and U23374 (N_23374,N_21912,N_21435);
and U23375 (N_23375,N_22330,N_22398);
nor U23376 (N_23376,N_22103,N_22424);
nor U23377 (N_23377,N_22054,N_21948);
and U23378 (N_23378,N_21995,N_21666);
nor U23379 (N_23379,N_21298,N_21902);
nand U23380 (N_23380,N_22480,N_21657);
or U23381 (N_23381,N_21688,N_21403);
or U23382 (N_23382,N_21477,N_21308);
nand U23383 (N_23383,N_22280,N_22492);
nor U23384 (N_23384,N_21455,N_22207);
xor U23385 (N_23385,N_22200,N_22116);
nand U23386 (N_23386,N_21943,N_22372);
xor U23387 (N_23387,N_21654,N_21633);
xor U23388 (N_23388,N_21431,N_22279);
xor U23389 (N_23389,N_21281,N_22348);
nor U23390 (N_23390,N_22047,N_21844);
or U23391 (N_23391,N_21549,N_21522);
nor U23392 (N_23392,N_21556,N_21655);
nand U23393 (N_23393,N_22367,N_22141);
nand U23394 (N_23394,N_22277,N_21354);
xor U23395 (N_23395,N_21928,N_22140);
nand U23396 (N_23396,N_22320,N_22335);
xor U23397 (N_23397,N_21699,N_22177);
and U23398 (N_23398,N_21477,N_21726);
nor U23399 (N_23399,N_21307,N_22073);
nand U23400 (N_23400,N_21997,N_22336);
xor U23401 (N_23401,N_21955,N_21946);
and U23402 (N_23402,N_21754,N_21485);
nor U23403 (N_23403,N_22105,N_21325);
or U23404 (N_23404,N_21285,N_21287);
nand U23405 (N_23405,N_21800,N_22368);
xnor U23406 (N_23406,N_21446,N_22100);
xnor U23407 (N_23407,N_21977,N_22359);
and U23408 (N_23408,N_21412,N_21342);
or U23409 (N_23409,N_22234,N_21454);
and U23410 (N_23410,N_21310,N_21351);
nor U23411 (N_23411,N_22069,N_21941);
nand U23412 (N_23412,N_21992,N_21929);
xor U23413 (N_23413,N_22299,N_21735);
and U23414 (N_23414,N_21784,N_21800);
nand U23415 (N_23415,N_21864,N_21800);
nand U23416 (N_23416,N_22269,N_21259);
nor U23417 (N_23417,N_22432,N_22060);
xnor U23418 (N_23418,N_21350,N_21940);
nand U23419 (N_23419,N_21367,N_22078);
or U23420 (N_23420,N_21284,N_22365);
or U23421 (N_23421,N_21921,N_21770);
nor U23422 (N_23422,N_22071,N_21614);
nor U23423 (N_23423,N_21433,N_22180);
nand U23424 (N_23424,N_21730,N_21661);
or U23425 (N_23425,N_21921,N_22020);
or U23426 (N_23426,N_22002,N_21646);
or U23427 (N_23427,N_21438,N_21578);
or U23428 (N_23428,N_21601,N_22264);
xnor U23429 (N_23429,N_21569,N_21944);
xnor U23430 (N_23430,N_22357,N_22202);
xor U23431 (N_23431,N_21337,N_21390);
nor U23432 (N_23432,N_22217,N_21972);
nor U23433 (N_23433,N_21562,N_21612);
nand U23434 (N_23434,N_21618,N_21561);
nand U23435 (N_23435,N_22248,N_22227);
nor U23436 (N_23436,N_22433,N_22343);
or U23437 (N_23437,N_21966,N_21505);
xor U23438 (N_23438,N_21868,N_21719);
nor U23439 (N_23439,N_22344,N_22379);
nand U23440 (N_23440,N_21696,N_21555);
xnor U23441 (N_23441,N_21755,N_22480);
nand U23442 (N_23442,N_22348,N_21395);
or U23443 (N_23443,N_21359,N_22093);
nand U23444 (N_23444,N_21435,N_22080);
and U23445 (N_23445,N_22422,N_22008);
and U23446 (N_23446,N_21406,N_22499);
or U23447 (N_23447,N_22023,N_22198);
and U23448 (N_23448,N_21596,N_22437);
nand U23449 (N_23449,N_22082,N_22220);
nor U23450 (N_23450,N_21853,N_21882);
and U23451 (N_23451,N_22082,N_22173);
or U23452 (N_23452,N_21551,N_22356);
nand U23453 (N_23453,N_22437,N_21279);
nand U23454 (N_23454,N_21971,N_22421);
xor U23455 (N_23455,N_21276,N_22446);
xor U23456 (N_23456,N_22283,N_21950);
nand U23457 (N_23457,N_21741,N_21756);
and U23458 (N_23458,N_22490,N_22324);
nor U23459 (N_23459,N_21668,N_21941);
and U23460 (N_23460,N_22410,N_22045);
xor U23461 (N_23461,N_22498,N_22134);
nand U23462 (N_23462,N_22492,N_21584);
xnor U23463 (N_23463,N_21433,N_21863);
or U23464 (N_23464,N_21326,N_21969);
nor U23465 (N_23465,N_21437,N_21435);
or U23466 (N_23466,N_21606,N_21324);
nand U23467 (N_23467,N_21562,N_22433);
nand U23468 (N_23468,N_21872,N_22199);
xnor U23469 (N_23469,N_21419,N_21751);
or U23470 (N_23470,N_21321,N_22451);
nand U23471 (N_23471,N_22425,N_22034);
xor U23472 (N_23472,N_22410,N_21373);
nand U23473 (N_23473,N_22394,N_21993);
or U23474 (N_23474,N_22454,N_21573);
or U23475 (N_23475,N_21718,N_21858);
nand U23476 (N_23476,N_21763,N_21712);
nand U23477 (N_23477,N_21664,N_22443);
xor U23478 (N_23478,N_22417,N_22411);
and U23479 (N_23479,N_21897,N_21261);
nor U23480 (N_23480,N_21531,N_21974);
nor U23481 (N_23481,N_22367,N_21714);
xor U23482 (N_23482,N_21980,N_22172);
nand U23483 (N_23483,N_22051,N_21941);
nand U23484 (N_23484,N_22408,N_21509);
nor U23485 (N_23485,N_22262,N_22081);
nand U23486 (N_23486,N_21457,N_22486);
nand U23487 (N_23487,N_21703,N_21463);
and U23488 (N_23488,N_22304,N_22297);
xnor U23489 (N_23489,N_22303,N_22486);
or U23490 (N_23490,N_21941,N_21770);
or U23491 (N_23491,N_21350,N_22463);
nor U23492 (N_23492,N_21581,N_21304);
xnor U23493 (N_23493,N_22243,N_22280);
and U23494 (N_23494,N_21303,N_22111);
or U23495 (N_23495,N_21973,N_21707);
nand U23496 (N_23496,N_22330,N_22362);
and U23497 (N_23497,N_21443,N_21377);
nand U23498 (N_23498,N_21915,N_22104);
or U23499 (N_23499,N_21323,N_21377);
nand U23500 (N_23500,N_21928,N_22315);
xnor U23501 (N_23501,N_21316,N_21866);
or U23502 (N_23502,N_22226,N_22201);
nand U23503 (N_23503,N_21400,N_21350);
xor U23504 (N_23504,N_21393,N_21708);
nor U23505 (N_23505,N_21858,N_22218);
nor U23506 (N_23506,N_21423,N_21755);
xor U23507 (N_23507,N_22288,N_21767);
and U23508 (N_23508,N_22260,N_21555);
nand U23509 (N_23509,N_22377,N_21779);
or U23510 (N_23510,N_22186,N_21937);
or U23511 (N_23511,N_21699,N_22092);
nor U23512 (N_23512,N_22170,N_21673);
xnor U23513 (N_23513,N_21485,N_22294);
or U23514 (N_23514,N_21571,N_21986);
and U23515 (N_23515,N_21602,N_22191);
xnor U23516 (N_23516,N_21991,N_22206);
or U23517 (N_23517,N_22428,N_22431);
and U23518 (N_23518,N_21285,N_21605);
and U23519 (N_23519,N_21415,N_21501);
nand U23520 (N_23520,N_22136,N_21330);
nor U23521 (N_23521,N_21925,N_21863);
nor U23522 (N_23522,N_22416,N_22192);
xnor U23523 (N_23523,N_21559,N_21988);
nor U23524 (N_23524,N_21815,N_21513);
nor U23525 (N_23525,N_22249,N_21853);
nor U23526 (N_23526,N_22429,N_21756);
nand U23527 (N_23527,N_21936,N_21505);
or U23528 (N_23528,N_21674,N_21673);
xor U23529 (N_23529,N_21985,N_22100);
and U23530 (N_23530,N_22120,N_21980);
nor U23531 (N_23531,N_22165,N_21823);
xnor U23532 (N_23532,N_22137,N_21437);
nor U23533 (N_23533,N_21405,N_21717);
xnor U23534 (N_23534,N_21320,N_22249);
or U23535 (N_23535,N_22485,N_22061);
nand U23536 (N_23536,N_21704,N_22402);
or U23537 (N_23537,N_21806,N_21552);
nor U23538 (N_23538,N_21621,N_22378);
or U23539 (N_23539,N_22015,N_22191);
and U23540 (N_23540,N_21803,N_22409);
and U23541 (N_23541,N_21714,N_22282);
nand U23542 (N_23542,N_22251,N_21310);
nand U23543 (N_23543,N_21491,N_22310);
or U23544 (N_23544,N_22005,N_22041);
nor U23545 (N_23545,N_22401,N_21652);
nand U23546 (N_23546,N_21595,N_21664);
and U23547 (N_23547,N_21562,N_22370);
nor U23548 (N_23548,N_22277,N_22107);
nand U23549 (N_23549,N_22383,N_21935);
and U23550 (N_23550,N_21924,N_21810);
xor U23551 (N_23551,N_21620,N_21827);
and U23552 (N_23552,N_21497,N_21580);
xor U23553 (N_23553,N_21460,N_21796);
and U23554 (N_23554,N_22207,N_21964);
and U23555 (N_23555,N_21387,N_21301);
xor U23556 (N_23556,N_21387,N_21557);
nand U23557 (N_23557,N_22230,N_22291);
nand U23558 (N_23558,N_21920,N_22362);
or U23559 (N_23559,N_22064,N_21432);
nand U23560 (N_23560,N_21572,N_22304);
xnor U23561 (N_23561,N_22046,N_22086);
or U23562 (N_23562,N_21549,N_21752);
nand U23563 (N_23563,N_21428,N_21902);
or U23564 (N_23564,N_22192,N_21342);
nor U23565 (N_23565,N_21326,N_22116);
and U23566 (N_23566,N_21478,N_22186);
and U23567 (N_23567,N_22293,N_22043);
and U23568 (N_23568,N_21343,N_22070);
xor U23569 (N_23569,N_22093,N_21369);
nand U23570 (N_23570,N_21785,N_22483);
or U23571 (N_23571,N_22268,N_21463);
or U23572 (N_23572,N_22428,N_21429);
xnor U23573 (N_23573,N_21274,N_22481);
nor U23574 (N_23574,N_21696,N_22157);
or U23575 (N_23575,N_22488,N_21884);
nor U23576 (N_23576,N_21559,N_22390);
xnor U23577 (N_23577,N_21437,N_22321);
or U23578 (N_23578,N_22197,N_22138);
nand U23579 (N_23579,N_21288,N_22347);
or U23580 (N_23580,N_21440,N_21289);
nand U23581 (N_23581,N_21451,N_21780);
nor U23582 (N_23582,N_21279,N_21292);
and U23583 (N_23583,N_22220,N_21859);
nand U23584 (N_23584,N_22434,N_21845);
xnor U23585 (N_23585,N_22108,N_21531);
xnor U23586 (N_23586,N_21436,N_21469);
or U23587 (N_23587,N_21271,N_21416);
nor U23588 (N_23588,N_21979,N_21386);
and U23589 (N_23589,N_21266,N_22481);
xor U23590 (N_23590,N_22083,N_22367);
nand U23591 (N_23591,N_22345,N_22250);
xor U23592 (N_23592,N_21274,N_21439);
or U23593 (N_23593,N_21763,N_21553);
xor U23594 (N_23594,N_21279,N_21264);
nand U23595 (N_23595,N_22243,N_22069);
or U23596 (N_23596,N_21595,N_21974);
and U23597 (N_23597,N_21510,N_21741);
nand U23598 (N_23598,N_21608,N_21947);
xor U23599 (N_23599,N_22456,N_21859);
xnor U23600 (N_23600,N_21988,N_22227);
or U23601 (N_23601,N_21380,N_21640);
nor U23602 (N_23602,N_22219,N_22343);
or U23603 (N_23603,N_22470,N_22364);
nand U23604 (N_23604,N_21909,N_21957);
or U23605 (N_23605,N_21613,N_21869);
and U23606 (N_23606,N_21934,N_22470);
and U23607 (N_23607,N_21940,N_21404);
nor U23608 (N_23608,N_21303,N_21675);
or U23609 (N_23609,N_22453,N_21766);
nand U23610 (N_23610,N_21365,N_22230);
nor U23611 (N_23611,N_21510,N_22058);
nand U23612 (N_23612,N_21557,N_22313);
nor U23613 (N_23613,N_22291,N_21261);
and U23614 (N_23614,N_21691,N_22214);
or U23615 (N_23615,N_21360,N_22236);
nor U23616 (N_23616,N_22014,N_21681);
xnor U23617 (N_23617,N_22184,N_21918);
or U23618 (N_23618,N_22093,N_22117);
xor U23619 (N_23619,N_22348,N_22217);
and U23620 (N_23620,N_21676,N_21589);
and U23621 (N_23621,N_21597,N_21410);
xor U23622 (N_23622,N_21614,N_21710);
nand U23623 (N_23623,N_21559,N_21328);
xnor U23624 (N_23624,N_21320,N_22183);
nand U23625 (N_23625,N_22063,N_22195);
xnor U23626 (N_23626,N_21899,N_22447);
or U23627 (N_23627,N_22194,N_21590);
or U23628 (N_23628,N_22448,N_21356);
nand U23629 (N_23629,N_22217,N_21957);
xor U23630 (N_23630,N_21440,N_22465);
nor U23631 (N_23631,N_21827,N_22121);
or U23632 (N_23632,N_22341,N_21977);
or U23633 (N_23633,N_22173,N_22294);
and U23634 (N_23634,N_21842,N_21589);
xor U23635 (N_23635,N_21562,N_21423);
nor U23636 (N_23636,N_21646,N_21267);
and U23637 (N_23637,N_22153,N_21707);
xnor U23638 (N_23638,N_21423,N_22321);
xnor U23639 (N_23639,N_22327,N_21524);
xnor U23640 (N_23640,N_22015,N_22121);
or U23641 (N_23641,N_21965,N_22177);
or U23642 (N_23642,N_21960,N_21741);
or U23643 (N_23643,N_22037,N_22099);
nand U23644 (N_23644,N_21313,N_21549);
or U23645 (N_23645,N_21904,N_21918);
nor U23646 (N_23646,N_21418,N_22006);
xor U23647 (N_23647,N_21551,N_22458);
nand U23648 (N_23648,N_22186,N_21607);
nor U23649 (N_23649,N_21359,N_21370);
nor U23650 (N_23650,N_21866,N_21568);
and U23651 (N_23651,N_22423,N_22377);
xnor U23652 (N_23652,N_22410,N_21481);
and U23653 (N_23653,N_21687,N_21346);
or U23654 (N_23654,N_21419,N_21693);
nor U23655 (N_23655,N_21531,N_22458);
nand U23656 (N_23656,N_21981,N_22414);
nand U23657 (N_23657,N_22247,N_21468);
and U23658 (N_23658,N_21250,N_22079);
and U23659 (N_23659,N_21990,N_21661);
nor U23660 (N_23660,N_22071,N_21523);
xor U23661 (N_23661,N_21795,N_21955);
nand U23662 (N_23662,N_21937,N_21631);
nand U23663 (N_23663,N_21950,N_21901);
nor U23664 (N_23664,N_22472,N_21681);
nor U23665 (N_23665,N_21259,N_21286);
nand U23666 (N_23666,N_22080,N_21903);
nand U23667 (N_23667,N_21569,N_21873);
and U23668 (N_23668,N_21551,N_21608);
nand U23669 (N_23669,N_21438,N_21322);
nand U23670 (N_23670,N_22435,N_21614);
nor U23671 (N_23671,N_22484,N_22144);
or U23672 (N_23672,N_22283,N_21399);
nor U23673 (N_23673,N_22380,N_21979);
xor U23674 (N_23674,N_21402,N_22356);
nand U23675 (N_23675,N_22186,N_21789);
xnor U23676 (N_23676,N_21685,N_21857);
nand U23677 (N_23677,N_21821,N_22439);
and U23678 (N_23678,N_21828,N_21709);
or U23679 (N_23679,N_21682,N_22486);
or U23680 (N_23680,N_21866,N_21890);
nor U23681 (N_23681,N_22397,N_21583);
nand U23682 (N_23682,N_22193,N_21817);
nand U23683 (N_23683,N_22106,N_22027);
xnor U23684 (N_23684,N_22456,N_21935);
xor U23685 (N_23685,N_22392,N_21484);
nand U23686 (N_23686,N_21932,N_21738);
or U23687 (N_23687,N_21785,N_21952);
or U23688 (N_23688,N_22470,N_21447);
nand U23689 (N_23689,N_21858,N_21881);
nand U23690 (N_23690,N_21487,N_21253);
or U23691 (N_23691,N_22101,N_21972);
xor U23692 (N_23692,N_21417,N_21755);
nand U23693 (N_23693,N_22396,N_22304);
or U23694 (N_23694,N_21427,N_22379);
xor U23695 (N_23695,N_21590,N_21481);
nor U23696 (N_23696,N_21814,N_21611);
xor U23697 (N_23697,N_22104,N_21872);
nand U23698 (N_23698,N_22395,N_21296);
nand U23699 (N_23699,N_22332,N_21423);
nor U23700 (N_23700,N_21967,N_21690);
or U23701 (N_23701,N_22017,N_22085);
and U23702 (N_23702,N_22113,N_21563);
nand U23703 (N_23703,N_22072,N_21621);
or U23704 (N_23704,N_22295,N_22082);
nand U23705 (N_23705,N_22108,N_21802);
nand U23706 (N_23706,N_22262,N_21593);
or U23707 (N_23707,N_22062,N_21541);
nand U23708 (N_23708,N_21886,N_21987);
or U23709 (N_23709,N_22264,N_21419);
nor U23710 (N_23710,N_21328,N_21428);
xnor U23711 (N_23711,N_21562,N_22480);
nand U23712 (N_23712,N_21526,N_21606);
nand U23713 (N_23713,N_21420,N_21359);
xor U23714 (N_23714,N_22209,N_21282);
or U23715 (N_23715,N_22112,N_21427);
xnor U23716 (N_23716,N_21504,N_21510);
nand U23717 (N_23717,N_22487,N_21684);
nand U23718 (N_23718,N_21349,N_21619);
xor U23719 (N_23719,N_22053,N_21378);
or U23720 (N_23720,N_22035,N_21492);
or U23721 (N_23721,N_21384,N_21670);
nand U23722 (N_23722,N_22473,N_22023);
and U23723 (N_23723,N_21267,N_22074);
nand U23724 (N_23724,N_21259,N_22000);
or U23725 (N_23725,N_21385,N_21273);
nand U23726 (N_23726,N_21344,N_22130);
or U23727 (N_23727,N_22179,N_22447);
xor U23728 (N_23728,N_21983,N_22026);
or U23729 (N_23729,N_21793,N_21904);
nand U23730 (N_23730,N_21813,N_21866);
nand U23731 (N_23731,N_22163,N_21538);
nand U23732 (N_23732,N_22429,N_21419);
or U23733 (N_23733,N_21732,N_21548);
or U23734 (N_23734,N_21260,N_22403);
nand U23735 (N_23735,N_22201,N_22325);
and U23736 (N_23736,N_21308,N_21347);
nor U23737 (N_23737,N_21754,N_22293);
or U23738 (N_23738,N_21586,N_21425);
or U23739 (N_23739,N_21448,N_21666);
xnor U23740 (N_23740,N_21928,N_21736);
nand U23741 (N_23741,N_21957,N_21321);
nor U23742 (N_23742,N_22087,N_21739);
and U23743 (N_23743,N_21673,N_22293);
or U23744 (N_23744,N_21850,N_22424);
xor U23745 (N_23745,N_22020,N_22023);
nand U23746 (N_23746,N_21904,N_21272);
nand U23747 (N_23747,N_21768,N_21703);
xor U23748 (N_23748,N_21980,N_21852);
or U23749 (N_23749,N_22049,N_22091);
nand U23750 (N_23750,N_23109,N_23261);
and U23751 (N_23751,N_22782,N_23742);
nor U23752 (N_23752,N_23516,N_22941);
nand U23753 (N_23753,N_22584,N_22596);
nand U23754 (N_23754,N_22899,N_22965);
or U23755 (N_23755,N_23463,N_22910);
xor U23756 (N_23756,N_22845,N_22936);
nor U23757 (N_23757,N_22576,N_22582);
or U23758 (N_23758,N_22716,N_23552);
nor U23759 (N_23759,N_23720,N_22517);
nand U23760 (N_23760,N_22858,N_23195);
nor U23761 (N_23761,N_23290,N_23601);
or U23762 (N_23762,N_23030,N_23500);
nor U23763 (N_23763,N_23490,N_23431);
xor U23764 (N_23764,N_23162,N_23170);
nor U23765 (N_23765,N_22696,N_22616);
nand U23766 (N_23766,N_22760,N_23201);
or U23767 (N_23767,N_23114,N_22879);
nand U23768 (N_23768,N_23364,N_22556);
and U23769 (N_23769,N_23453,N_23724);
nor U23770 (N_23770,N_23040,N_22698);
or U23771 (N_23771,N_22786,N_22962);
and U23772 (N_23772,N_23477,N_22836);
nor U23773 (N_23773,N_23726,N_22945);
nand U23774 (N_23774,N_22662,N_23407);
xnor U23775 (N_23775,N_22923,N_23338);
nand U23776 (N_23776,N_22809,N_22885);
xor U23777 (N_23777,N_22881,N_22621);
xor U23778 (N_23778,N_23438,N_22915);
or U23779 (N_23779,N_23586,N_22762);
or U23780 (N_23780,N_22612,N_23445);
nand U23781 (N_23781,N_22999,N_22839);
and U23782 (N_23782,N_23672,N_23578);
and U23783 (N_23783,N_23384,N_22811);
xnor U23784 (N_23784,N_22701,N_22602);
and U23785 (N_23785,N_22613,N_23144);
nand U23786 (N_23786,N_23625,N_23447);
and U23787 (N_23787,N_22647,N_23713);
or U23788 (N_23788,N_22810,N_23243);
nor U23789 (N_23789,N_23482,N_23266);
nor U23790 (N_23790,N_23061,N_22976);
or U23791 (N_23791,N_22989,N_23164);
or U23792 (N_23792,N_23068,N_23539);
xnor U23793 (N_23793,N_23688,N_22623);
nand U23794 (N_23794,N_22951,N_23291);
and U23795 (N_23795,N_22635,N_23006);
nor U23796 (N_23796,N_22679,N_23715);
or U23797 (N_23797,N_23295,N_22715);
or U23798 (N_23798,N_22942,N_23611);
or U23799 (N_23799,N_23213,N_22966);
xor U23800 (N_23800,N_23512,N_23371);
nand U23801 (N_23801,N_23367,N_22659);
nor U23802 (N_23802,N_23383,N_23474);
and U23803 (N_23803,N_23632,N_22940);
nand U23804 (N_23804,N_23476,N_22683);
nor U23805 (N_23805,N_23662,N_23530);
and U23806 (N_23806,N_22513,N_23327);
or U23807 (N_23807,N_23260,N_23199);
or U23808 (N_23808,N_23323,N_23120);
nor U23809 (N_23809,N_22864,N_22756);
xnor U23810 (N_23810,N_23063,N_22888);
nor U23811 (N_23811,N_23262,N_23534);
and U23812 (N_23812,N_23169,N_23282);
nor U23813 (N_23813,N_23118,N_23635);
or U23814 (N_23814,N_23074,N_23087);
nor U23815 (N_23815,N_23422,N_22692);
nor U23816 (N_23816,N_23374,N_23200);
nand U23817 (N_23817,N_23234,N_22851);
nand U23818 (N_23818,N_23531,N_23108);
or U23819 (N_23819,N_22818,N_22672);
nor U23820 (N_23820,N_22639,N_23684);
nor U23821 (N_23821,N_22573,N_22977);
xnor U23822 (N_23822,N_22884,N_23370);
nor U23823 (N_23823,N_23461,N_23054);
nor U23824 (N_23824,N_23513,N_22955);
or U23825 (N_23825,N_23519,N_23137);
nand U23826 (N_23826,N_23712,N_23062);
nand U23827 (N_23827,N_23022,N_22925);
and U23828 (N_23828,N_23175,N_23640);
nand U23829 (N_23829,N_22935,N_22693);
and U23830 (N_23830,N_23096,N_22532);
and U23831 (N_23831,N_23280,N_23702);
and U23832 (N_23832,N_23723,N_23010);
xnor U23833 (N_23833,N_23523,N_23636);
xnor U23834 (N_23834,N_22800,N_23703);
and U23835 (N_23835,N_23650,N_22739);
xnor U23836 (N_23836,N_22606,N_23509);
nand U23837 (N_23837,N_23221,N_22644);
or U23838 (N_23838,N_23709,N_23669);
and U23839 (N_23839,N_23205,N_22958);
nand U23840 (N_23840,N_23112,N_23456);
and U23841 (N_23841,N_23434,N_23585);
xor U23842 (N_23842,N_23554,N_23599);
nand U23843 (N_23843,N_22719,N_22963);
and U23844 (N_23844,N_22569,N_23073);
nor U23845 (N_23845,N_23146,N_23608);
and U23846 (N_23846,N_23267,N_23612);
nand U23847 (N_23847,N_23239,N_23748);
and U23848 (N_23848,N_23457,N_22559);
and U23849 (N_23849,N_23522,N_23437);
or U23850 (N_23850,N_22819,N_22952);
xnor U23851 (N_23851,N_22831,N_22770);
and U23852 (N_23852,N_23587,N_23423);
or U23853 (N_23853,N_23240,N_22789);
xnor U23854 (N_23854,N_23397,N_23095);
xor U23855 (N_23855,N_23029,N_23592);
or U23856 (N_23856,N_23046,N_23244);
nor U23857 (N_23857,N_23580,N_23644);
and U23858 (N_23858,N_23499,N_23528);
nor U23859 (N_23859,N_23495,N_22993);
and U23860 (N_23860,N_22678,N_23679);
xor U23861 (N_23861,N_23518,N_23288);
xnor U23862 (N_23862,N_22540,N_22907);
and U23863 (N_23863,N_22593,N_23372);
xnor U23864 (N_23864,N_23100,N_23224);
and U23865 (N_23865,N_23363,N_23607);
xnor U23866 (N_23866,N_23634,N_22944);
nand U23867 (N_23867,N_23716,N_23107);
and U23868 (N_23868,N_22664,N_23188);
nand U23869 (N_23869,N_22790,N_22724);
nand U23870 (N_23870,N_23093,N_23223);
and U23871 (N_23871,N_22852,N_23717);
nand U23872 (N_23872,N_23392,N_22933);
and U23873 (N_23873,N_23119,N_22731);
nand U23874 (N_23874,N_22759,N_22954);
xnor U23875 (N_23875,N_22805,N_23140);
and U23876 (N_23876,N_22938,N_23511);
and U23877 (N_23877,N_23695,N_23336);
xnor U23878 (N_23878,N_22558,N_23049);
nor U23879 (N_23879,N_22533,N_23352);
nor U23880 (N_23880,N_22514,N_23744);
nor U23881 (N_23881,N_23572,N_23211);
nor U23882 (N_23882,N_23448,N_23517);
or U23883 (N_23883,N_23331,N_23203);
or U23884 (N_23884,N_23614,N_23685);
and U23885 (N_23885,N_23719,N_22974);
nand U23886 (N_23886,N_23590,N_23738);
and U23887 (N_23887,N_22837,N_23086);
nor U23888 (N_23888,N_23017,N_22791);
nor U23889 (N_23889,N_22971,N_23693);
nand U23890 (N_23890,N_22537,N_23160);
or U23891 (N_23891,N_22892,N_23013);
nand U23892 (N_23892,N_23193,N_23305);
nor U23893 (N_23893,N_23314,N_23268);
xor U23894 (N_23894,N_23273,N_23341);
and U23895 (N_23895,N_23402,N_22717);
or U23896 (N_23896,N_22661,N_23003);
xnor U23897 (N_23897,N_22516,N_22917);
and U23898 (N_23898,N_23251,N_23056);
or U23899 (N_23899,N_23181,N_23230);
xor U23900 (N_23900,N_22667,N_23393);
nor U23901 (N_23901,N_22640,N_23464);
and U23902 (N_23902,N_22721,N_23729);
xor U23903 (N_23903,N_23197,N_23706);
xor U23904 (N_23904,N_23092,N_22788);
nand U23905 (N_23905,N_22626,N_22707);
nand U23906 (N_23906,N_23105,N_23569);
xor U23907 (N_23907,N_23537,N_22869);
nor U23908 (N_23908,N_23035,N_22987);
nor U23909 (N_23909,N_22651,N_23508);
and U23910 (N_23910,N_23192,N_23245);
or U23911 (N_23911,N_22953,N_23225);
and U23912 (N_23912,N_23025,N_22874);
and U23913 (N_23913,N_23130,N_22865);
nand U23914 (N_23914,N_23148,N_23173);
nor U23915 (N_23915,N_23649,N_23673);
xor U23916 (N_23916,N_22657,N_23440);
and U23917 (N_23917,N_23177,N_23089);
and U23918 (N_23918,N_22700,N_23031);
nand U23919 (N_23919,N_23237,N_22745);
nor U23920 (N_23920,N_22763,N_22758);
or U23921 (N_23921,N_22821,N_22685);
xnor U23922 (N_23922,N_23732,N_22650);
or U23923 (N_23923,N_23428,N_23106);
xnor U23924 (N_23924,N_22741,N_22894);
nand U23925 (N_23925,N_22547,N_22853);
nand U23926 (N_23926,N_23222,N_23627);
and U23927 (N_23927,N_22607,N_22960);
nand U23928 (N_23928,N_22748,N_22998);
or U23929 (N_23929,N_22620,N_22530);
and U23930 (N_23930,N_23568,N_22796);
nand U23931 (N_23931,N_22591,N_23481);
nor U23932 (N_23932,N_22824,N_22630);
and U23933 (N_23933,N_23694,N_22538);
nand U23934 (N_23934,N_23598,N_23666);
and U23935 (N_23935,N_22768,N_23227);
nand U23936 (N_23936,N_23353,N_23409);
nand U23937 (N_23937,N_23308,N_23345);
and U23938 (N_23938,N_22554,N_22946);
nand U23939 (N_23939,N_23027,N_22846);
xnor U23940 (N_23940,N_22841,N_22705);
nor U23941 (N_23941,N_23149,N_22889);
nor U23942 (N_23942,N_22978,N_23139);
nand U23943 (N_23943,N_22730,N_23104);
xor U23944 (N_23944,N_23659,N_22812);
nor U23945 (N_23945,N_23090,N_22857);
nand U23946 (N_23946,N_22862,N_23171);
nand U23947 (N_23947,N_23404,N_22511);
nor U23948 (N_23948,N_22787,N_22594);
or U23949 (N_23949,N_22743,N_23670);
and U23950 (N_23950,N_22872,N_23403);
nor U23951 (N_23951,N_23651,N_23645);
and U23952 (N_23952,N_22599,N_23265);
or U23953 (N_23953,N_22930,N_22927);
and U23954 (N_23954,N_22799,N_23721);
nand U23955 (N_23955,N_23385,N_23122);
nand U23956 (N_23956,N_22820,N_23487);
nor U23957 (N_23957,N_22746,N_23593);
or U23958 (N_23958,N_23001,N_22902);
xnor U23959 (N_23959,N_22914,N_23279);
nor U23960 (N_23960,N_23080,N_22783);
nand U23961 (N_23961,N_22854,N_22997);
nor U23962 (N_23962,N_22928,N_23451);
nor U23963 (N_23963,N_23527,N_22753);
nand U23964 (N_23964,N_23128,N_22570);
nand U23965 (N_23965,N_23182,N_23011);
nand U23966 (N_23966,N_23042,N_23136);
nand U23967 (N_23967,N_22757,N_22673);
nor U23968 (N_23968,N_23418,N_23621);
nor U23969 (N_23969,N_23624,N_22595);
nand U23970 (N_23970,N_23198,N_22994);
nand U23971 (N_23971,N_23299,N_23493);
or U23972 (N_23972,N_22877,N_22718);
or U23973 (N_23973,N_23497,N_22572);
nor U23974 (N_23974,N_23015,N_22519);
nand U23975 (N_23975,N_23283,N_23084);
or U23976 (N_23976,N_22658,N_22704);
nand U23977 (N_23977,N_23480,N_23613);
nand U23978 (N_23978,N_23462,N_23272);
nand U23979 (N_23979,N_23504,N_22979);
nor U23980 (N_23980,N_23322,N_23259);
xor U23981 (N_23981,N_22712,N_23184);
or U23982 (N_23982,N_22565,N_23329);
xnor U23983 (N_23983,N_23387,N_23014);
xnor U23984 (N_23984,N_22764,N_22991);
and U23985 (N_23985,N_22567,N_23135);
nor U23986 (N_23986,N_23432,N_23053);
nor U23987 (N_23987,N_22961,N_22702);
and U23988 (N_23988,N_22992,N_22550);
or U23989 (N_23989,N_22956,N_23124);
nor U23990 (N_23990,N_23667,N_22969);
nor U23991 (N_23991,N_22713,N_23631);
nand U23992 (N_23992,N_22777,N_22840);
and U23993 (N_23993,N_23735,N_22975);
or U23994 (N_23994,N_23389,N_22562);
or U23995 (N_23995,N_22523,N_22939);
xnor U23996 (N_23996,N_23313,N_22876);
and U23997 (N_23997,N_23264,N_23442);
and U23998 (N_23998,N_23340,N_22676);
or U23999 (N_23999,N_23465,N_22868);
and U24000 (N_24000,N_23386,N_22545);
nor U24001 (N_24001,N_23172,N_22897);
xnor U24002 (N_24002,N_23113,N_23577);
and U24003 (N_24003,N_23471,N_23707);
and U24004 (N_24004,N_22950,N_23357);
and U24005 (N_24005,N_22866,N_23215);
nand U24006 (N_24006,N_23714,N_22849);
xnor U24007 (N_24007,N_23343,N_23085);
and U24008 (N_24008,N_23110,N_22911);
or U24009 (N_24009,N_23533,N_23454);
nor U24010 (N_24010,N_23347,N_23398);
nor U24011 (N_24011,N_23176,N_23507);
xnor U24012 (N_24012,N_23615,N_23249);
or U24013 (N_24013,N_23286,N_23258);
or U24014 (N_24014,N_23020,N_23642);
or U24015 (N_24015,N_22856,N_23241);
and U24016 (N_24016,N_22903,N_22867);
nand U24017 (N_24017,N_23475,N_23315);
and U24018 (N_24018,N_23256,N_23235);
and U24019 (N_24019,N_23505,N_23102);
nor U24020 (N_24020,N_23485,N_22541);
and U24021 (N_24021,N_23028,N_23048);
nand U24022 (N_24022,N_23668,N_23316);
or U24023 (N_24023,N_22656,N_22668);
nor U24024 (N_24024,N_22909,N_23697);
nand U24025 (N_24025,N_23510,N_22531);
and U24026 (N_24026,N_22959,N_22674);
xor U24027 (N_24027,N_23333,N_22948);
and U24028 (N_24028,N_22870,N_23362);
nand U24029 (N_24029,N_22551,N_23351);
xnor U24030 (N_24030,N_22905,N_22699);
nand U24031 (N_24031,N_22742,N_23562);
xor U24032 (N_24032,N_22931,N_23247);
nand U24033 (N_24033,N_23604,N_23620);
or U24034 (N_24034,N_23538,N_23725);
nand U24035 (N_24035,N_23747,N_23097);
and U24036 (N_24036,N_22728,N_23705);
and U24037 (N_24037,N_22807,N_23421);
or U24038 (N_24038,N_23233,N_23276);
xor U24039 (N_24039,N_23318,N_23559);
or U24040 (N_24040,N_22826,N_22798);
nand U24041 (N_24041,N_23444,N_23154);
xor U24042 (N_24042,N_22848,N_23129);
xnor U24043 (N_24043,N_22827,N_23115);
or U24044 (N_24044,N_23180,N_23582);
and U24045 (N_24045,N_22813,N_23629);
nand U24046 (N_24046,N_23731,N_23525);
and U24047 (N_24047,N_23478,N_22614);
nand U24048 (N_24048,N_22703,N_23382);
nor U24049 (N_24049,N_22654,N_23255);
and U24050 (N_24050,N_23134,N_23220);
or U24051 (N_24051,N_23532,N_23745);
xnor U24052 (N_24052,N_23228,N_23066);
and U24053 (N_24053,N_22898,N_22611);
or U24054 (N_24054,N_22609,N_22887);
nor U24055 (N_24055,N_23596,N_23021);
and U24056 (N_24056,N_23473,N_22871);
xor U24057 (N_24057,N_23378,N_23459);
xor U24058 (N_24058,N_23346,N_23676);
or U24059 (N_24059,N_22795,N_23032);
or U24060 (N_24060,N_23064,N_22710);
nand U24061 (N_24061,N_22687,N_23242);
nand U24062 (N_24062,N_22920,N_23655);
xor U24063 (N_24063,N_23401,N_23069);
xor U24064 (N_24064,N_22643,N_23567);
nor U24065 (N_24065,N_23253,N_22502);
nand U24066 (N_24066,N_22528,N_22981);
nand U24067 (N_24067,N_22581,N_22906);
nand U24068 (N_24068,N_23167,N_22968);
xor U24069 (N_24069,N_22553,N_23565);
xor U24070 (N_24070,N_23257,N_22624);
xor U24071 (N_24071,N_22814,N_22843);
and U24072 (N_24072,N_23406,N_23236);
and U24073 (N_24073,N_22964,N_23541);
and U24074 (N_24074,N_23369,N_22566);
nor U24075 (N_24075,N_22904,N_23388);
nor U24076 (N_24076,N_22973,N_23639);
nand U24077 (N_24077,N_23289,N_22793);
or U24078 (N_24078,N_22586,N_23036);
and U24079 (N_24079,N_22901,N_22601);
or U24080 (N_24080,N_23012,N_22563);
and U24081 (N_24081,N_22524,N_23326);
nor U24082 (N_24082,N_23157,N_23166);
or U24083 (N_24083,N_23296,N_22855);
or U24084 (N_24084,N_22589,N_23573);
or U24085 (N_24085,N_23571,N_23652);
nand U24086 (N_24086,N_23252,N_23689);
nand U24087 (N_24087,N_22934,N_23526);
nor U24088 (N_24088,N_23678,N_22803);
nand U24089 (N_24089,N_23337,N_22766);
nor U24090 (N_24090,N_23151,N_22801);
and U24091 (N_24091,N_22750,N_22875);
nor U24092 (N_24092,N_22886,N_23628);
xor U24093 (N_24093,N_23656,N_23588);
nor U24094 (N_24094,N_23324,N_23502);
and U24095 (N_24095,N_22548,N_23396);
and U24096 (N_24096,N_22680,N_23007);
or U24097 (N_24097,N_23033,N_23165);
xnor U24098 (N_24098,N_23566,N_23359);
or U24099 (N_24099,N_23209,N_23037);
and U24100 (N_24100,N_22794,N_23647);
xnor U24101 (N_24101,N_23041,N_22631);
nor U24102 (N_24102,N_23285,N_22652);
nor U24103 (N_24103,N_23501,N_22600);
xnor U24104 (N_24104,N_23202,N_22629);
nor U24105 (N_24105,N_22633,N_23034);
or U24106 (N_24106,N_23619,N_22833);
nand U24107 (N_24107,N_23099,N_23414);
and U24108 (N_24108,N_23292,N_22937);
or U24109 (N_24109,N_23736,N_22949);
nor U24110 (N_24110,N_23680,N_23616);
nand U24111 (N_24111,N_23186,N_22546);
nor U24112 (N_24112,N_22891,N_23297);
nand U24113 (N_24113,N_22690,N_23179);
xnor U24114 (N_24114,N_22815,N_23116);
and U24115 (N_24115,N_23556,N_23605);
or U24116 (N_24116,N_23319,N_22564);
and U24117 (N_24117,N_23563,N_22618);
nand U24118 (N_24118,N_23681,N_22544);
nand U24119 (N_24119,N_23226,N_22832);
nor U24120 (N_24120,N_22555,N_22655);
and U24121 (N_24121,N_23366,N_23178);
or U24122 (N_24122,N_22665,N_23690);
or U24123 (N_24123,N_22785,N_22571);
or U24124 (N_24124,N_23091,N_23420);
nand U24125 (N_24125,N_23379,N_23741);
or U24126 (N_24126,N_22878,N_23399);
nor U24127 (N_24127,N_23094,N_23489);
nor U24128 (N_24128,N_22579,N_22515);
or U24129 (N_24129,N_22711,N_22649);
and U24130 (N_24130,N_23483,N_23310);
nor U24131 (N_24131,N_22781,N_23380);
xor U24132 (N_24132,N_23597,N_23138);
nor U24133 (N_24133,N_23433,N_23121);
xor U24134 (N_24134,N_23536,N_22714);
or U24135 (N_24135,N_23158,N_23708);
nand U24136 (N_24136,N_23131,N_22536);
nand U24137 (N_24137,N_22772,N_23743);
or U24138 (N_24138,N_23381,N_22587);
and U24139 (N_24139,N_22873,N_23558);
and U24140 (N_24140,N_22597,N_22642);
nand U24141 (N_24141,N_22808,N_23275);
nor U24142 (N_24142,N_23038,N_23412);
and U24143 (N_24143,N_23334,N_23060);
xor U24144 (N_24144,N_22980,N_23304);
nor U24145 (N_24145,N_23349,N_22771);
xor U24146 (N_24146,N_22529,N_22988);
and U24147 (N_24147,N_22535,N_23610);
and U24148 (N_24148,N_22984,N_23663);
xor U24149 (N_24149,N_23000,N_22996);
nand U24150 (N_24150,N_23698,N_23737);
nand U24151 (N_24151,N_23579,N_23147);
nor U24152 (N_24152,N_23687,N_23111);
nor U24153 (N_24153,N_23691,N_23692);
and U24154 (N_24154,N_22720,N_22776);
nand U24155 (N_24155,N_22592,N_23549);
nand U24156 (N_24156,N_23075,N_22924);
nor U24157 (N_24157,N_22972,N_23330);
and U24158 (N_24158,N_23638,N_23051);
and U24159 (N_24159,N_22695,N_23312);
nor U24160 (N_24160,N_23602,N_22842);
nand U24161 (N_24161,N_22706,N_23187);
nand U24162 (N_24162,N_22726,N_22986);
xnor U24163 (N_24163,N_23270,N_22522);
and U24164 (N_24164,N_22520,N_22542);
nand U24165 (N_24165,N_22723,N_22694);
xnor U24166 (N_24166,N_22893,N_22754);
xnor U24167 (N_24167,N_23545,N_22835);
xnor U24168 (N_24168,N_22580,N_22967);
nand U24169 (N_24169,N_23600,N_23293);
nand U24170 (N_24170,N_23699,N_22575);
xor U24171 (N_24171,N_23281,N_22637);
nand U24172 (N_24172,N_23492,N_23088);
nor U24173 (N_24173,N_23059,N_22709);
xnor U24174 (N_24174,N_22918,N_22834);
or U24175 (N_24175,N_22850,N_22778);
or U24176 (N_24176,N_23626,N_22863);
and U24177 (N_24177,N_23005,N_23443);
nand U24178 (N_24178,N_22929,N_22504);
xnor U24179 (N_24179,N_22751,N_23637);
nand U24180 (N_24180,N_23101,N_23133);
nand U24181 (N_24181,N_23643,N_23376);
or U24182 (N_24182,N_23077,N_23019);
or U24183 (N_24183,N_23039,N_22666);
and U24184 (N_24184,N_23561,N_23395);
and U24185 (N_24185,N_23302,N_23219);
nand U24186 (N_24186,N_22527,N_23163);
nor U24187 (N_24187,N_23328,N_23057);
or U24188 (N_24188,N_23439,N_22671);
or U24189 (N_24189,N_23229,N_22749);
nand U24190 (N_24190,N_23294,N_23425);
nor U24191 (N_24191,N_22895,N_23132);
nand U24192 (N_24192,N_22557,N_23496);
nor U24193 (N_24193,N_22500,N_23472);
or U24194 (N_24194,N_23682,N_23018);
nand U24195 (N_24195,N_23653,N_22779);
nand U24196 (N_24196,N_23467,N_23026);
nor U24197 (N_24197,N_23606,N_23045);
xnor U24198 (N_24198,N_22823,N_23739);
xor U24199 (N_24199,N_23514,N_23044);
nor U24200 (N_24200,N_23664,N_22510);
xor U24201 (N_24201,N_22646,N_22638);
nand U24202 (N_24202,N_23072,N_22932);
or U24203 (N_24203,N_23413,N_23400);
and U24204 (N_24204,N_23390,N_23591);
xnor U24205 (N_24205,N_23141,N_22825);
and U24206 (N_24206,N_22615,N_23441);
xor U24207 (N_24207,N_23491,N_23127);
nand U24208 (N_24208,N_23117,N_23557);
nor U24209 (N_24209,N_23658,N_23430);
xor U24210 (N_24210,N_23633,N_23191);
xor U24211 (N_24211,N_22521,N_23581);
and U24212 (N_24212,N_22560,N_22985);
or U24213 (N_24213,N_22585,N_22921);
and U24214 (N_24214,N_23231,N_23701);
xnor U24215 (N_24215,N_22681,N_22784);
or U24216 (N_24216,N_23161,N_22735);
or U24217 (N_24217,N_23583,N_23520);
nor U24218 (N_24218,N_22919,N_22608);
nand U24219 (N_24219,N_22675,N_22744);
nand U24220 (N_24220,N_23575,N_23544);
nand U24221 (N_24221,N_23189,N_23217);
xnor U24222 (N_24222,N_23551,N_23468);
or U24223 (N_24223,N_22619,N_23317);
or U24224 (N_24224,N_23617,N_22577);
xor U24225 (N_24225,N_23307,N_23123);
or U24226 (N_24226,N_23734,N_23446);
nor U24227 (N_24227,N_22830,N_23603);
xor U24228 (N_24228,N_22578,N_22755);
nor U24229 (N_24229,N_22908,N_22636);
nor U24230 (N_24230,N_23082,N_23070);
nor U24231 (N_24231,N_22583,N_23661);
or U24232 (N_24232,N_23419,N_23306);
xor U24233 (N_24233,N_23546,N_23067);
xnor U24234 (N_24234,N_23728,N_23065);
nor U24235 (N_24235,N_23553,N_22588);
xnor U24236 (N_24236,N_23309,N_23208);
xnor U24237 (N_24237,N_23429,N_23250);
nand U24238 (N_24238,N_22610,N_23426);
xor U24239 (N_24239,N_23550,N_23263);
nand U24240 (N_24240,N_23675,N_23004);
nand U24241 (N_24241,N_23354,N_23515);
xor U24242 (N_24242,N_23365,N_23641);
or U24243 (N_24243,N_22734,N_23740);
or U24244 (N_24244,N_22733,N_22844);
and U24245 (N_24245,N_22797,N_22663);
or U24246 (N_24246,N_23356,N_23190);
or U24247 (N_24247,N_22767,N_23325);
nand U24248 (N_24248,N_23078,N_22861);
or U24249 (N_24249,N_23646,N_23156);
or U24250 (N_24250,N_23271,N_22765);
or U24251 (N_24251,N_23623,N_23677);
or U24252 (N_24252,N_22732,N_22627);
or U24253 (N_24253,N_23023,N_22738);
xnor U24254 (N_24254,N_23071,N_23142);
and U24255 (N_24255,N_23730,N_23560);
or U24256 (N_24256,N_22922,N_23269);
xor U24257 (N_24257,N_22603,N_23047);
nand U24258 (N_24258,N_23206,N_22737);
nand U24259 (N_24259,N_22883,N_23435);
or U24260 (N_24260,N_22775,N_22604);
or U24261 (N_24261,N_23055,N_23564);
xnor U24262 (N_24262,N_23455,N_22617);
and U24263 (N_24263,N_22729,N_22983);
nand U24264 (N_24264,N_23076,N_22605);
and U24265 (N_24265,N_23452,N_22804);
nor U24266 (N_24266,N_23321,N_22970);
nor U24267 (N_24267,N_23368,N_23301);
xnor U24268 (N_24268,N_22686,N_22802);
xor U24269 (N_24269,N_23043,N_23150);
nand U24270 (N_24270,N_22598,N_23686);
nor U24271 (N_24271,N_23488,N_22990);
xnor U24272 (N_24272,N_22747,N_22660);
xor U24273 (N_24273,N_22761,N_23339);
xor U24274 (N_24274,N_23348,N_22645);
and U24275 (N_24275,N_22780,N_23630);
or U24276 (N_24276,N_23665,N_23574);
nand U24277 (N_24277,N_23427,N_22806);
nor U24278 (N_24278,N_23722,N_22689);
xor U24279 (N_24279,N_23284,N_23303);
and U24280 (N_24280,N_23424,N_23159);
xnor U24281 (N_24281,N_23350,N_23718);
nor U24282 (N_24282,N_23733,N_22822);
or U24283 (N_24283,N_23050,N_23595);
or U24284 (N_24284,N_23540,N_23524);
nand U24285 (N_24285,N_23212,N_23232);
and U24286 (N_24286,N_23470,N_22957);
xor U24287 (N_24287,N_23081,N_22501);
and U24288 (N_24288,N_23210,N_23469);
nand U24289 (N_24289,N_22670,N_23394);
xor U24290 (N_24290,N_22926,N_23727);
or U24291 (N_24291,N_22896,N_23449);
nand U24292 (N_24292,N_23373,N_23355);
or U24293 (N_24293,N_23408,N_23618);
xnor U24294 (N_24294,N_23589,N_23479);
xnor U24295 (N_24295,N_22882,N_22543);
and U24296 (N_24296,N_23332,N_23375);
or U24297 (N_24297,N_23168,N_23503);
and U24298 (N_24298,N_23683,N_23052);
or U24299 (N_24299,N_22549,N_22708);
or U24300 (N_24300,N_23710,N_22677);
and U24301 (N_24301,N_22792,N_22725);
or U24302 (N_24302,N_23335,N_22774);
nand U24303 (N_24303,N_23570,N_23529);
or U24304 (N_24304,N_23622,N_22503);
xor U24305 (N_24305,N_23711,N_23358);
nor U24306 (N_24306,N_23145,N_23547);
nand U24307 (N_24307,N_22568,N_23360);
nor U24308 (N_24308,N_23660,N_23125);
and U24309 (N_24309,N_23277,N_23002);
nor U24310 (N_24310,N_22561,N_23506);
nand U24311 (N_24311,N_23153,N_23486);
xnor U24312 (N_24312,N_22518,N_23704);
and U24313 (N_24313,N_23458,N_22653);
and U24314 (N_24314,N_22628,N_23555);
xor U24315 (N_24315,N_23584,N_22632);
xnor U24316 (N_24316,N_22622,N_23216);
nor U24317 (N_24317,N_22552,N_23436);
nand U24318 (N_24318,N_22913,N_23466);
xnor U24319 (N_24319,N_23204,N_23416);
nand U24320 (N_24320,N_23484,N_23749);
or U24321 (N_24321,N_23410,N_23174);
nand U24322 (N_24322,N_23417,N_23300);
nand U24323 (N_24323,N_22947,N_22526);
and U24324 (N_24324,N_22829,N_22534);
xnor U24325 (N_24325,N_23521,N_23535);
or U24326 (N_24326,N_23746,N_22817);
or U24327 (N_24327,N_23344,N_23654);
nor U24328 (N_24328,N_22740,N_22773);
nor U24329 (N_24329,N_23548,N_22880);
or U24330 (N_24330,N_23254,N_22682);
and U24331 (N_24331,N_23320,N_22507);
and U24332 (N_24332,N_22506,N_22769);
xor U24333 (N_24333,N_22574,N_23576);
or U24334 (N_24334,N_22982,N_22900);
and U24335 (N_24335,N_23126,N_23674);
xnor U24336 (N_24336,N_23361,N_23405);
xor U24337 (N_24337,N_22509,N_23183);
nand U24338 (N_24338,N_22641,N_23218);
nor U24339 (N_24339,N_22505,N_23196);
xnor U24340 (N_24340,N_23024,N_23700);
or U24341 (N_24341,N_22752,N_23542);
xor U24342 (N_24342,N_23155,N_23498);
or U24343 (N_24343,N_23657,N_22859);
nand U24344 (N_24344,N_23214,N_23450);
or U24345 (N_24345,N_22691,N_22512);
xor U24346 (N_24346,N_23207,N_22912);
nand U24347 (N_24347,N_23009,N_22890);
nand U24348 (N_24348,N_23696,N_22995);
nand U24349 (N_24349,N_23278,N_23415);
nand U24350 (N_24350,N_22590,N_23058);
nor U24351 (N_24351,N_23671,N_22525);
xnor U24352 (N_24352,N_23377,N_22847);
nand U24353 (N_24353,N_22539,N_22625);
xor U24354 (N_24354,N_23143,N_23016);
or U24355 (N_24355,N_23460,N_22684);
nand U24356 (N_24356,N_23391,N_23609);
nand U24357 (N_24357,N_22648,N_23287);
and U24358 (N_24358,N_23494,N_22669);
or U24359 (N_24359,N_22860,N_22727);
or U24360 (N_24360,N_23594,N_23008);
nor U24361 (N_24361,N_23298,N_23311);
xor U24362 (N_24362,N_23543,N_22916);
nand U24363 (N_24363,N_23238,N_22697);
nor U24364 (N_24364,N_23248,N_22838);
nor U24365 (N_24365,N_22816,N_23103);
and U24366 (N_24366,N_23342,N_22634);
nor U24367 (N_24367,N_23194,N_23098);
nor U24368 (N_24368,N_23083,N_22943);
or U24369 (N_24369,N_22722,N_23274);
and U24370 (N_24370,N_22688,N_23246);
and U24371 (N_24371,N_23079,N_23152);
nor U24372 (N_24372,N_22828,N_23185);
nand U24373 (N_24373,N_22508,N_23411);
or U24374 (N_24374,N_22736,N_23648);
or U24375 (N_24375,N_22613,N_22989);
and U24376 (N_24376,N_23263,N_23689);
nor U24377 (N_24377,N_23069,N_22806);
nand U24378 (N_24378,N_22780,N_22972);
and U24379 (N_24379,N_23061,N_23663);
or U24380 (N_24380,N_23327,N_22734);
nand U24381 (N_24381,N_23223,N_23256);
nor U24382 (N_24382,N_22904,N_22996);
nand U24383 (N_24383,N_22511,N_23194);
nor U24384 (N_24384,N_22971,N_23663);
nor U24385 (N_24385,N_23053,N_22581);
xor U24386 (N_24386,N_22821,N_23723);
nor U24387 (N_24387,N_23235,N_23091);
nor U24388 (N_24388,N_22903,N_23479);
or U24389 (N_24389,N_23713,N_23200);
or U24390 (N_24390,N_23248,N_23708);
nand U24391 (N_24391,N_23416,N_23249);
nand U24392 (N_24392,N_23010,N_23622);
xor U24393 (N_24393,N_22719,N_22502);
nor U24394 (N_24394,N_23265,N_22615);
xnor U24395 (N_24395,N_22768,N_22503);
or U24396 (N_24396,N_23680,N_23625);
nor U24397 (N_24397,N_23354,N_23195);
nor U24398 (N_24398,N_22939,N_23080);
and U24399 (N_24399,N_23308,N_23213);
or U24400 (N_24400,N_23562,N_22833);
nand U24401 (N_24401,N_23208,N_23494);
and U24402 (N_24402,N_23413,N_23615);
and U24403 (N_24403,N_23160,N_23450);
nand U24404 (N_24404,N_22735,N_22668);
xnor U24405 (N_24405,N_22716,N_23635);
nor U24406 (N_24406,N_23284,N_23718);
and U24407 (N_24407,N_23038,N_23442);
nor U24408 (N_24408,N_23306,N_23665);
xor U24409 (N_24409,N_23701,N_23175);
or U24410 (N_24410,N_23400,N_22514);
xor U24411 (N_24411,N_22937,N_22908);
nor U24412 (N_24412,N_23019,N_23379);
or U24413 (N_24413,N_23360,N_23569);
or U24414 (N_24414,N_22819,N_22995);
or U24415 (N_24415,N_23099,N_22643);
and U24416 (N_24416,N_22798,N_22933);
and U24417 (N_24417,N_23525,N_23092);
or U24418 (N_24418,N_23108,N_23158);
and U24419 (N_24419,N_23033,N_23120);
and U24420 (N_24420,N_23419,N_23165);
xnor U24421 (N_24421,N_22769,N_23541);
and U24422 (N_24422,N_22633,N_23380);
nor U24423 (N_24423,N_22738,N_22540);
nand U24424 (N_24424,N_22555,N_23682);
nor U24425 (N_24425,N_23322,N_22920);
or U24426 (N_24426,N_23348,N_23035);
xor U24427 (N_24427,N_22759,N_23423);
xnor U24428 (N_24428,N_22572,N_22893);
nand U24429 (N_24429,N_23306,N_23125);
xnor U24430 (N_24430,N_23136,N_22644);
nand U24431 (N_24431,N_23289,N_23173);
nand U24432 (N_24432,N_22880,N_23547);
and U24433 (N_24433,N_23474,N_23324);
or U24434 (N_24434,N_22660,N_22952);
xnor U24435 (N_24435,N_22901,N_23009);
and U24436 (N_24436,N_23011,N_23302);
or U24437 (N_24437,N_23507,N_22626);
nor U24438 (N_24438,N_23362,N_23220);
or U24439 (N_24439,N_22778,N_23562);
nand U24440 (N_24440,N_23375,N_23292);
or U24441 (N_24441,N_23463,N_22770);
or U24442 (N_24442,N_22856,N_23193);
nor U24443 (N_24443,N_23079,N_23163);
xnor U24444 (N_24444,N_23391,N_23129);
or U24445 (N_24445,N_22984,N_23007);
nor U24446 (N_24446,N_22918,N_23028);
xnor U24447 (N_24447,N_22512,N_22947);
nand U24448 (N_24448,N_23728,N_23156);
xnor U24449 (N_24449,N_23643,N_23571);
xor U24450 (N_24450,N_23152,N_22938);
xnor U24451 (N_24451,N_22818,N_23745);
xnor U24452 (N_24452,N_23031,N_22854);
or U24453 (N_24453,N_23222,N_23375);
or U24454 (N_24454,N_23298,N_23303);
or U24455 (N_24455,N_22896,N_23657);
nor U24456 (N_24456,N_23487,N_22575);
nand U24457 (N_24457,N_22831,N_22726);
nor U24458 (N_24458,N_22973,N_23667);
xor U24459 (N_24459,N_23703,N_23117);
nand U24460 (N_24460,N_23044,N_23145);
and U24461 (N_24461,N_23603,N_23535);
or U24462 (N_24462,N_23289,N_22811);
or U24463 (N_24463,N_23510,N_22863);
xor U24464 (N_24464,N_22790,N_22922);
nor U24465 (N_24465,N_22684,N_22676);
and U24466 (N_24466,N_23148,N_23648);
nand U24467 (N_24467,N_23350,N_22544);
and U24468 (N_24468,N_23010,N_23688);
or U24469 (N_24469,N_22812,N_23299);
and U24470 (N_24470,N_22854,N_22620);
or U24471 (N_24471,N_23250,N_23438);
xor U24472 (N_24472,N_22703,N_23028);
nand U24473 (N_24473,N_23123,N_23020);
xnor U24474 (N_24474,N_23379,N_23040);
nand U24475 (N_24475,N_22705,N_23524);
xor U24476 (N_24476,N_22948,N_23746);
or U24477 (N_24477,N_22876,N_22827);
and U24478 (N_24478,N_23625,N_23265);
nand U24479 (N_24479,N_23195,N_23392);
nand U24480 (N_24480,N_23174,N_22607);
or U24481 (N_24481,N_22759,N_23529);
and U24482 (N_24482,N_22856,N_23077);
xnor U24483 (N_24483,N_23404,N_23418);
and U24484 (N_24484,N_22887,N_23512);
nand U24485 (N_24485,N_22746,N_23405);
or U24486 (N_24486,N_23334,N_22835);
nand U24487 (N_24487,N_23380,N_22535);
or U24488 (N_24488,N_23581,N_23711);
or U24489 (N_24489,N_23213,N_22942);
nor U24490 (N_24490,N_22955,N_23112);
nand U24491 (N_24491,N_23282,N_23349);
xor U24492 (N_24492,N_22708,N_23388);
xnor U24493 (N_24493,N_22784,N_23606);
nand U24494 (N_24494,N_23148,N_22896);
or U24495 (N_24495,N_23517,N_23726);
nand U24496 (N_24496,N_23146,N_22643);
or U24497 (N_24497,N_22691,N_23557);
nand U24498 (N_24498,N_22830,N_22793);
nor U24499 (N_24499,N_22777,N_22505);
nand U24500 (N_24500,N_22960,N_23542);
or U24501 (N_24501,N_22863,N_23649);
or U24502 (N_24502,N_23678,N_22854);
xor U24503 (N_24503,N_23295,N_22542);
nor U24504 (N_24504,N_22525,N_23284);
and U24505 (N_24505,N_23043,N_23402);
nand U24506 (N_24506,N_23454,N_22839);
nand U24507 (N_24507,N_22961,N_22939);
nor U24508 (N_24508,N_23530,N_23567);
nand U24509 (N_24509,N_23536,N_23365);
nand U24510 (N_24510,N_23321,N_22923);
nand U24511 (N_24511,N_23129,N_23356);
xnor U24512 (N_24512,N_22714,N_22685);
nor U24513 (N_24513,N_22852,N_23401);
nor U24514 (N_24514,N_22808,N_22693);
or U24515 (N_24515,N_22625,N_23580);
xor U24516 (N_24516,N_22650,N_22801);
xnor U24517 (N_24517,N_22597,N_23425);
or U24518 (N_24518,N_22662,N_23227);
nand U24519 (N_24519,N_23503,N_23417);
or U24520 (N_24520,N_23073,N_23028);
and U24521 (N_24521,N_22505,N_22978);
or U24522 (N_24522,N_22756,N_23364);
xnor U24523 (N_24523,N_22971,N_22815);
or U24524 (N_24524,N_23463,N_23161);
xor U24525 (N_24525,N_22796,N_22625);
nor U24526 (N_24526,N_23254,N_23470);
nor U24527 (N_24527,N_23395,N_22663);
nand U24528 (N_24528,N_23262,N_23577);
xnor U24529 (N_24529,N_23574,N_22767);
nor U24530 (N_24530,N_22634,N_23748);
nor U24531 (N_24531,N_22735,N_23113);
nor U24532 (N_24532,N_23253,N_23587);
nor U24533 (N_24533,N_22754,N_23483);
xor U24534 (N_24534,N_23637,N_22589);
xor U24535 (N_24535,N_23546,N_23519);
and U24536 (N_24536,N_22879,N_23422);
nor U24537 (N_24537,N_23019,N_23179);
or U24538 (N_24538,N_22972,N_23429);
nand U24539 (N_24539,N_22865,N_23305);
nor U24540 (N_24540,N_23370,N_22921);
xnor U24541 (N_24541,N_22706,N_23173);
nor U24542 (N_24542,N_22892,N_23081);
nand U24543 (N_24543,N_22893,N_23507);
and U24544 (N_24544,N_22869,N_22532);
or U24545 (N_24545,N_23346,N_23161);
or U24546 (N_24546,N_22737,N_23622);
nor U24547 (N_24547,N_23380,N_23731);
or U24548 (N_24548,N_22960,N_23118);
xnor U24549 (N_24549,N_23094,N_22518);
nand U24550 (N_24550,N_23487,N_23307);
nor U24551 (N_24551,N_22553,N_22837);
or U24552 (N_24552,N_23665,N_23301);
nand U24553 (N_24553,N_22864,N_22760);
xor U24554 (N_24554,N_22565,N_23115);
nand U24555 (N_24555,N_23259,N_23131);
or U24556 (N_24556,N_22896,N_22648);
nor U24557 (N_24557,N_22626,N_22702);
and U24558 (N_24558,N_23733,N_23191);
nor U24559 (N_24559,N_23008,N_23721);
or U24560 (N_24560,N_22518,N_23338);
nand U24561 (N_24561,N_23098,N_23006);
xor U24562 (N_24562,N_22537,N_23264);
xor U24563 (N_24563,N_23392,N_23226);
xnor U24564 (N_24564,N_23288,N_23040);
nand U24565 (N_24565,N_22608,N_22537);
and U24566 (N_24566,N_23022,N_23457);
or U24567 (N_24567,N_22995,N_23085);
nor U24568 (N_24568,N_23671,N_23683);
and U24569 (N_24569,N_23700,N_23629);
xnor U24570 (N_24570,N_23478,N_23664);
nand U24571 (N_24571,N_23693,N_23566);
or U24572 (N_24572,N_23510,N_23524);
xor U24573 (N_24573,N_23475,N_22656);
or U24574 (N_24574,N_22721,N_22640);
or U24575 (N_24575,N_22573,N_23531);
xnor U24576 (N_24576,N_23196,N_23620);
or U24577 (N_24577,N_23575,N_22861);
xor U24578 (N_24578,N_23326,N_23282);
xor U24579 (N_24579,N_23603,N_23407);
xor U24580 (N_24580,N_23663,N_23377);
xor U24581 (N_24581,N_23690,N_23619);
nor U24582 (N_24582,N_22746,N_23095);
and U24583 (N_24583,N_23634,N_23496);
and U24584 (N_24584,N_23013,N_23376);
nor U24585 (N_24585,N_22723,N_22767);
nor U24586 (N_24586,N_22929,N_22837);
and U24587 (N_24587,N_22698,N_23398);
nor U24588 (N_24588,N_23491,N_23123);
and U24589 (N_24589,N_22520,N_22680);
nor U24590 (N_24590,N_23625,N_22858);
or U24591 (N_24591,N_23666,N_23739);
and U24592 (N_24592,N_23333,N_23162);
and U24593 (N_24593,N_22891,N_22910);
nor U24594 (N_24594,N_23293,N_22643);
nand U24595 (N_24595,N_23082,N_22873);
xnor U24596 (N_24596,N_23406,N_23635);
and U24597 (N_24597,N_22652,N_23141);
nand U24598 (N_24598,N_23491,N_22525);
and U24599 (N_24599,N_22973,N_23027);
nand U24600 (N_24600,N_22850,N_23130);
or U24601 (N_24601,N_23105,N_22699);
xor U24602 (N_24602,N_23254,N_23198);
or U24603 (N_24603,N_23589,N_23266);
nand U24604 (N_24604,N_23276,N_23526);
nor U24605 (N_24605,N_23714,N_23381);
and U24606 (N_24606,N_22627,N_23345);
and U24607 (N_24607,N_22571,N_23415);
nor U24608 (N_24608,N_23318,N_22968);
xor U24609 (N_24609,N_22816,N_23545);
nand U24610 (N_24610,N_23696,N_22762);
xnor U24611 (N_24611,N_22830,N_23451);
nor U24612 (N_24612,N_22997,N_22830);
and U24613 (N_24613,N_22516,N_22770);
xor U24614 (N_24614,N_22965,N_22777);
nor U24615 (N_24615,N_23725,N_22930);
xor U24616 (N_24616,N_23629,N_23251);
nand U24617 (N_24617,N_22842,N_23160);
xor U24618 (N_24618,N_23737,N_23648);
or U24619 (N_24619,N_23096,N_22655);
nand U24620 (N_24620,N_23729,N_22804);
xnor U24621 (N_24621,N_23109,N_22791);
nand U24622 (N_24622,N_22788,N_22721);
nand U24623 (N_24623,N_23599,N_22586);
and U24624 (N_24624,N_22759,N_23306);
nor U24625 (N_24625,N_23099,N_23357);
nand U24626 (N_24626,N_23613,N_23744);
xnor U24627 (N_24627,N_22815,N_22979);
xnor U24628 (N_24628,N_22664,N_23722);
xor U24629 (N_24629,N_23398,N_22600);
nor U24630 (N_24630,N_23147,N_23038);
and U24631 (N_24631,N_23060,N_23115);
nand U24632 (N_24632,N_23474,N_23636);
or U24633 (N_24633,N_23561,N_23411);
nand U24634 (N_24634,N_22933,N_22569);
nand U24635 (N_24635,N_23084,N_22574);
and U24636 (N_24636,N_23154,N_23382);
and U24637 (N_24637,N_23469,N_23199);
xor U24638 (N_24638,N_23361,N_22955);
and U24639 (N_24639,N_23035,N_22629);
nand U24640 (N_24640,N_22694,N_22713);
and U24641 (N_24641,N_23194,N_23598);
xnor U24642 (N_24642,N_22681,N_23552);
xnor U24643 (N_24643,N_22785,N_22753);
xor U24644 (N_24644,N_23205,N_23669);
nand U24645 (N_24645,N_23662,N_22844);
nor U24646 (N_24646,N_23023,N_23331);
or U24647 (N_24647,N_23410,N_23521);
nor U24648 (N_24648,N_22823,N_23484);
and U24649 (N_24649,N_22548,N_22641);
and U24650 (N_24650,N_23200,N_22715);
nor U24651 (N_24651,N_22608,N_23209);
nand U24652 (N_24652,N_23206,N_22882);
or U24653 (N_24653,N_23511,N_23061);
xor U24654 (N_24654,N_23067,N_23741);
nor U24655 (N_24655,N_22659,N_23335);
nor U24656 (N_24656,N_22628,N_23560);
xnor U24657 (N_24657,N_23666,N_22593);
or U24658 (N_24658,N_22651,N_23614);
nand U24659 (N_24659,N_23430,N_23516);
nor U24660 (N_24660,N_22880,N_23265);
nand U24661 (N_24661,N_23696,N_22578);
nor U24662 (N_24662,N_23644,N_23200);
nor U24663 (N_24663,N_23379,N_23467);
and U24664 (N_24664,N_22688,N_22945);
and U24665 (N_24665,N_23723,N_22853);
or U24666 (N_24666,N_22719,N_23582);
nand U24667 (N_24667,N_23116,N_23706);
nand U24668 (N_24668,N_23697,N_22614);
nand U24669 (N_24669,N_23268,N_22670);
nand U24670 (N_24670,N_23666,N_22888);
and U24671 (N_24671,N_23159,N_22712);
xor U24672 (N_24672,N_22721,N_22513);
or U24673 (N_24673,N_23102,N_22905);
or U24674 (N_24674,N_22969,N_23048);
xnor U24675 (N_24675,N_23477,N_23090);
nor U24676 (N_24676,N_22706,N_23392);
nor U24677 (N_24677,N_23711,N_23685);
xnor U24678 (N_24678,N_23549,N_22603);
or U24679 (N_24679,N_22743,N_23377);
and U24680 (N_24680,N_23418,N_23472);
nand U24681 (N_24681,N_23282,N_23637);
nor U24682 (N_24682,N_23348,N_23657);
nor U24683 (N_24683,N_23730,N_22707);
xor U24684 (N_24684,N_23137,N_23733);
or U24685 (N_24685,N_23075,N_23289);
xor U24686 (N_24686,N_22503,N_22796);
or U24687 (N_24687,N_23395,N_22930);
or U24688 (N_24688,N_23252,N_23714);
nand U24689 (N_24689,N_23003,N_22999);
nor U24690 (N_24690,N_23648,N_22817);
nand U24691 (N_24691,N_22858,N_23003);
xnor U24692 (N_24692,N_23624,N_23325);
xnor U24693 (N_24693,N_22638,N_23728);
nor U24694 (N_24694,N_22679,N_23742);
or U24695 (N_24695,N_22791,N_23014);
nand U24696 (N_24696,N_22742,N_22888);
nand U24697 (N_24697,N_22612,N_23548);
nand U24698 (N_24698,N_23113,N_23330);
nor U24699 (N_24699,N_23597,N_23052);
or U24700 (N_24700,N_22999,N_23449);
nor U24701 (N_24701,N_23475,N_23527);
and U24702 (N_24702,N_22544,N_23115);
nand U24703 (N_24703,N_23707,N_23251);
or U24704 (N_24704,N_22743,N_22896);
xnor U24705 (N_24705,N_22923,N_22613);
or U24706 (N_24706,N_23735,N_22777);
and U24707 (N_24707,N_23096,N_23690);
or U24708 (N_24708,N_22915,N_22739);
nand U24709 (N_24709,N_23281,N_22704);
and U24710 (N_24710,N_23107,N_22600);
xor U24711 (N_24711,N_23721,N_23610);
nor U24712 (N_24712,N_22516,N_23372);
nand U24713 (N_24713,N_23642,N_22719);
xor U24714 (N_24714,N_23445,N_23478);
xnor U24715 (N_24715,N_23209,N_23538);
xor U24716 (N_24716,N_22765,N_22879);
xor U24717 (N_24717,N_22867,N_23727);
and U24718 (N_24718,N_23233,N_23545);
and U24719 (N_24719,N_23621,N_23300);
or U24720 (N_24720,N_23481,N_22904);
xnor U24721 (N_24721,N_23345,N_23712);
nor U24722 (N_24722,N_22680,N_22600);
or U24723 (N_24723,N_23619,N_23324);
and U24724 (N_24724,N_22846,N_22560);
nand U24725 (N_24725,N_22872,N_22746);
or U24726 (N_24726,N_22531,N_23170);
nand U24727 (N_24727,N_22839,N_23620);
nor U24728 (N_24728,N_22966,N_22739);
xor U24729 (N_24729,N_22755,N_22663);
and U24730 (N_24730,N_23110,N_22877);
nand U24731 (N_24731,N_23196,N_23722);
and U24732 (N_24732,N_22967,N_23698);
or U24733 (N_24733,N_23439,N_23560);
and U24734 (N_24734,N_22714,N_22640);
nor U24735 (N_24735,N_23238,N_23741);
or U24736 (N_24736,N_23361,N_22675);
xor U24737 (N_24737,N_23551,N_23610);
xor U24738 (N_24738,N_22873,N_23088);
or U24739 (N_24739,N_22513,N_23605);
nor U24740 (N_24740,N_22869,N_22701);
xor U24741 (N_24741,N_22793,N_23268);
or U24742 (N_24742,N_23450,N_23317);
xor U24743 (N_24743,N_22748,N_22633);
or U24744 (N_24744,N_22820,N_23480);
or U24745 (N_24745,N_23676,N_22689);
and U24746 (N_24746,N_23025,N_23437);
xnor U24747 (N_24747,N_23380,N_23091);
xor U24748 (N_24748,N_23183,N_23046);
and U24749 (N_24749,N_22820,N_22697);
nand U24750 (N_24750,N_22852,N_22816);
xnor U24751 (N_24751,N_23236,N_23362);
or U24752 (N_24752,N_23123,N_22862);
and U24753 (N_24753,N_22630,N_23616);
xnor U24754 (N_24754,N_23380,N_22701);
xor U24755 (N_24755,N_23734,N_22652);
nand U24756 (N_24756,N_23340,N_22590);
xnor U24757 (N_24757,N_23460,N_22999);
nand U24758 (N_24758,N_23275,N_22860);
xor U24759 (N_24759,N_23011,N_23260);
nand U24760 (N_24760,N_23414,N_22541);
nor U24761 (N_24761,N_22793,N_23400);
and U24762 (N_24762,N_23385,N_23354);
and U24763 (N_24763,N_23629,N_23121);
nor U24764 (N_24764,N_23158,N_23166);
and U24765 (N_24765,N_22844,N_23340);
nand U24766 (N_24766,N_23515,N_23477);
xnor U24767 (N_24767,N_23747,N_22788);
and U24768 (N_24768,N_22650,N_23595);
or U24769 (N_24769,N_23480,N_23528);
nand U24770 (N_24770,N_23159,N_22914);
nand U24771 (N_24771,N_22542,N_22685);
nand U24772 (N_24772,N_23646,N_22736);
and U24773 (N_24773,N_23668,N_22747);
and U24774 (N_24774,N_23038,N_23456);
and U24775 (N_24775,N_22671,N_23010);
nand U24776 (N_24776,N_22792,N_23191);
xnor U24777 (N_24777,N_22679,N_22802);
or U24778 (N_24778,N_22873,N_23289);
nor U24779 (N_24779,N_22521,N_22688);
xor U24780 (N_24780,N_23274,N_23641);
or U24781 (N_24781,N_23631,N_23172);
nor U24782 (N_24782,N_22726,N_22622);
nand U24783 (N_24783,N_23450,N_22638);
nor U24784 (N_24784,N_23147,N_22614);
and U24785 (N_24785,N_23724,N_22645);
and U24786 (N_24786,N_23270,N_23075);
nand U24787 (N_24787,N_22979,N_22720);
and U24788 (N_24788,N_23598,N_23335);
or U24789 (N_24789,N_22933,N_22883);
nand U24790 (N_24790,N_22579,N_23727);
xor U24791 (N_24791,N_23631,N_23015);
and U24792 (N_24792,N_23131,N_22709);
and U24793 (N_24793,N_23495,N_23338);
xnor U24794 (N_24794,N_22936,N_23296);
nor U24795 (N_24795,N_22912,N_23634);
and U24796 (N_24796,N_23289,N_23611);
nor U24797 (N_24797,N_23692,N_22820);
xnor U24798 (N_24798,N_22876,N_23476);
and U24799 (N_24799,N_23608,N_22551);
xor U24800 (N_24800,N_23389,N_22881);
nor U24801 (N_24801,N_23194,N_23570);
xor U24802 (N_24802,N_23338,N_23387);
nor U24803 (N_24803,N_23651,N_23068);
nand U24804 (N_24804,N_23370,N_23407);
and U24805 (N_24805,N_22508,N_22595);
nand U24806 (N_24806,N_23079,N_23130);
nand U24807 (N_24807,N_23096,N_23578);
or U24808 (N_24808,N_23332,N_22618);
nor U24809 (N_24809,N_22883,N_23178);
or U24810 (N_24810,N_23684,N_22837);
nor U24811 (N_24811,N_22824,N_23709);
and U24812 (N_24812,N_23486,N_22779);
xnor U24813 (N_24813,N_23171,N_23053);
nand U24814 (N_24814,N_23052,N_22932);
or U24815 (N_24815,N_23491,N_23588);
nand U24816 (N_24816,N_22589,N_23267);
nand U24817 (N_24817,N_22727,N_23136);
and U24818 (N_24818,N_23728,N_23333);
nand U24819 (N_24819,N_23601,N_23528);
or U24820 (N_24820,N_22752,N_22916);
or U24821 (N_24821,N_23349,N_23137);
xor U24822 (N_24822,N_23433,N_23048);
nand U24823 (N_24823,N_23097,N_23037);
nor U24824 (N_24824,N_23057,N_22972);
nor U24825 (N_24825,N_23061,N_23137);
or U24826 (N_24826,N_22739,N_23376);
and U24827 (N_24827,N_23373,N_23159);
nor U24828 (N_24828,N_23689,N_22804);
xor U24829 (N_24829,N_23098,N_22951);
xnor U24830 (N_24830,N_23525,N_23615);
xor U24831 (N_24831,N_22999,N_23576);
nor U24832 (N_24832,N_23361,N_22856);
and U24833 (N_24833,N_22893,N_22802);
or U24834 (N_24834,N_23680,N_23730);
nand U24835 (N_24835,N_22722,N_23571);
and U24836 (N_24836,N_23105,N_22878);
nand U24837 (N_24837,N_23481,N_23721);
xnor U24838 (N_24838,N_23520,N_23243);
and U24839 (N_24839,N_22500,N_22820);
and U24840 (N_24840,N_23027,N_22877);
xor U24841 (N_24841,N_23449,N_22949);
nand U24842 (N_24842,N_23105,N_22654);
nor U24843 (N_24843,N_23034,N_23311);
and U24844 (N_24844,N_23004,N_23366);
xnor U24845 (N_24845,N_23618,N_23016);
or U24846 (N_24846,N_23141,N_23334);
or U24847 (N_24847,N_23395,N_22873);
nand U24848 (N_24848,N_22750,N_23523);
xor U24849 (N_24849,N_22986,N_23320);
xnor U24850 (N_24850,N_22809,N_23006);
nor U24851 (N_24851,N_22796,N_23010);
xor U24852 (N_24852,N_23500,N_22766);
xnor U24853 (N_24853,N_23549,N_22985);
nor U24854 (N_24854,N_23430,N_23299);
nor U24855 (N_24855,N_23176,N_22894);
and U24856 (N_24856,N_22908,N_23528);
nand U24857 (N_24857,N_23193,N_22724);
nand U24858 (N_24858,N_23297,N_23670);
nand U24859 (N_24859,N_22993,N_22773);
and U24860 (N_24860,N_23385,N_23198);
or U24861 (N_24861,N_23208,N_23249);
nor U24862 (N_24862,N_23114,N_23515);
nand U24863 (N_24863,N_22841,N_22776);
xnor U24864 (N_24864,N_23234,N_22506);
nand U24865 (N_24865,N_23072,N_23661);
and U24866 (N_24866,N_23623,N_23424);
nor U24867 (N_24867,N_22717,N_22760);
and U24868 (N_24868,N_22556,N_23581);
nand U24869 (N_24869,N_23364,N_22826);
xnor U24870 (N_24870,N_23374,N_23419);
xor U24871 (N_24871,N_22687,N_23594);
and U24872 (N_24872,N_23558,N_23540);
or U24873 (N_24873,N_23387,N_23139);
or U24874 (N_24874,N_23258,N_22630);
xor U24875 (N_24875,N_23011,N_23497);
nor U24876 (N_24876,N_22657,N_23563);
nor U24877 (N_24877,N_22597,N_22658);
and U24878 (N_24878,N_23525,N_23718);
nor U24879 (N_24879,N_23247,N_22869);
and U24880 (N_24880,N_23539,N_23645);
xor U24881 (N_24881,N_23651,N_23733);
and U24882 (N_24882,N_22731,N_23310);
nor U24883 (N_24883,N_22613,N_22981);
xor U24884 (N_24884,N_23229,N_23096);
and U24885 (N_24885,N_23454,N_23409);
and U24886 (N_24886,N_23722,N_22586);
and U24887 (N_24887,N_22742,N_22741);
and U24888 (N_24888,N_23514,N_23551);
nand U24889 (N_24889,N_23657,N_23118);
or U24890 (N_24890,N_23488,N_23000);
nor U24891 (N_24891,N_23006,N_23356);
and U24892 (N_24892,N_23013,N_23247);
xnor U24893 (N_24893,N_22526,N_23023);
nand U24894 (N_24894,N_22561,N_22533);
and U24895 (N_24895,N_22967,N_23379);
nand U24896 (N_24896,N_22916,N_22547);
and U24897 (N_24897,N_22586,N_23105);
xnor U24898 (N_24898,N_23115,N_23549);
nor U24899 (N_24899,N_22773,N_23113);
nand U24900 (N_24900,N_23271,N_23360);
xnor U24901 (N_24901,N_22547,N_22819);
nor U24902 (N_24902,N_23140,N_22999);
or U24903 (N_24903,N_23463,N_22735);
nand U24904 (N_24904,N_23592,N_22597);
xnor U24905 (N_24905,N_23100,N_23247);
or U24906 (N_24906,N_22622,N_23123);
and U24907 (N_24907,N_22779,N_22746);
nand U24908 (N_24908,N_22850,N_22767);
and U24909 (N_24909,N_23361,N_22720);
and U24910 (N_24910,N_22823,N_23618);
nor U24911 (N_24911,N_23589,N_23375);
nand U24912 (N_24912,N_23385,N_22610);
xor U24913 (N_24913,N_22530,N_23106);
nor U24914 (N_24914,N_23562,N_23185);
or U24915 (N_24915,N_23111,N_23520);
or U24916 (N_24916,N_22794,N_22911);
xor U24917 (N_24917,N_22825,N_23012);
nor U24918 (N_24918,N_23073,N_22617);
nor U24919 (N_24919,N_23021,N_23269);
nor U24920 (N_24920,N_23323,N_23689);
and U24921 (N_24921,N_23129,N_23590);
or U24922 (N_24922,N_23030,N_23676);
and U24923 (N_24923,N_23150,N_23529);
nor U24924 (N_24924,N_23402,N_23447);
and U24925 (N_24925,N_23672,N_23744);
or U24926 (N_24926,N_23389,N_23498);
nor U24927 (N_24927,N_23266,N_23507);
nand U24928 (N_24928,N_23580,N_23066);
xor U24929 (N_24929,N_23177,N_23019);
nor U24930 (N_24930,N_23088,N_23747);
or U24931 (N_24931,N_23442,N_23454);
xor U24932 (N_24932,N_22949,N_22615);
xor U24933 (N_24933,N_22899,N_22701);
nor U24934 (N_24934,N_23308,N_22612);
and U24935 (N_24935,N_22946,N_22806);
xnor U24936 (N_24936,N_22895,N_23629);
xnor U24937 (N_24937,N_23190,N_22841);
nand U24938 (N_24938,N_23139,N_23723);
nor U24939 (N_24939,N_22848,N_22849);
nand U24940 (N_24940,N_23662,N_23509);
nor U24941 (N_24941,N_23245,N_23470);
and U24942 (N_24942,N_23680,N_23354);
or U24943 (N_24943,N_23553,N_22568);
and U24944 (N_24944,N_23357,N_23450);
and U24945 (N_24945,N_23464,N_23265);
xnor U24946 (N_24946,N_22873,N_22624);
xor U24947 (N_24947,N_23256,N_22640);
nand U24948 (N_24948,N_23673,N_23378);
or U24949 (N_24949,N_22904,N_22882);
nor U24950 (N_24950,N_22527,N_23366);
xnor U24951 (N_24951,N_22896,N_23068);
and U24952 (N_24952,N_22621,N_22742);
nor U24953 (N_24953,N_23005,N_22922);
nor U24954 (N_24954,N_22902,N_23566);
nor U24955 (N_24955,N_23490,N_23359);
nor U24956 (N_24956,N_22928,N_23676);
or U24957 (N_24957,N_23513,N_23205);
nand U24958 (N_24958,N_23504,N_22800);
nor U24959 (N_24959,N_23556,N_23302);
or U24960 (N_24960,N_23184,N_23089);
and U24961 (N_24961,N_23097,N_23266);
xor U24962 (N_24962,N_22858,N_23713);
or U24963 (N_24963,N_22748,N_22950);
xor U24964 (N_24964,N_22597,N_23062);
or U24965 (N_24965,N_22888,N_22678);
and U24966 (N_24966,N_22713,N_22855);
nor U24967 (N_24967,N_22801,N_22520);
nor U24968 (N_24968,N_22531,N_22795);
xnor U24969 (N_24969,N_23046,N_22758);
xor U24970 (N_24970,N_23346,N_22704);
nor U24971 (N_24971,N_23232,N_22963);
nand U24972 (N_24972,N_23449,N_23038);
nand U24973 (N_24973,N_22790,N_23724);
xor U24974 (N_24974,N_22676,N_22808);
and U24975 (N_24975,N_23628,N_22890);
xor U24976 (N_24976,N_23170,N_23556);
nand U24977 (N_24977,N_22816,N_22917);
xnor U24978 (N_24978,N_23549,N_23074);
and U24979 (N_24979,N_23505,N_23006);
and U24980 (N_24980,N_23521,N_22774);
or U24981 (N_24981,N_22966,N_23683);
nor U24982 (N_24982,N_23702,N_22801);
nor U24983 (N_24983,N_22838,N_23471);
xor U24984 (N_24984,N_23510,N_23115);
or U24985 (N_24985,N_23301,N_22986);
nand U24986 (N_24986,N_23579,N_23363);
or U24987 (N_24987,N_23416,N_22908);
nand U24988 (N_24988,N_22739,N_22921);
nand U24989 (N_24989,N_23359,N_23524);
xor U24990 (N_24990,N_22614,N_23319);
nor U24991 (N_24991,N_22537,N_23269);
nor U24992 (N_24992,N_23150,N_22735);
nand U24993 (N_24993,N_23497,N_22659);
and U24994 (N_24994,N_23457,N_23395);
xor U24995 (N_24995,N_22690,N_22963);
nor U24996 (N_24996,N_23421,N_23261);
or U24997 (N_24997,N_22715,N_23257);
nand U24998 (N_24998,N_23646,N_23538);
and U24999 (N_24999,N_23485,N_22688);
xor UO_0 (O_0,N_24110,N_24924);
xor UO_1 (O_1,N_24186,N_24668);
and UO_2 (O_2,N_23775,N_24039);
nor UO_3 (O_3,N_24538,N_24262);
and UO_4 (O_4,N_24999,N_23793);
nand UO_5 (O_5,N_24631,N_24147);
nor UO_6 (O_6,N_24275,N_24265);
xnor UO_7 (O_7,N_24777,N_24701);
or UO_8 (O_8,N_24634,N_24439);
nand UO_9 (O_9,N_24004,N_24018);
or UO_10 (O_10,N_23870,N_24414);
nor UO_11 (O_11,N_23894,N_24406);
nor UO_12 (O_12,N_24712,N_24674);
or UO_13 (O_13,N_24301,N_24381);
xor UO_14 (O_14,N_24149,N_23835);
nor UO_15 (O_15,N_24917,N_24325);
xnor UO_16 (O_16,N_24798,N_23751);
xor UO_17 (O_17,N_23909,N_24692);
and UO_18 (O_18,N_24821,N_24020);
nand UO_19 (O_19,N_23821,N_24288);
xnor UO_20 (O_20,N_24533,N_24923);
or UO_21 (O_21,N_23954,N_24331);
nor UO_22 (O_22,N_23903,N_23759);
nand UO_23 (O_23,N_24160,N_24482);
nand UO_24 (O_24,N_24600,N_24783);
and UO_25 (O_25,N_24006,N_24138);
xor UO_26 (O_26,N_23784,N_24091);
or UO_27 (O_27,N_24475,N_24390);
xnor UO_28 (O_28,N_24738,N_24530);
or UO_29 (O_29,N_24983,N_24977);
nor UO_30 (O_30,N_23998,N_24435);
or UO_31 (O_31,N_24889,N_23970);
or UO_32 (O_32,N_24108,N_24744);
nand UO_33 (O_33,N_24412,N_24569);
nand UO_34 (O_34,N_24845,N_24419);
or UO_35 (O_35,N_24164,N_24469);
nand UO_36 (O_36,N_24661,N_24895);
nand UO_37 (O_37,N_23808,N_24825);
and UO_38 (O_38,N_24461,N_24894);
nand UO_39 (O_39,N_24540,N_24935);
or UO_40 (O_40,N_24552,N_24974);
xnor UO_41 (O_41,N_24396,N_24945);
and UO_42 (O_42,N_24684,N_24713);
nor UO_43 (O_43,N_24460,N_23755);
xor UO_44 (O_44,N_24636,N_24949);
nor UO_45 (O_45,N_24590,N_24840);
nand UO_46 (O_46,N_24034,N_24127);
or UO_47 (O_47,N_24446,N_23857);
and UO_48 (O_48,N_24306,N_24978);
or UO_49 (O_49,N_24191,N_24902);
xnor UO_50 (O_50,N_24335,N_24979);
or UO_51 (O_51,N_24341,N_24660);
nand UO_52 (O_52,N_24922,N_23763);
or UO_53 (O_53,N_24302,N_24354);
nand UO_54 (O_54,N_24383,N_24679);
and UO_55 (O_55,N_24471,N_23845);
xnor UO_56 (O_56,N_24221,N_24623);
nand UO_57 (O_57,N_24440,N_24157);
or UO_58 (O_58,N_24918,N_24070);
nor UO_59 (O_59,N_24520,N_24096);
nor UO_60 (O_60,N_24824,N_24787);
xor UO_61 (O_61,N_24338,N_24271);
nor UO_62 (O_62,N_23764,N_24180);
or UO_63 (O_63,N_23796,N_24179);
and UO_64 (O_64,N_24462,N_24937);
nand UO_65 (O_65,N_24342,N_24077);
or UO_66 (O_66,N_24316,N_24357);
or UO_67 (O_67,N_24167,N_24795);
nor UO_68 (O_68,N_24653,N_24364);
xnor UO_69 (O_69,N_23760,N_23914);
and UO_70 (O_70,N_24133,N_24496);
nor UO_71 (O_71,N_23789,N_24458);
nand UO_72 (O_72,N_24087,N_23818);
or UO_73 (O_73,N_24719,N_24499);
nor UO_74 (O_74,N_23897,N_24963);
or UO_75 (O_75,N_24046,N_24747);
xor UO_76 (O_76,N_23819,N_24075);
xnor UO_77 (O_77,N_24410,N_24346);
and UO_78 (O_78,N_23875,N_24907);
xnor UO_79 (O_79,N_24896,N_24916);
nor UO_80 (O_80,N_24480,N_24742);
nand UO_81 (O_81,N_24259,N_24545);
nor UO_82 (O_82,N_24099,N_24062);
nand UO_83 (O_83,N_24076,N_24151);
and UO_84 (O_84,N_23902,N_23790);
xor UO_85 (O_85,N_23913,N_24314);
nor UO_86 (O_86,N_23887,N_23920);
xnor UO_87 (O_87,N_24094,N_24558);
nand UO_88 (O_88,N_24064,N_24365);
nor UO_89 (O_89,N_24641,N_23817);
nand UO_90 (O_90,N_24502,N_24700);
nand UO_91 (O_91,N_23883,N_24154);
nor UO_92 (O_92,N_24348,N_24142);
nor UO_93 (O_93,N_24721,N_24337);
or UO_94 (O_94,N_23872,N_24685);
or UO_95 (O_95,N_24539,N_23921);
nand UO_96 (O_96,N_24613,N_24589);
nor UO_97 (O_97,N_24955,N_24417);
and UO_98 (O_98,N_24019,N_24557);
and UO_99 (O_99,N_24898,N_24696);
and UO_100 (O_100,N_24961,N_24804);
or UO_101 (O_101,N_23997,N_24788);
or UO_102 (O_102,N_24195,N_23839);
xor UO_103 (O_103,N_24194,N_23867);
nand UO_104 (O_104,N_24115,N_24843);
or UO_105 (O_105,N_24403,N_24758);
nand UO_106 (O_106,N_24678,N_24047);
nor UO_107 (O_107,N_24782,N_24362);
xor UO_108 (O_108,N_24145,N_23892);
xnor UO_109 (O_109,N_24465,N_24415);
and UO_110 (O_110,N_24053,N_24352);
or UO_111 (O_111,N_24165,N_23795);
nand UO_112 (O_112,N_23978,N_23855);
or UO_113 (O_113,N_23853,N_24866);
or UO_114 (O_114,N_23767,N_24009);
xor UO_115 (O_115,N_23823,N_24715);
nand UO_116 (O_116,N_24809,N_24510);
nand UO_117 (O_117,N_24617,N_24134);
xor UO_118 (O_118,N_24375,N_24002);
or UO_119 (O_119,N_24212,N_24041);
nor UO_120 (O_120,N_23915,N_24305);
xor UO_121 (O_121,N_24888,N_24449);
and UO_122 (O_122,N_24610,N_24242);
nor UO_123 (O_123,N_23959,N_24547);
nand UO_124 (O_124,N_23937,N_23791);
nor UO_125 (O_125,N_24579,N_24570);
or UO_126 (O_126,N_23905,N_24878);
and UO_127 (O_127,N_24119,N_23918);
nor UO_128 (O_128,N_24125,N_23911);
or UO_129 (O_129,N_24571,N_23856);
nand UO_130 (O_130,N_24445,N_24230);
xor UO_131 (O_131,N_24083,N_24694);
xnor UO_132 (O_132,N_24683,N_24799);
or UO_133 (O_133,N_24765,N_24677);
or UO_134 (O_134,N_23936,N_24444);
and UO_135 (O_135,N_24132,N_24013);
xnor UO_136 (O_136,N_24090,N_24920);
and UO_137 (O_137,N_24264,N_24771);
xnor UO_138 (O_138,N_24773,N_24048);
or UO_139 (O_139,N_24232,N_24508);
or UO_140 (O_140,N_24386,N_24527);
nand UO_141 (O_141,N_24481,N_23981);
xor UO_142 (O_142,N_23991,N_24231);
nand UO_143 (O_143,N_23885,N_23929);
or UO_144 (O_144,N_23972,N_24268);
xor UO_145 (O_145,N_24318,N_24521);
nor UO_146 (O_146,N_24309,N_24546);
xnor UO_147 (O_147,N_24792,N_24356);
and UO_148 (O_148,N_23977,N_24656);
nand UO_149 (O_149,N_24483,N_24594);
xnor UO_150 (O_150,N_24913,N_24796);
xnor UO_151 (O_151,N_24402,N_24463);
and UO_152 (O_152,N_24189,N_24226);
and UO_153 (O_153,N_24060,N_23891);
or UO_154 (O_154,N_24373,N_23908);
nand UO_155 (O_155,N_24903,N_24645);
xnor UO_156 (O_156,N_24856,N_23899);
and UO_157 (O_157,N_24926,N_24328);
nand UO_158 (O_158,N_24612,N_24411);
nor UO_159 (O_159,N_24644,N_24720);
and UO_160 (O_160,N_24181,N_24056);
nor UO_161 (O_161,N_24812,N_24274);
or UO_162 (O_162,N_23943,N_24097);
xor UO_163 (O_163,N_23901,N_24453);
nor UO_164 (O_164,N_24037,N_24972);
nand UO_165 (O_165,N_24861,N_24584);
nand UO_166 (O_166,N_24515,N_24437);
nor UO_167 (O_167,N_24892,N_24639);
nor UO_168 (O_168,N_24389,N_24772);
xor UO_169 (O_169,N_24178,N_24688);
nor UO_170 (O_170,N_24556,N_23838);
or UO_171 (O_171,N_24217,N_24849);
nor UO_172 (O_172,N_23946,N_24586);
and UO_173 (O_173,N_24256,N_24135);
and UO_174 (O_174,N_24248,N_24956);
xor UO_175 (O_175,N_24855,N_24535);
nor UO_176 (O_176,N_24879,N_24332);
or UO_177 (O_177,N_24223,N_24672);
xnor UO_178 (O_178,N_24627,N_24126);
and UO_179 (O_179,N_24371,N_24954);
nor UO_180 (O_180,N_24253,N_23849);
or UO_181 (O_181,N_24263,N_24366);
and UO_182 (O_182,N_23761,N_24830);
nand UO_183 (O_183,N_24958,N_23974);
xnor UO_184 (O_184,N_24632,N_24624);
or UO_185 (O_185,N_24575,N_24304);
or UO_186 (O_186,N_24750,N_24313);
xor UO_187 (O_187,N_23962,N_24484);
nor UO_188 (O_188,N_24485,N_24211);
nor UO_189 (O_189,N_24884,N_23843);
nand UO_190 (O_190,N_23851,N_24850);
and UO_191 (O_191,N_23890,N_23996);
xor UO_192 (O_192,N_24355,N_24940);
nand UO_193 (O_193,N_23985,N_24741);
and UO_194 (O_194,N_24580,N_24380);
nand UO_195 (O_195,N_23820,N_24838);
nand UO_196 (O_196,N_24786,N_24582);
nand UO_197 (O_197,N_24123,N_24592);
xnor UO_198 (O_198,N_24505,N_24139);
or UO_199 (O_199,N_24454,N_23932);
nor UO_200 (O_200,N_24511,N_24358);
and UO_201 (O_201,N_23874,N_23832);
and UO_202 (O_202,N_24984,N_24122);
or UO_203 (O_203,N_23935,N_24239);
xnor UO_204 (O_204,N_23800,N_24307);
nor UO_205 (O_205,N_24057,N_24597);
xor UO_206 (O_206,N_24835,N_24379);
or UO_207 (O_207,N_24395,N_24052);
and UO_208 (O_208,N_24012,N_24737);
or UO_209 (O_209,N_24686,N_24517);
or UO_210 (O_210,N_24093,N_23948);
xnor UO_211 (O_211,N_24904,N_23917);
nand UO_212 (O_212,N_23881,N_24982);
or UO_213 (O_213,N_23830,N_24368);
and UO_214 (O_214,N_23924,N_24144);
or UO_215 (O_215,N_24942,N_24962);
nor UO_216 (O_216,N_24699,N_24299);
or UO_217 (O_217,N_23926,N_24489);
and UO_218 (O_218,N_24303,N_23848);
xnor UO_219 (O_219,N_23827,N_24203);
nor UO_220 (O_220,N_24109,N_24294);
or UO_221 (O_221,N_24209,N_24021);
xor UO_222 (O_222,N_24664,N_24997);
and UO_223 (O_223,N_24030,N_23864);
or UO_224 (O_224,N_24168,N_24529);
and UO_225 (O_225,N_24662,N_24103);
nand UO_226 (O_226,N_24543,N_24351);
xnor UO_227 (O_227,N_24970,N_24257);
nand UO_228 (O_228,N_24646,N_23907);
and UO_229 (O_229,N_24757,N_24731);
and UO_230 (O_230,N_23834,N_24234);
and UO_231 (O_231,N_24184,N_24359);
nor UO_232 (O_232,N_24811,N_24973);
or UO_233 (O_233,N_23980,N_24576);
xor UO_234 (O_234,N_24710,N_24273);
or UO_235 (O_235,N_23785,N_24442);
and UO_236 (O_236,N_24790,N_24588);
or UO_237 (O_237,N_23801,N_23994);
nand UO_238 (O_238,N_24260,N_24560);
xor UO_239 (O_239,N_24908,N_24643);
nor UO_240 (O_240,N_24599,N_24620);
and UO_241 (O_241,N_24562,N_24844);
and UO_242 (O_242,N_24312,N_24397);
and UO_243 (O_243,N_24238,N_24503);
or UO_244 (O_244,N_24280,N_24289);
and UO_245 (O_245,N_24279,N_24969);
and UO_246 (O_246,N_24689,N_23960);
nand UO_247 (O_247,N_24652,N_24714);
nand UO_248 (O_248,N_24655,N_24549);
nand UO_249 (O_249,N_23797,N_24881);
xnor UO_250 (O_250,N_24113,N_24343);
or UO_251 (O_251,N_24407,N_24794);
or UO_252 (O_252,N_24010,N_24638);
or UO_253 (O_253,N_24198,N_24286);
and UO_254 (O_254,N_24367,N_24960);
xnor UO_255 (O_255,N_24036,N_23773);
nand UO_256 (O_256,N_24659,N_23792);
and UO_257 (O_257,N_24675,N_24893);
and UO_258 (O_258,N_24567,N_24088);
and UO_259 (O_259,N_24630,N_24427);
nor UO_260 (O_260,N_24282,N_24761);
nand UO_261 (O_261,N_24801,N_24158);
nor UO_262 (O_262,N_24376,N_24501);
or UO_263 (O_263,N_24345,N_24150);
or UO_264 (O_264,N_23869,N_24785);
nand UO_265 (O_265,N_24272,N_24323);
and UO_266 (O_266,N_24038,N_23871);
and UO_267 (O_267,N_23886,N_24528);
and UO_268 (O_268,N_24063,N_24491);
or UO_269 (O_269,N_23884,N_24625);
xnor UO_270 (O_270,N_24350,N_24073);
nor UO_271 (O_271,N_23811,N_24531);
xor UO_272 (O_272,N_24320,N_24116);
and UO_273 (O_273,N_24105,N_24258);
xnor UO_274 (O_274,N_24155,N_24204);
nor UO_275 (O_275,N_24162,N_23882);
and UO_276 (O_276,N_23840,N_24704);
xor UO_277 (O_277,N_24494,N_24957);
and UO_278 (O_278,N_24423,N_24474);
and UO_279 (O_279,N_23778,N_23923);
nor UO_280 (O_280,N_24754,N_24296);
nand UO_281 (O_281,N_24936,N_24055);
nand UO_282 (O_282,N_23966,N_23799);
and UO_283 (O_283,N_24219,N_24981);
or UO_284 (O_284,N_24793,N_24572);
nand UO_285 (O_285,N_24770,N_23950);
nor UO_286 (O_286,N_24618,N_24953);
nand UO_287 (O_287,N_24875,N_24544);
xnor UO_288 (O_288,N_23878,N_24829);
nand UO_289 (O_289,N_24550,N_24387);
nand UO_290 (O_290,N_23963,N_24431);
or UO_291 (O_291,N_24990,N_24665);
nor UO_292 (O_292,N_24255,N_24723);
nand UO_293 (O_293,N_23990,N_23782);
or UO_294 (O_294,N_24869,N_24947);
and UO_295 (O_295,N_24868,N_24749);
xnor UO_296 (O_296,N_24237,N_23916);
xor UO_297 (O_297,N_24228,N_24774);
and UO_298 (O_298,N_23988,N_24479);
and UO_299 (O_299,N_24732,N_24224);
or UO_300 (O_300,N_24581,N_24111);
and UO_301 (O_301,N_24506,N_24360);
and UO_302 (O_302,N_24814,N_24728);
or UO_303 (O_303,N_24089,N_24016);
and UO_304 (O_304,N_24416,N_24778);
nand UO_305 (O_305,N_24727,N_24252);
or UO_306 (O_306,N_23931,N_23898);
or UO_307 (O_307,N_24565,N_24218);
and UO_308 (O_308,N_23951,N_24946);
nand UO_309 (O_309,N_24240,N_24227);
or UO_310 (O_310,N_24175,N_24404);
or UO_311 (O_311,N_24196,N_24022);
xor UO_312 (O_312,N_24400,N_24270);
nand UO_313 (O_313,N_23927,N_24890);
and UO_314 (O_314,N_24608,N_24975);
xor UO_315 (O_315,N_24349,N_24595);
and UO_316 (O_316,N_23975,N_24472);
xor UO_317 (O_317,N_24910,N_24583);
or UO_318 (O_318,N_24803,N_24043);
xnor UO_319 (O_319,N_24311,N_24065);
nand UO_320 (O_320,N_24912,N_24059);
xor UO_321 (O_321,N_24611,N_24734);
xnor UO_322 (O_322,N_24098,N_24229);
nand UO_323 (O_323,N_24326,N_24032);
and UO_324 (O_324,N_24836,N_24278);
xnor UO_325 (O_325,N_24478,N_24806);
nand UO_326 (O_326,N_24779,N_24436);
nor UO_327 (O_327,N_23896,N_24837);
nand UO_328 (O_328,N_24300,N_24781);
xor UO_329 (O_329,N_24522,N_24339);
nand UO_330 (O_330,N_23982,N_24353);
and UO_331 (O_331,N_24319,N_24554);
nor UO_332 (O_332,N_24045,N_24939);
and UO_333 (O_333,N_24933,N_23910);
nand UO_334 (O_334,N_24764,N_24054);
and UO_335 (O_335,N_23812,N_23912);
nand UO_336 (O_336,N_23945,N_24998);
xnor UO_337 (O_337,N_24553,N_24249);
and UO_338 (O_338,N_24051,N_24438);
and UO_339 (O_339,N_24197,N_24745);
and UO_340 (O_340,N_23806,N_24159);
nor UO_341 (O_341,N_24828,N_24370);
nor UO_342 (O_342,N_23802,N_24329);
nand UO_343 (O_343,N_24810,N_24965);
and UO_344 (O_344,N_24340,N_23803);
and UO_345 (O_345,N_24996,N_23815);
and UO_346 (O_346,N_24932,N_24598);
xor UO_347 (O_347,N_23758,N_24883);
and UO_348 (O_348,N_23774,N_24459);
or UO_349 (O_349,N_24222,N_24388);
and UO_350 (O_350,N_24860,N_24267);
and UO_351 (O_351,N_24657,N_24137);
nor UO_352 (O_352,N_24372,N_23769);
nand UO_353 (O_353,N_24163,N_23889);
nand UO_354 (O_354,N_24452,N_24784);
or UO_355 (O_355,N_24061,N_23942);
and UO_356 (O_356,N_24780,N_24681);
or UO_357 (O_357,N_23964,N_24992);
and UO_358 (O_358,N_24711,N_24216);
xnor UO_359 (O_359,N_24080,N_24591);
nand UO_360 (O_360,N_24891,N_24141);
xor UO_361 (O_361,N_24493,N_24733);
and UO_362 (O_362,N_24315,N_23983);
nand UO_363 (O_363,N_24466,N_24951);
xnor UO_364 (O_364,N_24193,N_24470);
xnor UO_365 (O_365,N_24152,N_24867);
or UO_366 (O_366,N_24433,N_24832);
or UO_367 (O_367,N_24759,N_24601);
nand UO_368 (O_368,N_23859,N_24769);
or UO_369 (O_369,N_24669,N_23862);
nor UO_370 (O_370,N_24432,N_24200);
or UO_371 (O_371,N_24287,N_24626);
nor UO_372 (O_372,N_23955,N_24284);
xor UO_373 (O_373,N_23854,N_24106);
nor UO_374 (O_374,N_23939,N_24391);
and UO_375 (O_375,N_24680,N_24001);
or UO_376 (O_376,N_24900,N_24899);
or UO_377 (O_377,N_24512,N_24457);
xor UO_378 (O_378,N_24143,N_24188);
or UO_379 (O_379,N_24995,N_23961);
nor UO_380 (O_380,N_24207,N_23770);
and UO_381 (O_381,N_24994,N_24541);
xor UO_382 (O_382,N_24691,N_24698);
or UO_383 (O_383,N_23766,N_24606);
and UO_384 (O_384,N_24490,N_24235);
nor UO_385 (O_385,N_24763,N_23953);
and UO_386 (O_386,N_24455,N_23949);
nor UO_387 (O_387,N_24295,N_24676);
nand UO_388 (O_388,N_23968,N_24808);
nand UO_389 (O_389,N_23944,N_23816);
or UO_390 (O_390,N_24082,N_24418);
and UO_391 (O_391,N_24000,N_24324);
nand UO_392 (O_392,N_24044,N_24863);
xnor UO_393 (O_393,N_24693,N_24833);
xor UO_394 (O_394,N_24602,N_24716);
or UO_395 (O_395,N_24277,N_24938);
xnor UO_396 (O_396,N_24649,N_24635);
xnor UO_397 (O_397,N_23750,N_24604);
or UO_398 (O_398,N_23992,N_23873);
or UO_399 (O_399,N_23860,N_24950);
and UO_400 (O_400,N_24633,N_24118);
or UO_401 (O_401,N_24872,N_24344);
or UO_402 (O_402,N_24492,N_24847);
nand UO_403 (O_403,N_23858,N_24585);
xor UO_404 (O_404,N_23925,N_24401);
and UO_405 (O_405,N_24746,N_24202);
or UO_406 (O_406,N_24011,N_24842);
nor UO_407 (O_407,N_24690,N_24619);
xnor UO_408 (O_408,N_24399,N_24815);
xor UO_409 (O_409,N_24532,N_24031);
xor UO_410 (O_410,N_24526,N_24752);
or UO_411 (O_411,N_24298,N_24124);
nor UO_412 (O_412,N_24425,N_24254);
nor UO_413 (O_413,N_24524,N_23930);
nand UO_414 (O_414,N_24495,N_23781);
xor UO_415 (O_415,N_24851,N_24853);
nand UO_416 (O_416,N_24559,N_24839);
nand UO_417 (O_417,N_23976,N_24504);
nand UO_418 (O_418,N_24443,N_23779);
nor UO_419 (O_419,N_24991,N_23756);
nor UO_420 (O_420,N_24171,N_24886);
or UO_421 (O_421,N_24536,N_23846);
and UO_422 (O_422,N_23877,N_24233);
and UO_423 (O_423,N_24966,N_24276);
and UO_424 (O_424,N_23831,N_24921);
nand UO_425 (O_425,N_24753,N_24285);
xor UO_426 (O_426,N_24384,N_24885);
xor UO_427 (O_427,N_24967,N_24291);
xor UO_428 (O_428,N_24857,N_24434);
and UO_429 (O_429,N_24548,N_24568);
and UO_430 (O_430,N_23833,N_24642);
nand UO_431 (O_431,N_24813,N_24729);
nor UO_432 (O_432,N_24682,N_24650);
xor UO_433 (O_433,N_24247,N_24183);
nor UO_434 (O_434,N_24876,N_24897);
nor UO_435 (O_435,N_24614,N_23777);
xor UO_436 (O_436,N_24333,N_24709);
or UO_437 (O_437,N_24250,N_24555);
and UO_438 (O_438,N_24007,N_24708);
nor UO_439 (O_439,N_24042,N_23984);
nand UO_440 (O_440,N_24725,N_24605);
xnor UO_441 (O_441,N_24948,N_24706);
nor UO_442 (O_442,N_24500,N_24776);
nor UO_443 (O_443,N_24336,N_24578);
xnor UO_444 (O_444,N_24648,N_24718);
and UO_445 (O_445,N_23866,N_24015);
nor UO_446 (O_446,N_24663,N_24448);
nor UO_447 (O_447,N_24170,N_24382);
nand UO_448 (O_448,N_24671,N_24673);
xor UO_449 (O_449,N_24441,N_24146);
nand UO_450 (O_450,N_23919,N_24129);
nor UO_451 (O_451,N_23842,N_24182);
nor UO_452 (O_452,N_24166,N_24943);
nand UO_453 (O_453,N_24577,N_24827);
nor UO_454 (O_454,N_24596,N_24206);
and UO_455 (O_455,N_24498,N_23969);
or UO_456 (O_456,N_23965,N_24128);
nor UO_457 (O_457,N_24988,N_24927);
or UO_458 (O_458,N_24736,N_23989);
nand UO_459 (O_459,N_24456,N_24817);
nor UO_460 (O_460,N_24906,N_24887);
xor UO_461 (O_461,N_23879,N_24363);
xnor UO_462 (O_462,N_24327,N_23852);
and UO_463 (O_463,N_24871,N_24609);
and UO_464 (O_464,N_24074,N_24347);
or UO_465 (O_465,N_24518,N_23863);
nor UO_466 (O_466,N_24743,N_24236);
and UO_467 (O_467,N_24775,N_24451);
or UO_468 (O_468,N_24161,N_24187);
or UO_469 (O_469,N_23786,N_23822);
nand UO_470 (O_470,N_23906,N_24993);
and UO_471 (O_471,N_24846,N_24928);
nand UO_472 (O_472,N_24985,N_24424);
or UO_473 (O_473,N_24826,N_24797);
nand UO_474 (O_474,N_23825,N_24130);
and UO_475 (O_475,N_24762,N_24802);
nand UO_476 (O_476,N_24408,N_24081);
xnor UO_477 (O_477,N_24172,N_23798);
or UO_478 (O_478,N_24040,N_24789);
nor UO_479 (O_479,N_24330,N_24430);
and UO_480 (O_480,N_24756,N_23837);
nor UO_481 (O_481,N_24192,N_24067);
and UO_482 (O_482,N_23999,N_24877);
xnor UO_483 (O_483,N_24488,N_23995);
xor UO_484 (O_484,N_24467,N_24120);
xor UO_485 (O_485,N_24537,N_24587);
xor UO_486 (O_486,N_23933,N_24914);
xnor UO_487 (O_487,N_24628,N_24621);
nor UO_488 (O_488,N_24931,N_23783);
and UO_489 (O_489,N_24507,N_24140);
xor UO_490 (O_490,N_23973,N_24220);
or UO_491 (O_491,N_23772,N_24148);
or UO_492 (O_492,N_23958,N_24819);
nand UO_493 (O_493,N_23762,N_24117);
nand UO_494 (O_494,N_24551,N_24574);
xor UO_495 (O_495,N_24880,N_24058);
xnor UO_496 (O_496,N_24915,N_24266);
and UO_497 (O_497,N_24243,N_23880);
nand UO_498 (O_498,N_24486,N_24944);
xor UO_499 (O_499,N_24724,N_24862);
xor UO_500 (O_500,N_24176,N_24428);
and UO_501 (O_501,N_23754,N_24092);
or UO_502 (O_502,N_23895,N_24516);
nor UO_503 (O_503,N_24695,N_24023);
nand UO_504 (O_504,N_24952,N_24911);
nor UO_505 (O_505,N_23804,N_24473);
or UO_506 (O_506,N_24697,N_24101);
xor UO_507 (O_507,N_23940,N_24566);
or UO_508 (O_508,N_23826,N_24374);
nor UO_509 (O_509,N_23780,N_24385);
nand UO_510 (O_510,N_24210,N_24667);
or UO_511 (O_511,N_23841,N_24748);
xnor UO_512 (O_512,N_24476,N_24722);
xor UO_513 (O_513,N_24393,N_23971);
or UO_514 (O_514,N_24317,N_24637);
or UO_515 (O_515,N_23986,N_24095);
and UO_516 (O_516,N_24068,N_23752);
nor UO_517 (O_517,N_24687,N_24873);
nand UO_518 (O_518,N_24666,N_24169);
nand UO_519 (O_519,N_24131,N_23928);
nor UO_520 (O_520,N_23987,N_24409);
nand UO_521 (O_521,N_24800,N_24185);
nand UO_522 (O_522,N_24934,N_24865);
nor UO_523 (O_523,N_24859,N_23938);
or UO_524 (O_524,N_24870,N_23904);
nand UO_525 (O_525,N_24028,N_24703);
nor UO_526 (O_526,N_24959,N_24102);
nor UO_527 (O_527,N_24310,N_24214);
xnor UO_528 (O_528,N_24874,N_23957);
and UO_529 (O_529,N_23850,N_24654);
xnor UO_530 (O_530,N_24534,N_24702);
or UO_531 (O_531,N_24066,N_24807);
and UO_532 (O_532,N_24112,N_24730);
and UO_533 (O_533,N_24477,N_23807);
nor UO_534 (O_534,N_24173,N_24705);
nand UO_535 (O_535,N_24976,N_24153);
nor UO_536 (O_536,N_23771,N_23765);
or UO_537 (O_537,N_24003,N_24542);
nand UO_538 (O_538,N_24079,N_23993);
or UO_539 (O_539,N_23952,N_24269);
xnor UO_540 (O_540,N_24392,N_24739);
xor UO_541 (O_541,N_24201,N_24241);
or UO_542 (O_542,N_24293,N_24244);
nand UO_543 (O_543,N_24980,N_24468);
or UO_544 (O_544,N_23794,N_24525);
nor UO_545 (O_545,N_24322,N_24755);
or UO_546 (O_546,N_24069,N_24429);
nor UO_547 (O_547,N_24205,N_24086);
xnor UO_548 (O_548,N_23768,N_23810);
and UO_549 (O_549,N_24290,N_24820);
nor UO_550 (O_550,N_24413,N_24564);
and UO_551 (O_551,N_23861,N_24078);
nor UO_552 (O_552,N_23788,N_23814);
nand UO_553 (O_553,N_23956,N_24726);
xor UO_554 (O_554,N_24008,N_23836);
nand UO_555 (O_555,N_24717,N_24283);
xnor UO_556 (O_556,N_24027,N_24852);
xnor UO_557 (O_557,N_24805,N_24225);
nand UO_558 (O_558,N_24651,N_24640);
nor UO_559 (O_559,N_24369,N_23893);
or UO_560 (O_560,N_24024,N_24121);
nor UO_561 (O_561,N_24405,N_23922);
and UO_562 (O_562,N_24377,N_24622);
nor UO_563 (O_563,N_24816,N_24026);
and UO_564 (O_564,N_24049,N_24487);
or UO_565 (O_565,N_23824,N_24615);
or UO_566 (O_566,N_24281,N_24398);
nor UO_567 (O_567,N_24848,N_24930);
nand UO_568 (O_568,N_24104,N_24199);
or UO_569 (O_569,N_24014,N_24447);
xnor UO_570 (O_570,N_24834,N_24968);
or UO_571 (O_571,N_24941,N_23865);
and UO_572 (O_572,N_23787,N_24513);
and UO_573 (O_573,N_23757,N_24050);
nor UO_574 (O_574,N_24208,N_23809);
nand UO_575 (O_575,N_24905,N_23829);
xnor UO_576 (O_576,N_24760,N_24114);
nor UO_577 (O_577,N_24107,N_24136);
xnor UO_578 (O_578,N_24017,N_24563);
nor UO_579 (O_579,N_24177,N_23753);
nand UO_580 (O_580,N_24450,N_24925);
nor UO_581 (O_581,N_24514,N_24215);
nand UO_582 (O_582,N_24573,N_24292);
nand UO_583 (O_583,N_24426,N_24766);
or UO_584 (O_584,N_24308,N_24670);
and UO_585 (O_585,N_24818,N_23900);
or UO_586 (O_586,N_24005,N_24100);
and UO_587 (O_587,N_24593,N_24334);
and UO_588 (O_588,N_24882,N_23868);
and UO_589 (O_589,N_24822,N_24971);
xnor UO_590 (O_590,N_24740,N_23805);
xnor UO_591 (O_591,N_24658,N_23934);
and UO_592 (O_592,N_24791,N_24420);
nand UO_593 (O_593,N_23844,N_23876);
xnor UO_594 (O_594,N_24523,N_24174);
xnor UO_595 (O_595,N_24246,N_24864);
nand UO_596 (O_596,N_24629,N_23941);
nand UO_597 (O_597,N_24987,N_24603);
nor UO_598 (O_598,N_24854,N_24707);
or UO_599 (O_599,N_24901,N_24929);
and UO_600 (O_600,N_24964,N_24909);
or UO_601 (O_601,N_24989,N_24156);
xnor UO_602 (O_602,N_24422,N_24245);
nor UO_603 (O_603,N_24190,N_23776);
and UO_604 (O_604,N_24421,N_24919);
xnor UO_605 (O_605,N_24213,N_24029);
xnor UO_606 (O_606,N_24561,N_24261);
nor UO_607 (O_607,N_24464,N_24072);
and UO_608 (O_608,N_24735,N_24858);
xor UO_609 (O_609,N_24647,N_24841);
or UO_610 (O_610,N_23888,N_24025);
nor UO_611 (O_611,N_24378,N_23967);
and UO_612 (O_612,N_24768,N_23947);
and UO_613 (O_613,N_24831,N_24297);
and UO_614 (O_614,N_24071,N_24394);
nand UO_615 (O_615,N_24084,N_23813);
nor UO_616 (O_616,N_24616,N_24823);
or UO_617 (O_617,N_24321,N_24085);
nor UO_618 (O_618,N_24497,N_23847);
nor UO_619 (O_619,N_24361,N_24986);
and UO_620 (O_620,N_23828,N_24519);
xnor UO_621 (O_621,N_23979,N_24509);
xor UO_622 (O_622,N_24035,N_24033);
xnor UO_623 (O_623,N_24751,N_24251);
nor UO_624 (O_624,N_24767,N_24607);
nor UO_625 (O_625,N_24637,N_23843);
nor UO_626 (O_626,N_23783,N_24431);
nor UO_627 (O_627,N_23786,N_24095);
and UO_628 (O_628,N_23931,N_24885);
xnor UO_629 (O_629,N_24246,N_24826);
and UO_630 (O_630,N_24230,N_23778);
and UO_631 (O_631,N_23822,N_24895);
and UO_632 (O_632,N_24756,N_23881);
xnor UO_633 (O_633,N_23992,N_24541);
nor UO_634 (O_634,N_24059,N_23861);
xor UO_635 (O_635,N_24680,N_24512);
nand UO_636 (O_636,N_24539,N_24031);
nor UO_637 (O_637,N_24243,N_24635);
nor UO_638 (O_638,N_24712,N_24357);
xor UO_639 (O_639,N_24295,N_24577);
nor UO_640 (O_640,N_24928,N_24545);
xnor UO_641 (O_641,N_23985,N_24765);
or UO_642 (O_642,N_24233,N_23888);
nand UO_643 (O_643,N_24509,N_24175);
or UO_644 (O_644,N_24339,N_24158);
and UO_645 (O_645,N_24662,N_24846);
nor UO_646 (O_646,N_24112,N_24348);
or UO_647 (O_647,N_24992,N_23921);
nand UO_648 (O_648,N_24658,N_24398);
and UO_649 (O_649,N_24832,N_24973);
nor UO_650 (O_650,N_24673,N_24735);
nand UO_651 (O_651,N_24167,N_24841);
or UO_652 (O_652,N_24287,N_24029);
nand UO_653 (O_653,N_24576,N_23784);
xor UO_654 (O_654,N_24221,N_24478);
nand UO_655 (O_655,N_24501,N_24689);
or UO_656 (O_656,N_24615,N_23800);
or UO_657 (O_657,N_23856,N_23928);
nand UO_658 (O_658,N_24271,N_24086);
and UO_659 (O_659,N_24925,N_24447);
nand UO_660 (O_660,N_23846,N_24629);
and UO_661 (O_661,N_24594,N_24383);
nand UO_662 (O_662,N_24041,N_23977);
nand UO_663 (O_663,N_24279,N_24349);
nand UO_664 (O_664,N_24190,N_24262);
nand UO_665 (O_665,N_23789,N_24264);
and UO_666 (O_666,N_24202,N_24577);
xor UO_667 (O_667,N_24346,N_23857);
nand UO_668 (O_668,N_24774,N_24113);
and UO_669 (O_669,N_24867,N_24560);
nor UO_670 (O_670,N_23960,N_23976);
xor UO_671 (O_671,N_24002,N_24590);
nor UO_672 (O_672,N_24216,N_24592);
nor UO_673 (O_673,N_24899,N_24565);
and UO_674 (O_674,N_24701,N_24639);
or UO_675 (O_675,N_24848,N_24727);
and UO_676 (O_676,N_24105,N_24585);
and UO_677 (O_677,N_24955,N_24903);
xor UO_678 (O_678,N_24816,N_24674);
nand UO_679 (O_679,N_24091,N_24637);
nand UO_680 (O_680,N_23918,N_24827);
and UO_681 (O_681,N_24118,N_24718);
xor UO_682 (O_682,N_24548,N_24032);
and UO_683 (O_683,N_24860,N_24911);
xor UO_684 (O_684,N_23807,N_23782);
nand UO_685 (O_685,N_24958,N_24976);
nor UO_686 (O_686,N_24474,N_24433);
and UO_687 (O_687,N_24273,N_24657);
nor UO_688 (O_688,N_24390,N_24695);
xor UO_689 (O_689,N_23789,N_24281);
nor UO_690 (O_690,N_24229,N_24919);
nor UO_691 (O_691,N_24849,N_24753);
and UO_692 (O_692,N_24481,N_24903);
nor UO_693 (O_693,N_24643,N_24752);
xnor UO_694 (O_694,N_24646,N_24859);
nor UO_695 (O_695,N_23877,N_24582);
and UO_696 (O_696,N_24228,N_24536);
nor UO_697 (O_697,N_24300,N_24790);
or UO_698 (O_698,N_24333,N_24794);
xnor UO_699 (O_699,N_24726,N_23778);
xnor UO_700 (O_700,N_24628,N_24259);
nor UO_701 (O_701,N_24490,N_24404);
or UO_702 (O_702,N_23869,N_24578);
or UO_703 (O_703,N_24124,N_23762);
xnor UO_704 (O_704,N_24142,N_24789);
and UO_705 (O_705,N_24813,N_24396);
and UO_706 (O_706,N_24082,N_24030);
xor UO_707 (O_707,N_24283,N_23967);
or UO_708 (O_708,N_24085,N_24732);
and UO_709 (O_709,N_23863,N_24514);
nand UO_710 (O_710,N_24876,N_24509);
xor UO_711 (O_711,N_24576,N_24936);
nand UO_712 (O_712,N_24406,N_24914);
nor UO_713 (O_713,N_24185,N_23901);
and UO_714 (O_714,N_23911,N_24247);
or UO_715 (O_715,N_24202,N_24061);
nor UO_716 (O_716,N_24178,N_24577);
nor UO_717 (O_717,N_24263,N_23830);
nor UO_718 (O_718,N_24711,N_23924);
and UO_719 (O_719,N_23832,N_24030);
nand UO_720 (O_720,N_24421,N_24520);
and UO_721 (O_721,N_24056,N_23761);
and UO_722 (O_722,N_24513,N_24242);
and UO_723 (O_723,N_23841,N_23952);
or UO_724 (O_724,N_24893,N_24797);
and UO_725 (O_725,N_23851,N_24175);
and UO_726 (O_726,N_24524,N_23790);
nor UO_727 (O_727,N_24227,N_24460);
or UO_728 (O_728,N_24909,N_24183);
and UO_729 (O_729,N_24724,N_24221);
and UO_730 (O_730,N_24899,N_24109);
or UO_731 (O_731,N_24089,N_24945);
nor UO_732 (O_732,N_23761,N_23833);
nand UO_733 (O_733,N_24756,N_24624);
xor UO_734 (O_734,N_24629,N_24980);
xor UO_735 (O_735,N_24704,N_24775);
nor UO_736 (O_736,N_23820,N_24229);
and UO_737 (O_737,N_24029,N_24382);
xor UO_738 (O_738,N_24991,N_24249);
xnor UO_739 (O_739,N_24621,N_24915);
nand UO_740 (O_740,N_23902,N_24752);
nor UO_741 (O_741,N_24525,N_24006);
nor UO_742 (O_742,N_24244,N_24103);
nor UO_743 (O_743,N_24595,N_23954);
or UO_744 (O_744,N_24360,N_23823);
and UO_745 (O_745,N_24449,N_24670);
and UO_746 (O_746,N_24487,N_24118);
and UO_747 (O_747,N_24953,N_23873);
or UO_748 (O_748,N_24932,N_24643);
and UO_749 (O_749,N_23891,N_24794);
nor UO_750 (O_750,N_24096,N_24507);
or UO_751 (O_751,N_24373,N_24271);
nor UO_752 (O_752,N_24559,N_24102);
nor UO_753 (O_753,N_24310,N_23992);
xor UO_754 (O_754,N_24754,N_24442);
and UO_755 (O_755,N_23881,N_23813);
xnor UO_756 (O_756,N_24047,N_24819);
or UO_757 (O_757,N_24807,N_23901);
or UO_758 (O_758,N_24980,N_24357);
or UO_759 (O_759,N_24047,N_24068);
or UO_760 (O_760,N_24572,N_24874);
or UO_761 (O_761,N_24657,N_24407);
nand UO_762 (O_762,N_24501,N_24465);
and UO_763 (O_763,N_24684,N_24340);
xnor UO_764 (O_764,N_24886,N_24831);
xnor UO_765 (O_765,N_24427,N_23806);
nand UO_766 (O_766,N_24608,N_24671);
xor UO_767 (O_767,N_24052,N_23974);
nand UO_768 (O_768,N_23971,N_24913);
nand UO_769 (O_769,N_24580,N_24737);
nand UO_770 (O_770,N_23882,N_24410);
and UO_771 (O_771,N_24466,N_24866);
or UO_772 (O_772,N_24535,N_24814);
nor UO_773 (O_773,N_24801,N_24914);
xnor UO_774 (O_774,N_24530,N_24282);
xnor UO_775 (O_775,N_24043,N_24819);
nand UO_776 (O_776,N_24781,N_23765);
nor UO_777 (O_777,N_24358,N_24320);
and UO_778 (O_778,N_23779,N_24011);
xor UO_779 (O_779,N_24786,N_24380);
xor UO_780 (O_780,N_24267,N_24647);
xnor UO_781 (O_781,N_24725,N_24594);
or UO_782 (O_782,N_24223,N_24945);
and UO_783 (O_783,N_23758,N_23791);
nand UO_784 (O_784,N_24996,N_24447);
nor UO_785 (O_785,N_24228,N_24850);
or UO_786 (O_786,N_24814,N_23892);
or UO_787 (O_787,N_23891,N_24230);
xnor UO_788 (O_788,N_24821,N_24369);
or UO_789 (O_789,N_24265,N_24883);
and UO_790 (O_790,N_23775,N_24165);
nor UO_791 (O_791,N_23828,N_24326);
nand UO_792 (O_792,N_24842,N_24475);
or UO_793 (O_793,N_24093,N_24378);
nor UO_794 (O_794,N_24190,N_24638);
nor UO_795 (O_795,N_24424,N_24083);
nand UO_796 (O_796,N_24556,N_24833);
or UO_797 (O_797,N_24672,N_24087);
or UO_798 (O_798,N_24848,N_24915);
or UO_799 (O_799,N_24505,N_24248);
or UO_800 (O_800,N_23959,N_24687);
xnor UO_801 (O_801,N_24873,N_24693);
nand UO_802 (O_802,N_24714,N_23947);
nand UO_803 (O_803,N_24879,N_23955);
nor UO_804 (O_804,N_24345,N_24818);
nand UO_805 (O_805,N_24822,N_24777);
and UO_806 (O_806,N_24833,N_24686);
nand UO_807 (O_807,N_23988,N_24526);
xor UO_808 (O_808,N_24621,N_24425);
nand UO_809 (O_809,N_24579,N_23959);
nand UO_810 (O_810,N_24903,N_24679);
and UO_811 (O_811,N_24515,N_23899);
and UO_812 (O_812,N_23868,N_24551);
nand UO_813 (O_813,N_24776,N_24631);
nor UO_814 (O_814,N_24472,N_24047);
and UO_815 (O_815,N_24881,N_24065);
and UO_816 (O_816,N_24772,N_24218);
nand UO_817 (O_817,N_24874,N_24784);
and UO_818 (O_818,N_24141,N_24395);
nand UO_819 (O_819,N_24797,N_23810);
xor UO_820 (O_820,N_24214,N_24402);
xor UO_821 (O_821,N_24478,N_23967);
nand UO_822 (O_822,N_24053,N_24613);
nand UO_823 (O_823,N_24639,N_24871);
xor UO_824 (O_824,N_23951,N_24698);
nand UO_825 (O_825,N_24192,N_24484);
nand UO_826 (O_826,N_24031,N_24463);
or UO_827 (O_827,N_24847,N_24656);
xnor UO_828 (O_828,N_24083,N_24545);
nor UO_829 (O_829,N_24814,N_24156);
nand UO_830 (O_830,N_24098,N_23912);
and UO_831 (O_831,N_24463,N_24236);
nor UO_832 (O_832,N_23797,N_24906);
nor UO_833 (O_833,N_24033,N_24754);
or UO_834 (O_834,N_24826,N_24180);
nor UO_835 (O_835,N_23970,N_24523);
or UO_836 (O_836,N_24002,N_24105);
nand UO_837 (O_837,N_24292,N_23973);
xor UO_838 (O_838,N_24414,N_23874);
nand UO_839 (O_839,N_24418,N_24384);
nor UO_840 (O_840,N_24778,N_23862);
xnor UO_841 (O_841,N_24428,N_24787);
and UO_842 (O_842,N_24041,N_24033);
xor UO_843 (O_843,N_24142,N_24805);
and UO_844 (O_844,N_24898,N_24415);
nand UO_845 (O_845,N_24601,N_23772);
or UO_846 (O_846,N_24496,N_24054);
nor UO_847 (O_847,N_24224,N_23811);
xnor UO_848 (O_848,N_24293,N_23894);
nand UO_849 (O_849,N_24597,N_24922);
xor UO_850 (O_850,N_24016,N_23768);
or UO_851 (O_851,N_24791,N_24634);
or UO_852 (O_852,N_24048,N_24088);
nor UO_853 (O_853,N_24776,N_24065);
xnor UO_854 (O_854,N_24457,N_23792);
nand UO_855 (O_855,N_24632,N_24890);
or UO_856 (O_856,N_24543,N_23949);
nand UO_857 (O_857,N_24942,N_23856);
xor UO_858 (O_858,N_23873,N_24466);
or UO_859 (O_859,N_24598,N_24503);
or UO_860 (O_860,N_23871,N_24607);
xnor UO_861 (O_861,N_24361,N_24858);
nor UO_862 (O_862,N_23790,N_24858);
xor UO_863 (O_863,N_24194,N_23792);
and UO_864 (O_864,N_24948,N_24087);
xor UO_865 (O_865,N_24568,N_24042);
nor UO_866 (O_866,N_24342,N_24944);
or UO_867 (O_867,N_24161,N_24015);
and UO_868 (O_868,N_24008,N_23906);
nand UO_869 (O_869,N_24836,N_24442);
and UO_870 (O_870,N_24351,N_24940);
xor UO_871 (O_871,N_24419,N_24679);
or UO_872 (O_872,N_24625,N_23867);
xnor UO_873 (O_873,N_23844,N_24076);
nor UO_874 (O_874,N_24361,N_24052);
and UO_875 (O_875,N_24652,N_24360);
nor UO_876 (O_876,N_24466,N_24701);
nor UO_877 (O_877,N_24307,N_24052);
nand UO_878 (O_878,N_24665,N_24587);
nor UO_879 (O_879,N_24304,N_24065);
nor UO_880 (O_880,N_24284,N_24452);
nand UO_881 (O_881,N_24892,N_24514);
nor UO_882 (O_882,N_24530,N_23977);
or UO_883 (O_883,N_24561,N_24103);
xor UO_884 (O_884,N_24533,N_23987);
nor UO_885 (O_885,N_24045,N_24973);
nand UO_886 (O_886,N_23886,N_24535);
and UO_887 (O_887,N_24703,N_24921);
nand UO_888 (O_888,N_24142,N_24667);
nor UO_889 (O_889,N_24305,N_23847);
nor UO_890 (O_890,N_23896,N_24104);
or UO_891 (O_891,N_23892,N_24031);
nor UO_892 (O_892,N_24026,N_24741);
xnor UO_893 (O_893,N_24334,N_24953);
nand UO_894 (O_894,N_24194,N_24147);
xor UO_895 (O_895,N_23926,N_24345);
nand UO_896 (O_896,N_23828,N_23845);
or UO_897 (O_897,N_24216,N_24978);
xor UO_898 (O_898,N_24757,N_23997);
or UO_899 (O_899,N_24179,N_24036);
xor UO_900 (O_900,N_24469,N_24301);
and UO_901 (O_901,N_23818,N_23929);
nand UO_902 (O_902,N_24179,N_24044);
nand UO_903 (O_903,N_23820,N_24348);
xor UO_904 (O_904,N_24057,N_24603);
or UO_905 (O_905,N_24555,N_24387);
or UO_906 (O_906,N_23819,N_24503);
xor UO_907 (O_907,N_24414,N_23911);
or UO_908 (O_908,N_24519,N_23900);
or UO_909 (O_909,N_23847,N_24580);
or UO_910 (O_910,N_24250,N_24736);
nand UO_911 (O_911,N_24670,N_24744);
and UO_912 (O_912,N_24463,N_24586);
or UO_913 (O_913,N_24534,N_24911);
and UO_914 (O_914,N_24079,N_24212);
nand UO_915 (O_915,N_24333,N_24690);
or UO_916 (O_916,N_24991,N_24185);
and UO_917 (O_917,N_24145,N_24446);
nand UO_918 (O_918,N_23974,N_24198);
or UO_919 (O_919,N_24817,N_24393);
xnor UO_920 (O_920,N_23928,N_23881);
nor UO_921 (O_921,N_24555,N_24348);
and UO_922 (O_922,N_24707,N_23920);
and UO_923 (O_923,N_24739,N_24332);
or UO_924 (O_924,N_24320,N_24423);
and UO_925 (O_925,N_23921,N_23761);
xnor UO_926 (O_926,N_24086,N_24981);
xor UO_927 (O_927,N_24752,N_24947);
or UO_928 (O_928,N_24400,N_24908);
and UO_929 (O_929,N_23811,N_23952);
or UO_930 (O_930,N_24497,N_23960);
nor UO_931 (O_931,N_24380,N_23908);
nand UO_932 (O_932,N_23890,N_23887);
nand UO_933 (O_933,N_24834,N_24477);
and UO_934 (O_934,N_24698,N_24451);
nand UO_935 (O_935,N_24135,N_23766);
nand UO_936 (O_936,N_24248,N_24436);
nor UO_937 (O_937,N_24540,N_24719);
nor UO_938 (O_938,N_23937,N_24288);
and UO_939 (O_939,N_24083,N_24888);
nor UO_940 (O_940,N_24610,N_24440);
xnor UO_941 (O_941,N_24761,N_24828);
or UO_942 (O_942,N_24102,N_24930);
xor UO_943 (O_943,N_24118,N_24282);
and UO_944 (O_944,N_24954,N_24348);
nor UO_945 (O_945,N_24619,N_24232);
xnor UO_946 (O_946,N_24346,N_23901);
nand UO_947 (O_947,N_24946,N_23877);
and UO_948 (O_948,N_24182,N_24310);
or UO_949 (O_949,N_24542,N_24147);
nor UO_950 (O_950,N_24499,N_24128);
nor UO_951 (O_951,N_24294,N_24789);
or UO_952 (O_952,N_24960,N_24345);
or UO_953 (O_953,N_24832,N_24804);
nand UO_954 (O_954,N_23770,N_24714);
or UO_955 (O_955,N_24396,N_23992);
nor UO_956 (O_956,N_24074,N_23914);
xnor UO_957 (O_957,N_24251,N_24125);
or UO_958 (O_958,N_24989,N_24396);
xor UO_959 (O_959,N_24566,N_23987);
and UO_960 (O_960,N_23812,N_24754);
nand UO_961 (O_961,N_23764,N_23936);
and UO_962 (O_962,N_24566,N_24784);
or UO_963 (O_963,N_24757,N_24836);
nand UO_964 (O_964,N_24221,N_24051);
or UO_965 (O_965,N_24405,N_23998);
nor UO_966 (O_966,N_24779,N_24485);
nor UO_967 (O_967,N_24334,N_24192);
nand UO_968 (O_968,N_23793,N_24333);
xor UO_969 (O_969,N_24208,N_24696);
nand UO_970 (O_970,N_23788,N_23848);
nor UO_971 (O_971,N_24991,N_23849);
or UO_972 (O_972,N_24733,N_24586);
and UO_973 (O_973,N_24136,N_24461);
nor UO_974 (O_974,N_24701,N_24803);
or UO_975 (O_975,N_24585,N_24744);
xnor UO_976 (O_976,N_23894,N_24887);
nor UO_977 (O_977,N_23757,N_24160);
or UO_978 (O_978,N_24852,N_24322);
nor UO_979 (O_979,N_24338,N_23982);
nand UO_980 (O_980,N_24831,N_24106);
nand UO_981 (O_981,N_24017,N_23766);
xnor UO_982 (O_982,N_24586,N_24291);
and UO_983 (O_983,N_24112,N_23819);
and UO_984 (O_984,N_23924,N_23860);
and UO_985 (O_985,N_23900,N_24698);
nand UO_986 (O_986,N_24488,N_23806);
and UO_987 (O_987,N_24614,N_24000);
nor UO_988 (O_988,N_24134,N_24290);
nand UO_989 (O_989,N_24682,N_24838);
nor UO_990 (O_990,N_24724,N_24218);
xor UO_991 (O_991,N_24739,N_24469);
and UO_992 (O_992,N_24221,N_24361);
nor UO_993 (O_993,N_24386,N_24276);
or UO_994 (O_994,N_24377,N_24298);
nand UO_995 (O_995,N_23792,N_23888);
or UO_996 (O_996,N_24448,N_24944);
nand UO_997 (O_997,N_24097,N_24824);
nand UO_998 (O_998,N_24604,N_24300);
nor UO_999 (O_999,N_24476,N_24316);
or UO_1000 (O_1000,N_24594,N_24493);
or UO_1001 (O_1001,N_23778,N_24768);
xnor UO_1002 (O_1002,N_24595,N_24555);
nand UO_1003 (O_1003,N_24248,N_23877);
nor UO_1004 (O_1004,N_23935,N_24361);
and UO_1005 (O_1005,N_24470,N_23834);
nand UO_1006 (O_1006,N_24423,N_24304);
nand UO_1007 (O_1007,N_24405,N_24702);
nor UO_1008 (O_1008,N_24266,N_24714);
nor UO_1009 (O_1009,N_24491,N_24871);
nand UO_1010 (O_1010,N_24317,N_24470);
nand UO_1011 (O_1011,N_24378,N_23791);
nor UO_1012 (O_1012,N_24100,N_24312);
and UO_1013 (O_1013,N_23900,N_24574);
nand UO_1014 (O_1014,N_24281,N_24456);
or UO_1015 (O_1015,N_24541,N_24536);
nand UO_1016 (O_1016,N_24800,N_24318);
nand UO_1017 (O_1017,N_24530,N_23878);
and UO_1018 (O_1018,N_24880,N_24700);
xnor UO_1019 (O_1019,N_24419,N_24230);
and UO_1020 (O_1020,N_24145,N_24407);
xor UO_1021 (O_1021,N_24037,N_24977);
nor UO_1022 (O_1022,N_24285,N_24163);
nor UO_1023 (O_1023,N_24502,N_23857);
nor UO_1024 (O_1024,N_24840,N_24083);
nor UO_1025 (O_1025,N_24552,N_23936);
nor UO_1026 (O_1026,N_24636,N_24990);
xor UO_1027 (O_1027,N_24415,N_24831);
and UO_1028 (O_1028,N_24304,N_24876);
xor UO_1029 (O_1029,N_24193,N_24770);
or UO_1030 (O_1030,N_24914,N_24294);
or UO_1031 (O_1031,N_24818,N_24467);
or UO_1032 (O_1032,N_24742,N_24920);
nand UO_1033 (O_1033,N_24821,N_24764);
xor UO_1034 (O_1034,N_24364,N_23796);
and UO_1035 (O_1035,N_24323,N_24040);
and UO_1036 (O_1036,N_23835,N_23971);
nand UO_1037 (O_1037,N_24989,N_24057);
xnor UO_1038 (O_1038,N_24866,N_24199);
nor UO_1039 (O_1039,N_24193,N_24312);
and UO_1040 (O_1040,N_24095,N_24463);
nand UO_1041 (O_1041,N_23773,N_24051);
nor UO_1042 (O_1042,N_24068,N_24418);
and UO_1043 (O_1043,N_24672,N_24000);
and UO_1044 (O_1044,N_24430,N_24787);
or UO_1045 (O_1045,N_24050,N_24253);
or UO_1046 (O_1046,N_24314,N_24484);
nand UO_1047 (O_1047,N_24337,N_24247);
nor UO_1048 (O_1048,N_23862,N_24699);
or UO_1049 (O_1049,N_24175,N_24021);
and UO_1050 (O_1050,N_23840,N_24324);
xnor UO_1051 (O_1051,N_24411,N_24667);
nand UO_1052 (O_1052,N_23753,N_24610);
and UO_1053 (O_1053,N_24046,N_24222);
and UO_1054 (O_1054,N_24973,N_24141);
nor UO_1055 (O_1055,N_24457,N_24101);
nand UO_1056 (O_1056,N_24454,N_23785);
xor UO_1057 (O_1057,N_24615,N_24384);
nand UO_1058 (O_1058,N_24637,N_24448);
and UO_1059 (O_1059,N_23942,N_23868);
nor UO_1060 (O_1060,N_24041,N_24463);
xnor UO_1061 (O_1061,N_24794,N_23912);
nand UO_1062 (O_1062,N_24143,N_23887);
or UO_1063 (O_1063,N_24809,N_24557);
nand UO_1064 (O_1064,N_23970,N_23987);
and UO_1065 (O_1065,N_23755,N_24804);
nand UO_1066 (O_1066,N_24075,N_24693);
nor UO_1067 (O_1067,N_24399,N_24164);
or UO_1068 (O_1068,N_24891,N_24840);
nor UO_1069 (O_1069,N_24512,N_24808);
nand UO_1070 (O_1070,N_24721,N_24167);
nand UO_1071 (O_1071,N_24801,N_24284);
and UO_1072 (O_1072,N_24188,N_24933);
nor UO_1073 (O_1073,N_24626,N_24976);
and UO_1074 (O_1074,N_24981,N_24608);
nor UO_1075 (O_1075,N_24748,N_24989);
or UO_1076 (O_1076,N_24425,N_24987);
and UO_1077 (O_1077,N_24244,N_24966);
xor UO_1078 (O_1078,N_24274,N_23794);
nand UO_1079 (O_1079,N_24064,N_24234);
xor UO_1080 (O_1080,N_24813,N_23959);
nor UO_1081 (O_1081,N_24663,N_24609);
xnor UO_1082 (O_1082,N_23928,N_24998);
xnor UO_1083 (O_1083,N_24228,N_23959);
nand UO_1084 (O_1084,N_24181,N_23774);
or UO_1085 (O_1085,N_23813,N_24553);
and UO_1086 (O_1086,N_24120,N_23891);
or UO_1087 (O_1087,N_23772,N_24489);
nor UO_1088 (O_1088,N_24881,N_24655);
or UO_1089 (O_1089,N_24301,N_24711);
or UO_1090 (O_1090,N_24063,N_24056);
nand UO_1091 (O_1091,N_24481,N_24593);
and UO_1092 (O_1092,N_24631,N_24944);
or UO_1093 (O_1093,N_24528,N_23874);
and UO_1094 (O_1094,N_23789,N_24275);
and UO_1095 (O_1095,N_24814,N_24161);
nand UO_1096 (O_1096,N_24127,N_23849);
xnor UO_1097 (O_1097,N_23923,N_23849);
and UO_1098 (O_1098,N_24761,N_24050);
nand UO_1099 (O_1099,N_24650,N_24315);
xnor UO_1100 (O_1100,N_24189,N_24858);
nor UO_1101 (O_1101,N_23826,N_24560);
nand UO_1102 (O_1102,N_24303,N_23778);
and UO_1103 (O_1103,N_24663,N_24529);
or UO_1104 (O_1104,N_24180,N_24955);
and UO_1105 (O_1105,N_23760,N_23862);
nor UO_1106 (O_1106,N_23776,N_24392);
xor UO_1107 (O_1107,N_24826,N_24949);
nand UO_1108 (O_1108,N_23781,N_24226);
nand UO_1109 (O_1109,N_24285,N_23779);
or UO_1110 (O_1110,N_24722,N_24836);
nor UO_1111 (O_1111,N_24070,N_24245);
and UO_1112 (O_1112,N_24964,N_23874);
or UO_1113 (O_1113,N_24489,N_24461);
xor UO_1114 (O_1114,N_23836,N_24418);
nand UO_1115 (O_1115,N_24501,N_24695);
nor UO_1116 (O_1116,N_24383,N_23989);
nand UO_1117 (O_1117,N_24828,N_24474);
xor UO_1118 (O_1118,N_24074,N_24791);
or UO_1119 (O_1119,N_23945,N_24688);
nand UO_1120 (O_1120,N_24721,N_24048);
nor UO_1121 (O_1121,N_23888,N_24127);
or UO_1122 (O_1122,N_24959,N_24141);
and UO_1123 (O_1123,N_24430,N_24840);
xnor UO_1124 (O_1124,N_24128,N_23886);
xnor UO_1125 (O_1125,N_24805,N_23784);
and UO_1126 (O_1126,N_24474,N_24243);
and UO_1127 (O_1127,N_24250,N_23826);
and UO_1128 (O_1128,N_24155,N_24008);
or UO_1129 (O_1129,N_24909,N_24890);
or UO_1130 (O_1130,N_23789,N_24945);
xnor UO_1131 (O_1131,N_24553,N_24036);
or UO_1132 (O_1132,N_24347,N_24456);
or UO_1133 (O_1133,N_23829,N_24366);
nand UO_1134 (O_1134,N_23881,N_24474);
and UO_1135 (O_1135,N_24594,N_24663);
or UO_1136 (O_1136,N_24431,N_24061);
and UO_1137 (O_1137,N_24714,N_24165);
nand UO_1138 (O_1138,N_24565,N_23899);
nand UO_1139 (O_1139,N_24307,N_23804);
nand UO_1140 (O_1140,N_23899,N_24518);
nor UO_1141 (O_1141,N_24196,N_24883);
nor UO_1142 (O_1142,N_24807,N_23814);
nand UO_1143 (O_1143,N_24670,N_24830);
nor UO_1144 (O_1144,N_24815,N_24567);
or UO_1145 (O_1145,N_24959,N_24846);
nand UO_1146 (O_1146,N_24319,N_23872);
xnor UO_1147 (O_1147,N_24745,N_24021);
and UO_1148 (O_1148,N_23847,N_24988);
xor UO_1149 (O_1149,N_24931,N_24093);
nor UO_1150 (O_1150,N_23908,N_24497);
or UO_1151 (O_1151,N_24450,N_23869);
xor UO_1152 (O_1152,N_24446,N_24990);
xor UO_1153 (O_1153,N_24079,N_24476);
xnor UO_1154 (O_1154,N_24648,N_24772);
nor UO_1155 (O_1155,N_24287,N_24646);
xor UO_1156 (O_1156,N_24675,N_24560);
xnor UO_1157 (O_1157,N_23846,N_23807);
nor UO_1158 (O_1158,N_24774,N_24887);
or UO_1159 (O_1159,N_24182,N_24900);
and UO_1160 (O_1160,N_23852,N_24824);
nor UO_1161 (O_1161,N_24493,N_24592);
nand UO_1162 (O_1162,N_23833,N_23886);
xor UO_1163 (O_1163,N_24717,N_23773);
nor UO_1164 (O_1164,N_24251,N_24907);
nor UO_1165 (O_1165,N_24263,N_23888);
and UO_1166 (O_1166,N_24695,N_24641);
nor UO_1167 (O_1167,N_24304,N_23767);
nor UO_1168 (O_1168,N_24598,N_23873);
and UO_1169 (O_1169,N_24993,N_23838);
xnor UO_1170 (O_1170,N_23994,N_24682);
or UO_1171 (O_1171,N_23888,N_24949);
nor UO_1172 (O_1172,N_24849,N_24022);
nor UO_1173 (O_1173,N_24050,N_23752);
nand UO_1174 (O_1174,N_24970,N_24843);
xor UO_1175 (O_1175,N_23885,N_24483);
or UO_1176 (O_1176,N_23886,N_24816);
nand UO_1177 (O_1177,N_24939,N_24535);
nor UO_1178 (O_1178,N_24858,N_23904);
nor UO_1179 (O_1179,N_24264,N_24150);
nor UO_1180 (O_1180,N_24628,N_24839);
nor UO_1181 (O_1181,N_24516,N_24778);
nand UO_1182 (O_1182,N_24155,N_24253);
and UO_1183 (O_1183,N_24953,N_24285);
and UO_1184 (O_1184,N_23763,N_24254);
nor UO_1185 (O_1185,N_23970,N_24253);
nor UO_1186 (O_1186,N_24880,N_24857);
xor UO_1187 (O_1187,N_23824,N_23766);
nand UO_1188 (O_1188,N_23928,N_24454);
and UO_1189 (O_1189,N_24885,N_24716);
nand UO_1190 (O_1190,N_24563,N_24662);
and UO_1191 (O_1191,N_23917,N_24129);
or UO_1192 (O_1192,N_24403,N_24432);
and UO_1193 (O_1193,N_24657,N_24181);
and UO_1194 (O_1194,N_24792,N_24877);
nand UO_1195 (O_1195,N_24786,N_24222);
or UO_1196 (O_1196,N_24264,N_23800);
and UO_1197 (O_1197,N_24508,N_24261);
and UO_1198 (O_1198,N_23792,N_24859);
nor UO_1199 (O_1199,N_24252,N_24046);
or UO_1200 (O_1200,N_24430,N_24547);
nor UO_1201 (O_1201,N_24184,N_24717);
or UO_1202 (O_1202,N_24323,N_24532);
or UO_1203 (O_1203,N_23777,N_24958);
nor UO_1204 (O_1204,N_23962,N_24430);
nand UO_1205 (O_1205,N_24679,N_24656);
nand UO_1206 (O_1206,N_24548,N_24173);
or UO_1207 (O_1207,N_24334,N_23945);
or UO_1208 (O_1208,N_24528,N_24110);
or UO_1209 (O_1209,N_23948,N_24238);
nor UO_1210 (O_1210,N_24808,N_24716);
xor UO_1211 (O_1211,N_24158,N_24822);
xor UO_1212 (O_1212,N_24589,N_23979);
nand UO_1213 (O_1213,N_24545,N_24429);
xor UO_1214 (O_1214,N_24391,N_24836);
xnor UO_1215 (O_1215,N_23916,N_24046);
and UO_1216 (O_1216,N_24191,N_24309);
or UO_1217 (O_1217,N_24315,N_23805);
xnor UO_1218 (O_1218,N_24852,N_24063);
nor UO_1219 (O_1219,N_24436,N_24072);
xor UO_1220 (O_1220,N_23780,N_24094);
and UO_1221 (O_1221,N_24728,N_24905);
xor UO_1222 (O_1222,N_24782,N_24091);
nand UO_1223 (O_1223,N_23820,N_24742);
and UO_1224 (O_1224,N_24362,N_24335);
and UO_1225 (O_1225,N_24463,N_24659);
or UO_1226 (O_1226,N_24848,N_23839);
or UO_1227 (O_1227,N_24343,N_24729);
nand UO_1228 (O_1228,N_24808,N_24416);
xnor UO_1229 (O_1229,N_24321,N_24399);
nor UO_1230 (O_1230,N_24278,N_24421);
xor UO_1231 (O_1231,N_24505,N_23837);
xnor UO_1232 (O_1232,N_23845,N_24240);
nor UO_1233 (O_1233,N_24893,N_23917);
nand UO_1234 (O_1234,N_24791,N_23766);
and UO_1235 (O_1235,N_24371,N_24479);
xnor UO_1236 (O_1236,N_24483,N_24706);
nor UO_1237 (O_1237,N_23767,N_24836);
nor UO_1238 (O_1238,N_24828,N_23760);
and UO_1239 (O_1239,N_24338,N_24543);
and UO_1240 (O_1240,N_23928,N_24866);
or UO_1241 (O_1241,N_23798,N_24171);
xor UO_1242 (O_1242,N_24353,N_24916);
xor UO_1243 (O_1243,N_24635,N_23991);
xnor UO_1244 (O_1244,N_24470,N_24107);
nor UO_1245 (O_1245,N_24310,N_24456);
nor UO_1246 (O_1246,N_24939,N_24703);
and UO_1247 (O_1247,N_24622,N_23882);
and UO_1248 (O_1248,N_24175,N_24965);
nor UO_1249 (O_1249,N_24283,N_24145);
nand UO_1250 (O_1250,N_24278,N_24500);
nor UO_1251 (O_1251,N_23836,N_23871);
and UO_1252 (O_1252,N_24004,N_24192);
xor UO_1253 (O_1253,N_24896,N_24310);
and UO_1254 (O_1254,N_24990,N_24943);
xnor UO_1255 (O_1255,N_24811,N_24274);
or UO_1256 (O_1256,N_24219,N_24485);
xnor UO_1257 (O_1257,N_24607,N_24625);
and UO_1258 (O_1258,N_24188,N_24037);
xor UO_1259 (O_1259,N_24831,N_23902);
nor UO_1260 (O_1260,N_23929,N_24752);
xor UO_1261 (O_1261,N_24742,N_24163);
xnor UO_1262 (O_1262,N_23798,N_24111);
xnor UO_1263 (O_1263,N_24121,N_24197);
nor UO_1264 (O_1264,N_24356,N_24528);
nand UO_1265 (O_1265,N_24256,N_24745);
nor UO_1266 (O_1266,N_23902,N_23979);
or UO_1267 (O_1267,N_23964,N_24692);
nor UO_1268 (O_1268,N_24607,N_24592);
or UO_1269 (O_1269,N_24239,N_24810);
or UO_1270 (O_1270,N_24923,N_24708);
nand UO_1271 (O_1271,N_24950,N_23880);
nor UO_1272 (O_1272,N_24593,N_24971);
xnor UO_1273 (O_1273,N_24461,N_24640);
nand UO_1274 (O_1274,N_24350,N_24019);
xnor UO_1275 (O_1275,N_24726,N_24180);
and UO_1276 (O_1276,N_24853,N_24528);
and UO_1277 (O_1277,N_23752,N_24342);
xor UO_1278 (O_1278,N_24904,N_24081);
and UO_1279 (O_1279,N_24390,N_23856);
nand UO_1280 (O_1280,N_24146,N_23893);
nor UO_1281 (O_1281,N_23985,N_24247);
and UO_1282 (O_1282,N_23872,N_24015);
xor UO_1283 (O_1283,N_24758,N_24364);
and UO_1284 (O_1284,N_23877,N_24040);
nor UO_1285 (O_1285,N_24109,N_24017);
nor UO_1286 (O_1286,N_24383,N_24384);
nor UO_1287 (O_1287,N_24408,N_24035);
xor UO_1288 (O_1288,N_24367,N_24178);
xnor UO_1289 (O_1289,N_24966,N_24469);
xor UO_1290 (O_1290,N_24042,N_24324);
xnor UO_1291 (O_1291,N_24957,N_24390);
and UO_1292 (O_1292,N_24260,N_24376);
or UO_1293 (O_1293,N_24500,N_24168);
nor UO_1294 (O_1294,N_23811,N_23907);
nand UO_1295 (O_1295,N_24650,N_24060);
xnor UO_1296 (O_1296,N_24535,N_24042);
or UO_1297 (O_1297,N_24551,N_24133);
and UO_1298 (O_1298,N_24828,N_24932);
nor UO_1299 (O_1299,N_23965,N_24857);
or UO_1300 (O_1300,N_24712,N_24069);
or UO_1301 (O_1301,N_24838,N_24935);
nor UO_1302 (O_1302,N_24739,N_24191);
xnor UO_1303 (O_1303,N_24412,N_24952);
and UO_1304 (O_1304,N_24746,N_24894);
and UO_1305 (O_1305,N_24508,N_24864);
xor UO_1306 (O_1306,N_24142,N_24165);
or UO_1307 (O_1307,N_24722,N_24138);
xor UO_1308 (O_1308,N_24408,N_24924);
xor UO_1309 (O_1309,N_24865,N_24216);
nor UO_1310 (O_1310,N_24082,N_24192);
or UO_1311 (O_1311,N_24886,N_24457);
xor UO_1312 (O_1312,N_24477,N_23931);
and UO_1313 (O_1313,N_24424,N_24987);
xor UO_1314 (O_1314,N_24922,N_24205);
and UO_1315 (O_1315,N_24046,N_24229);
nand UO_1316 (O_1316,N_23987,N_24929);
and UO_1317 (O_1317,N_24275,N_24317);
or UO_1318 (O_1318,N_24913,N_24151);
nand UO_1319 (O_1319,N_24731,N_23888);
or UO_1320 (O_1320,N_23768,N_24451);
and UO_1321 (O_1321,N_24414,N_24970);
nor UO_1322 (O_1322,N_24946,N_23886);
and UO_1323 (O_1323,N_24354,N_23812);
nand UO_1324 (O_1324,N_24513,N_24640);
and UO_1325 (O_1325,N_24249,N_24127);
or UO_1326 (O_1326,N_23874,N_23899);
and UO_1327 (O_1327,N_24163,N_24282);
nand UO_1328 (O_1328,N_24078,N_24561);
nand UO_1329 (O_1329,N_24033,N_24707);
xnor UO_1330 (O_1330,N_24609,N_24184);
and UO_1331 (O_1331,N_24533,N_24630);
nand UO_1332 (O_1332,N_23873,N_24997);
nand UO_1333 (O_1333,N_24305,N_24655);
nor UO_1334 (O_1334,N_24795,N_24861);
or UO_1335 (O_1335,N_23795,N_24065);
xnor UO_1336 (O_1336,N_24887,N_24776);
nand UO_1337 (O_1337,N_23907,N_24272);
or UO_1338 (O_1338,N_24487,N_23966);
and UO_1339 (O_1339,N_23843,N_24472);
xor UO_1340 (O_1340,N_24864,N_24907);
xor UO_1341 (O_1341,N_24253,N_24933);
and UO_1342 (O_1342,N_23984,N_24191);
nand UO_1343 (O_1343,N_24338,N_24705);
xnor UO_1344 (O_1344,N_24789,N_24182);
nand UO_1345 (O_1345,N_24377,N_24417);
xnor UO_1346 (O_1346,N_24155,N_23929);
or UO_1347 (O_1347,N_24217,N_24696);
nand UO_1348 (O_1348,N_24070,N_23935);
nand UO_1349 (O_1349,N_24919,N_24574);
and UO_1350 (O_1350,N_24727,N_24090);
xor UO_1351 (O_1351,N_24896,N_24350);
or UO_1352 (O_1352,N_24637,N_24329);
xnor UO_1353 (O_1353,N_24994,N_24839);
xor UO_1354 (O_1354,N_24658,N_24518);
nand UO_1355 (O_1355,N_24233,N_24990);
nand UO_1356 (O_1356,N_24184,N_24860);
xor UO_1357 (O_1357,N_24564,N_23882);
or UO_1358 (O_1358,N_24839,N_23993);
xnor UO_1359 (O_1359,N_23942,N_24410);
nor UO_1360 (O_1360,N_24373,N_24248);
nand UO_1361 (O_1361,N_24532,N_24991);
nor UO_1362 (O_1362,N_23827,N_24022);
and UO_1363 (O_1363,N_24202,N_24667);
nand UO_1364 (O_1364,N_24395,N_24516);
xor UO_1365 (O_1365,N_24940,N_23815);
and UO_1366 (O_1366,N_24087,N_24524);
and UO_1367 (O_1367,N_23915,N_24154);
and UO_1368 (O_1368,N_24363,N_24325);
or UO_1369 (O_1369,N_24955,N_24413);
nor UO_1370 (O_1370,N_24006,N_24765);
or UO_1371 (O_1371,N_24071,N_24385);
nor UO_1372 (O_1372,N_24352,N_24547);
nor UO_1373 (O_1373,N_24886,N_24268);
nand UO_1374 (O_1374,N_24010,N_23932);
and UO_1375 (O_1375,N_23878,N_24657);
or UO_1376 (O_1376,N_24440,N_24145);
and UO_1377 (O_1377,N_23864,N_24076);
nor UO_1378 (O_1378,N_24836,N_23845);
or UO_1379 (O_1379,N_24430,N_24795);
nor UO_1380 (O_1380,N_24945,N_24054);
and UO_1381 (O_1381,N_24727,N_24891);
nand UO_1382 (O_1382,N_24910,N_23883);
nor UO_1383 (O_1383,N_23777,N_23770);
nand UO_1384 (O_1384,N_23783,N_24483);
or UO_1385 (O_1385,N_24557,N_24343);
nand UO_1386 (O_1386,N_24895,N_24749);
nor UO_1387 (O_1387,N_24822,N_24601);
nor UO_1388 (O_1388,N_24619,N_24347);
or UO_1389 (O_1389,N_24836,N_24303);
nand UO_1390 (O_1390,N_23827,N_24523);
or UO_1391 (O_1391,N_24617,N_24240);
xor UO_1392 (O_1392,N_24283,N_24835);
and UO_1393 (O_1393,N_24343,N_23961);
xnor UO_1394 (O_1394,N_24724,N_24932);
xor UO_1395 (O_1395,N_24554,N_24191);
or UO_1396 (O_1396,N_24359,N_24656);
and UO_1397 (O_1397,N_24440,N_24545);
or UO_1398 (O_1398,N_24863,N_24262);
nor UO_1399 (O_1399,N_24949,N_24434);
nand UO_1400 (O_1400,N_24506,N_24639);
xnor UO_1401 (O_1401,N_24640,N_24771);
or UO_1402 (O_1402,N_24495,N_24970);
nor UO_1403 (O_1403,N_23918,N_24058);
nand UO_1404 (O_1404,N_24918,N_24411);
xnor UO_1405 (O_1405,N_24678,N_24025);
and UO_1406 (O_1406,N_24509,N_24156);
xor UO_1407 (O_1407,N_24998,N_24100);
and UO_1408 (O_1408,N_24528,N_24513);
nand UO_1409 (O_1409,N_23929,N_23827);
nor UO_1410 (O_1410,N_23964,N_23783);
or UO_1411 (O_1411,N_24049,N_24693);
nand UO_1412 (O_1412,N_24146,N_24977);
nor UO_1413 (O_1413,N_24122,N_24818);
and UO_1414 (O_1414,N_23800,N_23770);
or UO_1415 (O_1415,N_24110,N_24309);
or UO_1416 (O_1416,N_23786,N_24407);
xnor UO_1417 (O_1417,N_24594,N_24283);
nor UO_1418 (O_1418,N_24569,N_24548);
xor UO_1419 (O_1419,N_24152,N_24335);
and UO_1420 (O_1420,N_23936,N_23878);
xnor UO_1421 (O_1421,N_23884,N_24901);
xnor UO_1422 (O_1422,N_24503,N_24308);
and UO_1423 (O_1423,N_23753,N_24157);
nand UO_1424 (O_1424,N_24914,N_24709);
nor UO_1425 (O_1425,N_24121,N_24443);
and UO_1426 (O_1426,N_24887,N_24466);
nand UO_1427 (O_1427,N_24459,N_24002);
nor UO_1428 (O_1428,N_24233,N_23984);
and UO_1429 (O_1429,N_23931,N_24715);
and UO_1430 (O_1430,N_24914,N_24822);
nor UO_1431 (O_1431,N_24241,N_23891);
xnor UO_1432 (O_1432,N_23752,N_24053);
or UO_1433 (O_1433,N_23849,N_24025);
nand UO_1434 (O_1434,N_24587,N_24935);
nor UO_1435 (O_1435,N_24163,N_24520);
nand UO_1436 (O_1436,N_24626,N_24589);
and UO_1437 (O_1437,N_24397,N_24937);
nor UO_1438 (O_1438,N_24034,N_23870);
nand UO_1439 (O_1439,N_24088,N_24221);
nand UO_1440 (O_1440,N_24998,N_24708);
nor UO_1441 (O_1441,N_23882,N_24925);
nand UO_1442 (O_1442,N_23901,N_24997);
nand UO_1443 (O_1443,N_24923,N_23871);
and UO_1444 (O_1444,N_23938,N_24586);
nor UO_1445 (O_1445,N_24420,N_24978);
nor UO_1446 (O_1446,N_23788,N_24039);
xor UO_1447 (O_1447,N_24105,N_24778);
and UO_1448 (O_1448,N_24447,N_24322);
xor UO_1449 (O_1449,N_24770,N_23975);
xor UO_1450 (O_1450,N_24996,N_24806);
or UO_1451 (O_1451,N_23791,N_23990);
nor UO_1452 (O_1452,N_24133,N_24369);
or UO_1453 (O_1453,N_24479,N_23954);
nand UO_1454 (O_1454,N_24916,N_23996);
nand UO_1455 (O_1455,N_24162,N_24592);
xor UO_1456 (O_1456,N_24941,N_24894);
nand UO_1457 (O_1457,N_24881,N_24180);
and UO_1458 (O_1458,N_23896,N_24504);
nor UO_1459 (O_1459,N_24330,N_24352);
nor UO_1460 (O_1460,N_23932,N_24343);
nor UO_1461 (O_1461,N_24359,N_24798);
nor UO_1462 (O_1462,N_23993,N_24338);
nor UO_1463 (O_1463,N_24408,N_24193);
xnor UO_1464 (O_1464,N_24361,N_24358);
nand UO_1465 (O_1465,N_24111,N_24436);
nand UO_1466 (O_1466,N_24464,N_24106);
nor UO_1467 (O_1467,N_24758,N_23988);
and UO_1468 (O_1468,N_23797,N_23760);
nand UO_1469 (O_1469,N_24070,N_24319);
nor UO_1470 (O_1470,N_24999,N_24463);
xnor UO_1471 (O_1471,N_23992,N_24508);
nand UO_1472 (O_1472,N_23821,N_24711);
nand UO_1473 (O_1473,N_24795,N_24926);
xnor UO_1474 (O_1474,N_23802,N_23823);
nor UO_1475 (O_1475,N_23953,N_24686);
or UO_1476 (O_1476,N_24119,N_23759);
and UO_1477 (O_1477,N_23897,N_24660);
or UO_1478 (O_1478,N_24353,N_24607);
or UO_1479 (O_1479,N_24830,N_24373);
or UO_1480 (O_1480,N_23785,N_24623);
and UO_1481 (O_1481,N_24493,N_24727);
nand UO_1482 (O_1482,N_24333,N_24174);
xor UO_1483 (O_1483,N_24593,N_24587);
xnor UO_1484 (O_1484,N_24327,N_24354);
or UO_1485 (O_1485,N_24504,N_24865);
nand UO_1486 (O_1486,N_23751,N_24148);
nand UO_1487 (O_1487,N_24895,N_24299);
nand UO_1488 (O_1488,N_23928,N_24415);
nand UO_1489 (O_1489,N_23798,N_23784);
nor UO_1490 (O_1490,N_24004,N_24884);
xor UO_1491 (O_1491,N_24226,N_24105);
nor UO_1492 (O_1492,N_24725,N_24207);
xor UO_1493 (O_1493,N_24737,N_24828);
or UO_1494 (O_1494,N_24607,N_24284);
and UO_1495 (O_1495,N_23939,N_24281);
nand UO_1496 (O_1496,N_24944,N_24383);
xnor UO_1497 (O_1497,N_24559,N_24630);
nand UO_1498 (O_1498,N_24036,N_24383);
nand UO_1499 (O_1499,N_24235,N_23957);
xor UO_1500 (O_1500,N_24731,N_24879);
nand UO_1501 (O_1501,N_24669,N_24668);
nor UO_1502 (O_1502,N_24965,N_24798);
nor UO_1503 (O_1503,N_24458,N_24522);
nor UO_1504 (O_1504,N_24429,N_24030);
or UO_1505 (O_1505,N_23993,N_24052);
nor UO_1506 (O_1506,N_23908,N_24298);
nor UO_1507 (O_1507,N_24301,N_24463);
or UO_1508 (O_1508,N_23905,N_24284);
nand UO_1509 (O_1509,N_24318,N_24437);
xor UO_1510 (O_1510,N_24274,N_24083);
and UO_1511 (O_1511,N_24580,N_24236);
or UO_1512 (O_1512,N_24712,N_24745);
or UO_1513 (O_1513,N_24478,N_24726);
or UO_1514 (O_1514,N_24048,N_23985);
xnor UO_1515 (O_1515,N_24048,N_24067);
xor UO_1516 (O_1516,N_24324,N_24090);
xor UO_1517 (O_1517,N_24668,N_24968);
nor UO_1518 (O_1518,N_23851,N_23882);
and UO_1519 (O_1519,N_24498,N_24375);
and UO_1520 (O_1520,N_23877,N_23835);
and UO_1521 (O_1521,N_24498,N_24017);
or UO_1522 (O_1522,N_24061,N_24028);
or UO_1523 (O_1523,N_24139,N_24445);
nand UO_1524 (O_1524,N_24024,N_24103);
or UO_1525 (O_1525,N_23842,N_24923);
or UO_1526 (O_1526,N_23877,N_24049);
nor UO_1527 (O_1527,N_24954,N_24320);
nor UO_1528 (O_1528,N_24781,N_23979);
nor UO_1529 (O_1529,N_24599,N_24690);
nor UO_1530 (O_1530,N_24446,N_24174);
or UO_1531 (O_1531,N_23898,N_24834);
xor UO_1532 (O_1532,N_24318,N_24695);
nor UO_1533 (O_1533,N_24452,N_24234);
and UO_1534 (O_1534,N_24712,N_24259);
nor UO_1535 (O_1535,N_23924,N_24408);
or UO_1536 (O_1536,N_24309,N_24529);
or UO_1537 (O_1537,N_24472,N_24256);
nand UO_1538 (O_1538,N_24034,N_24272);
or UO_1539 (O_1539,N_24032,N_24897);
or UO_1540 (O_1540,N_24860,N_24687);
nand UO_1541 (O_1541,N_24896,N_24125);
nand UO_1542 (O_1542,N_24700,N_24072);
nor UO_1543 (O_1543,N_23810,N_23951);
xnor UO_1544 (O_1544,N_24459,N_24807);
nand UO_1545 (O_1545,N_24822,N_24957);
xnor UO_1546 (O_1546,N_24536,N_24602);
or UO_1547 (O_1547,N_24444,N_23835);
nand UO_1548 (O_1548,N_24693,N_23811);
or UO_1549 (O_1549,N_24733,N_24328);
nand UO_1550 (O_1550,N_24844,N_24478);
or UO_1551 (O_1551,N_24373,N_23817);
xnor UO_1552 (O_1552,N_24205,N_24891);
and UO_1553 (O_1553,N_24814,N_24052);
and UO_1554 (O_1554,N_24967,N_24255);
nor UO_1555 (O_1555,N_23873,N_24661);
nor UO_1556 (O_1556,N_23785,N_24210);
nand UO_1557 (O_1557,N_24681,N_24331);
xor UO_1558 (O_1558,N_24366,N_24607);
and UO_1559 (O_1559,N_24033,N_24224);
nand UO_1560 (O_1560,N_24431,N_24340);
or UO_1561 (O_1561,N_24779,N_24245);
or UO_1562 (O_1562,N_24182,N_23920);
or UO_1563 (O_1563,N_23866,N_24598);
or UO_1564 (O_1564,N_24388,N_24851);
nor UO_1565 (O_1565,N_24167,N_24495);
nor UO_1566 (O_1566,N_24660,N_24359);
nand UO_1567 (O_1567,N_23989,N_24691);
nor UO_1568 (O_1568,N_24372,N_23885);
nand UO_1569 (O_1569,N_24529,N_24810);
nor UO_1570 (O_1570,N_24221,N_24543);
or UO_1571 (O_1571,N_24980,N_24863);
nand UO_1572 (O_1572,N_24925,N_23861);
and UO_1573 (O_1573,N_24639,N_23793);
xnor UO_1574 (O_1574,N_24440,N_24438);
xnor UO_1575 (O_1575,N_24960,N_24487);
nor UO_1576 (O_1576,N_24617,N_24780);
nand UO_1577 (O_1577,N_23934,N_24140);
or UO_1578 (O_1578,N_24014,N_24969);
xor UO_1579 (O_1579,N_24078,N_23758);
nor UO_1580 (O_1580,N_24052,N_24500);
nand UO_1581 (O_1581,N_24317,N_24343);
or UO_1582 (O_1582,N_24833,N_24065);
xnor UO_1583 (O_1583,N_24824,N_24224);
nor UO_1584 (O_1584,N_23822,N_24583);
and UO_1585 (O_1585,N_24079,N_24635);
xor UO_1586 (O_1586,N_23894,N_24282);
nand UO_1587 (O_1587,N_24608,N_24886);
or UO_1588 (O_1588,N_23901,N_24507);
or UO_1589 (O_1589,N_24483,N_24355);
or UO_1590 (O_1590,N_24530,N_24985);
or UO_1591 (O_1591,N_24495,N_24676);
nor UO_1592 (O_1592,N_24985,N_24026);
or UO_1593 (O_1593,N_24247,N_24479);
or UO_1594 (O_1594,N_24418,N_24057);
xnor UO_1595 (O_1595,N_24612,N_24862);
and UO_1596 (O_1596,N_24494,N_24006);
and UO_1597 (O_1597,N_24797,N_24791);
nor UO_1598 (O_1598,N_23906,N_24885);
nand UO_1599 (O_1599,N_24498,N_24503);
nor UO_1600 (O_1600,N_24734,N_23878);
nor UO_1601 (O_1601,N_24820,N_23811);
nor UO_1602 (O_1602,N_24513,N_24645);
and UO_1603 (O_1603,N_23883,N_24812);
or UO_1604 (O_1604,N_24693,N_24343);
nor UO_1605 (O_1605,N_24599,N_23899);
xnor UO_1606 (O_1606,N_24563,N_24230);
nor UO_1607 (O_1607,N_24519,N_24146);
xor UO_1608 (O_1608,N_23776,N_24533);
nor UO_1609 (O_1609,N_23809,N_24323);
and UO_1610 (O_1610,N_24715,N_24738);
or UO_1611 (O_1611,N_24840,N_24469);
xor UO_1612 (O_1612,N_24684,N_23875);
nand UO_1613 (O_1613,N_24206,N_24648);
or UO_1614 (O_1614,N_23867,N_24887);
nand UO_1615 (O_1615,N_24148,N_24980);
or UO_1616 (O_1616,N_24423,N_23764);
and UO_1617 (O_1617,N_24684,N_23786);
nor UO_1618 (O_1618,N_24707,N_24438);
nor UO_1619 (O_1619,N_24951,N_24111);
xnor UO_1620 (O_1620,N_24747,N_24402);
nor UO_1621 (O_1621,N_23864,N_24261);
or UO_1622 (O_1622,N_24619,N_23991);
nor UO_1623 (O_1623,N_24133,N_23825);
xor UO_1624 (O_1624,N_24529,N_24532);
and UO_1625 (O_1625,N_24634,N_24689);
and UO_1626 (O_1626,N_23934,N_24395);
xnor UO_1627 (O_1627,N_24227,N_24517);
xor UO_1628 (O_1628,N_24164,N_24954);
or UO_1629 (O_1629,N_24627,N_24505);
nand UO_1630 (O_1630,N_24640,N_24452);
nand UO_1631 (O_1631,N_24978,N_24788);
or UO_1632 (O_1632,N_24216,N_24365);
or UO_1633 (O_1633,N_24065,N_23774);
nor UO_1634 (O_1634,N_24455,N_24429);
or UO_1635 (O_1635,N_23871,N_24347);
and UO_1636 (O_1636,N_24458,N_23822);
nand UO_1637 (O_1637,N_24925,N_24537);
and UO_1638 (O_1638,N_24898,N_24559);
nand UO_1639 (O_1639,N_24216,N_24146);
or UO_1640 (O_1640,N_24237,N_24683);
xor UO_1641 (O_1641,N_24123,N_23814);
nor UO_1642 (O_1642,N_24943,N_24151);
and UO_1643 (O_1643,N_24323,N_24176);
and UO_1644 (O_1644,N_24240,N_24421);
xnor UO_1645 (O_1645,N_24520,N_24645);
nand UO_1646 (O_1646,N_23853,N_24192);
nand UO_1647 (O_1647,N_24160,N_24791);
or UO_1648 (O_1648,N_23765,N_23933);
xor UO_1649 (O_1649,N_24493,N_24328);
nor UO_1650 (O_1650,N_24387,N_24417);
nor UO_1651 (O_1651,N_24867,N_24720);
nor UO_1652 (O_1652,N_23778,N_24364);
or UO_1653 (O_1653,N_23762,N_24100);
or UO_1654 (O_1654,N_24041,N_24318);
nor UO_1655 (O_1655,N_23892,N_24946);
and UO_1656 (O_1656,N_23993,N_24898);
nor UO_1657 (O_1657,N_24594,N_24524);
xor UO_1658 (O_1658,N_24440,N_23883);
nor UO_1659 (O_1659,N_24973,N_24652);
and UO_1660 (O_1660,N_24703,N_24589);
nand UO_1661 (O_1661,N_23807,N_23827);
nor UO_1662 (O_1662,N_24387,N_24384);
and UO_1663 (O_1663,N_24623,N_24358);
nand UO_1664 (O_1664,N_23952,N_24968);
xor UO_1665 (O_1665,N_24577,N_24876);
xor UO_1666 (O_1666,N_23788,N_23774);
or UO_1667 (O_1667,N_24980,N_24969);
and UO_1668 (O_1668,N_24633,N_23985);
nor UO_1669 (O_1669,N_23867,N_24498);
nor UO_1670 (O_1670,N_24432,N_24463);
xnor UO_1671 (O_1671,N_24148,N_24769);
nor UO_1672 (O_1672,N_24480,N_24605);
nor UO_1673 (O_1673,N_24754,N_24608);
or UO_1674 (O_1674,N_24826,N_24067);
and UO_1675 (O_1675,N_24595,N_23752);
or UO_1676 (O_1676,N_24519,N_24558);
or UO_1677 (O_1677,N_23982,N_24982);
nand UO_1678 (O_1678,N_24319,N_23878);
and UO_1679 (O_1679,N_24805,N_24845);
nor UO_1680 (O_1680,N_24827,N_23874);
xor UO_1681 (O_1681,N_24083,N_24945);
nor UO_1682 (O_1682,N_24193,N_23996);
nand UO_1683 (O_1683,N_24756,N_24305);
and UO_1684 (O_1684,N_24666,N_24575);
xnor UO_1685 (O_1685,N_23871,N_24460);
nand UO_1686 (O_1686,N_23777,N_23842);
nand UO_1687 (O_1687,N_24203,N_24941);
nor UO_1688 (O_1688,N_24246,N_24055);
xor UO_1689 (O_1689,N_23808,N_24263);
or UO_1690 (O_1690,N_24496,N_24923);
and UO_1691 (O_1691,N_24989,N_24217);
xor UO_1692 (O_1692,N_24424,N_24399);
and UO_1693 (O_1693,N_24026,N_24369);
or UO_1694 (O_1694,N_24491,N_24242);
or UO_1695 (O_1695,N_24598,N_24422);
or UO_1696 (O_1696,N_24699,N_24306);
xor UO_1697 (O_1697,N_24535,N_24954);
or UO_1698 (O_1698,N_24666,N_24639);
nand UO_1699 (O_1699,N_23850,N_23787);
nor UO_1700 (O_1700,N_24222,N_24994);
nor UO_1701 (O_1701,N_24366,N_24165);
nor UO_1702 (O_1702,N_23785,N_24523);
or UO_1703 (O_1703,N_24326,N_24493);
or UO_1704 (O_1704,N_24127,N_23839);
nor UO_1705 (O_1705,N_24012,N_24030);
nand UO_1706 (O_1706,N_24086,N_24642);
nand UO_1707 (O_1707,N_24790,N_24569);
nor UO_1708 (O_1708,N_24754,N_24610);
xnor UO_1709 (O_1709,N_23815,N_24716);
nand UO_1710 (O_1710,N_24064,N_23971);
or UO_1711 (O_1711,N_23861,N_24112);
xnor UO_1712 (O_1712,N_24078,N_24409);
xnor UO_1713 (O_1713,N_23843,N_23839);
or UO_1714 (O_1714,N_23814,N_24665);
nand UO_1715 (O_1715,N_24520,N_24798);
nand UO_1716 (O_1716,N_24563,N_24313);
and UO_1717 (O_1717,N_24585,N_24679);
nor UO_1718 (O_1718,N_23840,N_24777);
nand UO_1719 (O_1719,N_24471,N_23911);
nor UO_1720 (O_1720,N_23901,N_24674);
and UO_1721 (O_1721,N_24231,N_24779);
nor UO_1722 (O_1722,N_24494,N_24256);
nand UO_1723 (O_1723,N_24384,N_23809);
xnor UO_1724 (O_1724,N_23948,N_23779);
nor UO_1725 (O_1725,N_24277,N_24970);
or UO_1726 (O_1726,N_24210,N_24369);
or UO_1727 (O_1727,N_24762,N_24368);
or UO_1728 (O_1728,N_24052,N_23926);
nor UO_1729 (O_1729,N_24248,N_23941);
nand UO_1730 (O_1730,N_23761,N_24217);
or UO_1731 (O_1731,N_24988,N_24443);
nor UO_1732 (O_1732,N_23906,N_24225);
nand UO_1733 (O_1733,N_24278,N_23827);
or UO_1734 (O_1734,N_24415,N_24503);
nor UO_1735 (O_1735,N_23946,N_24393);
nor UO_1736 (O_1736,N_24321,N_24333);
xor UO_1737 (O_1737,N_24845,N_24768);
xnor UO_1738 (O_1738,N_24748,N_24305);
or UO_1739 (O_1739,N_23839,N_24600);
nand UO_1740 (O_1740,N_24070,N_23887);
nand UO_1741 (O_1741,N_24923,N_24992);
or UO_1742 (O_1742,N_24531,N_24069);
or UO_1743 (O_1743,N_24995,N_24423);
and UO_1744 (O_1744,N_24809,N_24378);
nor UO_1745 (O_1745,N_23930,N_23944);
and UO_1746 (O_1746,N_24749,N_24386);
nor UO_1747 (O_1747,N_24513,N_23768);
or UO_1748 (O_1748,N_24060,N_24837);
nor UO_1749 (O_1749,N_24714,N_24550);
and UO_1750 (O_1750,N_23999,N_24958);
nor UO_1751 (O_1751,N_24839,N_24421);
nor UO_1752 (O_1752,N_24854,N_24387);
and UO_1753 (O_1753,N_24743,N_24343);
nand UO_1754 (O_1754,N_24966,N_24272);
or UO_1755 (O_1755,N_23916,N_23914);
or UO_1756 (O_1756,N_24434,N_24296);
nor UO_1757 (O_1757,N_23963,N_24094);
or UO_1758 (O_1758,N_24313,N_24959);
xor UO_1759 (O_1759,N_24031,N_24621);
nand UO_1760 (O_1760,N_24521,N_24641);
and UO_1761 (O_1761,N_24519,N_24598);
nor UO_1762 (O_1762,N_24440,N_23920);
nor UO_1763 (O_1763,N_24126,N_23912);
or UO_1764 (O_1764,N_24396,N_24240);
and UO_1765 (O_1765,N_24250,N_24792);
nor UO_1766 (O_1766,N_24268,N_24224);
nand UO_1767 (O_1767,N_24012,N_24394);
and UO_1768 (O_1768,N_24534,N_24177);
nor UO_1769 (O_1769,N_23890,N_24706);
and UO_1770 (O_1770,N_24986,N_24391);
xnor UO_1771 (O_1771,N_24311,N_24282);
or UO_1772 (O_1772,N_24966,N_24051);
nor UO_1773 (O_1773,N_24105,N_24839);
xor UO_1774 (O_1774,N_24455,N_24839);
or UO_1775 (O_1775,N_24673,N_24996);
xor UO_1776 (O_1776,N_24059,N_23787);
nor UO_1777 (O_1777,N_24021,N_24757);
nor UO_1778 (O_1778,N_24674,N_24021);
or UO_1779 (O_1779,N_23786,N_23770);
and UO_1780 (O_1780,N_24923,N_24192);
nor UO_1781 (O_1781,N_24468,N_24294);
or UO_1782 (O_1782,N_24557,N_24202);
or UO_1783 (O_1783,N_24248,N_24448);
xor UO_1784 (O_1784,N_23895,N_23971);
xnor UO_1785 (O_1785,N_24153,N_24724);
nor UO_1786 (O_1786,N_24376,N_24133);
nor UO_1787 (O_1787,N_24352,N_24436);
nand UO_1788 (O_1788,N_24518,N_23926);
or UO_1789 (O_1789,N_24865,N_24166);
xor UO_1790 (O_1790,N_24312,N_23853);
or UO_1791 (O_1791,N_24011,N_23992);
and UO_1792 (O_1792,N_24161,N_24777);
or UO_1793 (O_1793,N_24941,N_24642);
or UO_1794 (O_1794,N_24838,N_24744);
xor UO_1795 (O_1795,N_24663,N_24166);
nor UO_1796 (O_1796,N_24608,N_24310);
nor UO_1797 (O_1797,N_24749,N_24087);
and UO_1798 (O_1798,N_24629,N_24637);
or UO_1799 (O_1799,N_24028,N_24008);
nor UO_1800 (O_1800,N_24592,N_23912);
and UO_1801 (O_1801,N_24281,N_24761);
nor UO_1802 (O_1802,N_24104,N_24768);
or UO_1803 (O_1803,N_24590,N_24396);
xnor UO_1804 (O_1804,N_24856,N_24000);
xnor UO_1805 (O_1805,N_23806,N_24081);
or UO_1806 (O_1806,N_23995,N_23884);
nor UO_1807 (O_1807,N_24112,N_24110);
or UO_1808 (O_1808,N_24213,N_24242);
or UO_1809 (O_1809,N_23805,N_24772);
nand UO_1810 (O_1810,N_24792,N_24618);
nand UO_1811 (O_1811,N_24471,N_24312);
and UO_1812 (O_1812,N_23896,N_24042);
nor UO_1813 (O_1813,N_24198,N_24778);
nand UO_1814 (O_1814,N_24800,N_23791);
and UO_1815 (O_1815,N_24891,N_24547);
xor UO_1816 (O_1816,N_24463,N_23829);
or UO_1817 (O_1817,N_23761,N_24995);
nand UO_1818 (O_1818,N_24442,N_24007);
nand UO_1819 (O_1819,N_24391,N_24409);
nor UO_1820 (O_1820,N_24046,N_24638);
or UO_1821 (O_1821,N_24244,N_24018);
nor UO_1822 (O_1822,N_24799,N_24640);
and UO_1823 (O_1823,N_24170,N_24202);
xor UO_1824 (O_1824,N_24818,N_23870);
or UO_1825 (O_1825,N_24390,N_24016);
xor UO_1826 (O_1826,N_24466,N_24858);
nor UO_1827 (O_1827,N_24271,N_24698);
xor UO_1828 (O_1828,N_23963,N_24348);
nor UO_1829 (O_1829,N_23895,N_24063);
and UO_1830 (O_1830,N_23771,N_24990);
xor UO_1831 (O_1831,N_24143,N_24065);
and UO_1832 (O_1832,N_23806,N_24411);
nand UO_1833 (O_1833,N_23877,N_23992);
or UO_1834 (O_1834,N_24024,N_23889);
xor UO_1835 (O_1835,N_24115,N_24694);
or UO_1836 (O_1836,N_23927,N_24642);
or UO_1837 (O_1837,N_24757,N_24744);
nor UO_1838 (O_1838,N_24102,N_24055);
xor UO_1839 (O_1839,N_24744,N_23803);
nor UO_1840 (O_1840,N_24705,N_24260);
xnor UO_1841 (O_1841,N_24737,N_24586);
and UO_1842 (O_1842,N_24645,N_24611);
xnor UO_1843 (O_1843,N_23859,N_24857);
nor UO_1844 (O_1844,N_24179,N_24133);
and UO_1845 (O_1845,N_24920,N_23936);
and UO_1846 (O_1846,N_24848,N_23774);
nor UO_1847 (O_1847,N_24335,N_24190);
or UO_1848 (O_1848,N_23908,N_24281);
or UO_1849 (O_1849,N_23836,N_23837);
and UO_1850 (O_1850,N_24877,N_23820);
and UO_1851 (O_1851,N_24114,N_24326);
or UO_1852 (O_1852,N_24910,N_24876);
nand UO_1853 (O_1853,N_24650,N_24058);
nor UO_1854 (O_1854,N_24186,N_24088);
and UO_1855 (O_1855,N_24592,N_23957);
nor UO_1856 (O_1856,N_24808,N_23868);
nand UO_1857 (O_1857,N_24557,N_23910);
and UO_1858 (O_1858,N_24314,N_24322);
and UO_1859 (O_1859,N_24844,N_24434);
nor UO_1860 (O_1860,N_24418,N_24307);
xor UO_1861 (O_1861,N_24845,N_23994);
or UO_1862 (O_1862,N_24493,N_24741);
nand UO_1863 (O_1863,N_24220,N_24882);
and UO_1864 (O_1864,N_24058,N_24159);
and UO_1865 (O_1865,N_24237,N_24053);
xnor UO_1866 (O_1866,N_24157,N_24719);
nand UO_1867 (O_1867,N_23861,N_24921);
nor UO_1868 (O_1868,N_24333,N_24082);
nand UO_1869 (O_1869,N_24204,N_24854);
nor UO_1870 (O_1870,N_24145,N_24121);
nor UO_1871 (O_1871,N_24082,N_24668);
xnor UO_1872 (O_1872,N_24621,N_23905);
nor UO_1873 (O_1873,N_24021,N_23794);
nand UO_1874 (O_1874,N_24978,N_24876);
xor UO_1875 (O_1875,N_23871,N_24093);
nand UO_1876 (O_1876,N_24241,N_24134);
or UO_1877 (O_1877,N_23932,N_24961);
and UO_1878 (O_1878,N_24013,N_23893);
nor UO_1879 (O_1879,N_24205,N_24978);
xor UO_1880 (O_1880,N_24463,N_24923);
or UO_1881 (O_1881,N_24261,N_24003);
and UO_1882 (O_1882,N_24209,N_24530);
nor UO_1883 (O_1883,N_24507,N_23970);
xor UO_1884 (O_1884,N_24443,N_23913);
or UO_1885 (O_1885,N_24670,N_24567);
and UO_1886 (O_1886,N_24277,N_24935);
or UO_1887 (O_1887,N_24660,N_23901);
nor UO_1888 (O_1888,N_24025,N_24633);
xor UO_1889 (O_1889,N_24967,N_24846);
nand UO_1890 (O_1890,N_23956,N_24801);
or UO_1891 (O_1891,N_24116,N_24245);
xnor UO_1892 (O_1892,N_24137,N_24667);
or UO_1893 (O_1893,N_24080,N_24963);
xor UO_1894 (O_1894,N_24059,N_24956);
nand UO_1895 (O_1895,N_24984,N_24535);
xor UO_1896 (O_1896,N_23766,N_23834);
nor UO_1897 (O_1897,N_23895,N_24311);
nor UO_1898 (O_1898,N_24336,N_24031);
and UO_1899 (O_1899,N_24484,N_24558);
xnor UO_1900 (O_1900,N_24661,N_24331);
nand UO_1901 (O_1901,N_24942,N_24415);
xor UO_1902 (O_1902,N_24100,N_24449);
and UO_1903 (O_1903,N_23926,N_24564);
nor UO_1904 (O_1904,N_24178,N_24687);
and UO_1905 (O_1905,N_24115,N_24712);
nor UO_1906 (O_1906,N_24868,N_24179);
and UO_1907 (O_1907,N_24631,N_24175);
or UO_1908 (O_1908,N_24293,N_24479);
xnor UO_1909 (O_1909,N_23796,N_24778);
or UO_1910 (O_1910,N_24835,N_23890);
xor UO_1911 (O_1911,N_23860,N_24660);
nor UO_1912 (O_1912,N_24103,N_24142);
nor UO_1913 (O_1913,N_24718,N_24727);
and UO_1914 (O_1914,N_23817,N_24997);
nor UO_1915 (O_1915,N_23835,N_24866);
or UO_1916 (O_1916,N_24117,N_24601);
or UO_1917 (O_1917,N_24913,N_24416);
xor UO_1918 (O_1918,N_23850,N_23835);
xor UO_1919 (O_1919,N_24045,N_23832);
nor UO_1920 (O_1920,N_24300,N_24610);
and UO_1921 (O_1921,N_24520,N_23900);
nand UO_1922 (O_1922,N_24751,N_24942);
xnor UO_1923 (O_1923,N_24918,N_24132);
nor UO_1924 (O_1924,N_23887,N_24190);
nor UO_1925 (O_1925,N_24573,N_24315);
nor UO_1926 (O_1926,N_24871,N_24025);
xnor UO_1927 (O_1927,N_24626,N_24439);
xor UO_1928 (O_1928,N_24459,N_24826);
nor UO_1929 (O_1929,N_23935,N_23755);
xor UO_1930 (O_1930,N_24014,N_24070);
and UO_1931 (O_1931,N_24436,N_24204);
xnor UO_1932 (O_1932,N_24512,N_24327);
and UO_1933 (O_1933,N_24433,N_24655);
xor UO_1934 (O_1934,N_24736,N_23921);
xor UO_1935 (O_1935,N_24501,N_23954);
and UO_1936 (O_1936,N_24783,N_24920);
or UO_1937 (O_1937,N_24913,N_23928);
xor UO_1938 (O_1938,N_24439,N_24932);
nor UO_1939 (O_1939,N_24952,N_24163);
and UO_1940 (O_1940,N_24496,N_24916);
or UO_1941 (O_1941,N_23868,N_24897);
xnor UO_1942 (O_1942,N_23776,N_24956);
and UO_1943 (O_1943,N_24526,N_24913);
or UO_1944 (O_1944,N_24902,N_24284);
nand UO_1945 (O_1945,N_24648,N_24537);
nor UO_1946 (O_1946,N_23782,N_24248);
xor UO_1947 (O_1947,N_24021,N_24922);
nand UO_1948 (O_1948,N_24831,N_24673);
xor UO_1949 (O_1949,N_24488,N_23889);
and UO_1950 (O_1950,N_24004,N_24401);
xnor UO_1951 (O_1951,N_24999,N_23835);
and UO_1952 (O_1952,N_24710,N_24354);
xnor UO_1953 (O_1953,N_24026,N_24183);
or UO_1954 (O_1954,N_24299,N_23903);
nand UO_1955 (O_1955,N_24896,N_24606);
or UO_1956 (O_1956,N_24057,N_23845);
and UO_1957 (O_1957,N_24945,N_24781);
or UO_1958 (O_1958,N_24148,N_24697);
nand UO_1959 (O_1959,N_24718,N_23954);
nand UO_1960 (O_1960,N_24251,N_24591);
xnor UO_1961 (O_1961,N_23808,N_24378);
nor UO_1962 (O_1962,N_24255,N_24262);
nor UO_1963 (O_1963,N_23810,N_24752);
nand UO_1964 (O_1964,N_24045,N_24705);
nand UO_1965 (O_1965,N_23797,N_23753);
and UO_1966 (O_1966,N_24459,N_23760);
nor UO_1967 (O_1967,N_23913,N_24034);
nand UO_1968 (O_1968,N_24446,N_23820);
xor UO_1969 (O_1969,N_24451,N_24465);
nor UO_1970 (O_1970,N_23870,N_23880);
or UO_1971 (O_1971,N_24172,N_24586);
xor UO_1972 (O_1972,N_24556,N_24618);
and UO_1973 (O_1973,N_24012,N_23993);
nor UO_1974 (O_1974,N_24824,N_24326);
or UO_1975 (O_1975,N_23899,N_24172);
and UO_1976 (O_1976,N_24217,N_24211);
xnor UO_1977 (O_1977,N_24116,N_24814);
and UO_1978 (O_1978,N_24570,N_24224);
xor UO_1979 (O_1979,N_23920,N_24938);
xnor UO_1980 (O_1980,N_24536,N_23936);
xor UO_1981 (O_1981,N_24333,N_24263);
and UO_1982 (O_1982,N_23914,N_23770);
or UO_1983 (O_1983,N_24002,N_23949);
and UO_1984 (O_1984,N_24846,N_24955);
and UO_1985 (O_1985,N_24916,N_24874);
xor UO_1986 (O_1986,N_23952,N_24234);
and UO_1987 (O_1987,N_24855,N_24760);
xor UO_1988 (O_1988,N_24838,N_24049);
and UO_1989 (O_1989,N_24777,N_23996);
nand UO_1990 (O_1990,N_23879,N_24519);
and UO_1991 (O_1991,N_24705,N_24397);
nor UO_1992 (O_1992,N_24543,N_24004);
nor UO_1993 (O_1993,N_24294,N_24752);
and UO_1994 (O_1994,N_24337,N_24816);
nor UO_1995 (O_1995,N_23930,N_24511);
nand UO_1996 (O_1996,N_24579,N_24380);
xnor UO_1997 (O_1997,N_24795,N_24661);
and UO_1998 (O_1998,N_24874,N_24917);
nor UO_1999 (O_1999,N_24617,N_23834);
xnor UO_2000 (O_2000,N_24000,N_24323);
nor UO_2001 (O_2001,N_24185,N_24173);
nand UO_2002 (O_2002,N_24705,N_24467);
or UO_2003 (O_2003,N_24201,N_24940);
nand UO_2004 (O_2004,N_23865,N_24461);
xnor UO_2005 (O_2005,N_23920,N_24962);
or UO_2006 (O_2006,N_23803,N_24555);
nand UO_2007 (O_2007,N_24170,N_24534);
and UO_2008 (O_2008,N_24279,N_24483);
and UO_2009 (O_2009,N_24304,N_24004);
or UO_2010 (O_2010,N_24882,N_24977);
or UO_2011 (O_2011,N_24744,N_24283);
nand UO_2012 (O_2012,N_24075,N_24182);
nand UO_2013 (O_2013,N_24690,N_24662);
or UO_2014 (O_2014,N_23850,N_24678);
xnor UO_2015 (O_2015,N_24008,N_24157);
nand UO_2016 (O_2016,N_24526,N_24905);
and UO_2017 (O_2017,N_24514,N_24084);
nor UO_2018 (O_2018,N_23912,N_24029);
nand UO_2019 (O_2019,N_24755,N_23836);
xor UO_2020 (O_2020,N_24676,N_24521);
nand UO_2021 (O_2021,N_24508,N_24191);
nor UO_2022 (O_2022,N_24945,N_24544);
nor UO_2023 (O_2023,N_24563,N_24639);
nor UO_2024 (O_2024,N_24969,N_24620);
nand UO_2025 (O_2025,N_23834,N_24088);
nor UO_2026 (O_2026,N_24840,N_24093);
or UO_2027 (O_2027,N_24643,N_24614);
xnor UO_2028 (O_2028,N_24115,N_24222);
nand UO_2029 (O_2029,N_24815,N_24884);
nor UO_2030 (O_2030,N_24435,N_24273);
nor UO_2031 (O_2031,N_24725,N_24474);
or UO_2032 (O_2032,N_24365,N_24149);
and UO_2033 (O_2033,N_24546,N_23889);
xnor UO_2034 (O_2034,N_24351,N_24084);
nor UO_2035 (O_2035,N_24090,N_24017);
nand UO_2036 (O_2036,N_24855,N_24627);
xor UO_2037 (O_2037,N_24261,N_24495);
and UO_2038 (O_2038,N_24019,N_24096);
and UO_2039 (O_2039,N_24237,N_24374);
nand UO_2040 (O_2040,N_24998,N_24845);
and UO_2041 (O_2041,N_24642,N_24752);
xor UO_2042 (O_2042,N_24267,N_24219);
and UO_2043 (O_2043,N_24952,N_23907);
and UO_2044 (O_2044,N_24298,N_23917);
nor UO_2045 (O_2045,N_24511,N_23885);
nor UO_2046 (O_2046,N_24140,N_24228);
nor UO_2047 (O_2047,N_24782,N_24963);
nand UO_2048 (O_2048,N_24231,N_24409);
nand UO_2049 (O_2049,N_24983,N_23873);
or UO_2050 (O_2050,N_24121,N_23908);
xor UO_2051 (O_2051,N_23879,N_24389);
and UO_2052 (O_2052,N_24489,N_24305);
xor UO_2053 (O_2053,N_24982,N_24396);
nor UO_2054 (O_2054,N_23795,N_24212);
xnor UO_2055 (O_2055,N_24320,N_24417);
nor UO_2056 (O_2056,N_24425,N_24156);
or UO_2057 (O_2057,N_23929,N_23812);
nand UO_2058 (O_2058,N_24435,N_24915);
nand UO_2059 (O_2059,N_24686,N_24653);
nand UO_2060 (O_2060,N_24727,N_24712);
and UO_2061 (O_2061,N_24295,N_24808);
nor UO_2062 (O_2062,N_24969,N_24690);
or UO_2063 (O_2063,N_24202,N_23760);
and UO_2064 (O_2064,N_23831,N_24532);
nand UO_2065 (O_2065,N_24925,N_24604);
nor UO_2066 (O_2066,N_24852,N_23837);
xor UO_2067 (O_2067,N_24111,N_24527);
nand UO_2068 (O_2068,N_24860,N_24895);
nand UO_2069 (O_2069,N_24007,N_24290);
xnor UO_2070 (O_2070,N_24755,N_24841);
or UO_2071 (O_2071,N_24987,N_24280);
xor UO_2072 (O_2072,N_23912,N_24897);
nor UO_2073 (O_2073,N_24095,N_24375);
nand UO_2074 (O_2074,N_24005,N_24665);
and UO_2075 (O_2075,N_24334,N_23839);
xnor UO_2076 (O_2076,N_24246,N_24222);
or UO_2077 (O_2077,N_24836,N_24508);
nand UO_2078 (O_2078,N_23987,N_24957);
xnor UO_2079 (O_2079,N_24946,N_24131);
or UO_2080 (O_2080,N_24380,N_23817);
nor UO_2081 (O_2081,N_24100,N_24332);
and UO_2082 (O_2082,N_24949,N_24040);
nand UO_2083 (O_2083,N_24099,N_24838);
xnor UO_2084 (O_2084,N_23819,N_24447);
nor UO_2085 (O_2085,N_24302,N_24282);
and UO_2086 (O_2086,N_24638,N_24784);
nor UO_2087 (O_2087,N_24257,N_24636);
nor UO_2088 (O_2088,N_24771,N_23815);
nand UO_2089 (O_2089,N_24465,N_24911);
or UO_2090 (O_2090,N_24153,N_24176);
xor UO_2091 (O_2091,N_23752,N_24101);
xnor UO_2092 (O_2092,N_24143,N_24807);
nand UO_2093 (O_2093,N_24283,N_24002);
xor UO_2094 (O_2094,N_24423,N_24548);
xor UO_2095 (O_2095,N_24242,N_23994);
xor UO_2096 (O_2096,N_24335,N_24078);
nand UO_2097 (O_2097,N_24995,N_23769);
nor UO_2098 (O_2098,N_24948,N_24982);
xnor UO_2099 (O_2099,N_24133,N_24778);
nand UO_2100 (O_2100,N_24343,N_24941);
or UO_2101 (O_2101,N_23949,N_24702);
nor UO_2102 (O_2102,N_24403,N_24967);
or UO_2103 (O_2103,N_24105,N_24283);
xnor UO_2104 (O_2104,N_23876,N_24281);
and UO_2105 (O_2105,N_23947,N_23883);
and UO_2106 (O_2106,N_24256,N_24848);
nor UO_2107 (O_2107,N_24229,N_23785);
and UO_2108 (O_2108,N_23910,N_24259);
or UO_2109 (O_2109,N_24869,N_24977);
nor UO_2110 (O_2110,N_24336,N_23898);
or UO_2111 (O_2111,N_24534,N_23861);
or UO_2112 (O_2112,N_24984,N_24808);
xnor UO_2113 (O_2113,N_23849,N_24585);
or UO_2114 (O_2114,N_24961,N_23893);
xnor UO_2115 (O_2115,N_23988,N_24631);
xnor UO_2116 (O_2116,N_24532,N_24110);
and UO_2117 (O_2117,N_24615,N_24454);
or UO_2118 (O_2118,N_24646,N_24494);
or UO_2119 (O_2119,N_24993,N_24608);
xnor UO_2120 (O_2120,N_24335,N_23769);
nand UO_2121 (O_2121,N_24653,N_24441);
and UO_2122 (O_2122,N_23804,N_24265);
and UO_2123 (O_2123,N_24250,N_24806);
nor UO_2124 (O_2124,N_24972,N_24775);
and UO_2125 (O_2125,N_24600,N_23771);
or UO_2126 (O_2126,N_24530,N_23824);
or UO_2127 (O_2127,N_24280,N_24588);
nor UO_2128 (O_2128,N_24915,N_23765);
xnor UO_2129 (O_2129,N_24413,N_24811);
nand UO_2130 (O_2130,N_24919,N_24269);
xnor UO_2131 (O_2131,N_24154,N_24591);
xor UO_2132 (O_2132,N_24965,N_24870);
and UO_2133 (O_2133,N_24779,N_24441);
and UO_2134 (O_2134,N_23893,N_23927);
and UO_2135 (O_2135,N_24804,N_23984);
and UO_2136 (O_2136,N_24698,N_24552);
nand UO_2137 (O_2137,N_24423,N_24279);
xor UO_2138 (O_2138,N_24985,N_24462);
nor UO_2139 (O_2139,N_24486,N_24426);
nor UO_2140 (O_2140,N_24100,N_24518);
nor UO_2141 (O_2141,N_24015,N_24843);
nand UO_2142 (O_2142,N_23783,N_23961);
or UO_2143 (O_2143,N_23819,N_23817);
nor UO_2144 (O_2144,N_24536,N_24598);
nand UO_2145 (O_2145,N_24694,N_24763);
nor UO_2146 (O_2146,N_24266,N_24605);
or UO_2147 (O_2147,N_23853,N_24945);
xnor UO_2148 (O_2148,N_23765,N_24796);
nand UO_2149 (O_2149,N_24915,N_24645);
or UO_2150 (O_2150,N_24610,N_24144);
nor UO_2151 (O_2151,N_24125,N_23935);
or UO_2152 (O_2152,N_23933,N_23780);
xnor UO_2153 (O_2153,N_23839,N_24398);
and UO_2154 (O_2154,N_24368,N_24404);
nor UO_2155 (O_2155,N_24717,N_24985);
and UO_2156 (O_2156,N_24542,N_24634);
xor UO_2157 (O_2157,N_24600,N_24108);
xnor UO_2158 (O_2158,N_24046,N_24282);
nand UO_2159 (O_2159,N_24247,N_24698);
xor UO_2160 (O_2160,N_24218,N_24952);
xor UO_2161 (O_2161,N_24932,N_24990);
and UO_2162 (O_2162,N_24235,N_24191);
nand UO_2163 (O_2163,N_24331,N_24826);
or UO_2164 (O_2164,N_24447,N_24358);
or UO_2165 (O_2165,N_24552,N_23993);
xnor UO_2166 (O_2166,N_24743,N_24822);
nand UO_2167 (O_2167,N_24839,N_24774);
xor UO_2168 (O_2168,N_24063,N_24784);
and UO_2169 (O_2169,N_23832,N_23917);
nand UO_2170 (O_2170,N_24630,N_24354);
or UO_2171 (O_2171,N_23875,N_24241);
nor UO_2172 (O_2172,N_24067,N_24120);
nand UO_2173 (O_2173,N_24914,N_24263);
nand UO_2174 (O_2174,N_24241,N_23969);
nand UO_2175 (O_2175,N_24619,N_24968);
nor UO_2176 (O_2176,N_24648,N_24928);
nand UO_2177 (O_2177,N_24308,N_24004);
xor UO_2178 (O_2178,N_24096,N_24471);
nand UO_2179 (O_2179,N_24499,N_23779);
xnor UO_2180 (O_2180,N_24537,N_23990);
xnor UO_2181 (O_2181,N_24409,N_24925);
nor UO_2182 (O_2182,N_23958,N_24979);
nor UO_2183 (O_2183,N_23865,N_24676);
nor UO_2184 (O_2184,N_24566,N_24144);
or UO_2185 (O_2185,N_24574,N_24994);
nor UO_2186 (O_2186,N_24965,N_24056);
xnor UO_2187 (O_2187,N_24462,N_24722);
and UO_2188 (O_2188,N_24537,N_24424);
nor UO_2189 (O_2189,N_24425,N_24796);
and UO_2190 (O_2190,N_24690,N_24178);
or UO_2191 (O_2191,N_23991,N_24792);
nand UO_2192 (O_2192,N_24157,N_23878);
or UO_2193 (O_2193,N_24989,N_24853);
or UO_2194 (O_2194,N_24069,N_24883);
and UO_2195 (O_2195,N_24356,N_24878);
and UO_2196 (O_2196,N_24157,N_24018);
nand UO_2197 (O_2197,N_23782,N_24794);
nand UO_2198 (O_2198,N_24975,N_23949);
and UO_2199 (O_2199,N_24727,N_23811);
and UO_2200 (O_2200,N_24985,N_23914);
xnor UO_2201 (O_2201,N_24332,N_24319);
nand UO_2202 (O_2202,N_23833,N_24957);
xnor UO_2203 (O_2203,N_24905,N_24748);
nor UO_2204 (O_2204,N_24578,N_23944);
xor UO_2205 (O_2205,N_24473,N_24346);
nand UO_2206 (O_2206,N_24282,N_24266);
or UO_2207 (O_2207,N_24453,N_24811);
xor UO_2208 (O_2208,N_24135,N_24953);
nor UO_2209 (O_2209,N_24437,N_24265);
or UO_2210 (O_2210,N_24975,N_24350);
nor UO_2211 (O_2211,N_24279,N_24249);
or UO_2212 (O_2212,N_23981,N_24936);
or UO_2213 (O_2213,N_23772,N_23936);
or UO_2214 (O_2214,N_24958,N_24799);
nor UO_2215 (O_2215,N_23761,N_23782);
nor UO_2216 (O_2216,N_24983,N_24894);
nor UO_2217 (O_2217,N_24585,N_24852);
or UO_2218 (O_2218,N_24418,N_23770);
or UO_2219 (O_2219,N_24993,N_24890);
xnor UO_2220 (O_2220,N_24288,N_24335);
xor UO_2221 (O_2221,N_24232,N_24514);
nand UO_2222 (O_2222,N_24410,N_24171);
or UO_2223 (O_2223,N_24677,N_24679);
or UO_2224 (O_2224,N_23825,N_24442);
and UO_2225 (O_2225,N_23776,N_24906);
nand UO_2226 (O_2226,N_24745,N_24603);
and UO_2227 (O_2227,N_24462,N_24596);
or UO_2228 (O_2228,N_24007,N_23903);
and UO_2229 (O_2229,N_23842,N_24536);
nor UO_2230 (O_2230,N_24926,N_23956);
and UO_2231 (O_2231,N_24603,N_24086);
or UO_2232 (O_2232,N_24521,N_23811);
nor UO_2233 (O_2233,N_24958,N_24484);
or UO_2234 (O_2234,N_23851,N_24892);
or UO_2235 (O_2235,N_24537,N_24541);
nor UO_2236 (O_2236,N_24931,N_24747);
xor UO_2237 (O_2237,N_24638,N_24664);
nand UO_2238 (O_2238,N_24454,N_24693);
or UO_2239 (O_2239,N_24926,N_24888);
and UO_2240 (O_2240,N_24329,N_23866);
or UO_2241 (O_2241,N_24008,N_24459);
nor UO_2242 (O_2242,N_24952,N_23823);
nor UO_2243 (O_2243,N_24090,N_24279);
nor UO_2244 (O_2244,N_24016,N_24440);
and UO_2245 (O_2245,N_24546,N_24294);
nor UO_2246 (O_2246,N_23808,N_24468);
nand UO_2247 (O_2247,N_23916,N_24736);
or UO_2248 (O_2248,N_23934,N_24547);
nor UO_2249 (O_2249,N_23834,N_24735);
or UO_2250 (O_2250,N_24998,N_23947);
or UO_2251 (O_2251,N_24488,N_24733);
nand UO_2252 (O_2252,N_24748,N_24253);
or UO_2253 (O_2253,N_24591,N_24065);
nand UO_2254 (O_2254,N_24695,N_24058);
and UO_2255 (O_2255,N_24103,N_23865);
xor UO_2256 (O_2256,N_24723,N_24170);
and UO_2257 (O_2257,N_24290,N_24937);
xnor UO_2258 (O_2258,N_24090,N_24788);
xnor UO_2259 (O_2259,N_24107,N_24678);
nor UO_2260 (O_2260,N_24394,N_24210);
and UO_2261 (O_2261,N_23958,N_24576);
xor UO_2262 (O_2262,N_24252,N_24804);
and UO_2263 (O_2263,N_24899,N_24193);
nand UO_2264 (O_2264,N_24849,N_24508);
or UO_2265 (O_2265,N_23915,N_24814);
or UO_2266 (O_2266,N_24756,N_24898);
nand UO_2267 (O_2267,N_24423,N_24630);
xnor UO_2268 (O_2268,N_24398,N_24589);
nand UO_2269 (O_2269,N_24666,N_24588);
xor UO_2270 (O_2270,N_24606,N_24076);
nor UO_2271 (O_2271,N_23843,N_24381);
xor UO_2272 (O_2272,N_24384,N_24738);
nor UO_2273 (O_2273,N_24955,N_23837);
and UO_2274 (O_2274,N_23763,N_24123);
nand UO_2275 (O_2275,N_24094,N_24783);
nand UO_2276 (O_2276,N_24253,N_24352);
and UO_2277 (O_2277,N_24716,N_24705);
xor UO_2278 (O_2278,N_24841,N_24261);
xor UO_2279 (O_2279,N_24925,N_24451);
nand UO_2280 (O_2280,N_24344,N_24873);
nor UO_2281 (O_2281,N_24876,N_23781);
and UO_2282 (O_2282,N_24404,N_23758);
and UO_2283 (O_2283,N_24994,N_24450);
or UO_2284 (O_2284,N_23996,N_23975);
and UO_2285 (O_2285,N_23843,N_24895);
nand UO_2286 (O_2286,N_24145,N_24676);
and UO_2287 (O_2287,N_24109,N_24528);
nor UO_2288 (O_2288,N_24588,N_24327);
nand UO_2289 (O_2289,N_24764,N_24770);
xnor UO_2290 (O_2290,N_24703,N_24052);
nor UO_2291 (O_2291,N_24062,N_24572);
nand UO_2292 (O_2292,N_24777,N_24515);
xor UO_2293 (O_2293,N_24459,N_24265);
and UO_2294 (O_2294,N_24854,N_24025);
xnor UO_2295 (O_2295,N_24865,N_24790);
or UO_2296 (O_2296,N_24893,N_23791);
or UO_2297 (O_2297,N_23903,N_24074);
xnor UO_2298 (O_2298,N_24690,N_24065);
xor UO_2299 (O_2299,N_24038,N_24909);
nand UO_2300 (O_2300,N_24322,N_24112);
or UO_2301 (O_2301,N_24759,N_23889);
and UO_2302 (O_2302,N_23907,N_24970);
nand UO_2303 (O_2303,N_24367,N_23829);
and UO_2304 (O_2304,N_24338,N_24912);
and UO_2305 (O_2305,N_24980,N_24828);
xnor UO_2306 (O_2306,N_24230,N_24357);
and UO_2307 (O_2307,N_24549,N_23965);
or UO_2308 (O_2308,N_23898,N_23774);
and UO_2309 (O_2309,N_24109,N_23781);
nand UO_2310 (O_2310,N_23788,N_24228);
or UO_2311 (O_2311,N_24693,N_24699);
nor UO_2312 (O_2312,N_23807,N_24959);
or UO_2313 (O_2313,N_24155,N_24399);
nor UO_2314 (O_2314,N_24967,N_24705);
nor UO_2315 (O_2315,N_24929,N_24773);
xor UO_2316 (O_2316,N_24691,N_24630);
or UO_2317 (O_2317,N_24439,N_23921);
xor UO_2318 (O_2318,N_24478,N_24033);
xor UO_2319 (O_2319,N_24321,N_24487);
or UO_2320 (O_2320,N_24437,N_24685);
xnor UO_2321 (O_2321,N_24076,N_23959);
nor UO_2322 (O_2322,N_24690,N_24758);
xor UO_2323 (O_2323,N_23760,N_24151);
nand UO_2324 (O_2324,N_24263,N_24541);
and UO_2325 (O_2325,N_24342,N_24218);
or UO_2326 (O_2326,N_23778,N_24787);
or UO_2327 (O_2327,N_24641,N_24885);
and UO_2328 (O_2328,N_24104,N_24734);
or UO_2329 (O_2329,N_24785,N_24539);
and UO_2330 (O_2330,N_23766,N_24878);
and UO_2331 (O_2331,N_24964,N_24380);
and UO_2332 (O_2332,N_24583,N_24534);
or UO_2333 (O_2333,N_24733,N_24809);
and UO_2334 (O_2334,N_23927,N_24258);
xnor UO_2335 (O_2335,N_24548,N_24270);
xor UO_2336 (O_2336,N_24408,N_24959);
nand UO_2337 (O_2337,N_23833,N_24385);
nor UO_2338 (O_2338,N_24293,N_23834);
xor UO_2339 (O_2339,N_23975,N_24347);
nor UO_2340 (O_2340,N_24424,N_24706);
nand UO_2341 (O_2341,N_24093,N_24579);
and UO_2342 (O_2342,N_23830,N_24903);
nor UO_2343 (O_2343,N_24128,N_24683);
xor UO_2344 (O_2344,N_24664,N_24500);
or UO_2345 (O_2345,N_24235,N_24835);
xnor UO_2346 (O_2346,N_24574,N_24011);
or UO_2347 (O_2347,N_24914,N_23965);
and UO_2348 (O_2348,N_23830,N_24890);
or UO_2349 (O_2349,N_24048,N_24204);
xnor UO_2350 (O_2350,N_24992,N_24231);
nand UO_2351 (O_2351,N_24747,N_24155);
and UO_2352 (O_2352,N_24606,N_24824);
and UO_2353 (O_2353,N_23942,N_24119);
nand UO_2354 (O_2354,N_23754,N_24660);
or UO_2355 (O_2355,N_23762,N_23896);
and UO_2356 (O_2356,N_24741,N_24104);
nor UO_2357 (O_2357,N_24394,N_24168);
xor UO_2358 (O_2358,N_24329,N_24489);
xnor UO_2359 (O_2359,N_24147,N_24390);
and UO_2360 (O_2360,N_24576,N_24104);
xor UO_2361 (O_2361,N_24090,N_24249);
nor UO_2362 (O_2362,N_24374,N_24422);
xor UO_2363 (O_2363,N_24735,N_24641);
nand UO_2364 (O_2364,N_24707,N_24955);
xor UO_2365 (O_2365,N_23959,N_23823);
nand UO_2366 (O_2366,N_24551,N_23919);
xor UO_2367 (O_2367,N_24860,N_24650);
nor UO_2368 (O_2368,N_24521,N_24179);
xnor UO_2369 (O_2369,N_23930,N_24154);
and UO_2370 (O_2370,N_23957,N_23825);
nor UO_2371 (O_2371,N_24105,N_23929);
nand UO_2372 (O_2372,N_24415,N_24036);
xor UO_2373 (O_2373,N_23861,N_23910);
and UO_2374 (O_2374,N_24368,N_24339);
nor UO_2375 (O_2375,N_24840,N_24265);
nor UO_2376 (O_2376,N_24859,N_24005);
or UO_2377 (O_2377,N_24894,N_24510);
or UO_2378 (O_2378,N_24114,N_23971);
nand UO_2379 (O_2379,N_23821,N_23811);
nor UO_2380 (O_2380,N_24725,N_24641);
nand UO_2381 (O_2381,N_24602,N_24800);
nand UO_2382 (O_2382,N_24921,N_24376);
xnor UO_2383 (O_2383,N_24073,N_24981);
or UO_2384 (O_2384,N_23934,N_23793);
xnor UO_2385 (O_2385,N_24712,N_24530);
and UO_2386 (O_2386,N_24698,N_24063);
and UO_2387 (O_2387,N_24016,N_23864);
nor UO_2388 (O_2388,N_24107,N_24034);
xnor UO_2389 (O_2389,N_23973,N_24091);
xnor UO_2390 (O_2390,N_24693,N_24555);
nor UO_2391 (O_2391,N_24433,N_23797);
xnor UO_2392 (O_2392,N_23849,N_24633);
xnor UO_2393 (O_2393,N_23988,N_24698);
nor UO_2394 (O_2394,N_24190,N_24194);
nand UO_2395 (O_2395,N_24273,N_24555);
nor UO_2396 (O_2396,N_24424,N_24190);
xor UO_2397 (O_2397,N_24934,N_23794);
xnor UO_2398 (O_2398,N_24417,N_24402);
nand UO_2399 (O_2399,N_24500,N_24103);
nor UO_2400 (O_2400,N_24675,N_24178);
nor UO_2401 (O_2401,N_24693,N_23773);
and UO_2402 (O_2402,N_24081,N_24512);
nand UO_2403 (O_2403,N_24069,N_24041);
or UO_2404 (O_2404,N_23920,N_24614);
xor UO_2405 (O_2405,N_24317,N_24104);
or UO_2406 (O_2406,N_24331,N_24986);
nand UO_2407 (O_2407,N_23914,N_24729);
nand UO_2408 (O_2408,N_24373,N_23875);
nor UO_2409 (O_2409,N_23782,N_24782);
or UO_2410 (O_2410,N_24414,N_24925);
or UO_2411 (O_2411,N_24792,N_24915);
xnor UO_2412 (O_2412,N_24543,N_24533);
and UO_2413 (O_2413,N_24312,N_23899);
nand UO_2414 (O_2414,N_23854,N_24642);
and UO_2415 (O_2415,N_24285,N_24457);
nand UO_2416 (O_2416,N_24266,N_24061);
and UO_2417 (O_2417,N_24951,N_24107);
and UO_2418 (O_2418,N_24048,N_24424);
or UO_2419 (O_2419,N_23848,N_24977);
nand UO_2420 (O_2420,N_24822,N_24767);
xor UO_2421 (O_2421,N_24467,N_24202);
nand UO_2422 (O_2422,N_24634,N_23765);
nor UO_2423 (O_2423,N_24678,N_24403);
and UO_2424 (O_2424,N_24510,N_24845);
nor UO_2425 (O_2425,N_24877,N_24583);
nor UO_2426 (O_2426,N_24726,N_24662);
and UO_2427 (O_2427,N_24205,N_23794);
or UO_2428 (O_2428,N_24770,N_24785);
or UO_2429 (O_2429,N_24501,N_24385);
xor UO_2430 (O_2430,N_24064,N_24435);
or UO_2431 (O_2431,N_24382,N_24646);
or UO_2432 (O_2432,N_23954,N_24207);
nor UO_2433 (O_2433,N_24389,N_23896);
nand UO_2434 (O_2434,N_24205,N_24216);
and UO_2435 (O_2435,N_23819,N_24286);
nor UO_2436 (O_2436,N_24248,N_23896);
and UO_2437 (O_2437,N_24743,N_23971);
nor UO_2438 (O_2438,N_23888,N_24742);
nor UO_2439 (O_2439,N_24802,N_24689);
and UO_2440 (O_2440,N_24660,N_23760);
nor UO_2441 (O_2441,N_24283,N_24503);
nor UO_2442 (O_2442,N_24032,N_24306);
nand UO_2443 (O_2443,N_24671,N_23863);
or UO_2444 (O_2444,N_24486,N_24889);
xnor UO_2445 (O_2445,N_23878,N_24695);
nand UO_2446 (O_2446,N_24185,N_24163);
xor UO_2447 (O_2447,N_24243,N_24792);
xor UO_2448 (O_2448,N_24596,N_24509);
or UO_2449 (O_2449,N_24312,N_24578);
nor UO_2450 (O_2450,N_24904,N_24706);
nand UO_2451 (O_2451,N_24730,N_24638);
xnor UO_2452 (O_2452,N_24148,N_24198);
xnor UO_2453 (O_2453,N_24107,N_24121);
and UO_2454 (O_2454,N_24816,N_23809);
and UO_2455 (O_2455,N_24385,N_23899);
xnor UO_2456 (O_2456,N_24891,N_24817);
and UO_2457 (O_2457,N_23912,N_24688);
xnor UO_2458 (O_2458,N_23760,N_23940);
nand UO_2459 (O_2459,N_24199,N_24124);
nor UO_2460 (O_2460,N_24910,N_24420);
and UO_2461 (O_2461,N_24782,N_24851);
nand UO_2462 (O_2462,N_24554,N_24040);
and UO_2463 (O_2463,N_23916,N_24429);
and UO_2464 (O_2464,N_24039,N_24330);
and UO_2465 (O_2465,N_24471,N_24189);
nor UO_2466 (O_2466,N_24324,N_23814);
xor UO_2467 (O_2467,N_24239,N_24370);
nor UO_2468 (O_2468,N_24561,N_24035);
xnor UO_2469 (O_2469,N_24455,N_24412);
nand UO_2470 (O_2470,N_23791,N_24075);
nand UO_2471 (O_2471,N_24443,N_24574);
xor UO_2472 (O_2472,N_23922,N_24494);
xor UO_2473 (O_2473,N_23774,N_24260);
nand UO_2474 (O_2474,N_24973,N_24960);
and UO_2475 (O_2475,N_24682,N_23806);
nor UO_2476 (O_2476,N_23754,N_24276);
nand UO_2477 (O_2477,N_24417,N_23752);
or UO_2478 (O_2478,N_24087,N_24621);
nor UO_2479 (O_2479,N_23935,N_24802);
xnor UO_2480 (O_2480,N_23864,N_23860);
nor UO_2481 (O_2481,N_24168,N_24182);
and UO_2482 (O_2482,N_23878,N_24086);
nor UO_2483 (O_2483,N_24757,N_24190);
nand UO_2484 (O_2484,N_24347,N_24772);
nand UO_2485 (O_2485,N_24935,N_23846);
nor UO_2486 (O_2486,N_24600,N_23904);
nor UO_2487 (O_2487,N_24050,N_24256);
xnor UO_2488 (O_2488,N_23857,N_24501);
nand UO_2489 (O_2489,N_24977,N_24383);
and UO_2490 (O_2490,N_24896,N_24168);
or UO_2491 (O_2491,N_24603,N_24634);
xnor UO_2492 (O_2492,N_23774,N_24571);
and UO_2493 (O_2493,N_23909,N_23998);
and UO_2494 (O_2494,N_24888,N_24602);
and UO_2495 (O_2495,N_24672,N_24327);
xnor UO_2496 (O_2496,N_24987,N_24089);
and UO_2497 (O_2497,N_23824,N_23853);
nor UO_2498 (O_2498,N_24131,N_24057);
nor UO_2499 (O_2499,N_24422,N_23939);
xor UO_2500 (O_2500,N_24761,N_24774);
and UO_2501 (O_2501,N_24176,N_24895);
nor UO_2502 (O_2502,N_23821,N_24241);
nand UO_2503 (O_2503,N_24517,N_24468);
xor UO_2504 (O_2504,N_24415,N_24886);
nor UO_2505 (O_2505,N_24706,N_23798);
nor UO_2506 (O_2506,N_24495,N_24260);
nand UO_2507 (O_2507,N_23887,N_24872);
nor UO_2508 (O_2508,N_24255,N_24762);
or UO_2509 (O_2509,N_23774,N_23831);
xnor UO_2510 (O_2510,N_23805,N_24030);
xor UO_2511 (O_2511,N_24892,N_24240);
and UO_2512 (O_2512,N_24461,N_24365);
and UO_2513 (O_2513,N_23810,N_23923);
nor UO_2514 (O_2514,N_24729,N_23870);
and UO_2515 (O_2515,N_24979,N_24055);
and UO_2516 (O_2516,N_24734,N_23886);
or UO_2517 (O_2517,N_23885,N_24573);
nor UO_2518 (O_2518,N_24749,N_23862);
nand UO_2519 (O_2519,N_24397,N_24123);
xor UO_2520 (O_2520,N_23914,N_24776);
nor UO_2521 (O_2521,N_24627,N_24686);
xnor UO_2522 (O_2522,N_24420,N_24280);
and UO_2523 (O_2523,N_24142,N_23827);
nand UO_2524 (O_2524,N_24801,N_24985);
and UO_2525 (O_2525,N_24510,N_24338);
nor UO_2526 (O_2526,N_23856,N_24621);
and UO_2527 (O_2527,N_24773,N_24353);
or UO_2528 (O_2528,N_24738,N_24153);
xor UO_2529 (O_2529,N_24498,N_23858);
nand UO_2530 (O_2530,N_24538,N_24101);
or UO_2531 (O_2531,N_24865,N_24079);
nor UO_2532 (O_2532,N_24464,N_24096);
xor UO_2533 (O_2533,N_24754,N_24880);
nor UO_2534 (O_2534,N_24425,N_24287);
nand UO_2535 (O_2535,N_24155,N_24164);
nor UO_2536 (O_2536,N_24643,N_23775);
or UO_2537 (O_2537,N_24259,N_24082);
or UO_2538 (O_2538,N_24137,N_24392);
and UO_2539 (O_2539,N_24670,N_24574);
nand UO_2540 (O_2540,N_24847,N_24588);
nand UO_2541 (O_2541,N_24889,N_24558);
and UO_2542 (O_2542,N_23995,N_24524);
nand UO_2543 (O_2543,N_24460,N_23783);
xor UO_2544 (O_2544,N_24495,N_24128);
and UO_2545 (O_2545,N_24099,N_23796);
and UO_2546 (O_2546,N_24781,N_24192);
nand UO_2547 (O_2547,N_23976,N_24954);
nor UO_2548 (O_2548,N_24684,N_24009);
nor UO_2549 (O_2549,N_24784,N_24119);
nor UO_2550 (O_2550,N_24869,N_24303);
and UO_2551 (O_2551,N_24482,N_24500);
nor UO_2552 (O_2552,N_24455,N_24674);
nor UO_2553 (O_2553,N_24881,N_24258);
nor UO_2554 (O_2554,N_24269,N_24544);
nand UO_2555 (O_2555,N_24699,N_23794);
nand UO_2556 (O_2556,N_24741,N_24064);
nor UO_2557 (O_2557,N_24392,N_24577);
or UO_2558 (O_2558,N_24069,N_23950);
and UO_2559 (O_2559,N_24883,N_24066);
nor UO_2560 (O_2560,N_23976,N_24048);
xor UO_2561 (O_2561,N_24229,N_24203);
and UO_2562 (O_2562,N_24105,N_24695);
nor UO_2563 (O_2563,N_23875,N_24554);
nand UO_2564 (O_2564,N_24435,N_24942);
xor UO_2565 (O_2565,N_24453,N_24473);
and UO_2566 (O_2566,N_24528,N_24175);
nand UO_2567 (O_2567,N_24556,N_24196);
nor UO_2568 (O_2568,N_24667,N_23777);
or UO_2569 (O_2569,N_24015,N_23884);
or UO_2570 (O_2570,N_24786,N_24644);
or UO_2571 (O_2571,N_24232,N_24036);
or UO_2572 (O_2572,N_24433,N_24191);
nand UO_2573 (O_2573,N_24285,N_24238);
nand UO_2574 (O_2574,N_24147,N_24326);
nand UO_2575 (O_2575,N_24778,N_24640);
xnor UO_2576 (O_2576,N_23823,N_23858);
and UO_2577 (O_2577,N_24631,N_24260);
xor UO_2578 (O_2578,N_23998,N_23871);
nand UO_2579 (O_2579,N_24579,N_23921);
xnor UO_2580 (O_2580,N_24343,N_24176);
or UO_2581 (O_2581,N_24736,N_24104);
nand UO_2582 (O_2582,N_24586,N_24508);
and UO_2583 (O_2583,N_24520,N_24381);
and UO_2584 (O_2584,N_24699,N_24359);
xor UO_2585 (O_2585,N_24915,N_24214);
or UO_2586 (O_2586,N_23777,N_23875);
and UO_2587 (O_2587,N_24011,N_24638);
nor UO_2588 (O_2588,N_24416,N_24679);
or UO_2589 (O_2589,N_24513,N_24746);
or UO_2590 (O_2590,N_23830,N_24069);
nor UO_2591 (O_2591,N_24015,N_24971);
nor UO_2592 (O_2592,N_23822,N_24710);
xor UO_2593 (O_2593,N_23826,N_24923);
or UO_2594 (O_2594,N_24108,N_23976);
or UO_2595 (O_2595,N_24448,N_24209);
nand UO_2596 (O_2596,N_24810,N_23887);
nand UO_2597 (O_2597,N_24793,N_24271);
or UO_2598 (O_2598,N_24811,N_24911);
nor UO_2599 (O_2599,N_24304,N_24316);
nand UO_2600 (O_2600,N_24854,N_23875);
nand UO_2601 (O_2601,N_24797,N_24727);
xor UO_2602 (O_2602,N_23900,N_24738);
xnor UO_2603 (O_2603,N_24081,N_23996);
or UO_2604 (O_2604,N_24327,N_24389);
and UO_2605 (O_2605,N_23824,N_24488);
nand UO_2606 (O_2606,N_24128,N_24345);
nand UO_2607 (O_2607,N_24608,N_23754);
xor UO_2608 (O_2608,N_24990,N_24160);
and UO_2609 (O_2609,N_24642,N_24274);
xnor UO_2610 (O_2610,N_24164,N_24566);
nor UO_2611 (O_2611,N_24177,N_24642);
and UO_2612 (O_2612,N_24984,N_24032);
xnor UO_2613 (O_2613,N_24944,N_24546);
xnor UO_2614 (O_2614,N_24816,N_24672);
and UO_2615 (O_2615,N_24840,N_24569);
and UO_2616 (O_2616,N_24917,N_24947);
nand UO_2617 (O_2617,N_23841,N_24166);
or UO_2618 (O_2618,N_24562,N_24758);
xor UO_2619 (O_2619,N_24550,N_24761);
xnor UO_2620 (O_2620,N_24560,N_24407);
nor UO_2621 (O_2621,N_24436,N_24610);
and UO_2622 (O_2622,N_24516,N_24190);
nor UO_2623 (O_2623,N_24389,N_23814);
and UO_2624 (O_2624,N_24994,N_23752);
nand UO_2625 (O_2625,N_24507,N_24039);
nand UO_2626 (O_2626,N_23981,N_24540);
or UO_2627 (O_2627,N_24022,N_24740);
nand UO_2628 (O_2628,N_23980,N_24540);
nor UO_2629 (O_2629,N_23768,N_24999);
or UO_2630 (O_2630,N_24168,N_24334);
xnor UO_2631 (O_2631,N_23836,N_24169);
nor UO_2632 (O_2632,N_24130,N_23846);
and UO_2633 (O_2633,N_24408,N_23800);
and UO_2634 (O_2634,N_24448,N_24572);
nor UO_2635 (O_2635,N_24950,N_24829);
nand UO_2636 (O_2636,N_24412,N_24738);
and UO_2637 (O_2637,N_24147,N_24217);
or UO_2638 (O_2638,N_24778,N_24996);
nand UO_2639 (O_2639,N_24802,N_24607);
xnor UO_2640 (O_2640,N_24115,N_24432);
or UO_2641 (O_2641,N_24134,N_23827);
nand UO_2642 (O_2642,N_24848,N_24245);
xnor UO_2643 (O_2643,N_24112,N_24002);
or UO_2644 (O_2644,N_24142,N_24967);
xnor UO_2645 (O_2645,N_24284,N_24568);
nand UO_2646 (O_2646,N_23827,N_24768);
nor UO_2647 (O_2647,N_24184,N_23858);
or UO_2648 (O_2648,N_24745,N_24978);
and UO_2649 (O_2649,N_24211,N_23802);
nor UO_2650 (O_2650,N_24091,N_24717);
nand UO_2651 (O_2651,N_24081,N_24647);
nand UO_2652 (O_2652,N_24409,N_23937);
and UO_2653 (O_2653,N_24317,N_24848);
and UO_2654 (O_2654,N_24962,N_23938);
xnor UO_2655 (O_2655,N_24752,N_24866);
nand UO_2656 (O_2656,N_24309,N_24068);
or UO_2657 (O_2657,N_24906,N_24450);
nor UO_2658 (O_2658,N_24590,N_24019);
xnor UO_2659 (O_2659,N_24272,N_24377);
nor UO_2660 (O_2660,N_24091,N_23842);
xnor UO_2661 (O_2661,N_24629,N_23765);
or UO_2662 (O_2662,N_24324,N_24512);
xor UO_2663 (O_2663,N_24982,N_24370);
and UO_2664 (O_2664,N_24488,N_24786);
and UO_2665 (O_2665,N_24518,N_24725);
and UO_2666 (O_2666,N_24595,N_24495);
xnor UO_2667 (O_2667,N_23796,N_24755);
nor UO_2668 (O_2668,N_24038,N_24994);
or UO_2669 (O_2669,N_24049,N_24930);
xor UO_2670 (O_2670,N_24232,N_24415);
nor UO_2671 (O_2671,N_24524,N_24762);
and UO_2672 (O_2672,N_24290,N_24677);
or UO_2673 (O_2673,N_24276,N_24427);
nor UO_2674 (O_2674,N_24867,N_24529);
nor UO_2675 (O_2675,N_24780,N_24128);
and UO_2676 (O_2676,N_24997,N_24743);
xnor UO_2677 (O_2677,N_23791,N_23873);
or UO_2678 (O_2678,N_24441,N_24290);
xnor UO_2679 (O_2679,N_24116,N_23956);
nor UO_2680 (O_2680,N_24752,N_23823);
or UO_2681 (O_2681,N_24821,N_24953);
and UO_2682 (O_2682,N_24310,N_24034);
xnor UO_2683 (O_2683,N_24718,N_24744);
or UO_2684 (O_2684,N_23919,N_24665);
nor UO_2685 (O_2685,N_24263,N_24239);
and UO_2686 (O_2686,N_24716,N_23938);
nor UO_2687 (O_2687,N_24645,N_24634);
or UO_2688 (O_2688,N_24684,N_24781);
nand UO_2689 (O_2689,N_23841,N_24915);
xor UO_2690 (O_2690,N_24673,N_24179);
xnor UO_2691 (O_2691,N_23896,N_24429);
nand UO_2692 (O_2692,N_23826,N_24887);
nor UO_2693 (O_2693,N_24665,N_24305);
xnor UO_2694 (O_2694,N_24838,N_24092);
nor UO_2695 (O_2695,N_24522,N_24040);
xnor UO_2696 (O_2696,N_23946,N_24721);
xor UO_2697 (O_2697,N_24227,N_23969);
nor UO_2698 (O_2698,N_24210,N_24030);
nand UO_2699 (O_2699,N_24135,N_24659);
nor UO_2700 (O_2700,N_24248,N_24167);
or UO_2701 (O_2701,N_24551,N_23772);
xor UO_2702 (O_2702,N_24797,N_23936);
or UO_2703 (O_2703,N_24078,N_24607);
and UO_2704 (O_2704,N_24009,N_24435);
and UO_2705 (O_2705,N_24713,N_24507);
nor UO_2706 (O_2706,N_23967,N_24529);
xor UO_2707 (O_2707,N_24640,N_24505);
and UO_2708 (O_2708,N_23949,N_24270);
or UO_2709 (O_2709,N_24124,N_24085);
nor UO_2710 (O_2710,N_24297,N_24015);
nand UO_2711 (O_2711,N_24471,N_24814);
xnor UO_2712 (O_2712,N_24548,N_23904);
nand UO_2713 (O_2713,N_24878,N_23771);
nor UO_2714 (O_2714,N_24964,N_24406);
and UO_2715 (O_2715,N_23984,N_23815);
xnor UO_2716 (O_2716,N_24949,N_23813);
and UO_2717 (O_2717,N_24733,N_24253);
or UO_2718 (O_2718,N_24221,N_24732);
and UO_2719 (O_2719,N_24775,N_23899);
xor UO_2720 (O_2720,N_24315,N_24467);
xor UO_2721 (O_2721,N_24082,N_24558);
or UO_2722 (O_2722,N_24789,N_23941);
or UO_2723 (O_2723,N_24154,N_24519);
and UO_2724 (O_2724,N_24193,N_24737);
or UO_2725 (O_2725,N_23873,N_23933);
nor UO_2726 (O_2726,N_23970,N_23997);
nor UO_2727 (O_2727,N_24798,N_24067);
and UO_2728 (O_2728,N_24356,N_24621);
nor UO_2729 (O_2729,N_23911,N_24307);
and UO_2730 (O_2730,N_23821,N_24801);
nor UO_2731 (O_2731,N_24263,N_23956);
nor UO_2732 (O_2732,N_24852,N_24906);
nand UO_2733 (O_2733,N_24332,N_24888);
xor UO_2734 (O_2734,N_24420,N_24132);
or UO_2735 (O_2735,N_24457,N_24970);
or UO_2736 (O_2736,N_24347,N_23755);
or UO_2737 (O_2737,N_24439,N_24868);
nand UO_2738 (O_2738,N_24842,N_24300);
and UO_2739 (O_2739,N_24716,N_24647);
or UO_2740 (O_2740,N_24070,N_24826);
and UO_2741 (O_2741,N_23832,N_23784);
nand UO_2742 (O_2742,N_24242,N_23759);
and UO_2743 (O_2743,N_24367,N_24999);
nand UO_2744 (O_2744,N_24753,N_23787);
nand UO_2745 (O_2745,N_24677,N_24346);
and UO_2746 (O_2746,N_24354,N_24477);
nor UO_2747 (O_2747,N_24217,N_24624);
and UO_2748 (O_2748,N_23795,N_24995);
nor UO_2749 (O_2749,N_24786,N_24329);
nand UO_2750 (O_2750,N_24913,N_24349);
nor UO_2751 (O_2751,N_24283,N_24708);
and UO_2752 (O_2752,N_24883,N_24311);
and UO_2753 (O_2753,N_24794,N_24686);
nor UO_2754 (O_2754,N_23751,N_24514);
xnor UO_2755 (O_2755,N_23859,N_24156);
or UO_2756 (O_2756,N_24509,N_24686);
xor UO_2757 (O_2757,N_24036,N_24588);
xor UO_2758 (O_2758,N_24092,N_24637);
and UO_2759 (O_2759,N_24713,N_24170);
nor UO_2760 (O_2760,N_23928,N_24103);
or UO_2761 (O_2761,N_24768,N_23871);
xor UO_2762 (O_2762,N_24986,N_24517);
or UO_2763 (O_2763,N_23772,N_23795);
nor UO_2764 (O_2764,N_24026,N_24911);
xnor UO_2765 (O_2765,N_24053,N_24586);
or UO_2766 (O_2766,N_24282,N_24937);
nor UO_2767 (O_2767,N_23853,N_23871);
and UO_2768 (O_2768,N_24197,N_24207);
nor UO_2769 (O_2769,N_24968,N_24736);
nor UO_2770 (O_2770,N_24649,N_23817);
xnor UO_2771 (O_2771,N_24916,N_24946);
nor UO_2772 (O_2772,N_23948,N_24803);
and UO_2773 (O_2773,N_24850,N_24473);
nand UO_2774 (O_2774,N_24697,N_24887);
nand UO_2775 (O_2775,N_24389,N_24575);
nor UO_2776 (O_2776,N_24832,N_24661);
and UO_2777 (O_2777,N_24406,N_24974);
xnor UO_2778 (O_2778,N_24456,N_23930);
xnor UO_2779 (O_2779,N_24908,N_24930);
and UO_2780 (O_2780,N_23907,N_24254);
nand UO_2781 (O_2781,N_24792,N_24764);
nor UO_2782 (O_2782,N_23754,N_24765);
nand UO_2783 (O_2783,N_24646,N_24457);
or UO_2784 (O_2784,N_23985,N_24433);
and UO_2785 (O_2785,N_24431,N_23926);
nand UO_2786 (O_2786,N_24584,N_24855);
nand UO_2787 (O_2787,N_24062,N_24868);
or UO_2788 (O_2788,N_24658,N_23785);
nand UO_2789 (O_2789,N_24352,N_24955);
xor UO_2790 (O_2790,N_24661,N_23992);
nor UO_2791 (O_2791,N_24426,N_23938);
or UO_2792 (O_2792,N_24512,N_24797);
and UO_2793 (O_2793,N_23842,N_24250);
nand UO_2794 (O_2794,N_24114,N_24715);
xnor UO_2795 (O_2795,N_24448,N_24942);
nor UO_2796 (O_2796,N_23858,N_23995);
xnor UO_2797 (O_2797,N_24310,N_23968);
nand UO_2798 (O_2798,N_24016,N_24934);
and UO_2799 (O_2799,N_24535,N_23928);
xor UO_2800 (O_2800,N_24676,N_24226);
or UO_2801 (O_2801,N_23768,N_23791);
nand UO_2802 (O_2802,N_24461,N_24352);
nor UO_2803 (O_2803,N_23784,N_24986);
and UO_2804 (O_2804,N_24605,N_24419);
or UO_2805 (O_2805,N_24246,N_23857);
xor UO_2806 (O_2806,N_24060,N_23814);
nor UO_2807 (O_2807,N_24410,N_23844);
xnor UO_2808 (O_2808,N_24713,N_24607);
nor UO_2809 (O_2809,N_24175,N_24302);
nand UO_2810 (O_2810,N_24607,N_24966);
and UO_2811 (O_2811,N_24918,N_24187);
nor UO_2812 (O_2812,N_24199,N_24223);
or UO_2813 (O_2813,N_24824,N_24760);
or UO_2814 (O_2814,N_24096,N_24277);
nor UO_2815 (O_2815,N_24997,N_24042);
and UO_2816 (O_2816,N_24942,N_24909);
xor UO_2817 (O_2817,N_24435,N_24994);
or UO_2818 (O_2818,N_24193,N_24930);
nand UO_2819 (O_2819,N_24751,N_23887);
xnor UO_2820 (O_2820,N_24965,N_24364);
or UO_2821 (O_2821,N_24112,N_23871);
and UO_2822 (O_2822,N_24225,N_24675);
xnor UO_2823 (O_2823,N_24412,N_24048);
nand UO_2824 (O_2824,N_24431,N_24854);
nand UO_2825 (O_2825,N_24818,N_24739);
and UO_2826 (O_2826,N_24958,N_24629);
or UO_2827 (O_2827,N_23937,N_24424);
and UO_2828 (O_2828,N_24157,N_24298);
xnor UO_2829 (O_2829,N_24943,N_24593);
nand UO_2830 (O_2830,N_23994,N_24374);
and UO_2831 (O_2831,N_24884,N_24771);
or UO_2832 (O_2832,N_23835,N_23806);
and UO_2833 (O_2833,N_24766,N_24428);
nand UO_2834 (O_2834,N_24123,N_24272);
nand UO_2835 (O_2835,N_24710,N_23790);
nor UO_2836 (O_2836,N_24533,N_23809);
and UO_2837 (O_2837,N_24898,N_24389);
nor UO_2838 (O_2838,N_24418,N_24986);
nor UO_2839 (O_2839,N_24084,N_24023);
or UO_2840 (O_2840,N_24571,N_24762);
nand UO_2841 (O_2841,N_24464,N_24828);
or UO_2842 (O_2842,N_24043,N_24481);
or UO_2843 (O_2843,N_24767,N_24220);
nand UO_2844 (O_2844,N_24933,N_24329);
xor UO_2845 (O_2845,N_24424,N_24633);
and UO_2846 (O_2846,N_24982,N_24197);
and UO_2847 (O_2847,N_24169,N_24464);
nand UO_2848 (O_2848,N_24533,N_24160);
and UO_2849 (O_2849,N_24237,N_24540);
nand UO_2850 (O_2850,N_24344,N_24375);
and UO_2851 (O_2851,N_24021,N_24031);
nand UO_2852 (O_2852,N_24372,N_24345);
nor UO_2853 (O_2853,N_24969,N_24958);
or UO_2854 (O_2854,N_24551,N_23977);
and UO_2855 (O_2855,N_24626,N_24134);
xor UO_2856 (O_2856,N_24289,N_24075);
nor UO_2857 (O_2857,N_24782,N_24317);
nor UO_2858 (O_2858,N_24313,N_23754);
nor UO_2859 (O_2859,N_24065,N_24972);
nor UO_2860 (O_2860,N_24422,N_24997);
xnor UO_2861 (O_2861,N_23865,N_23803);
nand UO_2862 (O_2862,N_24466,N_23939);
or UO_2863 (O_2863,N_23763,N_23909);
or UO_2864 (O_2864,N_23858,N_24188);
nor UO_2865 (O_2865,N_24065,N_24806);
and UO_2866 (O_2866,N_24946,N_23945);
xnor UO_2867 (O_2867,N_23984,N_23832);
nand UO_2868 (O_2868,N_24471,N_23895);
nor UO_2869 (O_2869,N_24029,N_23923);
and UO_2870 (O_2870,N_23982,N_24049);
nand UO_2871 (O_2871,N_23933,N_24267);
xor UO_2872 (O_2872,N_24356,N_24393);
nand UO_2873 (O_2873,N_24001,N_24714);
nand UO_2874 (O_2874,N_24516,N_24037);
nand UO_2875 (O_2875,N_24952,N_24336);
and UO_2876 (O_2876,N_24572,N_23936);
and UO_2877 (O_2877,N_24627,N_24023);
or UO_2878 (O_2878,N_23981,N_23820);
or UO_2879 (O_2879,N_24588,N_24001);
xnor UO_2880 (O_2880,N_24220,N_24077);
nor UO_2881 (O_2881,N_24560,N_24988);
xnor UO_2882 (O_2882,N_23827,N_24409);
xor UO_2883 (O_2883,N_24083,N_24409);
xor UO_2884 (O_2884,N_24692,N_24280);
or UO_2885 (O_2885,N_24523,N_23826);
or UO_2886 (O_2886,N_24205,N_24590);
nor UO_2887 (O_2887,N_24649,N_24917);
nor UO_2888 (O_2888,N_24706,N_24158);
or UO_2889 (O_2889,N_24025,N_24283);
xor UO_2890 (O_2890,N_24640,N_23877);
xor UO_2891 (O_2891,N_24514,N_24175);
or UO_2892 (O_2892,N_24631,N_24445);
nor UO_2893 (O_2893,N_23802,N_24302);
nor UO_2894 (O_2894,N_23958,N_23857);
xnor UO_2895 (O_2895,N_24654,N_23881);
nand UO_2896 (O_2896,N_24634,N_24781);
or UO_2897 (O_2897,N_23842,N_24941);
nor UO_2898 (O_2898,N_24254,N_24158);
nor UO_2899 (O_2899,N_24528,N_24165);
nand UO_2900 (O_2900,N_24477,N_24749);
nand UO_2901 (O_2901,N_24892,N_24040);
nand UO_2902 (O_2902,N_24160,N_24794);
xnor UO_2903 (O_2903,N_23874,N_24225);
or UO_2904 (O_2904,N_24465,N_24217);
nand UO_2905 (O_2905,N_24921,N_24316);
nand UO_2906 (O_2906,N_23914,N_24527);
nand UO_2907 (O_2907,N_24226,N_23940);
and UO_2908 (O_2908,N_23785,N_23880);
nor UO_2909 (O_2909,N_24847,N_24598);
xnor UO_2910 (O_2910,N_24044,N_24663);
xor UO_2911 (O_2911,N_24411,N_24670);
and UO_2912 (O_2912,N_24434,N_24457);
nor UO_2913 (O_2913,N_24509,N_24838);
and UO_2914 (O_2914,N_23969,N_23773);
xor UO_2915 (O_2915,N_24358,N_24481);
or UO_2916 (O_2916,N_24282,N_24324);
or UO_2917 (O_2917,N_24362,N_24385);
xnor UO_2918 (O_2918,N_24231,N_24168);
nand UO_2919 (O_2919,N_24020,N_24900);
and UO_2920 (O_2920,N_24960,N_24368);
xnor UO_2921 (O_2921,N_24142,N_23931);
xnor UO_2922 (O_2922,N_24078,N_23799);
nor UO_2923 (O_2923,N_24448,N_24503);
and UO_2924 (O_2924,N_24606,N_24067);
or UO_2925 (O_2925,N_23866,N_24906);
or UO_2926 (O_2926,N_24252,N_24537);
and UO_2927 (O_2927,N_24055,N_24220);
nor UO_2928 (O_2928,N_24429,N_24747);
nor UO_2929 (O_2929,N_24722,N_24310);
or UO_2930 (O_2930,N_23968,N_24688);
xnor UO_2931 (O_2931,N_23844,N_24594);
or UO_2932 (O_2932,N_23920,N_24464);
and UO_2933 (O_2933,N_24255,N_23819);
nor UO_2934 (O_2934,N_24027,N_24325);
and UO_2935 (O_2935,N_24648,N_24259);
nor UO_2936 (O_2936,N_24195,N_24005);
or UO_2937 (O_2937,N_23763,N_24395);
xor UO_2938 (O_2938,N_24659,N_24179);
or UO_2939 (O_2939,N_24076,N_24345);
and UO_2940 (O_2940,N_23917,N_23935);
nor UO_2941 (O_2941,N_24148,N_24932);
and UO_2942 (O_2942,N_24321,N_24577);
nor UO_2943 (O_2943,N_24364,N_24852);
or UO_2944 (O_2944,N_24848,N_23868);
nand UO_2945 (O_2945,N_24288,N_24014);
nor UO_2946 (O_2946,N_23794,N_24083);
and UO_2947 (O_2947,N_24346,N_24926);
xnor UO_2948 (O_2948,N_24092,N_24047);
or UO_2949 (O_2949,N_23940,N_24147);
xor UO_2950 (O_2950,N_24027,N_24468);
nand UO_2951 (O_2951,N_24169,N_24813);
nand UO_2952 (O_2952,N_24016,N_24809);
nor UO_2953 (O_2953,N_24448,N_24197);
nand UO_2954 (O_2954,N_24981,N_24177);
and UO_2955 (O_2955,N_24848,N_24592);
or UO_2956 (O_2956,N_24527,N_23765);
nor UO_2957 (O_2957,N_24801,N_23991);
xnor UO_2958 (O_2958,N_23871,N_23972);
xor UO_2959 (O_2959,N_24841,N_23835);
nor UO_2960 (O_2960,N_24530,N_24860);
nor UO_2961 (O_2961,N_24548,N_23942);
and UO_2962 (O_2962,N_24272,N_24774);
or UO_2963 (O_2963,N_24685,N_24585);
or UO_2964 (O_2964,N_24821,N_24182);
nand UO_2965 (O_2965,N_24640,N_23772);
nand UO_2966 (O_2966,N_24609,N_24945);
xor UO_2967 (O_2967,N_24713,N_24165);
nor UO_2968 (O_2968,N_24152,N_24247);
nor UO_2969 (O_2969,N_23789,N_23831);
xor UO_2970 (O_2970,N_24644,N_23863);
xor UO_2971 (O_2971,N_24708,N_24933);
or UO_2972 (O_2972,N_24461,N_24893);
nor UO_2973 (O_2973,N_24385,N_24592);
xor UO_2974 (O_2974,N_24066,N_24958);
or UO_2975 (O_2975,N_24969,N_24873);
nand UO_2976 (O_2976,N_23777,N_23840);
or UO_2977 (O_2977,N_24638,N_23789);
nor UO_2978 (O_2978,N_24147,N_24385);
and UO_2979 (O_2979,N_24638,N_24043);
xnor UO_2980 (O_2980,N_24489,N_24097);
nor UO_2981 (O_2981,N_23756,N_24104);
xnor UO_2982 (O_2982,N_24122,N_23752);
or UO_2983 (O_2983,N_24797,N_24015);
nor UO_2984 (O_2984,N_24285,N_24371);
or UO_2985 (O_2985,N_23916,N_24612);
nand UO_2986 (O_2986,N_23843,N_24959);
and UO_2987 (O_2987,N_23781,N_23839);
nor UO_2988 (O_2988,N_24110,N_24170);
nor UO_2989 (O_2989,N_23847,N_24756);
nor UO_2990 (O_2990,N_24408,N_23939);
xnor UO_2991 (O_2991,N_23896,N_23909);
xnor UO_2992 (O_2992,N_23901,N_24808);
and UO_2993 (O_2993,N_23800,N_24374);
nand UO_2994 (O_2994,N_24060,N_24068);
nand UO_2995 (O_2995,N_24106,N_24027);
xnor UO_2996 (O_2996,N_24611,N_23889);
nand UO_2997 (O_2997,N_23870,N_23820);
and UO_2998 (O_2998,N_24765,N_23891);
nor UO_2999 (O_2999,N_24193,N_23759);
endmodule