module basic_750_5000_1000_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_631,In_256);
xor U1 (N_1,In_593,In_367);
and U2 (N_2,In_204,In_446);
xor U3 (N_3,In_507,In_230);
nor U4 (N_4,In_660,In_48);
and U5 (N_5,In_186,In_749);
and U6 (N_6,In_23,In_592);
xnor U7 (N_7,In_199,In_375);
or U8 (N_8,In_328,In_474);
or U9 (N_9,In_545,In_203);
or U10 (N_10,In_667,In_700);
or U11 (N_11,In_222,In_188);
xor U12 (N_12,In_527,In_440);
xor U13 (N_13,In_513,In_502);
xor U14 (N_14,In_308,In_82);
nor U15 (N_15,In_649,In_601);
xnor U16 (N_16,In_466,In_81);
nor U17 (N_17,In_694,In_60);
nor U18 (N_18,In_63,In_118);
xor U19 (N_19,In_143,In_457);
xor U20 (N_20,In_445,In_427);
or U21 (N_21,In_242,In_9);
xnor U22 (N_22,In_268,In_119);
nand U23 (N_23,In_448,In_486);
and U24 (N_24,In_595,In_290);
or U25 (N_25,In_438,In_506);
xor U26 (N_26,In_79,In_471);
or U27 (N_27,In_183,In_740);
xor U28 (N_28,In_106,In_152);
nand U29 (N_29,In_169,In_621);
or U30 (N_30,In_100,In_662);
xor U31 (N_31,In_389,In_373);
and U32 (N_32,In_167,In_391);
nor U33 (N_33,In_158,In_163);
and U34 (N_34,In_463,In_668);
xnor U35 (N_35,In_735,In_295);
nor U36 (N_36,In_741,In_363);
xnor U37 (N_37,In_742,In_408);
xnor U38 (N_38,In_539,In_386);
nand U39 (N_39,In_399,In_586);
or U40 (N_40,In_24,In_229);
xor U41 (N_41,In_569,In_615);
nor U42 (N_42,In_334,In_115);
or U43 (N_43,In_5,In_336);
xor U44 (N_44,In_33,In_747);
nor U45 (N_45,In_546,In_355);
nor U46 (N_46,In_73,In_514);
xnor U47 (N_47,In_429,In_257);
xor U48 (N_48,In_715,In_622);
xor U49 (N_49,In_589,In_42);
xnor U50 (N_50,In_383,In_164);
or U51 (N_51,In_263,In_642);
nand U52 (N_52,In_40,In_208);
or U53 (N_53,In_364,In_55);
xnor U54 (N_54,In_231,In_479);
or U55 (N_55,In_721,In_184);
or U56 (N_56,In_273,In_542);
or U57 (N_57,In_746,In_0);
or U58 (N_58,In_619,In_266);
or U59 (N_59,In_217,In_65);
nand U60 (N_60,In_254,In_430);
or U61 (N_61,In_543,In_585);
nor U62 (N_62,In_674,In_117);
or U63 (N_63,In_180,In_142);
nor U64 (N_64,In_25,In_602);
xor U65 (N_65,In_38,In_96);
and U66 (N_66,In_11,In_415);
and U67 (N_67,In_561,In_531);
and U68 (N_68,In_663,In_44);
nor U69 (N_69,In_47,In_551);
nand U70 (N_70,In_719,In_197);
and U71 (N_71,In_381,In_15);
xor U72 (N_72,In_594,In_282);
xor U73 (N_73,In_144,In_504);
nand U74 (N_74,In_179,In_573);
nand U75 (N_75,In_736,In_43);
or U76 (N_76,In_613,In_76);
and U77 (N_77,In_372,In_554);
and U78 (N_78,In_330,In_260);
xor U79 (N_79,In_567,In_552);
xor U80 (N_80,In_270,In_534);
nor U81 (N_81,In_600,In_181);
nand U82 (N_82,In_124,In_512);
xnor U83 (N_83,In_394,In_459);
nand U84 (N_84,In_718,In_174);
nor U85 (N_85,In_299,In_332);
nand U86 (N_86,In_85,In_313);
nor U87 (N_87,In_198,In_583);
and U88 (N_88,In_467,In_3);
nor U89 (N_89,In_650,In_220);
nand U90 (N_90,In_434,In_587);
nand U91 (N_91,In_251,In_666);
or U92 (N_92,In_210,In_262);
nor U93 (N_93,In_553,In_572);
nand U94 (N_94,In_664,In_245);
nand U95 (N_95,In_105,In_215);
nand U96 (N_96,In_702,In_192);
xnor U97 (N_97,In_352,In_101);
and U98 (N_98,In_249,In_46);
nor U99 (N_99,In_175,In_547);
nor U100 (N_100,In_291,In_303);
xor U101 (N_101,In_378,In_22);
nand U102 (N_102,In_120,In_521);
or U103 (N_103,In_219,In_345);
nand U104 (N_104,In_456,In_316);
or U105 (N_105,In_398,In_89);
nor U106 (N_106,In_239,In_691);
and U107 (N_107,In_97,In_522);
nand U108 (N_108,In_342,In_423);
or U109 (N_109,In_671,In_509);
nor U110 (N_110,In_558,In_454);
nand U111 (N_111,In_689,In_307);
or U112 (N_112,In_550,In_238);
nand U113 (N_113,In_370,In_125);
or U114 (N_114,In_200,In_116);
nor U115 (N_115,In_354,In_21);
nor U116 (N_116,In_726,In_397);
nor U117 (N_117,In_194,In_409);
nand U118 (N_118,In_647,In_114);
nor U119 (N_119,In_253,In_629);
nor U120 (N_120,In_108,In_744);
xnor U121 (N_121,In_733,In_218);
or U122 (N_122,In_693,In_669);
and U123 (N_123,In_289,In_310);
nor U124 (N_124,In_30,In_155);
nand U125 (N_125,In_7,In_732);
nor U126 (N_126,In_157,In_722);
xor U127 (N_127,In_562,In_297);
xor U128 (N_128,In_280,In_248);
and U129 (N_129,In_433,In_528);
nor U130 (N_130,In_641,In_505);
xor U131 (N_131,In_340,In_435);
or U132 (N_132,In_576,In_94);
nor U133 (N_133,In_609,In_258);
or U134 (N_134,In_444,In_275);
and U135 (N_135,In_465,In_491);
or U136 (N_136,In_503,In_317);
nand U137 (N_137,In_196,In_516);
or U138 (N_138,In_489,In_533);
or U139 (N_139,In_255,In_300);
and U140 (N_140,In_329,In_61);
and U141 (N_141,In_86,In_72);
xnor U142 (N_142,In_580,In_520);
nand U143 (N_143,In_374,In_637);
nand U144 (N_144,In_57,In_278);
and U145 (N_145,In_421,In_78);
and U146 (N_146,In_406,In_577);
and U147 (N_147,In_630,In_306);
xor U148 (N_148,In_298,In_476);
nand U149 (N_149,In_511,In_645);
xor U150 (N_150,In_682,In_632);
nand U151 (N_151,In_154,In_95);
or U152 (N_152,In_523,In_274);
nor U153 (N_153,In_214,In_627);
or U154 (N_154,In_341,In_131);
xor U155 (N_155,In_233,In_205);
nor U156 (N_156,In_49,In_697);
nor U157 (N_157,In_56,In_172);
xnor U158 (N_158,In_54,In_714);
xor U159 (N_159,In_481,In_243);
nor U160 (N_160,In_318,In_309);
nand U161 (N_161,In_128,In_395);
nor U162 (N_162,In_327,In_487);
nand U163 (N_163,In_51,In_344);
nand U164 (N_164,In_193,In_734);
or U165 (N_165,In_655,In_713);
nor U166 (N_166,In_599,In_261);
or U167 (N_167,In_292,In_638);
or U168 (N_168,In_234,In_166);
nand U169 (N_169,In_515,In_469);
or U170 (N_170,In_416,In_12);
or U171 (N_171,In_449,In_141);
and U172 (N_172,In_566,In_276);
nor U173 (N_173,In_482,In_623);
nand U174 (N_174,In_111,In_259);
nand U175 (N_175,In_675,In_343);
nor U176 (N_176,In_696,In_745);
nand U177 (N_177,In_490,In_92);
nand U178 (N_178,In_360,In_296);
nor U179 (N_179,In_35,In_392);
nand U180 (N_180,In_676,In_347);
xnor U181 (N_181,In_451,In_703);
and U182 (N_182,In_563,In_739);
and U183 (N_183,In_147,In_688);
nand U184 (N_184,In_314,In_530);
xor U185 (N_185,In_730,In_425);
xor U186 (N_186,In_350,In_137);
or U187 (N_187,In_62,In_387);
or U188 (N_188,In_109,In_657);
nor U189 (N_189,In_346,In_351);
nor U190 (N_190,In_652,In_401);
and U191 (N_191,In_335,In_711);
or U192 (N_192,In_312,In_685);
and U193 (N_193,In_302,In_134);
xnor U194 (N_194,In_283,In_692);
xor U195 (N_195,In_556,In_162);
and U196 (N_196,In_738,In_485);
nor U197 (N_197,In_83,In_160);
and U198 (N_198,In_411,In_420);
nand U199 (N_199,In_221,In_525);
xor U200 (N_200,In_37,In_6);
and U201 (N_201,In_470,In_548);
or U202 (N_202,In_428,In_705);
nand U203 (N_203,In_99,In_450);
and U204 (N_204,In_150,In_13);
nand U205 (N_205,In_709,In_322);
and U206 (N_206,In_31,In_368);
nor U207 (N_207,In_447,In_468);
or U208 (N_208,In_492,In_604);
nand U209 (N_209,In_182,In_698);
nor U210 (N_210,In_75,In_455);
and U211 (N_211,In_417,In_555);
and U212 (N_212,In_236,In_517);
and U213 (N_213,In_337,In_149);
xor U214 (N_214,In_396,In_442);
nand U215 (N_215,In_497,In_460);
and U216 (N_216,In_107,In_603);
nand U217 (N_217,In_384,In_178);
or U218 (N_218,In_670,In_737);
nand U219 (N_219,In_281,In_494);
nor U220 (N_220,In_356,In_213);
and U221 (N_221,In_70,In_661);
xnor U222 (N_222,In_541,In_206);
or U223 (N_223,In_358,In_265);
xnor U224 (N_224,In_320,In_45);
xnor U225 (N_225,In_480,In_87);
and U226 (N_226,In_635,In_605);
and U227 (N_227,In_185,In_598);
xor U228 (N_228,In_584,In_235);
nor U229 (N_229,In_385,In_161);
xor U230 (N_230,In_612,In_319);
xor U231 (N_231,In_339,In_64);
xnor U232 (N_232,In_410,In_267);
or U233 (N_233,In_404,In_201);
nor U234 (N_234,In_225,In_103);
nand U235 (N_235,In_110,In_699);
xnor U236 (N_236,In_723,In_640);
nor U237 (N_237,In_148,In_653);
nand U238 (N_238,In_366,In_681);
and U239 (N_239,In_654,In_237);
nand U240 (N_240,In_496,In_93);
and U241 (N_241,In_50,In_701);
nand U242 (N_242,In_683,In_228);
xnor U243 (N_243,In_269,In_597);
or U244 (N_244,In_91,In_126);
nor U245 (N_245,In_359,In_628);
or U246 (N_246,In_400,In_393);
or U247 (N_247,In_211,In_311);
nand U248 (N_248,In_287,In_538);
or U249 (N_249,In_643,In_644);
and U250 (N_250,In_2,In_146);
nand U251 (N_251,In_684,In_241);
and U252 (N_252,In_98,In_177);
and U253 (N_253,In_560,In_568);
nand U254 (N_254,In_607,In_532);
xnor U255 (N_255,In_582,In_74);
and U256 (N_256,In_659,In_365);
and U257 (N_257,In_729,In_41);
nand U258 (N_258,In_570,In_357);
nand U259 (N_259,In_176,In_537);
and U260 (N_260,In_136,In_324);
and U261 (N_261,In_325,In_695);
or U262 (N_262,In_677,In_724);
or U263 (N_263,In_540,In_611);
or U264 (N_264,In_422,In_461);
nand U265 (N_265,In_708,In_191);
and U266 (N_266,In_590,In_680);
or U267 (N_267,In_443,In_66);
and U268 (N_268,In_535,In_588);
or U269 (N_269,In_113,In_71);
xnor U270 (N_270,In_333,In_707);
or U271 (N_271,In_294,In_403);
nor U272 (N_272,In_493,In_690);
or U273 (N_273,In_304,In_1);
xor U274 (N_274,In_68,In_575);
or U275 (N_275,In_526,In_606);
and U276 (N_276,In_122,In_727);
xor U277 (N_277,In_686,In_288);
and U278 (N_278,In_4,In_501);
xnor U279 (N_279,In_250,In_651);
or U280 (N_280,In_704,In_478);
nor U281 (N_281,In_69,In_338);
nor U282 (N_282,In_227,In_376);
or U283 (N_283,In_18,In_321);
or U284 (N_284,In_656,In_315);
xor U285 (N_285,In_153,In_748);
nor U286 (N_286,In_39,In_135);
xnor U287 (N_287,In_633,In_151);
and U288 (N_288,In_59,In_578);
xnor U289 (N_289,In_518,In_488);
and U290 (N_290,In_710,In_725);
or U291 (N_291,In_564,In_139);
nand U292 (N_292,In_679,In_247);
nand U293 (N_293,In_286,In_8);
and U294 (N_294,In_130,In_610);
xor U295 (N_295,In_90,In_67);
xor U296 (N_296,In_17,In_648);
nand U297 (N_297,In_508,In_439);
nand U298 (N_298,In_596,In_323);
nor U299 (N_299,In_559,In_140);
nor U300 (N_300,In_84,In_731);
nor U301 (N_301,In_209,In_138);
nor U302 (N_302,In_716,In_240);
and U303 (N_303,In_424,In_102);
nor U304 (N_304,In_743,In_207);
nor U305 (N_305,In_519,In_171);
or U306 (N_306,In_168,In_305);
or U307 (N_307,In_706,In_436);
or U308 (N_308,In_616,In_264);
or U309 (N_309,In_571,In_301);
xnor U310 (N_310,In_624,In_202);
xnor U311 (N_311,In_687,In_14);
nor U312 (N_312,In_495,In_382);
xnor U313 (N_313,In_58,In_88);
and U314 (N_314,In_379,In_53);
nor U315 (N_315,In_10,In_591);
xnor U316 (N_316,In_380,In_190);
nand U317 (N_317,In_349,In_665);
nor U318 (N_318,In_499,In_472);
xor U319 (N_319,In_20,In_159);
xnor U320 (N_320,In_636,In_565);
nand U321 (N_321,In_614,In_32);
nand U322 (N_322,In_617,In_272);
or U323 (N_323,In_34,In_544);
nand U324 (N_324,In_326,In_170);
nor U325 (N_325,In_361,In_419);
xnor U326 (N_326,In_413,In_529);
and U327 (N_327,In_464,In_244);
xor U328 (N_328,In_672,In_536);
or U329 (N_329,In_618,In_189);
nor U330 (N_330,In_484,In_121);
nand U331 (N_331,In_717,In_388);
xnor U332 (N_332,In_279,In_16);
nor U333 (N_333,In_165,In_483);
xor U334 (N_334,In_293,In_19);
nor U335 (N_335,In_720,In_414);
nor U336 (N_336,In_452,In_27);
and U337 (N_337,In_104,In_36);
and U338 (N_338,In_271,In_646);
xor U339 (N_339,In_348,In_285);
xor U340 (N_340,In_625,In_639);
nor U341 (N_341,In_549,In_232);
xnor U342 (N_342,In_477,In_626);
nand U343 (N_343,In_195,In_673);
or U344 (N_344,In_123,In_458);
or U345 (N_345,In_246,In_473);
nor U346 (N_346,In_432,In_112);
nand U347 (N_347,In_252,In_132);
and U348 (N_348,In_407,In_426);
and U349 (N_349,In_212,In_441);
nor U350 (N_350,In_462,In_453);
xor U351 (N_351,In_127,In_223);
nand U352 (N_352,In_431,In_524);
nand U353 (N_353,In_510,In_728);
xor U354 (N_354,In_412,In_579);
and U355 (N_355,In_475,In_129);
or U356 (N_356,In_29,In_658);
or U357 (N_357,In_557,In_712);
xnor U358 (N_358,In_418,In_369);
nor U359 (N_359,In_581,In_437);
nor U360 (N_360,In_620,In_634);
nand U361 (N_361,In_405,In_224);
nor U362 (N_362,In_574,In_133);
or U363 (N_363,In_187,In_331);
or U364 (N_364,In_77,In_284);
or U365 (N_365,In_500,In_156);
and U366 (N_366,In_26,In_353);
nand U367 (N_367,In_678,In_390);
nor U368 (N_368,In_362,In_28);
xor U369 (N_369,In_52,In_216);
xor U370 (N_370,In_498,In_173);
nand U371 (N_371,In_145,In_80);
nand U372 (N_372,In_377,In_371);
xor U373 (N_373,In_277,In_608);
and U374 (N_374,In_402,In_226);
nor U375 (N_375,In_48,In_251);
and U376 (N_376,In_123,In_515);
nor U377 (N_377,In_279,In_463);
or U378 (N_378,In_574,In_301);
and U379 (N_379,In_488,In_388);
or U380 (N_380,In_106,In_314);
nand U381 (N_381,In_278,In_741);
nand U382 (N_382,In_585,In_421);
and U383 (N_383,In_515,In_138);
nor U384 (N_384,In_206,In_290);
or U385 (N_385,In_326,In_660);
xnor U386 (N_386,In_39,In_617);
nor U387 (N_387,In_378,In_466);
and U388 (N_388,In_579,In_93);
nor U389 (N_389,In_728,In_451);
xnor U390 (N_390,In_126,In_542);
xor U391 (N_391,In_525,In_65);
or U392 (N_392,In_96,In_18);
nor U393 (N_393,In_555,In_631);
xor U394 (N_394,In_101,In_294);
nor U395 (N_395,In_606,In_351);
xnor U396 (N_396,In_669,In_61);
or U397 (N_397,In_701,In_237);
and U398 (N_398,In_42,In_364);
or U399 (N_399,In_601,In_123);
or U400 (N_400,In_620,In_690);
nor U401 (N_401,In_294,In_8);
nand U402 (N_402,In_586,In_423);
nand U403 (N_403,In_47,In_601);
xnor U404 (N_404,In_163,In_410);
or U405 (N_405,In_353,In_27);
nor U406 (N_406,In_664,In_603);
or U407 (N_407,In_559,In_595);
xor U408 (N_408,In_557,In_126);
and U409 (N_409,In_173,In_473);
xor U410 (N_410,In_209,In_670);
and U411 (N_411,In_531,In_415);
nor U412 (N_412,In_84,In_124);
and U413 (N_413,In_517,In_609);
nor U414 (N_414,In_319,In_556);
or U415 (N_415,In_10,In_691);
and U416 (N_416,In_116,In_624);
and U417 (N_417,In_730,In_170);
nand U418 (N_418,In_444,In_73);
nand U419 (N_419,In_364,In_68);
xor U420 (N_420,In_485,In_242);
or U421 (N_421,In_451,In_356);
nor U422 (N_422,In_283,In_18);
nand U423 (N_423,In_663,In_732);
and U424 (N_424,In_370,In_702);
xnor U425 (N_425,In_245,In_309);
nand U426 (N_426,In_152,In_253);
nor U427 (N_427,In_314,In_125);
nand U428 (N_428,In_199,In_481);
and U429 (N_429,In_702,In_99);
or U430 (N_430,In_342,In_214);
xor U431 (N_431,In_623,In_110);
and U432 (N_432,In_588,In_566);
and U433 (N_433,In_139,In_403);
nor U434 (N_434,In_336,In_312);
xnor U435 (N_435,In_739,In_327);
nor U436 (N_436,In_683,In_470);
nand U437 (N_437,In_650,In_442);
nand U438 (N_438,In_251,In_390);
nand U439 (N_439,In_516,In_445);
or U440 (N_440,In_170,In_240);
nor U441 (N_441,In_390,In_615);
and U442 (N_442,In_722,In_417);
or U443 (N_443,In_655,In_697);
or U444 (N_444,In_628,In_706);
and U445 (N_445,In_575,In_554);
nand U446 (N_446,In_108,In_468);
nand U447 (N_447,In_264,In_25);
xnor U448 (N_448,In_178,In_36);
or U449 (N_449,In_693,In_468);
and U450 (N_450,In_724,In_276);
or U451 (N_451,In_540,In_703);
nand U452 (N_452,In_114,In_743);
nand U453 (N_453,In_126,In_11);
and U454 (N_454,In_185,In_352);
nand U455 (N_455,In_412,In_317);
and U456 (N_456,In_673,In_253);
nand U457 (N_457,In_568,In_621);
or U458 (N_458,In_542,In_589);
or U459 (N_459,In_247,In_256);
xnor U460 (N_460,In_274,In_296);
nand U461 (N_461,In_155,In_404);
xnor U462 (N_462,In_101,In_364);
nand U463 (N_463,In_312,In_20);
nand U464 (N_464,In_288,In_498);
nor U465 (N_465,In_521,In_435);
or U466 (N_466,In_532,In_735);
nor U467 (N_467,In_463,In_706);
xnor U468 (N_468,In_561,In_689);
nand U469 (N_469,In_540,In_164);
nand U470 (N_470,In_198,In_239);
nand U471 (N_471,In_80,In_20);
and U472 (N_472,In_332,In_333);
and U473 (N_473,In_42,In_653);
xor U474 (N_474,In_40,In_331);
xnor U475 (N_475,In_413,In_549);
xnor U476 (N_476,In_707,In_356);
and U477 (N_477,In_377,In_133);
or U478 (N_478,In_618,In_146);
xnor U479 (N_479,In_618,In_720);
nand U480 (N_480,In_153,In_348);
xnor U481 (N_481,In_40,In_656);
and U482 (N_482,In_497,In_509);
or U483 (N_483,In_28,In_678);
or U484 (N_484,In_444,In_191);
or U485 (N_485,In_736,In_51);
nand U486 (N_486,In_620,In_644);
nor U487 (N_487,In_579,In_616);
or U488 (N_488,In_433,In_659);
and U489 (N_489,In_26,In_531);
nor U490 (N_490,In_7,In_584);
xor U491 (N_491,In_161,In_56);
xor U492 (N_492,In_557,In_52);
nor U493 (N_493,In_73,In_534);
nor U494 (N_494,In_489,In_228);
nand U495 (N_495,In_580,In_604);
and U496 (N_496,In_228,In_735);
nor U497 (N_497,In_383,In_102);
xnor U498 (N_498,In_288,In_210);
nor U499 (N_499,In_476,In_177);
nor U500 (N_500,In_151,In_181);
xor U501 (N_501,In_331,In_535);
and U502 (N_502,In_329,In_646);
nand U503 (N_503,In_317,In_270);
xnor U504 (N_504,In_574,In_101);
nor U505 (N_505,In_558,In_487);
nor U506 (N_506,In_488,In_652);
and U507 (N_507,In_67,In_281);
nand U508 (N_508,In_482,In_210);
and U509 (N_509,In_260,In_620);
xor U510 (N_510,In_665,In_0);
xor U511 (N_511,In_183,In_479);
nand U512 (N_512,In_278,In_671);
nor U513 (N_513,In_223,In_296);
or U514 (N_514,In_140,In_346);
and U515 (N_515,In_357,In_133);
and U516 (N_516,In_681,In_450);
xor U517 (N_517,In_206,In_501);
or U518 (N_518,In_509,In_427);
and U519 (N_519,In_40,In_441);
and U520 (N_520,In_113,In_462);
and U521 (N_521,In_580,In_703);
nor U522 (N_522,In_75,In_2);
or U523 (N_523,In_606,In_623);
nand U524 (N_524,In_636,In_255);
nor U525 (N_525,In_515,In_134);
or U526 (N_526,In_341,In_92);
or U527 (N_527,In_614,In_487);
and U528 (N_528,In_461,In_552);
xnor U529 (N_529,In_114,In_221);
xor U530 (N_530,In_364,In_161);
and U531 (N_531,In_453,In_40);
nor U532 (N_532,In_431,In_229);
and U533 (N_533,In_647,In_155);
and U534 (N_534,In_724,In_22);
xnor U535 (N_535,In_402,In_630);
nor U536 (N_536,In_541,In_480);
nor U537 (N_537,In_505,In_664);
or U538 (N_538,In_109,In_312);
xnor U539 (N_539,In_45,In_213);
nor U540 (N_540,In_494,In_200);
and U541 (N_541,In_123,In_67);
nand U542 (N_542,In_706,In_569);
nor U543 (N_543,In_69,In_589);
or U544 (N_544,In_336,In_225);
and U545 (N_545,In_102,In_191);
and U546 (N_546,In_484,In_520);
nand U547 (N_547,In_680,In_101);
nand U548 (N_548,In_432,In_74);
nand U549 (N_549,In_632,In_716);
xnor U550 (N_550,In_211,In_148);
nor U551 (N_551,In_609,In_351);
nor U552 (N_552,In_46,In_377);
and U553 (N_553,In_142,In_739);
xnor U554 (N_554,In_192,In_537);
xnor U555 (N_555,In_83,In_648);
and U556 (N_556,In_686,In_531);
nor U557 (N_557,In_145,In_493);
or U558 (N_558,In_436,In_174);
or U559 (N_559,In_26,In_124);
or U560 (N_560,In_58,In_505);
and U561 (N_561,In_284,In_169);
or U562 (N_562,In_391,In_372);
nand U563 (N_563,In_441,In_299);
or U564 (N_564,In_281,In_192);
nor U565 (N_565,In_339,In_156);
nand U566 (N_566,In_559,In_221);
or U567 (N_567,In_531,In_631);
or U568 (N_568,In_617,In_507);
nor U569 (N_569,In_611,In_175);
nand U570 (N_570,In_386,In_412);
nand U571 (N_571,In_368,In_569);
and U572 (N_572,In_429,In_498);
and U573 (N_573,In_299,In_254);
xor U574 (N_574,In_204,In_546);
xor U575 (N_575,In_290,In_344);
and U576 (N_576,In_487,In_415);
xnor U577 (N_577,In_87,In_219);
nor U578 (N_578,In_515,In_282);
nand U579 (N_579,In_274,In_394);
or U580 (N_580,In_81,In_97);
and U581 (N_581,In_359,In_395);
nand U582 (N_582,In_505,In_733);
nor U583 (N_583,In_252,In_646);
or U584 (N_584,In_701,In_102);
and U585 (N_585,In_519,In_46);
nand U586 (N_586,In_9,In_178);
nor U587 (N_587,In_313,In_286);
xnor U588 (N_588,In_494,In_710);
nand U589 (N_589,In_341,In_589);
nand U590 (N_590,In_113,In_170);
xor U591 (N_591,In_611,In_418);
xnor U592 (N_592,In_560,In_740);
nor U593 (N_593,In_61,In_205);
nand U594 (N_594,In_377,In_384);
and U595 (N_595,In_388,In_78);
and U596 (N_596,In_655,In_265);
or U597 (N_597,In_489,In_557);
nor U598 (N_598,In_249,In_283);
nand U599 (N_599,In_618,In_740);
nor U600 (N_600,In_6,In_77);
nor U601 (N_601,In_51,In_413);
and U602 (N_602,In_373,In_533);
xor U603 (N_603,In_548,In_436);
or U604 (N_604,In_134,In_518);
and U605 (N_605,In_336,In_430);
nor U606 (N_606,In_627,In_408);
or U607 (N_607,In_512,In_257);
xnor U608 (N_608,In_77,In_452);
and U609 (N_609,In_628,In_81);
and U610 (N_610,In_626,In_392);
xnor U611 (N_611,In_372,In_400);
nor U612 (N_612,In_731,In_543);
or U613 (N_613,In_656,In_724);
xor U614 (N_614,In_120,In_564);
nand U615 (N_615,In_364,In_435);
nor U616 (N_616,In_305,In_475);
nor U617 (N_617,In_450,In_8);
xnor U618 (N_618,In_423,In_19);
xnor U619 (N_619,In_399,In_544);
xnor U620 (N_620,In_45,In_375);
nand U621 (N_621,In_33,In_181);
and U622 (N_622,In_614,In_441);
nor U623 (N_623,In_514,In_183);
nand U624 (N_624,In_388,In_401);
nand U625 (N_625,In_1,In_39);
nand U626 (N_626,In_395,In_290);
nor U627 (N_627,In_746,In_178);
nor U628 (N_628,In_621,In_52);
or U629 (N_629,In_464,In_59);
or U630 (N_630,In_92,In_554);
xor U631 (N_631,In_401,In_182);
or U632 (N_632,In_340,In_660);
xnor U633 (N_633,In_276,In_78);
or U634 (N_634,In_631,In_705);
xnor U635 (N_635,In_525,In_591);
or U636 (N_636,In_730,In_493);
or U637 (N_637,In_330,In_623);
nand U638 (N_638,In_156,In_574);
xor U639 (N_639,In_371,In_643);
nor U640 (N_640,In_470,In_246);
xnor U641 (N_641,In_580,In_428);
and U642 (N_642,In_524,In_6);
nand U643 (N_643,In_431,In_592);
xnor U644 (N_644,In_220,In_80);
nor U645 (N_645,In_604,In_294);
or U646 (N_646,In_149,In_351);
nand U647 (N_647,In_489,In_150);
nand U648 (N_648,In_372,In_563);
xor U649 (N_649,In_395,In_239);
or U650 (N_650,In_462,In_67);
and U651 (N_651,In_286,In_53);
or U652 (N_652,In_376,In_695);
nand U653 (N_653,In_162,In_133);
and U654 (N_654,In_523,In_711);
xnor U655 (N_655,In_672,In_733);
or U656 (N_656,In_722,In_83);
xor U657 (N_657,In_21,In_219);
nand U658 (N_658,In_680,In_642);
nand U659 (N_659,In_157,In_422);
or U660 (N_660,In_746,In_63);
nor U661 (N_661,In_377,In_585);
nor U662 (N_662,In_554,In_739);
and U663 (N_663,In_314,In_628);
or U664 (N_664,In_551,In_243);
xnor U665 (N_665,In_231,In_13);
or U666 (N_666,In_255,In_279);
nor U667 (N_667,In_507,In_64);
xor U668 (N_668,In_262,In_655);
xnor U669 (N_669,In_475,In_539);
xor U670 (N_670,In_332,In_93);
and U671 (N_671,In_572,In_435);
nor U672 (N_672,In_488,In_100);
xor U673 (N_673,In_737,In_26);
or U674 (N_674,In_25,In_454);
xnor U675 (N_675,In_227,In_523);
nor U676 (N_676,In_365,In_116);
nand U677 (N_677,In_597,In_606);
nand U678 (N_678,In_31,In_669);
nor U679 (N_679,In_313,In_514);
and U680 (N_680,In_293,In_639);
xor U681 (N_681,In_161,In_412);
or U682 (N_682,In_311,In_121);
or U683 (N_683,In_675,In_372);
nand U684 (N_684,In_553,In_384);
nand U685 (N_685,In_27,In_157);
xnor U686 (N_686,In_230,In_125);
and U687 (N_687,In_734,In_315);
xor U688 (N_688,In_738,In_192);
or U689 (N_689,In_663,In_344);
xnor U690 (N_690,In_345,In_190);
and U691 (N_691,In_280,In_373);
and U692 (N_692,In_160,In_514);
or U693 (N_693,In_256,In_345);
nand U694 (N_694,In_373,In_338);
or U695 (N_695,In_5,In_329);
nor U696 (N_696,In_110,In_465);
and U697 (N_697,In_36,In_516);
or U698 (N_698,In_280,In_242);
xnor U699 (N_699,In_301,In_596);
xor U700 (N_700,In_459,In_172);
xor U701 (N_701,In_317,In_637);
and U702 (N_702,In_231,In_205);
and U703 (N_703,In_449,In_50);
and U704 (N_704,In_492,In_489);
nand U705 (N_705,In_157,In_547);
and U706 (N_706,In_68,In_40);
and U707 (N_707,In_185,In_49);
nand U708 (N_708,In_576,In_455);
and U709 (N_709,In_702,In_540);
or U710 (N_710,In_579,In_566);
or U711 (N_711,In_589,In_557);
or U712 (N_712,In_245,In_303);
and U713 (N_713,In_456,In_280);
or U714 (N_714,In_98,In_39);
and U715 (N_715,In_436,In_226);
or U716 (N_716,In_74,In_274);
or U717 (N_717,In_319,In_136);
nor U718 (N_718,In_75,In_445);
nand U719 (N_719,In_395,In_717);
or U720 (N_720,In_40,In_401);
nor U721 (N_721,In_584,In_24);
or U722 (N_722,In_407,In_395);
xor U723 (N_723,In_67,In_300);
nand U724 (N_724,In_617,In_391);
xnor U725 (N_725,In_384,In_149);
xnor U726 (N_726,In_489,In_675);
xnor U727 (N_727,In_636,In_323);
nor U728 (N_728,In_428,In_249);
nand U729 (N_729,In_80,In_101);
nor U730 (N_730,In_504,In_409);
nor U731 (N_731,In_376,In_70);
xor U732 (N_732,In_258,In_67);
nand U733 (N_733,In_178,In_713);
nand U734 (N_734,In_502,In_343);
xnor U735 (N_735,In_196,In_713);
xnor U736 (N_736,In_661,In_354);
nand U737 (N_737,In_586,In_121);
nor U738 (N_738,In_528,In_543);
or U739 (N_739,In_83,In_476);
and U740 (N_740,In_116,In_697);
and U741 (N_741,In_417,In_21);
or U742 (N_742,In_229,In_635);
or U743 (N_743,In_343,In_538);
nand U744 (N_744,In_77,In_737);
and U745 (N_745,In_381,In_169);
xor U746 (N_746,In_337,In_508);
or U747 (N_747,In_461,In_702);
or U748 (N_748,In_586,In_293);
nor U749 (N_749,In_502,In_163);
and U750 (N_750,In_544,In_624);
nand U751 (N_751,In_336,In_4);
and U752 (N_752,In_31,In_393);
and U753 (N_753,In_177,In_356);
nand U754 (N_754,In_658,In_719);
or U755 (N_755,In_573,In_608);
nor U756 (N_756,In_739,In_581);
nand U757 (N_757,In_419,In_404);
or U758 (N_758,In_133,In_336);
xnor U759 (N_759,In_191,In_630);
xnor U760 (N_760,In_666,In_165);
nand U761 (N_761,In_395,In_676);
nor U762 (N_762,In_644,In_430);
nor U763 (N_763,In_613,In_567);
and U764 (N_764,In_251,In_55);
or U765 (N_765,In_458,In_113);
xor U766 (N_766,In_647,In_37);
nor U767 (N_767,In_558,In_150);
nand U768 (N_768,In_477,In_366);
xor U769 (N_769,In_251,In_507);
nor U770 (N_770,In_24,In_371);
xnor U771 (N_771,In_535,In_124);
xnor U772 (N_772,In_484,In_360);
xor U773 (N_773,In_147,In_482);
or U774 (N_774,In_507,In_48);
xnor U775 (N_775,In_260,In_515);
xnor U776 (N_776,In_553,In_708);
xor U777 (N_777,In_206,In_706);
nand U778 (N_778,In_450,In_610);
and U779 (N_779,In_629,In_94);
xnor U780 (N_780,In_363,In_674);
nor U781 (N_781,In_611,In_384);
and U782 (N_782,In_714,In_370);
and U783 (N_783,In_717,In_507);
nor U784 (N_784,In_517,In_258);
xor U785 (N_785,In_609,In_115);
or U786 (N_786,In_72,In_696);
and U787 (N_787,In_673,In_4);
or U788 (N_788,In_414,In_221);
and U789 (N_789,In_364,In_395);
and U790 (N_790,In_660,In_227);
xnor U791 (N_791,In_478,In_141);
xnor U792 (N_792,In_96,In_335);
xor U793 (N_793,In_686,In_748);
xor U794 (N_794,In_289,In_504);
nand U795 (N_795,In_132,In_678);
or U796 (N_796,In_339,In_504);
and U797 (N_797,In_748,In_558);
nand U798 (N_798,In_528,In_654);
and U799 (N_799,In_195,In_748);
xor U800 (N_800,In_212,In_309);
nor U801 (N_801,In_290,In_716);
or U802 (N_802,In_107,In_198);
nand U803 (N_803,In_352,In_537);
and U804 (N_804,In_79,In_344);
nand U805 (N_805,In_207,In_185);
or U806 (N_806,In_610,In_291);
nand U807 (N_807,In_395,In_240);
or U808 (N_808,In_476,In_402);
and U809 (N_809,In_507,In_748);
nor U810 (N_810,In_242,In_623);
or U811 (N_811,In_253,In_82);
or U812 (N_812,In_438,In_43);
nand U813 (N_813,In_382,In_62);
nor U814 (N_814,In_492,In_152);
xor U815 (N_815,In_165,In_202);
xor U816 (N_816,In_134,In_105);
xor U817 (N_817,In_638,In_686);
and U818 (N_818,In_426,In_224);
xnor U819 (N_819,In_539,In_121);
or U820 (N_820,In_190,In_489);
xor U821 (N_821,In_42,In_99);
nor U822 (N_822,In_300,In_477);
xnor U823 (N_823,In_38,In_418);
nor U824 (N_824,In_738,In_190);
and U825 (N_825,In_397,In_554);
nand U826 (N_826,In_396,In_252);
xnor U827 (N_827,In_234,In_497);
xnor U828 (N_828,In_429,In_608);
xor U829 (N_829,In_421,In_411);
and U830 (N_830,In_173,In_34);
and U831 (N_831,In_280,In_18);
nor U832 (N_832,In_481,In_106);
or U833 (N_833,In_143,In_334);
or U834 (N_834,In_608,In_219);
or U835 (N_835,In_423,In_30);
or U836 (N_836,In_173,In_277);
nand U837 (N_837,In_657,In_423);
xnor U838 (N_838,In_671,In_491);
nand U839 (N_839,In_448,In_351);
xnor U840 (N_840,In_459,In_504);
or U841 (N_841,In_432,In_13);
nor U842 (N_842,In_601,In_539);
or U843 (N_843,In_439,In_473);
and U844 (N_844,In_656,In_177);
xnor U845 (N_845,In_482,In_85);
and U846 (N_846,In_167,In_608);
nor U847 (N_847,In_105,In_630);
and U848 (N_848,In_658,In_512);
xor U849 (N_849,In_4,In_415);
xor U850 (N_850,In_37,In_631);
nand U851 (N_851,In_103,In_180);
nor U852 (N_852,In_749,In_453);
xor U853 (N_853,In_337,In_601);
xnor U854 (N_854,In_315,In_409);
or U855 (N_855,In_689,In_257);
nor U856 (N_856,In_683,In_463);
or U857 (N_857,In_259,In_103);
or U858 (N_858,In_526,In_431);
or U859 (N_859,In_421,In_184);
nand U860 (N_860,In_10,In_198);
and U861 (N_861,In_21,In_373);
xnor U862 (N_862,In_405,In_308);
xor U863 (N_863,In_41,In_699);
and U864 (N_864,In_6,In_377);
nor U865 (N_865,In_702,In_200);
xor U866 (N_866,In_749,In_448);
nand U867 (N_867,In_47,In_497);
nand U868 (N_868,In_627,In_123);
nor U869 (N_869,In_661,In_24);
and U870 (N_870,In_184,In_724);
nor U871 (N_871,In_687,In_475);
nor U872 (N_872,In_530,In_358);
or U873 (N_873,In_488,In_364);
nor U874 (N_874,In_528,In_660);
or U875 (N_875,In_51,In_127);
nand U876 (N_876,In_457,In_180);
and U877 (N_877,In_413,In_8);
nor U878 (N_878,In_70,In_675);
nand U879 (N_879,In_402,In_134);
xnor U880 (N_880,In_154,In_336);
and U881 (N_881,In_172,In_494);
and U882 (N_882,In_78,In_417);
xor U883 (N_883,In_523,In_609);
or U884 (N_884,In_572,In_316);
or U885 (N_885,In_630,In_94);
xor U886 (N_886,In_283,In_559);
xnor U887 (N_887,In_137,In_657);
or U888 (N_888,In_45,In_412);
nor U889 (N_889,In_457,In_192);
or U890 (N_890,In_567,In_518);
or U891 (N_891,In_457,In_475);
and U892 (N_892,In_583,In_50);
xor U893 (N_893,In_276,In_304);
and U894 (N_894,In_481,In_459);
xnor U895 (N_895,In_356,In_47);
and U896 (N_896,In_136,In_278);
nor U897 (N_897,In_398,In_456);
nor U898 (N_898,In_669,In_367);
and U899 (N_899,In_651,In_606);
nand U900 (N_900,In_479,In_632);
xnor U901 (N_901,In_503,In_529);
and U902 (N_902,In_344,In_218);
and U903 (N_903,In_531,In_394);
and U904 (N_904,In_507,In_604);
nor U905 (N_905,In_647,In_320);
and U906 (N_906,In_738,In_608);
xnor U907 (N_907,In_107,In_214);
and U908 (N_908,In_729,In_373);
nand U909 (N_909,In_165,In_248);
and U910 (N_910,In_222,In_321);
nand U911 (N_911,In_408,In_41);
and U912 (N_912,In_56,In_663);
and U913 (N_913,In_680,In_59);
and U914 (N_914,In_210,In_124);
and U915 (N_915,In_746,In_566);
nand U916 (N_916,In_743,In_557);
and U917 (N_917,In_245,In_74);
nand U918 (N_918,In_82,In_425);
nor U919 (N_919,In_488,In_6);
xor U920 (N_920,In_108,In_119);
or U921 (N_921,In_70,In_554);
nand U922 (N_922,In_613,In_558);
or U923 (N_923,In_74,In_150);
and U924 (N_924,In_351,In_135);
nand U925 (N_925,In_334,In_374);
xor U926 (N_926,In_748,In_432);
nor U927 (N_927,In_450,In_41);
or U928 (N_928,In_351,In_391);
or U929 (N_929,In_311,In_447);
nand U930 (N_930,In_322,In_193);
nor U931 (N_931,In_582,In_684);
xnor U932 (N_932,In_305,In_711);
and U933 (N_933,In_658,In_228);
nand U934 (N_934,In_534,In_11);
nor U935 (N_935,In_55,In_357);
nor U936 (N_936,In_606,In_543);
xnor U937 (N_937,In_309,In_295);
nor U938 (N_938,In_57,In_492);
xnor U939 (N_939,In_587,In_125);
or U940 (N_940,In_331,In_267);
nor U941 (N_941,In_705,In_650);
nand U942 (N_942,In_333,In_635);
nand U943 (N_943,In_211,In_449);
xnor U944 (N_944,In_511,In_736);
nor U945 (N_945,In_204,In_473);
nor U946 (N_946,In_105,In_217);
nand U947 (N_947,In_334,In_619);
nand U948 (N_948,In_196,In_17);
xor U949 (N_949,In_353,In_485);
nor U950 (N_950,In_699,In_371);
xnor U951 (N_951,In_10,In_459);
xnor U952 (N_952,In_250,In_235);
nand U953 (N_953,In_499,In_623);
or U954 (N_954,In_176,In_97);
nor U955 (N_955,In_248,In_574);
xor U956 (N_956,In_634,In_303);
nand U957 (N_957,In_106,In_740);
or U958 (N_958,In_307,In_650);
and U959 (N_959,In_644,In_657);
and U960 (N_960,In_235,In_391);
nor U961 (N_961,In_172,In_311);
nor U962 (N_962,In_749,In_688);
and U963 (N_963,In_409,In_707);
xor U964 (N_964,In_499,In_537);
nor U965 (N_965,In_747,In_576);
or U966 (N_966,In_514,In_254);
xor U967 (N_967,In_687,In_439);
or U968 (N_968,In_412,In_74);
and U969 (N_969,In_199,In_643);
nand U970 (N_970,In_526,In_307);
or U971 (N_971,In_441,In_453);
nor U972 (N_972,In_287,In_4);
nor U973 (N_973,In_654,In_584);
xnor U974 (N_974,In_362,In_663);
or U975 (N_975,In_339,In_572);
nand U976 (N_976,In_202,In_615);
or U977 (N_977,In_80,In_58);
and U978 (N_978,In_337,In_49);
or U979 (N_979,In_479,In_382);
and U980 (N_980,In_512,In_604);
nand U981 (N_981,In_221,In_465);
xnor U982 (N_982,In_389,In_22);
nand U983 (N_983,In_683,In_299);
xor U984 (N_984,In_7,In_4);
xnor U985 (N_985,In_715,In_190);
xnor U986 (N_986,In_253,In_519);
nand U987 (N_987,In_246,In_489);
xnor U988 (N_988,In_49,In_474);
nand U989 (N_989,In_13,In_704);
nor U990 (N_990,In_99,In_0);
or U991 (N_991,In_97,In_453);
or U992 (N_992,In_397,In_600);
nand U993 (N_993,In_3,In_315);
and U994 (N_994,In_228,In_719);
nor U995 (N_995,In_142,In_452);
nor U996 (N_996,In_185,In_348);
nand U997 (N_997,In_521,In_520);
or U998 (N_998,In_582,In_150);
and U999 (N_999,In_715,In_697);
nand U1000 (N_1000,N_46,N_635);
nor U1001 (N_1001,N_947,N_442);
nor U1002 (N_1002,N_272,N_330);
nand U1003 (N_1003,N_132,N_350);
nand U1004 (N_1004,N_900,N_924);
nor U1005 (N_1005,N_627,N_555);
or U1006 (N_1006,N_3,N_233);
or U1007 (N_1007,N_164,N_224);
nor U1008 (N_1008,N_691,N_539);
nand U1009 (N_1009,N_389,N_798);
and U1010 (N_1010,N_421,N_343);
or U1011 (N_1011,N_835,N_60);
xnor U1012 (N_1012,N_746,N_415);
and U1013 (N_1013,N_865,N_206);
nand U1014 (N_1014,N_55,N_657);
and U1015 (N_1015,N_459,N_834);
and U1016 (N_1016,N_198,N_280);
and U1017 (N_1017,N_916,N_688);
nor U1018 (N_1018,N_370,N_252);
or U1019 (N_1019,N_884,N_380);
and U1020 (N_1020,N_180,N_679);
nor U1021 (N_1021,N_148,N_464);
xor U1022 (N_1022,N_583,N_636);
and U1023 (N_1023,N_931,N_446);
nand U1024 (N_1024,N_376,N_122);
and U1025 (N_1025,N_162,N_830);
and U1026 (N_1026,N_845,N_215);
and U1027 (N_1027,N_611,N_396);
and U1028 (N_1028,N_126,N_155);
nor U1029 (N_1029,N_800,N_142);
and U1030 (N_1030,N_842,N_293);
nor U1031 (N_1031,N_944,N_456);
xnor U1032 (N_1032,N_129,N_500);
or U1033 (N_1033,N_922,N_153);
or U1034 (N_1034,N_738,N_868);
or U1035 (N_1035,N_656,N_686);
nor U1036 (N_1036,N_440,N_581);
nor U1037 (N_1037,N_196,N_239);
nor U1038 (N_1038,N_347,N_402);
nor U1039 (N_1039,N_466,N_386);
or U1040 (N_1040,N_664,N_538);
and U1041 (N_1041,N_905,N_86);
xor U1042 (N_1042,N_369,N_474);
and U1043 (N_1043,N_625,N_600);
or U1044 (N_1044,N_10,N_626);
nand U1045 (N_1045,N_286,N_229);
and U1046 (N_1046,N_751,N_308);
nand U1047 (N_1047,N_222,N_297);
nand U1048 (N_1048,N_225,N_195);
nor U1049 (N_1049,N_57,N_431);
nor U1050 (N_1050,N_313,N_384);
xor U1051 (N_1051,N_356,N_712);
xnor U1052 (N_1052,N_217,N_56);
nor U1053 (N_1053,N_317,N_91);
or U1054 (N_1054,N_84,N_183);
xor U1055 (N_1055,N_346,N_698);
xnor U1056 (N_1056,N_75,N_913);
xnor U1057 (N_1057,N_750,N_536);
or U1058 (N_1058,N_78,N_637);
nand U1059 (N_1059,N_27,N_899);
nand U1060 (N_1060,N_99,N_933);
and U1061 (N_1061,N_266,N_717);
and U1062 (N_1062,N_935,N_364);
nand U1063 (N_1063,N_392,N_146);
or U1064 (N_1064,N_400,N_687);
nor U1065 (N_1065,N_508,N_173);
xor U1066 (N_1066,N_537,N_274);
and U1067 (N_1067,N_952,N_878);
or U1068 (N_1068,N_739,N_966);
nor U1069 (N_1069,N_486,N_200);
xor U1070 (N_1070,N_190,N_377);
or U1071 (N_1071,N_619,N_33);
nor U1072 (N_1072,N_419,N_136);
xor U1073 (N_1073,N_475,N_320);
and U1074 (N_1074,N_919,N_938);
nand U1075 (N_1075,N_915,N_765);
or U1076 (N_1076,N_478,N_490);
nand U1077 (N_1077,N_673,N_325);
and U1078 (N_1078,N_454,N_862);
xor U1079 (N_1079,N_177,N_911);
xor U1080 (N_1080,N_199,N_801);
xnor U1081 (N_1081,N_340,N_453);
xor U1082 (N_1082,N_826,N_125);
and U1083 (N_1083,N_113,N_850);
xnor U1084 (N_1084,N_609,N_836);
xnor U1085 (N_1085,N_394,N_816);
nand U1086 (N_1086,N_398,N_886);
nor U1087 (N_1087,N_560,N_957);
or U1088 (N_1088,N_334,N_448);
nor U1089 (N_1089,N_964,N_22);
xnor U1090 (N_1090,N_852,N_734);
nand U1091 (N_1091,N_928,N_268);
xnor U1092 (N_1092,N_974,N_759);
or U1093 (N_1093,N_288,N_283);
xnor U1094 (N_1094,N_418,N_708);
nand U1095 (N_1095,N_832,N_769);
and U1096 (N_1096,N_417,N_458);
and U1097 (N_1097,N_624,N_169);
nor U1098 (N_1098,N_485,N_756);
and U1099 (N_1099,N_871,N_940);
and U1100 (N_1100,N_178,N_117);
or U1101 (N_1101,N_408,N_705);
nor U1102 (N_1102,N_445,N_322);
xor U1103 (N_1103,N_6,N_156);
or U1104 (N_1104,N_110,N_867);
nand U1105 (N_1105,N_306,N_773);
or U1106 (N_1106,N_41,N_812);
nand U1107 (N_1107,N_427,N_405);
or U1108 (N_1108,N_279,N_715);
nand U1109 (N_1109,N_608,N_888);
nand U1110 (N_1110,N_647,N_336);
xnor U1111 (N_1111,N_690,N_477);
nor U1112 (N_1112,N_425,N_988);
and U1113 (N_1113,N_612,N_668);
or U1114 (N_1114,N_105,N_666);
xor U1115 (N_1115,N_585,N_163);
nand U1116 (N_1116,N_228,N_589);
and U1117 (N_1117,N_365,N_783);
nor U1118 (N_1118,N_315,N_861);
nor U1119 (N_1119,N_559,N_391);
xnor U1120 (N_1120,N_923,N_753);
or U1121 (N_1121,N_643,N_806);
and U1122 (N_1122,N_603,N_363);
or U1123 (N_1123,N_81,N_532);
and U1124 (N_1124,N_423,N_997);
nand U1125 (N_1125,N_621,N_790);
or U1126 (N_1126,N_482,N_604);
nand U1127 (N_1127,N_287,N_497);
and U1128 (N_1128,N_502,N_106);
or U1129 (N_1129,N_259,N_109);
or U1130 (N_1130,N_28,N_985);
and U1131 (N_1131,N_282,N_702);
and U1132 (N_1132,N_975,N_260);
nor U1133 (N_1133,N_675,N_755);
xor U1134 (N_1134,N_709,N_145);
or U1135 (N_1135,N_158,N_362);
nor U1136 (N_1136,N_186,N_713);
nor U1137 (N_1137,N_669,N_171);
xor U1138 (N_1138,N_0,N_236);
and U1139 (N_1139,N_776,N_614);
and U1140 (N_1140,N_823,N_662);
and U1141 (N_1141,N_566,N_891);
xnor U1142 (N_1142,N_367,N_332);
nand U1143 (N_1143,N_847,N_700);
nand U1144 (N_1144,N_978,N_789);
xor U1145 (N_1145,N_23,N_311);
and U1146 (N_1146,N_525,N_455);
nor U1147 (N_1147,N_895,N_295);
xor U1148 (N_1148,N_472,N_552);
and U1149 (N_1149,N_616,N_1);
xnor U1150 (N_1150,N_920,N_925);
nor U1151 (N_1151,N_615,N_275);
nand U1152 (N_1152,N_617,N_694);
nor U1153 (N_1153,N_981,N_395);
or U1154 (N_1154,N_413,N_192);
nor U1155 (N_1155,N_889,N_810);
nor U1156 (N_1156,N_52,N_121);
nand U1157 (N_1157,N_660,N_159);
and U1158 (N_1158,N_493,N_735);
and U1159 (N_1159,N_98,N_452);
or U1160 (N_1160,N_752,N_214);
or U1161 (N_1161,N_557,N_563);
nor U1162 (N_1162,N_593,N_761);
and U1163 (N_1163,N_181,N_299);
or U1164 (N_1164,N_729,N_654);
or U1165 (N_1165,N_963,N_794);
xor U1166 (N_1166,N_529,N_646);
and U1167 (N_1167,N_762,N_201);
xnor U1168 (N_1168,N_914,N_212);
nand U1169 (N_1169,N_469,N_953);
nor U1170 (N_1170,N_207,N_590);
xnor U1171 (N_1171,N_726,N_831);
nor U1172 (N_1172,N_620,N_528);
nor U1173 (N_1173,N_820,N_242);
xnor U1174 (N_1174,N_489,N_904);
xnor U1175 (N_1175,N_727,N_586);
nand U1176 (N_1176,N_788,N_618);
and U1177 (N_1177,N_167,N_813);
nand U1178 (N_1178,N_986,N_235);
nor U1179 (N_1179,N_663,N_4);
nand U1180 (N_1180,N_166,N_674);
nand U1181 (N_1181,N_987,N_141);
nand U1182 (N_1182,N_232,N_79);
xor U1183 (N_1183,N_994,N_331);
xor U1184 (N_1184,N_504,N_373);
nor U1185 (N_1185,N_689,N_917);
nor U1186 (N_1186,N_246,N_594);
or U1187 (N_1187,N_284,N_730);
nor U1188 (N_1188,N_292,N_574);
xor U1189 (N_1189,N_378,N_111);
and U1190 (N_1190,N_747,N_152);
nor U1191 (N_1191,N_678,N_337);
and U1192 (N_1192,N_573,N_64);
nand U1193 (N_1193,N_515,N_95);
nor U1194 (N_1194,N_18,N_443);
nor U1195 (N_1195,N_19,N_87);
and U1196 (N_1196,N_855,N_348);
xnor U1197 (N_1197,N_21,N_194);
and U1198 (N_1198,N_32,N_345);
and U1199 (N_1199,N_704,N_307);
xnor U1200 (N_1200,N_818,N_366);
and U1201 (N_1201,N_409,N_172);
and U1202 (N_1202,N_226,N_932);
nor U1203 (N_1203,N_736,N_516);
nor U1204 (N_1204,N_843,N_447);
or U1205 (N_1205,N_498,N_541);
xor U1206 (N_1206,N_771,N_805);
xor U1207 (N_1207,N_133,N_602);
and U1208 (N_1208,N_896,N_351);
nor U1209 (N_1209,N_718,N_219);
nor U1210 (N_1210,N_333,N_969);
nor U1211 (N_1211,N_197,N_781);
nand U1212 (N_1212,N_505,N_856);
xor U1213 (N_1213,N_534,N_150);
nand U1214 (N_1214,N_587,N_564);
or U1215 (N_1215,N_846,N_758);
and U1216 (N_1216,N_467,N_520);
and U1217 (N_1217,N_303,N_5);
and U1218 (N_1218,N_639,N_606);
nor U1219 (N_1219,N_763,N_680);
nand U1220 (N_1220,N_770,N_271);
xnor U1221 (N_1221,N_123,N_841);
nand U1222 (N_1222,N_630,N_184);
nor U1223 (N_1223,N_115,N_745);
xor U1224 (N_1224,N_909,N_479);
or U1225 (N_1225,N_906,N_149);
nand U1226 (N_1226,N_393,N_213);
or U1227 (N_1227,N_278,N_772);
xor U1228 (N_1228,N_744,N_607);
xnor U1229 (N_1229,N_848,N_277);
nand U1230 (N_1230,N_576,N_30);
or U1231 (N_1231,N_48,N_410);
nand U1232 (N_1232,N_96,N_995);
and U1233 (N_1233,N_494,N_645);
nand U1234 (N_1234,N_558,N_492);
nor U1235 (N_1235,N_706,N_483);
or U1236 (N_1236,N_261,N_210);
or U1237 (N_1237,N_468,N_665);
and U1238 (N_1238,N_872,N_480);
xnor U1239 (N_1239,N_926,N_894);
and U1240 (N_1240,N_359,N_305);
xor U1241 (N_1241,N_962,N_73);
nand U1242 (N_1242,N_316,N_294);
nor U1243 (N_1243,N_991,N_821);
nor U1244 (N_1244,N_154,N_866);
and U1245 (N_1245,N_354,N_601);
nand U1246 (N_1246,N_707,N_556);
nor U1247 (N_1247,N_757,N_36);
xor U1248 (N_1248,N_103,N_509);
or U1249 (N_1249,N_329,N_451);
or U1250 (N_1250,N_774,N_677);
nor U1251 (N_1251,N_649,N_24);
xnor U1252 (N_1252,N_561,N_53);
xor U1253 (N_1253,N_102,N_240);
xnor U1254 (N_1254,N_94,N_12);
or U1255 (N_1255,N_631,N_439);
xor U1256 (N_1256,N_642,N_39);
or U1257 (N_1257,N_2,N_910);
and U1258 (N_1258,N_179,N_716);
and U1259 (N_1259,N_151,N_732);
nand U1260 (N_1260,N_265,N_858);
or U1261 (N_1261,N_959,N_51);
nor U1262 (N_1262,N_724,N_465);
and U1263 (N_1263,N_319,N_946);
or U1264 (N_1264,N_257,N_681);
or U1265 (N_1265,N_484,N_877);
and U1266 (N_1266,N_281,N_353);
or U1267 (N_1267,N_754,N_107);
xor U1268 (N_1268,N_428,N_569);
nand U1269 (N_1269,N_811,N_571);
nor U1270 (N_1270,N_50,N_720);
nand U1271 (N_1271,N_85,N_548);
xor U1272 (N_1272,N_567,N_499);
or U1273 (N_1273,N_839,N_941);
nand U1274 (N_1274,N_628,N_450);
or U1275 (N_1275,N_513,N_591);
xnor U1276 (N_1276,N_870,N_565);
or U1277 (N_1277,N_787,N_887);
nor U1278 (N_1278,N_175,N_535);
and U1279 (N_1279,N_289,N_339);
xor U1280 (N_1280,N_936,N_92);
or U1281 (N_1281,N_385,N_245);
nor U1282 (N_1282,N_542,N_651);
nand U1283 (N_1283,N_244,N_948);
xnor U1284 (N_1284,N_815,N_568);
nand U1285 (N_1285,N_420,N_945);
or U1286 (N_1286,N_989,N_824);
xnor U1287 (N_1287,N_89,N_227);
nand U1288 (N_1288,N_728,N_863);
nand U1289 (N_1289,N_360,N_929);
and U1290 (N_1290,N_785,N_444);
nor U1291 (N_1291,N_661,N_135);
nand U1292 (N_1292,N_634,N_797);
nand U1293 (N_1293,N_851,N_838);
nand U1294 (N_1294,N_971,N_840);
nand U1295 (N_1295,N_633,N_312);
xnor U1296 (N_1296,N_640,N_723);
and U1297 (N_1297,N_880,N_550);
or U1298 (N_1298,N_209,N_131);
nor U1299 (N_1299,N_481,N_791);
nor U1300 (N_1300,N_216,N_66);
nor U1301 (N_1301,N_967,N_208);
nand U1302 (N_1302,N_983,N_328);
nor U1303 (N_1303,N_503,N_185);
nand U1304 (N_1304,N_270,N_290);
nand U1305 (N_1305,N_854,N_368);
nor U1306 (N_1306,N_203,N_890);
and U1307 (N_1307,N_249,N_780);
xor U1308 (N_1308,N_438,N_83);
and U1309 (N_1309,N_432,N_42);
xor U1310 (N_1310,N_338,N_580);
or U1311 (N_1311,N_379,N_956);
and U1312 (N_1312,N_97,N_256);
nor U1313 (N_1313,N_908,N_323);
nor U1314 (N_1314,N_531,N_300);
and U1315 (N_1315,N_719,N_588);
or U1316 (N_1316,N_255,N_999);
nand U1317 (N_1317,N_934,N_976);
and U1318 (N_1318,N_74,N_114);
nor U1319 (N_1319,N_685,N_683);
xnor U1320 (N_1320,N_374,N_701);
nand U1321 (N_1321,N_61,N_523);
and U1322 (N_1322,N_375,N_958);
nand U1323 (N_1323,N_864,N_309);
nor U1324 (N_1324,N_9,N_961);
nor U1325 (N_1325,N_189,N_80);
nor U1326 (N_1326,N_488,N_157);
or U1327 (N_1327,N_128,N_766);
xor U1328 (N_1328,N_460,N_161);
nand U1329 (N_1329,N_285,N_549);
nor U1330 (N_1330,N_301,N_692);
and U1331 (N_1331,N_584,N_572);
nor U1332 (N_1332,N_112,N_204);
xnor U1333 (N_1333,N_814,N_29);
and U1334 (N_1334,N_786,N_422);
or U1335 (N_1335,N_258,N_44);
xnor U1336 (N_1336,N_247,N_116);
nand U1337 (N_1337,N_104,N_387);
xnor U1338 (N_1338,N_551,N_424);
nor U1339 (N_1339,N_623,N_596);
and U1340 (N_1340,N_613,N_950);
and U1341 (N_1341,N_998,N_960);
and U1342 (N_1342,N_127,N_314);
xnor U1343 (N_1343,N_828,N_696);
nor U1344 (N_1344,N_599,N_760);
xor U1345 (N_1345,N_433,N_38);
nor U1346 (N_1346,N_598,N_276);
xor U1347 (N_1347,N_349,N_530);
nand U1348 (N_1348,N_837,N_737);
nor U1349 (N_1349,N_965,N_461);
nor U1350 (N_1350,N_388,N_462);
nand U1351 (N_1351,N_970,N_7);
or U1352 (N_1352,N_34,N_120);
xnor U1353 (N_1353,N_658,N_11);
nor U1354 (N_1354,N_907,N_491);
nand U1355 (N_1355,N_638,N_648);
xnor U1356 (N_1356,N_90,N_912);
xnor U1357 (N_1357,N_243,N_218);
nor U1358 (N_1358,N_223,N_412);
xor U1359 (N_1359,N_230,N_429);
or U1360 (N_1360,N_533,N_951);
or U1361 (N_1361,N_100,N_108);
xor U1362 (N_1362,N_65,N_361);
xnor U1363 (N_1363,N_76,N_982);
and U1364 (N_1364,N_250,N_984);
or U1365 (N_1365,N_802,N_143);
xor U1366 (N_1366,N_799,N_968);
nor U1367 (N_1367,N_202,N_733);
xnor U1368 (N_1368,N_344,N_434);
xnor U1369 (N_1369,N_544,N_833);
nand U1370 (N_1370,N_859,N_426);
and U1371 (N_1371,N_205,N_942);
or U1372 (N_1372,N_372,N_578);
nand U1373 (N_1373,N_653,N_546);
or U1374 (N_1374,N_68,N_874);
xnor U1375 (N_1375,N_355,N_807);
nor U1376 (N_1376,N_174,N_82);
xor U1377 (N_1377,N_191,N_775);
nor U1378 (N_1378,N_436,N_416);
or U1379 (N_1379,N_804,N_939);
nor U1380 (N_1380,N_595,N_570);
nor U1381 (N_1381,N_321,N_873);
nand U1382 (N_1382,N_43,N_514);
and U1383 (N_1383,N_629,N_844);
nand U1384 (N_1384,N_435,N_411);
and U1385 (N_1385,N_902,N_193);
xnor U1386 (N_1386,N_803,N_238);
nor U1387 (N_1387,N_262,N_672);
xor U1388 (N_1388,N_139,N_211);
or U1389 (N_1389,N_695,N_597);
or U1390 (N_1390,N_40,N_954);
xor U1391 (N_1391,N_487,N_977);
xor U1392 (N_1392,N_881,N_809);
nor U1393 (N_1393,N_949,N_170);
nor U1394 (N_1394,N_298,N_575);
and U1395 (N_1395,N_993,N_918);
nand U1396 (N_1396,N_93,N_31);
and U1397 (N_1397,N_682,N_693);
and U1398 (N_1398,N_898,N_140);
and U1399 (N_1399,N_883,N_722);
and U1400 (N_1400,N_699,N_16);
or U1401 (N_1401,N_793,N_980);
xor U1402 (N_1402,N_784,N_441);
or U1403 (N_1403,N_15,N_187);
nor U1404 (N_1404,N_930,N_511);
or U1405 (N_1405,N_8,N_20);
xnor U1406 (N_1406,N_644,N_562);
nand U1407 (N_1407,N_822,N_554);
and U1408 (N_1408,N_901,N_540);
nand U1409 (N_1409,N_71,N_437);
and U1410 (N_1410,N_341,N_518);
and U1411 (N_1411,N_748,N_955);
and U1412 (N_1412,N_582,N_470);
or U1413 (N_1413,N_296,N_13);
and U1414 (N_1414,N_937,N_670);
nor U1415 (N_1415,N_547,N_35);
or U1416 (N_1416,N_605,N_69);
nor U1417 (N_1417,N_371,N_49);
or U1418 (N_1418,N_324,N_326);
nand U1419 (N_1419,N_742,N_857);
nand U1420 (N_1420,N_510,N_404);
or U1421 (N_1421,N_973,N_545);
nor U1422 (N_1422,N_383,N_382);
and U1423 (N_1423,N_676,N_269);
nor U1424 (N_1424,N_253,N_342);
nor U1425 (N_1425,N_168,N_471);
or U1426 (N_1426,N_77,N_592);
nor U1427 (N_1427,N_782,N_519);
nand U1428 (N_1428,N_463,N_496);
xor U1429 (N_1429,N_652,N_767);
xnor U1430 (N_1430,N_327,N_241);
nand U1431 (N_1431,N_248,N_819);
and U1432 (N_1432,N_990,N_796);
or U1433 (N_1433,N_358,N_495);
xor U1434 (N_1434,N_579,N_251);
and U1435 (N_1435,N_473,N_263);
or U1436 (N_1436,N_72,N_543);
xor U1437 (N_1437,N_352,N_632);
or U1438 (N_1438,N_273,N_414);
or U1439 (N_1439,N_817,N_524);
nor U1440 (N_1440,N_119,N_47);
xor U1441 (N_1441,N_875,N_138);
nor U1442 (N_1442,N_893,N_725);
nor U1443 (N_1443,N_808,N_684);
nand U1444 (N_1444,N_45,N_318);
nand U1445 (N_1445,N_650,N_972);
or U1446 (N_1446,N_610,N_144);
and U1447 (N_1447,N_903,N_449);
nor U1448 (N_1448,N_622,N_892);
xnor U1449 (N_1449,N_130,N_743);
or U1450 (N_1450,N_527,N_740);
or U1451 (N_1451,N_231,N_943);
and U1452 (N_1452,N_26,N_234);
nor U1453 (N_1453,N_302,N_58);
and U1454 (N_1454,N_67,N_710);
or U1455 (N_1455,N_667,N_147);
or U1456 (N_1456,N_927,N_778);
and U1457 (N_1457,N_876,N_777);
nand U1458 (N_1458,N_749,N_476);
nand U1459 (N_1459,N_335,N_517);
xor U1460 (N_1460,N_176,N_827);
nand U1461 (N_1461,N_731,N_671);
or U1462 (N_1462,N_897,N_267);
and U1463 (N_1463,N_992,N_304);
xor U1464 (N_1464,N_521,N_407);
or U1465 (N_1465,N_577,N_137);
nor U1466 (N_1466,N_768,N_860);
and U1467 (N_1467,N_711,N_403);
and U1468 (N_1468,N_882,N_221);
xor U1469 (N_1469,N_291,N_641);
xnor U1470 (N_1470,N_921,N_220);
nand U1471 (N_1471,N_697,N_54);
and U1472 (N_1472,N_996,N_512);
nor U1473 (N_1473,N_17,N_655);
or U1474 (N_1474,N_390,N_714);
and U1475 (N_1475,N_795,N_979);
nor U1476 (N_1476,N_703,N_310);
xor U1477 (N_1477,N_507,N_825);
or U1478 (N_1478,N_188,N_829);
xor U1479 (N_1479,N_124,N_553);
nor U1480 (N_1480,N_381,N_182);
and U1481 (N_1481,N_522,N_62);
and U1482 (N_1482,N_406,N_63);
nor U1483 (N_1483,N_399,N_101);
xnor U1484 (N_1484,N_501,N_134);
and U1485 (N_1485,N_118,N_506);
or U1486 (N_1486,N_659,N_397);
and U1487 (N_1487,N_457,N_37);
xnor U1488 (N_1488,N_237,N_779);
nand U1489 (N_1489,N_25,N_741);
xnor U1490 (N_1490,N_869,N_14);
and U1491 (N_1491,N_70,N_401);
nor U1492 (N_1492,N_764,N_165);
nor U1493 (N_1493,N_357,N_792);
and U1494 (N_1494,N_849,N_430);
xnor U1495 (N_1495,N_88,N_853);
nor U1496 (N_1496,N_264,N_160);
nand U1497 (N_1497,N_59,N_254);
and U1498 (N_1498,N_879,N_721);
and U1499 (N_1499,N_526,N_885);
or U1500 (N_1500,N_925,N_627);
nor U1501 (N_1501,N_786,N_864);
nand U1502 (N_1502,N_927,N_631);
nand U1503 (N_1503,N_405,N_671);
and U1504 (N_1504,N_966,N_875);
and U1505 (N_1505,N_136,N_548);
nand U1506 (N_1506,N_653,N_541);
and U1507 (N_1507,N_841,N_392);
and U1508 (N_1508,N_757,N_994);
nand U1509 (N_1509,N_143,N_160);
xnor U1510 (N_1510,N_115,N_789);
nand U1511 (N_1511,N_655,N_619);
nor U1512 (N_1512,N_727,N_801);
nor U1513 (N_1513,N_160,N_797);
xor U1514 (N_1514,N_225,N_334);
nand U1515 (N_1515,N_428,N_214);
nand U1516 (N_1516,N_491,N_138);
or U1517 (N_1517,N_92,N_601);
nand U1518 (N_1518,N_937,N_660);
nand U1519 (N_1519,N_325,N_494);
or U1520 (N_1520,N_600,N_542);
or U1521 (N_1521,N_317,N_132);
and U1522 (N_1522,N_391,N_501);
or U1523 (N_1523,N_136,N_244);
nor U1524 (N_1524,N_856,N_531);
nor U1525 (N_1525,N_13,N_526);
or U1526 (N_1526,N_691,N_351);
or U1527 (N_1527,N_98,N_47);
and U1528 (N_1528,N_935,N_831);
or U1529 (N_1529,N_952,N_802);
or U1530 (N_1530,N_958,N_550);
nor U1531 (N_1531,N_403,N_766);
or U1532 (N_1532,N_908,N_879);
nand U1533 (N_1533,N_126,N_242);
or U1534 (N_1534,N_46,N_736);
and U1535 (N_1535,N_476,N_136);
nand U1536 (N_1536,N_598,N_765);
xor U1537 (N_1537,N_881,N_883);
nor U1538 (N_1538,N_849,N_828);
nand U1539 (N_1539,N_334,N_840);
or U1540 (N_1540,N_564,N_265);
xnor U1541 (N_1541,N_972,N_96);
and U1542 (N_1542,N_80,N_368);
xnor U1543 (N_1543,N_723,N_71);
or U1544 (N_1544,N_205,N_202);
nor U1545 (N_1545,N_313,N_887);
nand U1546 (N_1546,N_561,N_337);
nor U1547 (N_1547,N_435,N_848);
and U1548 (N_1548,N_25,N_705);
or U1549 (N_1549,N_84,N_940);
and U1550 (N_1550,N_126,N_18);
nand U1551 (N_1551,N_1,N_634);
nor U1552 (N_1552,N_465,N_156);
nor U1553 (N_1553,N_912,N_80);
nor U1554 (N_1554,N_797,N_724);
nor U1555 (N_1555,N_639,N_142);
or U1556 (N_1556,N_419,N_281);
nand U1557 (N_1557,N_337,N_722);
or U1558 (N_1558,N_181,N_602);
xor U1559 (N_1559,N_358,N_769);
nand U1560 (N_1560,N_443,N_996);
xor U1561 (N_1561,N_323,N_569);
xor U1562 (N_1562,N_493,N_891);
or U1563 (N_1563,N_761,N_597);
nand U1564 (N_1564,N_89,N_356);
nand U1565 (N_1565,N_643,N_256);
nand U1566 (N_1566,N_237,N_987);
xor U1567 (N_1567,N_830,N_422);
nor U1568 (N_1568,N_167,N_101);
nand U1569 (N_1569,N_838,N_854);
or U1570 (N_1570,N_421,N_643);
xor U1571 (N_1571,N_641,N_926);
and U1572 (N_1572,N_881,N_138);
and U1573 (N_1573,N_587,N_669);
xnor U1574 (N_1574,N_108,N_762);
xnor U1575 (N_1575,N_352,N_242);
xnor U1576 (N_1576,N_920,N_943);
nand U1577 (N_1577,N_910,N_446);
nor U1578 (N_1578,N_505,N_838);
or U1579 (N_1579,N_204,N_392);
nor U1580 (N_1580,N_599,N_501);
xor U1581 (N_1581,N_364,N_620);
nor U1582 (N_1582,N_236,N_535);
nand U1583 (N_1583,N_760,N_24);
or U1584 (N_1584,N_366,N_99);
and U1585 (N_1585,N_5,N_886);
and U1586 (N_1586,N_614,N_400);
nand U1587 (N_1587,N_431,N_697);
nand U1588 (N_1588,N_673,N_810);
and U1589 (N_1589,N_28,N_744);
or U1590 (N_1590,N_75,N_541);
or U1591 (N_1591,N_198,N_210);
or U1592 (N_1592,N_466,N_556);
and U1593 (N_1593,N_572,N_181);
or U1594 (N_1594,N_285,N_401);
xor U1595 (N_1595,N_71,N_789);
xnor U1596 (N_1596,N_297,N_382);
and U1597 (N_1597,N_0,N_187);
nand U1598 (N_1598,N_854,N_379);
or U1599 (N_1599,N_586,N_166);
xnor U1600 (N_1600,N_310,N_719);
or U1601 (N_1601,N_223,N_453);
or U1602 (N_1602,N_786,N_167);
nand U1603 (N_1603,N_661,N_57);
or U1604 (N_1604,N_136,N_954);
and U1605 (N_1605,N_394,N_826);
nand U1606 (N_1606,N_545,N_855);
xnor U1607 (N_1607,N_970,N_649);
or U1608 (N_1608,N_616,N_69);
nor U1609 (N_1609,N_170,N_609);
or U1610 (N_1610,N_199,N_166);
nor U1611 (N_1611,N_943,N_559);
nand U1612 (N_1612,N_738,N_454);
or U1613 (N_1613,N_735,N_20);
nor U1614 (N_1614,N_640,N_866);
nand U1615 (N_1615,N_536,N_408);
nand U1616 (N_1616,N_702,N_102);
or U1617 (N_1617,N_425,N_711);
nand U1618 (N_1618,N_989,N_140);
nor U1619 (N_1619,N_244,N_549);
and U1620 (N_1620,N_927,N_575);
nand U1621 (N_1621,N_225,N_403);
and U1622 (N_1622,N_919,N_824);
and U1623 (N_1623,N_821,N_47);
or U1624 (N_1624,N_857,N_66);
nand U1625 (N_1625,N_772,N_23);
xor U1626 (N_1626,N_81,N_436);
nor U1627 (N_1627,N_315,N_956);
xnor U1628 (N_1628,N_561,N_991);
xnor U1629 (N_1629,N_495,N_97);
xor U1630 (N_1630,N_166,N_849);
nor U1631 (N_1631,N_106,N_820);
xor U1632 (N_1632,N_777,N_404);
nand U1633 (N_1633,N_680,N_90);
xnor U1634 (N_1634,N_890,N_324);
xnor U1635 (N_1635,N_661,N_888);
or U1636 (N_1636,N_744,N_221);
nor U1637 (N_1637,N_745,N_797);
and U1638 (N_1638,N_573,N_289);
xor U1639 (N_1639,N_243,N_503);
and U1640 (N_1640,N_471,N_290);
nand U1641 (N_1641,N_417,N_211);
nand U1642 (N_1642,N_206,N_455);
and U1643 (N_1643,N_989,N_481);
nand U1644 (N_1644,N_46,N_346);
nand U1645 (N_1645,N_652,N_120);
xor U1646 (N_1646,N_814,N_493);
nor U1647 (N_1647,N_515,N_974);
or U1648 (N_1648,N_757,N_16);
nor U1649 (N_1649,N_426,N_466);
nor U1650 (N_1650,N_491,N_610);
and U1651 (N_1651,N_360,N_182);
nand U1652 (N_1652,N_797,N_633);
nand U1653 (N_1653,N_129,N_478);
and U1654 (N_1654,N_960,N_873);
and U1655 (N_1655,N_201,N_168);
and U1656 (N_1656,N_187,N_526);
or U1657 (N_1657,N_103,N_680);
and U1658 (N_1658,N_109,N_0);
nand U1659 (N_1659,N_148,N_457);
and U1660 (N_1660,N_889,N_446);
xor U1661 (N_1661,N_763,N_734);
or U1662 (N_1662,N_826,N_870);
or U1663 (N_1663,N_954,N_91);
nor U1664 (N_1664,N_126,N_690);
xor U1665 (N_1665,N_681,N_678);
xnor U1666 (N_1666,N_332,N_456);
xnor U1667 (N_1667,N_190,N_233);
or U1668 (N_1668,N_586,N_955);
nand U1669 (N_1669,N_880,N_600);
or U1670 (N_1670,N_738,N_993);
nor U1671 (N_1671,N_693,N_259);
nor U1672 (N_1672,N_254,N_137);
or U1673 (N_1673,N_217,N_980);
or U1674 (N_1674,N_159,N_576);
nand U1675 (N_1675,N_116,N_306);
nand U1676 (N_1676,N_335,N_657);
xor U1677 (N_1677,N_844,N_956);
xnor U1678 (N_1678,N_613,N_744);
and U1679 (N_1679,N_571,N_517);
nor U1680 (N_1680,N_755,N_464);
nor U1681 (N_1681,N_780,N_184);
nand U1682 (N_1682,N_229,N_153);
nand U1683 (N_1683,N_554,N_955);
or U1684 (N_1684,N_979,N_425);
nand U1685 (N_1685,N_807,N_528);
xor U1686 (N_1686,N_904,N_919);
or U1687 (N_1687,N_249,N_96);
xor U1688 (N_1688,N_358,N_855);
or U1689 (N_1689,N_341,N_998);
nor U1690 (N_1690,N_899,N_215);
nor U1691 (N_1691,N_387,N_112);
or U1692 (N_1692,N_712,N_153);
and U1693 (N_1693,N_158,N_132);
nor U1694 (N_1694,N_208,N_345);
nor U1695 (N_1695,N_166,N_287);
or U1696 (N_1696,N_867,N_870);
xor U1697 (N_1697,N_495,N_469);
nor U1698 (N_1698,N_447,N_702);
nand U1699 (N_1699,N_200,N_766);
and U1700 (N_1700,N_573,N_655);
or U1701 (N_1701,N_391,N_377);
or U1702 (N_1702,N_211,N_152);
nor U1703 (N_1703,N_590,N_511);
xnor U1704 (N_1704,N_721,N_374);
nand U1705 (N_1705,N_228,N_928);
or U1706 (N_1706,N_910,N_707);
xnor U1707 (N_1707,N_241,N_788);
xnor U1708 (N_1708,N_706,N_764);
nand U1709 (N_1709,N_779,N_883);
xor U1710 (N_1710,N_555,N_111);
nand U1711 (N_1711,N_705,N_588);
and U1712 (N_1712,N_255,N_854);
or U1713 (N_1713,N_660,N_787);
and U1714 (N_1714,N_752,N_312);
and U1715 (N_1715,N_808,N_782);
or U1716 (N_1716,N_403,N_650);
xor U1717 (N_1717,N_6,N_500);
nand U1718 (N_1718,N_954,N_211);
and U1719 (N_1719,N_933,N_850);
xor U1720 (N_1720,N_338,N_552);
nor U1721 (N_1721,N_134,N_377);
nor U1722 (N_1722,N_572,N_58);
nand U1723 (N_1723,N_383,N_581);
and U1724 (N_1724,N_725,N_193);
nand U1725 (N_1725,N_422,N_582);
nor U1726 (N_1726,N_519,N_913);
nand U1727 (N_1727,N_495,N_317);
or U1728 (N_1728,N_858,N_304);
nand U1729 (N_1729,N_220,N_797);
nand U1730 (N_1730,N_125,N_130);
and U1731 (N_1731,N_873,N_869);
nand U1732 (N_1732,N_366,N_598);
and U1733 (N_1733,N_625,N_786);
nor U1734 (N_1734,N_635,N_807);
nand U1735 (N_1735,N_978,N_157);
nand U1736 (N_1736,N_84,N_990);
or U1737 (N_1737,N_308,N_113);
and U1738 (N_1738,N_730,N_181);
xor U1739 (N_1739,N_587,N_624);
or U1740 (N_1740,N_186,N_514);
nand U1741 (N_1741,N_661,N_458);
nor U1742 (N_1742,N_606,N_271);
xor U1743 (N_1743,N_271,N_56);
or U1744 (N_1744,N_342,N_795);
or U1745 (N_1745,N_301,N_893);
and U1746 (N_1746,N_844,N_359);
or U1747 (N_1747,N_522,N_868);
or U1748 (N_1748,N_89,N_754);
nor U1749 (N_1749,N_494,N_27);
nand U1750 (N_1750,N_670,N_634);
xnor U1751 (N_1751,N_242,N_521);
nor U1752 (N_1752,N_320,N_878);
nor U1753 (N_1753,N_373,N_908);
nor U1754 (N_1754,N_36,N_641);
or U1755 (N_1755,N_448,N_58);
or U1756 (N_1756,N_935,N_680);
nand U1757 (N_1757,N_3,N_273);
nand U1758 (N_1758,N_512,N_845);
nand U1759 (N_1759,N_876,N_993);
or U1760 (N_1760,N_485,N_504);
nor U1761 (N_1761,N_652,N_34);
nor U1762 (N_1762,N_1,N_842);
xor U1763 (N_1763,N_329,N_823);
nand U1764 (N_1764,N_418,N_182);
nor U1765 (N_1765,N_692,N_586);
nor U1766 (N_1766,N_374,N_376);
xor U1767 (N_1767,N_672,N_581);
nor U1768 (N_1768,N_30,N_950);
and U1769 (N_1769,N_305,N_264);
nor U1770 (N_1770,N_295,N_1);
nor U1771 (N_1771,N_683,N_71);
or U1772 (N_1772,N_309,N_689);
nor U1773 (N_1773,N_938,N_751);
xnor U1774 (N_1774,N_604,N_540);
or U1775 (N_1775,N_352,N_610);
and U1776 (N_1776,N_744,N_441);
and U1777 (N_1777,N_549,N_69);
and U1778 (N_1778,N_545,N_616);
or U1779 (N_1779,N_936,N_131);
nor U1780 (N_1780,N_653,N_319);
or U1781 (N_1781,N_624,N_316);
nor U1782 (N_1782,N_89,N_263);
nor U1783 (N_1783,N_571,N_432);
and U1784 (N_1784,N_60,N_207);
xnor U1785 (N_1785,N_487,N_998);
xor U1786 (N_1786,N_97,N_960);
and U1787 (N_1787,N_459,N_774);
nand U1788 (N_1788,N_219,N_917);
and U1789 (N_1789,N_982,N_985);
nand U1790 (N_1790,N_409,N_495);
xor U1791 (N_1791,N_861,N_712);
xor U1792 (N_1792,N_244,N_279);
nand U1793 (N_1793,N_40,N_66);
or U1794 (N_1794,N_547,N_954);
xor U1795 (N_1795,N_27,N_583);
nor U1796 (N_1796,N_459,N_596);
nor U1797 (N_1797,N_849,N_626);
xor U1798 (N_1798,N_357,N_136);
xnor U1799 (N_1799,N_697,N_732);
or U1800 (N_1800,N_391,N_562);
or U1801 (N_1801,N_347,N_16);
or U1802 (N_1802,N_529,N_553);
and U1803 (N_1803,N_50,N_740);
xnor U1804 (N_1804,N_862,N_284);
or U1805 (N_1805,N_385,N_664);
xnor U1806 (N_1806,N_40,N_22);
nand U1807 (N_1807,N_476,N_131);
xnor U1808 (N_1808,N_512,N_19);
xnor U1809 (N_1809,N_149,N_29);
and U1810 (N_1810,N_232,N_713);
or U1811 (N_1811,N_455,N_51);
xnor U1812 (N_1812,N_976,N_277);
nor U1813 (N_1813,N_574,N_392);
nand U1814 (N_1814,N_92,N_569);
or U1815 (N_1815,N_609,N_159);
xnor U1816 (N_1816,N_987,N_955);
or U1817 (N_1817,N_314,N_641);
and U1818 (N_1818,N_989,N_304);
and U1819 (N_1819,N_426,N_385);
or U1820 (N_1820,N_418,N_449);
nand U1821 (N_1821,N_932,N_584);
nand U1822 (N_1822,N_332,N_953);
xnor U1823 (N_1823,N_344,N_267);
or U1824 (N_1824,N_904,N_825);
xnor U1825 (N_1825,N_559,N_816);
xnor U1826 (N_1826,N_479,N_91);
xor U1827 (N_1827,N_854,N_667);
or U1828 (N_1828,N_589,N_331);
nor U1829 (N_1829,N_990,N_128);
or U1830 (N_1830,N_745,N_385);
nand U1831 (N_1831,N_765,N_689);
or U1832 (N_1832,N_449,N_729);
nand U1833 (N_1833,N_481,N_163);
nand U1834 (N_1834,N_242,N_790);
nor U1835 (N_1835,N_900,N_456);
and U1836 (N_1836,N_209,N_922);
or U1837 (N_1837,N_552,N_451);
nand U1838 (N_1838,N_936,N_57);
or U1839 (N_1839,N_30,N_292);
or U1840 (N_1840,N_769,N_817);
xor U1841 (N_1841,N_576,N_980);
and U1842 (N_1842,N_351,N_812);
or U1843 (N_1843,N_571,N_495);
nor U1844 (N_1844,N_171,N_200);
nand U1845 (N_1845,N_162,N_118);
nand U1846 (N_1846,N_365,N_382);
nand U1847 (N_1847,N_776,N_88);
nor U1848 (N_1848,N_250,N_205);
nand U1849 (N_1849,N_491,N_685);
nor U1850 (N_1850,N_880,N_109);
and U1851 (N_1851,N_977,N_761);
nand U1852 (N_1852,N_934,N_543);
or U1853 (N_1853,N_598,N_883);
nor U1854 (N_1854,N_723,N_749);
or U1855 (N_1855,N_541,N_440);
and U1856 (N_1856,N_667,N_884);
or U1857 (N_1857,N_491,N_392);
or U1858 (N_1858,N_358,N_598);
nor U1859 (N_1859,N_416,N_961);
nor U1860 (N_1860,N_89,N_917);
nor U1861 (N_1861,N_180,N_171);
nand U1862 (N_1862,N_821,N_956);
or U1863 (N_1863,N_110,N_522);
and U1864 (N_1864,N_228,N_744);
nand U1865 (N_1865,N_246,N_417);
nor U1866 (N_1866,N_380,N_532);
nor U1867 (N_1867,N_963,N_886);
or U1868 (N_1868,N_42,N_263);
nor U1869 (N_1869,N_572,N_286);
nor U1870 (N_1870,N_431,N_996);
nand U1871 (N_1871,N_528,N_297);
xnor U1872 (N_1872,N_551,N_995);
and U1873 (N_1873,N_670,N_3);
and U1874 (N_1874,N_327,N_753);
nand U1875 (N_1875,N_753,N_290);
xnor U1876 (N_1876,N_777,N_757);
nor U1877 (N_1877,N_523,N_768);
or U1878 (N_1878,N_581,N_770);
and U1879 (N_1879,N_497,N_597);
nand U1880 (N_1880,N_843,N_888);
or U1881 (N_1881,N_223,N_509);
xor U1882 (N_1882,N_223,N_685);
or U1883 (N_1883,N_487,N_943);
or U1884 (N_1884,N_213,N_830);
or U1885 (N_1885,N_322,N_806);
and U1886 (N_1886,N_861,N_797);
nand U1887 (N_1887,N_258,N_325);
or U1888 (N_1888,N_403,N_247);
and U1889 (N_1889,N_60,N_824);
and U1890 (N_1890,N_67,N_406);
nand U1891 (N_1891,N_657,N_23);
nor U1892 (N_1892,N_479,N_287);
and U1893 (N_1893,N_40,N_93);
nor U1894 (N_1894,N_877,N_631);
and U1895 (N_1895,N_747,N_971);
or U1896 (N_1896,N_48,N_977);
xnor U1897 (N_1897,N_300,N_902);
and U1898 (N_1898,N_835,N_439);
nand U1899 (N_1899,N_950,N_410);
nand U1900 (N_1900,N_917,N_98);
xor U1901 (N_1901,N_415,N_121);
xnor U1902 (N_1902,N_361,N_896);
nand U1903 (N_1903,N_974,N_308);
or U1904 (N_1904,N_357,N_335);
and U1905 (N_1905,N_737,N_238);
nor U1906 (N_1906,N_973,N_32);
and U1907 (N_1907,N_651,N_78);
and U1908 (N_1908,N_897,N_78);
or U1909 (N_1909,N_350,N_675);
or U1910 (N_1910,N_495,N_154);
and U1911 (N_1911,N_562,N_598);
or U1912 (N_1912,N_704,N_939);
nor U1913 (N_1913,N_56,N_123);
or U1914 (N_1914,N_81,N_823);
and U1915 (N_1915,N_722,N_654);
and U1916 (N_1916,N_385,N_117);
xor U1917 (N_1917,N_443,N_222);
or U1918 (N_1918,N_991,N_829);
nand U1919 (N_1919,N_187,N_377);
xnor U1920 (N_1920,N_70,N_19);
xnor U1921 (N_1921,N_182,N_226);
and U1922 (N_1922,N_254,N_919);
xnor U1923 (N_1923,N_677,N_651);
or U1924 (N_1924,N_539,N_35);
or U1925 (N_1925,N_263,N_803);
nand U1926 (N_1926,N_824,N_251);
xnor U1927 (N_1927,N_6,N_534);
nor U1928 (N_1928,N_246,N_274);
and U1929 (N_1929,N_935,N_720);
xor U1930 (N_1930,N_186,N_678);
or U1931 (N_1931,N_808,N_846);
xor U1932 (N_1932,N_432,N_528);
or U1933 (N_1933,N_746,N_946);
xor U1934 (N_1934,N_40,N_129);
nor U1935 (N_1935,N_815,N_453);
nand U1936 (N_1936,N_485,N_435);
and U1937 (N_1937,N_781,N_895);
nor U1938 (N_1938,N_394,N_324);
nor U1939 (N_1939,N_495,N_86);
or U1940 (N_1940,N_341,N_50);
and U1941 (N_1941,N_66,N_207);
xor U1942 (N_1942,N_590,N_37);
nand U1943 (N_1943,N_558,N_59);
and U1944 (N_1944,N_284,N_946);
nor U1945 (N_1945,N_911,N_316);
and U1946 (N_1946,N_997,N_584);
nand U1947 (N_1947,N_659,N_312);
or U1948 (N_1948,N_880,N_699);
and U1949 (N_1949,N_699,N_586);
nor U1950 (N_1950,N_128,N_504);
and U1951 (N_1951,N_721,N_403);
and U1952 (N_1952,N_239,N_121);
nor U1953 (N_1953,N_179,N_798);
nand U1954 (N_1954,N_502,N_117);
and U1955 (N_1955,N_763,N_945);
and U1956 (N_1956,N_938,N_17);
nor U1957 (N_1957,N_176,N_681);
xnor U1958 (N_1958,N_677,N_15);
or U1959 (N_1959,N_893,N_387);
nand U1960 (N_1960,N_598,N_89);
nand U1961 (N_1961,N_749,N_132);
nor U1962 (N_1962,N_966,N_414);
nor U1963 (N_1963,N_893,N_958);
and U1964 (N_1964,N_165,N_281);
nand U1965 (N_1965,N_131,N_747);
nor U1966 (N_1966,N_80,N_526);
nand U1967 (N_1967,N_356,N_785);
xnor U1968 (N_1968,N_188,N_642);
nand U1969 (N_1969,N_999,N_420);
xnor U1970 (N_1970,N_358,N_142);
nor U1971 (N_1971,N_869,N_970);
and U1972 (N_1972,N_351,N_964);
and U1973 (N_1973,N_660,N_939);
nor U1974 (N_1974,N_39,N_861);
nor U1975 (N_1975,N_587,N_886);
or U1976 (N_1976,N_833,N_575);
xor U1977 (N_1977,N_364,N_65);
nand U1978 (N_1978,N_989,N_453);
xnor U1979 (N_1979,N_704,N_488);
and U1980 (N_1980,N_694,N_997);
or U1981 (N_1981,N_436,N_521);
nor U1982 (N_1982,N_144,N_959);
and U1983 (N_1983,N_76,N_841);
or U1984 (N_1984,N_518,N_205);
nand U1985 (N_1985,N_531,N_814);
or U1986 (N_1986,N_342,N_814);
nor U1987 (N_1987,N_443,N_522);
nand U1988 (N_1988,N_132,N_566);
or U1989 (N_1989,N_755,N_895);
nand U1990 (N_1990,N_59,N_141);
and U1991 (N_1991,N_946,N_475);
nand U1992 (N_1992,N_98,N_729);
or U1993 (N_1993,N_457,N_816);
nor U1994 (N_1994,N_345,N_93);
nand U1995 (N_1995,N_877,N_537);
nand U1996 (N_1996,N_214,N_70);
nor U1997 (N_1997,N_669,N_783);
nor U1998 (N_1998,N_389,N_294);
and U1999 (N_1999,N_721,N_687);
or U2000 (N_2000,N_1962,N_1079);
and U2001 (N_2001,N_1842,N_1355);
nand U2002 (N_2002,N_1626,N_1811);
or U2003 (N_2003,N_1189,N_1571);
xnor U2004 (N_2004,N_1767,N_1375);
and U2005 (N_2005,N_1239,N_1966);
and U2006 (N_2006,N_1756,N_1337);
or U2007 (N_2007,N_1955,N_1059);
nor U2008 (N_2008,N_1875,N_1323);
xnor U2009 (N_2009,N_1096,N_1160);
xnor U2010 (N_2010,N_1789,N_1569);
or U2011 (N_2011,N_1070,N_1702);
nor U2012 (N_2012,N_1975,N_1991);
nand U2013 (N_2013,N_1914,N_1940);
or U2014 (N_2014,N_1572,N_1827);
xor U2015 (N_2015,N_1683,N_1410);
and U2016 (N_2016,N_1293,N_1573);
xor U2017 (N_2017,N_1530,N_1656);
nor U2018 (N_2018,N_1093,N_1772);
xnor U2019 (N_2019,N_1603,N_1556);
nand U2020 (N_2020,N_1668,N_1947);
nor U2021 (N_2021,N_1590,N_1317);
and U2022 (N_2022,N_1432,N_1696);
and U2023 (N_2023,N_1402,N_1779);
nor U2024 (N_2024,N_1716,N_1318);
or U2025 (N_2025,N_1970,N_1983);
xor U2026 (N_2026,N_1340,N_1253);
xnor U2027 (N_2027,N_1594,N_1254);
nor U2028 (N_2028,N_1431,N_1113);
and U2029 (N_2029,N_1188,N_1926);
xnor U2030 (N_2030,N_1904,N_1047);
nand U2031 (N_2031,N_1846,N_1880);
nand U2032 (N_2032,N_1540,N_1619);
and U2033 (N_2033,N_1324,N_1841);
xnor U2034 (N_2034,N_1497,N_1061);
xnor U2035 (N_2035,N_1416,N_1051);
and U2036 (N_2036,N_1479,N_1447);
nor U2037 (N_2037,N_1934,N_1232);
xor U2038 (N_2038,N_1197,N_1622);
nand U2039 (N_2039,N_1660,N_1397);
or U2040 (N_2040,N_1374,N_1555);
nand U2041 (N_2041,N_1194,N_1078);
and U2042 (N_2042,N_1316,N_1993);
or U2043 (N_2043,N_1033,N_1972);
and U2044 (N_2044,N_1272,N_1579);
or U2045 (N_2045,N_1399,N_1215);
and U2046 (N_2046,N_1528,N_1210);
and U2047 (N_2047,N_1670,N_1029);
and U2048 (N_2048,N_1167,N_1109);
xnor U2049 (N_2049,N_1040,N_1710);
nand U2050 (N_2050,N_1472,N_1786);
or U2051 (N_2051,N_1110,N_1884);
nand U2052 (N_2052,N_1956,N_1417);
nor U2053 (N_2053,N_1627,N_1192);
nor U2054 (N_2054,N_1299,N_1055);
nor U2055 (N_2055,N_1149,N_1831);
nand U2056 (N_2056,N_1730,N_1224);
nand U2057 (N_2057,N_1435,N_1760);
xnor U2058 (N_2058,N_1478,N_1689);
nand U2059 (N_2059,N_1283,N_1180);
nand U2060 (N_2060,N_1761,N_1373);
nor U2061 (N_2061,N_1853,N_1607);
nor U2062 (N_2062,N_1837,N_1644);
xor U2063 (N_2063,N_1217,N_1143);
or U2064 (N_2064,N_1963,N_1502);
or U2065 (N_2065,N_1225,N_1064);
or U2066 (N_2066,N_1581,N_1218);
xor U2067 (N_2067,N_1279,N_1521);
xnor U2068 (N_2068,N_1680,N_1146);
and U2069 (N_2069,N_1771,N_1357);
xnor U2070 (N_2070,N_1000,N_1764);
xor U2071 (N_2071,N_1142,N_1383);
and U2072 (N_2072,N_1558,N_1231);
nor U2073 (N_2073,N_1861,N_1129);
xnor U2074 (N_2074,N_1288,N_1939);
xnor U2075 (N_2075,N_1102,N_1511);
xor U2076 (N_2076,N_1200,N_1412);
nand U2077 (N_2077,N_1913,N_1049);
nor U2078 (N_2078,N_1004,N_1437);
or U2079 (N_2079,N_1308,N_1025);
and U2080 (N_2080,N_1698,N_1862);
nor U2081 (N_2081,N_1931,N_1953);
and U2082 (N_2082,N_1128,N_1929);
or U2083 (N_2083,N_1672,N_1391);
or U2084 (N_2084,N_1264,N_1669);
or U2085 (N_2085,N_1041,N_1695);
nand U2086 (N_2086,N_1867,N_1667);
nor U2087 (N_2087,N_1038,N_1507);
xor U2088 (N_2088,N_1274,N_1851);
nor U2089 (N_2089,N_1836,N_1957);
or U2090 (N_2090,N_1759,N_1312);
and U2091 (N_2091,N_1099,N_1276);
xor U2092 (N_2092,N_1723,N_1858);
nand U2093 (N_2093,N_1780,N_1612);
xor U2094 (N_2094,N_1782,N_1944);
xor U2095 (N_2095,N_1291,N_1985);
and U2096 (N_2096,N_1671,N_1525);
and U2097 (N_2097,N_1635,N_1187);
xor U2098 (N_2098,N_1908,N_1817);
or U2099 (N_2099,N_1075,N_1788);
or U2100 (N_2100,N_1092,N_1731);
and U2101 (N_2101,N_1453,N_1045);
nand U2102 (N_2102,N_1116,N_1509);
nor U2103 (N_2103,N_1292,N_1169);
and U2104 (N_2104,N_1170,N_1686);
and U2105 (N_2105,N_1023,N_1275);
and U2106 (N_2106,N_1943,N_1544);
and U2107 (N_2107,N_1824,N_1426);
nand U2108 (N_2108,N_1857,N_1928);
nor U2109 (N_2109,N_1120,N_1313);
xor U2110 (N_2110,N_1341,N_1655);
or U2111 (N_2111,N_1673,N_1514);
or U2112 (N_2112,N_1945,N_1582);
xnor U2113 (N_2113,N_1461,N_1968);
xor U2114 (N_2114,N_1442,N_1766);
xnor U2115 (N_2115,N_1922,N_1707);
or U2116 (N_2116,N_1958,N_1633);
nor U2117 (N_2117,N_1223,N_1071);
or U2118 (N_2118,N_1523,N_1758);
or U2119 (N_2119,N_1449,N_1744);
and U2120 (N_2120,N_1665,N_1577);
nand U2121 (N_2121,N_1826,N_1650);
or U2122 (N_2122,N_1153,N_1515);
and U2123 (N_2123,N_1897,N_1542);
nand U2124 (N_2124,N_1560,N_1924);
nand U2125 (N_2125,N_1420,N_1259);
or U2126 (N_2126,N_1812,N_1257);
or U2127 (N_2127,N_1407,N_1531);
xor U2128 (N_2128,N_1951,N_1765);
xor U2129 (N_2129,N_1158,N_1302);
nor U2130 (N_2130,N_1139,N_1735);
nand U2131 (N_2131,N_1591,N_1690);
nor U2132 (N_2132,N_1843,N_1809);
nor U2133 (N_2133,N_1948,N_1728);
xnor U2134 (N_2134,N_1002,N_1433);
or U2135 (N_2135,N_1992,N_1161);
or U2136 (N_2136,N_1877,N_1422);
xnor U2137 (N_2137,N_1322,N_1775);
or U2138 (N_2138,N_1762,N_1082);
and U2139 (N_2139,N_1713,N_1181);
nand U2140 (N_2140,N_1198,N_1740);
xnor U2141 (N_2141,N_1830,N_1026);
or U2142 (N_2142,N_1778,N_1840);
nor U2143 (N_2143,N_1251,N_1358);
xor U2144 (N_2144,N_1553,N_1097);
and U2145 (N_2145,N_1722,N_1803);
and U2146 (N_2146,N_1307,N_1865);
nand U2147 (N_2147,N_1294,N_1136);
xnor U2148 (N_2148,N_1783,N_1781);
nor U2149 (N_2149,N_1651,N_1798);
nand U2150 (N_2150,N_1380,N_1286);
xor U2151 (N_2151,N_1042,N_1459);
xor U2152 (N_2152,N_1193,N_1583);
xor U2153 (N_2153,N_1753,N_1236);
and U2154 (N_2154,N_1489,N_1729);
and U2155 (N_2155,N_1899,N_1098);
xnor U2156 (N_2156,N_1462,N_1452);
and U2157 (N_2157,N_1454,N_1411);
or U2158 (N_2158,N_1937,N_1131);
or U2159 (N_2159,N_1705,N_1403);
and U2160 (N_2160,N_1296,N_1003);
or U2161 (N_2161,N_1821,N_1141);
xor U2162 (N_2162,N_1652,N_1838);
xor U2163 (N_2163,N_1896,N_1886);
nand U2164 (N_2164,N_1328,N_1233);
or U2165 (N_2165,N_1398,N_1242);
xor U2166 (N_2166,N_1371,N_1360);
nand U2167 (N_2167,N_1263,N_1325);
or U2168 (N_2168,N_1868,N_1848);
and U2169 (N_2169,N_1065,N_1628);
or U2170 (N_2170,N_1155,N_1386);
and U2171 (N_2171,N_1845,N_1145);
nor U2172 (N_2172,N_1751,N_1587);
nor U2173 (N_2173,N_1228,N_1195);
nand U2174 (N_2174,N_1213,N_1494);
or U2175 (N_2175,N_1216,N_1290);
or U2176 (N_2176,N_1094,N_1476);
nand U2177 (N_2177,N_1396,N_1640);
and U2178 (N_2178,N_1832,N_1630);
nor U2179 (N_2179,N_1306,N_1874);
or U2180 (N_2180,N_1395,N_1477);
or U2181 (N_2181,N_1889,N_1256);
nand U2182 (N_2182,N_1847,N_1387);
and U2183 (N_2183,N_1935,N_1986);
xnor U2184 (N_2184,N_1164,N_1471);
nor U2185 (N_2185,N_1902,N_1208);
xnor U2186 (N_2186,N_1601,N_1586);
nand U2187 (N_2187,N_1885,N_1895);
or U2188 (N_2188,N_1295,N_1615);
or U2189 (N_2189,N_1769,N_1101);
or U2190 (N_2190,N_1829,N_1481);
or U2191 (N_2191,N_1500,N_1372);
nand U2192 (N_2192,N_1855,N_1872);
nor U2193 (N_2193,N_1600,N_1529);
nor U2194 (N_2194,N_1717,N_1973);
nand U2195 (N_2195,N_1984,N_1304);
or U2196 (N_2196,N_1384,N_1068);
or U2197 (N_2197,N_1954,N_1916);
or U2198 (N_2198,N_1390,N_1551);
nand U2199 (N_2199,N_1921,N_1941);
or U2200 (N_2200,N_1527,N_1332);
or U2201 (N_2201,N_1903,N_1260);
xnor U2202 (N_2202,N_1697,N_1785);
xor U2203 (N_2203,N_1608,N_1008);
nor U2204 (N_2204,N_1750,N_1353);
nor U2205 (N_2205,N_1297,N_1891);
xor U2206 (N_2206,N_1314,N_1270);
nand U2207 (N_2207,N_1566,N_1154);
xor U2208 (N_2208,N_1133,N_1550);
nand U2209 (N_2209,N_1988,N_1691);
xor U2210 (N_2210,N_1876,N_1563);
and U2211 (N_2211,N_1850,N_1870);
and U2212 (N_2212,N_1179,N_1382);
nand U2213 (N_2213,N_1498,N_1757);
nand U2214 (N_2214,N_1265,N_1733);
nand U2215 (N_2215,N_1054,N_1898);
nand U2216 (N_2216,N_1599,N_1122);
nor U2217 (N_2217,N_1346,N_1634);
nor U2218 (N_2218,N_1414,N_1281);
xor U2219 (N_2219,N_1754,N_1927);
and U2220 (N_2220,N_1980,N_1156);
and U2221 (N_2221,N_1726,N_1474);
nor U2222 (N_2222,N_1245,N_1457);
or U2223 (N_2223,N_1510,N_1117);
nor U2224 (N_2224,N_1632,N_1585);
xor U2225 (N_2225,N_1795,N_1349);
nand U2226 (N_2226,N_1535,N_1906);
and U2227 (N_2227,N_1370,N_1706);
nand U2228 (N_2228,N_1207,N_1364);
and U2229 (N_2229,N_1907,N_1226);
and U2230 (N_2230,N_1790,N_1369);
xnor U2231 (N_2231,N_1718,N_1742);
nor U2232 (N_2232,N_1379,N_1725);
nor U2233 (N_2233,N_1890,N_1401);
xor U2234 (N_2234,N_1524,N_1408);
nand U2235 (N_2235,N_1430,N_1801);
nor U2236 (N_2236,N_1506,N_1559);
and U2237 (N_2237,N_1770,N_1828);
or U2238 (N_2238,N_1835,N_1115);
nand U2239 (N_2239,N_1277,N_1177);
nor U2240 (N_2240,N_1543,N_1910);
or U2241 (N_2241,N_1969,N_1879);
or U2242 (N_2242,N_1088,N_1184);
and U2243 (N_2243,N_1694,N_1359);
or U2244 (N_2244,N_1567,N_1367);
nor U2245 (N_2245,N_1621,N_1007);
nand U2246 (N_2246,N_1912,N_1165);
or U2247 (N_2247,N_1252,N_1611);
or U2248 (N_2248,N_1077,N_1268);
nor U2249 (N_2249,N_1773,N_1491);
and U2250 (N_2250,N_1645,N_1990);
nand U2251 (N_2251,N_1043,N_1012);
and U2252 (N_2252,N_1923,N_1649);
and U2253 (N_2253,N_1784,N_1873);
or U2254 (N_2254,N_1799,N_1704);
xor U2255 (N_2255,N_1483,N_1159);
nor U2256 (N_2256,N_1244,N_1333);
nor U2257 (N_2257,N_1863,N_1894);
nor U2258 (N_2258,N_1925,N_1496);
xnor U2259 (N_2259,N_1114,N_1942);
nor U2260 (N_2260,N_1526,N_1887);
or U2261 (N_2261,N_1421,N_1278);
and U2262 (N_2262,N_1930,N_1214);
nor U2263 (N_2263,N_1063,N_1792);
and U2264 (N_2264,N_1202,N_1013);
and U2265 (N_2265,N_1011,N_1084);
or U2266 (N_2266,N_1106,N_1413);
nor U2267 (N_2267,N_1810,N_1878);
nor U2268 (N_2268,N_1825,N_1503);
xor U2269 (N_2269,N_1345,N_1605);
xor U2270 (N_2270,N_1456,N_1032);
xnor U2271 (N_2271,N_1152,N_1593);
and U2272 (N_2272,N_1377,N_1518);
or U2273 (N_2273,N_1964,N_1310);
and U2274 (N_2274,N_1173,N_1804);
nor U2275 (N_2275,N_1205,N_1001);
xnor U2276 (N_2276,N_1748,N_1182);
xnor U2277 (N_2277,N_1624,N_1178);
or U2278 (N_2278,N_1949,N_1900);
and U2279 (N_2279,N_1057,N_1201);
nor U2280 (N_2280,N_1220,N_1864);
and U2281 (N_2281,N_1654,N_1743);
xnor U2282 (N_2282,N_1440,N_1548);
xor U2283 (N_2283,N_1952,N_1091);
nor U2284 (N_2284,N_1805,N_1151);
nor U2285 (N_2285,N_1334,N_1467);
xnor U2286 (N_2286,N_1674,N_1693);
nand U2287 (N_2287,N_1493,N_1163);
or U2288 (N_2288,N_1918,N_1807);
and U2289 (N_2289,N_1246,N_1352);
nand U2290 (N_2290,N_1343,N_1534);
or U2291 (N_2291,N_1678,N_1485);
nor U2292 (N_2292,N_1589,N_1501);
or U2293 (N_2293,N_1185,N_1653);
and U2294 (N_2294,N_1137,N_1981);
xor U2295 (N_2295,N_1125,N_1708);
nand U2296 (N_2296,N_1961,N_1347);
nor U2297 (N_2297,N_1381,N_1794);
or U2298 (N_2298,N_1666,N_1028);
nand U2299 (N_2299,N_1516,N_1034);
xor U2300 (N_2300,N_1856,N_1176);
or U2301 (N_2301,N_1056,N_1933);
xor U2302 (N_2302,N_1869,N_1020);
or U2303 (N_2303,N_1679,N_1776);
nand U2304 (N_2304,N_1017,N_1237);
nand U2305 (N_2305,N_1280,N_1919);
nor U2306 (N_2306,N_1112,N_1363);
and U2307 (N_2307,N_1446,N_1974);
nor U2308 (N_2308,N_1504,N_1121);
and U2309 (N_2309,N_1844,N_1892);
nand U2310 (N_2310,N_1250,N_1211);
or U2311 (N_2311,N_1648,N_1319);
nor U2312 (N_2312,N_1598,N_1087);
xnor U2313 (N_2313,N_1796,N_1473);
nor U2314 (N_2314,N_1617,N_1044);
and U2315 (N_2315,N_1888,N_1118);
xor U2316 (N_2316,N_1734,N_1190);
or U2317 (N_2317,N_1338,N_1797);
nor U2318 (N_2318,N_1859,N_1344);
nor U2319 (N_2319,N_1326,N_1642);
or U2320 (N_2320,N_1238,N_1450);
or U2321 (N_2321,N_1575,N_1685);
and U2322 (N_2322,N_1737,N_1557);
and U2323 (N_2323,N_1639,N_1971);
nor U2324 (N_2324,N_1267,N_1549);
and U2325 (N_2325,N_1348,N_1736);
or U2326 (N_2326,N_1808,N_1212);
or U2327 (N_2327,N_1675,N_1597);
nor U2328 (N_2328,N_1860,N_1823);
and U2329 (N_2329,N_1715,N_1016);
nor U2330 (N_2330,N_1486,N_1901);
and U2331 (N_2331,N_1724,N_1266);
nand U2332 (N_2332,N_1625,N_1174);
and U2333 (N_2333,N_1458,N_1273);
or U2334 (N_2334,N_1932,N_1261);
and U2335 (N_2335,N_1946,N_1108);
nand U2336 (N_2336,N_1532,N_1168);
nand U2337 (N_2337,N_1460,N_1030);
nor U2338 (N_2338,N_1010,N_1989);
or U2339 (N_2339,N_1657,N_1606);
and U2340 (N_2340,N_1721,N_1335);
nor U2341 (N_2341,N_1741,N_1822);
and U2342 (N_2342,N_1005,N_1090);
nand U2343 (N_2343,N_1388,N_1183);
or U2344 (N_2344,N_1562,N_1443);
nand U2345 (N_2345,N_1763,N_1019);
xor U2346 (N_2346,N_1701,N_1229);
nand U2347 (N_2347,N_1438,N_1085);
nand U2348 (N_2348,N_1732,N_1578);
xnor U2349 (N_2349,N_1994,N_1699);
or U2350 (N_2350,N_1464,N_1482);
nand U2351 (N_2351,N_1618,N_1234);
nor U2352 (N_2352,N_1366,N_1802);
xnor U2353 (N_2353,N_1365,N_1738);
or U2354 (N_2354,N_1191,N_1915);
or U2355 (N_2355,N_1979,N_1052);
nand U2356 (N_2356,N_1469,N_1768);
nor U2357 (N_2357,N_1463,N_1282);
or U2358 (N_2358,N_1499,N_1613);
and U2359 (N_2359,N_1816,N_1774);
and U2360 (N_2360,N_1230,N_1074);
nor U2361 (N_2361,N_1646,N_1987);
nor U2362 (N_2362,N_1752,N_1662);
xor U2363 (N_2363,N_1419,N_1977);
nand U2364 (N_2364,N_1062,N_1227);
and U2365 (N_2365,N_1107,N_1135);
and U2366 (N_2366,N_1162,N_1787);
nand U2367 (N_2367,N_1311,N_1998);
xor U2368 (N_2368,N_1123,N_1262);
and U2369 (N_2369,N_1709,N_1997);
nor U2370 (N_2370,N_1470,N_1631);
nor U2371 (N_2371,N_1203,N_1248);
xnor U2372 (N_2372,N_1127,N_1893);
or U2373 (N_2373,N_1186,N_1058);
and U2374 (N_2374,N_1405,N_1455);
xor U2375 (N_2375,N_1409,N_1539);
nor U2376 (N_2376,N_1580,N_1546);
nor U2377 (N_2377,N_1637,N_1537);
xnor U2378 (N_2378,N_1342,N_1965);
or U2379 (N_2379,N_1967,N_1745);
or U2380 (N_2380,N_1565,N_1519);
nor U2381 (N_2381,N_1999,N_1545);
or U2382 (N_2382,N_1920,N_1100);
and U2383 (N_2383,N_1982,N_1031);
xnor U2384 (N_2384,N_1643,N_1909);
nand U2385 (N_2385,N_1222,N_1303);
and U2386 (N_2386,N_1661,N_1429);
and U2387 (N_2387,N_1330,N_1144);
nand U2388 (N_2388,N_1616,N_1076);
and U2389 (N_2389,N_1066,N_1623);
xor U2390 (N_2390,N_1755,N_1451);
or U2391 (N_2391,N_1561,N_1719);
xnor U2392 (N_2392,N_1434,N_1350);
or U2393 (N_2393,N_1243,N_1475);
or U2394 (N_2394,N_1659,N_1720);
xnor U2395 (N_2395,N_1105,N_1354);
xnor U2396 (N_2396,N_1554,N_1445);
nand U2397 (N_2397,N_1484,N_1911);
xnor U2398 (N_2398,N_1495,N_1356);
and U2399 (N_2399,N_1520,N_1406);
or U2400 (N_2400,N_1287,N_1351);
nor U2401 (N_2401,N_1849,N_1428);
nand U2402 (N_2402,N_1777,N_1852);
xnor U2403 (N_2403,N_1048,N_1368);
xnor U2404 (N_2404,N_1298,N_1271);
nand U2405 (N_2405,N_1487,N_1588);
nor U2406 (N_2406,N_1818,N_1604);
or U2407 (N_2407,N_1854,N_1018);
and U2408 (N_2408,N_1046,N_1219);
or U2409 (N_2409,N_1321,N_1791);
nor U2410 (N_2410,N_1331,N_1576);
nand U2411 (N_2411,N_1130,N_1552);
and U2412 (N_2412,N_1050,N_1833);
and U2413 (N_2413,N_1037,N_1547);
and U2414 (N_2414,N_1439,N_1418);
or U2415 (N_2415,N_1692,N_1072);
nand U2416 (N_2416,N_1309,N_1073);
xnor U2417 (N_2417,N_1385,N_1389);
or U2418 (N_2418,N_1006,N_1466);
or U2419 (N_2419,N_1541,N_1664);
xor U2420 (N_2420,N_1950,N_1103);
nand U2421 (N_2421,N_1688,N_1508);
nand U2422 (N_2422,N_1305,N_1638);
nand U2423 (N_2423,N_1839,N_1480);
and U2424 (N_2424,N_1727,N_1241);
nor U2425 (N_2425,N_1517,N_1564);
or U2426 (N_2426,N_1677,N_1235);
nor U2427 (N_2427,N_1658,N_1711);
xor U2428 (N_2428,N_1682,N_1570);
nand U2429 (N_2429,N_1148,N_1595);
nand U2430 (N_2430,N_1035,N_1425);
nand U2431 (N_2431,N_1104,N_1714);
xnor U2432 (N_2432,N_1240,N_1027);
xnor U2433 (N_2433,N_1448,N_1086);
nand U2434 (N_2434,N_1647,N_1444);
xor U2435 (N_2435,N_1024,N_1636);
nand U2436 (N_2436,N_1684,N_1996);
nand U2437 (N_2437,N_1676,N_1036);
nand U2438 (N_2438,N_1592,N_1749);
xor U2439 (N_2439,N_1400,N_1393);
nand U2440 (N_2440,N_1255,N_1505);
nor U2441 (N_2441,N_1739,N_1014);
or U2442 (N_2442,N_1301,N_1039);
and U2443 (N_2443,N_1015,N_1806);
xnor U2444 (N_2444,N_1147,N_1329);
xnor U2445 (N_2445,N_1053,N_1536);
xor U2446 (N_2446,N_1157,N_1111);
nand U2447 (N_2447,N_1315,N_1339);
or U2448 (N_2448,N_1378,N_1602);
xnor U2449 (N_2449,N_1820,N_1793);
nand U2450 (N_2450,N_1285,N_1132);
and U2451 (N_2451,N_1289,N_1150);
nor U2452 (N_2452,N_1171,N_1703);
and U2453 (N_2453,N_1938,N_1700);
and U2454 (N_2454,N_1392,N_1204);
or U2455 (N_2455,N_1881,N_1009);
xnor U2456 (N_2456,N_1814,N_1465);
or U2457 (N_2457,N_1140,N_1067);
xor U2458 (N_2458,N_1522,N_1568);
or U2459 (N_2459,N_1614,N_1021);
and U2460 (N_2460,N_1813,N_1960);
nor U2461 (N_2461,N_1641,N_1533);
and U2462 (N_2462,N_1427,N_1468);
or U2463 (N_2463,N_1687,N_1083);
and U2464 (N_2464,N_1361,N_1209);
nor U2465 (N_2465,N_1394,N_1134);
xor U2466 (N_2466,N_1905,N_1681);
nor U2467 (N_2467,N_1376,N_1022);
nand U2468 (N_2468,N_1415,N_1206);
nor U2469 (N_2469,N_1336,N_1300);
nor U2470 (N_2470,N_1138,N_1269);
and U2471 (N_2471,N_1959,N_1404);
or U2472 (N_2472,N_1196,N_1746);
xor U2473 (N_2473,N_1424,N_1819);
xnor U2474 (N_2474,N_1917,N_1441);
nor U2475 (N_2475,N_1490,N_1124);
nor U2476 (N_2476,N_1247,N_1800);
nand U2477 (N_2477,N_1199,N_1119);
nand U2478 (N_2478,N_1976,N_1488);
nor U2479 (N_2479,N_1258,N_1069);
nor U2480 (N_2480,N_1609,N_1538);
xor U2481 (N_2481,N_1423,N_1284);
xor U2482 (N_2482,N_1081,N_1172);
xor U2483 (N_2483,N_1362,N_1747);
nand U2484 (N_2484,N_1978,N_1584);
xnor U2485 (N_2485,N_1327,N_1574);
nor U2486 (N_2486,N_1492,N_1712);
nand U2487 (N_2487,N_1512,N_1320);
nand U2488 (N_2488,N_1126,N_1883);
and U2489 (N_2489,N_1080,N_1629);
nor U2490 (N_2490,N_1882,N_1620);
nand U2491 (N_2491,N_1936,N_1166);
or U2492 (N_2492,N_1596,N_1089);
or U2493 (N_2493,N_1249,N_1815);
and U2494 (N_2494,N_1175,N_1513);
and U2495 (N_2495,N_1060,N_1995);
and U2496 (N_2496,N_1436,N_1221);
nand U2497 (N_2497,N_1834,N_1095);
and U2498 (N_2498,N_1866,N_1871);
and U2499 (N_2499,N_1610,N_1663);
nand U2500 (N_2500,N_1159,N_1250);
or U2501 (N_2501,N_1626,N_1776);
nand U2502 (N_2502,N_1958,N_1744);
nor U2503 (N_2503,N_1775,N_1151);
nand U2504 (N_2504,N_1706,N_1790);
nor U2505 (N_2505,N_1943,N_1528);
xor U2506 (N_2506,N_1235,N_1124);
nand U2507 (N_2507,N_1332,N_1375);
xor U2508 (N_2508,N_1489,N_1776);
or U2509 (N_2509,N_1338,N_1445);
nor U2510 (N_2510,N_1060,N_1231);
xor U2511 (N_2511,N_1928,N_1141);
and U2512 (N_2512,N_1417,N_1822);
or U2513 (N_2513,N_1447,N_1821);
nor U2514 (N_2514,N_1520,N_1525);
nor U2515 (N_2515,N_1543,N_1291);
nand U2516 (N_2516,N_1348,N_1725);
and U2517 (N_2517,N_1344,N_1982);
or U2518 (N_2518,N_1084,N_1677);
nand U2519 (N_2519,N_1992,N_1861);
nor U2520 (N_2520,N_1457,N_1474);
or U2521 (N_2521,N_1422,N_1509);
nor U2522 (N_2522,N_1272,N_1146);
nor U2523 (N_2523,N_1491,N_1436);
or U2524 (N_2524,N_1103,N_1597);
and U2525 (N_2525,N_1897,N_1178);
nand U2526 (N_2526,N_1833,N_1442);
xnor U2527 (N_2527,N_1482,N_1034);
or U2528 (N_2528,N_1143,N_1354);
or U2529 (N_2529,N_1667,N_1404);
xnor U2530 (N_2530,N_1684,N_1372);
nor U2531 (N_2531,N_1331,N_1579);
or U2532 (N_2532,N_1302,N_1048);
nor U2533 (N_2533,N_1370,N_1122);
or U2534 (N_2534,N_1187,N_1899);
nor U2535 (N_2535,N_1862,N_1733);
and U2536 (N_2536,N_1785,N_1886);
and U2537 (N_2537,N_1078,N_1641);
nand U2538 (N_2538,N_1862,N_1731);
or U2539 (N_2539,N_1120,N_1773);
nor U2540 (N_2540,N_1569,N_1222);
xor U2541 (N_2541,N_1144,N_1825);
xnor U2542 (N_2542,N_1017,N_1209);
nor U2543 (N_2543,N_1265,N_1840);
and U2544 (N_2544,N_1744,N_1072);
or U2545 (N_2545,N_1484,N_1979);
and U2546 (N_2546,N_1883,N_1921);
or U2547 (N_2547,N_1354,N_1026);
nor U2548 (N_2548,N_1282,N_1933);
nand U2549 (N_2549,N_1533,N_1208);
or U2550 (N_2550,N_1985,N_1723);
nand U2551 (N_2551,N_1942,N_1868);
xor U2552 (N_2552,N_1974,N_1061);
and U2553 (N_2553,N_1617,N_1800);
nor U2554 (N_2554,N_1996,N_1102);
nor U2555 (N_2555,N_1772,N_1546);
nand U2556 (N_2556,N_1836,N_1000);
xnor U2557 (N_2557,N_1897,N_1786);
and U2558 (N_2558,N_1288,N_1349);
nand U2559 (N_2559,N_1910,N_1452);
nor U2560 (N_2560,N_1939,N_1015);
and U2561 (N_2561,N_1950,N_1745);
nand U2562 (N_2562,N_1884,N_1655);
or U2563 (N_2563,N_1859,N_1984);
xor U2564 (N_2564,N_1805,N_1917);
or U2565 (N_2565,N_1914,N_1964);
xor U2566 (N_2566,N_1726,N_1334);
and U2567 (N_2567,N_1031,N_1885);
or U2568 (N_2568,N_1386,N_1012);
nor U2569 (N_2569,N_1696,N_1480);
and U2570 (N_2570,N_1520,N_1118);
nand U2571 (N_2571,N_1124,N_1852);
xor U2572 (N_2572,N_1895,N_1932);
xor U2573 (N_2573,N_1695,N_1030);
nor U2574 (N_2574,N_1261,N_1263);
or U2575 (N_2575,N_1582,N_1245);
or U2576 (N_2576,N_1800,N_1036);
nand U2577 (N_2577,N_1648,N_1192);
xor U2578 (N_2578,N_1686,N_1953);
or U2579 (N_2579,N_1297,N_1993);
or U2580 (N_2580,N_1919,N_1028);
xnor U2581 (N_2581,N_1189,N_1179);
nand U2582 (N_2582,N_1232,N_1881);
nand U2583 (N_2583,N_1941,N_1912);
or U2584 (N_2584,N_1769,N_1750);
or U2585 (N_2585,N_1619,N_1403);
or U2586 (N_2586,N_1378,N_1083);
xnor U2587 (N_2587,N_1960,N_1723);
and U2588 (N_2588,N_1633,N_1167);
and U2589 (N_2589,N_1037,N_1281);
nand U2590 (N_2590,N_1391,N_1196);
and U2591 (N_2591,N_1953,N_1577);
and U2592 (N_2592,N_1109,N_1404);
xnor U2593 (N_2593,N_1571,N_1769);
xnor U2594 (N_2594,N_1827,N_1720);
or U2595 (N_2595,N_1606,N_1390);
nor U2596 (N_2596,N_1394,N_1786);
nand U2597 (N_2597,N_1685,N_1368);
xnor U2598 (N_2598,N_1747,N_1347);
or U2599 (N_2599,N_1287,N_1732);
or U2600 (N_2600,N_1881,N_1284);
or U2601 (N_2601,N_1665,N_1757);
xor U2602 (N_2602,N_1303,N_1626);
and U2603 (N_2603,N_1875,N_1658);
and U2604 (N_2604,N_1375,N_1925);
xor U2605 (N_2605,N_1219,N_1171);
nand U2606 (N_2606,N_1190,N_1122);
or U2607 (N_2607,N_1001,N_1047);
nor U2608 (N_2608,N_1757,N_1705);
nand U2609 (N_2609,N_1992,N_1899);
nor U2610 (N_2610,N_1020,N_1028);
xnor U2611 (N_2611,N_1351,N_1068);
and U2612 (N_2612,N_1485,N_1520);
xor U2613 (N_2613,N_1872,N_1818);
or U2614 (N_2614,N_1635,N_1643);
nor U2615 (N_2615,N_1672,N_1897);
or U2616 (N_2616,N_1779,N_1627);
xnor U2617 (N_2617,N_1537,N_1996);
nand U2618 (N_2618,N_1343,N_1768);
nor U2619 (N_2619,N_1451,N_1627);
xnor U2620 (N_2620,N_1232,N_1984);
nor U2621 (N_2621,N_1979,N_1010);
and U2622 (N_2622,N_1387,N_1050);
nor U2623 (N_2623,N_1219,N_1195);
or U2624 (N_2624,N_1178,N_1866);
nor U2625 (N_2625,N_1821,N_1187);
and U2626 (N_2626,N_1482,N_1014);
and U2627 (N_2627,N_1792,N_1472);
xnor U2628 (N_2628,N_1965,N_1570);
xnor U2629 (N_2629,N_1007,N_1913);
and U2630 (N_2630,N_1293,N_1200);
and U2631 (N_2631,N_1373,N_1920);
nor U2632 (N_2632,N_1974,N_1629);
nand U2633 (N_2633,N_1096,N_1407);
and U2634 (N_2634,N_1358,N_1323);
and U2635 (N_2635,N_1739,N_1848);
xor U2636 (N_2636,N_1914,N_1166);
and U2637 (N_2637,N_1024,N_1755);
or U2638 (N_2638,N_1939,N_1135);
xor U2639 (N_2639,N_1765,N_1918);
nand U2640 (N_2640,N_1210,N_1480);
or U2641 (N_2641,N_1348,N_1607);
and U2642 (N_2642,N_1901,N_1491);
nor U2643 (N_2643,N_1686,N_1889);
nor U2644 (N_2644,N_1661,N_1392);
and U2645 (N_2645,N_1817,N_1785);
nor U2646 (N_2646,N_1625,N_1388);
nand U2647 (N_2647,N_1179,N_1434);
xnor U2648 (N_2648,N_1234,N_1625);
or U2649 (N_2649,N_1989,N_1574);
or U2650 (N_2650,N_1569,N_1827);
xnor U2651 (N_2651,N_1642,N_1838);
nand U2652 (N_2652,N_1217,N_1103);
nor U2653 (N_2653,N_1811,N_1214);
nor U2654 (N_2654,N_1600,N_1750);
or U2655 (N_2655,N_1726,N_1316);
nand U2656 (N_2656,N_1985,N_1559);
xor U2657 (N_2657,N_1746,N_1316);
xor U2658 (N_2658,N_1909,N_1094);
and U2659 (N_2659,N_1976,N_1862);
or U2660 (N_2660,N_1137,N_1408);
and U2661 (N_2661,N_1167,N_1638);
nand U2662 (N_2662,N_1238,N_1160);
nor U2663 (N_2663,N_1921,N_1861);
or U2664 (N_2664,N_1172,N_1430);
xor U2665 (N_2665,N_1119,N_1708);
nand U2666 (N_2666,N_1912,N_1296);
or U2667 (N_2667,N_1010,N_1188);
and U2668 (N_2668,N_1660,N_1188);
xor U2669 (N_2669,N_1556,N_1217);
or U2670 (N_2670,N_1974,N_1479);
or U2671 (N_2671,N_1321,N_1853);
nor U2672 (N_2672,N_1866,N_1200);
and U2673 (N_2673,N_1723,N_1682);
nor U2674 (N_2674,N_1217,N_1105);
nor U2675 (N_2675,N_1519,N_1414);
nor U2676 (N_2676,N_1419,N_1103);
nand U2677 (N_2677,N_1416,N_1851);
and U2678 (N_2678,N_1817,N_1669);
nor U2679 (N_2679,N_1228,N_1443);
xor U2680 (N_2680,N_1301,N_1938);
or U2681 (N_2681,N_1391,N_1499);
and U2682 (N_2682,N_1797,N_1150);
xnor U2683 (N_2683,N_1481,N_1401);
nand U2684 (N_2684,N_1334,N_1905);
nor U2685 (N_2685,N_1483,N_1367);
nand U2686 (N_2686,N_1175,N_1523);
xor U2687 (N_2687,N_1674,N_1282);
nand U2688 (N_2688,N_1407,N_1338);
nor U2689 (N_2689,N_1066,N_1750);
nand U2690 (N_2690,N_1869,N_1280);
or U2691 (N_2691,N_1808,N_1683);
and U2692 (N_2692,N_1692,N_1909);
and U2693 (N_2693,N_1540,N_1597);
and U2694 (N_2694,N_1863,N_1672);
and U2695 (N_2695,N_1734,N_1639);
xnor U2696 (N_2696,N_1732,N_1556);
or U2697 (N_2697,N_1284,N_1149);
or U2698 (N_2698,N_1913,N_1944);
or U2699 (N_2699,N_1149,N_1161);
xnor U2700 (N_2700,N_1826,N_1366);
xor U2701 (N_2701,N_1522,N_1860);
xor U2702 (N_2702,N_1241,N_1844);
nand U2703 (N_2703,N_1562,N_1926);
nor U2704 (N_2704,N_1013,N_1085);
xor U2705 (N_2705,N_1419,N_1831);
or U2706 (N_2706,N_1877,N_1224);
xor U2707 (N_2707,N_1916,N_1447);
and U2708 (N_2708,N_1017,N_1348);
nor U2709 (N_2709,N_1037,N_1232);
xnor U2710 (N_2710,N_1893,N_1001);
and U2711 (N_2711,N_1994,N_1993);
xnor U2712 (N_2712,N_1665,N_1688);
xnor U2713 (N_2713,N_1715,N_1284);
or U2714 (N_2714,N_1252,N_1946);
and U2715 (N_2715,N_1096,N_1491);
xnor U2716 (N_2716,N_1135,N_1699);
and U2717 (N_2717,N_1920,N_1988);
and U2718 (N_2718,N_1758,N_1624);
nand U2719 (N_2719,N_1612,N_1939);
or U2720 (N_2720,N_1572,N_1301);
or U2721 (N_2721,N_1377,N_1929);
nor U2722 (N_2722,N_1549,N_1241);
and U2723 (N_2723,N_1999,N_1475);
nand U2724 (N_2724,N_1364,N_1614);
xnor U2725 (N_2725,N_1648,N_1751);
nor U2726 (N_2726,N_1921,N_1963);
nor U2727 (N_2727,N_1521,N_1280);
or U2728 (N_2728,N_1487,N_1311);
nand U2729 (N_2729,N_1499,N_1115);
and U2730 (N_2730,N_1138,N_1618);
nor U2731 (N_2731,N_1136,N_1130);
and U2732 (N_2732,N_1493,N_1633);
xnor U2733 (N_2733,N_1905,N_1910);
nand U2734 (N_2734,N_1408,N_1916);
nand U2735 (N_2735,N_1242,N_1484);
nor U2736 (N_2736,N_1734,N_1345);
or U2737 (N_2737,N_1194,N_1754);
nor U2738 (N_2738,N_1875,N_1825);
xor U2739 (N_2739,N_1509,N_1939);
and U2740 (N_2740,N_1998,N_1980);
and U2741 (N_2741,N_1797,N_1438);
nor U2742 (N_2742,N_1584,N_1742);
nor U2743 (N_2743,N_1023,N_1726);
or U2744 (N_2744,N_1844,N_1113);
nor U2745 (N_2745,N_1517,N_1778);
and U2746 (N_2746,N_1507,N_1255);
nor U2747 (N_2747,N_1311,N_1344);
xnor U2748 (N_2748,N_1273,N_1803);
and U2749 (N_2749,N_1147,N_1613);
or U2750 (N_2750,N_1437,N_1489);
or U2751 (N_2751,N_1481,N_1681);
nand U2752 (N_2752,N_1068,N_1739);
nor U2753 (N_2753,N_1654,N_1913);
and U2754 (N_2754,N_1584,N_1092);
and U2755 (N_2755,N_1723,N_1471);
xnor U2756 (N_2756,N_1166,N_1000);
nor U2757 (N_2757,N_1302,N_1878);
or U2758 (N_2758,N_1435,N_1421);
and U2759 (N_2759,N_1160,N_1656);
xnor U2760 (N_2760,N_1437,N_1393);
and U2761 (N_2761,N_1970,N_1579);
nor U2762 (N_2762,N_1245,N_1496);
nor U2763 (N_2763,N_1410,N_1081);
nor U2764 (N_2764,N_1522,N_1970);
nand U2765 (N_2765,N_1591,N_1073);
nor U2766 (N_2766,N_1023,N_1816);
or U2767 (N_2767,N_1575,N_1814);
and U2768 (N_2768,N_1062,N_1724);
nor U2769 (N_2769,N_1986,N_1756);
nor U2770 (N_2770,N_1203,N_1309);
or U2771 (N_2771,N_1009,N_1283);
nor U2772 (N_2772,N_1656,N_1451);
or U2773 (N_2773,N_1851,N_1356);
nand U2774 (N_2774,N_1685,N_1897);
nand U2775 (N_2775,N_1902,N_1420);
or U2776 (N_2776,N_1013,N_1516);
or U2777 (N_2777,N_1116,N_1966);
nor U2778 (N_2778,N_1382,N_1209);
or U2779 (N_2779,N_1433,N_1787);
nand U2780 (N_2780,N_1539,N_1115);
xnor U2781 (N_2781,N_1831,N_1051);
nand U2782 (N_2782,N_1071,N_1072);
nor U2783 (N_2783,N_1806,N_1214);
xor U2784 (N_2784,N_1870,N_1756);
and U2785 (N_2785,N_1266,N_1707);
nand U2786 (N_2786,N_1184,N_1995);
nor U2787 (N_2787,N_1776,N_1318);
and U2788 (N_2788,N_1376,N_1814);
and U2789 (N_2789,N_1844,N_1154);
or U2790 (N_2790,N_1830,N_1103);
or U2791 (N_2791,N_1104,N_1420);
nor U2792 (N_2792,N_1273,N_1336);
xor U2793 (N_2793,N_1517,N_1491);
nor U2794 (N_2794,N_1200,N_1815);
nand U2795 (N_2795,N_1071,N_1855);
xnor U2796 (N_2796,N_1142,N_1628);
or U2797 (N_2797,N_1208,N_1386);
or U2798 (N_2798,N_1573,N_1207);
or U2799 (N_2799,N_1135,N_1304);
and U2800 (N_2800,N_1151,N_1408);
nor U2801 (N_2801,N_1892,N_1362);
or U2802 (N_2802,N_1051,N_1330);
or U2803 (N_2803,N_1432,N_1620);
or U2804 (N_2804,N_1251,N_1734);
xnor U2805 (N_2805,N_1260,N_1377);
and U2806 (N_2806,N_1989,N_1655);
and U2807 (N_2807,N_1021,N_1869);
and U2808 (N_2808,N_1215,N_1150);
or U2809 (N_2809,N_1552,N_1795);
nor U2810 (N_2810,N_1991,N_1877);
or U2811 (N_2811,N_1438,N_1924);
or U2812 (N_2812,N_1882,N_1166);
nand U2813 (N_2813,N_1327,N_1884);
nor U2814 (N_2814,N_1564,N_1170);
nand U2815 (N_2815,N_1914,N_1247);
and U2816 (N_2816,N_1962,N_1236);
and U2817 (N_2817,N_1202,N_1707);
xor U2818 (N_2818,N_1961,N_1425);
xnor U2819 (N_2819,N_1842,N_1402);
and U2820 (N_2820,N_1548,N_1889);
xnor U2821 (N_2821,N_1680,N_1331);
nand U2822 (N_2822,N_1822,N_1563);
nand U2823 (N_2823,N_1642,N_1235);
nor U2824 (N_2824,N_1422,N_1449);
nand U2825 (N_2825,N_1121,N_1653);
and U2826 (N_2826,N_1716,N_1356);
xor U2827 (N_2827,N_1506,N_1796);
or U2828 (N_2828,N_1166,N_1557);
nor U2829 (N_2829,N_1142,N_1017);
xnor U2830 (N_2830,N_1378,N_1341);
xnor U2831 (N_2831,N_1638,N_1033);
xnor U2832 (N_2832,N_1992,N_1966);
and U2833 (N_2833,N_1167,N_1108);
nand U2834 (N_2834,N_1338,N_1939);
and U2835 (N_2835,N_1739,N_1489);
and U2836 (N_2836,N_1573,N_1056);
or U2837 (N_2837,N_1280,N_1196);
nor U2838 (N_2838,N_1363,N_1509);
xnor U2839 (N_2839,N_1395,N_1538);
and U2840 (N_2840,N_1497,N_1638);
and U2841 (N_2841,N_1368,N_1477);
and U2842 (N_2842,N_1254,N_1763);
xor U2843 (N_2843,N_1040,N_1452);
and U2844 (N_2844,N_1997,N_1714);
nor U2845 (N_2845,N_1614,N_1387);
or U2846 (N_2846,N_1716,N_1064);
nand U2847 (N_2847,N_1932,N_1911);
xor U2848 (N_2848,N_1643,N_1690);
nand U2849 (N_2849,N_1697,N_1726);
nand U2850 (N_2850,N_1562,N_1664);
xor U2851 (N_2851,N_1885,N_1447);
xor U2852 (N_2852,N_1767,N_1091);
nand U2853 (N_2853,N_1194,N_1593);
and U2854 (N_2854,N_1894,N_1536);
and U2855 (N_2855,N_1046,N_1925);
xnor U2856 (N_2856,N_1091,N_1107);
or U2857 (N_2857,N_1269,N_1837);
or U2858 (N_2858,N_1781,N_1402);
or U2859 (N_2859,N_1458,N_1151);
or U2860 (N_2860,N_1140,N_1046);
xor U2861 (N_2861,N_1311,N_1214);
nand U2862 (N_2862,N_1447,N_1923);
nand U2863 (N_2863,N_1894,N_1455);
or U2864 (N_2864,N_1717,N_1242);
xnor U2865 (N_2865,N_1490,N_1174);
xor U2866 (N_2866,N_1421,N_1553);
nor U2867 (N_2867,N_1142,N_1375);
and U2868 (N_2868,N_1834,N_1708);
or U2869 (N_2869,N_1703,N_1045);
and U2870 (N_2870,N_1698,N_1689);
xnor U2871 (N_2871,N_1697,N_1008);
nand U2872 (N_2872,N_1083,N_1184);
xnor U2873 (N_2873,N_1608,N_1882);
xnor U2874 (N_2874,N_1434,N_1207);
or U2875 (N_2875,N_1067,N_1916);
and U2876 (N_2876,N_1401,N_1835);
nand U2877 (N_2877,N_1848,N_1095);
nor U2878 (N_2878,N_1732,N_1491);
or U2879 (N_2879,N_1816,N_1208);
nand U2880 (N_2880,N_1805,N_1028);
or U2881 (N_2881,N_1681,N_1844);
and U2882 (N_2882,N_1610,N_1147);
or U2883 (N_2883,N_1369,N_1992);
or U2884 (N_2884,N_1920,N_1196);
and U2885 (N_2885,N_1516,N_1193);
nor U2886 (N_2886,N_1498,N_1627);
xor U2887 (N_2887,N_1856,N_1592);
xor U2888 (N_2888,N_1753,N_1191);
nor U2889 (N_2889,N_1095,N_1468);
or U2890 (N_2890,N_1466,N_1289);
nand U2891 (N_2891,N_1978,N_1096);
nor U2892 (N_2892,N_1721,N_1259);
and U2893 (N_2893,N_1878,N_1837);
and U2894 (N_2894,N_1082,N_1276);
xnor U2895 (N_2895,N_1678,N_1040);
and U2896 (N_2896,N_1358,N_1595);
or U2897 (N_2897,N_1758,N_1204);
and U2898 (N_2898,N_1723,N_1478);
nor U2899 (N_2899,N_1841,N_1941);
or U2900 (N_2900,N_1284,N_1249);
or U2901 (N_2901,N_1265,N_1547);
or U2902 (N_2902,N_1422,N_1007);
xnor U2903 (N_2903,N_1577,N_1138);
xnor U2904 (N_2904,N_1716,N_1846);
or U2905 (N_2905,N_1053,N_1852);
nand U2906 (N_2906,N_1576,N_1680);
nor U2907 (N_2907,N_1153,N_1002);
nor U2908 (N_2908,N_1682,N_1315);
nor U2909 (N_2909,N_1841,N_1510);
and U2910 (N_2910,N_1951,N_1247);
or U2911 (N_2911,N_1750,N_1163);
nand U2912 (N_2912,N_1703,N_1415);
and U2913 (N_2913,N_1205,N_1865);
nand U2914 (N_2914,N_1391,N_1012);
nand U2915 (N_2915,N_1362,N_1920);
xnor U2916 (N_2916,N_1300,N_1911);
or U2917 (N_2917,N_1838,N_1251);
and U2918 (N_2918,N_1451,N_1146);
or U2919 (N_2919,N_1393,N_1291);
or U2920 (N_2920,N_1790,N_1149);
xor U2921 (N_2921,N_1533,N_1431);
xnor U2922 (N_2922,N_1500,N_1173);
xor U2923 (N_2923,N_1714,N_1200);
nand U2924 (N_2924,N_1650,N_1165);
and U2925 (N_2925,N_1221,N_1336);
nor U2926 (N_2926,N_1211,N_1502);
xor U2927 (N_2927,N_1769,N_1891);
xor U2928 (N_2928,N_1229,N_1580);
xor U2929 (N_2929,N_1066,N_1860);
nor U2930 (N_2930,N_1047,N_1034);
nand U2931 (N_2931,N_1197,N_1151);
nor U2932 (N_2932,N_1762,N_1493);
or U2933 (N_2933,N_1526,N_1188);
or U2934 (N_2934,N_1059,N_1866);
nor U2935 (N_2935,N_1149,N_1741);
and U2936 (N_2936,N_1845,N_1881);
and U2937 (N_2937,N_1536,N_1165);
or U2938 (N_2938,N_1502,N_1443);
or U2939 (N_2939,N_1848,N_1234);
or U2940 (N_2940,N_1456,N_1428);
xnor U2941 (N_2941,N_1910,N_1717);
xor U2942 (N_2942,N_1303,N_1261);
nor U2943 (N_2943,N_1246,N_1005);
nand U2944 (N_2944,N_1159,N_1743);
nor U2945 (N_2945,N_1486,N_1987);
and U2946 (N_2946,N_1653,N_1521);
or U2947 (N_2947,N_1827,N_1437);
and U2948 (N_2948,N_1209,N_1354);
xnor U2949 (N_2949,N_1871,N_1783);
and U2950 (N_2950,N_1499,N_1975);
or U2951 (N_2951,N_1905,N_1106);
nand U2952 (N_2952,N_1594,N_1452);
and U2953 (N_2953,N_1200,N_1835);
nor U2954 (N_2954,N_1893,N_1210);
and U2955 (N_2955,N_1787,N_1699);
or U2956 (N_2956,N_1513,N_1189);
xor U2957 (N_2957,N_1005,N_1798);
xnor U2958 (N_2958,N_1860,N_1244);
and U2959 (N_2959,N_1711,N_1762);
xor U2960 (N_2960,N_1912,N_1958);
nor U2961 (N_2961,N_1627,N_1819);
xor U2962 (N_2962,N_1481,N_1103);
and U2963 (N_2963,N_1838,N_1615);
or U2964 (N_2964,N_1156,N_1994);
nand U2965 (N_2965,N_1618,N_1177);
and U2966 (N_2966,N_1487,N_1246);
or U2967 (N_2967,N_1368,N_1803);
xor U2968 (N_2968,N_1966,N_1913);
nand U2969 (N_2969,N_1091,N_1414);
or U2970 (N_2970,N_1368,N_1968);
and U2971 (N_2971,N_1258,N_1106);
or U2972 (N_2972,N_1977,N_1509);
or U2973 (N_2973,N_1766,N_1845);
nand U2974 (N_2974,N_1651,N_1983);
xor U2975 (N_2975,N_1751,N_1576);
or U2976 (N_2976,N_1452,N_1879);
or U2977 (N_2977,N_1694,N_1811);
xor U2978 (N_2978,N_1239,N_1365);
or U2979 (N_2979,N_1778,N_1217);
or U2980 (N_2980,N_1114,N_1045);
xor U2981 (N_2981,N_1906,N_1097);
xor U2982 (N_2982,N_1512,N_1436);
xor U2983 (N_2983,N_1860,N_1388);
xnor U2984 (N_2984,N_1074,N_1092);
nor U2985 (N_2985,N_1643,N_1590);
or U2986 (N_2986,N_1973,N_1868);
nand U2987 (N_2987,N_1686,N_1073);
nand U2988 (N_2988,N_1779,N_1904);
xor U2989 (N_2989,N_1065,N_1793);
nor U2990 (N_2990,N_1056,N_1805);
xnor U2991 (N_2991,N_1777,N_1715);
nor U2992 (N_2992,N_1539,N_1006);
and U2993 (N_2993,N_1141,N_1756);
or U2994 (N_2994,N_1226,N_1664);
nand U2995 (N_2995,N_1935,N_1614);
nor U2996 (N_2996,N_1066,N_1397);
xnor U2997 (N_2997,N_1267,N_1791);
xor U2998 (N_2998,N_1851,N_1059);
xnor U2999 (N_2999,N_1029,N_1513);
nor U3000 (N_3000,N_2001,N_2046);
nand U3001 (N_3001,N_2210,N_2692);
nand U3002 (N_3002,N_2599,N_2181);
or U3003 (N_3003,N_2035,N_2578);
xor U3004 (N_3004,N_2176,N_2879);
or U3005 (N_3005,N_2389,N_2028);
nand U3006 (N_3006,N_2308,N_2466);
xnor U3007 (N_3007,N_2496,N_2677);
or U3008 (N_3008,N_2188,N_2169);
xnor U3009 (N_3009,N_2849,N_2699);
xnor U3010 (N_3010,N_2768,N_2420);
and U3011 (N_3011,N_2970,N_2938);
xnor U3012 (N_3012,N_2174,N_2593);
or U3013 (N_3013,N_2780,N_2353);
nand U3014 (N_3014,N_2981,N_2041);
nor U3015 (N_3015,N_2914,N_2653);
or U3016 (N_3016,N_2221,N_2450);
nor U3017 (N_3017,N_2425,N_2663);
nand U3018 (N_3018,N_2477,N_2982);
and U3019 (N_3019,N_2608,N_2817);
xor U3020 (N_3020,N_2661,N_2963);
nor U3021 (N_3021,N_2340,N_2871);
and U3022 (N_3022,N_2183,N_2317);
xnor U3023 (N_3023,N_2994,N_2170);
xnor U3024 (N_3024,N_2305,N_2259);
nor U3025 (N_3025,N_2552,N_2918);
or U3026 (N_3026,N_2762,N_2057);
nor U3027 (N_3027,N_2920,N_2048);
nand U3028 (N_3028,N_2104,N_2157);
nand U3029 (N_3029,N_2084,N_2294);
nor U3030 (N_3030,N_2555,N_2063);
or U3031 (N_3031,N_2098,N_2650);
or U3032 (N_3032,N_2953,N_2708);
or U3033 (N_3033,N_2932,N_2944);
nor U3034 (N_3034,N_2710,N_2492);
nand U3035 (N_3035,N_2824,N_2907);
nor U3036 (N_3036,N_2457,N_2255);
nor U3037 (N_3037,N_2628,N_2546);
nor U3038 (N_3038,N_2795,N_2217);
xnor U3039 (N_3039,N_2204,N_2783);
xnor U3040 (N_3040,N_2229,N_2742);
or U3041 (N_3041,N_2293,N_2219);
or U3042 (N_3042,N_2580,N_2805);
nor U3043 (N_3043,N_2822,N_2671);
and U3044 (N_3044,N_2445,N_2139);
and U3045 (N_3045,N_2566,N_2286);
and U3046 (N_3046,N_2825,N_2648);
nor U3047 (N_3047,N_2560,N_2670);
and U3048 (N_3048,N_2263,N_2326);
nor U3049 (N_3049,N_2410,N_2534);
xnor U3050 (N_3050,N_2085,N_2521);
nand U3051 (N_3051,N_2226,N_2960);
nand U3052 (N_3052,N_2527,N_2331);
and U3053 (N_3053,N_2725,N_2744);
nor U3054 (N_3054,N_2830,N_2022);
and U3055 (N_3055,N_2592,N_2922);
nand U3056 (N_3056,N_2644,N_2548);
or U3057 (N_3057,N_2062,N_2270);
nand U3058 (N_3058,N_2213,N_2590);
nor U3059 (N_3059,N_2921,N_2375);
and U3060 (N_3060,N_2327,N_2614);
xnor U3061 (N_3061,N_2987,N_2823);
nand U3062 (N_3062,N_2646,N_2809);
nor U3063 (N_3063,N_2814,N_2924);
and U3064 (N_3064,N_2693,N_2686);
nor U3065 (N_3065,N_2208,N_2471);
and U3066 (N_3066,N_2930,N_2218);
nand U3067 (N_3067,N_2741,N_2258);
nand U3068 (N_3068,N_2969,N_2050);
or U3069 (N_3069,N_2411,N_2165);
xnor U3070 (N_3070,N_2266,N_2113);
nand U3071 (N_3071,N_2443,N_2915);
or U3072 (N_3072,N_2321,N_2382);
xor U3073 (N_3073,N_2985,N_2890);
xnor U3074 (N_3074,N_2612,N_2379);
nor U3075 (N_3075,N_2083,N_2381);
or U3076 (N_3076,N_2297,N_2983);
xor U3077 (N_3077,N_2417,N_2877);
nand U3078 (N_3078,N_2968,N_2225);
or U3079 (N_3079,N_2134,N_2544);
or U3080 (N_3080,N_2554,N_2908);
and U3081 (N_3081,N_2137,N_2750);
xor U3082 (N_3082,N_2336,N_2077);
xnor U3083 (N_3083,N_2127,N_2793);
and U3084 (N_3084,N_2607,N_2964);
xor U3085 (N_3085,N_2860,N_2060);
xnor U3086 (N_3086,N_2843,N_2383);
nand U3087 (N_3087,N_2965,N_2882);
or U3088 (N_3088,N_2299,N_2341);
nand U3089 (N_3089,N_2883,N_2595);
and U3090 (N_3090,N_2110,N_2058);
xor U3091 (N_3091,N_2800,N_2951);
or U3092 (N_3092,N_2702,N_2132);
or U3093 (N_3093,N_2832,N_2281);
xnor U3094 (N_3094,N_2515,N_2867);
and U3095 (N_3095,N_2941,N_2917);
or U3096 (N_3096,N_2704,N_2575);
xnor U3097 (N_3097,N_2666,N_2322);
nor U3098 (N_3098,N_2655,N_2950);
and U3099 (N_3099,N_2080,N_2769);
nand U3100 (N_3100,N_2540,N_2771);
or U3101 (N_3101,N_2014,N_2508);
xnor U3102 (N_3102,N_2449,N_2315);
nand U3103 (N_3103,N_2107,N_2333);
and U3104 (N_3104,N_2444,N_2790);
nor U3105 (N_3105,N_2000,N_2757);
or U3106 (N_3106,N_2818,N_2895);
nor U3107 (N_3107,N_2128,N_2966);
nand U3108 (N_3108,N_2470,N_2288);
nand U3109 (N_3109,N_2977,N_2412);
or U3110 (N_3110,N_2150,N_2533);
nor U3111 (N_3111,N_2786,N_2253);
or U3112 (N_3112,N_2474,N_2522);
nor U3113 (N_3113,N_2268,N_2545);
xnor U3114 (N_3114,N_2448,N_2668);
or U3115 (N_3115,N_2387,N_2638);
nand U3116 (N_3116,N_2397,N_2579);
nand U3117 (N_3117,N_2705,N_2469);
nor U3118 (N_3118,N_2992,N_2166);
nor U3119 (N_3119,N_2532,N_2919);
nand U3120 (N_3120,N_2452,N_2303);
and U3121 (N_3121,N_2282,N_2075);
xnor U3122 (N_3122,N_2766,N_2986);
nand U3123 (N_3123,N_2115,N_2759);
and U3124 (N_3124,N_2130,N_2633);
or U3125 (N_3125,N_2493,N_2119);
nand U3126 (N_3126,N_2989,N_2124);
xor U3127 (N_3127,N_2827,N_2662);
xor U3128 (N_3128,N_2838,N_2484);
xnor U3129 (N_3129,N_2975,N_2740);
nor U3130 (N_3130,N_2594,N_2858);
nand U3131 (N_3131,N_2179,N_2657);
xnor U3132 (N_3132,N_2839,N_2651);
and U3133 (N_3133,N_2993,N_2737);
and U3134 (N_3134,N_2433,N_2197);
xnor U3135 (N_3135,N_2031,N_2459);
or U3136 (N_3136,N_2467,N_2285);
nor U3137 (N_3137,N_2201,N_2419);
nor U3138 (N_3138,N_2461,N_2576);
nor U3139 (N_3139,N_2738,N_2880);
or U3140 (N_3140,N_2630,N_2356);
xor U3141 (N_3141,N_2367,N_2027);
nor U3142 (N_3142,N_2261,N_2088);
or U3143 (N_3143,N_2087,N_2841);
or U3144 (N_3144,N_2319,N_2763);
nor U3145 (N_3145,N_2019,N_2436);
xor U3146 (N_3146,N_2040,N_2585);
nor U3147 (N_3147,N_2034,N_2936);
or U3148 (N_3148,N_2010,N_2761);
nand U3149 (N_3149,N_2765,N_2377);
or U3150 (N_3150,N_2845,N_2894);
or U3151 (N_3151,N_2262,N_2898);
and U3152 (N_3152,N_2149,N_2220);
nor U3153 (N_3153,N_2338,N_2797);
nand U3154 (N_3154,N_2873,N_2352);
and U3155 (N_3155,N_2625,N_2151);
nor U3156 (N_3156,N_2365,N_2931);
xor U3157 (N_3157,N_2602,N_2510);
nand U3158 (N_3158,N_2980,N_2414);
nor U3159 (N_3159,N_2764,N_2067);
and U3160 (N_3160,N_2852,N_2792);
xnor U3161 (N_3161,N_2497,N_2660);
and U3162 (N_3162,N_2649,N_2309);
and U3163 (N_3163,N_2512,N_2007);
and U3164 (N_3164,N_2072,N_2289);
or U3165 (N_3165,N_2287,N_2231);
nor U3166 (N_3166,N_2501,N_2927);
nor U3167 (N_3167,N_2395,N_2161);
or U3168 (N_3168,N_2372,N_2222);
xor U3169 (N_3169,N_2730,N_2847);
nor U3170 (N_3170,N_2051,N_2721);
nor U3171 (N_3171,N_2854,N_2835);
nand U3172 (N_3172,N_2572,N_2009);
nand U3173 (N_3173,N_2587,N_2935);
or U3174 (N_3174,N_2910,N_2784);
xor U3175 (N_3175,N_2094,N_2519);
and U3176 (N_3176,N_2881,N_2836);
nand U3177 (N_3177,N_2652,N_2252);
xnor U3178 (N_3178,N_2206,N_2246);
xor U3179 (N_3179,N_2952,N_2772);
nor U3180 (N_3180,N_2047,N_2480);
nor U3181 (N_3181,N_2974,N_2717);
nand U3182 (N_3182,N_2198,N_2335);
and U3183 (N_3183,N_2549,N_2312);
xor U3184 (N_3184,N_2889,N_2984);
or U3185 (N_3185,N_2209,N_2520);
nor U3186 (N_3186,N_2487,N_2604);
or U3187 (N_3187,N_2866,N_2695);
nor U3188 (N_3188,N_2581,N_2189);
nor U3189 (N_3189,N_2106,N_2362);
or U3190 (N_3190,N_2112,N_2366);
nor U3191 (N_3191,N_2393,N_2925);
xnor U3192 (N_3192,N_2518,N_2082);
and U3193 (N_3193,N_2373,N_2829);
and U3194 (N_3194,N_2929,N_2846);
nor U3195 (N_3195,N_2946,N_2709);
or U3196 (N_3196,N_2167,N_2776);
nand U3197 (N_3197,N_2690,N_2096);
nand U3198 (N_3198,N_2430,N_2878);
nor U3199 (N_3199,N_2066,N_2943);
and U3200 (N_3200,N_2314,N_2525);
xnor U3201 (N_3201,N_2437,N_2739);
and U3202 (N_3202,N_2307,N_2090);
nor U3203 (N_3203,N_2909,N_2736);
and U3204 (N_3204,N_2862,N_2408);
xnor U3205 (N_3205,N_2103,N_2079);
nor U3206 (N_3206,N_2945,N_2828);
nand U3207 (N_3207,N_2834,N_2207);
nor U3208 (N_3208,N_2277,N_2758);
nand U3209 (N_3209,N_2683,N_2215);
nand U3210 (N_3210,N_2928,N_2248);
xor U3211 (N_3211,N_2647,N_2320);
and U3212 (N_3212,N_2329,N_2528);
and U3213 (N_3213,N_2271,N_2260);
nor U3214 (N_3214,N_2146,N_2626);
nand U3215 (N_3215,N_2004,N_2689);
xnor U3216 (N_3216,N_2117,N_2872);
and U3217 (N_3217,N_2426,N_2147);
nor U3218 (N_3218,N_2654,N_2745);
and U3219 (N_3219,N_2685,N_2820);
nand U3220 (N_3220,N_2888,N_2775);
nor U3221 (N_3221,N_2129,N_2301);
and U3222 (N_3222,N_2482,N_2158);
and U3223 (N_3223,N_2177,N_2245);
nand U3224 (N_3224,N_2465,N_2506);
or U3225 (N_3225,N_2617,N_2244);
nand U3226 (N_3226,N_2727,N_2354);
nand U3227 (N_3227,N_2012,N_2276);
or U3228 (N_3228,N_2937,N_2423);
xor U3229 (N_3229,N_2588,N_2233);
or U3230 (N_3230,N_2171,N_2008);
xnor U3231 (N_3231,N_2956,N_2205);
nor U3232 (N_3232,N_2211,N_2391);
xor U3233 (N_3233,N_2324,N_2184);
nor U3234 (N_3234,N_2716,N_2250);
xor U3235 (N_3235,N_2489,N_2400);
nand U3236 (N_3236,N_2837,N_2995);
and U3237 (N_3237,N_2388,N_2154);
xor U3238 (N_3238,N_2316,N_2441);
nor U3239 (N_3239,N_2615,N_2200);
nand U3240 (N_3240,N_2120,N_2409);
nor U3241 (N_3241,N_2337,N_2696);
and U3242 (N_3242,N_2280,N_2893);
and U3243 (N_3243,N_2194,N_2796);
or U3244 (N_3244,N_2573,N_2099);
or U3245 (N_3245,N_2723,N_2609);
xor U3246 (N_3246,N_2947,N_2160);
nor U3247 (N_3247,N_2756,N_2586);
or U3248 (N_3248,N_2070,N_2691);
and U3249 (N_3249,N_2567,N_2483);
or U3250 (N_3250,N_2767,N_2733);
and U3251 (N_3251,N_2688,N_2998);
xor U3252 (N_3252,N_2749,N_2939);
or U3253 (N_3253,N_2111,N_2714);
and U3254 (N_3254,N_2464,N_2643);
nor U3255 (N_3255,N_2190,N_2230);
nand U3256 (N_3256,N_2698,N_2196);
nand U3257 (N_3257,N_2539,N_2017);
nor U3258 (N_3258,N_2529,N_2906);
nor U3259 (N_3259,N_2892,N_2788);
and U3260 (N_3260,N_2264,N_2473);
nand U3261 (N_3261,N_2224,N_2274);
xor U3262 (N_3262,N_2346,N_2620);
nor U3263 (N_3263,N_2360,N_2886);
xnor U3264 (N_3264,N_2494,N_2163);
xor U3265 (N_3265,N_2538,N_2435);
or U3266 (N_3266,N_2491,N_2249);
nor U3267 (N_3267,N_2876,N_2524);
xor U3268 (N_3268,N_2658,N_2957);
nor U3269 (N_3269,N_2095,N_2642);
and U3270 (N_3270,N_2348,N_2514);
nor U3271 (N_3271,N_2342,N_2803);
or U3272 (N_3272,N_2634,N_2141);
and U3273 (N_3273,N_2347,N_2875);
or U3274 (N_3274,N_2054,N_2600);
or U3275 (N_3275,N_2632,N_2156);
xor U3276 (N_3276,N_2061,N_2254);
nor U3277 (N_3277,N_2751,N_2855);
or U3278 (N_3278,N_2967,N_2005);
nand U3279 (N_3279,N_2896,N_2454);
nand U3280 (N_3280,N_2603,N_2451);
and U3281 (N_3281,N_2973,N_2256);
xor U3282 (N_3282,N_2640,N_2731);
and U3283 (N_3283,N_2453,N_2396);
nand U3284 (N_3284,N_2142,N_2678);
and U3285 (N_3285,N_2782,N_2296);
xor U3286 (N_3286,N_2155,N_2350);
or U3287 (N_3287,N_2378,N_2446);
nand U3288 (N_3288,N_2840,N_2002);
xnor U3289 (N_3289,N_2804,N_2926);
nor U3290 (N_3290,N_2416,N_2583);
nand U3291 (N_3291,N_2853,N_2053);
nand U3292 (N_3292,N_2065,N_2162);
and U3293 (N_3293,N_2232,N_2463);
nand U3294 (N_3294,N_2026,N_2861);
or U3295 (N_3295,N_2178,N_2523);
nor U3296 (N_3296,N_2675,N_2310);
and U3297 (N_3297,N_2770,N_2193);
xnor U3298 (N_3298,N_2175,N_2236);
and U3299 (N_3299,N_2240,N_2385);
or U3300 (N_3300,N_2558,N_2623);
and U3301 (N_3301,N_2455,N_2344);
xor U3302 (N_3302,N_2798,N_2015);
nand U3303 (N_3303,N_2298,N_2682);
nor U3304 (N_3304,N_2049,N_2475);
or U3305 (N_3305,N_2187,N_2754);
xor U3306 (N_3306,N_2891,N_2006);
nor U3307 (N_3307,N_2021,N_2025);
xnor U3308 (N_3308,N_2864,N_2799);
nor U3309 (N_3309,N_2507,N_2536);
nand U3310 (N_3310,N_2773,N_2976);
and U3311 (N_3311,N_2753,N_2811);
and U3312 (N_3312,N_2306,N_2887);
nor U3313 (N_3313,N_2369,N_2961);
nor U3314 (N_3314,N_2789,N_2042);
nor U3315 (N_3315,N_2399,N_2684);
or U3316 (N_3316,N_2227,N_2334);
nor U3317 (N_3317,N_2904,N_2752);
or U3318 (N_3318,N_2064,N_2173);
nand U3319 (N_3319,N_2114,N_2153);
and U3320 (N_3320,N_2509,N_2398);
or U3321 (N_3321,N_2092,N_2641);
or U3322 (N_3322,N_2239,N_2903);
and U3323 (N_3323,N_2223,N_2343);
nand U3324 (N_3324,N_2313,N_2624);
nand U3325 (N_3325,N_2561,N_2850);
and U3326 (N_3326,N_2267,N_2667);
xnor U3327 (N_3327,N_2311,N_2029);
nand U3328 (N_3328,N_2582,N_2884);
or U3329 (N_3329,N_2370,N_2923);
or U3330 (N_3330,N_2030,N_2808);
nand U3331 (N_3331,N_2868,N_2897);
or U3332 (N_3332,N_2553,N_2332);
xor U3333 (N_3333,N_2713,N_2318);
nor U3334 (N_3334,N_2720,N_2499);
and U3335 (N_3335,N_2551,N_2136);
nor U3336 (N_3336,N_2364,N_2038);
nor U3337 (N_3337,N_2300,N_2043);
nor U3338 (N_3338,N_2556,N_2037);
xor U3339 (N_3339,N_2363,N_2456);
nand U3340 (N_3340,N_2785,N_2133);
nand U3341 (N_3341,N_2606,N_2724);
nand U3342 (N_3342,N_2024,N_2152);
nor U3343 (N_3343,N_2384,N_2371);
and U3344 (N_3344,N_2091,N_2349);
or U3345 (N_3345,N_2089,N_2290);
nand U3346 (N_3346,N_2781,N_2505);
nand U3347 (N_3347,N_2056,N_2774);
or U3348 (N_3348,N_2086,N_2991);
nor U3349 (N_3349,N_2562,N_2629);
nand U3350 (N_3350,N_2202,N_2905);
xor U3351 (N_3351,N_2068,N_2700);
xnor U3352 (N_3352,N_2901,N_2948);
nand U3353 (N_3353,N_2637,N_2237);
and U3354 (N_3354,N_2674,N_2097);
nor U3355 (N_3355,N_2328,N_2707);
nor U3356 (N_3356,N_2591,N_2971);
nand U3357 (N_3357,N_2447,N_2302);
nand U3358 (N_3358,N_2422,N_2357);
or U3359 (N_3359,N_2760,N_2857);
xor U3360 (N_3360,N_2032,N_2192);
nand U3361 (N_3361,N_2777,N_2413);
or U3362 (N_3362,N_2726,N_2279);
and U3363 (N_3363,N_2269,N_2794);
or U3364 (N_3364,N_2870,N_2656);
nor U3365 (N_3365,N_2504,N_2531);
or U3366 (N_3366,N_2990,N_2123);
nand U3367 (N_3367,N_2530,N_2039);
or U3368 (N_3368,N_2404,N_2517);
nand U3369 (N_3369,N_2673,N_2071);
and U3370 (N_3370,N_2622,N_2011);
or U3371 (N_3371,N_2735,N_2078);
xnor U3372 (N_3372,N_2568,N_2743);
or U3373 (N_3373,N_2486,N_2359);
nor U3374 (N_3374,N_2093,N_2182);
xor U3375 (N_3375,N_2495,N_2500);
xor U3376 (N_3376,N_2711,N_2074);
nor U3377 (N_3377,N_2164,N_2869);
or U3378 (N_3378,N_2863,N_2597);
and U3379 (N_3379,N_2569,N_2787);
nor U3380 (N_3380,N_2427,N_2610);
and U3381 (N_3381,N_2619,N_2899);
xor U3382 (N_3382,N_2358,N_2681);
and U3383 (N_3383,N_2541,N_2016);
nor U3384 (N_3384,N_2535,N_2601);
or U3385 (N_3385,N_2664,N_2415);
nand U3386 (N_3386,N_2791,N_2747);
nand U3387 (N_3387,N_2076,N_2406);
nor U3388 (N_3388,N_2498,N_2885);
nand U3389 (N_3389,N_2748,N_2680);
and U3390 (N_3390,N_2513,N_2728);
and U3391 (N_3391,N_2468,N_2330);
xor U3392 (N_3392,N_2186,N_2842);
xnor U3393 (N_3393,N_2584,N_2865);
and U3394 (N_3394,N_2421,N_2131);
or U3395 (N_3395,N_2003,N_2418);
xor U3396 (N_3396,N_2844,N_2669);
nor U3397 (N_3397,N_2605,N_2687);
xnor U3398 (N_3398,N_2826,N_2503);
nor U3399 (N_3399,N_2479,N_2325);
nand U3400 (N_3400,N_2676,N_2118);
or U3401 (N_3401,N_2949,N_2547);
nor U3402 (N_3402,N_2424,N_2801);
and U3403 (N_3403,N_2511,N_2933);
nand U3404 (N_3404,N_2778,N_2168);
or U3405 (N_3405,N_2972,N_2023);
and U3406 (N_3406,N_2143,N_2434);
and U3407 (N_3407,N_2185,N_2018);
and U3408 (N_3408,N_2485,N_2526);
and U3409 (N_3409,N_2069,N_2942);
xor U3410 (N_3410,N_2402,N_2251);
xor U3411 (N_3411,N_2833,N_2645);
or U3412 (N_3412,N_2394,N_2257);
nand U3413 (N_3413,N_2214,N_2543);
nand U3414 (N_3414,N_2428,N_2323);
xnor U3415 (N_3415,N_2100,N_2490);
nor U3416 (N_3416,N_2911,N_2283);
and U3417 (N_3417,N_2458,N_2559);
or U3418 (N_3418,N_2272,N_2679);
nand U3419 (N_3419,N_2407,N_2988);
and U3420 (N_3420,N_2962,N_2565);
nand U3421 (N_3421,N_2589,N_2275);
nor U3422 (N_3422,N_2339,N_2665);
and U3423 (N_3423,N_2631,N_2036);
and U3424 (N_3424,N_2802,N_2958);
and U3425 (N_3425,N_2719,N_2241);
and U3426 (N_3426,N_2916,N_2235);
nand U3427 (N_3427,N_2295,N_2627);
and U3428 (N_3428,N_2148,N_2557);
and U3429 (N_3429,N_2819,N_2304);
xor U3430 (N_3430,N_2460,N_2374);
and U3431 (N_3431,N_2571,N_2439);
xor U3432 (N_3432,N_2816,N_2125);
nor U3433 (N_3433,N_2831,N_2734);
xor U3434 (N_3434,N_2564,N_2821);
nand U3435 (N_3435,N_2807,N_2101);
and U3436 (N_3436,N_2020,N_2712);
and U3437 (N_3437,N_2563,N_2345);
nor U3438 (N_3438,N_2126,N_2108);
and U3439 (N_3439,N_2755,N_2902);
nor U3440 (N_3440,N_2746,N_2913);
xor U3441 (N_3441,N_2292,N_2247);
and U3442 (N_3442,N_2234,N_2476);
xnor U3443 (N_3443,N_2542,N_2228);
and U3444 (N_3444,N_2488,N_2613);
xor U3445 (N_3445,N_2122,N_2191);
xor U3446 (N_3446,N_2172,N_2856);
or U3447 (N_3447,N_2145,N_2238);
nand U3448 (N_3448,N_2195,N_2574);
nor U3449 (N_3449,N_2999,N_2537);
and U3450 (N_3450,N_2621,N_2138);
and U3451 (N_3451,N_2355,N_2577);
and U3452 (N_3452,N_2874,N_2934);
xor U3453 (N_3453,N_2438,N_2073);
and U3454 (N_3454,N_2978,N_2596);
nor U3455 (N_3455,N_2848,N_2815);
nor U3456 (N_3456,N_2081,N_2718);
or U3457 (N_3457,N_2109,N_2159);
nand U3458 (N_3458,N_2812,N_2284);
and U3459 (N_3459,N_2703,N_2806);
nor U3460 (N_3460,N_2203,N_2442);
xor U3461 (N_3461,N_2706,N_2900);
xor U3462 (N_3462,N_2013,N_2694);
and U3463 (N_3463,N_2401,N_2550);
xor U3464 (N_3464,N_2940,N_2729);
nand U3465 (N_3465,N_2472,N_2055);
or U3466 (N_3466,N_2598,N_2212);
or U3467 (N_3467,N_2105,N_2715);
or U3468 (N_3468,N_2361,N_2672);
and U3469 (N_3469,N_2959,N_2265);
and U3470 (N_3470,N_2502,N_2116);
xnor U3471 (N_3471,N_2462,N_2376);
or U3472 (N_3472,N_2997,N_2697);
and U3473 (N_3473,N_2351,N_2440);
xor U3474 (N_3474,N_2052,N_2996);
and U3475 (N_3475,N_2635,N_2639);
xnor U3476 (N_3476,N_2851,N_2368);
or U3477 (N_3477,N_2722,N_2701);
nor U3478 (N_3478,N_2429,N_2403);
xor U3479 (N_3479,N_2033,N_2779);
nor U3480 (N_3480,N_2431,N_2481);
nor U3481 (N_3481,N_2659,N_2616);
or U3482 (N_3482,N_2618,N_2121);
xnor U3483 (N_3483,N_2392,N_2242);
xnor U3484 (N_3484,N_2570,N_2979);
nor U3485 (N_3485,N_2291,N_2045);
or U3486 (N_3486,N_2243,N_2180);
or U3487 (N_3487,N_2432,N_2810);
and U3488 (N_3488,N_2636,N_2044);
xnor U3489 (N_3489,N_2380,N_2611);
nand U3490 (N_3490,N_2059,N_2273);
xor U3491 (N_3491,N_2199,N_2278);
xor U3492 (N_3492,N_2102,N_2405);
and U3493 (N_3493,N_2859,N_2386);
or U3494 (N_3494,N_2516,N_2140);
nand U3495 (N_3495,N_2135,N_2912);
xnor U3496 (N_3496,N_2216,N_2954);
or U3497 (N_3497,N_2144,N_2955);
nor U3498 (N_3498,N_2813,N_2390);
and U3499 (N_3499,N_2478,N_2732);
nor U3500 (N_3500,N_2166,N_2818);
xor U3501 (N_3501,N_2859,N_2256);
and U3502 (N_3502,N_2761,N_2088);
and U3503 (N_3503,N_2055,N_2846);
xor U3504 (N_3504,N_2765,N_2323);
nor U3505 (N_3505,N_2475,N_2135);
xor U3506 (N_3506,N_2979,N_2770);
nor U3507 (N_3507,N_2038,N_2219);
xnor U3508 (N_3508,N_2166,N_2699);
nor U3509 (N_3509,N_2666,N_2986);
or U3510 (N_3510,N_2012,N_2634);
nand U3511 (N_3511,N_2818,N_2927);
or U3512 (N_3512,N_2385,N_2162);
nor U3513 (N_3513,N_2727,N_2654);
nand U3514 (N_3514,N_2217,N_2394);
xnor U3515 (N_3515,N_2958,N_2559);
xor U3516 (N_3516,N_2740,N_2188);
nand U3517 (N_3517,N_2512,N_2961);
or U3518 (N_3518,N_2212,N_2609);
xnor U3519 (N_3519,N_2993,N_2006);
or U3520 (N_3520,N_2429,N_2163);
and U3521 (N_3521,N_2361,N_2408);
or U3522 (N_3522,N_2810,N_2576);
or U3523 (N_3523,N_2399,N_2529);
xnor U3524 (N_3524,N_2462,N_2006);
xnor U3525 (N_3525,N_2977,N_2379);
xnor U3526 (N_3526,N_2954,N_2101);
xnor U3527 (N_3527,N_2170,N_2454);
and U3528 (N_3528,N_2199,N_2122);
nor U3529 (N_3529,N_2365,N_2664);
nand U3530 (N_3530,N_2664,N_2761);
nand U3531 (N_3531,N_2554,N_2536);
xnor U3532 (N_3532,N_2622,N_2236);
nor U3533 (N_3533,N_2837,N_2339);
nor U3534 (N_3534,N_2264,N_2054);
nand U3535 (N_3535,N_2694,N_2884);
or U3536 (N_3536,N_2133,N_2306);
nand U3537 (N_3537,N_2835,N_2499);
nor U3538 (N_3538,N_2040,N_2793);
nand U3539 (N_3539,N_2997,N_2961);
nand U3540 (N_3540,N_2348,N_2536);
nand U3541 (N_3541,N_2763,N_2185);
nor U3542 (N_3542,N_2738,N_2597);
xor U3543 (N_3543,N_2362,N_2350);
nor U3544 (N_3544,N_2838,N_2483);
and U3545 (N_3545,N_2340,N_2164);
or U3546 (N_3546,N_2142,N_2704);
and U3547 (N_3547,N_2852,N_2687);
or U3548 (N_3548,N_2187,N_2538);
nor U3549 (N_3549,N_2723,N_2155);
and U3550 (N_3550,N_2965,N_2673);
nor U3551 (N_3551,N_2820,N_2842);
xnor U3552 (N_3552,N_2829,N_2620);
xnor U3553 (N_3553,N_2983,N_2526);
nor U3554 (N_3554,N_2690,N_2014);
xnor U3555 (N_3555,N_2268,N_2856);
and U3556 (N_3556,N_2602,N_2986);
xor U3557 (N_3557,N_2289,N_2759);
and U3558 (N_3558,N_2020,N_2480);
nand U3559 (N_3559,N_2612,N_2993);
nor U3560 (N_3560,N_2070,N_2968);
or U3561 (N_3561,N_2194,N_2449);
nor U3562 (N_3562,N_2915,N_2521);
nand U3563 (N_3563,N_2343,N_2435);
xnor U3564 (N_3564,N_2876,N_2303);
xor U3565 (N_3565,N_2112,N_2287);
nand U3566 (N_3566,N_2983,N_2628);
xor U3567 (N_3567,N_2151,N_2227);
and U3568 (N_3568,N_2543,N_2314);
and U3569 (N_3569,N_2205,N_2570);
nor U3570 (N_3570,N_2366,N_2704);
xor U3571 (N_3571,N_2849,N_2484);
xnor U3572 (N_3572,N_2018,N_2254);
nand U3573 (N_3573,N_2596,N_2007);
or U3574 (N_3574,N_2177,N_2558);
xor U3575 (N_3575,N_2538,N_2716);
or U3576 (N_3576,N_2991,N_2137);
or U3577 (N_3577,N_2198,N_2800);
xor U3578 (N_3578,N_2916,N_2509);
nor U3579 (N_3579,N_2875,N_2781);
nand U3580 (N_3580,N_2350,N_2308);
or U3581 (N_3581,N_2027,N_2256);
nand U3582 (N_3582,N_2516,N_2661);
nand U3583 (N_3583,N_2894,N_2723);
nand U3584 (N_3584,N_2152,N_2434);
xor U3585 (N_3585,N_2084,N_2903);
xnor U3586 (N_3586,N_2404,N_2293);
xor U3587 (N_3587,N_2836,N_2724);
and U3588 (N_3588,N_2411,N_2232);
xor U3589 (N_3589,N_2145,N_2424);
xor U3590 (N_3590,N_2249,N_2910);
nor U3591 (N_3591,N_2023,N_2923);
or U3592 (N_3592,N_2140,N_2688);
nand U3593 (N_3593,N_2303,N_2788);
xnor U3594 (N_3594,N_2936,N_2831);
nand U3595 (N_3595,N_2434,N_2359);
xor U3596 (N_3596,N_2727,N_2496);
nand U3597 (N_3597,N_2741,N_2324);
nor U3598 (N_3598,N_2624,N_2857);
xnor U3599 (N_3599,N_2969,N_2838);
or U3600 (N_3600,N_2282,N_2473);
nand U3601 (N_3601,N_2915,N_2480);
and U3602 (N_3602,N_2984,N_2210);
nor U3603 (N_3603,N_2043,N_2261);
xor U3604 (N_3604,N_2543,N_2653);
nor U3605 (N_3605,N_2508,N_2240);
nor U3606 (N_3606,N_2650,N_2948);
nand U3607 (N_3607,N_2119,N_2736);
nand U3608 (N_3608,N_2554,N_2329);
nand U3609 (N_3609,N_2485,N_2906);
or U3610 (N_3610,N_2887,N_2814);
nand U3611 (N_3611,N_2670,N_2574);
nand U3612 (N_3612,N_2553,N_2968);
xor U3613 (N_3613,N_2213,N_2546);
and U3614 (N_3614,N_2425,N_2570);
nor U3615 (N_3615,N_2523,N_2398);
xnor U3616 (N_3616,N_2558,N_2787);
nor U3617 (N_3617,N_2321,N_2595);
and U3618 (N_3618,N_2765,N_2476);
or U3619 (N_3619,N_2214,N_2088);
and U3620 (N_3620,N_2632,N_2570);
nor U3621 (N_3621,N_2800,N_2564);
or U3622 (N_3622,N_2725,N_2111);
or U3623 (N_3623,N_2516,N_2137);
nor U3624 (N_3624,N_2193,N_2050);
nand U3625 (N_3625,N_2472,N_2912);
nor U3626 (N_3626,N_2305,N_2522);
nand U3627 (N_3627,N_2633,N_2605);
xor U3628 (N_3628,N_2644,N_2820);
or U3629 (N_3629,N_2177,N_2333);
and U3630 (N_3630,N_2319,N_2393);
nand U3631 (N_3631,N_2687,N_2974);
xor U3632 (N_3632,N_2053,N_2425);
nor U3633 (N_3633,N_2862,N_2658);
nand U3634 (N_3634,N_2264,N_2785);
or U3635 (N_3635,N_2951,N_2860);
nand U3636 (N_3636,N_2981,N_2075);
xor U3637 (N_3637,N_2914,N_2952);
or U3638 (N_3638,N_2541,N_2869);
nand U3639 (N_3639,N_2058,N_2696);
and U3640 (N_3640,N_2686,N_2066);
xnor U3641 (N_3641,N_2146,N_2694);
nand U3642 (N_3642,N_2453,N_2001);
nor U3643 (N_3643,N_2200,N_2326);
nor U3644 (N_3644,N_2091,N_2036);
nor U3645 (N_3645,N_2518,N_2276);
and U3646 (N_3646,N_2449,N_2595);
xor U3647 (N_3647,N_2308,N_2106);
or U3648 (N_3648,N_2789,N_2738);
or U3649 (N_3649,N_2941,N_2151);
nand U3650 (N_3650,N_2027,N_2446);
or U3651 (N_3651,N_2503,N_2377);
and U3652 (N_3652,N_2882,N_2788);
nand U3653 (N_3653,N_2639,N_2774);
or U3654 (N_3654,N_2497,N_2068);
xnor U3655 (N_3655,N_2091,N_2998);
nand U3656 (N_3656,N_2863,N_2518);
xor U3657 (N_3657,N_2483,N_2264);
or U3658 (N_3658,N_2419,N_2933);
xor U3659 (N_3659,N_2070,N_2538);
nand U3660 (N_3660,N_2121,N_2263);
nor U3661 (N_3661,N_2502,N_2431);
and U3662 (N_3662,N_2371,N_2850);
or U3663 (N_3663,N_2204,N_2877);
nand U3664 (N_3664,N_2964,N_2301);
xnor U3665 (N_3665,N_2906,N_2554);
nor U3666 (N_3666,N_2164,N_2023);
and U3667 (N_3667,N_2840,N_2837);
nand U3668 (N_3668,N_2313,N_2097);
nand U3669 (N_3669,N_2915,N_2970);
or U3670 (N_3670,N_2421,N_2879);
xnor U3671 (N_3671,N_2508,N_2641);
nor U3672 (N_3672,N_2788,N_2183);
nor U3673 (N_3673,N_2063,N_2243);
or U3674 (N_3674,N_2137,N_2876);
nor U3675 (N_3675,N_2709,N_2356);
or U3676 (N_3676,N_2323,N_2930);
or U3677 (N_3677,N_2731,N_2120);
nand U3678 (N_3678,N_2387,N_2447);
or U3679 (N_3679,N_2198,N_2419);
nand U3680 (N_3680,N_2332,N_2202);
xnor U3681 (N_3681,N_2426,N_2556);
and U3682 (N_3682,N_2079,N_2780);
xnor U3683 (N_3683,N_2504,N_2862);
or U3684 (N_3684,N_2581,N_2081);
nand U3685 (N_3685,N_2835,N_2890);
nor U3686 (N_3686,N_2736,N_2403);
nor U3687 (N_3687,N_2761,N_2670);
or U3688 (N_3688,N_2047,N_2720);
xnor U3689 (N_3689,N_2250,N_2656);
and U3690 (N_3690,N_2364,N_2451);
and U3691 (N_3691,N_2544,N_2205);
nor U3692 (N_3692,N_2759,N_2528);
and U3693 (N_3693,N_2936,N_2105);
nor U3694 (N_3694,N_2844,N_2451);
nor U3695 (N_3695,N_2503,N_2346);
and U3696 (N_3696,N_2410,N_2653);
and U3697 (N_3697,N_2651,N_2060);
xor U3698 (N_3698,N_2381,N_2327);
or U3699 (N_3699,N_2623,N_2502);
xor U3700 (N_3700,N_2034,N_2489);
nor U3701 (N_3701,N_2065,N_2401);
or U3702 (N_3702,N_2603,N_2443);
and U3703 (N_3703,N_2464,N_2298);
or U3704 (N_3704,N_2437,N_2259);
nand U3705 (N_3705,N_2391,N_2681);
or U3706 (N_3706,N_2415,N_2243);
nand U3707 (N_3707,N_2132,N_2568);
nand U3708 (N_3708,N_2662,N_2297);
or U3709 (N_3709,N_2244,N_2292);
xnor U3710 (N_3710,N_2686,N_2506);
nor U3711 (N_3711,N_2893,N_2202);
xor U3712 (N_3712,N_2872,N_2073);
nor U3713 (N_3713,N_2813,N_2427);
or U3714 (N_3714,N_2838,N_2543);
nand U3715 (N_3715,N_2387,N_2791);
nor U3716 (N_3716,N_2056,N_2544);
xnor U3717 (N_3717,N_2445,N_2722);
or U3718 (N_3718,N_2061,N_2086);
and U3719 (N_3719,N_2354,N_2374);
nor U3720 (N_3720,N_2263,N_2744);
or U3721 (N_3721,N_2601,N_2949);
nand U3722 (N_3722,N_2625,N_2199);
xnor U3723 (N_3723,N_2842,N_2110);
or U3724 (N_3724,N_2844,N_2474);
nor U3725 (N_3725,N_2370,N_2381);
and U3726 (N_3726,N_2708,N_2824);
or U3727 (N_3727,N_2464,N_2194);
and U3728 (N_3728,N_2826,N_2412);
xor U3729 (N_3729,N_2188,N_2659);
nand U3730 (N_3730,N_2989,N_2869);
nand U3731 (N_3731,N_2093,N_2996);
nor U3732 (N_3732,N_2117,N_2984);
xnor U3733 (N_3733,N_2416,N_2685);
nand U3734 (N_3734,N_2230,N_2263);
and U3735 (N_3735,N_2386,N_2566);
or U3736 (N_3736,N_2551,N_2895);
and U3737 (N_3737,N_2615,N_2390);
and U3738 (N_3738,N_2970,N_2509);
and U3739 (N_3739,N_2591,N_2163);
nand U3740 (N_3740,N_2586,N_2785);
or U3741 (N_3741,N_2494,N_2534);
or U3742 (N_3742,N_2608,N_2776);
and U3743 (N_3743,N_2798,N_2653);
nor U3744 (N_3744,N_2264,N_2362);
nand U3745 (N_3745,N_2035,N_2718);
nor U3746 (N_3746,N_2442,N_2905);
and U3747 (N_3747,N_2748,N_2400);
nand U3748 (N_3748,N_2133,N_2089);
or U3749 (N_3749,N_2221,N_2586);
or U3750 (N_3750,N_2094,N_2194);
nor U3751 (N_3751,N_2883,N_2990);
xnor U3752 (N_3752,N_2082,N_2703);
and U3753 (N_3753,N_2872,N_2285);
nor U3754 (N_3754,N_2053,N_2908);
nand U3755 (N_3755,N_2112,N_2300);
and U3756 (N_3756,N_2493,N_2225);
and U3757 (N_3757,N_2251,N_2396);
xor U3758 (N_3758,N_2669,N_2978);
nor U3759 (N_3759,N_2445,N_2304);
nand U3760 (N_3760,N_2726,N_2562);
nand U3761 (N_3761,N_2763,N_2875);
or U3762 (N_3762,N_2941,N_2764);
or U3763 (N_3763,N_2310,N_2540);
nor U3764 (N_3764,N_2373,N_2681);
or U3765 (N_3765,N_2196,N_2041);
or U3766 (N_3766,N_2646,N_2476);
nor U3767 (N_3767,N_2214,N_2684);
xor U3768 (N_3768,N_2003,N_2822);
xnor U3769 (N_3769,N_2276,N_2287);
and U3770 (N_3770,N_2668,N_2547);
and U3771 (N_3771,N_2257,N_2341);
or U3772 (N_3772,N_2758,N_2197);
nor U3773 (N_3773,N_2721,N_2153);
and U3774 (N_3774,N_2126,N_2654);
nor U3775 (N_3775,N_2912,N_2060);
and U3776 (N_3776,N_2106,N_2306);
nand U3777 (N_3777,N_2586,N_2719);
and U3778 (N_3778,N_2666,N_2001);
nand U3779 (N_3779,N_2914,N_2961);
nor U3780 (N_3780,N_2098,N_2032);
nand U3781 (N_3781,N_2269,N_2652);
or U3782 (N_3782,N_2971,N_2058);
or U3783 (N_3783,N_2977,N_2416);
xnor U3784 (N_3784,N_2236,N_2364);
and U3785 (N_3785,N_2340,N_2997);
nand U3786 (N_3786,N_2221,N_2615);
nor U3787 (N_3787,N_2253,N_2813);
nor U3788 (N_3788,N_2249,N_2503);
and U3789 (N_3789,N_2993,N_2474);
nand U3790 (N_3790,N_2574,N_2086);
or U3791 (N_3791,N_2745,N_2543);
or U3792 (N_3792,N_2443,N_2988);
xor U3793 (N_3793,N_2828,N_2226);
xnor U3794 (N_3794,N_2540,N_2562);
or U3795 (N_3795,N_2990,N_2621);
xnor U3796 (N_3796,N_2609,N_2117);
nor U3797 (N_3797,N_2704,N_2103);
nand U3798 (N_3798,N_2013,N_2919);
and U3799 (N_3799,N_2482,N_2837);
xnor U3800 (N_3800,N_2849,N_2295);
nand U3801 (N_3801,N_2152,N_2844);
nand U3802 (N_3802,N_2965,N_2244);
or U3803 (N_3803,N_2902,N_2359);
xnor U3804 (N_3804,N_2435,N_2282);
nand U3805 (N_3805,N_2528,N_2322);
or U3806 (N_3806,N_2544,N_2899);
xnor U3807 (N_3807,N_2778,N_2634);
or U3808 (N_3808,N_2186,N_2383);
nor U3809 (N_3809,N_2135,N_2341);
or U3810 (N_3810,N_2964,N_2358);
nor U3811 (N_3811,N_2526,N_2330);
nand U3812 (N_3812,N_2479,N_2243);
and U3813 (N_3813,N_2960,N_2035);
and U3814 (N_3814,N_2102,N_2076);
nand U3815 (N_3815,N_2873,N_2718);
nand U3816 (N_3816,N_2286,N_2583);
and U3817 (N_3817,N_2733,N_2777);
xor U3818 (N_3818,N_2535,N_2845);
and U3819 (N_3819,N_2776,N_2989);
nand U3820 (N_3820,N_2536,N_2834);
and U3821 (N_3821,N_2542,N_2240);
and U3822 (N_3822,N_2820,N_2861);
and U3823 (N_3823,N_2605,N_2009);
and U3824 (N_3824,N_2383,N_2606);
nand U3825 (N_3825,N_2726,N_2332);
nand U3826 (N_3826,N_2810,N_2101);
nand U3827 (N_3827,N_2626,N_2431);
or U3828 (N_3828,N_2410,N_2727);
nand U3829 (N_3829,N_2178,N_2797);
xnor U3830 (N_3830,N_2738,N_2904);
or U3831 (N_3831,N_2333,N_2399);
and U3832 (N_3832,N_2021,N_2305);
or U3833 (N_3833,N_2183,N_2007);
or U3834 (N_3834,N_2904,N_2274);
and U3835 (N_3835,N_2193,N_2502);
or U3836 (N_3836,N_2855,N_2300);
xnor U3837 (N_3837,N_2495,N_2365);
or U3838 (N_3838,N_2471,N_2090);
nor U3839 (N_3839,N_2484,N_2209);
or U3840 (N_3840,N_2951,N_2115);
nand U3841 (N_3841,N_2727,N_2583);
xor U3842 (N_3842,N_2524,N_2287);
and U3843 (N_3843,N_2502,N_2168);
nand U3844 (N_3844,N_2588,N_2698);
xnor U3845 (N_3845,N_2903,N_2338);
or U3846 (N_3846,N_2047,N_2871);
and U3847 (N_3847,N_2588,N_2914);
and U3848 (N_3848,N_2676,N_2377);
nand U3849 (N_3849,N_2393,N_2356);
nand U3850 (N_3850,N_2727,N_2052);
nor U3851 (N_3851,N_2665,N_2142);
nand U3852 (N_3852,N_2624,N_2872);
and U3853 (N_3853,N_2323,N_2554);
and U3854 (N_3854,N_2076,N_2474);
and U3855 (N_3855,N_2910,N_2816);
and U3856 (N_3856,N_2281,N_2516);
nand U3857 (N_3857,N_2044,N_2619);
or U3858 (N_3858,N_2871,N_2169);
and U3859 (N_3859,N_2370,N_2739);
and U3860 (N_3860,N_2612,N_2984);
or U3861 (N_3861,N_2004,N_2039);
and U3862 (N_3862,N_2527,N_2522);
and U3863 (N_3863,N_2805,N_2771);
nand U3864 (N_3864,N_2242,N_2389);
or U3865 (N_3865,N_2495,N_2268);
nand U3866 (N_3866,N_2731,N_2975);
or U3867 (N_3867,N_2017,N_2469);
and U3868 (N_3868,N_2033,N_2903);
nor U3869 (N_3869,N_2411,N_2805);
or U3870 (N_3870,N_2421,N_2522);
nor U3871 (N_3871,N_2158,N_2599);
nand U3872 (N_3872,N_2574,N_2210);
or U3873 (N_3873,N_2152,N_2025);
or U3874 (N_3874,N_2085,N_2422);
nor U3875 (N_3875,N_2968,N_2454);
and U3876 (N_3876,N_2879,N_2773);
nor U3877 (N_3877,N_2173,N_2853);
or U3878 (N_3878,N_2027,N_2023);
or U3879 (N_3879,N_2412,N_2531);
xor U3880 (N_3880,N_2099,N_2247);
xor U3881 (N_3881,N_2544,N_2355);
and U3882 (N_3882,N_2718,N_2639);
and U3883 (N_3883,N_2256,N_2353);
nor U3884 (N_3884,N_2397,N_2032);
xnor U3885 (N_3885,N_2138,N_2532);
or U3886 (N_3886,N_2799,N_2611);
xnor U3887 (N_3887,N_2115,N_2268);
xnor U3888 (N_3888,N_2838,N_2169);
nand U3889 (N_3889,N_2928,N_2751);
and U3890 (N_3890,N_2768,N_2062);
nand U3891 (N_3891,N_2607,N_2997);
xnor U3892 (N_3892,N_2012,N_2886);
xnor U3893 (N_3893,N_2705,N_2004);
or U3894 (N_3894,N_2884,N_2686);
or U3895 (N_3895,N_2487,N_2801);
nor U3896 (N_3896,N_2038,N_2794);
or U3897 (N_3897,N_2040,N_2415);
and U3898 (N_3898,N_2151,N_2563);
xnor U3899 (N_3899,N_2552,N_2456);
nor U3900 (N_3900,N_2251,N_2023);
and U3901 (N_3901,N_2169,N_2380);
nand U3902 (N_3902,N_2887,N_2889);
xor U3903 (N_3903,N_2981,N_2524);
and U3904 (N_3904,N_2238,N_2747);
or U3905 (N_3905,N_2135,N_2171);
and U3906 (N_3906,N_2900,N_2090);
xor U3907 (N_3907,N_2627,N_2036);
nor U3908 (N_3908,N_2555,N_2067);
and U3909 (N_3909,N_2211,N_2515);
or U3910 (N_3910,N_2480,N_2946);
and U3911 (N_3911,N_2119,N_2183);
xor U3912 (N_3912,N_2361,N_2746);
xor U3913 (N_3913,N_2666,N_2699);
and U3914 (N_3914,N_2771,N_2467);
and U3915 (N_3915,N_2184,N_2107);
or U3916 (N_3916,N_2353,N_2566);
nand U3917 (N_3917,N_2630,N_2380);
xor U3918 (N_3918,N_2663,N_2630);
xor U3919 (N_3919,N_2348,N_2056);
xnor U3920 (N_3920,N_2886,N_2041);
and U3921 (N_3921,N_2074,N_2068);
nor U3922 (N_3922,N_2746,N_2784);
nand U3923 (N_3923,N_2284,N_2323);
or U3924 (N_3924,N_2002,N_2477);
nand U3925 (N_3925,N_2129,N_2720);
nand U3926 (N_3926,N_2745,N_2211);
nand U3927 (N_3927,N_2969,N_2667);
or U3928 (N_3928,N_2500,N_2110);
nand U3929 (N_3929,N_2284,N_2438);
and U3930 (N_3930,N_2691,N_2039);
and U3931 (N_3931,N_2698,N_2754);
xnor U3932 (N_3932,N_2550,N_2195);
xnor U3933 (N_3933,N_2654,N_2580);
nand U3934 (N_3934,N_2992,N_2858);
xor U3935 (N_3935,N_2374,N_2405);
and U3936 (N_3936,N_2790,N_2975);
and U3937 (N_3937,N_2905,N_2464);
or U3938 (N_3938,N_2853,N_2691);
nor U3939 (N_3939,N_2440,N_2724);
and U3940 (N_3940,N_2286,N_2962);
and U3941 (N_3941,N_2447,N_2027);
and U3942 (N_3942,N_2513,N_2224);
xnor U3943 (N_3943,N_2944,N_2141);
or U3944 (N_3944,N_2921,N_2475);
xnor U3945 (N_3945,N_2594,N_2169);
and U3946 (N_3946,N_2385,N_2360);
or U3947 (N_3947,N_2307,N_2052);
or U3948 (N_3948,N_2470,N_2728);
nand U3949 (N_3949,N_2913,N_2101);
and U3950 (N_3950,N_2635,N_2561);
nor U3951 (N_3951,N_2435,N_2407);
and U3952 (N_3952,N_2730,N_2540);
nand U3953 (N_3953,N_2749,N_2827);
nand U3954 (N_3954,N_2469,N_2405);
and U3955 (N_3955,N_2331,N_2340);
nand U3956 (N_3956,N_2606,N_2013);
xor U3957 (N_3957,N_2177,N_2048);
or U3958 (N_3958,N_2155,N_2536);
nand U3959 (N_3959,N_2670,N_2810);
nor U3960 (N_3960,N_2585,N_2050);
xor U3961 (N_3961,N_2004,N_2865);
or U3962 (N_3962,N_2956,N_2076);
nand U3963 (N_3963,N_2333,N_2839);
and U3964 (N_3964,N_2199,N_2462);
or U3965 (N_3965,N_2227,N_2862);
nor U3966 (N_3966,N_2533,N_2160);
nor U3967 (N_3967,N_2132,N_2963);
xor U3968 (N_3968,N_2274,N_2817);
and U3969 (N_3969,N_2985,N_2628);
and U3970 (N_3970,N_2897,N_2448);
or U3971 (N_3971,N_2735,N_2607);
nand U3972 (N_3972,N_2457,N_2418);
and U3973 (N_3973,N_2287,N_2283);
nand U3974 (N_3974,N_2619,N_2607);
and U3975 (N_3975,N_2190,N_2879);
and U3976 (N_3976,N_2589,N_2628);
xor U3977 (N_3977,N_2460,N_2696);
or U3978 (N_3978,N_2405,N_2384);
xor U3979 (N_3979,N_2181,N_2499);
nand U3980 (N_3980,N_2019,N_2455);
xor U3981 (N_3981,N_2743,N_2235);
xnor U3982 (N_3982,N_2128,N_2405);
and U3983 (N_3983,N_2544,N_2595);
or U3984 (N_3984,N_2021,N_2357);
and U3985 (N_3985,N_2139,N_2672);
or U3986 (N_3986,N_2144,N_2923);
xor U3987 (N_3987,N_2071,N_2050);
nor U3988 (N_3988,N_2082,N_2737);
xor U3989 (N_3989,N_2468,N_2471);
or U3990 (N_3990,N_2425,N_2901);
nor U3991 (N_3991,N_2810,N_2165);
xnor U3992 (N_3992,N_2971,N_2309);
nand U3993 (N_3993,N_2078,N_2206);
nor U3994 (N_3994,N_2744,N_2527);
nand U3995 (N_3995,N_2238,N_2197);
xor U3996 (N_3996,N_2498,N_2261);
or U3997 (N_3997,N_2983,N_2805);
or U3998 (N_3998,N_2759,N_2172);
xnor U3999 (N_3999,N_2222,N_2270);
or U4000 (N_4000,N_3194,N_3617);
nor U4001 (N_4001,N_3302,N_3761);
nand U4002 (N_4002,N_3718,N_3815);
or U4003 (N_4003,N_3583,N_3265);
nor U4004 (N_4004,N_3851,N_3945);
nand U4005 (N_4005,N_3448,N_3844);
xor U4006 (N_4006,N_3504,N_3779);
or U4007 (N_4007,N_3573,N_3404);
xor U4008 (N_4008,N_3665,N_3219);
nor U4009 (N_4009,N_3966,N_3681);
nand U4010 (N_4010,N_3956,N_3258);
and U4011 (N_4011,N_3816,N_3238);
xor U4012 (N_4012,N_3633,N_3214);
or U4013 (N_4013,N_3123,N_3324);
nor U4014 (N_4014,N_3057,N_3402);
and U4015 (N_4015,N_3961,N_3884);
or U4016 (N_4016,N_3616,N_3730);
nor U4017 (N_4017,N_3889,N_3874);
xnor U4018 (N_4018,N_3944,N_3178);
nor U4019 (N_4019,N_3352,N_3044);
and U4020 (N_4020,N_3077,N_3382);
nor U4021 (N_4021,N_3498,N_3133);
xnor U4022 (N_4022,N_3541,N_3016);
nand U4023 (N_4023,N_3818,N_3901);
or U4024 (N_4024,N_3054,N_3577);
nand U4025 (N_4025,N_3950,N_3925);
or U4026 (N_4026,N_3769,N_3872);
and U4027 (N_4027,N_3842,N_3042);
nand U4028 (N_4028,N_3393,N_3459);
and U4029 (N_4029,N_3273,N_3856);
or U4030 (N_4030,N_3240,N_3553);
and U4031 (N_4031,N_3788,N_3341);
or U4032 (N_4032,N_3752,N_3614);
xor U4033 (N_4033,N_3875,N_3415);
and U4034 (N_4034,N_3892,N_3557);
or U4035 (N_4035,N_3538,N_3795);
and U4036 (N_4036,N_3934,N_3174);
or U4037 (N_4037,N_3387,N_3430);
and U4038 (N_4038,N_3490,N_3411);
and U4039 (N_4039,N_3051,N_3540);
xor U4040 (N_4040,N_3787,N_3532);
or U4041 (N_4041,N_3671,N_3928);
xnor U4042 (N_4042,N_3218,N_3050);
or U4043 (N_4043,N_3331,N_3649);
and U4044 (N_4044,N_3880,N_3256);
xor U4045 (N_4045,N_3918,N_3740);
xor U4046 (N_4046,N_3068,N_3994);
nor U4047 (N_4047,N_3989,N_3590);
nand U4048 (N_4048,N_3386,N_3034);
and U4049 (N_4049,N_3786,N_3191);
nor U4050 (N_4050,N_3491,N_3919);
nand U4051 (N_4051,N_3987,N_3377);
xnor U4052 (N_4052,N_3164,N_3097);
and U4053 (N_4053,N_3328,N_3513);
nor U4054 (N_4054,N_3162,N_3579);
xnor U4055 (N_4055,N_3615,N_3335);
and U4056 (N_4056,N_3465,N_3172);
and U4057 (N_4057,N_3832,N_3243);
xnor U4058 (N_4058,N_3674,N_3713);
nor U4059 (N_4059,N_3467,N_3435);
xor U4060 (N_4060,N_3785,N_3609);
nand U4061 (N_4061,N_3252,N_3970);
or U4062 (N_4062,N_3662,N_3890);
nor U4063 (N_4063,N_3395,N_3206);
nand U4064 (N_4064,N_3018,N_3141);
nand U4065 (N_4065,N_3727,N_3200);
and U4066 (N_4066,N_3893,N_3486);
nand U4067 (N_4067,N_3547,N_3942);
nand U4068 (N_4068,N_3293,N_3575);
xnor U4069 (N_4069,N_3793,N_3555);
or U4070 (N_4070,N_3933,N_3120);
or U4071 (N_4071,N_3841,N_3332);
or U4072 (N_4072,N_3858,N_3298);
xnor U4073 (N_4073,N_3783,N_3110);
nor U4074 (N_4074,N_3263,N_3564);
or U4075 (N_4075,N_3909,N_3254);
xor U4076 (N_4076,N_3722,N_3804);
nand U4077 (N_4077,N_3952,N_3660);
nand U4078 (N_4078,N_3037,N_3518);
nand U4079 (N_4079,N_3572,N_3308);
and U4080 (N_4080,N_3007,N_3149);
xnor U4081 (N_4081,N_3439,N_3452);
or U4082 (N_4082,N_3210,N_3943);
nor U4083 (N_4083,N_3744,N_3669);
xor U4084 (N_4084,N_3724,N_3494);
nor U4085 (N_4085,N_3144,N_3843);
and U4086 (N_4086,N_3923,N_3554);
and U4087 (N_4087,N_3128,N_3005);
nor U4088 (N_4088,N_3136,N_3780);
nor U4089 (N_4089,N_3232,N_3963);
and U4090 (N_4090,N_3457,N_3319);
or U4091 (N_4091,N_3147,N_3087);
xor U4092 (N_4092,N_3536,N_3275);
or U4093 (N_4093,N_3621,N_3228);
xor U4094 (N_4094,N_3476,N_3433);
xnor U4095 (N_4095,N_3157,N_3589);
nor U4096 (N_4096,N_3262,N_3455);
nand U4097 (N_4097,N_3768,N_3221);
nor U4098 (N_4098,N_3215,N_3535);
xor U4099 (N_4099,N_3092,N_3188);
xnor U4100 (N_4100,N_3175,N_3721);
xor U4101 (N_4101,N_3608,N_3101);
nor U4102 (N_4102,N_3957,N_3654);
nor U4103 (N_4103,N_3114,N_3625);
or U4104 (N_4104,N_3138,N_3601);
xnor U4105 (N_4105,N_3686,N_3014);
xnor U4106 (N_4106,N_3571,N_3389);
nor U4107 (N_4107,N_3281,N_3846);
xor U4108 (N_4108,N_3807,N_3326);
nand U4109 (N_4109,N_3216,N_3205);
or U4110 (N_4110,N_3965,N_3720);
nand U4111 (N_4111,N_3260,N_3074);
xnor U4112 (N_4112,N_3552,N_3550);
nor U4113 (N_4113,N_3388,N_3269);
xor U4114 (N_4114,N_3531,N_3605);
nor U4115 (N_4115,N_3915,N_3775);
and U4116 (N_4116,N_3482,N_3090);
or U4117 (N_4117,N_3820,N_3480);
xor U4118 (N_4118,N_3829,N_3463);
and U4119 (N_4119,N_3121,N_3784);
nand U4120 (N_4120,N_3417,N_3597);
xnor U4121 (N_4121,N_3938,N_3198);
nor U4122 (N_4122,N_3249,N_3211);
nor U4123 (N_4123,N_3733,N_3567);
nand U4124 (N_4124,N_3351,N_3071);
xor U4125 (N_4125,N_3270,N_3861);
and U4126 (N_4126,N_3599,N_3237);
and U4127 (N_4127,N_3305,N_3049);
xnor U4128 (N_4128,N_3641,N_3380);
or U4129 (N_4129,N_3363,N_3119);
nand U4130 (N_4130,N_3209,N_3073);
and U4131 (N_4131,N_3821,N_3137);
nand U4132 (N_4132,N_3409,N_3507);
nor U4133 (N_4133,N_3063,N_3481);
xnor U4134 (N_4134,N_3863,N_3008);
or U4135 (N_4135,N_3544,N_3698);
nand U4136 (N_4136,N_3406,N_3062);
nor U4137 (N_4137,N_3977,N_3171);
or U4138 (N_4138,N_3568,N_3080);
and U4139 (N_4139,N_3757,N_3383);
nor U4140 (N_4140,N_3003,N_3358);
and U4141 (N_4141,N_3349,N_3885);
and U4142 (N_4142,N_3125,N_3810);
nand U4143 (N_4143,N_3290,N_3212);
xor U4144 (N_4144,N_3093,N_3576);
nand U4145 (N_4145,N_3401,N_3551);
nand U4146 (N_4146,N_3700,N_3109);
nand U4147 (N_4147,N_3496,N_3562);
nand U4148 (N_4148,N_3581,N_3372);
and U4149 (N_4149,N_3196,N_3508);
or U4150 (N_4150,N_3244,N_3190);
nor U4151 (N_4151,N_3545,N_3759);
or U4152 (N_4152,N_3017,N_3585);
nand U4153 (N_4153,N_3607,N_3202);
and U4154 (N_4154,N_3524,N_3279);
nor U4155 (N_4155,N_3794,N_3366);
and U4156 (N_4156,N_3808,N_3195);
nand U4157 (N_4157,N_3767,N_3812);
or U4158 (N_4158,N_3189,N_3484);
nor U4159 (N_4159,N_3865,N_3587);
or U4160 (N_4160,N_3748,N_3542);
nand U4161 (N_4161,N_3822,N_3135);
or U4162 (N_4162,N_3170,N_3280);
nand U4163 (N_4163,N_3651,N_3830);
xnor U4164 (N_4164,N_3592,N_3058);
xnor U4165 (N_4165,N_3040,N_3847);
or U4166 (N_4166,N_3334,N_3983);
xnor U4167 (N_4167,N_3255,N_3056);
or U4168 (N_4168,N_3461,N_3353);
xnor U4169 (N_4169,N_3303,N_3514);
and U4170 (N_4170,N_3320,N_3610);
nand U4171 (N_4171,N_3558,N_3711);
nor U4172 (N_4172,N_3339,N_3373);
and U4173 (N_4173,N_3392,N_3053);
nor U4174 (N_4174,N_3168,N_3760);
and U4175 (N_4175,N_3796,N_3870);
nand U4176 (N_4176,N_3248,N_3647);
or U4177 (N_4177,N_3356,N_3828);
or U4178 (N_4178,N_3852,N_3012);
or U4179 (N_4179,N_3111,N_3520);
xnor U4180 (N_4180,N_3338,N_3414);
and U4181 (N_4181,N_3595,N_3370);
or U4182 (N_4182,N_3580,N_3732);
or U4183 (N_4183,N_3112,N_3864);
nand U4184 (N_4184,N_3150,N_3337);
and U4185 (N_4185,N_3396,N_3464);
xor U4186 (N_4186,N_3516,N_3035);
and U4187 (N_4187,N_3611,N_3505);
and U4188 (N_4188,N_3530,N_3526);
or U4189 (N_4189,N_3510,N_3905);
and U4190 (N_4190,N_3735,N_3483);
or U4191 (N_4191,N_3184,N_3407);
xor U4192 (N_4192,N_3327,N_3503);
xnor U4193 (N_4193,N_3365,N_3563);
or U4194 (N_4194,N_3898,N_3878);
and U4195 (N_4195,N_3183,N_3257);
nand U4196 (N_4196,N_3418,N_3177);
and U4197 (N_4197,N_3499,N_3475);
and U4198 (N_4198,N_3038,N_3517);
or U4199 (N_4199,N_3441,N_3911);
or U4200 (N_4200,N_3083,N_3466);
and U4201 (N_4201,N_3811,N_3291);
or U4202 (N_4202,N_3375,N_3586);
nand U4203 (N_4203,N_3770,N_3271);
nor U4204 (N_4204,N_3102,N_3048);
xnor U4205 (N_4205,N_3225,N_3741);
or U4206 (N_4206,N_3648,N_3222);
nand U4207 (N_4207,N_3296,N_3376);
nor U4208 (N_4208,N_3019,N_3817);
xnor U4209 (N_4209,N_3234,N_3330);
and U4210 (N_4210,N_3468,N_3207);
or U4211 (N_4211,N_3569,N_3653);
nor U4212 (N_4212,N_3106,N_3941);
xor U4213 (N_4213,N_3477,N_3329);
and U4214 (N_4214,N_3004,N_3310);
nor U4215 (N_4215,N_3699,N_3714);
or U4216 (N_4216,N_3831,N_3716);
nand U4217 (N_4217,N_3313,N_3600);
and U4218 (N_4218,N_3130,N_3511);
nor U4219 (N_4219,N_3955,N_3186);
nand U4220 (N_4220,N_3076,N_3251);
nor U4221 (N_4221,N_3447,N_3061);
nand U4222 (N_4222,N_3519,N_3914);
and U4223 (N_4223,N_3845,N_3619);
and U4224 (N_4224,N_3277,N_3922);
nor U4225 (N_4225,N_3677,N_3999);
nand U4226 (N_4226,N_3613,N_3436);
and U4227 (N_4227,N_3990,N_3984);
nand U4228 (N_4228,N_3782,N_3322);
and U4229 (N_4229,N_3937,N_3045);
nor U4230 (N_4230,N_3756,N_3837);
and U4231 (N_4231,N_3242,N_3294);
nor U4232 (N_4232,N_3738,N_3179);
and U4233 (N_4233,N_3927,N_3932);
nor U4234 (N_4234,N_3646,N_3412);
and U4235 (N_4235,N_3778,N_3947);
nor U4236 (N_4236,N_3013,N_3838);
nor U4237 (N_4237,N_3458,N_3917);
nor U4238 (N_4238,N_3088,N_3960);
nor U4239 (N_4239,N_3082,N_3622);
and U4240 (N_4240,N_3113,N_3070);
nand U4241 (N_4241,N_3105,N_3543);
or U4242 (N_4242,N_3336,N_3318);
nor U4243 (N_4243,N_3390,N_3340);
xnor U4244 (N_4244,N_3728,N_3166);
nor U4245 (N_4245,N_3416,N_3187);
and U4246 (N_4246,N_3247,N_3980);
xnor U4247 (N_4247,N_3301,N_3284);
nand U4248 (N_4248,N_3185,N_3848);
or U4249 (N_4249,N_3169,N_3156);
nor U4250 (N_4250,N_3855,N_3378);
or U4251 (N_4251,N_3427,N_3763);
xor U4252 (N_4252,N_3515,N_3497);
nand U4253 (N_4253,N_3897,N_3473);
and U4254 (N_4254,N_3895,N_3274);
xnor U4255 (N_4255,N_3684,N_3454);
nand U4256 (N_4256,N_3635,N_3286);
xnor U4257 (N_4257,N_3143,N_3501);
or U4258 (N_4258,N_3276,N_3537);
nand U4259 (N_4259,N_3866,N_3750);
or U4260 (N_4260,N_3814,N_3470);
xnor U4261 (N_4261,N_3574,N_3687);
nand U4262 (N_4262,N_3636,N_3432);
xnor U4263 (N_4263,N_3835,N_3694);
and U4264 (N_4264,N_3367,N_3624);
xnor U4265 (N_4265,N_3086,N_3420);
xor U4266 (N_4266,N_3869,N_3239);
nand U4267 (N_4267,N_3026,N_3797);
nor U4268 (N_4268,N_3798,N_3643);
xnor U4269 (N_4269,N_3072,N_3949);
nor U4270 (N_4270,N_3772,N_3827);
nor U4271 (N_4271,N_3596,N_3776);
nor U4272 (N_4272,N_3158,N_3962);
or U4273 (N_4273,N_3904,N_3145);
or U4274 (N_4274,N_3116,N_3066);
nand U4275 (N_4275,N_3493,N_3295);
nand U4276 (N_4276,N_3031,N_3246);
nor U4277 (N_4277,N_3731,N_3361);
or U4278 (N_4278,N_3055,N_3556);
nor U4279 (N_4279,N_3697,N_3737);
and U4280 (N_4280,N_3023,N_3431);
xnor U4281 (N_4281,N_3449,N_3032);
nand U4282 (N_4282,N_3217,N_3405);
nor U4283 (N_4283,N_3836,N_3472);
xor U4284 (N_4284,N_3523,N_3098);
xnor U4285 (N_4285,N_3900,N_3969);
xnor U4286 (N_4286,N_3314,N_3781);
or U4287 (N_4287,N_3444,N_3774);
nor U4288 (N_4288,N_3434,N_3509);
nor U4289 (N_4289,N_3132,N_3566);
nand U4290 (N_4290,N_3877,N_3385);
xnor U4291 (N_4291,N_3203,N_3959);
nor U4292 (N_4292,N_3020,N_3084);
nand U4293 (N_4293,N_3789,N_3879);
or U4294 (N_4294,N_3805,N_3312);
nand U4295 (N_4295,N_3115,N_3299);
nand U4296 (N_4296,N_3939,N_3549);
and U4297 (N_4297,N_3655,N_3139);
xor U4298 (N_4298,N_3024,N_3039);
and U4299 (N_4299,N_3025,N_3134);
and U4300 (N_4300,N_3495,N_3471);
and U4301 (N_4301,N_3940,N_3899);
nand U4302 (N_4302,N_3428,N_3771);
or U4303 (N_4303,N_3155,N_3002);
nor U4304 (N_4304,N_3642,N_3272);
or U4305 (N_4305,N_3675,N_3445);
nor U4306 (N_4306,N_3381,N_3717);
and U4307 (N_4307,N_3981,N_3148);
nand U4308 (N_4308,N_3803,N_3704);
or U4309 (N_4309,N_3854,N_3991);
or U4310 (N_4310,N_3930,N_3951);
and U4311 (N_4311,N_3165,N_3259);
and U4312 (N_4312,N_3403,N_3231);
nand U4313 (N_4313,N_3400,N_3664);
nor U4314 (N_4314,N_3423,N_3751);
or U4315 (N_4315,N_3973,N_3637);
nand U4316 (N_4316,N_3287,N_3588);
xnor U4317 (N_4317,N_3348,N_3935);
or U4318 (N_4318,N_3146,N_3690);
nand U4319 (N_4319,N_3089,N_3630);
xor U4320 (N_4320,N_3891,N_3657);
nand U4321 (N_4321,N_3982,N_3634);
nor U4322 (N_4322,N_3626,N_3350);
and U4323 (N_4323,N_3343,N_3456);
xor U4324 (N_4324,N_3371,N_3443);
nand U4325 (N_4325,N_3819,N_3369);
xnor U4326 (N_4326,N_3708,N_3230);
xor U4327 (N_4327,N_3000,N_3355);
nor U4328 (N_4328,N_3297,N_3691);
and U4329 (N_4329,N_3606,N_3236);
or U4330 (N_4330,N_3670,N_3809);
nand U4331 (N_4331,N_3006,N_3422);
xnor U4332 (N_4332,N_3309,N_3478);
or U4333 (N_4333,N_3469,N_3502);
nand U4334 (N_4334,N_3992,N_3739);
nand U4335 (N_4335,N_3201,N_3027);
or U4336 (N_4336,N_3283,N_3176);
or U4337 (N_4337,N_3902,N_3565);
nor U4338 (N_4338,N_3632,N_3644);
and U4339 (N_4339,N_3397,N_3096);
nand U4340 (N_4340,N_3753,N_3548);
and U4341 (N_4341,N_3362,N_3533);
or U4342 (N_4342,N_3612,N_3292);
nor U4343 (N_4343,N_3791,N_3103);
nand U4344 (N_4344,N_3224,N_3010);
or U4345 (N_4345,N_3603,N_3715);
or U4346 (N_4346,N_3180,N_3873);
and U4347 (N_4347,N_3824,N_3823);
or U4348 (N_4348,N_3140,N_3451);
nand U4349 (N_4349,N_3075,N_3223);
nand U4350 (N_4350,N_3325,N_3527);
and U4351 (N_4351,N_3680,N_3976);
nand U4352 (N_4352,N_3594,N_3289);
and U4353 (N_4353,N_3931,N_3755);
xor U4354 (N_4354,N_3792,N_3682);
nand U4355 (N_4355,N_3220,N_3883);
or U4356 (N_4356,N_3163,N_3399);
nor U4357 (N_4357,N_3546,N_3153);
nor U4358 (N_4358,N_3182,N_3489);
nor U4359 (N_4359,N_3921,N_3894);
nor U4360 (N_4360,N_3410,N_3208);
nor U4361 (N_4361,N_3813,N_3602);
nor U4362 (N_4362,N_3881,N_3344);
xnor U4363 (N_4363,N_3316,N_3702);
and U4364 (N_4364,N_3656,N_3029);
and U4365 (N_4365,N_3910,N_3627);
nand U4366 (N_4366,N_3154,N_3867);
and U4367 (N_4367,N_3300,N_3342);
xnor U4368 (N_4368,N_3995,N_3620);
and U4369 (N_4369,N_3692,N_3913);
and U4370 (N_4370,N_3379,N_3001);
xnor U4371 (N_4371,N_3307,N_3850);
nand U4372 (N_4372,N_3623,N_3022);
nand U4373 (N_4373,N_3746,N_3181);
nor U4374 (N_4374,N_3802,N_3974);
xnor U4375 (N_4375,N_3317,N_3946);
or U4376 (N_4376,N_3213,N_3777);
nand U4377 (N_4377,N_3266,N_3512);
nand U4378 (N_4378,N_3161,N_3685);
and U4379 (N_4379,N_3559,N_3888);
xor U4380 (N_4380,N_3398,N_3360);
nand U4381 (N_4381,N_3639,N_3354);
xnor U4382 (N_4382,N_3368,N_3253);
and U4383 (N_4383,N_3081,N_3652);
or U4384 (N_4384,N_3985,N_3100);
nor U4385 (N_4385,N_3964,N_3359);
nor U4386 (N_4386,N_3673,N_3726);
nand U4387 (N_4387,N_3453,N_3167);
or U4388 (N_4388,N_3046,N_3764);
and U4389 (N_4389,N_3064,N_3906);
xor U4390 (N_4390,N_3226,N_3429);
and U4391 (N_4391,N_3345,N_3506);
nand U4392 (N_4392,N_3041,N_3015);
and U4393 (N_4393,N_3241,N_3678);
nand U4394 (N_4394,N_3446,N_3725);
and U4395 (N_4395,N_3419,N_3306);
and U4396 (N_4396,N_3790,N_3159);
nor U4397 (N_4397,N_3107,N_3800);
or U4398 (N_4398,N_3578,N_3408);
and U4399 (N_4399,N_3268,N_3421);
nand U4400 (N_4400,N_3672,N_3570);
nand U4401 (N_4401,N_3975,N_3347);
or U4402 (N_4402,N_3640,N_3924);
or U4403 (N_4403,N_3009,N_3912);
nand U4404 (N_4404,N_3229,N_3839);
or U4405 (N_4405,N_3043,N_3127);
nand U4406 (N_4406,N_3747,N_3060);
nand U4407 (N_4407,N_3122,N_3525);
nand U4408 (N_4408,N_3849,N_3696);
xor U4409 (N_4409,N_3374,N_3108);
nand U4410 (N_4410,N_3245,N_3462);
nor U4411 (N_4411,N_3709,N_3560);
and U4412 (N_4412,N_3719,N_3773);
or U4413 (N_4413,N_3492,N_3591);
and U4414 (N_4414,N_3998,N_3742);
nand U4415 (N_4415,N_3668,N_3069);
or U4416 (N_4416,N_3500,N_3391);
nand U4417 (N_4417,N_3199,N_3903);
xnor U4418 (N_4418,N_3065,N_3971);
nor U4419 (N_4419,N_3124,N_3754);
xor U4420 (N_4420,N_3264,N_3979);
or U4421 (N_4421,N_3749,N_3118);
and U4422 (N_4422,N_3978,N_3126);
xor U4423 (N_4423,N_3826,N_3907);
and U4424 (N_4424,N_3871,N_3896);
and U4425 (N_4425,N_3047,N_3765);
xnor U4426 (N_4426,N_3701,N_3059);
xnor U4427 (N_4427,N_3233,N_3658);
or U4428 (N_4428,N_3703,N_3676);
nor U4429 (N_4429,N_3321,N_3085);
nand U4430 (N_4430,N_3645,N_3629);
nor U4431 (N_4431,N_3282,N_3598);
xnor U4432 (N_4432,N_3972,N_3986);
and U4433 (N_4433,N_3679,N_3650);
nand U4434 (N_4434,N_3534,N_3887);
xnor U4435 (N_4435,N_3099,N_3712);
xnor U4436 (N_4436,N_3384,N_3235);
nand U4437 (N_4437,N_3173,N_3033);
nor U4438 (N_4438,N_3474,N_3323);
nor U4439 (N_4439,N_3425,N_3996);
and U4440 (N_4440,N_3707,N_3160);
nand U4441 (N_4441,N_3584,N_3857);
xnor U4442 (N_4442,N_3723,N_3993);
xor U4443 (N_4443,N_3052,N_3197);
and U4444 (N_4444,N_3091,N_3346);
nand U4445 (N_4445,N_3736,N_3364);
xor U4446 (N_4446,N_3604,N_3860);
xor U4447 (N_4447,N_3104,N_3948);
nand U4448 (N_4448,N_3193,N_3333);
xor U4449 (N_4449,N_3840,N_3710);
nor U4450 (N_4450,N_3442,N_3485);
and U4451 (N_4451,N_3638,N_3954);
nand U4452 (N_4452,N_3862,N_3689);
xor U4453 (N_4453,N_3488,N_3916);
xor U4454 (N_4454,N_3868,N_3582);
nand U4455 (N_4455,N_3859,N_3997);
or U4456 (N_4456,N_3036,N_3618);
nor U4457 (N_4457,N_3521,N_3304);
nand U4458 (N_4458,N_3278,N_3967);
xor U4459 (N_4459,N_3762,N_3394);
and U4460 (N_4460,N_3631,N_3659);
or U4461 (N_4461,N_3683,N_3729);
or U4462 (N_4462,N_3357,N_3920);
xnor U4463 (N_4463,N_3479,N_3663);
or U4464 (N_4464,N_3825,N_3834);
nor U4465 (N_4465,N_3021,N_3250);
xor U4466 (N_4466,N_3288,N_3261);
nor U4467 (N_4467,N_3926,N_3094);
nor U4468 (N_4468,N_3267,N_3539);
nor U4469 (N_4469,N_3745,N_3666);
xor U4470 (N_4470,N_3882,N_3192);
and U4471 (N_4471,N_3437,N_3936);
nor U4472 (N_4472,N_3438,N_3953);
nand U4473 (N_4473,N_3311,N_3667);
nand U4474 (N_4474,N_3929,N_3011);
nand U4475 (N_4475,N_3853,N_3030);
xor U4476 (N_4476,N_3426,N_3988);
and U4477 (N_4477,N_3450,N_3695);
and U4478 (N_4478,N_3152,N_3522);
nor U4479 (N_4479,N_3529,N_3628);
xor U4480 (N_4480,N_3028,N_3705);
nor U4481 (N_4481,N_3285,N_3413);
nand U4482 (N_4482,N_3706,N_3688);
nand U4483 (N_4483,N_3693,N_3886);
and U4484 (N_4484,N_3460,N_3440);
nor U4485 (N_4485,N_3131,N_3315);
nor U4486 (N_4486,N_3151,N_3129);
and U4487 (N_4487,N_3876,N_3801);
and U4488 (N_4488,N_3117,N_3799);
nand U4489 (N_4489,N_3528,N_3078);
nor U4490 (N_4490,N_3067,N_3734);
nand U4491 (N_4491,N_3095,N_3833);
xnor U4492 (N_4492,N_3758,N_3424);
nand U4493 (N_4493,N_3661,N_3743);
xor U4494 (N_4494,N_3487,N_3227);
xnor U4495 (N_4495,N_3958,N_3561);
or U4496 (N_4496,N_3079,N_3766);
xnor U4497 (N_4497,N_3806,N_3204);
or U4498 (N_4498,N_3968,N_3908);
nand U4499 (N_4499,N_3142,N_3593);
nand U4500 (N_4500,N_3324,N_3861);
and U4501 (N_4501,N_3146,N_3028);
xnor U4502 (N_4502,N_3584,N_3112);
or U4503 (N_4503,N_3244,N_3019);
and U4504 (N_4504,N_3809,N_3285);
xnor U4505 (N_4505,N_3870,N_3299);
and U4506 (N_4506,N_3063,N_3741);
or U4507 (N_4507,N_3728,N_3269);
nor U4508 (N_4508,N_3723,N_3022);
nand U4509 (N_4509,N_3014,N_3077);
or U4510 (N_4510,N_3788,N_3273);
nand U4511 (N_4511,N_3505,N_3317);
nor U4512 (N_4512,N_3484,N_3422);
nand U4513 (N_4513,N_3621,N_3425);
nand U4514 (N_4514,N_3653,N_3360);
and U4515 (N_4515,N_3698,N_3804);
nand U4516 (N_4516,N_3664,N_3849);
xor U4517 (N_4517,N_3400,N_3058);
xnor U4518 (N_4518,N_3893,N_3105);
nor U4519 (N_4519,N_3715,N_3553);
nand U4520 (N_4520,N_3550,N_3450);
xnor U4521 (N_4521,N_3721,N_3641);
and U4522 (N_4522,N_3744,N_3281);
or U4523 (N_4523,N_3048,N_3358);
nand U4524 (N_4524,N_3163,N_3395);
and U4525 (N_4525,N_3455,N_3186);
and U4526 (N_4526,N_3619,N_3030);
or U4527 (N_4527,N_3374,N_3176);
nor U4528 (N_4528,N_3492,N_3933);
nor U4529 (N_4529,N_3282,N_3093);
xnor U4530 (N_4530,N_3313,N_3805);
xnor U4531 (N_4531,N_3040,N_3825);
nand U4532 (N_4532,N_3039,N_3767);
xor U4533 (N_4533,N_3727,N_3882);
xnor U4534 (N_4534,N_3309,N_3143);
or U4535 (N_4535,N_3690,N_3790);
and U4536 (N_4536,N_3650,N_3338);
nor U4537 (N_4537,N_3052,N_3813);
xnor U4538 (N_4538,N_3805,N_3373);
or U4539 (N_4539,N_3033,N_3114);
and U4540 (N_4540,N_3492,N_3972);
nand U4541 (N_4541,N_3396,N_3617);
xnor U4542 (N_4542,N_3104,N_3170);
and U4543 (N_4543,N_3035,N_3673);
nor U4544 (N_4544,N_3244,N_3419);
nand U4545 (N_4545,N_3980,N_3865);
nor U4546 (N_4546,N_3610,N_3598);
xnor U4547 (N_4547,N_3796,N_3233);
or U4548 (N_4548,N_3172,N_3031);
xor U4549 (N_4549,N_3828,N_3533);
nor U4550 (N_4550,N_3223,N_3670);
nand U4551 (N_4551,N_3022,N_3087);
or U4552 (N_4552,N_3806,N_3382);
nor U4553 (N_4553,N_3292,N_3153);
or U4554 (N_4554,N_3468,N_3133);
nand U4555 (N_4555,N_3071,N_3664);
nor U4556 (N_4556,N_3476,N_3347);
nand U4557 (N_4557,N_3201,N_3123);
and U4558 (N_4558,N_3827,N_3835);
xnor U4559 (N_4559,N_3998,N_3918);
or U4560 (N_4560,N_3636,N_3858);
and U4561 (N_4561,N_3744,N_3737);
nand U4562 (N_4562,N_3094,N_3610);
and U4563 (N_4563,N_3521,N_3913);
nor U4564 (N_4564,N_3336,N_3622);
xnor U4565 (N_4565,N_3164,N_3265);
nor U4566 (N_4566,N_3641,N_3338);
xnor U4567 (N_4567,N_3268,N_3555);
or U4568 (N_4568,N_3968,N_3854);
or U4569 (N_4569,N_3144,N_3230);
and U4570 (N_4570,N_3552,N_3962);
nor U4571 (N_4571,N_3398,N_3352);
nand U4572 (N_4572,N_3875,N_3662);
nand U4573 (N_4573,N_3754,N_3405);
or U4574 (N_4574,N_3435,N_3930);
and U4575 (N_4575,N_3594,N_3253);
or U4576 (N_4576,N_3992,N_3492);
and U4577 (N_4577,N_3182,N_3934);
and U4578 (N_4578,N_3428,N_3606);
xnor U4579 (N_4579,N_3614,N_3935);
xor U4580 (N_4580,N_3168,N_3871);
xnor U4581 (N_4581,N_3759,N_3784);
xor U4582 (N_4582,N_3349,N_3117);
nor U4583 (N_4583,N_3221,N_3138);
xnor U4584 (N_4584,N_3317,N_3112);
nand U4585 (N_4585,N_3302,N_3452);
and U4586 (N_4586,N_3658,N_3567);
and U4587 (N_4587,N_3087,N_3049);
nand U4588 (N_4588,N_3906,N_3566);
nor U4589 (N_4589,N_3223,N_3140);
xnor U4590 (N_4590,N_3509,N_3349);
xnor U4591 (N_4591,N_3478,N_3859);
and U4592 (N_4592,N_3247,N_3406);
and U4593 (N_4593,N_3331,N_3021);
or U4594 (N_4594,N_3270,N_3399);
nand U4595 (N_4595,N_3583,N_3252);
and U4596 (N_4596,N_3170,N_3109);
and U4597 (N_4597,N_3481,N_3824);
nand U4598 (N_4598,N_3145,N_3479);
or U4599 (N_4599,N_3621,N_3679);
xnor U4600 (N_4600,N_3883,N_3672);
nor U4601 (N_4601,N_3882,N_3927);
xnor U4602 (N_4602,N_3818,N_3898);
nor U4603 (N_4603,N_3625,N_3453);
nand U4604 (N_4604,N_3668,N_3346);
xnor U4605 (N_4605,N_3019,N_3125);
or U4606 (N_4606,N_3096,N_3317);
nand U4607 (N_4607,N_3455,N_3719);
nand U4608 (N_4608,N_3675,N_3658);
nor U4609 (N_4609,N_3162,N_3356);
or U4610 (N_4610,N_3604,N_3508);
xor U4611 (N_4611,N_3516,N_3152);
xor U4612 (N_4612,N_3156,N_3189);
xnor U4613 (N_4613,N_3672,N_3086);
nor U4614 (N_4614,N_3787,N_3697);
nand U4615 (N_4615,N_3885,N_3090);
or U4616 (N_4616,N_3613,N_3490);
or U4617 (N_4617,N_3828,N_3006);
and U4618 (N_4618,N_3312,N_3814);
or U4619 (N_4619,N_3764,N_3941);
nor U4620 (N_4620,N_3456,N_3623);
and U4621 (N_4621,N_3842,N_3564);
and U4622 (N_4622,N_3035,N_3011);
nor U4623 (N_4623,N_3420,N_3589);
and U4624 (N_4624,N_3352,N_3451);
xnor U4625 (N_4625,N_3505,N_3700);
or U4626 (N_4626,N_3551,N_3122);
nor U4627 (N_4627,N_3563,N_3786);
nand U4628 (N_4628,N_3492,N_3450);
xor U4629 (N_4629,N_3340,N_3926);
nand U4630 (N_4630,N_3029,N_3104);
or U4631 (N_4631,N_3186,N_3154);
xor U4632 (N_4632,N_3444,N_3186);
or U4633 (N_4633,N_3312,N_3081);
nor U4634 (N_4634,N_3060,N_3214);
nor U4635 (N_4635,N_3382,N_3673);
nor U4636 (N_4636,N_3908,N_3177);
or U4637 (N_4637,N_3426,N_3356);
nor U4638 (N_4638,N_3148,N_3280);
nor U4639 (N_4639,N_3159,N_3634);
nand U4640 (N_4640,N_3887,N_3239);
xor U4641 (N_4641,N_3808,N_3291);
and U4642 (N_4642,N_3647,N_3835);
nand U4643 (N_4643,N_3526,N_3965);
and U4644 (N_4644,N_3247,N_3011);
nand U4645 (N_4645,N_3863,N_3191);
and U4646 (N_4646,N_3643,N_3323);
nor U4647 (N_4647,N_3844,N_3453);
xnor U4648 (N_4648,N_3124,N_3823);
nand U4649 (N_4649,N_3193,N_3099);
and U4650 (N_4650,N_3877,N_3185);
nand U4651 (N_4651,N_3911,N_3645);
nand U4652 (N_4652,N_3080,N_3540);
xnor U4653 (N_4653,N_3736,N_3899);
and U4654 (N_4654,N_3143,N_3747);
or U4655 (N_4655,N_3342,N_3487);
xor U4656 (N_4656,N_3007,N_3581);
xor U4657 (N_4657,N_3716,N_3262);
nor U4658 (N_4658,N_3589,N_3703);
or U4659 (N_4659,N_3159,N_3344);
and U4660 (N_4660,N_3647,N_3593);
nor U4661 (N_4661,N_3143,N_3564);
nor U4662 (N_4662,N_3870,N_3087);
nor U4663 (N_4663,N_3996,N_3990);
or U4664 (N_4664,N_3757,N_3927);
xnor U4665 (N_4665,N_3159,N_3963);
nor U4666 (N_4666,N_3599,N_3066);
or U4667 (N_4667,N_3332,N_3124);
xor U4668 (N_4668,N_3588,N_3698);
nand U4669 (N_4669,N_3154,N_3345);
nand U4670 (N_4670,N_3579,N_3058);
nand U4671 (N_4671,N_3909,N_3620);
xor U4672 (N_4672,N_3684,N_3398);
nand U4673 (N_4673,N_3147,N_3593);
nand U4674 (N_4674,N_3077,N_3207);
nand U4675 (N_4675,N_3132,N_3900);
and U4676 (N_4676,N_3861,N_3878);
nor U4677 (N_4677,N_3556,N_3237);
or U4678 (N_4678,N_3924,N_3917);
nand U4679 (N_4679,N_3968,N_3508);
or U4680 (N_4680,N_3514,N_3067);
or U4681 (N_4681,N_3688,N_3740);
nand U4682 (N_4682,N_3026,N_3742);
nand U4683 (N_4683,N_3080,N_3264);
nor U4684 (N_4684,N_3650,N_3080);
or U4685 (N_4685,N_3937,N_3075);
and U4686 (N_4686,N_3696,N_3412);
nor U4687 (N_4687,N_3073,N_3460);
nor U4688 (N_4688,N_3184,N_3357);
or U4689 (N_4689,N_3470,N_3885);
or U4690 (N_4690,N_3254,N_3987);
xnor U4691 (N_4691,N_3682,N_3311);
or U4692 (N_4692,N_3810,N_3349);
and U4693 (N_4693,N_3390,N_3305);
xor U4694 (N_4694,N_3239,N_3341);
nor U4695 (N_4695,N_3537,N_3057);
xnor U4696 (N_4696,N_3281,N_3277);
nor U4697 (N_4697,N_3370,N_3138);
or U4698 (N_4698,N_3529,N_3083);
xnor U4699 (N_4699,N_3373,N_3177);
or U4700 (N_4700,N_3445,N_3748);
xor U4701 (N_4701,N_3390,N_3568);
xnor U4702 (N_4702,N_3277,N_3440);
and U4703 (N_4703,N_3371,N_3324);
xnor U4704 (N_4704,N_3416,N_3695);
nand U4705 (N_4705,N_3934,N_3112);
xnor U4706 (N_4706,N_3564,N_3305);
nor U4707 (N_4707,N_3891,N_3086);
xnor U4708 (N_4708,N_3956,N_3636);
nor U4709 (N_4709,N_3612,N_3326);
or U4710 (N_4710,N_3966,N_3525);
nor U4711 (N_4711,N_3237,N_3445);
nand U4712 (N_4712,N_3378,N_3586);
nor U4713 (N_4713,N_3126,N_3729);
nor U4714 (N_4714,N_3289,N_3972);
or U4715 (N_4715,N_3358,N_3252);
xnor U4716 (N_4716,N_3387,N_3605);
nor U4717 (N_4717,N_3510,N_3936);
nor U4718 (N_4718,N_3961,N_3752);
or U4719 (N_4719,N_3361,N_3577);
nor U4720 (N_4720,N_3206,N_3686);
xnor U4721 (N_4721,N_3654,N_3025);
xor U4722 (N_4722,N_3788,N_3602);
nor U4723 (N_4723,N_3022,N_3244);
nor U4724 (N_4724,N_3434,N_3664);
nor U4725 (N_4725,N_3006,N_3868);
nor U4726 (N_4726,N_3037,N_3466);
or U4727 (N_4727,N_3143,N_3714);
xor U4728 (N_4728,N_3514,N_3866);
and U4729 (N_4729,N_3662,N_3941);
nand U4730 (N_4730,N_3234,N_3576);
and U4731 (N_4731,N_3668,N_3741);
nor U4732 (N_4732,N_3954,N_3733);
and U4733 (N_4733,N_3142,N_3839);
or U4734 (N_4734,N_3161,N_3028);
and U4735 (N_4735,N_3805,N_3118);
nor U4736 (N_4736,N_3373,N_3740);
nand U4737 (N_4737,N_3909,N_3749);
nand U4738 (N_4738,N_3822,N_3041);
xnor U4739 (N_4739,N_3144,N_3860);
or U4740 (N_4740,N_3422,N_3068);
or U4741 (N_4741,N_3707,N_3397);
xnor U4742 (N_4742,N_3648,N_3229);
and U4743 (N_4743,N_3897,N_3010);
or U4744 (N_4744,N_3448,N_3646);
xor U4745 (N_4745,N_3799,N_3589);
or U4746 (N_4746,N_3982,N_3082);
nand U4747 (N_4747,N_3334,N_3516);
nor U4748 (N_4748,N_3420,N_3925);
or U4749 (N_4749,N_3942,N_3816);
or U4750 (N_4750,N_3316,N_3383);
nor U4751 (N_4751,N_3204,N_3250);
nand U4752 (N_4752,N_3073,N_3962);
xor U4753 (N_4753,N_3034,N_3147);
or U4754 (N_4754,N_3360,N_3647);
or U4755 (N_4755,N_3530,N_3025);
and U4756 (N_4756,N_3588,N_3185);
nand U4757 (N_4757,N_3462,N_3115);
and U4758 (N_4758,N_3979,N_3320);
and U4759 (N_4759,N_3133,N_3614);
nor U4760 (N_4760,N_3063,N_3211);
nand U4761 (N_4761,N_3157,N_3184);
nor U4762 (N_4762,N_3243,N_3798);
or U4763 (N_4763,N_3865,N_3411);
xor U4764 (N_4764,N_3436,N_3283);
or U4765 (N_4765,N_3425,N_3985);
and U4766 (N_4766,N_3374,N_3085);
nor U4767 (N_4767,N_3125,N_3091);
xor U4768 (N_4768,N_3867,N_3421);
xnor U4769 (N_4769,N_3551,N_3273);
or U4770 (N_4770,N_3207,N_3056);
and U4771 (N_4771,N_3733,N_3810);
nor U4772 (N_4772,N_3964,N_3147);
or U4773 (N_4773,N_3150,N_3126);
or U4774 (N_4774,N_3907,N_3707);
nand U4775 (N_4775,N_3958,N_3525);
xnor U4776 (N_4776,N_3073,N_3411);
or U4777 (N_4777,N_3068,N_3091);
xnor U4778 (N_4778,N_3308,N_3318);
xor U4779 (N_4779,N_3672,N_3052);
nand U4780 (N_4780,N_3680,N_3059);
or U4781 (N_4781,N_3768,N_3937);
nand U4782 (N_4782,N_3392,N_3913);
and U4783 (N_4783,N_3549,N_3992);
or U4784 (N_4784,N_3305,N_3090);
or U4785 (N_4785,N_3048,N_3080);
or U4786 (N_4786,N_3603,N_3541);
nand U4787 (N_4787,N_3858,N_3095);
xor U4788 (N_4788,N_3481,N_3455);
nand U4789 (N_4789,N_3105,N_3962);
and U4790 (N_4790,N_3379,N_3041);
and U4791 (N_4791,N_3623,N_3084);
xor U4792 (N_4792,N_3653,N_3164);
or U4793 (N_4793,N_3343,N_3067);
nor U4794 (N_4794,N_3565,N_3864);
nand U4795 (N_4795,N_3378,N_3093);
xor U4796 (N_4796,N_3533,N_3697);
xnor U4797 (N_4797,N_3482,N_3637);
or U4798 (N_4798,N_3159,N_3320);
nand U4799 (N_4799,N_3484,N_3690);
and U4800 (N_4800,N_3584,N_3618);
and U4801 (N_4801,N_3839,N_3384);
xnor U4802 (N_4802,N_3191,N_3103);
and U4803 (N_4803,N_3375,N_3783);
nand U4804 (N_4804,N_3012,N_3504);
nor U4805 (N_4805,N_3018,N_3279);
nor U4806 (N_4806,N_3002,N_3346);
or U4807 (N_4807,N_3765,N_3665);
xor U4808 (N_4808,N_3750,N_3807);
nand U4809 (N_4809,N_3340,N_3952);
and U4810 (N_4810,N_3938,N_3615);
nor U4811 (N_4811,N_3472,N_3178);
nand U4812 (N_4812,N_3458,N_3375);
and U4813 (N_4813,N_3472,N_3463);
nand U4814 (N_4814,N_3102,N_3638);
xnor U4815 (N_4815,N_3135,N_3985);
and U4816 (N_4816,N_3500,N_3134);
nor U4817 (N_4817,N_3210,N_3619);
nor U4818 (N_4818,N_3119,N_3146);
nor U4819 (N_4819,N_3719,N_3461);
and U4820 (N_4820,N_3847,N_3549);
nor U4821 (N_4821,N_3988,N_3284);
xor U4822 (N_4822,N_3999,N_3149);
or U4823 (N_4823,N_3164,N_3358);
xnor U4824 (N_4824,N_3004,N_3480);
and U4825 (N_4825,N_3045,N_3998);
xor U4826 (N_4826,N_3507,N_3097);
xnor U4827 (N_4827,N_3530,N_3043);
xnor U4828 (N_4828,N_3925,N_3959);
nor U4829 (N_4829,N_3459,N_3012);
xor U4830 (N_4830,N_3036,N_3188);
xnor U4831 (N_4831,N_3917,N_3106);
nor U4832 (N_4832,N_3385,N_3348);
nand U4833 (N_4833,N_3171,N_3927);
nand U4834 (N_4834,N_3295,N_3624);
and U4835 (N_4835,N_3092,N_3034);
xor U4836 (N_4836,N_3292,N_3941);
and U4837 (N_4837,N_3831,N_3471);
or U4838 (N_4838,N_3770,N_3860);
nand U4839 (N_4839,N_3624,N_3774);
nand U4840 (N_4840,N_3133,N_3306);
and U4841 (N_4841,N_3759,N_3665);
and U4842 (N_4842,N_3601,N_3538);
xnor U4843 (N_4843,N_3024,N_3677);
and U4844 (N_4844,N_3348,N_3134);
nor U4845 (N_4845,N_3944,N_3590);
nand U4846 (N_4846,N_3016,N_3337);
nor U4847 (N_4847,N_3328,N_3279);
xor U4848 (N_4848,N_3001,N_3104);
and U4849 (N_4849,N_3257,N_3659);
nor U4850 (N_4850,N_3557,N_3524);
or U4851 (N_4851,N_3789,N_3059);
nand U4852 (N_4852,N_3920,N_3717);
or U4853 (N_4853,N_3045,N_3060);
xor U4854 (N_4854,N_3819,N_3389);
nand U4855 (N_4855,N_3258,N_3815);
xor U4856 (N_4856,N_3548,N_3878);
nor U4857 (N_4857,N_3885,N_3335);
nor U4858 (N_4858,N_3335,N_3006);
nor U4859 (N_4859,N_3815,N_3868);
nor U4860 (N_4860,N_3288,N_3182);
nor U4861 (N_4861,N_3143,N_3079);
nand U4862 (N_4862,N_3967,N_3456);
nand U4863 (N_4863,N_3677,N_3428);
nor U4864 (N_4864,N_3916,N_3113);
and U4865 (N_4865,N_3551,N_3591);
or U4866 (N_4866,N_3322,N_3895);
or U4867 (N_4867,N_3615,N_3073);
xor U4868 (N_4868,N_3647,N_3923);
nand U4869 (N_4869,N_3457,N_3123);
nor U4870 (N_4870,N_3548,N_3798);
and U4871 (N_4871,N_3651,N_3626);
and U4872 (N_4872,N_3924,N_3041);
or U4873 (N_4873,N_3530,N_3552);
xnor U4874 (N_4874,N_3491,N_3832);
or U4875 (N_4875,N_3719,N_3761);
and U4876 (N_4876,N_3953,N_3898);
nor U4877 (N_4877,N_3163,N_3139);
xnor U4878 (N_4878,N_3091,N_3247);
and U4879 (N_4879,N_3032,N_3041);
xor U4880 (N_4880,N_3818,N_3554);
nor U4881 (N_4881,N_3646,N_3907);
nand U4882 (N_4882,N_3093,N_3025);
xnor U4883 (N_4883,N_3507,N_3420);
or U4884 (N_4884,N_3060,N_3946);
xor U4885 (N_4885,N_3769,N_3196);
xor U4886 (N_4886,N_3848,N_3511);
nor U4887 (N_4887,N_3339,N_3522);
or U4888 (N_4888,N_3988,N_3998);
nor U4889 (N_4889,N_3244,N_3053);
nand U4890 (N_4890,N_3919,N_3689);
nand U4891 (N_4891,N_3870,N_3741);
xnor U4892 (N_4892,N_3685,N_3321);
or U4893 (N_4893,N_3859,N_3330);
or U4894 (N_4894,N_3263,N_3342);
nand U4895 (N_4895,N_3208,N_3259);
and U4896 (N_4896,N_3013,N_3336);
nor U4897 (N_4897,N_3065,N_3442);
xnor U4898 (N_4898,N_3222,N_3708);
or U4899 (N_4899,N_3525,N_3073);
nand U4900 (N_4900,N_3549,N_3386);
nand U4901 (N_4901,N_3833,N_3869);
xor U4902 (N_4902,N_3418,N_3475);
or U4903 (N_4903,N_3109,N_3096);
nor U4904 (N_4904,N_3339,N_3776);
nand U4905 (N_4905,N_3682,N_3946);
xnor U4906 (N_4906,N_3228,N_3547);
xor U4907 (N_4907,N_3329,N_3216);
or U4908 (N_4908,N_3476,N_3052);
nor U4909 (N_4909,N_3880,N_3393);
nand U4910 (N_4910,N_3861,N_3548);
or U4911 (N_4911,N_3157,N_3659);
and U4912 (N_4912,N_3403,N_3569);
and U4913 (N_4913,N_3515,N_3330);
and U4914 (N_4914,N_3338,N_3515);
nand U4915 (N_4915,N_3089,N_3699);
and U4916 (N_4916,N_3975,N_3684);
xor U4917 (N_4917,N_3931,N_3322);
xnor U4918 (N_4918,N_3389,N_3860);
nor U4919 (N_4919,N_3061,N_3642);
nor U4920 (N_4920,N_3164,N_3953);
or U4921 (N_4921,N_3909,N_3743);
xor U4922 (N_4922,N_3000,N_3174);
nor U4923 (N_4923,N_3196,N_3480);
nor U4924 (N_4924,N_3279,N_3142);
nand U4925 (N_4925,N_3034,N_3677);
xor U4926 (N_4926,N_3560,N_3505);
and U4927 (N_4927,N_3006,N_3718);
or U4928 (N_4928,N_3482,N_3257);
nand U4929 (N_4929,N_3583,N_3366);
xor U4930 (N_4930,N_3638,N_3919);
xnor U4931 (N_4931,N_3204,N_3879);
or U4932 (N_4932,N_3442,N_3394);
nand U4933 (N_4933,N_3872,N_3728);
nor U4934 (N_4934,N_3969,N_3059);
nand U4935 (N_4935,N_3300,N_3714);
and U4936 (N_4936,N_3834,N_3948);
nor U4937 (N_4937,N_3457,N_3208);
nor U4938 (N_4938,N_3827,N_3219);
nor U4939 (N_4939,N_3231,N_3983);
and U4940 (N_4940,N_3287,N_3901);
and U4941 (N_4941,N_3142,N_3604);
and U4942 (N_4942,N_3085,N_3070);
nor U4943 (N_4943,N_3889,N_3579);
and U4944 (N_4944,N_3636,N_3961);
or U4945 (N_4945,N_3354,N_3446);
or U4946 (N_4946,N_3785,N_3084);
nand U4947 (N_4947,N_3693,N_3520);
nor U4948 (N_4948,N_3132,N_3827);
nand U4949 (N_4949,N_3926,N_3946);
or U4950 (N_4950,N_3883,N_3481);
or U4951 (N_4951,N_3216,N_3061);
xor U4952 (N_4952,N_3674,N_3295);
nor U4953 (N_4953,N_3407,N_3935);
and U4954 (N_4954,N_3320,N_3093);
xnor U4955 (N_4955,N_3119,N_3616);
nor U4956 (N_4956,N_3936,N_3726);
xor U4957 (N_4957,N_3087,N_3557);
nand U4958 (N_4958,N_3057,N_3968);
or U4959 (N_4959,N_3601,N_3018);
and U4960 (N_4960,N_3310,N_3703);
or U4961 (N_4961,N_3671,N_3939);
and U4962 (N_4962,N_3460,N_3266);
nor U4963 (N_4963,N_3079,N_3751);
xnor U4964 (N_4964,N_3651,N_3374);
or U4965 (N_4965,N_3866,N_3353);
nand U4966 (N_4966,N_3431,N_3248);
xnor U4967 (N_4967,N_3827,N_3446);
nand U4968 (N_4968,N_3281,N_3497);
nor U4969 (N_4969,N_3781,N_3536);
nor U4970 (N_4970,N_3298,N_3978);
xnor U4971 (N_4971,N_3862,N_3076);
or U4972 (N_4972,N_3758,N_3997);
nand U4973 (N_4973,N_3292,N_3090);
nor U4974 (N_4974,N_3532,N_3687);
nor U4975 (N_4975,N_3665,N_3094);
xnor U4976 (N_4976,N_3928,N_3168);
and U4977 (N_4977,N_3161,N_3394);
nor U4978 (N_4978,N_3085,N_3782);
or U4979 (N_4979,N_3401,N_3642);
or U4980 (N_4980,N_3285,N_3308);
nor U4981 (N_4981,N_3639,N_3801);
xnor U4982 (N_4982,N_3313,N_3478);
and U4983 (N_4983,N_3767,N_3904);
xor U4984 (N_4984,N_3121,N_3027);
or U4985 (N_4985,N_3434,N_3944);
nor U4986 (N_4986,N_3579,N_3169);
or U4987 (N_4987,N_3995,N_3216);
xor U4988 (N_4988,N_3522,N_3700);
and U4989 (N_4989,N_3037,N_3241);
nor U4990 (N_4990,N_3281,N_3819);
or U4991 (N_4991,N_3407,N_3371);
nor U4992 (N_4992,N_3216,N_3223);
nor U4993 (N_4993,N_3529,N_3236);
xor U4994 (N_4994,N_3411,N_3543);
nand U4995 (N_4995,N_3220,N_3158);
and U4996 (N_4996,N_3708,N_3532);
xor U4997 (N_4997,N_3848,N_3483);
and U4998 (N_4998,N_3280,N_3893);
and U4999 (N_4999,N_3200,N_3193);
xor UO_0 (O_0,N_4592,N_4653);
nand UO_1 (O_1,N_4510,N_4294);
nor UO_2 (O_2,N_4332,N_4953);
xor UO_3 (O_3,N_4360,N_4888);
nand UO_4 (O_4,N_4496,N_4193);
or UO_5 (O_5,N_4788,N_4630);
nand UO_6 (O_6,N_4388,N_4734);
nand UO_7 (O_7,N_4257,N_4752);
nor UO_8 (O_8,N_4603,N_4454);
or UO_9 (O_9,N_4112,N_4292);
nand UO_10 (O_10,N_4606,N_4965);
or UO_11 (O_11,N_4746,N_4990);
xor UO_12 (O_12,N_4167,N_4500);
nor UO_13 (O_13,N_4816,N_4088);
or UO_14 (O_14,N_4674,N_4456);
nor UO_15 (O_15,N_4955,N_4376);
or UO_16 (O_16,N_4906,N_4024);
nand UO_17 (O_17,N_4714,N_4331);
nor UO_18 (O_18,N_4980,N_4662);
and UO_19 (O_19,N_4511,N_4197);
nor UO_20 (O_20,N_4975,N_4179);
xnor UO_21 (O_21,N_4673,N_4609);
xnor UO_22 (O_22,N_4043,N_4684);
nor UO_23 (O_23,N_4896,N_4401);
xnor UO_24 (O_24,N_4512,N_4622);
and UO_25 (O_25,N_4080,N_4085);
nor UO_26 (O_26,N_4514,N_4260);
and UO_27 (O_27,N_4134,N_4803);
or UO_28 (O_28,N_4768,N_4950);
or UO_29 (O_29,N_4231,N_4423);
or UO_30 (O_30,N_4006,N_4730);
nor UO_31 (O_31,N_4474,N_4656);
nand UO_32 (O_32,N_4517,N_4051);
xnor UO_33 (O_33,N_4974,N_4163);
xnor UO_34 (O_34,N_4407,N_4537);
and UO_35 (O_35,N_4605,N_4543);
or UO_36 (O_36,N_4610,N_4305);
or UO_37 (O_37,N_4594,N_4560);
and UO_38 (O_38,N_4307,N_4201);
and UO_39 (O_39,N_4072,N_4859);
or UO_40 (O_40,N_4289,N_4922);
xor UO_41 (O_41,N_4410,N_4183);
and UO_42 (O_42,N_4831,N_4427);
nand UO_43 (O_43,N_4329,N_4569);
xnor UO_44 (O_44,N_4437,N_4604);
xnor UO_45 (O_45,N_4936,N_4524);
xnor UO_46 (O_46,N_4216,N_4009);
nand UO_47 (O_47,N_4719,N_4219);
or UO_48 (O_48,N_4189,N_4280);
nor UO_49 (O_49,N_4494,N_4618);
nand UO_50 (O_50,N_4599,N_4534);
or UO_51 (O_51,N_4177,N_4228);
nor UO_52 (O_52,N_4882,N_4481);
or UO_53 (O_53,N_4866,N_4453);
xnor UO_54 (O_54,N_4636,N_4647);
and UO_55 (O_55,N_4196,N_4880);
and UO_56 (O_56,N_4264,N_4834);
and UO_57 (O_57,N_4995,N_4272);
and UO_58 (O_58,N_4550,N_4504);
nor UO_59 (O_59,N_4891,N_4690);
or UO_60 (O_60,N_4760,N_4602);
nand UO_61 (O_61,N_4152,N_4860);
and UO_62 (O_62,N_4055,N_4931);
or UO_63 (O_63,N_4877,N_4519);
xnor UO_64 (O_64,N_4027,N_4379);
or UO_65 (O_65,N_4439,N_4070);
nand UO_66 (O_66,N_4142,N_4246);
and UO_67 (O_67,N_4467,N_4290);
nor UO_68 (O_68,N_4670,N_4149);
and UO_69 (O_69,N_4729,N_4977);
nand UO_70 (O_70,N_4659,N_4047);
xnor UO_71 (O_71,N_4374,N_4476);
xnor UO_72 (O_72,N_4062,N_4774);
xor UO_73 (O_73,N_4966,N_4230);
or UO_74 (O_74,N_4155,N_4804);
and UO_75 (O_75,N_4801,N_4205);
xnor UO_76 (O_76,N_4204,N_4683);
or UO_77 (O_77,N_4417,N_4358);
nor UO_78 (O_78,N_4191,N_4981);
and UO_79 (O_79,N_4276,N_4371);
or UO_80 (O_80,N_4827,N_4722);
nand UO_81 (O_81,N_4778,N_4991);
xor UO_82 (O_82,N_4472,N_4459);
nor UO_83 (O_83,N_4930,N_4796);
and UO_84 (O_84,N_4387,N_4902);
nand UO_85 (O_85,N_4020,N_4852);
xnor UO_86 (O_86,N_4172,N_4297);
nand UO_87 (O_87,N_4635,N_4114);
and UO_88 (O_88,N_4727,N_4074);
and UO_89 (O_89,N_4435,N_4222);
nand UO_90 (O_90,N_4352,N_4631);
or UO_91 (O_91,N_4279,N_4701);
nand UO_92 (O_92,N_4198,N_4584);
nand UO_93 (O_93,N_4909,N_4724);
nand UO_94 (O_94,N_4935,N_4354);
or UO_95 (O_95,N_4612,N_4215);
xnor UO_96 (O_96,N_4516,N_4098);
nor UO_97 (O_97,N_4252,N_4840);
nor UO_98 (O_98,N_4824,N_4706);
nor UO_99 (O_99,N_4864,N_4747);
or UO_100 (O_100,N_4182,N_4751);
nor UO_101 (O_101,N_4259,N_4220);
or UO_102 (O_102,N_4773,N_4806);
or UO_103 (O_103,N_4726,N_4994);
nor UO_104 (O_104,N_4870,N_4945);
xnor UO_105 (O_105,N_4551,N_4238);
or UO_106 (O_106,N_4836,N_4025);
nor UO_107 (O_107,N_4503,N_4132);
or UO_108 (O_108,N_4996,N_4739);
or UO_109 (O_109,N_4780,N_4643);
xnor UO_110 (O_110,N_4745,N_4758);
nand UO_111 (O_111,N_4213,N_4968);
nor UO_112 (O_112,N_4807,N_4601);
or UO_113 (O_113,N_4478,N_4446);
nor UO_114 (O_114,N_4320,N_4750);
and UO_115 (O_115,N_4185,N_4023);
nand UO_116 (O_116,N_4949,N_4367);
xnor UO_117 (O_117,N_4812,N_4066);
nand UO_118 (O_118,N_4110,N_4833);
and UO_119 (O_119,N_4444,N_4717);
nand UO_120 (O_120,N_4288,N_4666);
nor UO_121 (O_121,N_4287,N_4923);
or UO_122 (O_122,N_4792,N_4771);
xnor UO_123 (O_123,N_4638,N_4413);
or UO_124 (O_124,N_4992,N_4822);
or UO_125 (O_125,N_4588,N_4925);
xor UO_126 (O_126,N_4421,N_4430);
and UO_127 (O_127,N_4460,N_4939);
nor UO_128 (O_128,N_4957,N_4581);
nor UO_129 (O_129,N_4687,N_4267);
nand UO_130 (O_130,N_4572,N_4349);
nand UO_131 (O_131,N_4497,N_4203);
nor UO_132 (O_132,N_4251,N_4910);
nor UO_133 (O_133,N_4766,N_4558);
and UO_134 (O_134,N_4702,N_4124);
and UO_135 (O_135,N_4914,N_4723);
xnor UO_136 (O_136,N_4785,N_4502);
nor UO_137 (O_137,N_4060,N_4944);
nand UO_138 (O_138,N_4099,N_4044);
and UO_139 (O_139,N_4976,N_4141);
nor UO_140 (O_140,N_4339,N_4528);
or UO_141 (O_141,N_4972,N_4495);
nor UO_142 (O_142,N_4616,N_4056);
or UO_143 (O_143,N_4614,N_4715);
xor UO_144 (O_144,N_4372,N_4895);
nand UO_145 (O_145,N_4082,N_4590);
nor UO_146 (O_146,N_4698,N_4225);
and UO_147 (O_147,N_4591,N_4743);
nor UO_148 (O_148,N_4458,N_4987);
and UO_149 (O_149,N_4400,N_4022);
or UO_150 (O_150,N_4844,N_4736);
nor UO_151 (O_151,N_4383,N_4818);
nand UO_152 (O_152,N_4820,N_4837);
xnor UO_153 (O_153,N_4823,N_4414);
nor UO_154 (O_154,N_4641,N_4032);
and UO_155 (O_155,N_4583,N_4915);
and UO_156 (O_156,N_4657,N_4784);
nand UO_157 (O_157,N_4688,N_4946);
nand UO_158 (O_158,N_4933,N_4003);
xnor UO_159 (O_159,N_4171,N_4274);
nor UO_160 (O_160,N_4889,N_4962);
nand UO_161 (O_161,N_4317,N_4620);
and UO_162 (O_162,N_4180,N_4951);
xnor UO_163 (O_163,N_4471,N_4059);
or UO_164 (O_164,N_4057,N_4244);
nand UO_165 (O_165,N_4808,N_4542);
nand UO_166 (O_166,N_4874,N_4243);
and UO_167 (O_167,N_4529,N_4181);
nor UO_168 (O_168,N_4680,N_4640);
xor UO_169 (O_169,N_4553,N_4342);
and UO_170 (O_170,N_4559,N_4095);
xnor UO_171 (O_171,N_4391,N_4042);
nand UO_172 (O_172,N_4985,N_4999);
xor UO_173 (O_173,N_4079,N_4821);
and UO_174 (O_174,N_4862,N_4286);
nand UO_175 (O_175,N_4703,N_4782);
nor UO_176 (O_176,N_4691,N_4646);
or UO_177 (O_177,N_4767,N_4798);
nor UO_178 (O_178,N_4355,N_4685);
or UO_179 (O_179,N_4654,N_4819);
nor UO_180 (O_180,N_4749,N_4893);
nor UO_181 (O_181,N_4942,N_4166);
nand UO_182 (O_182,N_4802,N_4786);
and UO_183 (O_183,N_4119,N_4855);
nand UO_184 (O_184,N_4755,N_4316);
xor UO_185 (O_185,N_4664,N_4211);
or UO_186 (O_186,N_4757,N_4068);
xnor UO_187 (O_187,N_4932,N_4732);
xor UO_188 (O_188,N_4487,N_4593);
nand UO_189 (O_189,N_4483,N_4012);
and UO_190 (O_190,N_4411,N_4389);
nand UO_191 (O_191,N_4200,N_4111);
nand UO_192 (O_192,N_4711,N_4318);
nor UO_193 (O_193,N_4623,N_4904);
nand UO_194 (O_194,N_4829,N_4894);
and UO_195 (O_195,N_4035,N_4105);
xor UO_196 (O_196,N_4291,N_4261);
and UO_197 (O_197,N_4769,N_4629);
or UO_198 (O_198,N_4563,N_4348);
and UO_199 (O_199,N_4489,N_4164);
xor UO_200 (O_200,N_4544,N_4063);
nand UO_201 (O_201,N_4508,N_4113);
xor UO_202 (O_202,N_4426,N_4916);
nor UO_203 (O_203,N_4102,N_4578);
and UO_204 (O_204,N_4109,N_4469);
and UO_205 (O_205,N_4740,N_4682);
or UO_206 (O_206,N_4327,N_4394);
nor UO_207 (O_207,N_4312,N_4507);
nor UO_208 (O_208,N_4983,N_4839);
nand UO_209 (O_209,N_4465,N_4323);
nand UO_210 (O_210,N_4143,N_4952);
and UO_211 (O_211,N_4709,N_4589);
nand UO_212 (O_212,N_4160,N_4648);
nor UO_213 (O_213,N_4908,N_4315);
xor UO_214 (O_214,N_4223,N_4368);
xnor UO_215 (O_215,N_4301,N_4013);
nor UO_216 (O_216,N_4262,N_4628);
nor UO_217 (O_217,N_4525,N_4169);
and UO_218 (O_218,N_4665,N_4378);
and UO_219 (O_219,N_4096,N_4236);
xnor UO_220 (O_220,N_4370,N_4303);
xnor UO_221 (O_221,N_4997,N_4775);
and UO_222 (O_222,N_4790,N_4725);
and UO_223 (O_223,N_4577,N_4308);
or UO_224 (O_224,N_4486,N_4029);
nand UO_225 (O_225,N_4548,N_4359);
nor UO_226 (O_226,N_4979,N_4284);
or UO_227 (O_227,N_4395,N_4364);
or UO_228 (O_228,N_4135,N_4067);
or UO_229 (O_229,N_4644,N_4853);
or UO_230 (O_230,N_4536,N_4233);
or UO_231 (O_231,N_4737,N_4676);
nor UO_232 (O_232,N_4106,N_4744);
nand UO_233 (O_233,N_4552,N_4720);
or UO_234 (O_234,N_4281,N_4718);
nand UO_235 (O_235,N_4772,N_4187);
nand UO_236 (O_236,N_4344,N_4127);
nor UO_237 (O_237,N_4340,N_4422);
or UO_238 (O_238,N_4762,N_4137);
nand UO_239 (O_239,N_4741,N_4712);
and UO_240 (O_240,N_4770,N_4879);
nand UO_241 (O_241,N_4186,N_4002);
xnor UO_242 (O_242,N_4438,N_4325);
xor UO_243 (O_243,N_4271,N_4199);
nand UO_244 (O_244,N_4168,N_4101);
nand UO_245 (O_245,N_4832,N_4268);
nor UO_246 (O_246,N_4457,N_4861);
nor UO_247 (O_247,N_4011,N_4522);
nor UO_248 (O_248,N_4753,N_4018);
and UO_249 (O_249,N_4026,N_4139);
or UO_250 (O_250,N_4607,N_4429);
and UO_251 (O_251,N_4091,N_4580);
nand UO_252 (O_252,N_4296,N_4781);
and UO_253 (O_253,N_4016,N_4689);
xor UO_254 (O_254,N_4385,N_4667);
xnor UO_255 (O_255,N_4224,N_4302);
nor UO_256 (O_256,N_4254,N_4655);
nand UO_257 (O_257,N_4380,N_4412);
or UO_258 (O_258,N_4993,N_4961);
and UO_259 (O_259,N_4535,N_4652);
or UO_260 (O_260,N_4505,N_4566);
nor UO_261 (O_261,N_4131,N_4697);
or UO_262 (O_262,N_4540,N_4948);
nand UO_263 (O_263,N_4897,N_4695);
nand UO_264 (O_264,N_4565,N_4420);
or UO_265 (O_265,N_4324,N_4087);
nand UO_266 (O_266,N_4779,N_4392);
nor UO_267 (O_267,N_4595,N_4813);
xnor UO_268 (O_268,N_4428,N_4892);
and UO_269 (O_269,N_4868,N_4998);
nand UO_270 (O_270,N_4313,N_4576);
nand UO_271 (O_271,N_4184,N_4473);
xor UO_272 (O_272,N_4436,N_4463);
nand UO_273 (O_273,N_4396,N_4869);
nor UO_274 (O_274,N_4513,N_4165);
xnor UO_275 (O_275,N_4937,N_4278);
and UO_276 (O_276,N_4447,N_4140);
nor UO_277 (O_277,N_4207,N_4075);
xor UO_278 (O_278,N_4579,N_4479);
or UO_279 (O_279,N_4466,N_4034);
nand UO_280 (O_280,N_4694,N_4545);
or UO_281 (O_281,N_4617,N_4398);
or UO_282 (O_282,N_4899,N_4731);
nor UO_283 (O_283,N_4245,N_4570);
nand UO_284 (O_284,N_4651,N_4943);
and UO_285 (O_285,N_4761,N_4600);
xnor UO_286 (O_286,N_4624,N_4843);
or UO_287 (O_287,N_4763,N_4174);
and UO_288 (O_288,N_4582,N_4250);
and UO_289 (O_289,N_4488,N_4547);
nor UO_290 (O_290,N_4309,N_4619);
xnor UO_291 (O_291,N_4650,N_4482);
nor UO_292 (O_292,N_4273,N_4206);
or UO_293 (O_293,N_4954,N_4492);
nand UO_294 (O_294,N_4875,N_4815);
and UO_295 (O_295,N_4065,N_4735);
nor UO_296 (O_296,N_4842,N_4856);
nor UO_297 (O_297,N_4728,N_4121);
nand UO_298 (O_298,N_4585,N_4887);
or UO_299 (O_299,N_4156,N_4865);
or UO_300 (O_300,N_4293,N_4061);
nand UO_301 (O_301,N_4351,N_4863);
nor UO_302 (O_302,N_4014,N_4054);
nand UO_303 (O_303,N_4402,N_4940);
nor UO_304 (O_304,N_4133,N_4108);
and UO_305 (O_305,N_4001,N_4345);
xnor UO_306 (O_306,N_4337,N_4800);
nor UO_307 (O_307,N_4506,N_4649);
xnor UO_308 (O_308,N_4120,N_4128);
xor UO_309 (O_309,N_4967,N_4326);
nand UO_310 (O_310,N_4192,N_4586);
nor UO_311 (O_311,N_4443,N_4625);
and UO_312 (O_312,N_4848,N_4509);
xnor UO_313 (O_313,N_4615,N_4369);
nand UO_314 (O_314,N_4554,N_4058);
or UO_315 (O_315,N_4239,N_4092);
and UO_316 (O_316,N_4037,N_4425);
or UO_317 (O_317,N_4217,N_4677);
xor UO_318 (O_318,N_4632,N_4408);
xor UO_319 (O_319,N_4162,N_4658);
nand UO_320 (O_320,N_4721,N_4464);
or UO_321 (O_321,N_4626,N_4237);
nand UO_322 (O_322,N_4964,N_4538);
or UO_323 (O_323,N_4248,N_4485);
and UO_324 (O_324,N_4365,N_4776);
nand UO_325 (O_325,N_4050,N_4161);
or UO_326 (O_326,N_4136,N_4300);
nor UO_327 (O_327,N_4270,N_4053);
or UO_328 (O_328,N_4826,N_4283);
or UO_329 (O_329,N_4357,N_4052);
xor UO_330 (O_330,N_4253,N_4696);
or UO_331 (O_331,N_4692,N_4825);
nor UO_332 (O_332,N_4247,N_4126);
and UO_333 (O_333,N_4947,N_4461);
nand UO_334 (O_334,N_4007,N_4963);
nor UO_335 (O_335,N_4918,N_4518);
nand UO_336 (O_336,N_4448,N_4138);
nand UO_337 (O_337,N_4613,N_4188);
and UO_338 (O_338,N_4299,N_4275);
xnor UO_339 (O_339,N_4639,N_4406);
or UO_340 (O_340,N_4989,N_4107);
nor UO_341 (O_341,N_4266,N_4970);
nor UO_342 (O_342,N_4830,N_4708);
and UO_343 (O_343,N_4671,N_4285);
nand UO_344 (O_344,N_4710,N_4078);
or UO_345 (O_345,N_4175,N_4934);
nand UO_346 (O_346,N_4928,N_4145);
or UO_347 (O_347,N_4218,N_4828);
nand UO_348 (O_348,N_4153,N_4019);
xor UO_349 (O_349,N_4546,N_4100);
nor UO_350 (O_350,N_4575,N_4384);
or UO_351 (O_351,N_4382,N_4346);
nor UO_352 (O_352,N_4450,N_4221);
or UO_353 (O_353,N_4147,N_4883);
nor UO_354 (O_354,N_4347,N_4873);
and UO_355 (O_355,N_4424,N_4885);
and UO_356 (O_356,N_4797,N_4634);
and UO_357 (O_357,N_4386,N_4452);
or UO_358 (O_358,N_4841,N_4125);
nor UO_359 (O_359,N_4811,N_4549);
or UO_360 (O_360,N_4679,N_4898);
or UO_361 (O_361,N_4433,N_4971);
nor UO_362 (O_362,N_4491,N_4097);
nand UO_363 (O_363,N_4700,N_4415);
xor UO_364 (O_364,N_4036,N_4912);
nand UO_365 (O_365,N_4048,N_4645);
nor UO_366 (O_366,N_4960,N_4442);
or UO_367 (O_367,N_4116,N_4986);
nand UO_368 (O_368,N_4190,N_4334);
or UO_369 (O_369,N_4038,N_4094);
nor UO_370 (O_370,N_4462,N_4817);
xnor UO_371 (O_371,N_4490,N_4501);
nand UO_372 (O_372,N_4556,N_4319);
xor UO_373 (O_373,N_4969,N_4567);
nor UO_374 (O_374,N_4350,N_4277);
and UO_375 (O_375,N_4765,N_4269);
and UO_376 (O_376,N_4255,N_4907);
or UO_377 (O_377,N_4377,N_4212);
xnor UO_378 (O_378,N_4678,N_4927);
nand UO_379 (O_379,N_4982,N_4039);
nand UO_380 (O_380,N_4333,N_4077);
nor UO_381 (O_381,N_4046,N_4498);
xor UO_382 (O_382,N_4903,N_4045);
nor UO_383 (O_383,N_4104,N_4115);
nor UO_384 (O_384,N_4526,N_4202);
xor UO_385 (O_385,N_4304,N_4532);
nand UO_386 (O_386,N_4335,N_4851);
xnor UO_387 (O_387,N_4445,N_4157);
nor UO_388 (O_388,N_4089,N_4004);
nand UO_389 (O_389,N_4929,N_4226);
xor UO_390 (O_390,N_4809,N_4693);
or UO_391 (O_391,N_4361,N_4672);
xor UO_392 (O_392,N_4049,N_4028);
xor UO_393 (O_393,N_4884,N_4170);
nand UO_394 (O_394,N_4733,N_4030);
or UO_395 (O_395,N_4926,N_4093);
or UO_396 (O_396,N_4633,N_4878);
nor UO_397 (O_397,N_4010,N_4924);
xnor UO_398 (O_398,N_4176,N_4681);
nor UO_399 (O_399,N_4799,N_4314);
or UO_400 (O_400,N_4064,N_4984);
or UO_401 (O_401,N_4521,N_4081);
and UO_402 (O_402,N_4938,N_4660);
nand UO_403 (O_403,N_4675,N_4144);
or UO_404 (O_404,N_4330,N_4210);
and UO_405 (O_405,N_4084,N_4341);
nand UO_406 (O_406,N_4791,N_4431);
xnor UO_407 (O_407,N_4338,N_4838);
nand UO_408 (O_408,N_4040,N_4794);
or UO_409 (O_409,N_4130,N_4403);
nor UO_410 (O_410,N_4493,N_4759);
nand UO_411 (O_411,N_4470,N_4611);
and UO_412 (O_412,N_4310,N_4748);
nand UO_413 (O_413,N_4911,N_4699);
and UO_414 (O_414,N_4008,N_4397);
nor UO_415 (O_415,N_4103,N_4195);
nor UO_416 (O_416,N_4441,N_4520);
and UO_417 (O_417,N_4857,N_4561);
nor UO_418 (O_418,N_4241,N_4416);
and UO_419 (O_419,N_4956,N_4587);
xnor UO_420 (O_420,N_4076,N_4738);
xor UO_421 (O_421,N_4322,N_4083);
nor UO_422 (O_422,N_4480,N_4835);
and UO_423 (O_423,N_4871,N_4178);
nor UO_424 (O_424,N_4890,N_4901);
and UO_425 (O_425,N_4298,N_4704);
xor UO_426 (O_426,N_4455,N_4913);
and UO_427 (O_427,N_4867,N_4214);
xor UO_428 (O_428,N_4573,N_4959);
or UO_429 (O_429,N_4263,N_4146);
xor UO_430 (O_430,N_4336,N_4854);
xnor UO_431 (O_431,N_4475,N_4846);
xor UO_432 (O_432,N_4432,N_4571);
xor UO_433 (O_433,N_4086,N_4713);
nor UO_434 (O_434,N_4021,N_4539);
and UO_435 (O_435,N_4258,N_4265);
xor UO_436 (O_436,N_4921,N_4282);
nand UO_437 (O_437,N_4235,N_4158);
xnor UO_438 (O_438,N_4663,N_4596);
xor UO_439 (O_439,N_4117,N_4232);
nor UO_440 (O_440,N_4366,N_4850);
xnor UO_441 (O_441,N_4686,N_4849);
or UO_442 (O_442,N_4716,N_4742);
and UO_443 (O_443,N_4256,N_4564);
nor UO_444 (O_444,N_4754,N_4876);
nand UO_445 (O_445,N_4194,N_4306);
nand UO_446 (O_446,N_4249,N_4661);
and UO_447 (O_447,N_4390,N_4608);
or UO_448 (O_448,N_4642,N_4440);
xnor UO_449 (O_449,N_4150,N_4527);
nand UO_450 (O_450,N_4523,N_4154);
nand UO_451 (O_451,N_4705,N_4033);
and UO_452 (O_452,N_4707,N_4515);
or UO_453 (O_453,N_4451,N_4353);
nand UO_454 (O_454,N_4847,N_4404);
and UO_455 (O_455,N_4533,N_4783);
xnor UO_456 (O_456,N_4941,N_4555);
nor UO_457 (O_457,N_4311,N_4845);
xor UO_458 (O_458,N_4668,N_4363);
or UO_459 (O_459,N_4499,N_4574);
and UO_460 (O_460,N_4041,N_4234);
nor UO_461 (O_461,N_4793,N_4118);
or UO_462 (O_462,N_4777,N_4920);
xnor UO_463 (O_463,N_4405,N_4343);
nand UO_464 (O_464,N_4399,N_4484);
xnor UO_465 (O_465,N_4795,N_4393);
nand UO_466 (O_466,N_4409,N_4129);
xnor UO_467 (O_467,N_4227,N_4858);
xnor UO_468 (O_468,N_4814,N_4148);
nor UO_469 (O_469,N_4637,N_4373);
and UO_470 (O_470,N_4240,N_4090);
and UO_471 (O_471,N_4419,N_4789);
nor UO_472 (O_472,N_4621,N_4900);
and UO_473 (O_473,N_4434,N_4886);
nand UO_474 (O_474,N_4764,N_4151);
nand UO_475 (O_475,N_4017,N_4031);
nand UO_476 (O_476,N_4669,N_4597);
xor UO_477 (O_477,N_4756,N_4562);
nand UO_478 (O_478,N_4598,N_4375);
or UO_479 (O_479,N_4362,N_4905);
nor UO_480 (O_480,N_4787,N_4627);
nor UO_481 (O_481,N_4541,N_4000);
nand UO_482 (O_482,N_4978,N_4069);
and UO_483 (O_483,N_4530,N_4122);
nor UO_484 (O_484,N_4988,N_4973);
and UO_485 (O_485,N_4881,N_4005);
and UO_486 (O_486,N_4557,N_4159);
nor UO_487 (O_487,N_4242,N_4328);
and UO_488 (O_488,N_4468,N_4173);
xnor UO_489 (O_489,N_4418,N_4805);
and UO_490 (O_490,N_4295,N_4568);
xor UO_491 (O_491,N_4015,N_4958);
and UO_492 (O_492,N_4356,N_4919);
or UO_493 (O_493,N_4208,N_4321);
or UO_494 (O_494,N_4381,N_4449);
xor UO_495 (O_495,N_4209,N_4071);
nor UO_496 (O_496,N_4123,N_4917);
and UO_497 (O_497,N_4531,N_4073);
xor UO_498 (O_498,N_4477,N_4872);
nand UO_499 (O_499,N_4229,N_4810);
nor UO_500 (O_500,N_4586,N_4255);
nor UO_501 (O_501,N_4667,N_4007);
nand UO_502 (O_502,N_4289,N_4364);
nand UO_503 (O_503,N_4967,N_4862);
or UO_504 (O_504,N_4383,N_4837);
nand UO_505 (O_505,N_4843,N_4379);
nor UO_506 (O_506,N_4585,N_4641);
nand UO_507 (O_507,N_4610,N_4916);
nor UO_508 (O_508,N_4625,N_4222);
nor UO_509 (O_509,N_4137,N_4554);
nand UO_510 (O_510,N_4619,N_4751);
and UO_511 (O_511,N_4646,N_4210);
and UO_512 (O_512,N_4559,N_4778);
xor UO_513 (O_513,N_4240,N_4376);
nand UO_514 (O_514,N_4774,N_4964);
nor UO_515 (O_515,N_4960,N_4107);
and UO_516 (O_516,N_4100,N_4792);
or UO_517 (O_517,N_4348,N_4534);
nand UO_518 (O_518,N_4475,N_4042);
or UO_519 (O_519,N_4343,N_4793);
nand UO_520 (O_520,N_4150,N_4567);
and UO_521 (O_521,N_4986,N_4298);
and UO_522 (O_522,N_4926,N_4366);
and UO_523 (O_523,N_4993,N_4233);
nor UO_524 (O_524,N_4069,N_4125);
and UO_525 (O_525,N_4117,N_4274);
nor UO_526 (O_526,N_4365,N_4207);
nand UO_527 (O_527,N_4850,N_4005);
nand UO_528 (O_528,N_4295,N_4586);
and UO_529 (O_529,N_4879,N_4345);
nor UO_530 (O_530,N_4635,N_4666);
and UO_531 (O_531,N_4147,N_4284);
and UO_532 (O_532,N_4195,N_4812);
nor UO_533 (O_533,N_4459,N_4057);
and UO_534 (O_534,N_4629,N_4984);
nand UO_535 (O_535,N_4078,N_4647);
or UO_536 (O_536,N_4408,N_4424);
xnor UO_537 (O_537,N_4931,N_4033);
and UO_538 (O_538,N_4840,N_4163);
or UO_539 (O_539,N_4771,N_4628);
or UO_540 (O_540,N_4259,N_4604);
nor UO_541 (O_541,N_4741,N_4696);
nor UO_542 (O_542,N_4620,N_4741);
nor UO_543 (O_543,N_4392,N_4913);
xor UO_544 (O_544,N_4716,N_4453);
xnor UO_545 (O_545,N_4440,N_4645);
nand UO_546 (O_546,N_4068,N_4286);
or UO_547 (O_547,N_4568,N_4723);
xor UO_548 (O_548,N_4666,N_4200);
xnor UO_549 (O_549,N_4568,N_4454);
nand UO_550 (O_550,N_4964,N_4837);
nor UO_551 (O_551,N_4007,N_4198);
nand UO_552 (O_552,N_4567,N_4817);
nor UO_553 (O_553,N_4719,N_4726);
and UO_554 (O_554,N_4487,N_4154);
or UO_555 (O_555,N_4268,N_4641);
nand UO_556 (O_556,N_4410,N_4131);
nor UO_557 (O_557,N_4100,N_4204);
xnor UO_558 (O_558,N_4726,N_4592);
or UO_559 (O_559,N_4430,N_4186);
xnor UO_560 (O_560,N_4611,N_4465);
nand UO_561 (O_561,N_4274,N_4682);
and UO_562 (O_562,N_4573,N_4792);
nor UO_563 (O_563,N_4690,N_4948);
and UO_564 (O_564,N_4970,N_4090);
or UO_565 (O_565,N_4456,N_4320);
and UO_566 (O_566,N_4104,N_4863);
nor UO_567 (O_567,N_4577,N_4230);
nand UO_568 (O_568,N_4921,N_4647);
nor UO_569 (O_569,N_4443,N_4062);
and UO_570 (O_570,N_4930,N_4087);
and UO_571 (O_571,N_4485,N_4869);
and UO_572 (O_572,N_4221,N_4963);
and UO_573 (O_573,N_4093,N_4490);
xor UO_574 (O_574,N_4437,N_4385);
and UO_575 (O_575,N_4766,N_4394);
and UO_576 (O_576,N_4798,N_4308);
xnor UO_577 (O_577,N_4443,N_4720);
or UO_578 (O_578,N_4095,N_4514);
or UO_579 (O_579,N_4686,N_4044);
xnor UO_580 (O_580,N_4923,N_4700);
nor UO_581 (O_581,N_4756,N_4495);
nor UO_582 (O_582,N_4606,N_4705);
nand UO_583 (O_583,N_4538,N_4164);
xor UO_584 (O_584,N_4774,N_4235);
xnor UO_585 (O_585,N_4504,N_4884);
or UO_586 (O_586,N_4338,N_4689);
nand UO_587 (O_587,N_4318,N_4639);
nor UO_588 (O_588,N_4164,N_4153);
xor UO_589 (O_589,N_4156,N_4475);
or UO_590 (O_590,N_4623,N_4998);
or UO_591 (O_591,N_4523,N_4483);
and UO_592 (O_592,N_4556,N_4760);
nand UO_593 (O_593,N_4340,N_4695);
xor UO_594 (O_594,N_4715,N_4661);
xor UO_595 (O_595,N_4980,N_4866);
nor UO_596 (O_596,N_4202,N_4164);
and UO_597 (O_597,N_4522,N_4420);
nor UO_598 (O_598,N_4770,N_4398);
xnor UO_599 (O_599,N_4266,N_4167);
and UO_600 (O_600,N_4028,N_4740);
nand UO_601 (O_601,N_4548,N_4778);
and UO_602 (O_602,N_4684,N_4865);
and UO_603 (O_603,N_4352,N_4861);
nor UO_604 (O_604,N_4134,N_4339);
nand UO_605 (O_605,N_4255,N_4503);
nor UO_606 (O_606,N_4557,N_4274);
nor UO_607 (O_607,N_4089,N_4565);
or UO_608 (O_608,N_4600,N_4823);
and UO_609 (O_609,N_4007,N_4577);
and UO_610 (O_610,N_4520,N_4765);
xor UO_611 (O_611,N_4872,N_4022);
nand UO_612 (O_612,N_4365,N_4351);
nor UO_613 (O_613,N_4225,N_4562);
or UO_614 (O_614,N_4681,N_4931);
xnor UO_615 (O_615,N_4596,N_4084);
and UO_616 (O_616,N_4313,N_4560);
and UO_617 (O_617,N_4054,N_4586);
nand UO_618 (O_618,N_4646,N_4433);
nor UO_619 (O_619,N_4170,N_4499);
and UO_620 (O_620,N_4215,N_4448);
nand UO_621 (O_621,N_4455,N_4003);
nand UO_622 (O_622,N_4469,N_4215);
and UO_623 (O_623,N_4729,N_4473);
and UO_624 (O_624,N_4933,N_4675);
nor UO_625 (O_625,N_4962,N_4597);
and UO_626 (O_626,N_4677,N_4024);
nor UO_627 (O_627,N_4290,N_4088);
or UO_628 (O_628,N_4107,N_4906);
and UO_629 (O_629,N_4759,N_4933);
nor UO_630 (O_630,N_4230,N_4825);
xor UO_631 (O_631,N_4256,N_4710);
nor UO_632 (O_632,N_4308,N_4007);
nor UO_633 (O_633,N_4550,N_4671);
xor UO_634 (O_634,N_4742,N_4132);
xnor UO_635 (O_635,N_4235,N_4506);
xnor UO_636 (O_636,N_4729,N_4113);
nand UO_637 (O_637,N_4962,N_4370);
or UO_638 (O_638,N_4064,N_4259);
nand UO_639 (O_639,N_4085,N_4942);
and UO_640 (O_640,N_4549,N_4260);
or UO_641 (O_641,N_4607,N_4913);
or UO_642 (O_642,N_4501,N_4554);
or UO_643 (O_643,N_4593,N_4665);
and UO_644 (O_644,N_4693,N_4893);
nand UO_645 (O_645,N_4225,N_4003);
nor UO_646 (O_646,N_4590,N_4309);
nand UO_647 (O_647,N_4820,N_4041);
nand UO_648 (O_648,N_4415,N_4497);
xnor UO_649 (O_649,N_4505,N_4090);
and UO_650 (O_650,N_4250,N_4050);
and UO_651 (O_651,N_4779,N_4369);
nand UO_652 (O_652,N_4939,N_4809);
nand UO_653 (O_653,N_4896,N_4258);
nand UO_654 (O_654,N_4607,N_4923);
and UO_655 (O_655,N_4078,N_4985);
nand UO_656 (O_656,N_4995,N_4278);
or UO_657 (O_657,N_4588,N_4692);
xnor UO_658 (O_658,N_4208,N_4488);
and UO_659 (O_659,N_4400,N_4263);
xnor UO_660 (O_660,N_4295,N_4632);
and UO_661 (O_661,N_4714,N_4610);
nor UO_662 (O_662,N_4323,N_4760);
xnor UO_663 (O_663,N_4603,N_4305);
nand UO_664 (O_664,N_4262,N_4692);
and UO_665 (O_665,N_4114,N_4002);
nor UO_666 (O_666,N_4322,N_4197);
or UO_667 (O_667,N_4853,N_4403);
and UO_668 (O_668,N_4990,N_4367);
nor UO_669 (O_669,N_4310,N_4664);
or UO_670 (O_670,N_4156,N_4835);
nor UO_671 (O_671,N_4984,N_4096);
nor UO_672 (O_672,N_4405,N_4857);
and UO_673 (O_673,N_4600,N_4868);
xnor UO_674 (O_674,N_4831,N_4869);
nor UO_675 (O_675,N_4495,N_4907);
nand UO_676 (O_676,N_4845,N_4576);
or UO_677 (O_677,N_4302,N_4072);
and UO_678 (O_678,N_4202,N_4567);
nor UO_679 (O_679,N_4869,N_4281);
or UO_680 (O_680,N_4969,N_4617);
xnor UO_681 (O_681,N_4321,N_4026);
and UO_682 (O_682,N_4771,N_4761);
xnor UO_683 (O_683,N_4319,N_4821);
nor UO_684 (O_684,N_4497,N_4889);
and UO_685 (O_685,N_4757,N_4570);
and UO_686 (O_686,N_4912,N_4679);
or UO_687 (O_687,N_4041,N_4447);
nand UO_688 (O_688,N_4878,N_4837);
or UO_689 (O_689,N_4393,N_4279);
nor UO_690 (O_690,N_4137,N_4371);
nor UO_691 (O_691,N_4446,N_4202);
or UO_692 (O_692,N_4482,N_4941);
nand UO_693 (O_693,N_4191,N_4834);
or UO_694 (O_694,N_4493,N_4816);
or UO_695 (O_695,N_4657,N_4839);
and UO_696 (O_696,N_4057,N_4684);
nand UO_697 (O_697,N_4070,N_4601);
nand UO_698 (O_698,N_4584,N_4128);
nand UO_699 (O_699,N_4032,N_4257);
xor UO_700 (O_700,N_4044,N_4815);
and UO_701 (O_701,N_4042,N_4827);
xnor UO_702 (O_702,N_4469,N_4075);
nor UO_703 (O_703,N_4763,N_4244);
nor UO_704 (O_704,N_4424,N_4731);
nor UO_705 (O_705,N_4409,N_4018);
or UO_706 (O_706,N_4637,N_4655);
nor UO_707 (O_707,N_4408,N_4820);
or UO_708 (O_708,N_4482,N_4943);
or UO_709 (O_709,N_4934,N_4578);
nor UO_710 (O_710,N_4914,N_4298);
nor UO_711 (O_711,N_4038,N_4211);
nor UO_712 (O_712,N_4035,N_4181);
xnor UO_713 (O_713,N_4930,N_4478);
nand UO_714 (O_714,N_4866,N_4571);
xor UO_715 (O_715,N_4669,N_4714);
or UO_716 (O_716,N_4521,N_4139);
xor UO_717 (O_717,N_4771,N_4586);
or UO_718 (O_718,N_4608,N_4386);
or UO_719 (O_719,N_4053,N_4328);
and UO_720 (O_720,N_4944,N_4343);
nand UO_721 (O_721,N_4588,N_4385);
and UO_722 (O_722,N_4607,N_4080);
nand UO_723 (O_723,N_4630,N_4653);
nand UO_724 (O_724,N_4787,N_4335);
nor UO_725 (O_725,N_4589,N_4453);
nor UO_726 (O_726,N_4654,N_4941);
or UO_727 (O_727,N_4013,N_4404);
xnor UO_728 (O_728,N_4966,N_4146);
nand UO_729 (O_729,N_4694,N_4410);
xor UO_730 (O_730,N_4247,N_4111);
or UO_731 (O_731,N_4102,N_4949);
xor UO_732 (O_732,N_4262,N_4171);
nand UO_733 (O_733,N_4069,N_4533);
nor UO_734 (O_734,N_4791,N_4507);
or UO_735 (O_735,N_4305,N_4580);
nor UO_736 (O_736,N_4112,N_4103);
or UO_737 (O_737,N_4332,N_4210);
nand UO_738 (O_738,N_4519,N_4061);
nand UO_739 (O_739,N_4160,N_4292);
nor UO_740 (O_740,N_4184,N_4862);
or UO_741 (O_741,N_4836,N_4411);
nor UO_742 (O_742,N_4757,N_4226);
or UO_743 (O_743,N_4509,N_4652);
nand UO_744 (O_744,N_4192,N_4338);
nor UO_745 (O_745,N_4270,N_4152);
nor UO_746 (O_746,N_4224,N_4033);
xor UO_747 (O_747,N_4566,N_4562);
xor UO_748 (O_748,N_4087,N_4111);
nand UO_749 (O_749,N_4547,N_4706);
nor UO_750 (O_750,N_4799,N_4536);
and UO_751 (O_751,N_4467,N_4178);
or UO_752 (O_752,N_4373,N_4873);
nor UO_753 (O_753,N_4979,N_4167);
and UO_754 (O_754,N_4006,N_4038);
nor UO_755 (O_755,N_4133,N_4164);
xnor UO_756 (O_756,N_4695,N_4764);
nand UO_757 (O_757,N_4866,N_4065);
or UO_758 (O_758,N_4713,N_4488);
xnor UO_759 (O_759,N_4848,N_4006);
xnor UO_760 (O_760,N_4903,N_4719);
or UO_761 (O_761,N_4921,N_4439);
xor UO_762 (O_762,N_4030,N_4226);
or UO_763 (O_763,N_4275,N_4015);
nor UO_764 (O_764,N_4381,N_4781);
nor UO_765 (O_765,N_4998,N_4990);
nand UO_766 (O_766,N_4286,N_4563);
xnor UO_767 (O_767,N_4149,N_4855);
xnor UO_768 (O_768,N_4637,N_4235);
nor UO_769 (O_769,N_4771,N_4454);
and UO_770 (O_770,N_4770,N_4602);
xnor UO_771 (O_771,N_4449,N_4737);
xor UO_772 (O_772,N_4109,N_4815);
nand UO_773 (O_773,N_4348,N_4193);
nand UO_774 (O_774,N_4922,N_4697);
and UO_775 (O_775,N_4952,N_4130);
and UO_776 (O_776,N_4919,N_4304);
xnor UO_777 (O_777,N_4588,N_4034);
nand UO_778 (O_778,N_4179,N_4620);
nor UO_779 (O_779,N_4951,N_4796);
nand UO_780 (O_780,N_4671,N_4660);
xor UO_781 (O_781,N_4403,N_4160);
nor UO_782 (O_782,N_4965,N_4157);
and UO_783 (O_783,N_4368,N_4137);
or UO_784 (O_784,N_4995,N_4270);
xnor UO_785 (O_785,N_4562,N_4909);
or UO_786 (O_786,N_4535,N_4519);
xnor UO_787 (O_787,N_4207,N_4851);
and UO_788 (O_788,N_4806,N_4473);
nor UO_789 (O_789,N_4685,N_4988);
nand UO_790 (O_790,N_4857,N_4441);
nand UO_791 (O_791,N_4310,N_4056);
or UO_792 (O_792,N_4964,N_4610);
or UO_793 (O_793,N_4987,N_4576);
nand UO_794 (O_794,N_4891,N_4662);
or UO_795 (O_795,N_4052,N_4005);
xnor UO_796 (O_796,N_4903,N_4911);
nor UO_797 (O_797,N_4435,N_4634);
nor UO_798 (O_798,N_4551,N_4646);
nand UO_799 (O_799,N_4300,N_4869);
and UO_800 (O_800,N_4447,N_4592);
nor UO_801 (O_801,N_4299,N_4037);
xor UO_802 (O_802,N_4026,N_4450);
xnor UO_803 (O_803,N_4589,N_4175);
or UO_804 (O_804,N_4817,N_4256);
nor UO_805 (O_805,N_4016,N_4610);
and UO_806 (O_806,N_4038,N_4435);
xor UO_807 (O_807,N_4210,N_4663);
nor UO_808 (O_808,N_4625,N_4702);
and UO_809 (O_809,N_4825,N_4738);
xnor UO_810 (O_810,N_4157,N_4809);
xor UO_811 (O_811,N_4581,N_4050);
nand UO_812 (O_812,N_4434,N_4591);
or UO_813 (O_813,N_4178,N_4069);
nand UO_814 (O_814,N_4300,N_4821);
xnor UO_815 (O_815,N_4905,N_4759);
and UO_816 (O_816,N_4230,N_4615);
xor UO_817 (O_817,N_4761,N_4017);
or UO_818 (O_818,N_4726,N_4396);
nor UO_819 (O_819,N_4649,N_4751);
or UO_820 (O_820,N_4012,N_4206);
nand UO_821 (O_821,N_4003,N_4356);
and UO_822 (O_822,N_4321,N_4437);
nor UO_823 (O_823,N_4364,N_4679);
nor UO_824 (O_824,N_4064,N_4317);
or UO_825 (O_825,N_4674,N_4255);
nand UO_826 (O_826,N_4164,N_4711);
or UO_827 (O_827,N_4529,N_4172);
xnor UO_828 (O_828,N_4736,N_4404);
xor UO_829 (O_829,N_4098,N_4911);
xor UO_830 (O_830,N_4971,N_4509);
nand UO_831 (O_831,N_4374,N_4219);
and UO_832 (O_832,N_4605,N_4363);
xnor UO_833 (O_833,N_4747,N_4509);
nor UO_834 (O_834,N_4611,N_4511);
nand UO_835 (O_835,N_4400,N_4271);
and UO_836 (O_836,N_4776,N_4289);
nand UO_837 (O_837,N_4647,N_4260);
nand UO_838 (O_838,N_4339,N_4366);
nand UO_839 (O_839,N_4645,N_4117);
and UO_840 (O_840,N_4323,N_4186);
or UO_841 (O_841,N_4729,N_4464);
nor UO_842 (O_842,N_4823,N_4365);
and UO_843 (O_843,N_4338,N_4329);
and UO_844 (O_844,N_4765,N_4441);
xnor UO_845 (O_845,N_4495,N_4683);
nor UO_846 (O_846,N_4274,N_4554);
xnor UO_847 (O_847,N_4010,N_4789);
and UO_848 (O_848,N_4920,N_4092);
and UO_849 (O_849,N_4780,N_4740);
or UO_850 (O_850,N_4122,N_4349);
xor UO_851 (O_851,N_4077,N_4305);
nor UO_852 (O_852,N_4263,N_4620);
and UO_853 (O_853,N_4813,N_4408);
or UO_854 (O_854,N_4248,N_4718);
xnor UO_855 (O_855,N_4363,N_4229);
nor UO_856 (O_856,N_4549,N_4581);
nand UO_857 (O_857,N_4539,N_4994);
xor UO_858 (O_858,N_4498,N_4749);
nor UO_859 (O_859,N_4778,N_4858);
nand UO_860 (O_860,N_4040,N_4716);
or UO_861 (O_861,N_4545,N_4245);
nand UO_862 (O_862,N_4869,N_4315);
nor UO_863 (O_863,N_4500,N_4653);
xnor UO_864 (O_864,N_4143,N_4068);
nand UO_865 (O_865,N_4828,N_4301);
or UO_866 (O_866,N_4816,N_4792);
nand UO_867 (O_867,N_4192,N_4250);
xnor UO_868 (O_868,N_4138,N_4687);
xnor UO_869 (O_869,N_4245,N_4751);
nor UO_870 (O_870,N_4099,N_4888);
or UO_871 (O_871,N_4186,N_4118);
xnor UO_872 (O_872,N_4069,N_4062);
and UO_873 (O_873,N_4528,N_4017);
nand UO_874 (O_874,N_4481,N_4750);
xnor UO_875 (O_875,N_4186,N_4022);
nand UO_876 (O_876,N_4852,N_4737);
xnor UO_877 (O_877,N_4701,N_4104);
and UO_878 (O_878,N_4736,N_4194);
nor UO_879 (O_879,N_4420,N_4925);
and UO_880 (O_880,N_4849,N_4490);
nor UO_881 (O_881,N_4501,N_4774);
xnor UO_882 (O_882,N_4751,N_4452);
nor UO_883 (O_883,N_4884,N_4755);
xor UO_884 (O_884,N_4095,N_4272);
and UO_885 (O_885,N_4967,N_4828);
xnor UO_886 (O_886,N_4964,N_4240);
xor UO_887 (O_887,N_4773,N_4622);
and UO_888 (O_888,N_4621,N_4646);
nand UO_889 (O_889,N_4482,N_4302);
nand UO_890 (O_890,N_4664,N_4979);
or UO_891 (O_891,N_4031,N_4460);
nor UO_892 (O_892,N_4228,N_4014);
or UO_893 (O_893,N_4602,N_4386);
or UO_894 (O_894,N_4664,N_4400);
nor UO_895 (O_895,N_4080,N_4023);
nand UO_896 (O_896,N_4629,N_4122);
xor UO_897 (O_897,N_4577,N_4762);
xor UO_898 (O_898,N_4481,N_4936);
nand UO_899 (O_899,N_4043,N_4468);
nor UO_900 (O_900,N_4249,N_4003);
nor UO_901 (O_901,N_4592,N_4138);
nor UO_902 (O_902,N_4376,N_4139);
nor UO_903 (O_903,N_4984,N_4860);
or UO_904 (O_904,N_4495,N_4095);
xnor UO_905 (O_905,N_4666,N_4778);
and UO_906 (O_906,N_4617,N_4931);
or UO_907 (O_907,N_4689,N_4065);
nor UO_908 (O_908,N_4233,N_4216);
or UO_909 (O_909,N_4395,N_4513);
nand UO_910 (O_910,N_4200,N_4767);
or UO_911 (O_911,N_4135,N_4021);
or UO_912 (O_912,N_4099,N_4085);
or UO_913 (O_913,N_4015,N_4083);
nand UO_914 (O_914,N_4811,N_4006);
and UO_915 (O_915,N_4631,N_4390);
and UO_916 (O_916,N_4676,N_4718);
and UO_917 (O_917,N_4892,N_4415);
or UO_918 (O_918,N_4698,N_4932);
and UO_919 (O_919,N_4338,N_4432);
nor UO_920 (O_920,N_4738,N_4906);
and UO_921 (O_921,N_4882,N_4890);
nand UO_922 (O_922,N_4163,N_4927);
nand UO_923 (O_923,N_4105,N_4983);
nor UO_924 (O_924,N_4330,N_4545);
xor UO_925 (O_925,N_4028,N_4032);
nor UO_926 (O_926,N_4246,N_4228);
xor UO_927 (O_927,N_4205,N_4892);
nor UO_928 (O_928,N_4353,N_4045);
nor UO_929 (O_929,N_4805,N_4522);
nand UO_930 (O_930,N_4092,N_4478);
nor UO_931 (O_931,N_4048,N_4012);
nand UO_932 (O_932,N_4981,N_4713);
nand UO_933 (O_933,N_4048,N_4311);
and UO_934 (O_934,N_4931,N_4133);
xor UO_935 (O_935,N_4238,N_4367);
or UO_936 (O_936,N_4531,N_4765);
and UO_937 (O_937,N_4408,N_4543);
and UO_938 (O_938,N_4447,N_4946);
or UO_939 (O_939,N_4747,N_4361);
nor UO_940 (O_940,N_4973,N_4022);
nand UO_941 (O_941,N_4353,N_4478);
and UO_942 (O_942,N_4880,N_4889);
and UO_943 (O_943,N_4303,N_4085);
xor UO_944 (O_944,N_4833,N_4342);
and UO_945 (O_945,N_4984,N_4744);
nand UO_946 (O_946,N_4706,N_4136);
nor UO_947 (O_947,N_4388,N_4611);
nand UO_948 (O_948,N_4106,N_4263);
xnor UO_949 (O_949,N_4578,N_4970);
and UO_950 (O_950,N_4152,N_4871);
and UO_951 (O_951,N_4560,N_4008);
nand UO_952 (O_952,N_4265,N_4001);
nor UO_953 (O_953,N_4849,N_4475);
xor UO_954 (O_954,N_4088,N_4417);
nor UO_955 (O_955,N_4697,N_4275);
nand UO_956 (O_956,N_4592,N_4541);
nand UO_957 (O_957,N_4239,N_4703);
nand UO_958 (O_958,N_4151,N_4564);
xnor UO_959 (O_959,N_4804,N_4648);
nor UO_960 (O_960,N_4898,N_4370);
and UO_961 (O_961,N_4512,N_4479);
nand UO_962 (O_962,N_4319,N_4260);
nor UO_963 (O_963,N_4405,N_4135);
nand UO_964 (O_964,N_4138,N_4888);
nor UO_965 (O_965,N_4854,N_4656);
nor UO_966 (O_966,N_4628,N_4378);
nor UO_967 (O_967,N_4236,N_4749);
xnor UO_968 (O_968,N_4473,N_4683);
or UO_969 (O_969,N_4777,N_4253);
or UO_970 (O_970,N_4585,N_4387);
nand UO_971 (O_971,N_4190,N_4290);
xnor UO_972 (O_972,N_4810,N_4683);
nor UO_973 (O_973,N_4759,N_4352);
nor UO_974 (O_974,N_4817,N_4805);
nand UO_975 (O_975,N_4514,N_4463);
or UO_976 (O_976,N_4659,N_4385);
and UO_977 (O_977,N_4826,N_4148);
xor UO_978 (O_978,N_4660,N_4108);
xnor UO_979 (O_979,N_4932,N_4658);
nand UO_980 (O_980,N_4118,N_4976);
and UO_981 (O_981,N_4984,N_4175);
nand UO_982 (O_982,N_4622,N_4035);
or UO_983 (O_983,N_4358,N_4278);
and UO_984 (O_984,N_4999,N_4810);
xor UO_985 (O_985,N_4608,N_4823);
xnor UO_986 (O_986,N_4452,N_4685);
or UO_987 (O_987,N_4178,N_4464);
and UO_988 (O_988,N_4643,N_4109);
and UO_989 (O_989,N_4676,N_4008);
or UO_990 (O_990,N_4129,N_4441);
nand UO_991 (O_991,N_4425,N_4564);
or UO_992 (O_992,N_4879,N_4937);
nand UO_993 (O_993,N_4452,N_4239);
or UO_994 (O_994,N_4384,N_4885);
or UO_995 (O_995,N_4604,N_4198);
nand UO_996 (O_996,N_4416,N_4792);
xnor UO_997 (O_997,N_4642,N_4828);
nor UO_998 (O_998,N_4887,N_4359);
nor UO_999 (O_999,N_4358,N_4846);
endmodule