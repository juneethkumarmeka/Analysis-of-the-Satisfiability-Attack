module basic_1000_10000_1500_50_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_301,In_161);
nor U1 (N_1,In_936,In_984);
or U2 (N_2,In_30,In_295);
or U3 (N_3,In_189,In_364);
xor U4 (N_4,In_365,In_659);
or U5 (N_5,In_347,In_491);
nor U6 (N_6,In_709,In_706);
nand U7 (N_7,In_985,In_44);
nor U8 (N_8,In_929,In_316);
and U9 (N_9,In_11,In_93);
nor U10 (N_10,In_398,In_819);
xor U11 (N_11,In_426,In_27);
and U12 (N_12,In_256,In_235);
and U13 (N_13,In_852,In_163);
or U14 (N_14,In_568,In_176);
and U15 (N_15,In_26,In_296);
xor U16 (N_16,In_278,In_68);
and U17 (N_17,In_135,In_81);
nand U18 (N_18,In_995,In_197);
xor U19 (N_19,In_841,In_905);
and U20 (N_20,In_320,In_818);
or U21 (N_21,In_540,In_638);
nor U22 (N_22,In_720,In_875);
nand U23 (N_23,In_39,In_501);
and U24 (N_24,In_116,In_331);
or U25 (N_25,In_496,In_721);
nor U26 (N_26,In_591,In_505);
nor U27 (N_27,In_752,In_503);
or U28 (N_28,In_140,In_238);
nand U29 (N_29,In_959,In_784);
or U30 (N_30,In_334,In_722);
and U31 (N_31,In_631,In_242);
nor U32 (N_32,In_408,In_147);
or U33 (N_33,In_732,In_343);
or U34 (N_34,In_705,In_53);
or U35 (N_35,In_828,In_155);
xnor U36 (N_36,In_356,In_225);
nor U37 (N_37,In_166,In_739);
and U38 (N_38,In_461,In_774);
nor U39 (N_39,In_867,In_223);
or U40 (N_40,In_972,In_891);
or U41 (N_41,In_648,In_727);
or U42 (N_42,In_282,In_847);
xnor U43 (N_43,In_96,In_649);
and U44 (N_44,In_178,In_59);
xor U45 (N_45,In_872,In_866);
and U46 (N_46,In_766,In_547);
or U47 (N_47,In_824,In_629);
or U48 (N_48,In_719,In_634);
nand U49 (N_49,In_779,In_133);
or U50 (N_50,In_758,In_640);
nand U51 (N_51,In_661,In_536);
xor U52 (N_52,In_506,In_160);
nand U53 (N_53,In_453,In_676);
nor U54 (N_54,In_77,In_479);
and U55 (N_55,In_437,In_3);
xor U56 (N_56,In_978,In_548);
or U57 (N_57,In_761,In_152);
or U58 (N_58,In_252,In_965);
and U59 (N_59,In_181,In_558);
or U60 (N_60,In_877,In_300);
nor U61 (N_61,In_478,In_74);
nand U62 (N_62,In_336,In_968);
nor U63 (N_63,In_401,In_349);
or U64 (N_64,In_931,In_693);
or U65 (N_65,In_352,In_864);
or U66 (N_66,In_2,In_660);
and U67 (N_67,In_345,In_517);
nand U68 (N_68,In_645,In_470);
nand U69 (N_69,In_246,In_249);
and U70 (N_70,In_962,In_359);
xnor U71 (N_71,In_725,In_159);
or U72 (N_72,In_520,In_707);
and U73 (N_73,In_441,In_70);
nor U74 (N_74,In_753,In_554);
nand U75 (N_75,In_283,In_613);
and U76 (N_76,In_534,In_251);
xor U77 (N_77,In_66,In_512);
xor U78 (N_78,In_783,In_52);
and U79 (N_79,In_432,In_179);
nand U80 (N_80,In_342,In_610);
and U81 (N_81,In_583,In_887);
xor U82 (N_82,In_522,In_746);
xor U83 (N_83,In_333,In_620);
or U84 (N_84,In_876,In_101);
nand U85 (N_85,In_107,In_786);
nor U86 (N_86,In_371,In_997);
xnor U87 (N_87,In_628,In_466);
or U88 (N_88,In_400,In_712);
and U89 (N_89,In_763,In_217);
nand U90 (N_90,In_399,In_48);
nand U91 (N_91,In_357,In_942);
and U92 (N_92,In_190,In_324);
and U93 (N_93,In_0,In_102);
nor U94 (N_94,In_148,In_290);
nor U95 (N_95,In_224,In_380);
or U96 (N_96,In_288,In_539);
or U97 (N_97,In_430,In_406);
nor U98 (N_98,In_618,In_92);
or U99 (N_99,In_105,In_913);
and U100 (N_100,In_428,In_254);
and U101 (N_101,In_790,In_695);
xor U102 (N_102,In_553,In_668);
or U103 (N_103,In_464,In_142);
nand U104 (N_104,In_797,In_507);
nor U105 (N_105,In_270,In_384);
nor U106 (N_106,In_767,In_210);
or U107 (N_107,In_827,In_173);
or U108 (N_108,In_346,In_260);
and U109 (N_109,In_80,In_396);
xor U110 (N_110,In_622,In_986);
nand U111 (N_111,In_976,In_216);
or U112 (N_112,In_945,In_938);
nand U113 (N_113,In_355,In_136);
or U114 (N_114,In_188,In_897);
and U115 (N_115,In_459,In_287);
and U116 (N_116,In_570,In_61);
or U117 (N_117,In_647,In_344);
and U118 (N_118,In_76,In_350);
or U119 (N_119,In_171,In_861);
nand U120 (N_120,In_374,In_574);
and U121 (N_121,In_881,In_332);
xnor U122 (N_122,In_185,In_996);
or U123 (N_123,In_89,In_741);
nand U124 (N_124,In_697,In_497);
and U125 (N_125,In_234,In_12);
or U126 (N_126,In_530,In_502);
or U127 (N_127,In_9,In_838);
nor U128 (N_128,In_713,In_311);
or U129 (N_129,In_259,In_604);
nor U130 (N_130,In_429,In_751);
nand U131 (N_131,In_499,In_5);
nand U132 (N_132,In_184,In_199);
or U133 (N_133,In_131,In_949);
nand U134 (N_134,In_918,In_851);
xor U135 (N_135,In_928,In_327);
nand U136 (N_136,In_518,In_277);
and U137 (N_137,In_800,In_420);
nor U138 (N_138,In_941,In_271);
nor U139 (N_139,In_439,In_337);
and U140 (N_140,In_36,In_34);
xor U141 (N_141,In_360,In_273);
or U142 (N_142,In_383,In_314);
or U143 (N_143,In_636,In_873);
xnor U144 (N_144,In_33,In_267);
and U145 (N_145,In_966,In_586);
nand U146 (N_146,In_961,In_381);
nor U147 (N_147,In_25,In_672);
and U148 (N_148,In_681,In_58);
nor U149 (N_149,In_389,In_51);
or U150 (N_150,In_750,In_983);
or U151 (N_151,In_494,In_504);
and U152 (N_152,In_122,In_35);
nor U153 (N_153,In_233,In_117);
nor U154 (N_154,In_963,In_885);
nand U155 (N_155,In_291,In_729);
nor U156 (N_156,In_444,In_943);
and U157 (N_157,In_987,In_994);
nor U158 (N_158,In_403,In_262);
nor U159 (N_159,In_687,In_696);
or U160 (N_160,In_509,In_261);
nand U161 (N_161,In_734,In_702);
nor U162 (N_162,In_169,In_286);
nand U163 (N_163,In_576,In_829);
nand U164 (N_164,In_678,In_351);
and U165 (N_165,In_328,In_47);
nand U166 (N_166,In_607,In_85);
xor U167 (N_167,In_674,In_840);
nor U168 (N_168,In_368,In_15);
nor U169 (N_169,In_529,In_258);
nand U170 (N_170,In_498,In_95);
nand U171 (N_171,In_546,In_206);
nand U172 (N_172,In_888,In_665);
nand U173 (N_173,In_569,In_410);
or U174 (N_174,In_572,In_728);
nand U175 (N_175,In_652,In_526);
or U176 (N_176,In_532,In_198);
or U177 (N_177,In_407,In_375);
nor U178 (N_178,In_670,In_780);
or U179 (N_179,In_550,In_99);
xor U180 (N_180,In_632,In_192);
or U181 (N_181,In_757,In_402);
and U182 (N_182,In_462,In_513);
nor U183 (N_183,In_606,In_880);
nor U184 (N_184,In_874,In_971);
xnor U185 (N_185,In_748,In_203);
or U186 (N_186,In_807,In_10);
and U187 (N_187,In_998,In_157);
or U188 (N_188,In_635,In_730);
nor U189 (N_189,In_377,In_394);
nand U190 (N_190,In_326,In_165);
nor U191 (N_191,In_71,In_643);
nand U192 (N_192,In_870,In_717);
nand U193 (N_193,In_651,In_759);
nand U194 (N_194,In_822,In_97);
nand U195 (N_195,In_538,In_280);
nand U196 (N_196,In_685,In_654);
and U197 (N_197,In_7,In_611);
xnor U198 (N_198,In_162,In_213);
or U199 (N_199,In_833,In_57);
and U200 (N_200,N_40,N_193);
nand U201 (N_201,In_603,In_835);
nor U202 (N_202,In_832,N_86);
xnor U203 (N_203,In_901,In_979);
nor U204 (N_204,N_1,N_95);
or U205 (N_205,In_912,In_955);
and U206 (N_206,In_825,In_718);
and U207 (N_207,In_49,In_125);
nand U208 (N_208,N_184,In_521);
and U209 (N_209,N_165,In_202);
nand U210 (N_210,In_883,In_531);
and U211 (N_211,In_372,In_698);
or U212 (N_212,In_682,In_970);
nand U213 (N_213,In_699,In_329);
or U214 (N_214,N_70,In_805);
nor U215 (N_215,N_187,In_17);
nor U216 (N_216,N_147,N_34);
or U217 (N_217,In_898,In_303);
xnor U218 (N_218,In_473,N_136);
xnor U219 (N_219,N_125,In_78);
and U220 (N_220,In_793,N_115);
and U221 (N_221,In_804,In_341);
nand U222 (N_222,In_519,In_83);
and U223 (N_223,N_83,N_109);
and U224 (N_224,In_951,In_692);
nor U225 (N_225,In_795,In_680);
and U226 (N_226,N_75,In_386);
nand U227 (N_227,N_188,In_879);
xnor U228 (N_228,In_777,N_120);
xnor U229 (N_229,In_361,In_156);
nor U230 (N_230,N_92,In_967);
and U231 (N_231,In_541,In_16);
and U232 (N_232,In_416,In_222);
or U233 (N_233,N_38,In_743);
nand U234 (N_234,N_174,N_194);
or U235 (N_235,In_684,N_69);
nor U236 (N_236,N_51,In_299);
or U237 (N_237,In_164,N_94);
and U238 (N_238,In_485,In_425);
or U239 (N_239,N_41,N_107);
or U240 (N_240,In_481,In_276);
nand U241 (N_241,In_714,N_55);
or U242 (N_242,In_281,In_561);
nor U243 (N_243,N_185,In_592);
nand U244 (N_244,In_476,In_193);
or U245 (N_245,In_307,N_84);
nor U246 (N_246,In_373,In_88);
nand U247 (N_247,In_305,N_143);
or U248 (N_248,N_71,N_133);
and U249 (N_249,N_131,In_239);
or U250 (N_250,In_627,In_863);
nand U251 (N_251,N_35,In_977);
and U252 (N_252,N_42,N_47);
nor U253 (N_253,In_150,In_397);
xor U254 (N_254,In_419,N_58);
or U255 (N_255,N_171,N_2);
or U256 (N_256,N_130,In_735);
nor U257 (N_257,In_960,In_435);
nand U258 (N_258,In_23,In_91);
nor U259 (N_259,In_447,N_192);
or U260 (N_260,In_808,N_112);
nor U261 (N_261,In_220,In_657);
xor U262 (N_262,N_161,In_289);
nand U263 (N_263,In_796,In_694);
and U264 (N_264,N_46,N_148);
nand U265 (N_265,In_310,In_500);
and U266 (N_266,In_566,In_230);
or U267 (N_267,In_975,N_50);
nand U268 (N_268,In_658,In_857);
or U269 (N_269,In_988,In_268);
or U270 (N_270,In_826,N_106);
or U271 (N_271,N_72,N_65);
nor U272 (N_272,In_686,In_475);
nand U273 (N_273,In_940,N_9);
nor U274 (N_274,In_323,N_162);
and U275 (N_275,In_191,N_199);
and U276 (N_276,In_846,In_134);
or U277 (N_277,N_26,In_791);
nor U278 (N_278,N_63,N_186);
nand U279 (N_279,In_882,In_815);
nor U280 (N_280,In_151,N_167);
xor U281 (N_281,In_950,In_257);
and U282 (N_282,In_524,In_322);
nor U283 (N_283,In_411,In_992);
and U284 (N_284,In_892,In_528);
nand U285 (N_285,In_132,In_584);
nor U286 (N_286,In_449,N_93);
nor U287 (N_287,In_820,In_465);
and U288 (N_288,In_590,In_409);
nand U289 (N_289,In_123,In_72);
nand U290 (N_290,N_15,N_8);
nand U291 (N_291,In_656,In_294);
nor U292 (N_292,In_902,In_480);
nor U293 (N_293,In_226,In_585);
nand U294 (N_294,In_460,In_770);
or U295 (N_295,In_515,In_608);
nand U296 (N_296,N_88,In_196);
nor U297 (N_297,In_218,N_110);
nand U298 (N_298,In_798,In_842);
and U299 (N_299,In_919,N_138);
or U300 (N_300,In_339,In_382);
nand U301 (N_301,N_96,In_803);
or U302 (N_302,In_121,In_204);
nand U303 (N_303,N_52,In_571);
xor U304 (N_304,In_456,In_124);
nand U305 (N_305,In_20,In_890);
xnor U306 (N_306,In_306,In_544);
or U307 (N_307,In_236,N_191);
and U308 (N_308,In_392,In_492);
nor U309 (N_309,In_947,N_16);
nand U310 (N_310,In_688,In_4);
and U311 (N_311,In_921,N_183);
and U312 (N_312,In_338,In_231);
or U313 (N_313,In_981,N_166);
nand U314 (N_314,In_84,In_484);
and U315 (N_315,N_5,In_565);
and U316 (N_316,In_293,In_559);
nand U317 (N_317,In_600,In_415);
xor U318 (N_318,N_179,In_340);
or U319 (N_319,In_785,In_749);
xor U320 (N_320,N_173,In_733);
nor U321 (N_321,N_78,In_922);
nor U322 (N_322,In_555,In_811);
nor U323 (N_323,In_745,In_272);
nor U324 (N_324,In_621,In_809);
or U325 (N_325,In_445,In_208);
or U326 (N_326,N_198,In_109);
nor U327 (N_327,N_49,In_302);
and U328 (N_328,In_335,In_45);
or U329 (N_329,In_508,N_87);
or U330 (N_330,In_209,In_557);
and U331 (N_331,N_27,In_40);
nor U332 (N_332,In_450,In_358);
and U333 (N_333,In_917,In_724);
and U334 (N_334,In_391,In_510);
and U335 (N_335,N_14,In_683);
and U336 (N_336,In_599,N_104);
and U337 (N_337,In_247,In_556);
nand U338 (N_338,In_738,In_212);
nor U339 (N_339,In_655,In_630);
and U340 (N_340,In_637,In_845);
and U341 (N_341,In_639,In_653);
or U342 (N_342,N_66,In_442);
and U343 (N_343,In_756,N_150);
and U344 (N_344,In_137,In_22);
and U345 (N_345,In_830,In_642);
nor U346 (N_346,N_175,N_168);
nor U347 (N_347,In_810,N_141);
nand U348 (N_348,N_29,In_103);
and U349 (N_349,In_376,In_413);
nand U350 (N_350,In_646,In_228);
nor U351 (N_351,N_157,N_44);
xnor U352 (N_352,N_23,N_81);
or U353 (N_353,In_390,In_769);
nor U354 (N_354,N_25,In_274);
nor U355 (N_355,In_595,In_205);
nand U356 (N_356,In_55,N_56);
or U357 (N_357,In_250,In_726);
nor U358 (N_358,In_38,In_862);
xnor U359 (N_359,In_284,In_100);
and U360 (N_360,In_991,In_982);
nand U361 (N_361,N_164,In_241);
or U362 (N_362,In_207,In_31);
nand U363 (N_363,In_737,N_32);
nor U364 (N_364,In_754,In_113);
or U365 (N_365,In_127,In_596);
and U366 (N_366,In_904,N_24);
and U367 (N_367,In_836,In_736);
xor U368 (N_368,In_602,In_666);
xor U369 (N_369,In_29,N_82);
and U370 (N_370,In_889,In_703);
xor U371 (N_371,In_926,In_317);
and U372 (N_372,N_118,In_451);
nand U373 (N_373,In_412,In_187);
or U374 (N_374,In_363,N_31);
or U375 (N_375,In_138,N_61);
xor U376 (N_376,In_446,In_844);
nand U377 (N_377,In_141,In_46);
and U378 (N_378,N_169,N_33);
nor U379 (N_379,N_181,In_298);
or U380 (N_380,In_248,In_860);
nand U381 (N_381,In_952,In_90);
or U382 (N_382,In_186,N_64);
and U383 (N_383,In_395,In_60);
and U384 (N_384,In_579,In_495);
or U385 (N_385,N_36,N_13);
nor U386 (N_386,In_581,In_549);
nand U387 (N_387,N_43,In_909);
xor U388 (N_388,In_839,In_969);
and U389 (N_389,In_886,In_980);
and U390 (N_390,N_48,In_14);
xor U391 (N_391,N_105,In_41);
xnor U392 (N_392,In_454,In_617);
xor U393 (N_393,N_12,In_716);
and U394 (N_394,In_935,In_848);
and U395 (N_395,In_62,N_177);
nor U396 (N_396,N_128,In_482);
xnor U397 (N_397,In_812,N_60);
or U398 (N_398,In_823,In_414);
nor U399 (N_399,In_417,In_474);
nand U400 (N_400,N_6,N_159);
nand U401 (N_401,In_689,In_787);
or U402 (N_402,N_242,In_675);
or U403 (N_403,N_277,N_151);
nand U404 (N_404,In_43,In_219);
nor U405 (N_405,N_3,In_993);
or U406 (N_406,In_370,In_195);
or U407 (N_407,N_114,N_222);
nand U408 (N_408,N_360,In_575);
and U409 (N_409,N_202,N_366);
nor U410 (N_410,N_170,In_948);
or U411 (N_411,N_37,In_463);
or U412 (N_412,N_137,N_227);
nor U413 (N_413,In_667,In_623);
and U414 (N_414,N_234,N_388);
nand U415 (N_415,In_990,N_196);
or U416 (N_416,In_799,N_383);
nor U417 (N_417,In_782,In_330);
or U418 (N_418,N_250,In_94);
or U419 (N_419,In_69,N_211);
or U420 (N_420,In_180,In_167);
nor U421 (N_421,In_120,In_850);
nor U422 (N_422,N_97,In_292);
or U423 (N_423,In_564,In_143);
nand U424 (N_424,N_190,N_89);
xor U425 (N_425,N_356,N_375);
and U426 (N_426,N_99,N_284);
and U427 (N_427,In_663,N_342);
nand U428 (N_428,In_469,In_149);
and U429 (N_429,N_270,N_321);
xnor U430 (N_430,N_397,In_854);
and U431 (N_431,N_243,N_180);
nand U432 (N_432,In_255,In_42);
or U433 (N_433,In_582,In_768);
or U434 (N_434,In_128,In_910);
nor U435 (N_435,In_900,N_272);
nor U436 (N_436,In_457,In_269);
and U437 (N_437,In_934,In_243);
nor U438 (N_438,In_440,N_382);
nor U439 (N_439,N_280,N_304);
nor U440 (N_440,N_100,N_214);
nor U441 (N_441,N_11,N_252);
or U442 (N_442,In_755,In_514);
and U443 (N_443,In_894,N_249);
and U444 (N_444,In_899,In_711);
or U445 (N_445,In_831,N_379);
xnor U446 (N_446,In_858,In_221);
nand U447 (N_447,In_773,In_616);
or U448 (N_448,In_421,N_163);
or U449 (N_449,In_263,In_488);
nor U450 (N_450,In_625,In_563);
or U451 (N_451,In_775,In_816);
and U452 (N_452,In_609,In_79);
nor U453 (N_453,In_927,N_343);
or U454 (N_454,In_789,N_45);
nor U455 (N_455,N_248,N_74);
nand U456 (N_456,N_232,In_664);
nand U457 (N_457,In_974,In_232);
and U458 (N_458,In_778,N_331);
or U459 (N_459,N_158,N_153);
nor U460 (N_460,N_327,N_390);
and U461 (N_461,N_309,In_455);
nand U462 (N_462,In_601,In_244);
or U463 (N_463,In_8,In_423);
and U464 (N_464,N_355,In_170);
nor U465 (N_465,In_129,In_126);
or U466 (N_466,In_366,In_379);
and U467 (N_467,N_296,In_597);
xor U468 (N_468,In_434,N_119);
and U469 (N_469,In_710,N_73);
or U470 (N_470,N_189,In_806);
nor U471 (N_471,In_471,N_123);
nor U472 (N_472,N_79,In_953);
nand U473 (N_473,N_121,In_859);
xor U474 (N_474,N_365,N_98);
and U475 (N_475,N_377,N_67);
and U476 (N_476,N_253,N_329);
nor U477 (N_477,N_347,In_431);
and U478 (N_478,N_283,N_62);
nor U479 (N_479,In_1,N_221);
nand U480 (N_480,N_247,N_350);
nand U481 (N_481,In_545,In_916);
or U482 (N_482,In_662,N_129);
or U483 (N_483,N_57,N_320);
or U484 (N_484,In_452,In_427);
and U485 (N_485,In_318,In_615);
or U486 (N_486,N_391,N_257);
nand U487 (N_487,In_158,In_624);
or U488 (N_488,N_200,N_235);
and U489 (N_489,N_373,In_560);
and U490 (N_490,In_487,In_13);
nor U491 (N_491,In_468,In_868);
and U492 (N_492,N_259,N_28);
nor U493 (N_493,N_239,N_325);
and U494 (N_494,In_849,In_747);
xnor U495 (N_495,N_231,N_18);
nand U496 (N_496,N_359,N_140);
xor U497 (N_497,In_201,In_884);
and U498 (N_498,In_211,In_56);
nor U499 (N_499,In_325,In_106);
xnor U500 (N_500,N_240,In_920);
or U501 (N_501,N_274,In_587);
and U502 (N_502,In_788,N_357);
and U503 (N_503,In_973,In_650);
nand U504 (N_504,In_438,N_364);
or U505 (N_505,N_363,In_297);
nand U506 (N_506,N_335,In_855);
and U507 (N_507,In_939,In_312);
nand U508 (N_508,In_145,In_893);
xor U509 (N_509,In_673,In_764);
or U510 (N_510,In_153,N_127);
and U511 (N_511,In_865,In_144);
or U512 (N_512,N_381,In_633);
or U513 (N_513,In_177,N_340);
and U514 (N_514,In_37,N_220);
nor U515 (N_515,N_156,N_53);
nand U516 (N_516,In_906,N_288);
and U517 (N_517,In_229,In_467);
nor U518 (N_518,N_395,N_113);
nand U519 (N_519,In_75,In_580);
nand U520 (N_520,N_228,N_217);
or U521 (N_521,In_516,In_458);
nand U522 (N_522,In_6,In_19);
xor U523 (N_523,In_598,In_869);
or U524 (N_524,N_116,In_619);
or U525 (N_525,N_351,N_68);
nor U526 (N_526,N_368,In_265);
and U527 (N_527,N_144,In_527);
nor U528 (N_528,N_339,In_551);
nor U529 (N_529,In_112,N_205);
or U530 (N_530,N_367,In_393);
or U531 (N_531,N_254,In_802);
nand U532 (N_532,N_142,In_511);
nand U533 (N_533,N_337,In_175);
or U534 (N_534,N_178,N_393);
or U535 (N_535,N_302,In_944);
and U536 (N_536,N_17,In_63);
or U537 (N_537,N_374,In_24);
or U538 (N_538,N_91,N_260);
xor U539 (N_539,In_933,N_307);
and U540 (N_540,In_237,In_701);
nor U541 (N_541,In_543,In_275);
xor U542 (N_542,N_349,In_813);
xor U543 (N_543,In_227,N_384);
nor U544 (N_544,In_50,N_385);
and U545 (N_545,In_154,N_266);
or U546 (N_546,N_286,In_264);
and U547 (N_547,In_958,N_297);
nand U548 (N_548,In_28,N_273);
or U549 (N_549,In_490,N_216);
or U550 (N_550,N_230,N_258);
or U551 (N_551,N_263,N_103);
nor U552 (N_552,In_486,In_573);
or U553 (N_553,N_326,In_82);
xor U554 (N_554,N_264,N_241);
or U555 (N_555,N_275,In_614);
and U556 (N_556,N_224,In_925);
xor U557 (N_557,N_305,In_433);
nor U558 (N_558,In_535,In_385);
nand U559 (N_559,N_208,N_330);
nand U560 (N_560,In_567,N_289);
xor U561 (N_561,In_215,In_723);
nand U562 (N_562,N_358,N_352);
nand U563 (N_563,N_149,In_304);
nand U564 (N_564,N_346,N_313);
or U565 (N_565,N_197,In_525);
and U566 (N_566,In_362,N_21);
nor U567 (N_567,In_168,In_146);
or U568 (N_568,N_262,N_246);
nand U569 (N_569,In_448,In_483);
and U570 (N_570,In_436,N_396);
or U571 (N_571,In_989,N_212);
xnor U572 (N_572,In_878,In_86);
or U573 (N_573,In_915,In_700);
xor U574 (N_574,In_605,In_671);
or U575 (N_575,In_588,In_577);
and U576 (N_576,N_244,In_73);
and U577 (N_577,In_908,N_182);
and U578 (N_578,N_176,N_236);
and U579 (N_579,In_776,In_87);
or U580 (N_580,N_267,N_387);
nor U581 (N_581,In_139,In_64);
nor U582 (N_582,In_896,N_206);
nor U583 (N_583,N_344,In_315);
or U584 (N_584,In_489,In_856);
nand U585 (N_585,In_194,In_612);
and U586 (N_586,N_10,N_237);
xnor U587 (N_587,N_299,In_477);
xnor U588 (N_588,N_317,N_281);
and U589 (N_589,N_392,In_279);
and U590 (N_590,In_378,In_321);
and U591 (N_591,N_345,N_152);
nor U592 (N_592,N_295,In_253);
nand U593 (N_593,N_315,N_19);
or U594 (N_594,In_794,N_308);
or U595 (N_595,In_914,In_937);
or U596 (N_596,N_255,In_443);
or U597 (N_597,N_135,N_7);
or U598 (N_598,In_814,N_332);
nand U599 (N_599,N_324,N_245);
and U600 (N_600,N_515,In_110);
nand U601 (N_601,In_593,N_77);
nand U602 (N_602,In_367,N_204);
or U603 (N_603,In_911,In_245);
nand U604 (N_604,N_334,N_425);
nor U605 (N_605,In_626,N_565);
nand U606 (N_606,In_762,N_400);
nand U607 (N_607,In_744,N_533);
and U608 (N_608,N_432,N_539);
and U609 (N_609,N_469,In_853);
and U610 (N_610,N_428,N_207);
nand U611 (N_611,In_98,N_416);
nand U612 (N_612,N_54,N_585);
nor U613 (N_613,N_434,N_333);
or U614 (N_614,N_422,N_209);
nand U615 (N_615,N_303,N_453);
xor U616 (N_616,N_80,In_932);
nand U617 (N_617,N_146,In_353);
nor U618 (N_618,N_338,N_477);
and U619 (N_619,N_459,N_445);
nand U620 (N_620,N_436,N_537);
nand U621 (N_621,N_456,N_22);
nor U622 (N_622,N_420,N_446);
and U623 (N_623,N_160,N_215);
and U624 (N_624,N_501,N_386);
and U625 (N_625,N_348,N_201);
xnor U626 (N_626,In_533,N_462);
and U627 (N_627,N_59,N_576);
and U628 (N_628,N_291,N_450);
nor U629 (N_629,N_492,In_319);
xor U630 (N_630,N_490,N_117);
nand U631 (N_631,N_361,N_418);
nand U632 (N_632,N_398,In_404);
nand U633 (N_633,N_526,N_323);
nor U634 (N_634,N_582,N_485);
nand U635 (N_635,N_172,N_213);
or U636 (N_636,N_573,N_543);
nor U637 (N_637,In_200,N_592);
nor U638 (N_638,N_455,N_522);
nand U639 (N_639,In_114,N_285);
xnor U640 (N_640,N_558,N_440);
nand U641 (N_641,N_591,In_895);
and U642 (N_642,N_225,N_532);
and U643 (N_643,N_85,N_541);
xnor U644 (N_644,In_907,N_486);
and U645 (N_645,In_641,N_403);
or U646 (N_646,N_139,In_523);
nand U647 (N_647,In_309,N_473);
xnor U648 (N_648,In_313,N_513);
nor U649 (N_649,N_101,N_482);
and U650 (N_650,N_419,N_322);
or U651 (N_651,N_540,N_569);
nand U652 (N_652,N_427,In_32);
xor U653 (N_653,In_183,N_354);
nand U654 (N_654,N_538,N_238);
nand U655 (N_655,In_837,N_406);
nor U656 (N_656,N_411,In_537);
and U657 (N_657,N_475,N_504);
nor U658 (N_658,In_957,N_488);
nor U659 (N_659,N_512,N_546);
or U660 (N_660,N_404,N_226);
nor U661 (N_661,N_598,In_104);
nor U662 (N_662,N_536,N_219);
nand U663 (N_663,N_528,In_493);
and U664 (N_664,In_115,N_506);
and U665 (N_665,N_353,N_568);
and U666 (N_666,N_531,N_424);
nor U667 (N_667,N_124,N_499);
nand U668 (N_668,N_479,N_596);
xor U669 (N_669,N_559,N_447);
or U670 (N_670,N_122,N_4);
nand U671 (N_671,N_599,N_437);
or U672 (N_672,N_502,N_414);
and U673 (N_673,N_500,In_21);
nand U674 (N_674,N_561,N_282);
or U675 (N_675,N_497,N_401);
nor U676 (N_676,N_464,N_76);
or U677 (N_677,N_594,N_495);
nor U678 (N_678,In_821,In_424);
or U679 (N_679,N_318,In_964);
nor U680 (N_680,N_514,N_20);
and U681 (N_681,In_387,N_0);
and U682 (N_682,In_817,In_308);
nand U683 (N_683,N_470,N_567);
nor U684 (N_684,N_218,N_452);
xnor U685 (N_685,N_589,N_465);
and U686 (N_686,In_644,N_442);
nand U687 (N_687,In_801,N_430);
nor U688 (N_688,N_265,In_214);
nand U689 (N_689,In_552,N_145);
xor U690 (N_690,N_544,In_108);
or U691 (N_691,In_130,In_781);
and U692 (N_692,N_566,N_505);
or U693 (N_693,N_410,N_551);
and U694 (N_694,N_341,N_578);
or U695 (N_695,N_510,N_300);
nand U696 (N_696,N_271,N_287);
nor U697 (N_697,N_223,N_461);
and U698 (N_698,N_278,N_586);
nor U699 (N_699,N_517,In_871);
nand U700 (N_700,N_39,N_523);
nor U701 (N_701,N_376,N_463);
nand U702 (N_702,N_203,N_415);
nand U703 (N_703,N_380,In_354);
xor U704 (N_704,In_930,N_597);
and U705 (N_705,In_388,N_412);
nand U706 (N_706,N_555,N_328);
or U707 (N_707,N_579,N_507);
or U708 (N_708,N_549,N_583);
xor U709 (N_709,N_575,N_493);
nand U710 (N_710,N_229,N_562);
nand U711 (N_711,N_276,In_348);
and U712 (N_712,N_316,N_574);
nor U713 (N_713,N_30,N_441);
nand U714 (N_714,In_946,N_298);
and U715 (N_715,N_134,N_449);
nor U716 (N_716,N_268,N_476);
nor U717 (N_717,In_118,N_108);
nor U718 (N_718,N_256,N_571);
nor U719 (N_719,In_111,N_496);
or U720 (N_720,N_433,N_478);
or U721 (N_721,N_483,In_999);
and U722 (N_722,N_511,In_669);
and U723 (N_723,In_172,In_18);
xor U724 (N_724,N_527,N_155);
nand U725 (N_725,N_399,N_516);
nand U726 (N_726,In_679,In_174);
nand U727 (N_727,In_765,N_314);
nor U728 (N_728,N_491,N_269);
xor U729 (N_729,In_715,In_405);
nor U730 (N_730,N_439,N_294);
nor U731 (N_731,In_690,N_293);
or U732 (N_732,N_407,N_154);
nor U733 (N_733,N_458,In_266);
and U734 (N_734,N_556,N_413);
and U735 (N_735,N_448,N_372);
or U736 (N_736,In_119,In_677);
or U737 (N_737,In_67,N_306);
and U738 (N_738,N_560,N_443);
or U739 (N_739,N_311,N_519);
or U740 (N_740,N_261,N_534);
xor U741 (N_741,In_542,N_529);
and U742 (N_742,N_292,In_691);
nand U743 (N_743,N_570,N_487);
xnor U744 (N_744,In_954,N_467);
nor U745 (N_745,N_279,In_742);
nor U746 (N_746,N_409,In_472);
or U747 (N_747,N_417,N_378);
xor U748 (N_748,N_498,N_548);
nor U749 (N_749,N_588,In_771);
nor U750 (N_750,N_474,N_429);
nor U751 (N_751,N_550,In_903);
nor U752 (N_752,N_484,N_444);
nand U753 (N_753,N_290,In_731);
nand U754 (N_754,N_369,N_545);
or U755 (N_755,N_584,N_389);
nand U756 (N_756,N_521,N_195);
nor U757 (N_757,N_251,N_454);
and U758 (N_758,N_563,N_408);
and U759 (N_759,N_564,N_435);
nand U760 (N_760,N_319,N_489);
and U761 (N_761,N_553,In_54);
nand U762 (N_762,N_402,In_369);
nor U763 (N_763,N_595,In_418);
or U764 (N_764,N_233,N_587);
or U765 (N_765,N_210,N_301);
nand U766 (N_766,N_480,In_578);
xor U767 (N_767,N_472,N_310);
nor U768 (N_768,N_431,N_370);
or U769 (N_769,N_468,N_593);
nor U770 (N_770,N_312,In_65);
and U771 (N_771,In_834,N_508);
nand U772 (N_772,N_518,N_394);
nor U773 (N_773,In_704,N_132);
or U774 (N_774,N_552,N_426);
xnor U775 (N_775,In_562,N_451);
or U776 (N_776,N_466,N_471);
nor U777 (N_777,N_577,In_708);
and U778 (N_778,N_530,N_581);
and U779 (N_779,N_503,In_792);
nand U780 (N_780,N_362,N_547);
nor U781 (N_781,In_240,N_90);
or U782 (N_782,N_520,N_580);
nand U783 (N_783,N_524,N_590);
nor U784 (N_784,In_589,N_336);
nand U785 (N_785,In_772,N_535);
and U786 (N_786,In_760,N_557);
nand U787 (N_787,N_405,In_956);
nor U788 (N_788,N_542,N_572);
nand U789 (N_789,N_126,N_457);
or U790 (N_790,N_494,N_371);
nor U791 (N_791,N_421,N_509);
nand U792 (N_792,In_843,N_111);
nor U793 (N_793,N_423,N_525);
nand U794 (N_794,N_460,N_438);
and U795 (N_795,In_594,In_740);
nand U796 (N_796,In_182,N_102);
nand U797 (N_797,In_422,In_285);
nor U798 (N_798,In_923,N_481);
or U799 (N_799,N_554,In_924);
nor U800 (N_800,N_718,N_700);
nand U801 (N_801,N_731,N_641);
nor U802 (N_802,N_760,N_741);
xnor U803 (N_803,N_695,N_603);
nor U804 (N_804,N_656,N_638);
or U805 (N_805,N_605,N_694);
and U806 (N_806,N_787,N_683);
nor U807 (N_807,N_721,N_708);
nand U808 (N_808,N_793,N_719);
or U809 (N_809,N_771,N_658);
or U810 (N_810,N_697,N_701);
xor U811 (N_811,N_753,N_630);
xnor U812 (N_812,N_729,N_690);
and U813 (N_813,N_685,N_672);
or U814 (N_814,N_657,N_779);
xnor U815 (N_815,N_670,N_674);
xnor U816 (N_816,N_791,N_659);
nand U817 (N_817,N_777,N_742);
and U818 (N_818,N_649,N_611);
or U819 (N_819,N_631,N_768);
nand U820 (N_820,N_639,N_712);
xor U821 (N_821,N_636,N_696);
nor U822 (N_822,N_752,N_673);
nand U823 (N_823,N_681,N_754);
nor U824 (N_824,N_734,N_788);
or U825 (N_825,N_775,N_646);
or U826 (N_826,N_786,N_666);
nor U827 (N_827,N_780,N_746);
nor U828 (N_828,N_743,N_660);
xor U829 (N_829,N_747,N_702);
nand U830 (N_830,N_765,N_751);
nand U831 (N_831,N_644,N_615);
or U832 (N_832,N_625,N_614);
and U833 (N_833,N_798,N_653);
nor U834 (N_834,N_667,N_755);
nor U835 (N_835,N_668,N_604);
nand U836 (N_836,N_609,N_643);
xor U837 (N_837,N_610,N_759);
and U838 (N_838,N_774,N_781);
or U839 (N_839,N_637,N_738);
or U840 (N_840,N_632,N_762);
or U841 (N_841,N_664,N_623);
nor U842 (N_842,N_772,N_621);
or U843 (N_843,N_606,N_622);
or U844 (N_844,N_784,N_705);
nand U845 (N_845,N_613,N_703);
and U846 (N_846,N_725,N_642);
nor U847 (N_847,N_654,N_704);
and U848 (N_848,N_723,N_601);
nand U849 (N_849,N_739,N_722);
or U850 (N_850,N_727,N_715);
and U851 (N_851,N_740,N_679);
and U852 (N_852,N_776,N_651);
nor U853 (N_853,N_783,N_677);
nor U854 (N_854,N_635,N_761);
nand U855 (N_855,N_717,N_688);
xnor U856 (N_856,N_633,N_745);
nor U857 (N_857,N_707,N_647);
or U858 (N_858,N_699,N_634);
nand U859 (N_859,N_764,N_665);
or U860 (N_860,N_716,N_767);
or U861 (N_861,N_686,N_794);
xnor U862 (N_862,N_789,N_618);
nand U863 (N_863,N_676,N_769);
nand U864 (N_864,N_682,N_640);
xor U865 (N_865,N_795,N_608);
nor U866 (N_866,N_720,N_726);
and U867 (N_867,N_706,N_612);
and U868 (N_868,N_627,N_652);
or U869 (N_869,N_744,N_782);
nor U870 (N_870,N_790,N_617);
xnor U871 (N_871,N_773,N_709);
nor U872 (N_872,N_711,N_691);
nor U873 (N_873,N_778,N_600);
or U874 (N_874,N_616,N_710);
or U875 (N_875,N_737,N_678);
xor U876 (N_876,N_785,N_624);
nand U877 (N_877,N_607,N_766);
or U878 (N_878,N_713,N_650);
and U879 (N_879,N_756,N_698);
or U880 (N_880,N_645,N_661);
and U881 (N_881,N_602,N_792);
nand U882 (N_882,N_663,N_684);
nor U883 (N_883,N_749,N_714);
and U884 (N_884,N_689,N_799);
or U885 (N_885,N_758,N_669);
and U886 (N_886,N_797,N_735);
nor U887 (N_887,N_724,N_750);
or U888 (N_888,N_796,N_728);
nor U889 (N_889,N_620,N_757);
nor U890 (N_890,N_687,N_732);
nor U891 (N_891,N_736,N_628);
xor U892 (N_892,N_680,N_629);
and U893 (N_893,N_648,N_730);
nor U894 (N_894,N_733,N_655);
or U895 (N_895,N_671,N_693);
xor U896 (N_896,N_748,N_763);
and U897 (N_897,N_692,N_662);
nand U898 (N_898,N_675,N_770);
and U899 (N_899,N_619,N_626);
nand U900 (N_900,N_758,N_685);
or U901 (N_901,N_738,N_791);
nand U902 (N_902,N_650,N_688);
nand U903 (N_903,N_633,N_617);
xnor U904 (N_904,N_740,N_676);
or U905 (N_905,N_630,N_692);
and U906 (N_906,N_760,N_743);
nor U907 (N_907,N_601,N_653);
and U908 (N_908,N_743,N_677);
and U909 (N_909,N_767,N_790);
nor U910 (N_910,N_737,N_697);
or U911 (N_911,N_617,N_622);
nor U912 (N_912,N_773,N_706);
and U913 (N_913,N_745,N_753);
nor U914 (N_914,N_749,N_726);
nand U915 (N_915,N_616,N_663);
nand U916 (N_916,N_642,N_719);
or U917 (N_917,N_790,N_709);
and U918 (N_918,N_655,N_621);
and U919 (N_919,N_792,N_721);
nor U920 (N_920,N_777,N_697);
or U921 (N_921,N_680,N_695);
nand U922 (N_922,N_663,N_627);
and U923 (N_923,N_787,N_799);
nor U924 (N_924,N_709,N_766);
nor U925 (N_925,N_798,N_679);
and U926 (N_926,N_618,N_796);
xor U927 (N_927,N_707,N_747);
nor U928 (N_928,N_742,N_613);
nand U929 (N_929,N_785,N_662);
and U930 (N_930,N_613,N_702);
xnor U931 (N_931,N_624,N_722);
or U932 (N_932,N_713,N_653);
xnor U933 (N_933,N_611,N_601);
or U934 (N_934,N_718,N_670);
nand U935 (N_935,N_608,N_715);
nand U936 (N_936,N_767,N_679);
and U937 (N_937,N_783,N_700);
or U938 (N_938,N_731,N_796);
and U939 (N_939,N_686,N_699);
and U940 (N_940,N_631,N_610);
nor U941 (N_941,N_777,N_635);
or U942 (N_942,N_694,N_740);
nand U943 (N_943,N_709,N_673);
xnor U944 (N_944,N_727,N_631);
and U945 (N_945,N_773,N_669);
or U946 (N_946,N_755,N_764);
nor U947 (N_947,N_777,N_764);
xnor U948 (N_948,N_791,N_644);
xnor U949 (N_949,N_728,N_711);
or U950 (N_950,N_604,N_780);
nor U951 (N_951,N_692,N_781);
nor U952 (N_952,N_738,N_652);
xor U953 (N_953,N_692,N_703);
or U954 (N_954,N_609,N_739);
and U955 (N_955,N_721,N_692);
or U956 (N_956,N_627,N_681);
or U957 (N_957,N_641,N_715);
and U958 (N_958,N_713,N_622);
and U959 (N_959,N_743,N_756);
or U960 (N_960,N_605,N_697);
xor U961 (N_961,N_635,N_703);
nor U962 (N_962,N_723,N_622);
and U963 (N_963,N_707,N_783);
nand U964 (N_964,N_636,N_707);
nor U965 (N_965,N_738,N_610);
or U966 (N_966,N_649,N_749);
nand U967 (N_967,N_773,N_746);
xnor U968 (N_968,N_760,N_718);
nand U969 (N_969,N_770,N_684);
and U970 (N_970,N_623,N_674);
or U971 (N_971,N_652,N_765);
and U972 (N_972,N_738,N_675);
xor U973 (N_973,N_650,N_606);
and U974 (N_974,N_754,N_653);
or U975 (N_975,N_766,N_798);
xor U976 (N_976,N_739,N_626);
or U977 (N_977,N_725,N_784);
and U978 (N_978,N_725,N_781);
nand U979 (N_979,N_618,N_705);
nand U980 (N_980,N_759,N_720);
and U981 (N_981,N_771,N_724);
nand U982 (N_982,N_678,N_771);
xnor U983 (N_983,N_651,N_621);
or U984 (N_984,N_666,N_778);
nand U985 (N_985,N_662,N_699);
nand U986 (N_986,N_795,N_602);
or U987 (N_987,N_790,N_639);
nand U988 (N_988,N_741,N_778);
or U989 (N_989,N_750,N_791);
nand U990 (N_990,N_636,N_601);
xor U991 (N_991,N_658,N_736);
nor U992 (N_992,N_628,N_612);
and U993 (N_993,N_765,N_661);
or U994 (N_994,N_661,N_791);
nand U995 (N_995,N_771,N_615);
and U996 (N_996,N_670,N_628);
or U997 (N_997,N_648,N_741);
or U998 (N_998,N_795,N_639);
or U999 (N_999,N_722,N_707);
or U1000 (N_1000,N_906,N_916);
nor U1001 (N_1001,N_812,N_945);
nor U1002 (N_1002,N_902,N_888);
nand U1003 (N_1003,N_872,N_891);
xnor U1004 (N_1004,N_807,N_814);
or U1005 (N_1005,N_830,N_889);
or U1006 (N_1006,N_824,N_992);
xor U1007 (N_1007,N_986,N_931);
or U1008 (N_1008,N_882,N_983);
nor U1009 (N_1009,N_852,N_972);
or U1010 (N_1010,N_897,N_835);
nor U1011 (N_1011,N_991,N_933);
nor U1012 (N_1012,N_808,N_841);
nand U1013 (N_1013,N_976,N_903);
nor U1014 (N_1014,N_927,N_925);
nand U1015 (N_1015,N_887,N_947);
nand U1016 (N_1016,N_923,N_855);
nand U1017 (N_1017,N_910,N_833);
nand U1018 (N_1018,N_871,N_909);
nand U1019 (N_1019,N_998,N_846);
and U1020 (N_1020,N_896,N_858);
or U1021 (N_1021,N_985,N_980);
nand U1022 (N_1022,N_955,N_938);
or U1023 (N_1023,N_936,N_918);
or U1024 (N_1024,N_930,N_861);
or U1025 (N_1025,N_898,N_911);
and U1026 (N_1026,N_907,N_827);
or U1027 (N_1027,N_951,N_883);
nand U1028 (N_1028,N_966,N_843);
or U1029 (N_1029,N_993,N_820);
nand U1030 (N_1030,N_953,N_996);
or U1031 (N_1031,N_847,N_869);
and U1032 (N_1032,N_881,N_971);
or U1033 (N_1033,N_978,N_973);
xor U1034 (N_1034,N_950,N_832);
nand U1035 (N_1035,N_990,N_844);
nand U1036 (N_1036,N_863,N_817);
xnor U1037 (N_1037,N_974,N_922);
nand U1038 (N_1038,N_942,N_944);
and U1039 (N_1039,N_956,N_940);
nor U1040 (N_1040,N_860,N_994);
nor U1041 (N_1041,N_811,N_997);
nand U1042 (N_1042,N_849,N_919);
or U1043 (N_1043,N_874,N_873);
nand U1044 (N_1044,N_970,N_865);
and U1045 (N_1045,N_999,N_831);
and U1046 (N_1046,N_886,N_959);
and U1047 (N_1047,N_920,N_929);
xnor U1048 (N_1048,N_821,N_939);
nand U1049 (N_1049,N_908,N_984);
nor U1050 (N_1050,N_805,N_982);
xor U1051 (N_1051,N_880,N_957);
xor U1052 (N_1052,N_870,N_859);
nand U1053 (N_1053,N_937,N_822);
or U1054 (N_1054,N_829,N_815);
nor U1055 (N_1055,N_879,N_924);
nand U1056 (N_1056,N_813,N_946);
nand U1057 (N_1057,N_948,N_845);
xor U1058 (N_1058,N_857,N_884);
nor U1059 (N_1059,N_894,N_932);
and U1060 (N_1060,N_875,N_967);
nand U1061 (N_1061,N_941,N_803);
xor U1062 (N_1062,N_912,N_850);
and U1063 (N_1063,N_962,N_893);
xnor U1064 (N_1064,N_935,N_809);
or U1065 (N_1065,N_988,N_826);
or U1066 (N_1066,N_837,N_917);
or U1067 (N_1067,N_904,N_801);
nor U1068 (N_1068,N_842,N_840);
and U1069 (N_1069,N_878,N_943);
nand U1070 (N_1070,N_800,N_915);
nand U1071 (N_1071,N_928,N_804);
nor U1072 (N_1072,N_949,N_851);
nand U1073 (N_1073,N_877,N_828);
or U1074 (N_1074,N_995,N_862);
or U1075 (N_1075,N_979,N_838);
nor U1076 (N_1076,N_839,N_934);
nand U1077 (N_1077,N_987,N_866);
and U1078 (N_1078,N_914,N_892);
and U1079 (N_1079,N_864,N_834);
and U1080 (N_1080,N_868,N_876);
nand U1081 (N_1081,N_964,N_913);
or U1082 (N_1082,N_818,N_954);
nor U1083 (N_1083,N_853,N_989);
and U1084 (N_1084,N_825,N_836);
nand U1085 (N_1085,N_885,N_975);
xor U1086 (N_1086,N_819,N_968);
or U1087 (N_1087,N_981,N_952);
nand U1088 (N_1088,N_901,N_921);
nand U1089 (N_1089,N_900,N_905);
nand U1090 (N_1090,N_963,N_977);
or U1091 (N_1091,N_848,N_961);
nand U1092 (N_1092,N_895,N_810);
nand U1093 (N_1093,N_969,N_802);
xor U1094 (N_1094,N_823,N_867);
or U1095 (N_1095,N_965,N_899);
or U1096 (N_1096,N_960,N_816);
and U1097 (N_1097,N_806,N_854);
nor U1098 (N_1098,N_926,N_890);
and U1099 (N_1099,N_958,N_856);
nor U1100 (N_1100,N_912,N_978);
nand U1101 (N_1101,N_946,N_862);
or U1102 (N_1102,N_818,N_879);
or U1103 (N_1103,N_937,N_904);
nand U1104 (N_1104,N_926,N_900);
and U1105 (N_1105,N_945,N_822);
nand U1106 (N_1106,N_952,N_930);
nor U1107 (N_1107,N_945,N_836);
nor U1108 (N_1108,N_860,N_935);
nor U1109 (N_1109,N_990,N_874);
xor U1110 (N_1110,N_993,N_877);
or U1111 (N_1111,N_988,N_867);
or U1112 (N_1112,N_803,N_963);
and U1113 (N_1113,N_957,N_973);
or U1114 (N_1114,N_913,N_988);
xnor U1115 (N_1115,N_982,N_925);
nor U1116 (N_1116,N_848,N_924);
nor U1117 (N_1117,N_825,N_925);
and U1118 (N_1118,N_992,N_907);
xnor U1119 (N_1119,N_950,N_869);
and U1120 (N_1120,N_820,N_804);
or U1121 (N_1121,N_805,N_842);
and U1122 (N_1122,N_856,N_891);
nor U1123 (N_1123,N_865,N_895);
nand U1124 (N_1124,N_968,N_900);
and U1125 (N_1125,N_876,N_990);
nand U1126 (N_1126,N_864,N_880);
xor U1127 (N_1127,N_813,N_901);
and U1128 (N_1128,N_864,N_921);
nor U1129 (N_1129,N_842,N_822);
nor U1130 (N_1130,N_984,N_827);
and U1131 (N_1131,N_839,N_800);
nand U1132 (N_1132,N_871,N_961);
nand U1133 (N_1133,N_877,N_974);
nand U1134 (N_1134,N_867,N_977);
and U1135 (N_1135,N_852,N_891);
and U1136 (N_1136,N_808,N_818);
nor U1137 (N_1137,N_982,N_931);
nand U1138 (N_1138,N_966,N_940);
nand U1139 (N_1139,N_827,N_982);
or U1140 (N_1140,N_868,N_935);
nor U1141 (N_1141,N_840,N_834);
or U1142 (N_1142,N_854,N_916);
or U1143 (N_1143,N_886,N_988);
or U1144 (N_1144,N_889,N_872);
or U1145 (N_1145,N_998,N_977);
nand U1146 (N_1146,N_966,N_938);
and U1147 (N_1147,N_874,N_850);
nand U1148 (N_1148,N_814,N_852);
and U1149 (N_1149,N_911,N_813);
xnor U1150 (N_1150,N_940,N_943);
nand U1151 (N_1151,N_877,N_858);
xnor U1152 (N_1152,N_870,N_844);
and U1153 (N_1153,N_893,N_878);
or U1154 (N_1154,N_854,N_835);
nor U1155 (N_1155,N_971,N_818);
or U1156 (N_1156,N_969,N_824);
or U1157 (N_1157,N_907,N_813);
or U1158 (N_1158,N_854,N_857);
nand U1159 (N_1159,N_911,N_996);
nand U1160 (N_1160,N_812,N_828);
nand U1161 (N_1161,N_895,N_923);
and U1162 (N_1162,N_920,N_948);
or U1163 (N_1163,N_876,N_995);
nand U1164 (N_1164,N_922,N_878);
or U1165 (N_1165,N_904,N_805);
nor U1166 (N_1166,N_998,N_868);
and U1167 (N_1167,N_876,N_833);
or U1168 (N_1168,N_896,N_819);
or U1169 (N_1169,N_979,N_881);
nor U1170 (N_1170,N_807,N_928);
and U1171 (N_1171,N_972,N_947);
nand U1172 (N_1172,N_863,N_990);
or U1173 (N_1173,N_850,N_839);
nand U1174 (N_1174,N_937,N_906);
nor U1175 (N_1175,N_808,N_852);
nor U1176 (N_1176,N_844,N_824);
nor U1177 (N_1177,N_910,N_848);
nor U1178 (N_1178,N_831,N_865);
nor U1179 (N_1179,N_959,N_850);
xor U1180 (N_1180,N_827,N_854);
and U1181 (N_1181,N_972,N_901);
or U1182 (N_1182,N_896,N_937);
nand U1183 (N_1183,N_996,N_958);
xor U1184 (N_1184,N_937,N_953);
nand U1185 (N_1185,N_864,N_853);
nand U1186 (N_1186,N_898,N_998);
and U1187 (N_1187,N_960,N_880);
or U1188 (N_1188,N_899,N_972);
and U1189 (N_1189,N_929,N_967);
and U1190 (N_1190,N_846,N_925);
or U1191 (N_1191,N_903,N_812);
or U1192 (N_1192,N_894,N_983);
xnor U1193 (N_1193,N_877,N_838);
or U1194 (N_1194,N_812,N_961);
nand U1195 (N_1195,N_840,N_816);
nand U1196 (N_1196,N_826,N_866);
and U1197 (N_1197,N_984,N_863);
nand U1198 (N_1198,N_963,N_997);
xnor U1199 (N_1199,N_854,N_943);
nor U1200 (N_1200,N_1060,N_1121);
xnor U1201 (N_1201,N_1164,N_1078);
or U1202 (N_1202,N_1128,N_1014);
and U1203 (N_1203,N_1165,N_1080);
nor U1204 (N_1204,N_1067,N_1033);
nor U1205 (N_1205,N_1030,N_1048);
xor U1206 (N_1206,N_1143,N_1058);
and U1207 (N_1207,N_1189,N_1049);
xnor U1208 (N_1208,N_1101,N_1056);
nor U1209 (N_1209,N_1126,N_1004);
nor U1210 (N_1210,N_1179,N_1027);
and U1211 (N_1211,N_1031,N_1083);
and U1212 (N_1212,N_1180,N_1136);
nand U1213 (N_1213,N_1148,N_1187);
nor U1214 (N_1214,N_1061,N_1175);
and U1215 (N_1215,N_1108,N_1013);
nand U1216 (N_1216,N_1157,N_1096);
or U1217 (N_1217,N_1050,N_1020);
or U1218 (N_1218,N_1043,N_1012);
nor U1219 (N_1219,N_1059,N_1035);
nor U1220 (N_1220,N_1029,N_1094);
nor U1221 (N_1221,N_1086,N_1079);
nor U1222 (N_1222,N_1181,N_1168);
xor U1223 (N_1223,N_1045,N_1199);
or U1224 (N_1224,N_1127,N_1010);
xnor U1225 (N_1225,N_1169,N_1171);
and U1226 (N_1226,N_1075,N_1006);
or U1227 (N_1227,N_1142,N_1021);
nand U1228 (N_1228,N_1093,N_1115);
nand U1229 (N_1229,N_1134,N_1024);
xnor U1230 (N_1230,N_1019,N_1182);
nand U1231 (N_1231,N_1087,N_1112);
nor U1232 (N_1232,N_1170,N_1039);
and U1233 (N_1233,N_1002,N_1173);
or U1234 (N_1234,N_1057,N_1100);
nand U1235 (N_1235,N_1119,N_1018);
or U1236 (N_1236,N_1135,N_1007);
or U1237 (N_1237,N_1026,N_1129);
nor U1238 (N_1238,N_1118,N_1076);
xnor U1239 (N_1239,N_1036,N_1001);
nand U1240 (N_1240,N_1023,N_1124);
or U1241 (N_1241,N_1074,N_1120);
nor U1242 (N_1242,N_1161,N_1032);
or U1243 (N_1243,N_1196,N_1028);
nor U1244 (N_1244,N_1069,N_1103);
or U1245 (N_1245,N_1085,N_1177);
and U1246 (N_1246,N_1047,N_1153);
nand U1247 (N_1247,N_1197,N_1042);
and U1248 (N_1248,N_1186,N_1138);
or U1249 (N_1249,N_1194,N_1107);
xor U1250 (N_1250,N_1110,N_1117);
and U1251 (N_1251,N_1088,N_1044);
and U1252 (N_1252,N_1077,N_1071);
nand U1253 (N_1253,N_1151,N_1152);
or U1254 (N_1254,N_1091,N_1102);
or U1255 (N_1255,N_1131,N_1188);
or U1256 (N_1256,N_1166,N_1106);
xor U1257 (N_1257,N_1193,N_1015);
or U1258 (N_1258,N_1178,N_1065);
nand U1259 (N_1259,N_1053,N_1174);
and U1260 (N_1260,N_1062,N_1114);
nor U1261 (N_1261,N_1192,N_1072);
or U1262 (N_1262,N_1038,N_1104);
nand U1263 (N_1263,N_1172,N_1090);
nor U1264 (N_1264,N_1154,N_1167);
and U1265 (N_1265,N_1054,N_1016);
and U1266 (N_1266,N_1063,N_1022);
or U1267 (N_1267,N_1105,N_1125);
nand U1268 (N_1268,N_1040,N_1095);
nand U1269 (N_1269,N_1109,N_1132);
nand U1270 (N_1270,N_1025,N_1159);
and U1271 (N_1271,N_1017,N_1082);
and U1272 (N_1272,N_1160,N_1011);
or U1273 (N_1273,N_1113,N_1155);
or U1274 (N_1274,N_1111,N_1066);
nor U1275 (N_1275,N_1084,N_1009);
xor U1276 (N_1276,N_1191,N_1185);
and U1277 (N_1277,N_1092,N_1046);
nand U1278 (N_1278,N_1099,N_1176);
and U1279 (N_1279,N_1116,N_1034);
or U1280 (N_1280,N_1140,N_1183);
xnor U1281 (N_1281,N_1073,N_1144);
or U1282 (N_1282,N_1005,N_1149);
nor U1283 (N_1283,N_1123,N_1008);
xnor U1284 (N_1284,N_1139,N_1137);
and U1285 (N_1285,N_1098,N_1051);
nand U1286 (N_1286,N_1037,N_1156);
nor U1287 (N_1287,N_1146,N_1122);
or U1288 (N_1288,N_1003,N_1198);
nor U1289 (N_1289,N_1064,N_1163);
and U1290 (N_1290,N_1147,N_1130);
or U1291 (N_1291,N_1158,N_1089);
nor U1292 (N_1292,N_1150,N_1190);
nor U1293 (N_1293,N_1162,N_1133);
nand U1294 (N_1294,N_1052,N_1070);
xor U1295 (N_1295,N_1041,N_1195);
nand U1296 (N_1296,N_1068,N_1081);
and U1297 (N_1297,N_1141,N_1184);
or U1298 (N_1298,N_1000,N_1097);
nand U1299 (N_1299,N_1145,N_1055);
nand U1300 (N_1300,N_1004,N_1096);
and U1301 (N_1301,N_1173,N_1008);
nor U1302 (N_1302,N_1171,N_1088);
nand U1303 (N_1303,N_1150,N_1088);
xor U1304 (N_1304,N_1175,N_1035);
or U1305 (N_1305,N_1017,N_1141);
nor U1306 (N_1306,N_1082,N_1006);
nand U1307 (N_1307,N_1049,N_1027);
xor U1308 (N_1308,N_1192,N_1143);
xnor U1309 (N_1309,N_1150,N_1021);
nor U1310 (N_1310,N_1156,N_1196);
nand U1311 (N_1311,N_1172,N_1063);
nor U1312 (N_1312,N_1037,N_1157);
nand U1313 (N_1313,N_1002,N_1028);
or U1314 (N_1314,N_1044,N_1030);
nor U1315 (N_1315,N_1031,N_1126);
nor U1316 (N_1316,N_1152,N_1103);
nor U1317 (N_1317,N_1151,N_1191);
nor U1318 (N_1318,N_1045,N_1096);
nor U1319 (N_1319,N_1014,N_1028);
and U1320 (N_1320,N_1176,N_1134);
and U1321 (N_1321,N_1037,N_1052);
or U1322 (N_1322,N_1180,N_1017);
or U1323 (N_1323,N_1073,N_1068);
and U1324 (N_1324,N_1002,N_1192);
or U1325 (N_1325,N_1003,N_1113);
and U1326 (N_1326,N_1079,N_1032);
nor U1327 (N_1327,N_1073,N_1140);
and U1328 (N_1328,N_1188,N_1032);
and U1329 (N_1329,N_1181,N_1065);
or U1330 (N_1330,N_1107,N_1034);
nor U1331 (N_1331,N_1030,N_1197);
nand U1332 (N_1332,N_1104,N_1094);
xnor U1333 (N_1333,N_1104,N_1067);
nand U1334 (N_1334,N_1098,N_1058);
and U1335 (N_1335,N_1001,N_1163);
or U1336 (N_1336,N_1132,N_1162);
nand U1337 (N_1337,N_1129,N_1121);
or U1338 (N_1338,N_1192,N_1050);
and U1339 (N_1339,N_1183,N_1086);
nand U1340 (N_1340,N_1172,N_1087);
nor U1341 (N_1341,N_1113,N_1106);
and U1342 (N_1342,N_1042,N_1179);
nand U1343 (N_1343,N_1079,N_1199);
xnor U1344 (N_1344,N_1092,N_1133);
nor U1345 (N_1345,N_1077,N_1117);
xnor U1346 (N_1346,N_1014,N_1094);
and U1347 (N_1347,N_1186,N_1100);
nor U1348 (N_1348,N_1090,N_1135);
nand U1349 (N_1349,N_1191,N_1012);
nand U1350 (N_1350,N_1016,N_1160);
xor U1351 (N_1351,N_1110,N_1175);
or U1352 (N_1352,N_1103,N_1051);
xnor U1353 (N_1353,N_1165,N_1052);
or U1354 (N_1354,N_1188,N_1067);
nor U1355 (N_1355,N_1104,N_1016);
xor U1356 (N_1356,N_1161,N_1192);
nand U1357 (N_1357,N_1143,N_1098);
xor U1358 (N_1358,N_1061,N_1164);
and U1359 (N_1359,N_1038,N_1084);
nand U1360 (N_1360,N_1046,N_1076);
and U1361 (N_1361,N_1088,N_1055);
or U1362 (N_1362,N_1197,N_1171);
nor U1363 (N_1363,N_1146,N_1148);
nor U1364 (N_1364,N_1058,N_1189);
nand U1365 (N_1365,N_1192,N_1066);
and U1366 (N_1366,N_1089,N_1036);
xor U1367 (N_1367,N_1048,N_1060);
nor U1368 (N_1368,N_1130,N_1075);
and U1369 (N_1369,N_1094,N_1187);
and U1370 (N_1370,N_1070,N_1059);
nor U1371 (N_1371,N_1124,N_1145);
nand U1372 (N_1372,N_1123,N_1035);
nor U1373 (N_1373,N_1122,N_1155);
nor U1374 (N_1374,N_1141,N_1149);
or U1375 (N_1375,N_1076,N_1068);
nand U1376 (N_1376,N_1093,N_1040);
nor U1377 (N_1377,N_1147,N_1191);
nor U1378 (N_1378,N_1061,N_1145);
nand U1379 (N_1379,N_1086,N_1182);
nand U1380 (N_1380,N_1098,N_1044);
nand U1381 (N_1381,N_1015,N_1108);
xnor U1382 (N_1382,N_1044,N_1148);
and U1383 (N_1383,N_1056,N_1150);
nand U1384 (N_1384,N_1174,N_1176);
nor U1385 (N_1385,N_1060,N_1176);
or U1386 (N_1386,N_1076,N_1007);
nand U1387 (N_1387,N_1120,N_1098);
nand U1388 (N_1388,N_1073,N_1087);
or U1389 (N_1389,N_1185,N_1112);
nand U1390 (N_1390,N_1169,N_1070);
nor U1391 (N_1391,N_1007,N_1115);
xor U1392 (N_1392,N_1194,N_1038);
nand U1393 (N_1393,N_1187,N_1037);
nand U1394 (N_1394,N_1080,N_1043);
or U1395 (N_1395,N_1094,N_1095);
nor U1396 (N_1396,N_1056,N_1152);
xor U1397 (N_1397,N_1018,N_1031);
nor U1398 (N_1398,N_1094,N_1049);
xor U1399 (N_1399,N_1113,N_1012);
nor U1400 (N_1400,N_1206,N_1313);
and U1401 (N_1401,N_1221,N_1388);
and U1402 (N_1402,N_1330,N_1291);
and U1403 (N_1403,N_1215,N_1391);
or U1404 (N_1404,N_1256,N_1398);
nand U1405 (N_1405,N_1254,N_1369);
and U1406 (N_1406,N_1340,N_1351);
nor U1407 (N_1407,N_1207,N_1362);
or U1408 (N_1408,N_1203,N_1249);
nand U1409 (N_1409,N_1309,N_1368);
xor U1410 (N_1410,N_1218,N_1304);
and U1411 (N_1411,N_1287,N_1255);
nand U1412 (N_1412,N_1245,N_1342);
and U1413 (N_1413,N_1293,N_1297);
or U1414 (N_1414,N_1325,N_1341);
or U1415 (N_1415,N_1259,N_1360);
nand U1416 (N_1416,N_1200,N_1314);
and U1417 (N_1417,N_1209,N_1367);
or U1418 (N_1418,N_1366,N_1295);
and U1419 (N_1419,N_1361,N_1364);
nand U1420 (N_1420,N_1386,N_1260);
nand U1421 (N_1421,N_1339,N_1228);
nand U1422 (N_1422,N_1357,N_1355);
or U1423 (N_1423,N_1322,N_1269);
nor U1424 (N_1424,N_1212,N_1305);
nor U1425 (N_1425,N_1288,N_1264);
and U1426 (N_1426,N_1374,N_1237);
or U1427 (N_1427,N_1270,N_1382);
nand U1428 (N_1428,N_1292,N_1343);
and U1429 (N_1429,N_1267,N_1277);
nand U1430 (N_1430,N_1332,N_1290);
or U1431 (N_1431,N_1281,N_1217);
xnor U1432 (N_1432,N_1222,N_1211);
nand U1433 (N_1433,N_1282,N_1253);
nand U1434 (N_1434,N_1216,N_1328);
or U1435 (N_1435,N_1225,N_1334);
or U1436 (N_1436,N_1394,N_1315);
and U1437 (N_1437,N_1296,N_1335);
nor U1438 (N_1438,N_1306,N_1311);
nor U1439 (N_1439,N_1376,N_1385);
nand U1440 (N_1440,N_1219,N_1380);
or U1441 (N_1441,N_1379,N_1327);
and U1442 (N_1442,N_1383,N_1223);
nor U1443 (N_1443,N_1389,N_1248);
or U1444 (N_1444,N_1384,N_1210);
and U1445 (N_1445,N_1354,N_1301);
and U1446 (N_1446,N_1375,N_1370);
and U1447 (N_1447,N_1214,N_1331);
nand U1448 (N_1448,N_1299,N_1284);
nor U1449 (N_1449,N_1393,N_1224);
nand U1450 (N_1450,N_1300,N_1319);
nand U1451 (N_1451,N_1220,N_1344);
nand U1452 (N_1452,N_1234,N_1258);
and U1453 (N_1453,N_1387,N_1246);
or U1454 (N_1454,N_1227,N_1347);
or U1455 (N_1455,N_1232,N_1353);
nor U1456 (N_1456,N_1392,N_1337);
or U1457 (N_1457,N_1205,N_1352);
nand U1458 (N_1458,N_1266,N_1338);
xnor U1459 (N_1459,N_1323,N_1202);
or U1460 (N_1460,N_1321,N_1312);
and U1461 (N_1461,N_1250,N_1286);
nor U1462 (N_1462,N_1348,N_1244);
and U1463 (N_1463,N_1371,N_1276);
and U1464 (N_1464,N_1397,N_1233);
or U1465 (N_1465,N_1308,N_1285);
and U1466 (N_1466,N_1372,N_1350);
nor U1467 (N_1467,N_1365,N_1229);
or U1468 (N_1468,N_1345,N_1204);
nand U1469 (N_1469,N_1395,N_1236);
and U1470 (N_1470,N_1257,N_1302);
nor U1471 (N_1471,N_1377,N_1231);
nor U1472 (N_1472,N_1378,N_1275);
or U1473 (N_1473,N_1346,N_1310);
or U1474 (N_1474,N_1271,N_1226);
nor U1475 (N_1475,N_1268,N_1213);
and U1476 (N_1476,N_1278,N_1320);
nor U1477 (N_1477,N_1363,N_1356);
and U1478 (N_1478,N_1242,N_1241);
and U1479 (N_1479,N_1243,N_1294);
nand U1480 (N_1480,N_1263,N_1283);
and U1481 (N_1481,N_1262,N_1230);
or U1482 (N_1482,N_1317,N_1251);
nor U1483 (N_1483,N_1349,N_1316);
or U1484 (N_1484,N_1324,N_1238);
nand U1485 (N_1485,N_1247,N_1318);
nand U1486 (N_1486,N_1274,N_1235);
and U1487 (N_1487,N_1307,N_1298);
or U1488 (N_1488,N_1381,N_1280);
nand U1489 (N_1489,N_1279,N_1201);
nand U1490 (N_1490,N_1396,N_1359);
nand U1491 (N_1491,N_1265,N_1272);
and U1492 (N_1492,N_1303,N_1333);
or U1493 (N_1493,N_1326,N_1273);
or U1494 (N_1494,N_1261,N_1240);
or U1495 (N_1495,N_1208,N_1289);
nand U1496 (N_1496,N_1358,N_1336);
xnor U1497 (N_1497,N_1399,N_1329);
and U1498 (N_1498,N_1252,N_1390);
nand U1499 (N_1499,N_1373,N_1239);
or U1500 (N_1500,N_1303,N_1241);
xor U1501 (N_1501,N_1342,N_1224);
or U1502 (N_1502,N_1236,N_1264);
nor U1503 (N_1503,N_1226,N_1349);
or U1504 (N_1504,N_1371,N_1226);
nand U1505 (N_1505,N_1358,N_1290);
and U1506 (N_1506,N_1366,N_1262);
nor U1507 (N_1507,N_1341,N_1236);
or U1508 (N_1508,N_1301,N_1242);
nand U1509 (N_1509,N_1330,N_1385);
or U1510 (N_1510,N_1334,N_1388);
nor U1511 (N_1511,N_1319,N_1339);
or U1512 (N_1512,N_1214,N_1202);
or U1513 (N_1513,N_1377,N_1241);
xor U1514 (N_1514,N_1255,N_1322);
or U1515 (N_1515,N_1226,N_1381);
or U1516 (N_1516,N_1379,N_1309);
nor U1517 (N_1517,N_1315,N_1258);
nor U1518 (N_1518,N_1368,N_1201);
nor U1519 (N_1519,N_1202,N_1379);
nor U1520 (N_1520,N_1355,N_1318);
or U1521 (N_1521,N_1348,N_1353);
nor U1522 (N_1522,N_1317,N_1356);
nor U1523 (N_1523,N_1311,N_1210);
nor U1524 (N_1524,N_1351,N_1335);
nand U1525 (N_1525,N_1250,N_1222);
or U1526 (N_1526,N_1207,N_1204);
and U1527 (N_1527,N_1226,N_1322);
nor U1528 (N_1528,N_1251,N_1326);
nor U1529 (N_1529,N_1345,N_1340);
nor U1530 (N_1530,N_1304,N_1278);
nand U1531 (N_1531,N_1396,N_1284);
nor U1532 (N_1532,N_1323,N_1332);
nor U1533 (N_1533,N_1343,N_1282);
or U1534 (N_1534,N_1376,N_1291);
nand U1535 (N_1535,N_1330,N_1246);
and U1536 (N_1536,N_1220,N_1396);
nand U1537 (N_1537,N_1274,N_1205);
nor U1538 (N_1538,N_1371,N_1301);
nand U1539 (N_1539,N_1354,N_1267);
nor U1540 (N_1540,N_1370,N_1289);
nand U1541 (N_1541,N_1399,N_1327);
nand U1542 (N_1542,N_1280,N_1363);
or U1543 (N_1543,N_1367,N_1345);
and U1544 (N_1544,N_1271,N_1241);
nand U1545 (N_1545,N_1215,N_1300);
or U1546 (N_1546,N_1309,N_1267);
nand U1547 (N_1547,N_1217,N_1299);
xnor U1548 (N_1548,N_1331,N_1309);
xor U1549 (N_1549,N_1277,N_1309);
nor U1550 (N_1550,N_1213,N_1308);
and U1551 (N_1551,N_1352,N_1207);
nor U1552 (N_1552,N_1338,N_1203);
nor U1553 (N_1553,N_1352,N_1291);
nand U1554 (N_1554,N_1382,N_1378);
nor U1555 (N_1555,N_1338,N_1299);
nand U1556 (N_1556,N_1208,N_1246);
xor U1557 (N_1557,N_1306,N_1264);
nor U1558 (N_1558,N_1371,N_1225);
nand U1559 (N_1559,N_1341,N_1229);
xnor U1560 (N_1560,N_1367,N_1221);
nand U1561 (N_1561,N_1325,N_1383);
nand U1562 (N_1562,N_1274,N_1320);
nor U1563 (N_1563,N_1330,N_1387);
or U1564 (N_1564,N_1294,N_1339);
xor U1565 (N_1565,N_1309,N_1282);
nor U1566 (N_1566,N_1353,N_1345);
and U1567 (N_1567,N_1236,N_1271);
nand U1568 (N_1568,N_1315,N_1266);
nor U1569 (N_1569,N_1359,N_1265);
nand U1570 (N_1570,N_1374,N_1372);
nor U1571 (N_1571,N_1246,N_1328);
and U1572 (N_1572,N_1228,N_1246);
nand U1573 (N_1573,N_1284,N_1231);
nand U1574 (N_1574,N_1242,N_1268);
nand U1575 (N_1575,N_1394,N_1393);
or U1576 (N_1576,N_1274,N_1322);
or U1577 (N_1577,N_1263,N_1281);
and U1578 (N_1578,N_1358,N_1211);
nand U1579 (N_1579,N_1293,N_1305);
or U1580 (N_1580,N_1377,N_1238);
nand U1581 (N_1581,N_1358,N_1372);
nor U1582 (N_1582,N_1281,N_1379);
nand U1583 (N_1583,N_1356,N_1286);
and U1584 (N_1584,N_1345,N_1228);
and U1585 (N_1585,N_1337,N_1330);
nand U1586 (N_1586,N_1288,N_1226);
nand U1587 (N_1587,N_1340,N_1276);
nand U1588 (N_1588,N_1208,N_1397);
nand U1589 (N_1589,N_1224,N_1332);
and U1590 (N_1590,N_1270,N_1241);
xor U1591 (N_1591,N_1376,N_1349);
nand U1592 (N_1592,N_1247,N_1289);
nor U1593 (N_1593,N_1392,N_1320);
nor U1594 (N_1594,N_1278,N_1318);
nand U1595 (N_1595,N_1260,N_1289);
nand U1596 (N_1596,N_1345,N_1311);
and U1597 (N_1597,N_1220,N_1200);
nor U1598 (N_1598,N_1355,N_1251);
nand U1599 (N_1599,N_1230,N_1345);
nor U1600 (N_1600,N_1477,N_1564);
and U1601 (N_1601,N_1434,N_1519);
nand U1602 (N_1602,N_1472,N_1460);
xnor U1603 (N_1603,N_1567,N_1500);
nand U1604 (N_1604,N_1508,N_1407);
and U1605 (N_1605,N_1510,N_1503);
nor U1606 (N_1606,N_1416,N_1509);
nor U1607 (N_1607,N_1490,N_1478);
and U1608 (N_1608,N_1512,N_1532);
nor U1609 (N_1609,N_1431,N_1496);
nand U1610 (N_1610,N_1482,N_1438);
nand U1611 (N_1611,N_1565,N_1597);
nor U1612 (N_1612,N_1479,N_1572);
and U1613 (N_1613,N_1468,N_1596);
and U1614 (N_1614,N_1495,N_1497);
nor U1615 (N_1615,N_1439,N_1586);
and U1616 (N_1616,N_1540,N_1591);
and U1617 (N_1617,N_1590,N_1421);
nand U1618 (N_1618,N_1518,N_1547);
nand U1619 (N_1619,N_1530,N_1568);
nor U1620 (N_1620,N_1437,N_1528);
nand U1621 (N_1621,N_1511,N_1463);
xor U1622 (N_1622,N_1459,N_1442);
xnor U1623 (N_1623,N_1505,N_1577);
nor U1624 (N_1624,N_1402,N_1550);
nand U1625 (N_1625,N_1556,N_1413);
xnor U1626 (N_1626,N_1525,N_1487);
nand U1627 (N_1627,N_1446,N_1592);
and U1628 (N_1628,N_1598,N_1444);
nor U1629 (N_1629,N_1435,N_1406);
and U1630 (N_1630,N_1553,N_1411);
or U1631 (N_1631,N_1539,N_1589);
or U1632 (N_1632,N_1515,N_1533);
nand U1633 (N_1633,N_1448,N_1581);
nor U1634 (N_1634,N_1410,N_1473);
nand U1635 (N_1635,N_1569,N_1428);
xor U1636 (N_1636,N_1543,N_1425);
and U1637 (N_1637,N_1401,N_1422);
and U1638 (N_1638,N_1430,N_1455);
and U1639 (N_1639,N_1418,N_1563);
xor U1640 (N_1640,N_1475,N_1464);
or U1641 (N_1641,N_1560,N_1474);
nand U1642 (N_1642,N_1485,N_1587);
nor U1643 (N_1643,N_1492,N_1514);
nand U1644 (N_1644,N_1593,N_1449);
or U1645 (N_1645,N_1458,N_1441);
and U1646 (N_1646,N_1538,N_1555);
and U1647 (N_1647,N_1578,N_1486);
nor U1648 (N_1648,N_1452,N_1494);
or U1649 (N_1649,N_1404,N_1480);
and U1650 (N_1650,N_1462,N_1520);
or U1651 (N_1651,N_1419,N_1417);
nor U1652 (N_1652,N_1470,N_1599);
nand U1653 (N_1653,N_1522,N_1546);
nand U1654 (N_1654,N_1541,N_1551);
nand U1655 (N_1655,N_1471,N_1595);
nand U1656 (N_1656,N_1573,N_1554);
or U1657 (N_1657,N_1420,N_1423);
or U1658 (N_1658,N_1445,N_1493);
nor U1659 (N_1659,N_1488,N_1580);
nand U1660 (N_1660,N_1409,N_1524);
and U1661 (N_1661,N_1469,N_1466);
and U1662 (N_1662,N_1467,N_1570);
and U1663 (N_1663,N_1408,N_1403);
or U1664 (N_1664,N_1481,N_1517);
or U1665 (N_1665,N_1535,N_1484);
nor U1666 (N_1666,N_1531,N_1558);
nor U1667 (N_1667,N_1451,N_1414);
or U1668 (N_1668,N_1527,N_1594);
or U1669 (N_1669,N_1521,N_1454);
nor U1670 (N_1670,N_1584,N_1545);
xor U1671 (N_1671,N_1523,N_1499);
nand U1672 (N_1672,N_1534,N_1548);
and U1673 (N_1673,N_1429,N_1415);
and U1674 (N_1674,N_1440,N_1461);
or U1675 (N_1675,N_1582,N_1537);
or U1676 (N_1676,N_1507,N_1427);
nor U1677 (N_1677,N_1566,N_1552);
nand U1678 (N_1678,N_1529,N_1588);
nand U1679 (N_1679,N_1433,N_1504);
or U1680 (N_1680,N_1557,N_1502);
nor U1681 (N_1681,N_1457,N_1456);
or U1682 (N_1682,N_1574,N_1447);
or U1683 (N_1683,N_1405,N_1542);
nand U1684 (N_1684,N_1465,N_1506);
nand U1685 (N_1685,N_1585,N_1501);
and U1686 (N_1686,N_1571,N_1576);
nand U1687 (N_1687,N_1536,N_1424);
nand U1688 (N_1688,N_1559,N_1544);
nor U1689 (N_1689,N_1498,N_1426);
nor U1690 (N_1690,N_1483,N_1575);
nand U1691 (N_1691,N_1476,N_1561);
and U1692 (N_1692,N_1562,N_1583);
nor U1693 (N_1693,N_1436,N_1516);
and U1694 (N_1694,N_1489,N_1579);
nor U1695 (N_1695,N_1526,N_1400);
or U1696 (N_1696,N_1450,N_1491);
nor U1697 (N_1697,N_1443,N_1513);
or U1698 (N_1698,N_1549,N_1453);
or U1699 (N_1699,N_1412,N_1432);
and U1700 (N_1700,N_1540,N_1555);
nor U1701 (N_1701,N_1563,N_1436);
and U1702 (N_1702,N_1536,N_1527);
or U1703 (N_1703,N_1575,N_1478);
and U1704 (N_1704,N_1571,N_1444);
nor U1705 (N_1705,N_1590,N_1448);
or U1706 (N_1706,N_1518,N_1517);
nand U1707 (N_1707,N_1469,N_1412);
and U1708 (N_1708,N_1483,N_1527);
nand U1709 (N_1709,N_1423,N_1561);
and U1710 (N_1710,N_1491,N_1571);
and U1711 (N_1711,N_1491,N_1411);
nor U1712 (N_1712,N_1556,N_1417);
and U1713 (N_1713,N_1475,N_1588);
nor U1714 (N_1714,N_1424,N_1555);
or U1715 (N_1715,N_1447,N_1579);
and U1716 (N_1716,N_1544,N_1531);
and U1717 (N_1717,N_1441,N_1566);
nor U1718 (N_1718,N_1484,N_1540);
xor U1719 (N_1719,N_1429,N_1419);
and U1720 (N_1720,N_1513,N_1595);
xor U1721 (N_1721,N_1433,N_1488);
nand U1722 (N_1722,N_1482,N_1409);
xor U1723 (N_1723,N_1538,N_1587);
nor U1724 (N_1724,N_1553,N_1501);
and U1725 (N_1725,N_1510,N_1544);
or U1726 (N_1726,N_1495,N_1473);
xor U1727 (N_1727,N_1538,N_1442);
and U1728 (N_1728,N_1538,N_1424);
nor U1729 (N_1729,N_1484,N_1414);
and U1730 (N_1730,N_1404,N_1503);
nand U1731 (N_1731,N_1581,N_1454);
or U1732 (N_1732,N_1519,N_1415);
and U1733 (N_1733,N_1476,N_1438);
nor U1734 (N_1734,N_1545,N_1554);
nand U1735 (N_1735,N_1486,N_1439);
or U1736 (N_1736,N_1469,N_1576);
nor U1737 (N_1737,N_1427,N_1459);
nand U1738 (N_1738,N_1558,N_1588);
or U1739 (N_1739,N_1497,N_1517);
nor U1740 (N_1740,N_1407,N_1436);
or U1741 (N_1741,N_1593,N_1404);
or U1742 (N_1742,N_1584,N_1572);
nor U1743 (N_1743,N_1442,N_1481);
and U1744 (N_1744,N_1570,N_1591);
or U1745 (N_1745,N_1476,N_1594);
and U1746 (N_1746,N_1474,N_1513);
and U1747 (N_1747,N_1453,N_1531);
or U1748 (N_1748,N_1469,N_1597);
or U1749 (N_1749,N_1427,N_1595);
and U1750 (N_1750,N_1534,N_1536);
xor U1751 (N_1751,N_1513,N_1532);
nor U1752 (N_1752,N_1589,N_1596);
nor U1753 (N_1753,N_1526,N_1557);
nor U1754 (N_1754,N_1513,N_1439);
or U1755 (N_1755,N_1462,N_1515);
nand U1756 (N_1756,N_1594,N_1449);
xnor U1757 (N_1757,N_1497,N_1473);
nand U1758 (N_1758,N_1414,N_1598);
and U1759 (N_1759,N_1522,N_1488);
nand U1760 (N_1760,N_1556,N_1465);
nand U1761 (N_1761,N_1485,N_1430);
and U1762 (N_1762,N_1529,N_1591);
nor U1763 (N_1763,N_1574,N_1519);
nor U1764 (N_1764,N_1543,N_1597);
or U1765 (N_1765,N_1416,N_1591);
nand U1766 (N_1766,N_1412,N_1414);
nand U1767 (N_1767,N_1536,N_1532);
nand U1768 (N_1768,N_1427,N_1460);
or U1769 (N_1769,N_1544,N_1527);
xor U1770 (N_1770,N_1583,N_1526);
and U1771 (N_1771,N_1546,N_1523);
and U1772 (N_1772,N_1559,N_1528);
xnor U1773 (N_1773,N_1423,N_1556);
nor U1774 (N_1774,N_1599,N_1446);
xor U1775 (N_1775,N_1513,N_1573);
nor U1776 (N_1776,N_1445,N_1522);
nor U1777 (N_1777,N_1427,N_1498);
nor U1778 (N_1778,N_1429,N_1452);
nor U1779 (N_1779,N_1459,N_1540);
xnor U1780 (N_1780,N_1564,N_1576);
nand U1781 (N_1781,N_1598,N_1504);
nor U1782 (N_1782,N_1593,N_1445);
nand U1783 (N_1783,N_1560,N_1409);
nor U1784 (N_1784,N_1420,N_1583);
nor U1785 (N_1785,N_1406,N_1512);
and U1786 (N_1786,N_1408,N_1551);
nor U1787 (N_1787,N_1452,N_1568);
nand U1788 (N_1788,N_1557,N_1404);
nand U1789 (N_1789,N_1582,N_1414);
or U1790 (N_1790,N_1472,N_1544);
nand U1791 (N_1791,N_1498,N_1479);
nand U1792 (N_1792,N_1480,N_1516);
nand U1793 (N_1793,N_1548,N_1559);
xnor U1794 (N_1794,N_1471,N_1456);
or U1795 (N_1795,N_1550,N_1438);
nand U1796 (N_1796,N_1430,N_1403);
nor U1797 (N_1797,N_1540,N_1512);
nand U1798 (N_1798,N_1475,N_1508);
or U1799 (N_1799,N_1595,N_1482);
or U1800 (N_1800,N_1681,N_1754);
nand U1801 (N_1801,N_1664,N_1672);
nor U1802 (N_1802,N_1707,N_1758);
nand U1803 (N_1803,N_1764,N_1651);
nand U1804 (N_1804,N_1771,N_1718);
and U1805 (N_1805,N_1716,N_1603);
and U1806 (N_1806,N_1663,N_1790);
and U1807 (N_1807,N_1655,N_1784);
xor U1808 (N_1808,N_1647,N_1714);
nand U1809 (N_1809,N_1608,N_1751);
or U1810 (N_1810,N_1649,N_1621);
and U1811 (N_1811,N_1682,N_1633);
or U1812 (N_1812,N_1782,N_1620);
or U1813 (N_1813,N_1629,N_1759);
xnor U1814 (N_1814,N_1753,N_1648);
nand U1815 (N_1815,N_1729,N_1695);
or U1816 (N_1816,N_1610,N_1722);
or U1817 (N_1817,N_1615,N_1743);
or U1818 (N_1818,N_1618,N_1792);
nand U1819 (N_1819,N_1631,N_1746);
and U1820 (N_1820,N_1781,N_1727);
and U1821 (N_1821,N_1600,N_1774);
nor U1822 (N_1822,N_1616,N_1699);
and U1823 (N_1823,N_1795,N_1674);
or U1824 (N_1824,N_1796,N_1731);
and U1825 (N_1825,N_1778,N_1747);
and U1826 (N_1826,N_1680,N_1737);
nand U1827 (N_1827,N_1789,N_1770);
nor U1828 (N_1828,N_1734,N_1689);
or U1829 (N_1829,N_1656,N_1619);
or U1830 (N_1830,N_1617,N_1657);
nand U1831 (N_1831,N_1724,N_1611);
or U1832 (N_1832,N_1653,N_1632);
and U1833 (N_1833,N_1660,N_1690);
or U1834 (N_1834,N_1742,N_1721);
nor U1835 (N_1835,N_1696,N_1791);
nand U1836 (N_1836,N_1725,N_1735);
nand U1837 (N_1837,N_1624,N_1756);
and U1838 (N_1838,N_1773,N_1794);
nor U1839 (N_1839,N_1654,N_1744);
or U1840 (N_1840,N_1694,N_1785);
nand U1841 (N_1841,N_1645,N_1669);
xor U1842 (N_1842,N_1652,N_1708);
nand U1843 (N_1843,N_1769,N_1772);
nor U1844 (N_1844,N_1644,N_1609);
xor U1845 (N_1845,N_1709,N_1787);
nor U1846 (N_1846,N_1755,N_1728);
or U1847 (N_1847,N_1639,N_1606);
or U1848 (N_1848,N_1625,N_1641);
and U1849 (N_1849,N_1676,N_1786);
xnor U1850 (N_1850,N_1730,N_1749);
nor U1851 (N_1851,N_1767,N_1640);
and U1852 (N_1852,N_1630,N_1702);
and U1853 (N_1853,N_1698,N_1678);
or U1854 (N_1854,N_1777,N_1738);
or U1855 (N_1855,N_1717,N_1797);
and U1856 (N_1856,N_1634,N_1622);
nor U1857 (N_1857,N_1684,N_1661);
and U1858 (N_1858,N_1692,N_1761);
nand U1859 (N_1859,N_1799,N_1688);
xnor U1860 (N_1860,N_1750,N_1732);
nand U1861 (N_1861,N_1703,N_1776);
or U1862 (N_1862,N_1668,N_1704);
and U1863 (N_1863,N_1673,N_1670);
or U1864 (N_1864,N_1768,N_1710);
nor U1865 (N_1865,N_1706,N_1671);
nand U1866 (N_1866,N_1793,N_1604);
and U1867 (N_1867,N_1628,N_1745);
or U1868 (N_1868,N_1780,N_1642);
xor U1869 (N_1869,N_1605,N_1783);
and U1870 (N_1870,N_1677,N_1602);
and U1871 (N_1871,N_1798,N_1691);
xnor U1872 (N_1872,N_1765,N_1752);
or U1873 (N_1873,N_1686,N_1779);
nand U1874 (N_1874,N_1739,N_1766);
nor U1875 (N_1875,N_1614,N_1726);
xor U1876 (N_1876,N_1685,N_1713);
nor U1877 (N_1877,N_1757,N_1635);
or U1878 (N_1878,N_1623,N_1636);
or U1879 (N_1879,N_1650,N_1601);
nor U1880 (N_1880,N_1701,N_1658);
nor U1881 (N_1881,N_1687,N_1715);
nor U1882 (N_1882,N_1613,N_1665);
and U1883 (N_1883,N_1693,N_1763);
and U1884 (N_1884,N_1705,N_1607);
nand U1885 (N_1885,N_1683,N_1662);
nor U1886 (N_1886,N_1700,N_1740);
nor U1887 (N_1887,N_1646,N_1775);
nor U1888 (N_1888,N_1720,N_1667);
and U1889 (N_1889,N_1748,N_1679);
or U1890 (N_1890,N_1627,N_1659);
nor U1891 (N_1891,N_1697,N_1762);
or U1892 (N_1892,N_1736,N_1612);
xor U1893 (N_1893,N_1638,N_1711);
xnor U1894 (N_1894,N_1712,N_1741);
or U1895 (N_1895,N_1760,N_1643);
nor U1896 (N_1896,N_1719,N_1733);
and U1897 (N_1897,N_1675,N_1666);
nor U1898 (N_1898,N_1626,N_1788);
and U1899 (N_1899,N_1637,N_1723);
and U1900 (N_1900,N_1769,N_1768);
nor U1901 (N_1901,N_1642,N_1781);
or U1902 (N_1902,N_1618,N_1724);
or U1903 (N_1903,N_1617,N_1726);
xnor U1904 (N_1904,N_1777,N_1618);
nor U1905 (N_1905,N_1655,N_1758);
nand U1906 (N_1906,N_1619,N_1722);
xnor U1907 (N_1907,N_1725,N_1757);
and U1908 (N_1908,N_1714,N_1680);
or U1909 (N_1909,N_1628,N_1638);
and U1910 (N_1910,N_1682,N_1733);
or U1911 (N_1911,N_1633,N_1794);
nor U1912 (N_1912,N_1719,N_1775);
or U1913 (N_1913,N_1772,N_1677);
nor U1914 (N_1914,N_1780,N_1657);
and U1915 (N_1915,N_1743,N_1628);
or U1916 (N_1916,N_1614,N_1616);
and U1917 (N_1917,N_1792,N_1760);
nor U1918 (N_1918,N_1774,N_1715);
or U1919 (N_1919,N_1758,N_1732);
or U1920 (N_1920,N_1704,N_1606);
and U1921 (N_1921,N_1723,N_1665);
xnor U1922 (N_1922,N_1733,N_1720);
or U1923 (N_1923,N_1750,N_1798);
and U1924 (N_1924,N_1637,N_1714);
nor U1925 (N_1925,N_1628,N_1695);
nor U1926 (N_1926,N_1748,N_1606);
and U1927 (N_1927,N_1622,N_1657);
and U1928 (N_1928,N_1637,N_1721);
nor U1929 (N_1929,N_1618,N_1683);
and U1930 (N_1930,N_1745,N_1715);
and U1931 (N_1931,N_1630,N_1600);
nor U1932 (N_1932,N_1780,N_1674);
nor U1933 (N_1933,N_1769,N_1626);
nand U1934 (N_1934,N_1627,N_1786);
nand U1935 (N_1935,N_1608,N_1715);
xor U1936 (N_1936,N_1657,N_1648);
or U1937 (N_1937,N_1744,N_1646);
and U1938 (N_1938,N_1657,N_1799);
nor U1939 (N_1939,N_1638,N_1625);
or U1940 (N_1940,N_1742,N_1636);
nand U1941 (N_1941,N_1734,N_1629);
nand U1942 (N_1942,N_1727,N_1763);
or U1943 (N_1943,N_1676,N_1668);
nor U1944 (N_1944,N_1756,N_1754);
and U1945 (N_1945,N_1693,N_1713);
and U1946 (N_1946,N_1664,N_1797);
and U1947 (N_1947,N_1742,N_1758);
and U1948 (N_1948,N_1750,N_1767);
nor U1949 (N_1949,N_1774,N_1775);
xor U1950 (N_1950,N_1700,N_1673);
and U1951 (N_1951,N_1750,N_1754);
nand U1952 (N_1952,N_1626,N_1637);
nor U1953 (N_1953,N_1735,N_1622);
nor U1954 (N_1954,N_1759,N_1717);
nand U1955 (N_1955,N_1606,N_1781);
and U1956 (N_1956,N_1694,N_1653);
nand U1957 (N_1957,N_1674,N_1725);
xor U1958 (N_1958,N_1695,N_1775);
and U1959 (N_1959,N_1674,N_1700);
or U1960 (N_1960,N_1639,N_1652);
or U1961 (N_1961,N_1777,N_1640);
nor U1962 (N_1962,N_1633,N_1645);
nor U1963 (N_1963,N_1799,N_1786);
nor U1964 (N_1964,N_1601,N_1609);
nand U1965 (N_1965,N_1602,N_1640);
nand U1966 (N_1966,N_1656,N_1658);
or U1967 (N_1967,N_1642,N_1720);
nand U1968 (N_1968,N_1772,N_1722);
nand U1969 (N_1969,N_1647,N_1798);
nor U1970 (N_1970,N_1614,N_1653);
nand U1971 (N_1971,N_1677,N_1732);
nand U1972 (N_1972,N_1703,N_1659);
nand U1973 (N_1973,N_1629,N_1707);
nor U1974 (N_1974,N_1624,N_1612);
nor U1975 (N_1975,N_1786,N_1770);
and U1976 (N_1976,N_1621,N_1670);
nand U1977 (N_1977,N_1668,N_1743);
nand U1978 (N_1978,N_1673,N_1638);
or U1979 (N_1979,N_1695,N_1697);
or U1980 (N_1980,N_1628,N_1657);
and U1981 (N_1981,N_1627,N_1732);
and U1982 (N_1982,N_1799,N_1774);
and U1983 (N_1983,N_1795,N_1717);
and U1984 (N_1984,N_1661,N_1672);
nand U1985 (N_1985,N_1780,N_1614);
xor U1986 (N_1986,N_1643,N_1779);
or U1987 (N_1987,N_1770,N_1745);
nand U1988 (N_1988,N_1688,N_1653);
xnor U1989 (N_1989,N_1637,N_1796);
nor U1990 (N_1990,N_1736,N_1627);
xnor U1991 (N_1991,N_1733,N_1665);
and U1992 (N_1992,N_1741,N_1674);
nor U1993 (N_1993,N_1621,N_1690);
and U1994 (N_1994,N_1779,N_1664);
or U1995 (N_1995,N_1627,N_1604);
xor U1996 (N_1996,N_1611,N_1607);
nand U1997 (N_1997,N_1658,N_1789);
or U1998 (N_1998,N_1726,N_1698);
or U1999 (N_1999,N_1780,N_1799);
or U2000 (N_2000,N_1932,N_1829);
or U2001 (N_2001,N_1995,N_1843);
or U2002 (N_2002,N_1855,N_1884);
xor U2003 (N_2003,N_1980,N_1894);
nand U2004 (N_2004,N_1826,N_1989);
nor U2005 (N_2005,N_1975,N_1857);
nor U2006 (N_2006,N_1941,N_1981);
nor U2007 (N_2007,N_1946,N_1871);
or U2008 (N_2008,N_1830,N_1921);
and U2009 (N_2009,N_1860,N_1994);
xor U2010 (N_2010,N_1991,N_1922);
or U2011 (N_2011,N_1923,N_1859);
or U2012 (N_2012,N_1848,N_1863);
nand U2013 (N_2013,N_1920,N_1952);
nor U2014 (N_2014,N_1937,N_1891);
nand U2015 (N_2015,N_1953,N_1969);
or U2016 (N_2016,N_1962,N_1806);
and U2017 (N_2017,N_1868,N_1893);
nand U2018 (N_2018,N_1869,N_1899);
nor U2019 (N_2019,N_1892,N_1934);
nor U2020 (N_2020,N_1812,N_1943);
nor U2021 (N_2021,N_1822,N_1902);
nor U2022 (N_2022,N_1847,N_1842);
nor U2023 (N_2023,N_1909,N_1808);
nor U2024 (N_2024,N_1942,N_1963);
and U2025 (N_2025,N_1940,N_1901);
nand U2026 (N_2026,N_1992,N_1956);
nor U2027 (N_2027,N_1982,N_1895);
or U2028 (N_2028,N_1906,N_1972);
nand U2029 (N_2029,N_1861,N_1834);
nor U2030 (N_2030,N_1805,N_1957);
and U2031 (N_2031,N_1846,N_1927);
or U2032 (N_2032,N_1961,N_1947);
nor U2033 (N_2033,N_1880,N_1964);
or U2034 (N_2034,N_1827,N_1955);
nand U2035 (N_2035,N_1878,N_1944);
and U2036 (N_2036,N_1983,N_1910);
nor U2037 (N_2037,N_1973,N_1990);
and U2038 (N_2038,N_1925,N_1960);
and U2039 (N_2039,N_1959,N_1810);
xnor U2040 (N_2040,N_1974,N_1832);
xnor U2041 (N_2041,N_1851,N_1821);
nand U2042 (N_2042,N_1801,N_1837);
nand U2043 (N_2043,N_1881,N_1935);
nor U2044 (N_2044,N_1879,N_1800);
or U2045 (N_2045,N_1896,N_1933);
or U2046 (N_2046,N_1882,N_1874);
or U2047 (N_2047,N_1887,N_1915);
nand U2048 (N_2048,N_1838,N_1862);
or U2049 (N_2049,N_1905,N_1802);
nor U2050 (N_2050,N_1888,N_1954);
nor U2051 (N_2051,N_1841,N_1885);
or U2052 (N_2052,N_1967,N_1986);
or U2053 (N_2053,N_1819,N_1889);
xnor U2054 (N_2054,N_1886,N_1907);
and U2055 (N_2055,N_1870,N_1977);
nand U2056 (N_2056,N_1997,N_1850);
nand U2057 (N_2057,N_1976,N_1864);
nor U2058 (N_2058,N_1970,N_1823);
and U2059 (N_2059,N_1979,N_1856);
or U2060 (N_2060,N_1965,N_1996);
xnor U2061 (N_2061,N_1950,N_1936);
xor U2062 (N_2062,N_1814,N_1945);
or U2063 (N_2063,N_1903,N_1804);
or U2064 (N_2064,N_1833,N_1924);
nand U2065 (N_2065,N_1968,N_1825);
and U2066 (N_2066,N_1912,N_1914);
xnor U2067 (N_2067,N_1815,N_1985);
and U2068 (N_2068,N_1897,N_1807);
nor U2069 (N_2069,N_1858,N_1839);
and U2070 (N_2070,N_1877,N_1908);
and U2071 (N_2071,N_1811,N_1984);
or U2072 (N_2072,N_1873,N_1867);
nor U2073 (N_2073,N_1828,N_1958);
nand U2074 (N_2074,N_1844,N_1926);
nand U2075 (N_2075,N_1813,N_1809);
nor U2076 (N_2076,N_1883,N_1890);
and U2077 (N_2077,N_1951,N_1900);
or U2078 (N_2078,N_1816,N_1898);
xor U2079 (N_2079,N_1919,N_1872);
nand U2080 (N_2080,N_1918,N_1971);
xnor U2081 (N_2081,N_1803,N_1911);
nand U2082 (N_2082,N_1852,N_1917);
nand U2083 (N_2083,N_1948,N_1916);
nand U2084 (N_2084,N_1854,N_1820);
or U2085 (N_2085,N_1949,N_1939);
nand U2086 (N_2086,N_1929,N_1904);
nor U2087 (N_2087,N_1849,N_1865);
or U2088 (N_2088,N_1876,N_1836);
or U2089 (N_2089,N_1866,N_1824);
or U2090 (N_2090,N_1928,N_1978);
nor U2091 (N_2091,N_1930,N_1818);
xnor U2092 (N_2092,N_1913,N_1998);
or U2093 (N_2093,N_1999,N_1817);
and U2094 (N_2094,N_1966,N_1875);
nand U2095 (N_2095,N_1845,N_1853);
nand U2096 (N_2096,N_1831,N_1931);
nor U2097 (N_2097,N_1835,N_1987);
or U2098 (N_2098,N_1938,N_1988);
nor U2099 (N_2099,N_1840,N_1993);
nor U2100 (N_2100,N_1858,N_1916);
or U2101 (N_2101,N_1861,N_1859);
and U2102 (N_2102,N_1849,N_1896);
nor U2103 (N_2103,N_1808,N_1939);
nor U2104 (N_2104,N_1919,N_1884);
and U2105 (N_2105,N_1909,N_1880);
and U2106 (N_2106,N_1837,N_1954);
and U2107 (N_2107,N_1958,N_1961);
nor U2108 (N_2108,N_1959,N_1877);
nand U2109 (N_2109,N_1825,N_1870);
and U2110 (N_2110,N_1844,N_1906);
xnor U2111 (N_2111,N_1982,N_1907);
and U2112 (N_2112,N_1802,N_1930);
and U2113 (N_2113,N_1802,N_1949);
xnor U2114 (N_2114,N_1887,N_1877);
or U2115 (N_2115,N_1962,N_1940);
and U2116 (N_2116,N_1820,N_1895);
nand U2117 (N_2117,N_1818,N_1896);
and U2118 (N_2118,N_1920,N_1818);
or U2119 (N_2119,N_1979,N_1816);
and U2120 (N_2120,N_1938,N_1965);
xor U2121 (N_2121,N_1997,N_1828);
nand U2122 (N_2122,N_1819,N_1854);
and U2123 (N_2123,N_1830,N_1892);
nand U2124 (N_2124,N_1921,N_1944);
nand U2125 (N_2125,N_1938,N_1918);
nor U2126 (N_2126,N_1980,N_1836);
nand U2127 (N_2127,N_1958,N_1910);
and U2128 (N_2128,N_1891,N_1819);
xor U2129 (N_2129,N_1846,N_1930);
nor U2130 (N_2130,N_1939,N_1925);
nand U2131 (N_2131,N_1937,N_1876);
and U2132 (N_2132,N_1895,N_1886);
and U2133 (N_2133,N_1804,N_1966);
xor U2134 (N_2134,N_1893,N_1959);
and U2135 (N_2135,N_1951,N_1988);
nor U2136 (N_2136,N_1923,N_1845);
nand U2137 (N_2137,N_1806,N_1811);
or U2138 (N_2138,N_1872,N_1918);
nor U2139 (N_2139,N_1896,N_1962);
or U2140 (N_2140,N_1888,N_1851);
and U2141 (N_2141,N_1935,N_1985);
nand U2142 (N_2142,N_1917,N_1951);
nand U2143 (N_2143,N_1999,N_1854);
or U2144 (N_2144,N_1815,N_1885);
and U2145 (N_2145,N_1991,N_1978);
nand U2146 (N_2146,N_1913,N_1811);
nand U2147 (N_2147,N_1976,N_1809);
xnor U2148 (N_2148,N_1875,N_1810);
or U2149 (N_2149,N_1887,N_1994);
xor U2150 (N_2150,N_1977,N_1806);
nand U2151 (N_2151,N_1952,N_1882);
nand U2152 (N_2152,N_1902,N_1940);
and U2153 (N_2153,N_1951,N_1883);
nand U2154 (N_2154,N_1824,N_1899);
nor U2155 (N_2155,N_1895,N_1941);
nor U2156 (N_2156,N_1843,N_1960);
nand U2157 (N_2157,N_1871,N_1847);
nor U2158 (N_2158,N_1910,N_1900);
nor U2159 (N_2159,N_1850,N_1978);
nand U2160 (N_2160,N_1952,N_1823);
or U2161 (N_2161,N_1954,N_1980);
nand U2162 (N_2162,N_1876,N_1983);
and U2163 (N_2163,N_1829,N_1937);
nor U2164 (N_2164,N_1830,N_1992);
nor U2165 (N_2165,N_1883,N_1831);
nand U2166 (N_2166,N_1910,N_1985);
xnor U2167 (N_2167,N_1921,N_1994);
and U2168 (N_2168,N_1915,N_1850);
nand U2169 (N_2169,N_1914,N_1825);
or U2170 (N_2170,N_1989,N_1811);
nand U2171 (N_2171,N_1978,N_1981);
xor U2172 (N_2172,N_1874,N_1950);
and U2173 (N_2173,N_1824,N_1963);
and U2174 (N_2174,N_1862,N_1992);
xor U2175 (N_2175,N_1999,N_1988);
nand U2176 (N_2176,N_1801,N_1997);
and U2177 (N_2177,N_1989,N_1853);
nand U2178 (N_2178,N_1963,N_1950);
nor U2179 (N_2179,N_1852,N_1920);
nand U2180 (N_2180,N_1815,N_1913);
nor U2181 (N_2181,N_1921,N_1978);
or U2182 (N_2182,N_1980,N_1926);
nor U2183 (N_2183,N_1822,N_1988);
or U2184 (N_2184,N_1908,N_1951);
or U2185 (N_2185,N_1956,N_1846);
and U2186 (N_2186,N_1961,N_1825);
nor U2187 (N_2187,N_1979,N_1850);
or U2188 (N_2188,N_1964,N_1851);
and U2189 (N_2189,N_1823,N_1831);
nand U2190 (N_2190,N_1942,N_1968);
and U2191 (N_2191,N_1988,N_1831);
nand U2192 (N_2192,N_1989,N_1812);
nor U2193 (N_2193,N_1927,N_1823);
or U2194 (N_2194,N_1852,N_1938);
nor U2195 (N_2195,N_1957,N_1813);
and U2196 (N_2196,N_1966,N_1965);
and U2197 (N_2197,N_1846,N_1878);
or U2198 (N_2198,N_1867,N_1894);
and U2199 (N_2199,N_1920,N_1812);
nand U2200 (N_2200,N_2000,N_2047);
nor U2201 (N_2201,N_2018,N_2193);
and U2202 (N_2202,N_2188,N_2015);
or U2203 (N_2203,N_2100,N_2174);
xnor U2204 (N_2204,N_2008,N_2079);
nand U2205 (N_2205,N_2041,N_2032);
or U2206 (N_2206,N_2111,N_2068);
nand U2207 (N_2207,N_2140,N_2034);
and U2208 (N_2208,N_2120,N_2141);
and U2209 (N_2209,N_2148,N_2116);
xor U2210 (N_2210,N_2089,N_2164);
and U2211 (N_2211,N_2057,N_2064);
and U2212 (N_2212,N_2009,N_2092);
or U2213 (N_2213,N_2078,N_2155);
xnor U2214 (N_2214,N_2048,N_2112);
nand U2215 (N_2215,N_2090,N_2051);
or U2216 (N_2216,N_2022,N_2136);
xnor U2217 (N_2217,N_2172,N_2045);
nand U2218 (N_2218,N_2049,N_2102);
nand U2219 (N_2219,N_2131,N_2128);
nand U2220 (N_2220,N_2161,N_2012);
nor U2221 (N_2221,N_2184,N_2165);
nand U2222 (N_2222,N_2030,N_2042);
nand U2223 (N_2223,N_2087,N_2139);
or U2224 (N_2224,N_2154,N_2053);
nand U2225 (N_2225,N_2084,N_2010);
and U2226 (N_2226,N_2001,N_2098);
or U2227 (N_2227,N_2198,N_2007);
xor U2228 (N_2228,N_2138,N_2176);
or U2229 (N_2229,N_2003,N_2014);
and U2230 (N_2230,N_2150,N_2023);
or U2231 (N_2231,N_2028,N_2145);
nor U2232 (N_2232,N_2011,N_2126);
or U2233 (N_2233,N_2134,N_2059);
nand U2234 (N_2234,N_2113,N_2058);
or U2235 (N_2235,N_2072,N_2081);
nor U2236 (N_2236,N_2080,N_2189);
nor U2237 (N_2237,N_2105,N_2151);
and U2238 (N_2238,N_2152,N_2027);
xnor U2239 (N_2239,N_2135,N_2075);
and U2240 (N_2240,N_2107,N_2187);
or U2241 (N_2241,N_2196,N_2044);
or U2242 (N_2242,N_2061,N_2142);
xor U2243 (N_2243,N_2056,N_2195);
nor U2244 (N_2244,N_2173,N_2006);
or U2245 (N_2245,N_2181,N_2066);
and U2246 (N_2246,N_2117,N_2082);
or U2247 (N_2247,N_2017,N_2086);
or U2248 (N_2248,N_2185,N_2191);
and U2249 (N_2249,N_2088,N_2149);
nor U2250 (N_2250,N_2130,N_2095);
or U2251 (N_2251,N_2108,N_2115);
and U2252 (N_2252,N_2123,N_2192);
nand U2253 (N_2253,N_2124,N_2063);
nand U2254 (N_2254,N_2043,N_2016);
nand U2255 (N_2255,N_2067,N_2077);
nand U2256 (N_2256,N_2050,N_2157);
nor U2257 (N_2257,N_2166,N_2099);
nand U2258 (N_2258,N_2071,N_2167);
or U2259 (N_2259,N_2033,N_2055);
nor U2260 (N_2260,N_2175,N_2093);
and U2261 (N_2261,N_2036,N_2127);
or U2262 (N_2262,N_2073,N_2038);
or U2263 (N_2263,N_2106,N_2160);
nand U2264 (N_2264,N_2025,N_2026);
nand U2265 (N_2265,N_2162,N_2122);
and U2266 (N_2266,N_2013,N_2186);
nor U2267 (N_2267,N_2029,N_2020);
xnor U2268 (N_2268,N_2182,N_2133);
nor U2269 (N_2269,N_2132,N_2085);
and U2270 (N_2270,N_2158,N_2119);
nand U2271 (N_2271,N_2019,N_2060);
nand U2272 (N_2272,N_2171,N_2070);
xor U2273 (N_2273,N_2110,N_2194);
and U2274 (N_2274,N_2144,N_2004);
and U2275 (N_2275,N_2163,N_2125);
nor U2276 (N_2276,N_2104,N_2168);
or U2277 (N_2277,N_2180,N_2002);
nand U2278 (N_2278,N_2101,N_2052);
and U2279 (N_2279,N_2062,N_2199);
nand U2280 (N_2280,N_2159,N_2103);
and U2281 (N_2281,N_2083,N_2040);
and U2282 (N_2282,N_2021,N_2076);
and U2283 (N_2283,N_2109,N_2035);
and U2284 (N_2284,N_2096,N_2069);
nand U2285 (N_2285,N_2137,N_2065);
nand U2286 (N_2286,N_2114,N_2156);
nor U2287 (N_2287,N_2054,N_2005);
nor U2288 (N_2288,N_2153,N_2143);
nand U2289 (N_2289,N_2037,N_2183);
and U2290 (N_2290,N_2177,N_2190);
nand U2291 (N_2291,N_2031,N_2169);
nand U2292 (N_2292,N_2024,N_2129);
nor U2293 (N_2293,N_2074,N_2147);
or U2294 (N_2294,N_2046,N_2039);
nand U2295 (N_2295,N_2118,N_2094);
and U2296 (N_2296,N_2091,N_2197);
or U2297 (N_2297,N_2179,N_2170);
nand U2298 (N_2298,N_2097,N_2178);
nor U2299 (N_2299,N_2121,N_2146);
or U2300 (N_2300,N_2107,N_2017);
and U2301 (N_2301,N_2045,N_2115);
and U2302 (N_2302,N_2087,N_2186);
and U2303 (N_2303,N_2103,N_2114);
or U2304 (N_2304,N_2132,N_2163);
nor U2305 (N_2305,N_2015,N_2060);
or U2306 (N_2306,N_2133,N_2047);
and U2307 (N_2307,N_2120,N_2189);
nor U2308 (N_2308,N_2189,N_2006);
nand U2309 (N_2309,N_2109,N_2179);
and U2310 (N_2310,N_2062,N_2003);
and U2311 (N_2311,N_2159,N_2179);
or U2312 (N_2312,N_2038,N_2199);
or U2313 (N_2313,N_2180,N_2023);
or U2314 (N_2314,N_2057,N_2019);
nand U2315 (N_2315,N_2091,N_2060);
nand U2316 (N_2316,N_2020,N_2152);
nand U2317 (N_2317,N_2073,N_2032);
and U2318 (N_2318,N_2176,N_2104);
or U2319 (N_2319,N_2175,N_2023);
xnor U2320 (N_2320,N_2131,N_2024);
or U2321 (N_2321,N_2023,N_2189);
and U2322 (N_2322,N_2049,N_2168);
nor U2323 (N_2323,N_2162,N_2173);
nand U2324 (N_2324,N_2076,N_2029);
or U2325 (N_2325,N_2147,N_2120);
and U2326 (N_2326,N_2083,N_2137);
nand U2327 (N_2327,N_2015,N_2034);
xor U2328 (N_2328,N_2063,N_2040);
and U2329 (N_2329,N_2147,N_2056);
nor U2330 (N_2330,N_2155,N_2167);
nor U2331 (N_2331,N_2105,N_2135);
or U2332 (N_2332,N_2128,N_2155);
nand U2333 (N_2333,N_2147,N_2191);
and U2334 (N_2334,N_2014,N_2073);
and U2335 (N_2335,N_2048,N_2003);
and U2336 (N_2336,N_2069,N_2127);
xnor U2337 (N_2337,N_2076,N_2010);
xor U2338 (N_2338,N_2182,N_2025);
xnor U2339 (N_2339,N_2195,N_2006);
nor U2340 (N_2340,N_2097,N_2156);
nand U2341 (N_2341,N_2065,N_2088);
nor U2342 (N_2342,N_2040,N_2179);
nand U2343 (N_2343,N_2022,N_2151);
nand U2344 (N_2344,N_2173,N_2142);
or U2345 (N_2345,N_2106,N_2051);
and U2346 (N_2346,N_2020,N_2120);
xor U2347 (N_2347,N_2049,N_2010);
or U2348 (N_2348,N_2118,N_2027);
nand U2349 (N_2349,N_2197,N_2159);
or U2350 (N_2350,N_2149,N_2014);
or U2351 (N_2351,N_2176,N_2156);
and U2352 (N_2352,N_2101,N_2058);
or U2353 (N_2353,N_2093,N_2146);
xnor U2354 (N_2354,N_2031,N_2079);
nand U2355 (N_2355,N_2168,N_2056);
nor U2356 (N_2356,N_2016,N_2010);
or U2357 (N_2357,N_2148,N_2099);
and U2358 (N_2358,N_2185,N_2140);
or U2359 (N_2359,N_2164,N_2074);
or U2360 (N_2360,N_2040,N_2004);
nand U2361 (N_2361,N_2091,N_2078);
nor U2362 (N_2362,N_2015,N_2014);
or U2363 (N_2363,N_2051,N_2123);
and U2364 (N_2364,N_2188,N_2124);
and U2365 (N_2365,N_2018,N_2087);
and U2366 (N_2366,N_2155,N_2096);
and U2367 (N_2367,N_2189,N_2135);
nor U2368 (N_2368,N_2152,N_2168);
nor U2369 (N_2369,N_2157,N_2061);
and U2370 (N_2370,N_2016,N_2127);
nand U2371 (N_2371,N_2150,N_2189);
xnor U2372 (N_2372,N_2063,N_2169);
nand U2373 (N_2373,N_2089,N_2044);
or U2374 (N_2374,N_2016,N_2154);
or U2375 (N_2375,N_2171,N_2165);
xor U2376 (N_2376,N_2172,N_2121);
or U2377 (N_2377,N_2149,N_2054);
nand U2378 (N_2378,N_2087,N_2193);
or U2379 (N_2379,N_2136,N_2011);
xnor U2380 (N_2380,N_2141,N_2000);
or U2381 (N_2381,N_2126,N_2067);
or U2382 (N_2382,N_2193,N_2031);
nor U2383 (N_2383,N_2011,N_2183);
and U2384 (N_2384,N_2026,N_2077);
nand U2385 (N_2385,N_2088,N_2061);
or U2386 (N_2386,N_2158,N_2181);
or U2387 (N_2387,N_2103,N_2023);
nor U2388 (N_2388,N_2035,N_2017);
or U2389 (N_2389,N_2106,N_2105);
nand U2390 (N_2390,N_2170,N_2193);
nand U2391 (N_2391,N_2181,N_2134);
and U2392 (N_2392,N_2133,N_2073);
xor U2393 (N_2393,N_2165,N_2114);
nand U2394 (N_2394,N_2099,N_2126);
nand U2395 (N_2395,N_2095,N_2023);
xor U2396 (N_2396,N_2171,N_2120);
nor U2397 (N_2397,N_2123,N_2065);
nor U2398 (N_2398,N_2032,N_2085);
nor U2399 (N_2399,N_2101,N_2047);
and U2400 (N_2400,N_2251,N_2346);
nand U2401 (N_2401,N_2301,N_2385);
nor U2402 (N_2402,N_2286,N_2265);
nand U2403 (N_2403,N_2348,N_2354);
xnor U2404 (N_2404,N_2377,N_2389);
xor U2405 (N_2405,N_2374,N_2261);
nand U2406 (N_2406,N_2298,N_2368);
and U2407 (N_2407,N_2362,N_2337);
or U2408 (N_2408,N_2339,N_2322);
nor U2409 (N_2409,N_2342,N_2314);
and U2410 (N_2410,N_2370,N_2258);
or U2411 (N_2411,N_2231,N_2257);
and U2412 (N_2412,N_2280,N_2200);
nor U2413 (N_2413,N_2313,N_2390);
nor U2414 (N_2414,N_2387,N_2290);
nor U2415 (N_2415,N_2309,N_2204);
nand U2416 (N_2416,N_2276,N_2352);
or U2417 (N_2417,N_2376,N_2344);
and U2418 (N_2418,N_2287,N_2224);
or U2419 (N_2419,N_2304,N_2328);
nand U2420 (N_2420,N_2321,N_2266);
nand U2421 (N_2421,N_2243,N_2375);
or U2422 (N_2422,N_2356,N_2212);
nand U2423 (N_2423,N_2351,N_2210);
nand U2424 (N_2424,N_2310,N_2221);
or U2425 (N_2425,N_2383,N_2273);
or U2426 (N_2426,N_2215,N_2392);
nand U2427 (N_2427,N_2270,N_2271);
xnor U2428 (N_2428,N_2229,N_2399);
and U2429 (N_2429,N_2343,N_2317);
nor U2430 (N_2430,N_2358,N_2260);
xor U2431 (N_2431,N_2217,N_2359);
nor U2432 (N_2432,N_2253,N_2335);
nor U2433 (N_2433,N_2277,N_2203);
or U2434 (N_2434,N_2331,N_2325);
or U2435 (N_2435,N_2249,N_2233);
nor U2436 (N_2436,N_2275,N_2338);
or U2437 (N_2437,N_2380,N_2236);
xnor U2438 (N_2438,N_2207,N_2355);
and U2439 (N_2439,N_2361,N_2311);
nor U2440 (N_2440,N_2283,N_2213);
and U2441 (N_2441,N_2388,N_2255);
nand U2442 (N_2442,N_2391,N_2378);
nor U2443 (N_2443,N_2289,N_2206);
and U2444 (N_2444,N_2396,N_2244);
or U2445 (N_2445,N_2205,N_2272);
xnor U2446 (N_2446,N_2284,N_2336);
nor U2447 (N_2447,N_2295,N_2382);
or U2448 (N_2448,N_2240,N_2341);
nand U2449 (N_2449,N_2211,N_2237);
and U2450 (N_2450,N_2372,N_2208);
nor U2451 (N_2451,N_2293,N_2305);
and U2452 (N_2452,N_2230,N_2226);
and U2453 (N_2453,N_2278,N_2274);
nor U2454 (N_2454,N_2347,N_2345);
and U2455 (N_2455,N_2291,N_2294);
or U2456 (N_2456,N_2367,N_2246);
and U2457 (N_2457,N_2302,N_2220);
or U2458 (N_2458,N_2223,N_2364);
or U2459 (N_2459,N_2279,N_2299);
and U2460 (N_2460,N_2242,N_2259);
nand U2461 (N_2461,N_2235,N_2324);
nor U2462 (N_2462,N_2381,N_2268);
nor U2463 (N_2463,N_2267,N_2366);
and U2464 (N_2464,N_2334,N_2292);
nor U2465 (N_2465,N_2201,N_2239);
nand U2466 (N_2466,N_2363,N_2329);
nor U2467 (N_2467,N_2256,N_2319);
and U2468 (N_2468,N_2318,N_2357);
nor U2469 (N_2469,N_2252,N_2264);
nor U2470 (N_2470,N_2296,N_2225);
or U2471 (N_2471,N_2247,N_2269);
xor U2472 (N_2472,N_2369,N_2263);
or U2473 (N_2473,N_2397,N_2350);
nand U2474 (N_2474,N_2327,N_2326);
nor U2475 (N_2475,N_2306,N_2232);
nand U2476 (N_2476,N_2312,N_2282);
nand U2477 (N_2477,N_2218,N_2373);
nor U2478 (N_2478,N_2395,N_2332);
nor U2479 (N_2479,N_2297,N_2320);
nand U2480 (N_2480,N_2262,N_2254);
or U2481 (N_2481,N_2209,N_2227);
xor U2482 (N_2482,N_2379,N_2288);
or U2483 (N_2483,N_2222,N_2386);
nor U2484 (N_2484,N_2228,N_2308);
or U2485 (N_2485,N_2216,N_2315);
or U2486 (N_2486,N_2234,N_2371);
nand U2487 (N_2487,N_2333,N_2316);
and U2488 (N_2488,N_2365,N_2307);
nor U2489 (N_2489,N_2250,N_2394);
and U2490 (N_2490,N_2330,N_2281);
xor U2491 (N_2491,N_2202,N_2238);
nand U2492 (N_2492,N_2214,N_2398);
nand U2493 (N_2493,N_2245,N_2241);
nand U2494 (N_2494,N_2219,N_2303);
nor U2495 (N_2495,N_2340,N_2248);
and U2496 (N_2496,N_2285,N_2393);
nand U2497 (N_2497,N_2353,N_2323);
and U2498 (N_2498,N_2349,N_2300);
and U2499 (N_2499,N_2360,N_2384);
xnor U2500 (N_2500,N_2294,N_2381);
nand U2501 (N_2501,N_2273,N_2232);
nor U2502 (N_2502,N_2381,N_2344);
and U2503 (N_2503,N_2329,N_2392);
nor U2504 (N_2504,N_2265,N_2308);
and U2505 (N_2505,N_2217,N_2309);
nand U2506 (N_2506,N_2389,N_2284);
nor U2507 (N_2507,N_2282,N_2210);
or U2508 (N_2508,N_2201,N_2202);
and U2509 (N_2509,N_2249,N_2277);
or U2510 (N_2510,N_2329,N_2300);
and U2511 (N_2511,N_2348,N_2356);
xnor U2512 (N_2512,N_2302,N_2351);
or U2513 (N_2513,N_2330,N_2233);
or U2514 (N_2514,N_2224,N_2250);
and U2515 (N_2515,N_2212,N_2233);
nor U2516 (N_2516,N_2338,N_2395);
or U2517 (N_2517,N_2226,N_2398);
nor U2518 (N_2518,N_2219,N_2249);
nand U2519 (N_2519,N_2313,N_2289);
nor U2520 (N_2520,N_2331,N_2298);
or U2521 (N_2521,N_2334,N_2361);
nand U2522 (N_2522,N_2386,N_2389);
and U2523 (N_2523,N_2389,N_2249);
or U2524 (N_2524,N_2334,N_2222);
and U2525 (N_2525,N_2370,N_2243);
and U2526 (N_2526,N_2319,N_2259);
or U2527 (N_2527,N_2228,N_2345);
xor U2528 (N_2528,N_2384,N_2329);
xor U2529 (N_2529,N_2267,N_2293);
and U2530 (N_2530,N_2346,N_2363);
and U2531 (N_2531,N_2284,N_2256);
nand U2532 (N_2532,N_2247,N_2326);
or U2533 (N_2533,N_2300,N_2208);
xnor U2534 (N_2534,N_2310,N_2276);
nand U2535 (N_2535,N_2347,N_2290);
nand U2536 (N_2536,N_2397,N_2249);
and U2537 (N_2537,N_2229,N_2222);
and U2538 (N_2538,N_2248,N_2260);
and U2539 (N_2539,N_2207,N_2309);
and U2540 (N_2540,N_2201,N_2254);
nand U2541 (N_2541,N_2331,N_2320);
and U2542 (N_2542,N_2273,N_2228);
or U2543 (N_2543,N_2221,N_2342);
xor U2544 (N_2544,N_2262,N_2221);
nand U2545 (N_2545,N_2385,N_2222);
nor U2546 (N_2546,N_2232,N_2384);
and U2547 (N_2547,N_2206,N_2256);
and U2548 (N_2548,N_2281,N_2326);
and U2549 (N_2549,N_2245,N_2380);
nor U2550 (N_2550,N_2209,N_2236);
and U2551 (N_2551,N_2282,N_2253);
nand U2552 (N_2552,N_2295,N_2304);
nor U2553 (N_2553,N_2220,N_2316);
nor U2554 (N_2554,N_2251,N_2280);
nor U2555 (N_2555,N_2374,N_2359);
and U2556 (N_2556,N_2321,N_2297);
or U2557 (N_2557,N_2277,N_2259);
nand U2558 (N_2558,N_2251,N_2266);
nor U2559 (N_2559,N_2238,N_2326);
or U2560 (N_2560,N_2378,N_2331);
xor U2561 (N_2561,N_2395,N_2216);
nand U2562 (N_2562,N_2358,N_2284);
nor U2563 (N_2563,N_2323,N_2367);
and U2564 (N_2564,N_2234,N_2388);
nand U2565 (N_2565,N_2316,N_2364);
nand U2566 (N_2566,N_2255,N_2281);
nand U2567 (N_2567,N_2298,N_2336);
nand U2568 (N_2568,N_2289,N_2281);
or U2569 (N_2569,N_2201,N_2243);
nor U2570 (N_2570,N_2204,N_2398);
nand U2571 (N_2571,N_2237,N_2264);
and U2572 (N_2572,N_2222,N_2379);
or U2573 (N_2573,N_2309,N_2334);
and U2574 (N_2574,N_2289,N_2200);
xor U2575 (N_2575,N_2381,N_2242);
and U2576 (N_2576,N_2261,N_2208);
nor U2577 (N_2577,N_2344,N_2366);
and U2578 (N_2578,N_2365,N_2316);
or U2579 (N_2579,N_2204,N_2311);
xor U2580 (N_2580,N_2359,N_2211);
or U2581 (N_2581,N_2271,N_2292);
xnor U2582 (N_2582,N_2339,N_2311);
nand U2583 (N_2583,N_2365,N_2392);
nor U2584 (N_2584,N_2272,N_2282);
and U2585 (N_2585,N_2395,N_2324);
xnor U2586 (N_2586,N_2288,N_2329);
or U2587 (N_2587,N_2354,N_2366);
nor U2588 (N_2588,N_2393,N_2273);
nor U2589 (N_2589,N_2393,N_2358);
nand U2590 (N_2590,N_2359,N_2226);
nand U2591 (N_2591,N_2393,N_2361);
nand U2592 (N_2592,N_2285,N_2368);
and U2593 (N_2593,N_2276,N_2312);
nand U2594 (N_2594,N_2217,N_2328);
or U2595 (N_2595,N_2207,N_2351);
or U2596 (N_2596,N_2319,N_2223);
or U2597 (N_2597,N_2324,N_2242);
and U2598 (N_2598,N_2321,N_2206);
and U2599 (N_2599,N_2202,N_2397);
xor U2600 (N_2600,N_2481,N_2504);
xnor U2601 (N_2601,N_2598,N_2484);
nand U2602 (N_2602,N_2577,N_2459);
or U2603 (N_2603,N_2582,N_2525);
or U2604 (N_2604,N_2578,N_2559);
or U2605 (N_2605,N_2547,N_2439);
or U2606 (N_2606,N_2461,N_2499);
nand U2607 (N_2607,N_2520,N_2572);
or U2608 (N_2608,N_2514,N_2566);
or U2609 (N_2609,N_2418,N_2509);
nor U2610 (N_2610,N_2546,N_2553);
and U2611 (N_2611,N_2543,N_2466);
nor U2612 (N_2612,N_2527,N_2446);
nand U2613 (N_2613,N_2528,N_2417);
nand U2614 (N_2614,N_2469,N_2497);
or U2615 (N_2615,N_2565,N_2567);
or U2616 (N_2616,N_2533,N_2545);
nor U2617 (N_2617,N_2452,N_2456);
and U2618 (N_2618,N_2523,N_2573);
nor U2619 (N_2619,N_2472,N_2536);
nand U2620 (N_2620,N_2590,N_2453);
and U2621 (N_2621,N_2587,N_2447);
and U2622 (N_2622,N_2562,N_2425);
or U2623 (N_2623,N_2548,N_2423);
and U2624 (N_2624,N_2480,N_2414);
nand U2625 (N_2625,N_2554,N_2597);
nor U2626 (N_2626,N_2463,N_2556);
or U2627 (N_2627,N_2415,N_2529);
nor U2628 (N_2628,N_2460,N_2451);
and U2629 (N_2629,N_2454,N_2450);
or U2630 (N_2630,N_2494,N_2437);
nand U2631 (N_2631,N_2549,N_2405);
nand U2632 (N_2632,N_2441,N_2436);
and U2633 (N_2633,N_2524,N_2516);
or U2634 (N_2634,N_2487,N_2531);
nor U2635 (N_2635,N_2448,N_2455);
or U2636 (N_2636,N_2498,N_2443);
nand U2637 (N_2637,N_2408,N_2535);
xor U2638 (N_2638,N_2584,N_2512);
nand U2639 (N_2639,N_2478,N_2403);
nand U2640 (N_2640,N_2581,N_2552);
xnor U2641 (N_2641,N_2506,N_2410);
and U2642 (N_2642,N_2489,N_2541);
or U2643 (N_2643,N_2579,N_2493);
nand U2644 (N_2644,N_2558,N_2402);
nand U2645 (N_2645,N_2444,N_2409);
nand U2646 (N_2646,N_2411,N_2477);
nand U2647 (N_2647,N_2490,N_2530);
and U2648 (N_2648,N_2589,N_2534);
nor U2649 (N_2649,N_2413,N_2511);
and U2650 (N_2650,N_2569,N_2505);
nand U2651 (N_2651,N_2518,N_2500);
nor U2652 (N_2652,N_2420,N_2592);
and U2653 (N_2653,N_2485,N_2571);
nor U2654 (N_2654,N_2432,N_2429);
nor U2655 (N_2655,N_2501,N_2431);
nand U2656 (N_2656,N_2464,N_2519);
or U2657 (N_2657,N_2570,N_2449);
xnor U2658 (N_2658,N_2517,N_2526);
and U2659 (N_2659,N_2532,N_2422);
nor U2660 (N_2660,N_2557,N_2407);
or U2661 (N_2661,N_2561,N_2435);
or U2662 (N_2662,N_2496,N_2424);
nor U2663 (N_2663,N_2465,N_2588);
nor U2664 (N_2664,N_2521,N_2538);
or U2665 (N_2665,N_2555,N_2428);
or U2666 (N_2666,N_2438,N_2475);
and U2667 (N_2667,N_2599,N_2593);
or U2668 (N_2668,N_2551,N_2585);
xnor U2669 (N_2669,N_2482,N_2430);
nor U2670 (N_2670,N_2476,N_2586);
or U2671 (N_2671,N_2495,N_2479);
or U2672 (N_2672,N_2419,N_2522);
or U2673 (N_2673,N_2486,N_2560);
and U2674 (N_2674,N_2537,N_2404);
and U2675 (N_2675,N_2542,N_2483);
or U2676 (N_2676,N_2491,N_2594);
nor U2677 (N_2677,N_2440,N_2433);
nor U2678 (N_2678,N_2462,N_2507);
nand U2679 (N_2679,N_2458,N_2539);
and U2680 (N_2680,N_2544,N_2583);
nor U2681 (N_2681,N_2401,N_2427);
or U2682 (N_2682,N_2492,N_2503);
nand U2683 (N_2683,N_2457,N_2591);
nand U2684 (N_2684,N_2471,N_2468);
and U2685 (N_2685,N_2595,N_2574);
nand U2686 (N_2686,N_2575,N_2406);
or U2687 (N_2687,N_2473,N_2474);
or U2688 (N_2688,N_2564,N_2596);
xor U2689 (N_2689,N_2515,N_2502);
and U2690 (N_2690,N_2426,N_2488);
nor U2691 (N_2691,N_2416,N_2467);
xnor U2692 (N_2692,N_2445,N_2412);
or U2693 (N_2693,N_2442,N_2421);
and U2694 (N_2694,N_2550,N_2400);
and U2695 (N_2695,N_2513,N_2470);
nor U2696 (N_2696,N_2540,N_2510);
nand U2697 (N_2697,N_2508,N_2580);
nor U2698 (N_2698,N_2568,N_2434);
and U2699 (N_2699,N_2576,N_2563);
nand U2700 (N_2700,N_2472,N_2436);
nor U2701 (N_2701,N_2498,N_2414);
or U2702 (N_2702,N_2523,N_2496);
or U2703 (N_2703,N_2546,N_2458);
or U2704 (N_2704,N_2572,N_2444);
and U2705 (N_2705,N_2594,N_2587);
or U2706 (N_2706,N_2547,N_2513);
and U2707 (N_2707,N_2553,N_2557);
or U2708 (N_2708,N_2413,N_2434);
nor U2709 (N_2709,N_2573,N_2529);
or U2710 (N_2710,N_2509,N_2521);
and U2711 (N_2711,N_2599,N_2428);
and U2712 (N_2712,N_2496,N_2430);
or U2713 (N_2713,N_2593,N_2424);
nand U2714 (N_2714,N_2425,N_2511);
or U2715 (N_2715,N_2571,N_2596);
nand U2716 (N_2716,N_2585,N_2440);
or U2717 (N_2717,N_2487,N_2486);
nor U2718 (N_2718,N_2529,N_2597);
and U2719 (N_2719,N_2568,N_2446);
and U2720 (N_2720,N_2462,N_2526);
and U2721 (N_2721,N_2537,N_2555);
and U2722 (N_2722,N_2534,N_2596);
nor U2723 (N_2723,N_2434,N_2479);
nor U2724 (N_2724,N_2471,N_2424);
nor U2725 (N_2725,N_2479,N_2534);
or U2726 (N_2726,N_2560,N_2400);
nor U2727 (N_2727,N_2482,N_2559);
xnor U2728 (N_2728,N_2500,N_2481);
nor U2729 (N_2729,N_2537,N_2562);
and U2730 (N_2730,N_2572,N_2457);
nor U2731 (N_2731,N_2482,N_2578);
xnor U2732 (N_2732,N_2404,N_2478);
and U2733 (N_2733,N_2543,N_2582);
nor U2734 (N_2734,N_2421,N_2464);
nor U2735 (N_2735,N_2578,N_2573);
nand U2736 (N_2736,N_2530,N_2486);
or U2737 (N_2737,N_2411,N_2516);
nor U2738 (N_2738,N_2460,N_2400);
nor U2739 (N_2739,N_2527,N_2444);
or U2740 (N_2740,N_2414,N_2532);
nor U2741 (N_2741,N_2432,N_2537);
and U2742 (N_2742,N_2513,N_2497);
or U2743 (N_2743,N_2424,N_2546);
nor U2744 (N_2744,N_2598,N_2517);
or U2745 (N_2745,N_2511,N_2438);
nor U2746 (N_2746,N_2469,N_2437);
and U2747 (N_2747,N_2553,N_2472);
or U2748 (N_2748,N_2455,N_2599);
xnor U2749 (N_2749,N_2563,N_2545);
nor U2750 (N_2750,N_2419,N_2584);
and U2751 (N_2751,N_2556,N_2488);
nor U2752 (N_2752,N_2448,N_2562);
or U2753 (N_2753,N_2571,N_2569);
nor U2754 (N_2754,N_2559,N_2550);
nor U2755 (N_2755,N_2535,N_2572);
nor U2756 (N_2756,N_2587,N_2423);
and U2757 (N_2757,N_2574,N_2498);
nor U2758 (N_2758,N_2476,N_2428);
or U2759 (N_2759,N_2498,N_2476);
nand U2760 (N_2760,N_2532,N_2572);
or U2761 (N_2761,N_2511,N_2560);
and U2762 (N_2762,N_2434,N_2405);
nor U2763 (N_2763,N_2584,N_2516);
nor U2764 (N_2764,N_2463,N_2416);
nor U2765 (N_2765,N_2584,N_2434);
and U2766 (N_2766,N_2524,N_2434);
or U2767 (N_2767,N_2498,N_2553);
or U2768 (N_2768,N_2472,N_2422);
and U2769 (N_2769,N_2559,N_2529);
nand U2770 (N_2770,N_2454,N_2462);
or U2771 (N_2771,N_2528,N_2502);
xnor U2772 (N_2772,N_2428,N_2407);
nand U2773 (N_2773,N_2568,N_2404);
xnor U2774 (N_2774,N_2558,N_2424);
or U2775 (N_2775,N_2467,N_2435);
nand U2776 (N_2776,N_2404,N_2587);
nor U2777 (N_2777,N_2534,N_2483);
xor U2778 (N_2778,N_2472,N_2479);
and U2779 (N_2779,N_2529,N_2503);
nand U2780 (N_2780,N_2477,N_2584);
or U2781 (N_2781,N_2523,N_2403);
and U2782 (N_2782,N_2516,N_2485);
nor U2783 (N_2783,N_2568,N_2481);
or U2784 (N_2784,N_2593,N_2586);
or U2785 (N_2785,N_2596,N_2435);
xor U2786 (N_2786,N_2497,N_2572);
xnor U2787 (N_2787,N_2423,N_2546);
nand U2788 (N_2788,N_2421,N_2504);
nand U2789 (N_2789,N_2421,N_2536);
nand U2790 (N_2790,N_2431,N_2536);
nand U2791 (N_2791,N_2455,N_2522);
xor U2792 (N_2792,N_2554,N_2457);
nor U2793 (N_2793,N_2528,N_2514);
nor U2794 (N_2794,N_2490,N_2533);
nand U2795 (N_2795,N_2581,N_2509);
or U2796 (N_2796,N_2485,N_2542);
xor U2797 (N_2797,N_2465,N_2470);
nor U2798 (N_2798,N_2563,N_2488);
or U2799 (N_2799,N_2440,N_2499);
nand U2800 (N_2800,N_2796,N_2606);
nand U2801 (N_2801,N_2626,N_2716);
or U2802 (N_2802,N_2790,N_2718);
nor U2803 (N_2803,N_2689,N_2633);
and U2804 (N_2804,N_2726,N_2763);
or U2805 (N_2805,N_2745,N_2685);
nand U2806 (N_2806,N_2672,N_2659);
or U2807 (N_2807,N_2688,N_2629);
nor U2808 (N_2808,N_2694,N_2671);
and U2809 (N_2809,N_2732,N_2656);
nand U2810 (N_2810,N_2620,N_2644);
and U2811 (N_2811,N_2752,N_2622);
nor U2812 (N_2812,N_2693,N_2768);
or U2813 (N_2813,N_2653,N_2612);
and U2814 (N_2814,N_2794,N_2687);
xor U2815 (N_2815,N_2727,N_2733);
or U2816 (N_2816,N_2657,N_2686);
nor U2817 (N_2817,N_2711,N_2757);
nor U2818 (N_2818,N_2791,N_2634);
nand U2819 (N_2819,N_2746,N_2788);
xor U2820 (N_2820,N_2611,N_2616);
or U2821 (N_2821,N_2737,N_2731);
or U2822 (N_2822,N_2738,N_2661);
nand U2823 (N_2823,N_2628,N_2713);
and U2824 (N_2824,N_2720,N_2690);
and U2825 (N_2825,N_2742,N_2639);
and U2826 (N_2826,N_2717,N_2775);
and U2827 (N_2827,N_2723,N_2674);
nor U2828 (N_2828,N_2780,N_2765);
and U2829 (N_2829,N_2664,N_2662);
and U2830 (N_2830,N_2762,N_2767);
or U2831 (N_2831,N_2744,N_2692);
nor U2832 (N_2832,N_2701,N_2728);
or U2833 (N_2833,N_2614,N_2630);
nand U2834 (N_2834,N_2709,N_2755);
nor U2835 (N_2835,N_2681,N_2778);
or U2836 (N_2836,N_2605,N_2797);
nand U2837 (N_2837,N_2640,N_2787);
nor U2838 (N_2838,N_2624,N_2785);
and U2839 (N_2839,N_2714,N_2617);
nand U2840 (N_2840,N_2725,N_2679);
nand U2841 (N_2841,N_2627,N_2772);
or U2842 (N_2842,N_2750,N_2771);
and U2843 (N_2843,N_2719,N_2710);
or U2844 (N_2844,N_2631,N_2676);
nor U2845 (N_2845,N_2669,N_2609);
and U2846 (N_2846,N_2654,N_2702);
and U2847 (N_2847,N_2641,N_2670);
or U2848 (N_2848,N_2683,N_2766);
or U2849 (N_2849,N_2708,N_2740);
and U2850 (N_2850,N_2667,N_2779);
xor U2851 (N_2851,N_2721,N_2781);
nor U2852 (N_2852,N_2696,N_2715);
nor U2853 (N_2853,N_2646,N_2608);
or U2854 (N_2854,N_2795,N_2600);
xnor U2855 (N_2855,N_2743,N_2700);
xor U2856 (N_2856,N_2623,N_2649);
and U2857 (N_2857,N_2603,N_2632);
xor U2858 (N_2858,N_2789,N_2610);
or U2859 (N_2859,N_2776,N_2741);
and U2860 (N_2860,N_2777,N_2663);
nor U2861 (N_2861,N_2784,N_2799);
nor U2862 (N_2862,N_2658,N_2758);
nor U2863 (N_2863,N_2770,N_2783);
nand U2864 (N_2864,N_2734,N_2735);
or U2865 (N_2865,N_2602,N_2673);
xor U2866 (N_2866,N_2613,N_2650);
or U2867 (N_2867,N_2707,N_2645);
and U2868 (N_2868,N_2764,N_2792);
or U2869 (N_2869,N_2643,N_2722);
and U2870 (N_2870,N_2793,N_2642);
nor U2871 (N_2871,N_2668,N_2655);
and U2872 (N_2872,N_2601,N_2782);
and U2873 (N_2873,N_2698,N_2625);
xor U2874 (N_2874,N_2703,N_2604);
or U2875 (N_2875,N_2736,N_2635);
or U2876 (N_2876,N_2619,N_2695);
nor U2877 (N_2877,N_2724,N_2647);
and U2878 (N_2878,N_2749,N_2712);
and U2879 (N_2879,N_2730,N_2621);
nand U2880 (N_2880,N_2675,N_2748);
and U2881 (N_2881,N_2747,N_2773);
nand U2882 (N_2882,N_2618,N_2705);
or U2883 (N_2883,N_2729,N_2678);
or U2884 (N_2884,N_2697,N_2680);
nor U2885 (N_2885,N_2665,N_2739);
xor U2886 (N_2886,N_2706,N_2677);
or U2887 (N_2887,N_2652,N_2638);
nor U2888 (N_2888,N_2753,N_2666);
nor U2889 (N_2889,N_2704,N_2636);
nand U2890 (N_2890,N_2637,N_2751);
nor U2891 (N_2891,N_2760,N_2615);
nor U2892 (N_2892,N_2769,N_2607);
nand U2893 (N_2893,N_2651,N_2660);
and U2894 (N_2894,N_2684,N_2798);
and U2895 (N_2895,N_2691,N_2682);
nor U2896 (N_2896,N_2648,N_2754);
nor U2897 (N_2897,N_2761,N_2756);
and U2898 (N_2898,N_2774,N_2699);
or U2899 (N_2899,N_2786,N_2759);
or U2900 (N_2900,N_2790,N_2710);
or U2901 (N_2901,N_2614,N_2741);
nor U2902 (N_2902,N_2749,N_2651);
and U2903 (N_2903,N_2691,N_2786);
nor U2904 (N_2904,N_2778,N_2745);
or U2905 (N_2905,N_2613,N_2780);
or U2906 (N_2906,N_2626,N_2744);
xor U2907 (N_2907,N_2793,N_2627);
and U2908 (N_2908,N_2601,N_2605);
and U2909 (N_2909,N_2611,N_2658);
nor U2910 (N_2910,N_2605,N_2708);
or U2911 (N_2911,N_2665,N_2677);
and U2912 (N_2912,N_2667,N_2712);
nand U2913 (N_2913,N_2657,N_2600);
xnor U2914 (N_2914,N_2674,N_2644);
xor U2915 (N_2915,N_2689,N_2781);
nor U2916 (N_2916,N_2785,N_2758);
nor U2917 (N_2917,N_2710,N_2671);
nand U2918 (N_2918,N_2605,N_2667);
or U2919 (N_2919,N_2649,N_2706);
and U2920 (N_2920,N_2670,N_2733);
or U2921 (N_2921,N_2743,N_2739);
nand U2922 (N_2922,N_2760,N_2612);
nand U2923 (N_2923,N_2649,N_2682);
nor U2924 (N_2924,N_2756,N_2730);
nand U2925 (N_2925,N_2718,N_2611);
nor U2926 (N_2926,N_2677,N_2730);
and U2927 (N_2927,N_2602,N_2649);
or U2928 (N_2928,N_2663,N_2684);
and U2929 (N_2929,N_2701,N_2608);
or U2930 (N_2930,N_2694,N_2723);
xnor U2931 (N_2931,N_2685,N_2782);
xor U2932 (N_2932,N_2697,N_2780);
xor U2933 (N_2933,N_2745,N_2640);
nor U2934 (N_2934,N_2768,N_2769);
and U2935 (N_2935,N_2797,N_2668);
and U2936 (N_2936,N_2700,N_2611);
or U2937 (N_2937,N_2718,N_2702);
nor U2938 (N_2938,N_2623,N_2657);
or U2939 (N_2939,N_2603,N_2625);
or U2940 (N_2940,N_2690,N_2732);
or U2941 (N_2941,N_2737,N_2658);
xnor U2942 (N_2942,N_2717,N_2628);
and U2943 (N_2943,N_2619,N_2721);
nor U2944 (N_2944,N_2742,N_2618);
and U2945 (N_2945,N_2731,N_2743);
nand U2946 (N_2946,N_2617,N_2797);
or U2947 (N_2947,N_2768,N_2705);
xor U2948 (N_2948,N_2724,N_2785);
nor U2949 (N_2949,N_2770,N_2637);
and U2950 (N_2950,N_2669,N_2618);
and U2951 (N_2951,N_2729,N_2721);
and U2952 (N_2952,N_2683,N_2743);
xor U2953 (N_2953,N_2663,N_2673);
nand U2954 (N_2954,N_2766,N_2645);
nor U2955 (N_2955,N_2677,N_2718);
or U2956 (N_2956,N_2790,N_2704);
or U2957 (N_2957,N_2650,N_2646);
nor U2958 (N_2958,N_2701,N_2624);
nand U2959 (N_2959,N_2757,N_2639);
and U2960 (N_2960,N_2770,N_2714);
or U2961 (N_2961,N_2693,N_2645);
and U2962 (N_2962,N_2634,N_2758);
nand U2963 (N_2963,N_2774,N_2614);
or U2964 (N_2964,N_2662,N_2673);
nand U2965 (N_2965,N_2743,N_2668);
nor U2966 (N_2966,N_2700,N_2739);
and U2967 (N_2967,N_2779,N_2608);
xor U2968 (N_2968,N_2612,N_2714);
nor U2969 (N_2969,N_2721,N_2674);
nor U2970 (N_2970,N_2718,N_2606);
nand U2971 (N_2971,N_2661,N_2705);
xor U2972 (N_2972,N_2658,N_2689);
or U2973 (N_2973,N_2765,N_2637);
and U2974 (N_2974,N_2723,N_2785);
and U2975 (N_2975,N_2643,N_2682);
nand U2976 (N_2976,N_2780,N_2628);
or U2977 (N_2977,N_2776,N_2660);
or U2978 (N_2978,N_2704,N_2702);
nand U2979 (N_2979,N_2758,N_2685);
or U2980 (N_2980,N_2752,N_2745);
nor U2981 (N_2981,N_2627,N_2647);
nor U2982 (N_2982,N_2798,N_2796);
and U2983 (N_2983,N_2753,N_2689);
and U2984 (N_2984,N_2687,N_2655);
nand U2985 (N_2985,N_2713,N_2796);
and U2986 (N_2986,N_2774,N_2796);
xor U2987 (N_2987,N_2710,N_2722);
and U2988 (N_2988,N_2648,N_2788);
xor U2989 (N_2989,N_2775,N_2744);
nand U2990 (N_2990,N_2625,N_2761);
or U2991 (N_2991,N_2700,N_2692);
xnor U2992 (N_2992,N_2715,N_2746);
xnor U2993 (N_2993,N_2779,N_2677);
xor U2994 (N_2994,N_2785,N_2657);
and U2995 (N_2995,N_2753,N_2735);
or U2996 (N_2996,N_2754,N_2770);
or U2997 (N_2997,N_2621,N_2648);
or U2998 (N_2998,N_2799,N_2620);
and U2999 (N_2999,N_2608,N_2778);
xor U3000 (N_3000,N_2974,N_2976);
or U3001 (N_3001,N_2902,N_2893);
nand U3002 (N_3002,N_2815,N_2954);
and U3003 (N_3003,N_2844,N_2997);
nand U3004 (N_3004,N_2991,N_2874);
nor U3005 (N_3005,N_2956,N_2900);
xor U3006 (N_3006,N_2803,N_2988);
nand U3007 (N_3007,N_2965,N_2901);
and U3008 (N_3008,N_2957,N_2802);
nor U3009 (N_3009,N_2964,N_2853);
nor U3010 (N_3010,N_2973,N_2841);
nor U3011 (N_3011,N_2951,N_2903);
and U3012 (N_3012,N_2994,N_2938);
and U3013 (N_3013,N_2854,N_2940);
or U3014 (N_3014,N_2896,N_2935);
nor U3015 (N_3015,N_2837,N_2870);
xnor U3016 (N_3016,N_2818,N_2831);
or U3017 (N_3017,N_2967,N_2961);
or U3018 (N_3018,N_2911,N_2999);
nand U3019 (N_3019,N_2924,N_2933);
and U3020 (N_3020,N_2929,N_2848);
nand U3021 (N_3021,N_2958,N_2811);
or U3022 (N_3022,N_2836,N_2871);
or U3023 (N_3023,N_2814,N_2858);
and U3024 (N_3024,N_2895,N_2998);
xnor U3025 (N_3025,N_2812,N_2863);
and U3026 (N_3026,N_2907,N_2877);
or U3027 (N_3027,N_2806,N_2852);
or U3028 (N_3028,N_2857,N_2805);
nand U3029 (N_3029,N_2913,N_2916);
or U3030 (N_3030,N_2977,N_2843);
and U3031 (N_3031,N_2982,N_2910);
nand U3032 (N_3032,N_2834,N_2948);
or U3033 (N_3033,N_2838,N_2971);
or U3034 (N_3034,N_2921,N_2828);
nor U3035 (N_3035,N_2904,N_2840);
nor U3036 (N_3036,N_2936,N_2914);
and U3037 (N_3037,N_2810,N_2939);
or U3038 (N_3038,N_2882,N_2846);
nor U3039 (N_3039,N_2917,N_2866);
nand U3040 (N_3040,N_2920,N_2931);
nor U3041 (N_3041,N_2968,N_2885);
and U3042 (N_3042,N_2829,N_2868);
nor U3043 (N_3043,N_2962,N_2861);
nand U3044 (N_3044,N_2819,N_2970);
or U3045 (N_3045,N_2930,N_2922);
nand U3046 (N_3046,N_2884,N_2889);
nor U3047 (N_3047,N_2851,N_2947);
nand U3048 (N_3048,N_2946,N_2850);
nor U3049 (N_3049,N_2941,N_2950);
and U3050 (N_3050,N_2963,N_2886);
nand U3051 (N_3051,N_2942,N_2925);
nand U3052 (N_3052,N_2827,N_2821);
and U3053 (N_3053,N_2881,N_2880);
or U3054 (N_3054,N_2989,N_2912);
and U3055 (N_3055,N_2992,N_2807);
nor U3056 (N_3056,N_2926,N_2820);
nand U3057 (N_3057,N_2944,N_2856);
nand U3058 (N_3058,N_2873,N_2869);
nand U3059 (N_3059,N_2979,N_2978);
nor U3060 (N_3060,N_2878,N_2928);
nor U3061 (N_3061,N_2980,N_2876);
nand U3062 (N_3062,N_2859,N_2823);
or U3063 (N_3063,N_2960,N_2809);
xor U3064 (N_3064,N_2919,N_2953);
nand U3065 (N_3065,N_2855,N_2832);
and U3066 (N_3066,N_2845,N_2879);
nor U3067 (N_3067,N_2892,N_2993);
and U3068 (N_3068,N_2996,N_2891);
nor U3069 (N_3069,N_2972,N_2934);
xnor U3070 (N_3070,N_2865,N_2937);
or U3071 (N_3071,N_2883,N_2955);
and U3072 (N_3072,N_2987,N_2932);
or U3073 (N_3073,N_2986,N_2824);
nor U3074 (N_3074,N_2872,N_2890);
nor U3075 (N_3075,N_2830,N_2813);
and U3076 (N_3076,N_2816,N_2990);
xor U3077 (N_3077,N_2835,N_2898);
or U3078 (N_3078,N_2905,N_2804);
xnor U3079 (N_3079,N_2817,N_2995);
or U3080 (N_3080,N_2867,N_2949);
and U3081 (N_3081,N_2899,N_2808);
and U3082 (N_3082,N_2918,N_2826);
and U3083 (N_3083,N_2887,N_2945);
and U3084 (N_3084,N_2822,N_2966);
xor U3085 (N_3085,N_2842,N_2864);
nand U3086 (N_3086,N_2943,N_2862);
or U3087 (N_3087,N_2897,N_2860);
and U3088 (N_3088,N_2894,N_2915);
and U3089 (N_3089,N_2927,N_2952);
nand U3090 (N_3090,N_2923,N_2825);
or U3091 (N_3091,N_2985,N_2909);
nor U3092 (N_3092,N_2906,N_2984);
nor U3093 (N_3093,N_2888,N_2975);
nand U3094 (N_3094,N_2875,N_2983);
or U3095 (N_3095,N_2959,N_2969);
or U3096 (N_3096,N_2849,N_2839);
nor U3097 (N_3097,N_2833,N_2908);
nor U3098 (N_3098,N_2800,N_2801);
nor U3099 (N_3099,N_2981,N_2847);
nand U3100 (N_3100,N_2963,N_2925);
nand U3101 (N_3101,N_2824,N_2924);
nand U3102 (N_3102,N_2804,N_2989);
nand U3103 (N_3103,N_2947,N_2852);
nand U3104 (N_3104,N_2943,N_2814);
or U3105 (N_3105,N_2978,N_2969);
or U3106 (N_3106,N_2845,N_2805);
nor U3107 (N_3107,N_2979,N_2848);
nand U3108 (N_3108,N_2985,N_2959);
nand U3109 (N_3109,N_2866,N_2881);
or U3110 (N_3110,N_2849,N_2891);
or U3111 (N_3111,N_2874,N_2935);
or U3112 (N_3112,N_2961,N_2868);
nor U3113 (N_3113,N_2938,N_2919);
or U3114 (N_3114,N_2833,N_2887);
nor U3115 (N_3115,N_2969,N_2882);
nor U3116 (N_3116,N_2854,N_2957);
or U3117 (N_3117,N_2869,N_2899);
or U3118 (N_3118,N_2978,N_2955);
xor U3119 (N_3119,N_2985,N_2807);
or U3120 (N_3120,N_2975,N_2822);
or U3121 (N_3121,N_2988,N_2805);
or U3122 (N_3122,N_2825,N_2826);
nor U3123 (N_3123,N_2907,N_2912);
nand U3124 (N_3124,N_2981,N_2800);
or U3125 (N_3125,N_2832,N_2883);
or U3126 (N_3126,N_2950,N_2850);
nand U3127 (N_3127,N_2951,N_2813);
and U3128 (N_3128,N_2891,N_2883);
nor U3129 (N_3129,N_2849,N_2930);
nor U3130 (N_3130,N_2828,N_2942);
xor U3131 (N_3131,N_2925,N_2885);
and U3132 (N_3132,N_2925,N_2900);
or U3133 (N_3133,N_2901,N_2933);
or U3134 (N_3134,N_2989,N_2959);
nor U3135 (N_3135,N_2956,N_2935);
and U3136 (N_3136,N_2896,N_2901);
or U3137 (N_3137,N_2845,N_2844);
xnor U3138 (N_3138,N_2885,N_2819);
and U3139 (N_3139,N_2925,N_2984);
and U3140 (N_3140,N_2829,N_2987);
nor U3141 (N_3141,N_2868,N_2860);
nand U3142 (N_3142,N_2820,N_2950);
and U3143 (N_3143,N_2895,N_2959);
and U3144 (N_3144,N_2958,N_2918);
xor U3145 (N_3145,N_2842,N_2913);
nor U3146 (N_3146,N_2938,N_2872);
or U3147 (N_3147,N_2926,N_2936);
and U3148 (N_3148,N_2863,N_2931);
nor U3149 (N_3149,N_2947,N_2878);
xnor U3150 (N_3150,N_2954,N_2936);
and U3151 (N_3151,N_2871,N_2825);
and U3152 (N_3152,N_2958,N_2926);
nor U3153 (N_3153,N_2985,N_2952);
or U3154 (N_3154,N_2852,N_2835);
or U3155 (N_3155,N_2878,N_2872);
and U3156 (N_3156,N_2874,N_2878);
and U3157 (N_3157,N_2971,N_2954);
xor U3158 (N_3158,N_2803,N_2895);
nand U3159 (N_3159,N_2909,N_2834);
xnor U3160 (N_3160,N_2844,N_2926);
nand U3161 (N_3161,N_2994,N_2847);
or U3162 (N_3162,N_2845,N_2921);
nand U3163 (N_3163,N_2888,N_2801);
nor U3164 (N_3164,N_2946,N_2858);
nand U3165 (N_3165,N_2967,N_2843);
nor U3166 (N_3166,N_2865,N_2956);
and U3167 (N_3167,N_2853,N_2941);
nand U3168 (N_3168,N_2915,N_2821);
nand U3169 (N_3169,N_2895,N_2826);
or U3170 (N_3170,N_2963,N_2804);
or U3171 (N_3171,N_2846,N_2848);
and U3172 (N_3172,N_2859,N_2999);
nand U3173 (N_3173,N_2997,N_2932);
nand U3174 (N_3174,N_2877,N_2902);
nand U3175 (N_3175,N_2809,N_2875);
or U3176 (N_3176,N_2915,N_2847);
and U3177 (N_3177,N_2999,N_2939);
nor U3178 (N_3178,N_2832,N_2823);
or U3179 (N_3179,N_2872,N_2997);
and U3180 (N_3180,N_2924,N_2885);
nand U3181 (N_3181,N_2872,N_2935);
nand U3182 (N_3182,N_2854,N_2876);
xor U3183 (N_3183,N_2951,N_2958);
nor U3184 (N_3184,N_2838,N_2946);
xor U3185 (N_3185,N_2936,N_2811);
nor U3186 (N_3186,N_2968,N_2977);
or U3187 (N_3187,N_2980,N_2952);
or U3188 (N_3188,N_2955,N_2972);
nand U3189 (N_3189,N_2828,N_2867);
nand U3190 (N_3190,N_2939,N_2910);
xor U3191 (N_3191,N_2848,N_2958);
nor U3192 (N_3192,N_2846,N_2852);
nand U3193 (N_3193,N_2896,N_2868);
xnor U3194 (N_3194,N_2865,N_2867);
nor U3195 (N_3195,N_2928,N_2993);
nand U3196 (N_3196,N_2829,N_2828);
xnor U3197 (N_3197,N_2882,N_2974);
nor U3198 (N_3198,N_2877,N_2813);
and U3199 (N_3199,N_2825,N_2902);
nor U3200 (N_3200,N_3177,N_3117);
and U3201 (N_3201,N_3166,N_3129);
and U3202 (N_3202,N_3079,N_3170);
or U3203 (N_3203,N_3081,N_3151);
nor U3204 (N_3204,N_3152,N_3020);
nor U3205 (N_3205,N_3083,N_3164);
and U3206 (N_3206,N_3054,N_3182);
nand U3207 (N_3207,N_3198,N_3199);
nand U3208 (N_3208,N_3160,N_3140);
nand U3209 (N_3209,N_3141,N_3009);
xor U3210 (N_3210,N_3088,N_3183);
and U3211 (N_3211,N_3090,N_3155);
or U3212 (N_3212,N_3137,N_3100);
xor U3213 (N_3213,N_3189,N_3032);
and U3214 (N_3214,N_3131,N_3018);
and U3215 (N_3215,N_3028,N_3180);
xnor U3216 (N_3216,N_3098,N_3049);
nand U3217 (N_3217,N_3069,N_3135);
or U3218 (N_3218,N_3107,N_3133);
nand U3219 (N_3219,N_3165,N_3070);
or U3220 (N_3220,N_3041,N_3027);
or U3221 (N_3221,N_3138,N_3123);
or U3222 (N_3222,N_3071,N_3019);
nor U3223 (N_3223,N_3063,N_3108);
and U3224 (N_3224,N_3043,N_3175);
nor U3225 (N_3225,N_3021,N_3168);
and U3226 (N_3226,N_3084,N_3091);
and U3227 (N_3227,N_3060,N_3121);
or U3228 (N_3228,N_3147,N_3113);
and U3229 (N_3229,N_3195,N_3044);
and U3230 (N_3230,N_3076,N_3139);
nand U3231 (N_3231,N_3127,N_3013);
or U3232 (N_3232,N_3097,N_3089);
nor U3233 (N_3233,N_3053,N_3184);
nand U3234 (N_3234,N_3185,N_3125);
nand U3235 (N_3235,N_3072,N_3197);
nand U3236 (N_3236,N_3010,N_3030);
or U3237 (N_3237,N_3162,N_3024);
nand U3238 (N_3238,N_3025,N_3048);
nor U3239 (N_3239,N_3156,N_3066);
and U3240 (N_3240,N_3059,N_3033);
and U3241 (N_3241,N_3181,N_3096);
nand U3242 (N_3242,N_3011,N_3057);
nand U3243 (N_3243,N_3051,N_3082);
and U3244 (N_3244,N_3006,N_3154);
and U3245 (N_3245,N_3163,N_3086);
or U3246 (N_3246,N_3075,N_3050);
nand U3247 (N_3247,N_3179,N_3172);
nor U3248 (N_3248,N_3120,N_3102);
nand U3249 (N_3249,N_3146,N_3134);
nand U3250 (N_3250,N_3008,N_3023);
xor U3251 (N_3251,N_3007,N_3012);
or U3252 (N_3252,N_3073,N_3099);
and U3253 (N_3253,N_3029,N_3087);
nand U3254 (N_3254,N_3142,N_3085);
nor U3255 (N_3255,N_3064,N_3035);
nor U3256 (N_3256,N_3103,N_3101);
and U3257 (N_3257,N_3017,N_3000);
or U3258 (N_3258,N_3145,N_3015);
nand U3259 (N_3259,N_3052,N_3148);
and U3260 (N_3260,N_3034,N_3169);
nand U3261 (N_3261,N_3171,N_3161);
or U3262 (N_3262,N_3110,N_3065);
or U3263 (N_3263,N_3105,N_3157);
nand U3264 (N_3264,N_3176,N_3126);
nand U3265 (N_3265,N_3058,N_3014);
xnor U3266 (N_3266,N_3042,N_3038);
and U3267 (N_3267,N_3190,N_3116);
nand U3268 (N_3268,N_3192,N_3132);
nand U3269 (N_3269,N_3111,N_3104);
or U3270 (N_3270,N_3119,N_3095);
and U3271 (N_3271,N_3036,N_3045);
or U3272 (N_3272,N_3040,N_3109);
and U3273 (N_3273,N_3122,N_3136);
nand U3274 (N_3274,N_3055,N_3167);
nand U3275 (N_3275,N_3062,N_3118);
or U3276 (N_3276,N_3143,N_3037);
and U3277 (N_3277,N_3115,N_3068);
and U3278 (N_3278,N_3150,N_3173);
nor U3279 (N_3279,N_3153,N_3067);
or U3280 (N_3280,N_3130,N_3093);
and U3281 (N_3281,N_3078,N_3022);
and U3282 (N_3282,N_3191,N_3002);
nor U3283 (N_3283,N_3128,N_3188);
or U3284 (N_3284,N_3046,N_3106);
and U3285 (N_3285,N_3056,N_3047);
nor U3286 (N_3286,N_3187,N_3186);
or U3287 (N_3287,N_3124,N_3196);
and U3288 (N_3288,N_3016,N_3003);
nor U3289 (N_3289,N_3026,N_3178);
nand U3290 (N_3290,N_3112,N_3193);
nand U3291 (N_3291,N_3114,N_3077);
nand U3292 (N_3292,N_3004,N_3092);
and U3293 (N_3293,N_3159,N_3061);
xor U3294 (N_3294,N_3174,N_3074);
or U3295 (N_3295,N_3031,N_3005);
or U3296 (N_3296,N_3039,N_3194);
nand U3297 (N_3297,N_3094,N_3158);
and U3298 (N_3298,N_3149,N_3144);
or U3299 (N_3299,N_3001,N_3080);
and U3300 (N_3300,N_3020,N_3197);
nand U3301 (N_3301,N_3171,N_3120);
xor U3302 (N_3302,N_3103,N_3048);
or U3303 (N_3303,N_3004,N_3131);
xnor U3304 (N_3304,N_3120,N_3191);
nand U3305 (N_3305,N_3188,N_3124);
nor U3306 (N_3306,N_3115,N_3102);
nor U3307 (N_3307,N_3109,N_3172);
and U3308 (N_3308,N_3184,N_3003);
nand U3309 (N_3309,N_3095,N_3061);
nand U3310 (N_3310,N_3097,N_3166);
nand U3311 (N_3311,N_3042,N_3067);
nand U3312 (N_3312,N_3007,N_3042);
nand U3313 (N_3313,N_3124,N_3182);
and U3314 (N_3314,N_3098,N_3080);
or U3315 (N_3315,N_3153,N_3066);
or U3316 (N_3316,N_3117,N_3059);
nand U3317 (N_3317,N_3089,N_3074);
nand U3318 (N_3318,N_3135,N_3094);
nand U3319 (N_3319,N_3193,N_3119);
nor U3320 (N_3320,N_3115,N_3082);
and U3321 (N_3321,N_3122,N_3057);
nor U3322 (N_3322,N_3135,N_3019);
nor U3323 (N_3323,N_3071,N_3141);
and U3324 (N_3324,N_3168,N_3158);
and U3325 (N_3325,N_3123,N_3114);
or U3326 (N_3326,N_3154,N_3054);
nor U3327 (N_3327,N_3065,N_3106);
or U3328 (N_3328,N_3041,N_3187);
nor U3329 (N_3329,N_3133,N_3051);
nand U3330 (N_3330,N_3064,N_3112);
and U3331 (N_3331,N_3058,N_3077);
and U3332 (N_3332,N_3155,N_3093);
and U3333 (N_3333,N_3099,N_3106);
and U3334 (N_3334,N_3062,N_3169);
nor U3335 (N_3335,N_3165,N_3149);
or U3336 (N_3336,N_3043,N_3082);
or U3337 (N_3337,N_3022,N_3192);
and U3338 (N_3338,N_3025,N_3046);
and U3339 (N_3339,N_3019,N_3109);
or U3340 (N_3340,N_3069,N_3187);
or U3341 (N_3341,N_3087,N_3113);
or U3342 (N_3342,N_3009,N_3020);
nand U3343 (N_3343,N_3195,N_3042);
or U3344 (N_3344,N_3156,N_3055);
nand U3345 (N_3345,N_3160,N_3004);
nor U3346 (N_3346,N_3043,N_3048);
or U3347 (N_3347,N_3066,N_3161);
or U3348 (N_3348,N_3008,N_3085);
nor U3349 (N_3349,N_3092,N_3057);
or U3350 (N_3350,N_3008,N_3001);
or U3351 (N_3351,N_3123,N_3043);
nand U3352 (N_3352,N_3059,N_3178);
nor U3353 (N_3353,N_3175,N_3087);
nor U3354 (N_3354,N_3172,N_3110);
and U3355 (N_3355,N_3144,N_3111);
nand U3356 (N_3356,N_3088,N_3176);
and U3357 (N_3357,N_3071,N_3163);
and U3358 (N_3358,N_3029,N_3080);
or U3359 (N_3359,N_3166,N_3036);
nand U3360 (N_3360,N_3093,N_3196);
nand U3361 (N_3361,N_3118,N_3040);
nand U3362 (N_3362,N_3199,N_3128);
nor U3363 (N_3363,N_3067,N_3114);
nand U3364 (N_3364,N_3165,N_3025);
nand U3365 (N_3365,N_3010,N_3057);
or U3366 (N_3366,N_3079,N_3029);
nor U3367 (N_3367,N_3166,N_3172);
xnor U3368 (N_3368,N_3035,N_3074);
and U3369 (N_3369,N_3107,N_3130);
nand U3370 (N_3370,N_3144,N_3133);
or U3371 (N_3371,N_3080,N_3024);
nand U3372 (N_3372,N_3119,N_3034);
or U3373 (N_3373,N_3091,N_3062);
and U3374 (N_3374,N_3153,N_3148);
nand U3375 (N_3375,N_3002,N_3092);
nor U3376 (N_3376,N_3095,N_3135);
or U3377 (N_3377,N_3067,N_3007);
nand U3378 (N_3378,N_3194,N_3050);
or U3379 (N_3379,N_3133,N_3092);
nand U3380 (N_3380,N_3133,N_3100);
and U3381 (N_3381,N_3115,N_3163);
nand U3382 (N_3382,N_3093,N_3025);
and U3383 (N_3383,N_3003,N_3112);
and U3384 (N_3384,N_3087,N_3172);
or U3385 (N_3385,N_3066,N_3089);
or U3386 (N_3386,N_3029,N_3195);
nand U3387 (N_3387,N_3113,N_3199);
or U3388 (N_3388,N_3016,N_3117);
xor U3389 (N_3389,N_3046,N_3157);
and U3390 (N_3390,N_3104,N_3091);
nand U3391 (N_3391,N_3184,N_3192);
and U3392 (N_3392,N_3147,N_3100);
and U3393 (N_3393,N_3095,N_3151);
xnor U3394 (N_3394,N_3164,N_3017);
or U3395 (N_3395,N_3059,N_3008);
nand U3396 (N_3396,N_3015,N_3122);
or U3397 (N_3397,N_3168,N_3153);
or U3398 (N_3398,N_3120,N_3009);
xnor U3399 (N_3399,N_3040,N_3083);
and U3400 (N_3400,N_3281,N_3265);
nor U3401 (N_3401,N_3344,N_3351);
nand U3402 (N_3402,N_3392,N_3390);
nor U3403 (N_3403,N_3398,N_3228);
or U3404 (N_3404,N_3395,N_3242);
nand U3405 (N_3405,N_3232,N_3379);
nand U3406 (N_3406,N_3310,N_3234);
nor U3407 (N_3407,N_3261,N_3399);
or U3408 (N_3408,N_3313,N_3224);
nor U3409 (N_3409,N_3363,N_3223);
nor U3410 (N_3410,N_3365,N_3356);
xnor U3411 (N_3411,N_3294,N_3255);
and U3412 (N_3412,N_3364,N_3346);
or U3413 (N_3413,N_3316,N_3358);
or U3414 (N_3414,N_3256,N_3247);
xnor U3415 (N_3415,N_3250,N_3216);
or U3416 (N_3416,N_3241,N_3201);
and U3417 (N_3417,N_3374,N_3293);
nand U3418 (N_3418,N_3245,N_3209);
and U3419 (N_3419,N_3291,N_3384);
or U3420 (N_3420,N_3371,N_3299);
nor U3421 (N_3421,N_3202,N_3280);
and U3422 (N_3422,N_3325,N_3377);
nand U3423 (N_3423,N_3345,N_3264);
xnor U3424 (N_3424,N_3215,N_3305);
or U3425 (N_3425,N_3376,N_3372);
or U3426 (N_3426,N_3211,N_3394);
nor U3427 (N_3427,N_3360,N_3295);
xor U3428 (N_3428,N_3320,N_3221);
and U3429 (N_3429,N_3318,N_3375);
nand U3430 (N_3430,N_3230,N_3240);
nor U3431 (N_3431,N_3200,N_3322);
nor U3432 (N_3432,N_3288,N_3220);
nor U3433 (N_3433,N_3324,N_3270);
nand U3434 (N_3434,N_3350,N_3336);
and U3435 (N_3435,N_3297,N_3301);
xor U3436 (N_3436,N_3206,N_3355);
nand U3437 (N_3437,N_3269,N_3319);
nand U3438 (N_3438,N_3210,N_3385);
nor U3439 (N_3439,N_3370,N_3396);
and U3440 (N_3440,N_3382,N_3335);
and U3441 (N_3441,N_3284,N_3208);
or U3442 (N_3442,N_3323,N_3233);
nor U3443 (N_3443,N_3257,N_3378);
and U3444 (N_3444,N_3326,N_3267);
nor U3445 (N_3445,N_3292,N_3286);
nor U3446 (N_3446,N_3219,N_3283);
or U3447 (N_3447,N_3312,N_3214);
or U3448 (N_3448,N_3359,N_3285);
or U3449 (N_3449,N_3268,N_3327);
and U3450 (N_3450,N_3338,N_3321);
or U3451 (N_3451,N_3304,N_3388);
nand U3452 (N_3452,N_3254,N_3306);
and U3453 (N_3453,N_3236,N_3258);
nand U3454 (N_3454,N_3217,N_3341);
nand U3455 (N_3455,N_3354,N_3290);
nand U3456 (N_3456,N_3275,N_3383);
nor U3457 (N_3457,N_3277,N_3315);
nor U3458 (N_3458,N_3347,N_3243);
and U3459 (N_3459,N_3203,N_3337);
nand U3460 (N_3460,N_3252,N_3328);
or U3461 (N_3461,N_3367,N_3366);
nand U3462 (N_3462,N_3357,N_3259);
and U3463 (N_3463,N_3333,N_3373);
nand U3464 (N_3464,N_3266,N_3368);
and U3465 (N_3465,N_3207,N_3239);
nand U3466 (N_3466,N_3263,N_3246);
and U3467 (N_3467,N_3272,N_3340);
and U3468 (N_3468,N_3262,N_3225);
and U3469 (N_3469,N_3279,N_3317);
nor U3470 (N_3470,N_3229,N_3342);
xnor U3471 (N_3471,N_3330,N_3353);
nor U3472 (N_3472,N_3289,N_3300);
and U3473 (N_3473,N_3352,N_3361);
nand U3474 (N_3474,N_3362,N_3311);
nor U3475 (N_3475,N_3296,N_3222);
or U3476 (N_3476,N_3231,N_3282);
nor U3477 (N_3477,N_3393,N_3397);
or U3478 (N_3478,N_3212,N_3307);
and U3479 (N_3479,N_3235,N_3278);
nor U3480 (N_3480,N_3237,N_3389);
or U3481 (N_3481,N_3331,N_3339);
xor U3482 (N_3482,N_3276,N_3303);
nor U3483 (N_3483,N_3332,N_3227);
or U3484 (N_3484,N_3329,N_3308);
and U3485 (N_3485,N_3314,N_3387);
nand U3486 (N_3486,N_3380,N_3213);
and U3487 (N_3487,N_3244,N_3205);
xnor U3488 (N_3488,N_3302,N_3298);
nor U3489 (N_3489,N_3271,N_3386);
or U3490 (N_3490,N_3249,N_3251);
and U3491 (N_3491,N_3226,N_3204);
nor U3492 (N_3492,N_3369,N_3273);
nor U3493 (N_3493,N_3274,N_3309);
xnor U3494 (N_3494,N_3260,N_3334);
nand U3495 (N_3495,N_3248,N_3348);
nor U3496 (N_3496,N_3343,N_3381);
nor U3497 (N_3497,N_3391,N_3238);
and U3498 (N_3498,N_3253,N_3349);
nor U3499 (N_3499,N_3287,N_3218);
nand U3500 (N_3500,N_3240,N_3365);
xor U3501 (N_3501,N_3354,N_3321);
xnor U3502 (N_3502,N_3318,N_3264);
nor U3503 (N_3503,N_3203,N_3306);
and U3504 (N_3504,N_3266,N_3351);
or U3505 (N_3505,N_3257,N_3318);
and U3506 (N_3506,N_3239,N_3348);
nor U3507 (N_3507,N_3339,N_3378);
and U3508 (N_3508,N_3314,N_3219);
nand U3509 (N_3509,N_3288,N_3205);
or U3510 (N_3510,N_3397,N_3355);
and U3511 (N_3511,N_3332,N_3225);
and U3512 (N_3512,N_3290,N_3384);
or U3513 (N_3513,N_3237,N_3381);
nand U3514 (N_3514,N_3357,N_3277);
nand U3515 (N_3515,N_3282,N_3248);
nor U3516 (N_3516,N_3241,N_3314);
or U3517 (N_3517,N_3246,N_3327);
or U3518 (N_3518,N_3270,N_3217);
and U3519 (N_3519,N_3364,N_3386);
and U3520 (N_3520,N_3207,N_3395);
and U3521 (N_3521,N_3316,N_3222);
or U3522 (N_3522,N_3205,N_3270);
and U3523 (N_3523,N_3284,N_3339);
nor U3524 (N_3524,N_3340,N_3295);
nor U3525 (N_3525,N_3331,N_3368);
nor U3526 (N_3526,N_3211,N_3268);
nand U3527 (N_3527,N_3300,N_3248);
or U3528 (N_3528,N_3241,N_3341);
nor U3529 (N_3529,N_3278,N_3238);
nor U3530 (N_3530,N_3277,N_3387);
nor U3531 (N_3531,N_3219,N_3278);
and U3532 (N_3532,N_3286,N_3214);
nand U3533 (N_3533,N_3312,N_3354);
nor U3534 (N_3534,N_3255,N_3257);
nand U3535 (N_3535,N_3283,N_3267);
nor U3536 (N_3536,N_3240,N_3377);
or U3537 (N_3537,N_3201,N_3389);
nor U3538 (N_3538,N_3221,N_3373);
nand U3539 (N_3539,N_3287,N_3289);
xor U3540 (N_3540,N_3385,N_3363);
nor U3541 (N_3541,N_3294,N_3355);
nor U3542 (N_3542,N_3360,N_3392);
and U3543 (N_3543,N_3367,N_3350);
and U3544 (N_3544,N_3210,N_3337);
nand U3545 (N_3545,N_3287,N_3274);
or U3546 (N_3546,N_3277,N_3280);
xor U3547 (N_3547,N_3278,N_3251);
and U3548 (N_3548,N_3320,N_3341);
and U3549 (N_3549,N_3279,N_3278);
nand U3550 (N_3550,N_3298,N_3388);
nand U3551 (N_3551,N_3263,N_3386);
nor U3552 (N_3552,N_3381,N_3233);
or U3553 (N_3553,N_3366,N_3312);
nand U3554 (N_3554,N_3388,N_3252);
nand U3555 (N_3555,N_3308,N_3381);
nand U3556 (N_3556,N_3285,N_3234);
and U3557 (N_3557,N_3271,N_3323);
nand U3558 (N_3558,N_3380,N_3242);
and U3559 (N_3559,N_3239,N_3250);
and U3560 (N_3560,N_3320,N_3304);
and U3561 (N_3561,N_3347,N_3238);
nor U3562 (N_3562,N_3386,N_3276);
xnor U3563 (N_3563,N_3265,N_3220);
nor U3564 (N_3564,N_3344,N_3239);
nand U3565 (N_3565,N_3211,N_3274);
nand U3566 (N_3566,N_3265,N_3239);
nor U3567 (N_3567,N_3363,N_3398);
or U3568 (N_3568,N_3341,N_3229);
and U3569 (N_3569,N_3263,N_3341);
nand U3570 (N_3570,N_3323,N_3212);
or U3571 (N_3571,N_3237,N_3299);
and U3572 (N_3572,N_3281,N_3394);
nor U3573 (N_3573,N_3231,N_3220);
or U3574 (N_3574,N_3346,N_3322);
and U3575 (N_3575,N_3235,N_3333);
nor U3576 (N_3576,N_3301,N_3237);
xor U3577 (N_3577,N_3292,N_3287);
and U3578 (N_3578,N_3261,N_3378);
nor U3579 (N_3579,N_3293,N_3244);
or U3580 (N_3580,N_3285,N_3202);
or U3581 (N_3581,N_3364,N_3203);
nand U3582 (N_3582,N_3348,N_3338);
or U3583 (N_3583,N_3335,N_3323);
or U3584 (N_3584,N_3315,N_3237);
or U3585 (N_3585,N_3275,N_3313);
nor U3586 (N_3586,N_3321,N_3337);
nand U3587 (N_3587,N_3345,N_3394);
xnor U3588 (N_3588,N_3249,N_3397);
or U3589 (N_3589,N_3308,N_3301);
or U3590 (N_3590,N_3386,N_3223);
and U3591 (N_3591,N_3322,N_3215);
nor U3592 (N_3592,N_3274,N_3310);
nand U3593 (N_3593,N_3263,N_3360);
nand U3594 (N_3594,N_3365,N_3339);
nor U3595 (N_3595,N_3253,N_3233);
xor U3596 (N_3596,N_3234,N_3360);
and U3597 (N_3597,N_3323,N_3325);
xor U3598 (N_3598,N_3290,N_3311);
xnor U3599 (N_3599,N_3282,N_3363);
nor U3600 (N_3600,N_3462,N_3580);
nand U3601 (N_3601,N_3433,N_3441);
and U3602 (N_3602,N_3592,N_3477);
and U3603 (N_3603,N_3567,N_3550);
xor U3604 (N_3604,N_3436,N_3468);
nor U3605 (N_3605,N_3405,N_3479);
xnor U3606 (N_3606,N_3529,N_3475);
and U3607 (N_3607,N_3534,N_3419);
nor U3608 (N_3608,N_3552,N_3450);
and U3609 (N_3609,N_3571,N_3528);
nor U3610 (N_3610,N_3507,N_3482);
or U3611 (N_3611,N_3535,N_3515);
nor U3612 (N_3612,N_3533,N_3585);
and U3613 (N_3613,N_3538,N_3536);
nor U3614 (N_3614,N_3532,N_3467);
and U3615 (N_3615,N_3430,N_3444);
xor U3616 (N_3616,N_3478,N_3516);
or U3617 (N_3617,N_3502,N_3497);
xor U3618 (N_3618,N_3511,N_3434);
and U3619 (N_3619,N_3403,N_3593);
nor U3620 (N_3620,N_3411,N_3429);
nor U3621 (N_3621,N_3527,N_3442);
xnor U3622 (N_3622,N_3590,N_3579);
nor U3623 (N_3623,N_3447,N_3598);
nand U3624 (N_3624,N_3588,N_3481);
nand U3625 (N_3625,N_3406,N_3470);
and U3626 (N_3626,N_3489,N_3460);
nand U3627 (N_3627,N_3524,N_3424);
nand U3628 (N_3628,N_3546,N_3574);
nor U3629 (N_3629,N_3488,N_3586);
or U3630 (N_3630,N_3496,N_3408);
xor U3631 (N_3631,N_3576,N_3548);
xor U3632 (N_3632,N_3509,N_3565);
and U3633 (N_3633,N_3453,N_3578);
nor U3634 (N_3634,N_3404,N_3537);
and U3635 (N_3635,N_3540,N_3422);
or U3636 (N_3636,N_3438,N_3577);
or U3637 (N_3637,N_3506,N_3448);
and U3638 (N_3638,N_3541,N_3547);
nor U3639 (N_3639,N_3581,N_3484);
nor U3640 (N_3640,N_3530,N_3432);
nor U3641 (N_3641,N_3518,N_3415);
nand U3642 (N_3642,N_3495,N_3457);
nand U3643 (N_3643,N_3575,N_3491);
nand U3644 (N_3644,N_3525,N_3499);
and U3645 (N_3645,N_3560,N_3439);
or U3646 (N_3646,N_3522,N_3417);
nor U3647 (N_3647,N_3437,N_3519);
nor U3648 (N_3648,N_3517,N_3410);
nand U3649 (N_3649,N_3555,N_3568);
xnor U3650 (N_3650,N_3451,N_3458);
nand U3651 (N_3651,N_3539,N_3523);
and U3652 (N_3652,N_3583,N_3445);
nor U3653 (N_3653,N_3589,N_3493);
and U3654 (N_3654,N_3483,N_3423);
xnor U3655 (N_3655,N_3465,N_3513);
nor U3656 (N_3656,N_3510,N_3400);
nand U3657 (N_3657,N_3456,N_3485);
nand U3658 (N_3658,N_3553,N_3473);
nor U3659 (N_3659,N_3584,N_3492);
nor U3660 (N_3660,N_3596,N_3463);
nor U3661 (N_3661,N_3490,N_3431);
or U3662 (N_3662,N_3564,N_3542);
and U3663 (N_3663,N_3494,N_3500);
or U3664 (N_3664,N_3435,N_3472);
nand U3665 (N_3665,N_3428,N_3420);
nor U3666 (N_3666,N_3461,N_3591);
or U3667 (N_3667,N_3466,N_3498);
or U3668 (N_3668,N_3526,N_3427);
or U3669 (N_3669,N_3440,N_3508);
nand U3670 (N_3670,N_3401,N_3446);
nand U3671 (N_3671,N_3409,N_3595);
or U3672 (N_3672,N_3452,N_3426);
or U3673 (N_3673,N_3469,N_3531);
or U3674 (N_3674,N_3421,N_3474);
nor U3675 (N_3675,N_3521,N_3573);
nand U3676 (N_3676,N_3597,N_3558);
or U3677 (N_3677,N_3599,N_3569);
nor U3678 (N_3678,N_3505,N_3554);
and U3679 (N_3679,N_3594,N_3449);
nor U3680 (N_3680,N_3504,N_3563);
and U3681 (N_3681,N_3561,N_3459);
nor U3682 (N_3682,N_3545,N_3503);
or U3683 (N_3683,N_3486,N_3425);
or U3684 (N_3684,N_3556,N_3520);
nand U3685 (N_3685,N_3416,N_3471);
nand U3686 (N_3686,N_3476,N_3455);
or U3687 (N_3687,N_3566,N_3413);
or U3688 (N_3688,N_3549,N_3443);
or U3689 (N_3689,N_3582,N_3414);
nand U3690 (N_3690,N_3570,N_3544);
nor U3691 (N_3691,N_3514,N_3412);
nor U3692 (N_3692,N_3407,N_3418);
and U3693 (N_3693,N_3562,N_3464);
nor U3694 (N_3694,N_3543,N_3587);
and U3695 (N_3695,N_3402,N_3551);
and U3696 (N_3696,N_3487,N_3557);
and U3697 (N_3697,N_3501,N_3512);
nor U3698 (N_3698,N_3454,N_3480);
or U3699 (N_3699,N_3572,N_3559);
or U3700 (N_3700,N_3537,N_3423);
nor U3701 (N_3701,N_3515,N_3488);
and U3702 (N_3702,N_3515,N_3557);
or U3703 (N_3703,N_3594,N_3411);
nor U3704 (N_3704,N_3588,N_3519);
nor U3705 (N_3705,N_3491,N_3580);
and U3706 (N_3706,N_3569,N_3510);
and U3707 (N_3707,N_3455,N_3575);
and U3708 (N_3708,N_3407,N_3510);
and U3709 (N_3709,N_3490,N_3585);
nor U3710 (N_3710,N_3475,N_3471);
or U3711 (N_3711,N_3576,N_3413);
or U3712 (N_3712,N_3584,N_3528);
or U3713 (N_3713,N_3492,N_3400);
nand U3714 (N_3714,N_3490,N_3598);
nand U3715 (N_3715,N_3479,N_3477);
and U3716 (N_3716,N_3419,N_3413);
or U3717 (N_3717,N_3445,N_3571);
nand U3718 (N_3718,N_3532,N_3473);
and U3719 (N_3719,N_3554,N_3580);
and U3720 (N_3720,N_3598,N_3470);
nor U3721 (N_3721,N_3410,N_3596);
and U3722 (N_3722,N_3525,N_3502);
nand U3723 (N_3723,N_3580,N_3599);
nand U3724 (N_3724,N_3549,N_3405);
and U3725 (N_3725,N_3481,N_3411);
and U3726 (N_3726,N_3413,N_3556);
nand U3727 (N_3727,N_3564,N_3465);
xor U3728 (N_3728,N_3567,N_3523);
nand U3729 (N_3729,N_3435,N_3498);
xor U3730 (N_3730,N_3409,N_3590);
nor U3731 (N_3731,N_3526,N_3562);
nor U3732 (N_3732,N_3474,N_3540);
nand U3733 (N_3733,N_3536,N_3540);
and U3734 (N_3734,N_3429,N_3511);
nor U3735 (N_3735,N_3511,N_3574);
and U3736 (N_3736,N_3493,N_3598);
nor U3737 (N_3737,N_3430,N_3418);
xor U3738 (N_3738,N_3421,N_3551);
nor U3739 (N_3739,N_3532,N_3531);
xor U3740 (N_3740,N_3568,N_3411);
or U3741 (N_3741,N_3410,N_3491);
nand U3742 (N_3742,N_3594,N_3404);
nor U3743 (N_3743,N_3493,N_3532);
or U3744 (N_3744,N_3431,N_3416);
nand U3745 (N_3745,N_3501,N_3571);
nand U3746 (N_3746,N_3408,N_3526);
nor U3747 (N_3747,N_3467,N_3403);
nor U3748 (N_3748,N_3447,N_3584);
or U3749 (N_3749,N_3425,N_3428);
xnor U3750 (N_3750,N_3578,N_3586);
nor U3751 (N_3751,N_3542,N_3536);
nor U3752 (N_3752,N_3523,N_3482);
or U3753 (N_3753,N_3401,N_3591);
nor U3754 (N_3754,N_3476,N_3459);
and U3755 (N_3755,N_3481,N_3479);
nand U3756 (N_3756,N_3448,N_3531);
and U3757 (N_3757,N_3440,N_3519);
and U3758 (N_3758,N_3466,N_3562);
and U3759 (N_3759,N_3444,N_3461);
and U3760 (N_3760,N_3590,N_3403);
nor U3761 (N_3761,N_3549,N_3483);
nor U3762 (N_3762,N_3434,N_3420);
and U3763 (N_3763,N_3458,N_3548);
nand U3764 (N_3764,N_3541,N_3486);
or U3765 (N_3765,N_3492,N_3475);
nor U3766 (N_3766,N_3589,N_3509);
or U3767 (N_3767,N_3598,N_3565);
and U3768 (N_3768,N_3444,N_3522);
nand U3769 (N_3769,N_3524,N_3401);
nand U3770 (N_3770,N_3405,N_3592);
nor U3771 (N_3771,N_3492,N_3503);
nand U3772 (N_3772,N_3540,N_3599);
or U3773 (N_3773,N_3524,N_3483);
or U3774 (N_3774,N_3577,N_3423);
nand U3775 (N_3775,N_3594,N_3460);
and U3776 (N_3776,N_3562,N_3534);
and U3777 (N_3777,N_3408,N_3420);
nor U3778 (N_3778,N_3440,N_3545);
or U3779 (N_3779,N_3440,N_3567);
nor U3780 (N_3780,N_3420,N_3522);
nand U3781 (N_3781,N_3580,N_3432);
and U3782 (N_3782,N_3574,N_3471);
nand U3783 (N_3783,N_3412,N_3484);
nand U3784 (N_3784,N_3499,N_3553);
xor U3785 (N_3785,N_3418,N_3488);
xor U3786 (N_3786,N_3540,N_3504);
and U3787 (N_3787,N_3594,N_3415);
nand U3788 (N_3788,N_3415,N_3536);
nor U3789 (N_3789,N_3586,N_3553);
nand U3790 (N_3790,N_3554,N_3436);
or U3791 (N_3791,N_3427,N_3405);
nand U3792 (N_3792,N_3580,N_3412);
nand U3793 (N_3793,N_3536,N_3484);
nor U3794 (N_3794,N_3490,N_3519);
nand U3795 (N_3795,N_3439,N_3483);
nor U3796 (N_3796,N_3523,N_3424);
nand U3797 (N_3797,N_3406,N_3590);
nand U3798 (N_3798,N_3513,N_3595);
nand U3799 (N_3799,N_3415,N_3564);
and U3800 (N_3800,N_3672,N_3625);
or U3801 (N_3801,N_3737,N_3742);
or U3802 (N_3802,N_3622,N_3739);
nor U3803 (N_3803,N_3615,N_3600);
nand U3804 (N_3804,N_3634,N_3710);
nor U3805 (N_3805,N_3741,N_3692);
and U3806 (N_3806,N_3708,N_3635);
nand U3807 (N_3807,N_3650,N_3761);
or U3808 (N_3808,N_3711,N_3719);
and U3809 (N_3809,N_3674,N_3798);
nand U3810 (N_3810,N_3767,N_3725);
and U3811 (N_3811,N_3653,N_3628);
and U3812 (N_3812,N_3655,N_3639);
and U3813 (N_3813,N_3790,N_3651);
and U3814 (N_3814,N_3694,N_3661);
nor U3815 (N_3815,N_3733,N_3760);
nand U3816 (N_3816,N_3702,N_3676);
nand U3817 (N_3817,N_3657,N_3620);
and U3818 (N_3818,N_3648,N_3637);
or U3819 (N_3819,N_3675,N_3682);
xor U3820 (N_3820,N_3613,N_3605);
nand U3821 (N_3821,N_3736,N_3746);
nand U3822 (N_3822,N_3783,N_3602);
or U3823 (N_3823,N_3716,N_3751);
and U3824 (N_3824,N_3713,N_3645);
nand U3825 (N_3825,N_3734,N_3730);
nand U3826 (N_3826,N_3705,N_3792);
or U3827 (N_3827,N_3677,N_3723);
nor U3828 (N_3828,N_3771,N_3683);
nor U3829 (N_3829,N_3631,N_3784);
and U3830 (N_3830,N_3652,N_3757);
nand U3831 (N_3831,N_3765,N_3715);
and U3832 (N_3832,N_3781,N_3778);
or U3833 (N_3833,N_3772,N_3775);
xnor U3834 (N_3834,N_3685,N_3782);
nand U3835 (N_3835,N_3623,N_3680);
nand U3836 (N_3836,N_3799,N_3610);
nor U3837 (N_3837,N_3749,N_3614);
nand U3838 (N_3838,N_3754,N_3774);
nand U3839 (N_3839,N_3776,N_3649);
or U3840 (N_3840,N_3756,N_3670);
or U3841 (N_3841,N_3704,N_3750);
nand U3842 (N_3842,N_3681,N_3640);
nand U3843 (N_3843,N_3611,N_3633);
or U3844 (N_3844,N_3712,N_3687);
nand U3845 (N_3845,N_3696,N_3743);
nor U3846 (N_3846,N_3787,N_3709);
nand U3847 (N_3847,N_3607,N_3647);
nand U3848 (N_3848,N_3618,N_3797);
or U3849 (N_3849,N_3759,N_3728);
nand U3850 (N_3850,N_3752,N_3636);
and U3851 (N_3851,N_3724,N_3748);
nand U3852 (N_3852,N_3608,N_3662);
or U3853 (N_3853,N_3638,N_3766);
xnor U3854 (N_3854,N_3668,N_3617);
nand U3855 (N_3855,N_3789,N_3658);
and U3856 (N_3856,N_3673,N_3606);
nand U3857 (N_3857,N_3786,N_3745);
and U3858 (N_3858,N_3763,N_3769);
and U3859 (N_3859,N_3758,N_3735);
nand U3860 (N_3860,N_3768,N_3701);
xnor U3861 (N_3861,N_3744,N_3740);
nand U3862 (N_3862,N_3604,N_3779);
or U3863 (N_3863,N_3686,N_3732);
nand U3864 (N_3864,N_3679,N_3659);
and U3865 (N_3865,N_3664,N_3717);
or U3866 (N_3866,N_3678,N_3747);
or U3867 (N_3867,N_3770,N_3699);
and U3868 (N_3868,N_3643,N_3632);
nand U3869 (N_3869,N_3788,N_3738);
nand U3870 (N_3870,N_3684,N_3707);
and U3871 (N_3871,N_3718,N_3693);
nand U3872 (N_3872,N_3700,N_3698);
or U3873 (N_3873,N_3726,N_3729);
nor U3874 (N_3874,N_3644,N_3795);
and U3875 (N_3875,N_3642,N_3706);
nand U3876 (N_3876,N_3755,N_3663);
nand U3877 (N_3877,N_3601,N_3616);
and U3878 (N_3878,N_3689,N_3697);
nor U3879 (N_3879,N_3665,N_3609);
and U3880 (N_3880,N_3671,N_3654);
xor U3881 (N_3881,N_3780,N_3619);
nor U3882 (N_3882,N_3630,N_3731);
and U3883 (N_3883,N_3764,N_3753);
nand U3884 (N_3884,N_3688,N_3656);
xnor U3885 (N_3885,N_3669,N_3641);
and U3886 (N_3886,N_3785,N_3794);
or U3887 (N_3887,N_3612,N_3762);
nor U3888 (N_3888,N_3621,N_3690);
nor U3889 (N_3889,N_3626,N_3773);
or U3890 (N_3890,N_3720,N_3796);
or U3891 (N_3891,N_3646,N_3691);
nor U3892 (N_3892,N_3777,N_3791);
and U3893 (N_3893,N_3721,N_3627);
xor U3894 (N_3894,N_3667,N_3727);
or U3895 (N_3895,N_3722,N_3714);
and U3896 (N_3896,N_3660,N_3703);
or U3897 (N_3897,N_3629,N_3666);
or U3898 (N_3898,N_3695,N_3624);
nor U3899 (N_3899,N_3793,N_3603);
xor U3900 (N_3900,N_3609,N_3649);
nor U3901 (N_3901,N_3725,N_3713);
nand U3902 (N_3902,N_3745,N_3601);
nor U3903 (N_3903,N_3783,N_3740);
or U3904 (N_3904,N_3616,N_3642);
and U3905 (N_3905,N_3794,N_3749);
nor U3906 (N_3906,N_3712,N_3731);
nor U3907 (N_3907,N_3720,N_3664);
nor U3908 (N_3908,N_3685,N_3748);
xnor U3909 (N_3909,N_3748,N_3792);
xnor U3910 (N_3910,N_3747,N_3710);
nand U3911 (N_3911,N_3703,N_3700);
or U3912 (N_3912,N_3695,N_3750);
or U3913 (N_3913,N_3704,N_3743);
or U3914 (N_3914,N_3773,N_3653);
nor U3915 (N_3915,N_3748,N_3692);
and U3916 (N_3916,N_3621,N_3739);
nand U3917 (N_3917,N_3718,N_3628);
or U3918 (N_3918,N_3794,N_3780);
nand U3919 (N_3919,N_3732,N_3620);
nor U3920 (N_3920,N_3797,N_3633);
nand U3921 (N_3921,N_3638,N_3621);
and U3922 (N_3922,N_3621,N_3694);
nand U3923 (N_3923,N_3763,N_3781);
and U3924 (N_3924,N_3708,N_3780);
xor U3925 (N_3925,N_3641,N_3643);
or U3926 (N_3926,N_3756,N_3749);
or U3927 (N_3927,N_3602,N_3639);
xnor U3928 (N_3928,N_3729,N_3735);
and U3929 (N_3929,N_3771,N_3712);
nor U3930 (N_3930,N_3618,N_3770);
and U3931 (N_3931,N_3600,N_3670);
or U3932 (N_3932,N_3759,N_3633);
nor U3933 (N_3933,N_3713,N_3631);
nor U3934 (N_3934,N_3674,N_3669);
or U3935 (N_3935,N_3667,N_3654);
or U3936 (N_3936,N_3641,N_3640);
nand U3937 (N_3937,N_3727,N_3671);
and U3938 (N_3938,N_3694,N_3630);
nor U3939 (N_3939,N_3734,N_3714);
xnor U3940 (N_3940,N_3714,N_3660);
or U3941 (N_3941,N_3712,N_3726);
nand U3942 (N_3942,N_3674,N_3682);
and U3943 (N_3943,N_3656,N_3764);
or U3944 (N_3944,N_3741,N_3695);
xor U3945 (N_3945,N_3743,N_3707);
nand U3946 (N_3946,N_3709,N_3749);
or U3947 (N_3947,N_3639,N_3694);
or U3948 (N_3948,N_3691,N_3702);
or U3949 (N_3949,N_3639,N_3686);
nor U3950 (N_3950,N_3765,N_3680);
nor U3951 (N_3951,N_3641,N_3652);
nor U3952 (N_3952,N_3731,N_3667);
or U3953 (N_3953,N_3624,N_3629);
xor U3954 (N_3954,N_3696,N_3769);
or U3955 (N_3955,N_3768,N_3722);
and U3956 (N_3956,N_3616,N_3798);
and U3957 (N_3957,N_3624,N_3765);
nor U3958 (N_3958,N_3760,N_3691);
and U3959 (N_3959,N_3773,N_3795);
or U3960 (N_3960,N_3720,N_3644);
or U3961 (N_3961,N_3620,N_3729);
nand U3962 (N_3962,N_3644,N_3620);
nand U3963 (N_3963,N_3686,N_3695);
nor U3964 (N_3964,N_3656,N_3617);
nand U3965 (N_3965,N_3682,N_3742);
nand U3966 (N_3966,N_3698,N_3648);
nand U3967 (N_3967,N_3673,N_3687);
nand U3968 (N_3968,N_3654,N_3732);
nand U3969 (N_3969,N_3636,N_3788);
nor U3970 (N_3970,N_3626,N_3750);
or U3971 (N_3971,N_3723,N_3733);
and U3972 (N_3972,N_3753,N_3675);
nor U3973 (N_3973,N_3708,N_3718);
nand U3974 (N_3974,N_3645,N_3769);
or U3975 (N_3975,N_3618,N_3784);
nor U3976 (N_3976,N_3653,N_3703);
and U3977 (N_3977,N_3754,N_3786);
or U3978 (N_3978,N_3773,N_3657);
nor U3979 (N_3979,N_3671,N_3796);
xor U3980 (N_3980,N_3645,N_3784);
xnor U3981 (N_3981,N_3633,N_3645);
and U3982 (N_3982,N_3734,N_3727);
or U3983 (N_3983,N_3756,N_3730);
xor U3984 (N_3984,N_3680,N_3747);
or U3985 (N_3985,N_3772,N_3789);
nor U3986 (N_3986,N_3756,N_3701);
nor U3987 (N_3987,N_3782,N_3726);
and U3988 (N_3988,N_3645,N_3686);
nor U3989 (N_3989,N_3625,N_3660);
nor U3990 (N_3990,N_3604,N_3685);
xnor U3991 (N_3991,N_3778,N_3695);
and U3992 (N_3992,N_3600,N_3742);
and U3993 (N_3993,N_3706,N_3795);
and U3994 (N_3994,N_3776,N_3610);
or U3995 (N_3995,N_3653,N_3766);
or U3996 (N_3996,N_3664,N_3757);
nand U3997 (N_3997,N_3613,N_3620);
nand U3998 (N_3998,N_3732,N_3786);
nand U3999 (N_3999,N_3721,N_3693);
nand U4000 (N_4000,N_3925,N_3971);
nand U4001 (N_4001,N_3814,N_3897);
nor U4002 (N_4002,N_3819,N_3886);
or U4003 (N_4003,N_3860,N_3878);
or U4004 (N_4004,N_3845,N_3888);
nand U4005 (N_4005,N_3895,N_3879);
nand U4006 (N_4006,N_3913,N_3958);
and U4007 (N_4007,N_3944,N_3810);
xnor U4008 (N_4008,N_3893,N_3969);
nor U4009 (N_4009,N_3873,N_3880);
or U4010 (N_4010,N_3833,N_3919);
or U4011 (N_4011,N_3938,N_3986);
or U4012 (N_4012,N_3943,N_3800);
and U4013 (N_4013,N_3834,N_3826);
nor U4014 (N_4014,N_3941,N_3965);
xor U4015 (N_4015,N_3973,N_3920);
or U4016 (N_4016,N_3823,N_3989);
and U4017 (N_4017,N_3949,N_3927);
nand U4018 (N_4018,N_3948,N_3859);
and U4019 (N_4019,N_3945,N_3837);
or U4020 (N_4020,N_3858,N_3866);
or U4021 (N_4021,N_3975,N_3831);
or U4022 (N_4022,N_3882,N_3961);
nand U4023 (N_4023,N_3933,N_3898);
or U4024 (N_4024,N_3972,N_3850);
and U4025 (N_4025,N_3844,N_3853);
xnor U4026 (N_4026,N_3929,N_3952);
nand U4027 (N_4027,N_3906,N_3911);
xnor U4028 (N_4028,N_3870,N_3977);
or U4029 (N_4029,N_3835,N_3808);
or U4030 (N_4030,N_3852,N_3816);
nand U4031 (N_4031,N_3851,N_3841);
and U4032 (N_4032,N_3817,N_3926);
or U4033 (N_4033,N_3830,N_3918);
xnor U4034 (N_4034,N_3954,N_3802);
nand U4035 (N_4035,N_3909,N_3912);
and U4036 (N_4036,N_3946,N_3967);
nand U4037 (N_4037,N_3900,N_3891);
or U4038 (N_4038,N_3990,N_3923);
nor U4039 (N_4039,N_3963,N_3979);
nor U4040 (N_4040,N_3884,N_3983);
xnor U4041 (N_4041,N_3905,N_3924);
nand U4042 (N_4042,N_3892,N_3854);
or U4043 (N_4043,N_3931,N_3887);
nand U4044 (N_4044,N_3825,N_3863);
or U4045 (N_4045,N_3836,N_3857);
or U4046 (N_4046,N_3978,N_3970);
nand U4047 (N_4047,N_3827,N_3940);
nand U4048 (N_4048,N_3981,N_3984);
or U4049 (N_4049,N_3813,N_3822);
nor U4050 (N_4050,N_3801,N_3875);
or U4051 (N_4051,N_3997,N_3820);
nor U4052 (N_4052,N_3921,N_3957);
nor U4053 (N_4053,N_3914,N_3915);
or U4054 (N_4054,N_3907,N_3966);
nor U4055 (N_4055,N_3818,N_3987);
nand U4056 (N_4056,N_3992,N_3899);
or U4057 (N_4057,N_3876,N_3842);
or U4058 (N_4058,N_3885,N_3883);
and U4059 (N_4059,N_3824,N_3991);
and U4060 (N_4060,N_3934,N_3838);
or U4061 (N_4061,N_3947,N_3815);
nand U4062 (N_4062,N_3902,N_3894);
nor U4063 (N_4063,N_3917,N_3960);
nor U4064 (N_4064,N_3928,N_3910);
xor U4065 (N_4065,N_3829,N_3951);
and U4066 (N_4066,N_3889,N_3982);
and U4067 (N_4067,N_3994,N_3996);
or U4068 (N_4068,N_3806,N_3932);
xor U4069 (N_4069,N_3872,N_3890);
nor U4070 (N_4070,N_3867,N_3862);
nor U4071 (N_4071,N_3877,N_3896);
xnor U4072 (N_4072,N_3955,N_3936);
nand U4073 (N_4073,N_3803,N_3942);
and U4074 (N_4074,N_3956,N_3922);
or U4075 (N_4075,N_3950,N_3809);
xor U4076 (N_4076,N_3843,N_3935);
and U4077 (N_4077,N_3861,N_3839);
nor U4078 (N_4078,N_3937,N_3976);
nand U4079 (N_4079,N_3939,N_3856);
nor U4080 (N_4080,N_3901,N_3807);
nand U4081 (N_4081,N_3828,N_3821);
and U4082 (N_4082,N_3974,N_3964);
nor U4083 (N_4083,N_3832,N_3812);
nor U4084 (N_4084,N_3811,N_3999);
and U4085 (N_4085,N_3874,N_3988);
nor U4086 (N_4086,N_3908,N_3869);
or U4087 (N_4087,N_3930,N_3848);
nor U4088 (N_4088,N_3980,N_3953);
nand U4089 (N_4089,N_3849,N_3985);
nand U4090 (N_4090,N_3847,N_3962);
xor U4091 (N_4091,N_3855,N_3998);
nor U4092 (N_4092,N_3805,N_3868);
or U4093 (N_4093,N_3871,N_3993);
or U4094 (N_4094,N_3904,N_3968);
and U4095 (N_4095,N_3903,N_3881);
nor U4096 (N_4096,N_3916,N_3865);
or U4097 (N_4097,N_3804,N_3864);
or U4098 (N_4098,N_3995,N_3959);
and U4099 (N_4099,N_3840,N_3846);
nor U4100 (N_4100,N_3911,N_3878);
nand U4101 (N_4101,N_3888,N_3992);
nor U4102 (N_4102,N_3985,N_3919);
or U4103 (N_4103,N_3849,N_3923);
or U4104 (N_4104,N_3843,N_3802);
nand U4105 (N_4105,N_3840,N_3865);
nor U4106 (N_4106,N_3975,N_3921);
or U4107 (N_4107,N_3890,N_3899);
or U4108 (N_4108,N_3883,N_3908);
or U4109 (N_4109,N_3882,N_3938);
or U4110 (N_4110,N_3846,N_3891);
and U4111 (N_4111,N_3843,N_3815);
nor U4112 (N_4112,N_3895,N_3968);
or U4113 (N_4113,N_3961,N_3948);
or U4114 (N_4114,N_3922,N_3986);
xnor U4115 (N_4115,N_3876,N_3970);
or U4116 (N_4116,N_3845,N_3817);
nand U4117 (N_4117,N_3962,N_3837);
or U4118 (N_4118,N_3918,N_3898);
nand U4119 (N_4119,N_3885,N_3806);
and U4120 (N_4120,N_3820,N_3964);
or U4121 (N_4121,N_3824,N_3885);
nor U4122 (N_4122,N_3986,N_3873);
and U4123 (N_4123,N_3803,N_3921);
or U4124 (N_4124,N_3952,N_3867);
and U4125 (N_4125,N_3893,N_3868);
and U4126 (N_4126,N_3871,N_3865);
or U4127 (N_4127,N_3941,N_3966);
nand U4128 (N_4128,N_3908,N_3847);
nand U4129 (N_4129,N_3905,N_3982);
or U4130 (N_4130,N_3835,N_3978);
and U4131 (N_4131,N_3871,N_3955);
or U4132 (N_4132,N_3815,N_3966);
nand U4133 (N_4133,N_3992,N_3988);
and U4134 (N_4134,N_3978,N_3988);
and U4135 (N_4135,N_3802,N_3920);
xor U4136 (N_4136,N_3932,N_3886);
and U4137 (N_4137,N_3851,N_3800);
nor U4138 (N_4138,N_3877,N_3897);
nor U4139 (N_4139,N_3988,N_3964);
nor U4140 (N_4140,N_3904,N_3948);
nand U4141 (N_4141,N_3946,N_3888);
xor U4142 (N_4142,N_3803,N_3818);
nor U4143 (N_4143,N_3991,N_3896);
or U4144 (N_4144,N_3976,N_3842);
or U4145 (N_4145,N_3920,N_3815);
or U4146 (N_4146,N_3927,N_3966);
and U4147 (N_4147,N_3937,N_3852);
or U4148 (N_4148,N_3870,N_3988);
nor U4149 (N_4149,N_3859,N_3949);
nand U4150 (N_4150,N_3947,N_3913);
nand U4151 (N_4151,N_3990,N_3886);
nand U4152 (N_4152,N_3982,N_3800);
or U4153 (N_4153,N_3921,N_3889);
xnor U4154 (N_4154,N_3908,N_3910);
or U4155 (N_4155,N_3967,N_3952);
nand U4156 (N_4156,N_3808,N_3908);
nand U4157 (N_4157,N_3849,N_3852);
and U4158 (N_4158,N_3954,N_3890);
nand U4159 (N_4159,N_3932,N_3973);
and U4160 (N_4160,N_3886,N_3907);
and U4161 (N_4161,N_3876,N_3953);
nor U4162 (N_4162,N_3889,N_3989);
nor U4163 (N_4163,N_3892,N_3825);
nand U4164 (N_4164,N_3931,N_3879);
nand U4165 (N_4165,N_3894,N_3831);
and U4166 (N_4166,N_3852,N_3820);
or U4167 (N_4167,N_3958,N_3879);
xor U4168 (N_4168,N_3894,N_3806);
nor U4169 (N_4169,N_3994,N_3917);
or U4170 (N_4170,N_3998,N_3972);
and U4171 (N_4171,N_3994,N_3869);
and U4172 (N_4172,N_3931,N_3905);
nor U4173 (N_4173,N_3837,N_3801);
and U4174 (N_4174,N_3908,N_3981);
nor U4175 (N_4175,N_3813,N_3968);
nand U4176 (N_4176,N_3953,N_3912);
and U4177 (N_4177,N_3861,N_3811);
xor U4178 (N_4178,N_3893,N_3947);
nand U4179 (N_4179,N_3997,N_3933);
and U4180 (N_4180,N_3975,N_3966);
nand U4181 (N_4181,N_3987,N_3920);
and U4182 (N_4182,N_3860,N_3903);
nand U4183 (N_4183,N_3936,N_3938);
xnor U4184 (N_4184,N_3934,N_3844);
nand U4185 (N_4185,N_3905,N_3979);
and U4186 (N_4186,N_3810,N_3842);
nor U4187 (N_4187,N_3810,N_3920);
and U4188 (N_4188,N_3905,N_3970);
and U4189 (N_4189,N_3962,N_3823);
xor U4190 (N_4190,N_3953,N_3991);
or U4191 (N_4191,N_3876,N_3854);
nand U4192 (N_4192,N_3948,N_3929);
nand U4193 (N_4193,N_3885,N_3950);
nand U4194 (N_4194,N_3888,N_3909);
nand U4195 (N_4195,N_3957,N_3983);
or U4196 (N_4196,N_3904,N_3800);
nand U4197 (N_4197,N_3812,N_3827);
and U4198 (N_4198,N_3827,N_3892);
nor U4199 (N_4199,N_3930,N_3936);
and U4200 (N_4200,N_4154,N_4085);
or U4201 (N_4201,N_4128,N_4037);
or U4202 (N_4202,N_4108,N_4008);
nor U4203 (N_4203,N_4041,N_4179);
or U4204 (N_4204,N_4164,N_4029);
nor U4205 (N_4205,N_4073,N_4016);
or U4206 (N_4206,N_4076,N_4138);
and U4207 (N_4207,N_4094,N_4005);
or U4208 (N_4208,N_4100,N_4150);
nand U4209 (N_4209,N_4182,N_4056);
and U4210 (N_4210,N_4009,N_4066);
nand U4211 (N_4211,N_4007,N_4034);
and U4212 (N_4212,N_4134,N_4160);
or U4213 (N_4213,N_4099,N_4006);
or U4214 (N_4214,N_4199,N_4071);
and U4215 (N_4215,N_4000,N_4035);
nand U4216 (N_4216,N_4031,N_4090);
and U4217 (N_4217,N_4185,N_4119);
or U4218 (N_4218,N_4139,N_4170);
or U4219 (N_4219,N_4162,N_4125);
or U4220 (N_4220,N_4057,N_4093);
nor U4221 (N_4221,N_4190,N_4002);
nand U4222 (N_4222,N_4050,N_4054);
xor U4223 (N_4223,N_4178,N_4124);
or U4224 (N_4224,N_4149,N_4111);
and U4225 (N_4225,N_4055,N_4086);
and U4226 (N_4226,N_4053,N_4158);
nor U4227 (N_4227,N_4025,N_4147);
or U4228 (N_4228,N_4169,N_4188);
or U4229 (N_4229,N_4072,N_4001);
nand U4230 (N_4230,N_4081,N_4023);
or U4231 (N_4231,N_4064,N_4152);
nand U4232 (N_4232,N_4101,N_4137);
nand U4233 (N_4233,N_4194,N_4103);
xnor U4234 (N_4234,N_4112,N_4091);
and U4235 (N_4235,N_4187,N_4042);
and U4236 (N_4236,N_4095,N_4197);
or U4237 (N_4237,N_4051,N_4181);
and U4238 (N_4238,N_4084,N_4174);
nor U4239 (N_4239,N_4018,N_4166);
nand U4240 (N_4240,N_4087,N_4039);
or U4241 (N_4241,N_4156,N_4068);
or U4242 (N_4242,N_4048,N_4013);
nor U4243 (N_4243,N_4171,N_4104);
and U4244 (N_4244,N_4024,N_4049);
or U4245 (N_4245,N_4075,N_4184);
nor U4246 (N_4246,N_4074,N_4180);
or U4247 (N_4247,N_4019,N_4098);
xnor U4248 (N_4248,N_4129,N_4082);
nand U4249 (N_4249,N_4163,N_4140);
xnor U4250 (N_4250,N_4017,N_4172);
nor U4251 (N_4251,N_4153,N_4168);
xnor U4252 (N_4252,N_4047,N_4014);
xnor U4253 (N_4253,N_4126,N_4026);
nor U4254 (N_4254,N_4131,N_4012);
and U4255 (N_4255,N_4136,N_4141);
nand U4256 (N_4256,N_4117,N_4083);
nor U4257 (N_4257,N_4135,N_4148);
nand U4258 (N_4258,N_4105,N_4159);
xnor U4259 (N_4259,N_4130,N_4183);
and U4260 (N_4260,N_4033,N_4021);
and U4261 (N_4261,N_4122,N_4040);
nand U4262 (N_4262,N_4079,N_4062);
or U4263 (N_4263,N_4192,N_4109);
xor U4264 (N_4264,N_4102,N_4173);
xor U4265 (N_4265,N_4096,N_4186);
or U4266 (N_4266,N_4011,N_4092);
and U4267 (N_4267,N_4052,N_4046);
or U4268 (N_4268,N_4010,N_4132);
nor U4269 (N_4269,N_4088,N_4080);
xor U4270 (N_4270,N_4123,N_4195);
nand U4271 (N_4271,N_4198,N_4089);
and U4272 (N_4272,N_4045,N_4061);
and U4273 (N_4273,N_4155,N_4177);
and U4274 (N_4274,N_4028,N_4118);
nor U4275 (N_4275,N_4107,N_4044);
nor U4276 (N_4276,N_4110,N_4097);
and U4277 (N_4277,N_4176,N_4146);
nand U4278 (N_4278,N_4157,N_4127);
nand U4279 (N_4279,N_4106,N_4063);
nor U4280 (N_4280,N_4036,N_4116);
xnor U4281 (N_4281,N_4020,N_4003);
or U4282 (N_4282,N_4004,N_4043);
nand U4283 (N_4283,N_4142,N_4167);
xnor U4284 (N_4284,N_4058,N_4144);
nand U4285 (N_4285,N_4115,N_4196);
and U4286 (N_4286,N_4032,N_4191);
or U4287 (N_4287,N_4165,N_4151);
and U4288 (N_4288,N_4114,N_4065);
or U4289 (N_4289,N_4069,N_4161);
nor U4290 (N_4290,N_4067,N_4175);
or U4291 (N_4291,N_4121,N_4133);
xor U4292 (N_4292,N_4120,N_4145);
nor U4293 (N_4293,N_4078,N_4022);
or U4294 (N_4294,N_4070,N_4015);
xnor U4295 (N_4295,N_4027,N_4030);
xor U4296 (N_4296,N_4193,N_4059);
nor U4297 (N_4297,N_4189,N_4113);
and U4298 (N_4298,N_4143,N_4060);
nor U4299 (N_4299,N_4077,N_4038);
and U4300 (N_4300,N_4079,N_4156);
nor U4301 (N_4301,N_4018,N_4158);
nand U4302 (N_4302,N_4151,N_4083);
and U4303 (N_4303,N_4146,N_4068);
nor U4304 (N_4304,N_4143,N_4084);
nand U4305 (N_4305,N_4190,N_4092);
nor U4306 (N_4306,N_4170,N_4102);
xor U4307 (N_4307,N_4009,N_4173);
nor U4308 (N_4308,N_4102,N_4003);
nand U4309 (N_4309,N_4002,N_4005);
or U4310 (N_4310,N_4110,N_4076);
and U4311 (N_4311,N_4150,N_4037);
or U4312 (N_4312,N_4165,N_4169);
xor U4313 (N_4313,N_4007,N_4088);
nor U4314 (N_4314,N_4111,N_4076);
and U4315 (N_4315,N_4158,N_4020);
and U4316 (N_4316,N_4134,N_4161);
and U4317 (N_4317,N_4138,N_4038);
or U4318 (N_4318,N_4154,N_4062);
xnor U4319 (N_4319,N_4005,N_4179);
xor U4320 (N_4320,N_4194,N_4043);
or U4321 (N_4321,N_4162,N_4170);
or U4322 (N_4322,N_4059,N_4034);
xor U4323 (N_4323,N_4188,N_4141);
or U4324 (N_4324,N_4196,N_4068);
xnor U4325 (N_4325,N_4173,N_4134);
xnor U4326 (N_4326,N_4034,N_4046);
or U4327 (N_4327,N_4195,N_4027);
nand U4328 (N_4328,N_4141,N_4086);
nor U4329 (N_4329,N_4169,N_4177);
xor U4330 (N_4330,N_4013,N_4128);
nand U4331 (N_4331,N_4070,N_4026);
and U4332 (N_4332,N_4063,N_4104);
and U4333 (N_4333,N_4005,N_4024);
nor U4334 (N_4334,N_4128,N_4193);
nor U4335 (N_4335,N_4051,N_4132);
and U4336 (N_4336,N_4114,N_4005);
nor U4337 (N_4337,N_4129,N_4053);
and U4338 (N_4338,N_4159,N_4169);
or U4339 (N_4339,N_4169,N_4131);
or U4340 (N_4340,N_4179,N_4198);
nor U4341 (N_4341,N_4185,N_4037);
xor U4342 (N_4342,N_4053,N_4022);
nor U4343 (N_4343,N_4148,N_4184);
nor U4344 (N_4344,N_4129,N_4000);
or U4345 (N_4345,N_4047,N_4084);
nand U4346 (N_4346,N_4105,N_4029);
or U4347 (N_4347,N_4056,N_4144);
and U4348 (N_4348,N_4001,N_4116);
and U4349 (N_4349,N_4112,N_4140);
or U4350 (N_4350,N_4062,N_4150);
nand U4351 (N_4351,N_4188,N_4029);
nand U4352 (N_4352,N_4188,N_4032);
and U4353 (N_4353,N_4162,N_4133);
and U4354 (N_4354,N_4180,N_4085);
nand U4355 (N_4355,N_4059,N_4023);
nor U4356 (N_4356,N_4022,N_4051);
or U4357 (N_4357,N_4095,N_4104);
nand U4358 (N_4358,N_4109,N_4003);
or U4359 (N_4359,N_4041,N_4182);
or U4360 (N_4360,N_4120,N_4173);
nor U4361 (N_4361,N_4139,N_4012);
nand U4362 (N_4362,N_4039,N_4034);
nand U4363 (N_4363,N_4032,N_4041);
nor U4364 (N_4364,N_4100,N_4163);
or U4365 (N_4365,N_4186,N_4160);
nand U4366 (N_4366,N_4103,N_4135);
or U4367 (N_4367,N_4090,N_4116);
xnor U4368 (N_4368,N_4147,N_4051);
xnor U4369 (N_4369,N_4061,N_4043);
xor U4370 (N_4370,N_4155,N_4180);
nor U4371 (N_4371,N_4136,N_4183);
or U4372 (N_4372,N_4030,N_4052);
xor U4373 (N_4373,N_4106,N_4029);
nor U4374 (N_4374,N_4084,N_4094);
nor U4375 (N_4375,N_4175,N_4083);
nand U4376 (N_4376,N_4098,N_4191);
or U4377 (N_4377,N_4195,N_4048);
nor U4378 (N_4378,N_4133,N_4009);
nor U4379 (N_4379,N_4195,N_4119);
or U4380 (N_4380,N_4071,N_4188);
nor U4381 (N_4381,N_4059,N_4138);
or U4382 (N_4382,N_4159,N_4012);
or U4383 (N_4383,N_4064,N_4184);
nand U4384 (N_4384,N_4097,N_4072);
nand U4385 (N_4385,N_4130,N_4146);
or U4386 (N_4386,N_4057,N_4182);
and U4387 (N_4387,N_4009,N_4187);
nand U4388 (N_4388,N_4058,N_4094);
and U4389 (N_4389,N_4094,N_4109);
nor U4390 (N_4390,N_4096,N_4008);
nor U4391 (N_4391,N_4087,N_4086);
nor U4392 (N_4392,N_4115,N_4146);
nor U4393 (N_4393,N_4098,N_4065);
or U4394 (N_4394,N_4171,N_4071);
nand U4395 (N_4395,N_4046,N_4083);
or U4396 (N_4396,N_4081,N_4051);
nor U4397 (N_4397,N_4162,N_4031);
nor U4398 (N_4398,N_4058,N_4172);
nand U4399 (N_4399,N_4112,N_4169);
xnor U4400 (N_4400,N_4309,N_4396);
or U4401 (N_4401,N_4232,N_4277);
nand U4402 (N_4402,N_4275,N_4241);
nor U4403 (N_4403,N_4305,N_4391);
nor U4404 (N_4404,N_4372,N_4387);
nor U4405 (N_4405,N_4316,N_4299);
nand U4406 (N_4406,N_4226,N_4202);
or U4407 (N_4407,N_4326,N_4247);
or U4408 (N_4408,N_4356,N_4203);
or U4409 (N_4409,N_4369,N_4265);
nor U4410 (N_4410,N_4227,N_4392);
or U4411 (N_4411,N_4332,N_4243);
or U4412 (N_4412,N_4220,N_4231);
nand U4413 (N_4413,N_4298,N_4230);
nand U4414 (N_4414,N_4266,N_4293);
and U4415 (N_4415,N_4268,N_4279);
nand U4416 (N_4416,N_4329,N_4375);
or U4417 (N_4417,N_4288,N_4398);
nand U4418 (N_4418,N_4336,N_4290);
nor U4419 (N_4419,N_4322,N_4325);
nor U4420 (N_4420,N_4307,N_4393);
and U4421 (N_4421,N_4389,N_4378);
nand U4422 (N_4422,N_4364,N_4251);
nand U4423 (N_4423,N_4354,N_4271);
nor U4424 (N_4424,N_4286,N_4225);
and U4425 (N_4425,N_4291,N_4386);
xor U4426 (N_4426,N_4315,N_4201);
nor U4427 (N_4427,N_4260,N_4381);
nor U4428 (N_4428,N_4397,N_4211);
nand U4429 (N_4429,N_4330,N_4360);
nand U4430 (N_4430,N_4242,N_4347);
and U4431 (N_4431,N_4212,N_4344);
nand U4432 (N_4432,N_4294,N_4323);
or U4433 (N_4433,N_4320,N_4258);
and U4434 (N_4434,N_4333,N_4281);
or U4435 (N_4435,N_4215,N_4273);
nor U4436 (N_4436,N_4287,N_4246);
nand U4437 (N_4437,N_4341,N_4257);
nor U4438 (N_4438,N_4306,N_4269);
and U4439 (N_4439,N_4228,N_4334);
and U4440 (N_4440,N_4236,N_4350);
and U4441 (N_4441,N_4283,N_4224);
nand U4442 (N_4442,N_4346,N_4348);
nand U4443 (N_4443,N_4352,N_4342);
xor U4444 (N_4444,N_4249,N_4335);
and U4445 (N_4445,N_4217,N_4284);
or U4446 (N_4446,N_4376,N_4317);
nand U4447 (N_4447,N_4244,N_4245);
nand U4448 (N_4448,N_4355,N_4278);
nand U4449 (N_4449,N_4327,N_4351);
nor U4450 (N_4450,N_4235,N_4263);
nand U4451 (N_4451,N_4267,N_4382);
or U4452 (N_4452,N_4308,N_4264);
or U4453 (N_4453,N_4303,N_4373);
nand U4454 (N_4454,N_4312,N_4274);
nand U4455 (N_4455,N_4349,N_4248);
nand U4456 (N_4456,N_4216,N_4261);
nand U4457 (N_4457,N_4363,N_4318);
and U4458 (N_4458,N_4313,N_4328);
nand U4459 (N_4459,N_4256,N_4214);
and U4460 (N_4460,N_4365,N_4234);
nand U4461 (N_4461,N_4207,N_4395);
nand U4462 (N_4462,N_4210,N_4379);
nand U4463 (N_4463,N_4200,N_4361);
or U4464 (N_4464,N_4295,N_4221);
xnor U4465 (N_4465,N_4310,N_4345);
nand U4466 (N_4466,N_4304,N_4383);
nor U4467 (N_4467,N_4219,N_4205);
and U4468 (N_4468,N_4302,N_4292);
or U4469 (N_4469,N_4324,N_4358);
and U4470 (N_4470,N_4340,N_4223);
nor U4471 (N_4471,N_4370,N_4296);
nor U4472 (N_4472,N_4311,N_4321);
or U4473 (N_4473,N_4240,N_4255);
nor U4474 (N_4474,N_4394,N_4388);
or U4475 (N_4475,N_4367,N_4368);
nand U4476 (N_4476,N_4366,N_4384);
nand U4477 (N_4477,N_4331,N_4262);
or U4478 (N_4478,N_4390,N_4276);
nor U4479 (N_4479,N_4371,N_4314);
or U4480 (N_4480,N_4280,N_4222);
nor U4481 (N_4481,N_4319,N_4259);
nand U4482 (N_4482,N_4270,N_4239);
nor U4483 (N_4483,N_4377,N_4362);
nand U4484 (N_4484,N_4238,N_4233);
or U4485 (N_4485,N_4208,N_4209);
xnor U4486 (N_4486,N_4297,N_4254);
and U4487 (N_4487,N_4300,N_4237);
nor U4488 (N_4488,N_4204,N_4289);
xor U4489 (N_4489,N_4337,N_4218);
and U4490 (N_4490,N_4272,N_4285);
nor U4491 (N_4491,N_4338,N_4339);
nor U4492 (N_4492,N_4374,N_4353);
nand U4493 (N_4493,N_4282,N_4359);
nand U4494 (N_4494,N_4253,N_4343);
or U4495 (N_4495,N_4385,N_4229);
and U4496 (N_4496,N_4399,N_4206);
nand U4497 (N_4497,N_4357,N_4252);
xor U4498 (N_4498,N_4380,N_4250);
nand U4499 (N_4499,N_4213,N_4301);
or U4500 (N_4500,N_4284,N_4215);
nor U4501 (N_4501,N_4381,N_4348);
nor U4502 (N_4502,N_4313,N_4291);
and U4503 (N_4503,N_4348,N_4275);
nor U4504 (N_4504,N_4225,N_4233);
nor U4505 (N_4505,N_4239,N_4373);
nand U4506 (N_4506,N_4238,N_4201);
nand U4507 (N_4507,N_4307,N_4284);
or U4508 (N_4508,N_4277,N_4356);
nand U4509 (N_4509,N_4206,N_4374);
and U4510 (N_4510,N_4386,N_4311);
nand U4511 (N_4511,N_4365,N_4227);
xnor U4512 (N_4512,N_4206,N_4267);
and U4513 (N_4513,N_4279,N_4218);
nor U4514 (N_4514,N_4270,N_4317);
xor U4515 (N_4515,N_4273,N_4298);
xor U4516 (N_4516,N_4391,N_4331);
or U4517 (N_4517,N_4386,N_4210);
and U4518 (N_4518,N_4394,N_4337);
and U4519 (N_4519,N_4261,N_4350);
nor U4520 (N_4520,N_4245,N_4217);
or U4521 (N_4521,N_4310,N_4293);
nor U4522 (N_4522,N_4285,N_4337);
xor U4523 (N_4523,N_4334,N_4321);
nor U4524 (N_4524,N_4298,N_4290);
nor U4525 (N_4525,N_4325,N_4326);
or U4526 (N_4526,N_4397,N_4218);
or U4527 (N_4527,N_4308,N_4394);
or U4528 (N_4528,N_4287,N_4209);
and U4529 (N_4529,N_4329,N_4303);
nor U4530 (N_4530,N_4243,N_4216);
or U4531 (N_4531,N_4314,N_4327);
or U4532 (N_4532,N_4360,N_4348);
nor U4533 (N_4533,N_4320,N_4232);
nand U4534 (N_4534,N_4389,N_4285);
nand U4535 (N_4535,N_4390,N_4364);
and U4536 (N_4536,N_4393,N_4345);
and U4537 (N_4537,N_4227,N_4391);
or U4538 (N_4538,N_4382,N_4299);
nor U4539 (N_4539,N_4233,N_4321);
and U4540 (N_4540,N_4392,N_4246);
nor U4541 (N_4541,N_4344,N_4319);
or U4542 (N_4542,N_4236,N_4378);
nor U4543 (N_4543,N_4323,N_4293);
and U4544 (N_4544,N_4394,N_4353);
and U4545 (N_4545,N_4236,N_4220);
or U4546 (N_4546,N_4270,N_4378);
and U4547 (N_4547,N_4388,N_4322);
or U4548 (N_4548,N_4350,N_4322);
or U4549 (N_4549,N_4370,N_4326);
nor U4550 (N_4550,N_4263,N_4338);
and U4551 (N_4551,N_4379,N_4344);
nor U4552 (N_4552,N_4363,N_4231);
nor U4553 (N_4553,N_4277,N_4206);
nand U4554 (N_4554,N_4296,N_4295);
or U4555 (N_4555,N_4304,N_4305);
xor U4556 (N_4556,N_4230,N_4329);
nor U4557 (N_4557,N_4209,N_4291);
nor U4558 (N_4558,N_4230,N_4269);
nand U4559 (N_4559,N_4313,N_4379);
nor U4560 (N_4560,N_4361,N_4271);
nor U4561 (N_4561,N_4212,N_4304);
or U4562 (N_4562,N_4291,N_4369);
and U4563 (N_4563,N_4298,N_4362);
nand U4564 (N_4564,N_4306,N_4324);
and U4565 (N_4565,N_4277,N_4212);
and U4566 (N_4566,N_4295,N_4255);
and U4567 (N_4567,N_4287,N_4238);
nand U4568 (N_4568,N_4235,N_4211);
or U4569 (N_4569,N_4344,N_4313);
nor U4570 (N_4570,N_4387,N_4319);
nor U4571 (N_4571,N_4274,N_4324);
or U4572 (N_4572,N_4243,N_4246);
or U4573 (N_4573,N_4271,N_4283);
and U4574 (N_4574,N_4323,N_4267);
and U4575 (N_4575,N_4203,N_4242);
nand U4576 (N_4576,N_4278,N_4266);
nor U4577 (N_4577,N_4313,N_4270);
or U4578 (N_4578,N_4299,N_4342);
and U4579 (N_4579,N_4207,N_4364);
or U4580 (N_4580,N_4204,N_4377);
nor U4581 (N_4581,N_4271,N_4376);
or U4582 (N_4582,N_4230,N_4255);
nor U4583 (N_4583,N_4237,N_4314);
nor U4584 (N_4584,N_4248,N_4375);
and U4585 (N_4585,N_4379,N_4228);
or U4586 (N_4586,N_4247,N_4343);
or U4587 (N_4587,N_4391,N_4258);
and U4588 (N_4588,N_4376,N_4364);
xor U4589 (N_4589,N_4297,N_4265);
nand U4590 (N_4590,N_4237,N_4366);
or U4591 (N_4591,N_4399,N_4311);
nand U4592 (N_4592,N_4212,N_4251);
xnor U4593 (N_4593,N_4218,N_4214);
nor U4594 (N_4594,N_4323,N_4311);
or U4595 (N_4595,N_4357,N_4381);
nor U4596 (N_4596,N_4225,N_4314);
and U4597 (N_4597,N_4338,N_4354);
and U4598 (N_4598,N_4205,N_4375);
nand U4599 (N_4599,N_4238,N_4395);
nand U4600 (N_4600,N_4439,N_4457);
nor U4601 (N_4601,N_4442,N_4423);
nand U4602 (N_4602,N_4488,N_4407);
or U4603 (N_4603,N_4471,N_4489);
nor U4604 (N_4604,N_4593,N_4436);
xor U4605 (N_4605,N_4472,N_4557);
nor U4606 (N_4606,N_4404,N_4470);
nor U4607 (N_4607,N_4562,N_4441);
and U4608 (N_4608,N_4577,N_4554);
or U4609 (N_4609,N_4418,N_4569);
nand U4610 (N_4610,N_4549,N_4579);
nor U4611 (N_4611,N_4496,N_4513);
nor U4612 (N_4612,N_4455,N_4479);
and U4613 (N_4613,N_4448,N_4464);
xnor U4614 (N_4614,N_4490,N_4500);
nand U4615 (N_4615,N_4552,N_4403);
nand U4616 (N_4616,N_4440,N_4461);
nor U4617 (N_4617,N_4570,N_4486);
xor U4618 (N_4618,N_4466,N_4529);
nor U4619 (N_4619,N_4463,N_4447);
nor U4620 (N_4620,N_4428,N_4477);
nand U4621 (N_4621,N_4419,N_4583);
nand U4622 (N_4622,N_4484,N_4532);
nand U4623 (N_4623,N_4411,N_4521);
xor U4624 (N_4624,N_4481,N_4467);
xor U4625 (N_4625,N_4434,N_4528);
and U4626 (N_4626,N_4426,N_4497);
nor U4627 (N_4627,N_4543,N_4525);
or U4628 (N_4628,N_4491,N_4402);
nor U4629 (N_4629,N_4417,N_4582);
nand U4630 (N_4630,N_4526,N_4591);
nor U4631 (N_4631,N_4504,N_4433);
and U4632 (N_4632,N_4506,N_4572);
nor U4633 (N_4633,N_4546,N_4573);
nor U4634 (N_4634,N_4444,N_4533);
and U4635 (N_4635,N_4435,N_4553);
nand U4636 (N_4636,N_4548,N_4415);
nor U4637 (N_4637,N_4503,N_4469);
and U4638 (N_4638,N_4502,N_4421);
nor U4639 (N_4639,N_4587,N_4485);
and U4640 (N_4640,N_4564,N_4429);
nand U4641 (N_4641,N_4537,N_4509);
xor U4642 (N_4642,N_4483,N_4515);
and U4643 (N_4643,N_4589,N_4535);
nand U4644 (N_4644,N_4530,N_4517);
nand U4645 (N_4645,N_4556,N_4401);
or U4646 (N_4646,N_4598,N_4599);
or U4647 (N_4647,N_4539,N_4494);
and U4648 (N_4648,N_4476,N_4545);
nand U4649 (N_4649,N_4510,N_4406);
xor U4650 (N_4650,N_4422,N_4498);
nand U4651 (N_4651,N_4424,N_4427);
and U4652 (N_4652,N_4495,N_4409);
nand U4653 (N_4653,N_4516,N_4459);
nor U4654 (N_4654,N_4446,N_4437);
and U4655 (N_4655,N_4578,N_4473);
nand U4656 (N_4656,N_4452,N_4468);
xnor U4657 (N_4657,N_4478,N_4561);
xnor U4658 (N_4658,N_4514,N_4499);
or U4659 (N_4659,N_4487,N_4560);
and U4660 (N_4660,N_4534,N_4450);
nand U4661 (N_4661,N_4585,N_4453);
and U4662 (N_4662,N_4460,N_4522);
nand U4663 (N_4663,N_4462,N_4480);
xor U4664 (N_4664,N_4438,N_4527);
nor U4665 (N_4665,N_4400,N_4405);
xor U4666 (N_4666,N_4542,N_4474);
xor U4667 (N_4667,N_4465,N_4408);
and U4668 (N_4668,N_4568,N_4416);
nor U4669 (N_4669,N_4493,N_4508);
nand U4670 (N_4670,N_4586,N_4511);
xor U4671 (N_4671,N_4584,N_4596);
and U4672 (N_4672,N_4445,N_4576);
and U4673 (N_4673,N_4536,N_4443);
or U4674 (N_4674,N_4410,N_4482);
nand U4675 (N_4675,N_4430,N_4431);
nand U4676 (N_4676,N_4512,N_4524);
or U4677 (N_4677,N_4597,N_4432);
or U4678 (N_4678,N_4414,N_4551);
or U4679 (N_4679,N_4501,N_4425);
or U4680 (N_4680,N_4538,N_4592);
and U4681 (N_4681,N_4505,N_4567);
or U4682 (N_4682,N_4547,N_4531);
nand U4683 (N_4683,N_4594,N_4541);
nand U4684 (N_4684,N_4590,N_4550);
and U4685 (N_4685,N_4458,N_4523);
nor U4686 (N_4686,N_4575,N_4412);
nor U4687 (N_4687,N_4544,N_4580);
nor U4688 (N_4688,N_4571,N_4540);
or U4689 (N_4689,N_4475,N_4456);
nand U4690 (N_4690,N_4559,N_4492);
or U4691 (N_4691,N_4565,N_4588);
or U4692 (N_4692,N_4413,N_4581);
or U4693 (N_4693,N_4566,N_4449);
nand U4694 (N_4694,N_4574,N_4454);
xor U4695 (N_4695,N_4451,N_4520);
nand U4696 (N_4696,N_4595,N_4518);
nand U4697 (N_4697,N_4563,N_4558);
and U4698 (N_4698,N_4519,N_4555);
or U4699 (N_4699,N_4507,N_4420);
nand U4700 (N_4700,N_4574,N_4461);
nor U4701 (N_4701,N_4464,N_4414);
and U4702 (N_4702,N_4474,N_4520);
nor U4703 (N_4703,N_4405,N_4447);
nand U4704 (N_4704,N_4427,N_4444);
or U4705 (N_4705,N_4563,N_4415);
or U4706 (N_4706,N_4452,N_4579);
xnor U4707 (N_4707,N_4422,N_4559);
nor U4708 (N_4708,N_4526,N_4427);
nor U4709 (N_4709,N_4421,N_4423);
nand U4710 (N_4710,N_4458,N_4533);
or U4711 (N_4711,N_4443,N_4505);
nor U4712 (N_4712,N_4489,N_4531);
nor U4713 (N_4713,N_4510,N_4409);
and U4714 (N_4714,N_4426,N_4428);
or U4715 (N_4715,N_4434,N_4545);
xnor U4716 (N_4716,N_4430,N_4450);
or U4717 (N_4717,N_4550,N_4413);
or U4718 (N_4718,N_4540,N_4461);
or U4719 (N_4719,N_4475,N_4479);
or U4720 (N_4720,N_4539,N_4536);
nor U4721 (N_4721,N_4541,N_4575);
nor U4722 (N_4722,N_4540,N_4546);
xor U4723 (N_4723,N_4513,N_4453);
nor U4724 (N_4724,N_4501,N_4560);
nor U4725 (N_4725,N_4452,N_4560);
nor U4726 (N_4726,N_4519,N_4469);
nor U4727 (N_4727,N_4449,N_4483);
nand U4728 (N_4728,N_4542,N_4410);
and U4729 (N_4729,N_4501,N_4587);
nand U4730 (N_4730,N_4419,N_4496);
and U4731 (N_4731,N_4560,N_4442);
and U4732 (N_4732,N_4413,N_4419);
nand U4733 (N_4733,N_4550,N_4537);
or U4734 (N_4734,N_4440,N_4503);
nand U4735 (N_4735,N_4447,N_4473);
or U4736 (N_4736,N_4456,N_4438);
or U4737 (N_4737,N_4571,N_4498);
nor U4738 (N_4738,N_4592,N_4402);
and U4739 (N_4739,N_4494,N_4586);
nor U4740 (N_4740,N_4590,N_4441);
nor U4741 (N_4741,N_4476,N_4578);
nor U4742 (N_4742,N_4514,N_4533);
nand U4743 (N_4743,N_4585,N_4489);
and U4744 (N_4744,N_4564,N_4524);
and U4745 (N_4745,N_4596,N_4459);
nand U4746 (N_4746,N_4597,N_4498);
and U4747 (N_4747,N_4401,N_4509);
nor U4748 (N_4748,N_4416,N_4519);
xor U4749 (N_4749,N_4442,N_4430);
and U4750 (N_4750,N_4406,N_4455);
xor U4751 (N_4751,N_4539,N_4524);
and U4752 (N_4752,N_4404,N_4432);
xor U4753 (N_4753,N_4523,N_4405);
nand U4754 (N_4754,N_4455,N_4558);
nor U4755 (N_4755,N_4508,N_4528);
nand U4756 (N_4756,N_4476,N_4519);
or U4757 (N_4757,N_4468,N_4465);
or U4758 (N_4758,N_4432,N_4423);
nand U4759 (N_4759,N_4572,N_4531);
nand U4760 (N_4760,N_4542,N_4400);
or U4761 (N_4761,N_4448,N_4474);
or U4762 (N_4762,N_4580,N_4483);
or U4763 (N_4763,N_4513,N_4448);
or U4764 (N_4764,N_4554,N_4543);
and U4765 (N_4765,N_4484,N_4410);
or U4766 (N_4766,N_4500,N_4426);
nand U4767 (N_4767,N_4540,N_4460);
or U4768 (N_4768,N_4468,N_4426);
xnor U4769 (N_4769,N_4532,N_4512);
and U4770 (N_4770,N_4459,N_4410);
nand U4771 (N_4771,N_4540,N_4568);
nor U4772 (N_4772,N_4553,N_4495);
and U4773 (N_4773,N_4445,N_4439);
nand U4774 (N_4774,N_4410,N_4421);
nor U4775 (N_4775,N_4525,N_4479);
xnor U4776 (N_4776,N_4426,N_4415);
or U4777 (N_4777,N_4559,N_4582);
nand U4778 (N_4778,N_4562,N_4497);
nor U4779 (N_4779,N_4469,N_4450);
and U4780 (N_4780,N_4545,N_4549);
nand U4781 (N_4781,N_4566,N_4428);
nor U4782 (N_4782,N_4482,N_4495);
nor U4783 (N_4783,N_4431,N_4564);
or U4784 (N_4784,N_4483,N_4520);
xnor U4785 (N_4785,N_4425,N_4469);
or U4786 (N_4786,N_4541,N_4422);
nand U4787 (N_4787,N_4439,N_4492);
nor U4788 (N_4788,N_4521,N_4528);
or U4789 (N_4789,N_4477,N_4408);
or U4790 (N_4790,N_4522,N_4586);
or U4791 (N_4791,N_4421,N_4528);
nor U4792 (N_4792,N_4404,N_4521);
or U4793 (N_4793,N_4475,N_4536);
and U4794 (N_4794,N_4496,N_4491);
nand U4795 (N_4795,N_4508,N_4572);
nor U4796 (N_4796,N_4404,N_4549);
or U4797 (N_4797,N_4536,N_4483);
and U4798 (N_4798,N_4438,N_4469);
or U4799 (N_4799,N_4534,N_4440);
nor U4800 (N_4800,N_4745,N_4749);
xnor U4801 (N_4801,N_4698,N_4769);
or U4802 (N_4802,N_4623,N_4649);
nor U4803 (N_4803,N_4606,N_4638);
nor U4804 (N_4804,N_4776,N_4701);
or U4805 (N_4805,N_4619,N_4788);
or U4806 (N_4806,N_4716,N_4611);
or U4807 (N_4807,N_4637,N_4628);
and U4808 (N_4808,N_4683,N_4697);
and U4809 (N_4809,N_4641,N_4636);
nand U4810 (N_4810,N_4651,N_4672);
nand U4811 (N_4811,N_4746,N_4753);
or U4812 (N_4812,N_4705,N_4694);
or U4813 (N_4813,N_4614,N_4775);
nand U4814 (N_4814,N_4731,N_4740);
or U4815 (N_4815,N_4782,N_4799);
nand U4816 (N_4816,N_4603,N_4659);
or U4817 (N_4817,N_4626,N_4657);
nor U4818 (N_4818,N_4772,N_4765);
nand U4819 (N_4819,N_4787,N_4752);
or U4820 (N_4820,N_4653,N_4785);
and U4821 (N_4821,N_4722,N_4767);
or U4822 (N_4822,N_4681,N_4635);
or U4823 (N_4823,N_4784,N_4631);
and U4824 (N_4824,N_4660,N_4607);
nor U4825 (N_4825,N_4691,N_4711);
or U4826 (N_4826,N_4630,N_4728);
or U4827 (N_4827,N_4747,N_4674);
and U4828 (N_4828,N_4652,N_4664);
nor U4829 (N_4829,N_4758,N_4602);
or U4830 (N_4830,N_4629,N_4798);
or U4831 (N_4831,N_4646,N_4621);
xor U4832 (N_4832,N_4726,N_4710);
nand U4833 (N_4833,N_4750,N_4778);
and U4834 (N_4834,N_4755,N_4645);
nand U4835 (N_4835,N_4719,N_4790);
and U4836 (N_4836,N_4632,N_4610);
nor U4837 (N_4837,N_4791,N_4770);
or U4838 (N_4838,N_4690,N_4618);
nor U4839 (N_4839,N_4760,N_4712);
nor U4840 (N_4840,N_4612,N_4615);
or U4841 (N_4841,N_4634,N_4643);
or U4842 (N_4842,N_4763,N_4617);
and U4843 (N_4843,N_4721,N_4748);
nand U4844 (N_4844,N_4771,N_4642);
xor U4845 (N_4845,N_4743,N_4759);
or U4846 (N_4846,N_4756,N_4686);
or U4847 (N_4847,N_4700,N_4715);
and U4848 (N_4848,N_4727,N_4709);
or U4849 (N_4849,N_4673,N_4622);
nor U4850 (N_4850,N_4723,N_4666);
nand U4851 (N_4851,N_4768,N_4640);
or U4852 (N_4852,N_4609,N_4624);
or U4853 (N_4853,N_4796,N_4608);
nand U4854 (N_4854,N_4764,N_4704);
nand U4855 (N_4855,N_4786,N_4751);
and U4856 (N_4856,N_4739,N_4713);
or U4857 (N_4857,N_4761,N_4658);
nor U4858 (N_4858,N_4792,N_4601);
nand U4859 (N_4859,N_4669,N_4605);
and U4860 (N_4860,N_4766,N_4696);
nand U4861 (N_4861,N_4670,N_4708);
and U4862 (N_4862,N_4667,N_4647);
nand U4863 (N_4863,N_4780,N_4720);
nor U4864 (N_4864,N_4600,N_4692);
and U4865 (N_4865,N_4687,N_4794);
and U4866 (N_4866,N_4777,N_4702);
nor U4867 (N_4867,N_4736,N_4718);
nand U4868 (N_4868,N_4733,N_4774);
nand U4869 (N_4869,N_4644,N_4783);
nand U4870 (N_4870,N_4773,N_4685);
or U4871 (N_4871,N_4679,N_4734);
nand U4872 (N_4872,N_4724,N_4689);
and U4873 (N_4873,N_4677,N_4699);
or U4874 (N_4874,N_4789,N_4662);
nor U4875 (N_4875,N_4695,N_4671);
or U4876 (N_4876,N_4795,N_4714);
or U4877 (N_4877,N_4650,N_4735);
or U4878 (N_4878,N_4729,N_4633);
nand U4879 (N_4879,N_4741,N_4738);
or U4880 (N_4880,N_4604,N_4656);
xor U4881 (N_4881,N_4627,N_4639);
or U4882 (N_4882,N_4779,N_4693);
and U4883 (N_4883,N_4754,N_4676);
nand U4884 (N_4884,N_4616,N_4717);
nor U4885 (N_4885,N_4797,N_4668);
nor U4886 (N_4886,N_4757,N_4732);
nor U4887 (N_4887,N_4793,N_4625);
nand U4888 (N_4888,N_4707,N_4706);
nor U4889 (N_4889,N_4675,N_4688);
nor U4890 (N_4890,N_4737,N_4742);
xnor U4891 (N_4891,N_4648,N_4703);
and U4892 (N_4892,N_4663,N_4665);
nor U4893 (N_4893,N_4655,N_4620);
nand U4894 (N_4894,N_4682,N_4613);
nor U4895 (N_4895,N_4654,N_4762);
or U4896 (N_4896,N_4678,N_4730);
nor U4897 (N_4897,N_4661,N_4744);
xor U4898 (N_4898,N_4781,N_4680);
or U4899 (N_4899,N_4725,N_4684);
xor U4900 (N_4900,N_4699,N_4709);
nor U4901 (N_4901,N_4677,N_4642);
nor U4902 (N_4902,N_4761,N_4749);
nand U4903 (N_4903,N_4799,N_4779);
and U4904 (N_4904,N_4756,N_4770);
xor U4905 (N_4905,N_4705,N_4627);
and U4906 (N_4906,N_4723,N_4688);
xor U4907 (N_4907,N_4618,N_4727);
and U4908 (N_4908,N_4741,N_4674);
and U4909 (N_4909,N_4795,N_4653);
or U4910 (N_4910,N_4720,N_4705);
nand U4911 (N_4911,N_4761,N_4707);
xor U4912 (N_4912,N_4726,N_4684);
nor U4913 (N_4913,N_4716,N_4653);
or U4914 (N_4914,N_4720,N_4630);
and U4915 (N_4915,N_4757,N_4687);
nand U4916 (N_4916,N_4613,N_4655);
nand U4917 (N_4917,N_4701,N_4744);
nor U4918 (N_4918,N_4620,N_4731);
nand U4919 (N_4919,N_4662,N_4794);
and U4920 (N_4920,N_4605,N_4703);
nand U4921 (N_4921,N_4680,N_4762);
nor U4922 (N_4922,N_4717,N_4613);
nand U4923 (N_4923,N_4745,N_4728);
nor U4924 (N_4924,N_4745,N_4687);
and U4925 (N_4925,N_4777,N_4715);
xnor U4926 (N_4926,N_4709,N_4772);
and U4927 (N_4927,N_4628,N_4636);
nand U4928 (N_4928,N_4778,N_4793);
nand U4929 (N_4929,N_4712,N_4779);
nor U4930 (N_4930,N_4716,N_4605);
nand U4931 (N_4931,N_4646,N_4607);
nor U4932 (N_4932,N_4644,N_4743);
or U4933 (N_4933,N_4762,N_4684);
and U4934 (N_4934,N_4797,N_4657);
and U4935 (N_4935,N_4622,N_4732);
or U4936 (N_4936,N_4720,N_4743);
xor U4937 (N_4937,N_4777,N_4728);
nor U4938 (N_4938,N_4716,N_4683);
nor U4939 (N_4939,N_4611,N_4633);
nand U4940 (N_4940,N_4665,N_4684);
nand U4941 (N_4941,N_4693,N_4688);
nor U4942 (N_4942,N_4696,N_4611);
or U4943 (N_4943,N_4725,N_4788);
nand U4944 (N_4944,N_4781,N_4711);
or U4945 (N_4945,N_4622,N_4709);
nor U4946 (N_4946,N_4624,N_4762);
xor U4947 (N_4947,N_4786,N_4712);
and U4948 (N_4948,N_4771,N_4756);
xor U4949 (N_4949,N_4786,N_4777);
nand U4950 (N_4950,N_4693,N_4762);
xnor U4951 (N_4951,N_4634,N_4770);
nand U4952 (N_4952,N_4676,N_4625);
or U4953 (N_4953,N_4765,N_4687);
or U4954 (N_4954,N_4688,N_4742);
or U4955 (N_4955,N_4640,N_4737);
nand U4956 (N_4956,N_4677,N_4662);
nand U4957 (N_4957,N_4646,N_4623);
and U4958 (N_4958,N_4787,N_4692);
nand U4959 (N_4959,N_4740,N_4730);
or U4960 (N_4960,N_4759,N_4685);
or U4961 (N_4961,N_4752,N_4637);
nand U4962 (N_4962,N_4683,N_4767);
nand U4963 (N_4963,N_4704,N_4620);
or U4964 (N_4964,N_4652,N_4757);
nor U4965 (N_4965,N_4646,N_4709);
nand U4966 (N_4966,N_4708,N_4752);
nand U4967 (N_4967,N_4718,N_4609);
or U4968 (N_4968,N_4715,N_4607);
or U4969 (N_4969,N_4633,N_4734);
or U4970 (N_4970,N_4784,N_4728);
nor U4971 (N_4971,N_4660,N_4761);
nand U4972 (N_4972,N_4647,N_4686);
xnor U4973 (N_4973,N_4669,N_4699);
nand U4974 (N_4974,N_4792,N_4744);
or U4975 (N_4975,N_4633,N_4762);
or U4976 (N_4976,N_4632,N_4777);
xnor U4977 (N_4977,N_4741,N_4689);
nand U4978 (N_4978,N_4719,N_4752);
nor U4979 (N_4979,N_4723,N_4719);
and U4980 (N_4980,N_4722,N_4698);
nor U4981 (N_4981,N_4781,N_4749);
nand U4982 (N_4982,N_4628,N_4632);
and U4983 (N_4983,N_4604,N_4637);
and U4984 (N_4984,N_4701,N_4601);
or U4985 (N_4985,N_4683,N_4616);
xor U4986 (N_4986,N_4771,N_4628);
nand U4987 (N_4987,N_4758,N_4628);
nor U4988 (N_4988,N_4632,N_4734);
and U4989 (N_4989,N_4788,N_4773);
xnor U4990 (N_4990,N_4683,N_4605);
nand U4991 (N_4991,N_4777,N_4681);
xnor U4992 (N_4992,N_4752,N_4638);
nor U4993 (N_4993,N_4702,N_4648);
nand U4994 (N_4994,N_4688,N_4710);
xnor U4995 (N_4995,N_4737,N_4791);
or U4996 (N_4996,N_4644,N_4621);
xor U4997 (N_4997,N_4720,N_4611);
nor U4998 (N_4998,N_4708,N_4783);
nor U4999 (N_4999,N_4693,N_4626);
nor U5000 (N_5000,N_4835,N_4984);
nor U5001 (N_5001,N_4958,N_4902);
or U5002 (N_5002,N_4881,N_4855);
and U5003 (N_5003,N_4811,N_4986);
nor U5004 (N_5004,N_4901,N_4946);
nor U5005 (N_5005,N_4842,N_4845);
xnor U5006 (N_5006,N_4955,N_4972);
nand U5007 (N_5007,N_4915,N_4836);
nand U5008 (N_5008,N_4941,N_4945);
or U5009 (N_5009,N_4954,N_4913);
and U5010 (N_5010,N_4866,N_4854);
or U5011 (N_5011,N_4892,N_4921);
nand U5012 (N_5012,N_4805,N_4995);
xnor U5013 (N_5013,N_4815,N_4825);
nor U5014 (N_5014,N_4821,N_4844);
nand U5015 (N_5015,N_4814,N_4887);
and U5016 (N_5016,N_4977,N_4857);
xor U5017 (N_5017,N_4970,N_4834);
nand U5018 (N_5018,N_4940,N_4817);
or U5019 (N_5019,N_4904,N_4885);
nor U5020 (N_5020,N_4871,N_4883);
nor U5021 (N_5021,N_4917,N_4868);
nor U5022 (N_5022,N_4819,N_4846);
nand U5023 (N_5023,N_4994,N_4879);
or U5024 (N_5024,N_4967,N_4824);
or U5025 (N_5025,N_4907,N_4826);
and U5026 (N_5026,N_4830,N_4882);
nand U5027 (N_5027,N_4873,N_4850);
nor U5028 (N_5028,N_4959,N_4861);
nand U5029 (N_5029,N_4867,N_4912);
or U5030 (N_5030,N_4918,N_4849);
nand U5031 (N_5031,N_4804,N_4860);
nand U5032 (N_5032,N_4828,N_4953);
xnor U5033 (N_5033,N_4812,N_4999);
or U5034 (N_5034,N_4898,N_4943);
and U5035 (N_5035,N_4932,N_4859);
nand U5036 (N_5036,N_4964,N_4910);
nor U5037 (N_5037,N_4820,N_4878);
or U5038 (N_5038,N_4997,N_4916);
nand U5039 (N_5039,N_4848,N_4809);
nand U5040 (N_5040,N_4852,N_4800);
or U5041 (N_5041,N_4998,N_4890);
nor U5042 (N_5042,N_4993,N_4937);
nor U5043 (N_5043,N_4982,N_4990);
nor U5044 (N_5044,N_4831,N_4968);
nor U5045 (N_5045,N_4875,N_4876);
xnor U5046 (N_5046,N_4987,N_4919);
nor U5047 (N_5047,N_4864,N_4823);
or U5048 (N_5048,N_4971,N_4957);
xor U5049 (N_5049,N_4894,N_4837);
nand U5050 (N_5050,N_4806,N_4818);
nor U5051 (N_5051,N_4874,N_4951);
nor U5052 (N_5052,N_4988,N_4802);
or U5053 (N_5053,N_4803,N_4979);
or U5054 (N_5054,N_4838,N_4960);
nand U5055 (N_5055,N_4985,N_4925);
and U5056 (N_5056,N_4896,N_4923);
or U5057 (N_5057,N_4914,N_4851);
and U5058 (N_5058,N_4942,N_4980);
nand U5059 (N_5059,N_4939,N_4973);
nor U5060 (N_5060,N_4978,N_4862);
nor U5061 (N_5061,N_4928,N_4911);
xor U5062 (N_5062,N_4900,N_4930);
or U5063 (N_5063,N_4888,N_4889);
nor U5064 (N_5064,N_4975,N_4926);
xnor U5065 (N_5065,N_4807,N_4976);
nand U5066 (N_5066,N_4870,N_4922);
nand U5067 (N_5067,N_4991,N_4858);
nand U5068 (N_5068,N_4938,N_4969);
and U5069 (N_5069,N_4965,N_4880);
nor U5070 (N_5070,N_4933,N_4983);
nor U5071 (N_5071,N_4936,N_4853);
nor U5072 (N_5072,N_4952,N_4948);
nor U5073 (N_5073,N_4961,N_4865);
xor U5074 (N_5074,N_4956,N_4908);
nand U5075 (N_5075,N_4931,N_4839);
and U5076 (N_5076,N_4895,N_4863);
nand U5077 (N_5077,N_4877,N_4905);
nand U5078 (N_5078,N_4893,N_4927);
or U5079 (N_5079,N_4841,N_4899);
nor U5080 (N_5080,N_4884,N_4924);
or U5081 (N_5081,N_4929,N_4909);
or U5082 (N_5082,N_4816,N_4872);
nor U5083 (N_5083,N_4840,N_4974);
or U5084 (N_5084,N_4869,N_4810);
nand U5085 (N_5085,N_4963,N_4822);
and U5086 (N_5086,N_4833,N_4935);
xor U5087 (N_5087,N_4808,N_4934);
nor U5088 (N_5088,N_4920,N_4801);
nor U5089 (N_5089,N_4891,N_4856);
and U5090 (N_5090,N_4949,N_4832);
nor U5091 (N_5091,N_4847,N_4996);
or U5092 (N_5092,N_4813,N_4962);
or U5093 (N_5093,N_4897,N_4947);
or U5094 (N_5094,N_4944,N_4886);
nand U5095 (N_5095,N_4829,N_4906);
nand U5096 (N_5096,N_4981,N_4843);
and U5097 (N_5097,N_4827,N_4989);
or U5098 (N_5098,N_4950,N_4992);
nand U5099 (N_5099,N_4903,N_4966);
nand U5100 (N_5100,N_4917,N_4915);
or U5101 (N_5101,N_4913,N_4982);
and U5102 (N_5102,N_4849,N_4827);
and U5103 (N_5103,N_4951,N_4922);
nand U5104 (N_5104,N_4953,N_4980);
xor U5105 (N_5105,N_4805,N_4836);
and U5106 (N_5106,N_4977,N_4869);
nand U5107 (N_5107,N_4938,N_4930);
nor U5108 (N_5108,N_4966,N_4971);
or U5109 (N_5109,N_4930,N_4924);
nand U5110 (N_5110,N_4949,N_4962);
nand U5111 (N_5111,N_4836,N_4914);
or U5112 (N_5112,N_4820,N_4868);
nor U5113 (N_5113,N_4933,N_4998);
or U5114 (N_5114,N_4929,N_4838);
nand U5115 (N_5115,N_4844,N_4842);
and U5116 (N_5116,N_4976,N_4932);
or U5117 (N_5117,N_4886,N_4893);
nand U5118 (N_5118,N_4911,N_4949);
nor U5119 (N_5119,N_4919,N_4968);
xnor U5120 (N_5120,N_4904,N_4983);
and U5121 (N_5121,N_4884,N_4992);
or U5122 (N_5122,N_4866,N_4888);
and U5123 (N_5123,N_4989,N_4865);
or U5124 (N_5124,N_4958,N_4803);
or U5125 (N_5125,N_4918,N_4837);
xor U5126 (N_5126,N_4982,N_4932);
nor U5127 (N_5127,N_4811,N_4911);
nor U5128 (N_5128,N_4806,N_4805);
or U5129 (N_5129,N_4883,N_4947);
xor U5130 (N_5130,N_4924,N_4895);
or U5131 (N_5131,N_4924,N_4804);
nor U5132 (N_5132,N_4808,N_4811);
nand U5133 (N_5133,N_4879,N_4909);
and U5134 (N_5134,N_4953,N_4915);
nor U5135 (N_5135,N_4891,N_4992);
nor U5136 (N_5136,N_4893,N_4973);
and U5137 (N_5137,N_4938,N_4956);
or U5138 (N_5138,N_4831,N_4812);
xor U5139 (N_5139,N_4868,N_4927);
or U5140 (N_5140,N_4840,N_4812);
nand U5141 (N_5141,N_4954,N_4957);
nor U5142 (N_5142,N_4960,N_4978);
and U5143 (N_5143,N_4839,N_4892);
nor U5144 (N_5144,N_4977,N_4985);
nor U5145 (N_5145,N_4817,N_4910);
nand U5146 (N_5146,N_4988,N_4875);
and U5147 (N_5147,N_4864,N_4832);
xor U5148 (N_5148,N_4848,N_4801);
nor U5149 (N_5149,N_4976,N_4862);
and U5150 (N_5150,N_4899,N_4959);
and U5151 (N_5151,N_4864,N_4959);
or U5152 (N_5152,N_4961,N_4947);
nand U5153 (N_5153,N_4979,N_4982);
or U5154 (N_5154,N_4875,N_4949);
or U5155 (N_5155,N_4892,N_4882);
and U5156 (N_5156,N_4934,N_4886);
or U5157 (N_5157,N_4955,N_4855);
nand U5158 (N_5158,N_4986,N_4981);
or U5159 (N_5159,N_4854,N_4862);
xnor U5160 (N_5160,N_4963,N_4960);
or U5161 (N_5161,N_4882,N_4802);
nor U5162 (N_5162,N_4994,N_4801);
nand U5163 (N_5163,N_4804,N_4851);
nand U5164 (N_5164,N_4928,N_4868);
nor U5165 (N_5165,N_4810,N_4828);
and U5166 (N_5166,N_4951,N_4852);
and U5167 (N_5167,N_4829,N_4984);
nor U5168 (N_5168,N_4859,N_4861);
nand U5169 (N_5169,N_4857,N_4873);
or U5170 (N_5170,N_4955,N_4815);
nor U5171 (N_5171,N_4946,N_4925);
or U5172 (N_5172,N_4830,N_4870);
or U5173 (N_5173,N_4923,N_4961);
or U5174 (N_5174,N_4868,N_4932);
nand U5175 (N_5175,N_4904,N_4996);
nand U5176 (N_5176,N_4899,N_4988);
nand U5177 (N_5177,N_4957,N_4821);
nand U5178 (N_5178,N_4988,N_4800);
nor U5179 (N_5179,N_4968,N_4887);
or U5180 (N_5180,N_4870,N_4973);
nand U5181 (N_5181,N_4941,N_4970);
and U5182 (N_5182,N_4970,N_4898);
or U5183 (N_5183,N_4957,N_4881);
xnor U5184 (N_5184,N_4803,N_4981);
nand U5185 (N_5185,N_4804,N_4813);
nor U5186 (N_5186,N_4825,N_4866);
xnor U5187 (N_5187,N_4887,N_4800);
nand U5188 (N_5188,N_4921,N_4930);
nand U5189 (N_5189,N_4994,N_4850);
nor U5190 (N_5190,N_4935,N_4807);
or U5191 (N_5191,N_4866,N_4900);
xnor U5192 (N_5192,N_4892,N_4867);
nand U5193 (N_5193,N_4974,N_4819);
and U5194 (N_5194,N_4927,N_4985);
xor U5195 (N_5195,N_4902,N_4818);
xnor U5196 (N_5196,N_4984,N_4838);
nor U5197 (N_5197,N_4866,N_4818);
nand U5198 (N_5198,N_4983,N_4908);
and U5199 (N_5199,N_4846,N_4916);
or U5200 (N_5200,N_5168,N_5129);
and U5201 (N_5201,N_5182,N_5166);
nand U5202 (N_5202,N_5077,N_5091);
or U5203 (N_5203,N_5163,N_5178);
nand U5204 (N_5204,N_5044,N_5081);
nor U5205 (N_5205,N_5148,N_5058);
and U5206 (N_5206,N_5118,N_5007);
nand U5207 (N_5207,N_5169,N_5160);
or U5208 (N_5208,N_5053,N_5167);
nor U5209 (N_5209,N_5138,N_5088);
nor U5210 (N_5210,N_5135,N_5037);
xor U5211 (N_5211,N_5072,N_5032);
nand U5212 (N_5212,N_5100,N_5192);
nand U5213 (N_5213,N_5198,N_5185);
nor U5214 (N_5214,N_5063,N_5013);
xnor U5215 (N_5215,N_5019,N_5082);
nand U5216 (N_5216,N_5128,N_5174);
nand U5217 (N_5217,N_5045,N_5107);
and U5218 (N_5218,N_5051,N_5068);
nor U5219 (N_5219,N_5121,N_5078);
and U5220 (N_5220,N_5008,N_5193);
or U5221 (N_5221,N_5015,N_5035);
and U5222 (N_5222,N_5097,N_5086);
xnor U5223 (N_5223,N_5122,N_5130);
nor U5224 (N_5224,N_5162,N_5031);
nor U5225 (N_5225,N_5038,N_5009);
or U5226 (N_5226,N_5014,N_5164);
and U5227 (N_5227,N_5124,N_5188);
nand U5228 (N_5228,N_5036,N_5069);
nor U5229 (N_5229,N_5048,N_5143);
or U5230 (N_5230,N_5057,N_5012);
nand U5231 (N_5231,N_5060,N_5011);
nand U5232 (N_5232,N_5133,N_5020);
nand U5233 (N_5233,N_5150,N_5125);
xor U5234 (N_5234,N_5056,N_5040);
and U5235 (N_5235,N_5176,N_5158);
xnor U5236 (N_5236,N_5111,N_5093);
and U5237 (N_5237,N_5183,N_5004);
or U5238 (N_5238,N_5084,N_5054);
and U5239 (N_5239,N_5151,N_5195);
nand U5240 (N_5240,N_5017,N_5075);
nor U5241 (N_5241,N_5179,N_5165);
nor U5242 (N_5242,N_5094,N_5085);
nor U5243 (N_5243,N_5117,N_5073);
nand U5244 (N_5244,N_5005,N_5025);
or U5245 (N_5245,N_5096,N_5123);
or U5246 (N_5246,N_5028,N_5119);
nand U5247 (N_5247,N_5024,N_5027);
and U5248 (N_5248,N_5062,N_5052);
and U5249 (N_5249,N_5142,N_5153);
nor U5250 (N_5250,N_5147,N_5199);
and U5251 (N_5251,N_5099,N_5194);
or U5252 (N_5252,N_5071,N_5149);
nand U5253 (N_5253,N_5172,N_5104);
and U5254 (N_5254,N_5144,N_5187);
or U5255 (N_5255,N_5070,N_5112);
nand U5256 (N_5256,N_5110,N_5113);
and U5257 (N_5257,N_5065,N_5136);
or U5258 (N_5258,N_5139,N_5173);
nand U5259 (N_5259,N_5115,N_5180);
nand U5260 (N_5260,N_5171,N_5146);
nor U5261 (N_5261,N_5114,N_5186);
or U5262 (N_5262,N_5102,N_5018);
or U5263 (N_5263,N_5154,N_5010);
and U5264 (N_5264,N_5022,N_5103);
and U5265 (N_5265,N_5034,N_5092);
nand U5266 (N_5266,N_5016,N_5109);
nor U5267 (N_5267,N_5067,N_5043);
or U5268 (N_5268,N_5152,N_5079);
nor U5269 (N_5269,N_5002,N_5064);
nand U5270 (N_5270,N_5159,N_5170);
nor U5271 (N_5271,N_5066,N_5105);
and U5272 (N_5272,N_5061,N_5098);
and U5273 (N_5273,N_5197,N_5050);
or U5274 (N_5274,N_5021,N_5145);
or U5275 (N_5275,N_5131,N_5181);
xor U5276 (N_5276,N_5120,N_5074);
nand U5277 (N_5277,N_5080,N_5196);
nor U5278 (N_5278,N_5029,N_5116);
and U5279 (N_5279,N_5055,N_5132);
and U5280 (N_5280,N_5189,N_5087);
nor U5281 (N_5281,N_5134,N_5190);
and U5282 (N_5282,N_5089,N_5042);
nor U5283 (N_5283,N_5106,N_5000);
nor U5284 (N_5284,N_5177,N_5191);
nor U5285 (N_5285,N_5001,N_5046);
and U5286 (N_5286,N_5095,N_5049);
or U5287 (N_5287,N_5127,N_5030);
nor U5288 (N_5288,N_5175,N_5108);
and U5289 (N_5289,N_5140,N_5047);
and U5290 (N_5290,N_5157,N_5083);
or U5291 (N_5291,N_5006,N_5137);
nand U5292 (N_5292,N_5033,N_5059);
and U5293 (N_5293,N_5023,N_5184);
nand U5294 (N_5294,N_5041,N_5155);
and U5295 (N_5295,N_5101,N_5141);
nand U5296 (N_5296,N_5090,N_5039);
or U5297 (N_5297,N_5003,N_5126);
and U5298 (N_5298,N_5156,N_5026);
or U5299 (N_5299,N_5076,N_5161);
and U5300 (N_5300,N_5063,N_5081);
nand U5301 (N_5301,N_5147,N_5162);
and U5302 (N_5302,N_5074,N_5047);
nor U5303 (N_5303,N_5080,N_5087);
nor U5304 (N_5304,N_5047,N_5188);
and U5305 (N_5305,N_5047,N_5191);
xor U5306 (N_5306,N_5120,N_5053);
nor U5307 (N_5307,N_5034,N_5181);
nand U5308 (N_5308,N_5042,N_5093);
nor U5309 (N_5309,N_5195,N_5138);
or U5310 (N_5310,N_5076,N_5172);
and U5311 (N_5311,N_5035,N_5149);
nand U5312 (N_5312,N_5027,N_5052);
nand U5313 (N_5313,N_5087,N_5061);
or U5314 (N_5314,N_5076,N_5146);
nor U5315 (N_5315,N_5183,N_5022);
nand U5316 (N_5316,N_5060,N_5138);
nor U5317 (N_5317,N_5071,N_5008);
nor U5318 (N_5318,N_5033,N_5046);
or U5319 (N_5319,N_5126,N_5046);
nor U5320 (N_5320,N_5078,N_5150);
nand U5321 (N_5321,N_5006,N_5168);
nor U5322 (N_5322,N_5056,N_5172);
and U5323 (N_5323,N_5033,N_5007);
nand U5324 (N_5324,N_5173,N_5015);
xnor U5325 (N_5325,N_5079,N_5109);
nor U5326 (N_5326,N_5133,N_5000);
and U5327 (N_5327,N_5131,N_5133);
or U5328 (N_5328,N_5181,N_5112);
nand U5329 (N_5329,N_5146,N_5108);
nor U5330 (N_5330,N_5071,N_5094);
and U5331 (N_5331,N_5139,N_5049);
xor U5332 (N_5332,N_5153,N_5033);
nand U5333 (N_5333,N_5153,N_5014);
nor U5334 (N_5334,N_5052,N_5078);
or U5335 (N_5335,N_5173,N_5025);
nand U5336 (N_5336,N_5102,N_5014);
and U5337 (N_5337,N_5016,N_5178);
or U5338 (N_5338,N_5122,N_5096);
and U5339 (N_5339,N_5045,N_5069);
xor U5340 (N_5340,N_5169,N_5012);
or U5341 (N_5341,N_5088,N_5116);
or U5342 (N_5342,N_5005,N_5010);
nand U5343 (N_5343,N_5155,N_5124);
nand U5344 (N_5344,N_5006,N_5034);
nor U5345 (N_5345,N_5064,N_5127);
nand U5346 (N_5346,N_5002,N_5196);
nor U5347 (N_5347,N_5117,N_5087);
nand U5348 (N_5348,N_5077,N_5020);
nor U5349 (N_5349,N_5005,N_5020);
nand U5350 (N_5350,N_5108,N_5124);
and U5351 (N_5351,N_5014,N_5020);
nor U5352 (N_5352,N_5029,N_5141);
and U5353 (N_5353,N_5137,N_5036);
nor U5354 (N_5354,N_5040,N_5015);
nor U5355 (N_5355,N_5036,N_5165);
or U5356 (N_5356,N_5049,N_5036);
nor U5357 (N_5357,N_5176,N_5172);
nand U5358 (N_5358,N_5050,N_5162);
nor U5359 (N_5359,N_5123,N_5107);
nand U5360 (N_5360,N_5068,N_5067);
nor U5361 (N_5361,N_5166,N_5174);
xor U5362 (N_5362,N_5025,N_5000);
and U5363 (N_5363,N_5134,N_5012);
and U5364 (N_5364,N_5036,N_5077);
nand U5365 (N_5365,N_5167,N_5088);
nor U5366 (N_5366,N_5138,N_5035);
nor U5367 (N_5367,N_5059,N_5115);
or U5368 (N_5368,N_5117,N_5120);
nor U5369 (N_5369,N_5114,N_5131);
nor U5370 (N_5370,N_5073,N_5193);
and U5371 (N_5371,N_5083,N_5003);
and U5372 (N_5372,N_5133,N_5164);
nand U5373 (N_5373,N_5127,N_5146);
nand U5374 (N_5374,N_5024,N_5162);
nand U5375 (N_5375,N_5126,N_5193);
or U5376 (N_5376,N_5137,N_5144);
or U5377 (N_5377,N_5003,N_5054);
xnor U5378 (N_5378,N_5140,N_5191);
or U5379 (N_5379,N_5166,N_5193);
nor U5380 (N_5380,N_5159,N_5198);
xnor U5381 (N_5381,N_5119,N_5077);
nor U5382 (N_5382,N_5065,N_5162);
and U5383 (N_5383,N_5129,N_5005);
or U5384 (N_5384,N_5120,N_5064);
nor U5385 (N_5385,N_5050,N_5110);
nor U5386 (N_5386,N_5059,N_5069);
nor U5387 (N_5387,N_5065,N_5122);
or U5388 (N_5388,N_5039,N_5170);
and U5389 (N_5389,N_5022,N_5076);
and U5390 (N_5390,N_5190,N_5033);
xnor U5391 (N_5391,N_5069,N_5002);
nand U5392 (N_5392,N_5111,N_5087);
nand U5393 (N_5393,N_5148,N_5120);
nor U5394 (N_5394,N_5049,N_5135);
nor U5395 (N_5395,N_5189,N_5191);
nor U5396 (N_5396,N_5071,N_5087);
nand U5397 (N_5397,N_5106,N_5068);
nand U5398 (N_5398,N_5162,N_5082);
or U5399 (N_5399,N_5159,N_5197);
or U5400 (N_5400,N_5243,N_5274);
xor U5401 (N_5401,N_5270,N_5258);
or U5402 (N_5402,N_5298,N_5294);
and U5403 (N_5403,N_5305,N_5211);
and U5404 (N_5404,N_5226,N_5335);
or U5405 (N_5405,N_5350,N_5216);
and U5406 (N_5406,N_5221,N_5255);
nand U5407 (N_5407,N_5250,N_5222);
nand U5408 (N_5408,N_5267,N_5240);
nor U5409 (N_5409,N_5399,N_5382);
and U5410 (N_5410,N_5378,N_5287);
nand U5411 (N_5411,N_5374,N_5299);
nand U5412 (N_5412,N_5237,N_5276);
nor U5413 (N_5413,N_5202,N_5223);
nand U5414 (N_5414,N_5386,N_5387);
nand U5415 (N_5415,N_5277,N_5381);
and U5416 (N_5416,N_5310,N_5384);
nand U5417 (N_5417,N_5352,N_5213);
nand U5418 (N_5418,N_5329,N_5217);
xnor U5419 (N_5419,N_5224,N_5253);
xor U5420 (N_5420,N_5337,N_5201);
nor U5421 (N_5421,N_5319,N_5356);
nand U5422 (N_5422,N_5363,N_5364);
or U5423 (N_5423,N_5342,N_5260);
or U5424 (N_5424,N_5315,N_5295);
nor U5425 (N_5425,N_5355,N_5365);
nand U5426 (N_5426,N_5266,N_5314);
nor U5427 (N_5427,N_5333,N_5272);
nand U5428 (N_5428,N_5209,N_5293);
xor U5429 (N_5429,N_5351,N_5259);
nor U5430 (N_5430,N_5323,N_5245);
and U5431 (N_5431,N_5236,N_5206);
nor U5432 (N_5432,N_5361,N_5284);
and U5433 (N_5433,N_5300,N_5324);
xnor U5434 (N_5434,N_5358,N_5341);
nand U5435 (N_5435,N_5229,N_5385);
nor U5436 (N_5436,N_5207,N_5380);
nor U5437 (N_5437,N_5230,N_5247);
nand U5438 (N_5438,N_5311,N_5200);
and U5439 (N_5439,N_5330,N_5262);
nor U5440 (N_5440,N_5393,N_5347);
and U5441 (N_5441,N_5261,N_5228);
nor U5442 (N_5442,N_5291,N_5392);
nand U5443 (N_5443,N_5391,N_5215);
and U5444 (N_5444,N_5357,N_5322);
nor U5445 (N_5445,N_5268,N_5257);
and U5446 (N_5446,N_5340,N_5256);
nand U5447 (N_5447,N_5278,N_5346);
or U5448 (N_5448,N_5343,N_5344);
and U5449 (N_5449,N_5331,N_5264);
nor U5450 (N_5450,N_5366,N_5326);
nand U5451 (N_5451,N_5304,N_5210);
nor U5452 (N_5452,N_5377,N_5252);
xnor U5453 (N_5453,N_5204,N_5389);
xor U5454 (N_5454,N_5302,N_5368);
and U5455 (N_5455,N_5390,N_5325);
nand U5456 (N_5456,N_5388,N_5383);
nor U5457 (N_5457,N_5398,N_5376);
or U5458 (N_5458,N_5318,N_5312);
and U5459 (N_5459,N_5281,N_5327);
and U5460 (N_5460,N_5328,N_5233);
and U5461 (N_5461,N_5254,N_5301);
or U5462 (N_5462,N_5334,N_5395);
nand U5463 (N_5463,N_5321,N_5306);
nor U5464 (N_5464,N_5283,N_5289);
and U5465 (N_5465,N_5360,N_5338);
xnor U5466 (N_5466,N_5359,N_5227);
or U5467 (N_5467,N_5242,N_5394);
and U5468 (N_5468,N_5309,N_5203);
or U5469 (N_5469,N_5313,N_5280);
xor U5470 (N_5470,N_5219,N_5373);
xnor U5471 (N_5471,N_5225,N_5397);
nor U5472 (N_5472,N_5370,N_5308);
and U5473 (N_5473,N_5244,N_5212);
or U5474 (N_5474,N_5234,N_5263);
nand U5475 (N_5475,N_5275,N_5282);
and U5476 (N_5476,N_5371,N_5273);
or U5477 (N_5477,N_5214,N_5354);
and U5478 (N_5478,N_5290,N_5241);
nor U5479 (N_5479,N_5307,N_5265);
nand U5480 (N_5480,N_5396,N_5303);
or U5481 (N_5481,N_5251,N_5317);
nand U5482 (N_5482,N_5353,N_5372);
and U5483 (N_5483,N_5367,N_5362);
and U5484 (N_5484,N_5339,N_5279);
xor U5485 (N_5485,N_5246,N_5269);
nor U5486 (N_5486,N_5316,N_5286);
xnor U5487 (N_5487,N_5375,N_5379);
nand U5488 (N_5488,N_5349,N_5345);
or U5489 (N_5489,N_5232,N_5297);
and U5490 (N_5490,N_5332,N_5336);
xnor U5491 (N_5491,N_5288,N_5205);
and U5492 (N_5492,N_5239,N_5208);
nor U5493 (N_5493,N_5320,N_5348);
nand U5494 (N_5494,N_5249,N_5235);
and U5495 (N_5495,N_5369,N_5285);
xor U5496 (N_5496,N_5218,N_5238);
and U5497 (N_5497,N_5248,N_5271);
or U5498 (N_5498,N_5296,N_5220);
and U5499 (N_5499,N_5292,N_5231);
nor U5500 (N_5500,N_5306,N_5226);
nand U5501 (N_5501,N_5321,N_5262);
xor U5502 (N_5502,N_5356,N_5343);
and U5503 (N_5503,N_5386,N_5200);
or U5504 (N_5504,N_5330,N_5306);
nor U5505 (N_5505,N_5234,N_5397);
or U5506 (N_5506,N_5354,N_5288);
and U5507 (N_5507,N_5357,N_5371);
nor U5508 (N_5508,N_5227,N_5307);
xnor U5509 (N_5509,N_5390,N_5324);
or U5510 (N_5510,N_5384,N_5308);
nand U5511 (N_5511,N_5362,N_5265);
and U5512 (N_5512,N_5228,N_5219);
nor U5513 (N_5513,N_5266,N_5388);
xor U5514 (N_5514,N_5200,N_5337);
xnor U5515 (N_5515,N_5299,N_5326);
or U5516 (N_5516,N_5396,N_5366);
and U5517 (N_5517,N_5235,N_5204);
and U5518 (N_5518,N_5266,N_5343);
and U5519 (N_5519,N_5248,N_5294);
or U5520 (N_5520,N_5235,N_5371);
nor U5521 (N_5521,N_5242,N_5282);
nand U5522 (N_5522,N_5213,N_5225);
and U5523 (N_5523,N_5320,N_5316);
nand U5524 (N_5524,N_5321,N_5292);
or U5525 (N_5525,N_5287,N_5380);
nand U5526 (N_5526,N_5286,N_5337);
xor U5527 (N_5527,N_5317,N_5362);
and U5528 (N_5528,N_5388,N_5202);
and U5529 (N_5529,N_5226,N_5354);
and U5530 (N_5530,N_5325,N_5205);
or U5531 (N_5531,N_5371,N_5251);
and U5532 (N_5532,N_5322,N_5207);
or U5533 (N_5533,N_5212,N_5217);
xor U5534 (N_5534,N_5242,N_5349);
xnor U5535 (N_5535,N_5342,N_5377);
nand U5536 (N_5536,N_5298,N_5310);
nand U5537 (N_5537,N_5252,N_5201);
and U5538 (N_5538,N_5272,N_5399);
nand U5539 (N_5539,N_5301,N_5340);
and U5540 (N_5540,N_5257,N_5287);
and U5541 (N_5541,N_5213,N_5201);
nand U5542 (N_5542,N_5398,N_5332);
or U5543 (N_5543,N_5257,N_5225);
xnor U5544 (N_5544,N_5352,N_5251);
nor U5545 (N_5545,N_5304,N_5348);
xor U5546 (N_5546,N_5316,N_5344);
or U5547 (N_5547,N_5204,N_5287);
and U5548 (N_5548,N_5237,N_5339);
nor U5549 (N_5549,N_5230,N_5354);
nand U5550 (N_5550,N_5291,N_5372);
nor U5551 (N_5551,N_5391,N_5276);
and U5552 (N_5552,N_5220,N_5391);
or U5553 (N_5553,N_5379,N_5215);
and U5554 (N_5554,N_5324,N_5383);
nand U5555 (N_5555,N_5269,N_5241);
or U5556 (N_5556,N_5253,N_5316);
or U5557 (N_5557,N_5231,N_5384);
nand U5558 (N_5558,N_5238,N_5229);
nor U5559 (N_5559,N_5285,N_5238);
or U5560 (N_5560,N_5313,N_5231);
or U5561 (N_5561,N_5390,N_5308);
nand U5562 (N_5562,N_5250,N_5331);
xnor U5563 (N_5563,N_5302,N_5321);
nor U5564 (N_5564,N_5296,N_5233);
and U5565 (N_5565,N_5353,N_5304);
or U5566 (N_5566,N_5338,N_5370);
nand U5567 (N_5567,N_5384,N_5365);
xor U5568 (N_5568,N_5248,N_5225);
xnor U5569 (N_5569,N_5217,N_5396);
or U5570 (N_5570,N_5346,N_5259);
and U5571 (N_5571,N_5258,N_5376);
and U5572 (N_5572,N_5398,N_5212);
nand U5573 (N_5573,N_5382,N_5376);
and U5574 (N_5574,N_5263,N_5380);
and U5575 (N_5575,N_5310,N_5375);
nor U5576 (N_5576,N_5322,N_5365);
nor U5577 (N_5577,N_5324,N_5266);
or U5578 (N_5578,N_5222,N_5287);
nand U5579 (N_5579,N_5278,N_5331);
nand U5580 (N_5580,N_5225,N_5295);
or U5581 (N_5581,N_5284,N_5359);
nand U5582 (N_5582,N_5289,N_5216);
xor U5583 (N_5583,N_5359,N_5275);
or U5584 (N_5584,N_5398,N_5330);
xnor U5585 (N_5585,N_5269,N_5338);
nor U5586 (N_5586,N_5387,N_5354);
nand U5587 (N_5587,N_5214,N_5239);
nand U5588 (N_5588,N_5287,N_5250);
or U5589 (N_5589,N_5326,N_5388);
nor U5590 (N_5590,N_5292,N_5273);
nor U5591 (N_5591,N_5276,N_5308);
and U5592 (N_5592,N_5374,N_5202);
and U5593 (N_5593,N_5331,N_5299);
nor U5594 (N_5594,N_5229,N_5337);
nor U5595 (N_5595,N_5377,N_5261);
nand U5596 (N_5596,N_5234,N_5297);
or U5597 (N_5597,N_5349,N_5201);
or U5598 (N_5598,N_5361,N_5233);
and U5599 (N_5599,N_5260,N_5205);
and U5600 (N_5600,N_5501,N_5548);
nor U5601 (N_5601,N_5414,N_5456);
nand U5602 (N_5602,N_5515,N_5571);
nor U5603 (N_5603,N_5539,N_5541);
nor U5604 (N_5604,N_5527,N_5584);
nand U5605 (N_5605,N_5459,N_5556);
nor U5606 (N_5606,N_5519,N_5410);
nor U5607 (N_5607,N_5416,N_5413);
nor U5608 (N_5608,N_5421,N_5437);
or U5609 (N_5609,N_5407,N_5589);
and U5610 (N_5610,N_5559,N_5511);
nor U5611 (N_5611,N_5528,N_5512);
nor U5612 (N_5612,N_5406,N_5534);
nand U5613 (N_5613,N_5491,N_5498);
nor U5614 (N_5614,N_5466,N_5412);
nand U5615 (N_5615,N_5468,N_5486);
xor U5616 (N_5616,N_5572,N_5428);
nor U5617 (N_5617,N_5477,N_5596);
nor U5618 (N_5618,N_5505,N_5440);
nor U5619 (N_5619,N_5580,N_5582);
or U5620 (N_5620,N_5472,N_5591);
or U5621 (N_5621,N_5524,N_5436);
nand U5622 (N_5622,N_5403,N_5509);
nand U5623 (N_5623,N_5445,N_5508);
or U5624 (N_5624,N_5467,N_5404);
nor U5625 (N_5625,N_5418,N_5574);
nor U5626 (N_5626,N_5479,N_5578);
nand U5627 (N_5627,N_5441,N_5409);
and U5628 (N_5628,N_5438,N_5550);
or U5629 (N_5629,N_5518,N_5564);
or U5630 (N_5630,N_5478,N_5442);
nor U5631 (N_5631,N_5450,N_5411);
and U5632 (N_5632,N_5551,N_5533);
and U5633 (N_5633,N_5431,N_5536);
nand U5634 (N_5634,N_5542,N_5405);
or U5635 (N_5635,N_5487,N_5457);
or U5636 (N_5636,N_5588,N_5415);
and U5637 (N_5637,N_5446,N_5422);
nor U5638 (N_5638,N_5439,N_5543);
or U5639 (N_5639,N_5530,N_5433);
nand U5640 (N_5640,N_5461,N_5483);
nand U5641 (N_5641,N_5547,N_5400);
nand U5642 (N_5642,N_5570,N_5401);
and U5643 (N_5643,N_5417,N_5540);
nor U5644 (N_5644,N_5451,N_5531);
nand U5645 (N_5645,N_5581,N_5492);
or U5646 (N_5646,N_5599,N_5482);
nand U5647 (N_5647,N_5434,N_5430);
nand U5648 (N_5648,N_5544,N_5555);
nor U5649 (N_5649,N_5453,N_5480);
nand U5650 (N_5650,N_5552,N_5473);
xnor U5651 (N_5651,N_5429,N_5598);
nand U5652 (N_5652,N_5426,N_5546);
or U5653 (N_5653,N_5488,N_5537);
or U5654 (N_5654,N_5549,N_5579);
or U5655 (N_5655,N_5503,N_5490);
nor U5656 (N_5656,N_5448,N_5471);
xor U5657 (N_5657,N_5454,N_5424);
or U5658 (N_5658,N_5447,N_5408);
nor U5659 (N_5659,N_5567,N_5566);
nand U5660 (N_5660,N_5554,N_5425);
and U5661 (N_5661,N_5464,N_5526);
nor U5662 (N_5662,N_5583,N_5517);
or U5663 (N_5663,N_5558,N_5523);
nor U5664 (N_5664,N_5587,N_5506);
and U5665 (N_5665,N_5402,N_5520);
and U5666 (N_5666,N_5435,N_5484);
nand U5667 (N_5667,N_5463,N_5458);
xnor U5668 (N_5668,N_5476,N_5452);
xnor U5669 (N_5669,N_5474,N_5427);
and U5670 (N_5670,N_5593,N_5475);
or U5671 (N_5671,N_5590,N_5432);
nor U5672 (N_5672,N_5569,N_5455);
nand U5673 (N_5673,N_5470,N_5504);
and U5674 (N_5674,N_5493,N_5576);
xnor U5675 (N_5675,N_5465,N_5513);
nand U5676 (N_5676,N_5420,N_5419);
or U5677 (N_5677,N_5565,N_5495);
xnor U5678 (N_5678,N_5557,N_5423);
or U5679 (N_5679,N_5499,N_5525);
nand U5680 (N_5680,N_5500,N_5443);
nand U5681 (N_5681,N_5562,N_5577);
and U5682 (N_5682,N_5597,N_5497);
nand U5683 (N_5683,N_5516,N_5585);
or U5684 (N_5684,N_5545,N_5573);
or U5685 (N_5685,N_5460,N_5462);
nor U5686 (N_5686,N_5592,N_5469);
nor U5687 (N_5687,N_5535,N_5514);
nor U5688 (N_5688,N_5521,N_5563);
and U5689 (N_5689,N_5538,N_5586);
or U5690 (N_5690,N_5502,N_5522);
nor U5691 (N_5691,N_5553,N_5560);
and U5692 (N_5692,N_5568,N_5444);
or U5693 (N_5693,N_5575,N_5532);
and U5694 (N_5694,N_5489,N_5594);
and U5695 (N_5695,N_5494,N_5496);
and U5696 (N_5696,N_5481,N_5510);
nand U5697 (N_5697,N_5485,N_5595);
or U5698 (N_5698,N_5449,N_5529);
nand U5699 (N_5699,N_5561,N_5507);
nand U5700 (N_5700,N_5454,N_5419);
and U5701 (N_5701,N_5580,N_5489);
or U5702 (N_5702,N_5444,N_5421);
xnor U5703 (N_5703,N_5563,N_5443);
nand U5704 (N_5704,N_5473,N_5474);
xnor U5705 (N_5705,N_5520,N_5511);
or U5706 (N_5706,N_5546,N_5478);
nor U5707 (N_5707,N_5509,N_5449);
or U5708 (N_5708,N_5475,N_5401);
nor U5709 (N_5709,N_5497,N_5463);
nand U5710 (N_5710,N_5454,N_5430);
or U5711 (N_5711,N_5456,N_5574);
nand U5712 (N_5712,N_5481,N_5406);
xnor U5713 (N_5713,N_5446,N_5449);
or U5714 (N_5714,N_5472,N_5504);
nand U5715 (N_5715,N_5450,N_5437);
xor U5716 (N_5716,N_5528,N_5595);
nand U5717 (N_5717,N_5574,N_5445);
xnor U5718 (N_5718,N_5489,N_5554);
or U5719 (N_5719,N_5452,N_5527);
or U5720 (N_5720,N_5538,N_5510);
nor U5721 (N_5721,N_5433,N_5554);
nor U5722 (N_5722,N_5500,N_5594);
nor U5723 (N_5723,N_5505,N_5447);
and U5724 (N_5724,N_5430,N_5554);
or U5725 (N_5725,N_5541,N_5455);
and U5726 (N_5726,N_5594,N_5436);
xor U5727 (N_5727,N_5410,N_5508);
nand U5728 (N_5728,N_5598,N_5420);
and U5729 (N_5729,N_5566,N_5479);
nand U5730 (N_5730,N_5504,N_5466);
nand U5731 (N_5731,N_5523,N_5525);
nor U5732 (N_5732,N_5556,N_5525);
nand U5733 (N_5733,N_5588,N_5523);
nand U5734 (N_5734,N_5511,N_5594);
nor U5735 (N_5735,N_5427,N_5477);
and U5736 (N_5736,N_5461,N_5543);
nor U5737 (N_5737,N_5415,N_5519);
nor U5738 (N_5738,N_5410,N_5404);
and U5739 (N_5739,N_5459,N_5521);
nor U5740 (N_5740,N_5490,N_5579);
nand U5741 (N_5741,N_5428,N_5593);
nor U5742 (N_5742,N_5549,N_5574);
and U5743 (N_5743,N_5466,N_5445);
and U5744 (N_5744,N_5538,N_5528);
xor U5745 (N_5745,N_5577,N_5451);
or U5746 (N_5746,N_5490,N_5433);
and U5747 (N_5747,N_5549,N_5450);
or U5748 (N_5748,N_5575,N_5580);
nand U5749 (N_5749,N_5553,N_5479);
or U5750 (N_5750,N_5536,N_5442);
nor U5751 (N_5751,N_5447,N_5424);
and U5752 (N_5752,N_5491,N_5597);
xor U5753 (N_5753,N_5586,N_5414);
or U5754 (N_5754,N_5534,N_5590);
nor U5755 (N_5755,N_5487,N_5456);
xnor U5756 (N_5756,N_5431,N_5541);
nand U5757 (N_5757,N_5540,N_5442);
nor U5758 (N_5758,N_5443,N_5509);
nor U5759 (N_5759,N_5507,N_5483);
xnor U5760 (N_5760,N_5463,N_5591);
xnor U5761 (N_5761,N_5572,N_5473);
xor U5762 (N_5762,N_5549,N_5529);
or U5763 (N_5763,N_5589,N_5480);
nand U5764 (N_5764,N_5500,N_5412);
nor U5765 (N_5765,N_5484,N_5555);
nand U5766 (N_5766,N_5591,N_5427);
nor U5767 (N_5767,N_5418,N_5569);
nand U5768 (N_5768,N_5420,N_5518);
nor U5769 (N_5769,N_5580,N_5532);
nor U5770 (N_5770,N_5572,N_5490);
nand U5771 (N_5771,N_5411,N_5440);
nand U5772 (N_5772,N_5478,N_5576);
nand U5773 (N_5773,N_5484,N_5455);
and U5774 (N_5774,N_5417,N_5558);
and U5775 (N_5775,N_5402,N_5509);
and U5776 (N_5776,N_5446,N_5436);
or U5777 (N_5777,N_5449,N_5575);
xor U5778 (N_5778,N_5437,N_5513);
nand U5779 (N_5779,N_5499,N_5408);
nor U5780 (N_5780,N_5522,N_5458);
nand U5781 (N_5781,N_5516,N_5471);
nor U5782 (N_5782,N_5527,N_5546);
xor U5783 (N_5783,N_5567,N_5529);
and U5784 (N_5784,N_5566,N_5578);
nor U5785 (N_5785,N_5590,N_5541);
nor U5786 (N_5786,N_5512,N_5424);
and U5787 (N_5787,N_5447,N_5573);
xor U5788 (N_5788,N_5464,N_5595);
and U5789 (N_5789,N_5470,N_5532);
nor U5790 (N_5790,N_5549,N_5531);
nor U5791 (N_5791,N_5517,N_5537);
nand U5792 (N_5792,N_5479,N_5546);
nand U5793 (N_5793,N_5580,N_5419);
or U5794 (N_5794,N_5589,N_5416);
nand U5795 (N_5795,N_5540,N_5425);
xor U5796 (N_5796,N_5505,N_5595);
nor U5797 (N_5797,N_5509,N_5429);
and U5798 (N_5798,N_5468,N_5466);
nand U5799 (N_5799,N_5591,N_5456);
and U5800 (N_5800,N_5735,N_5788);
xor U5801 (N_5801,N_5652,N_5754);
nand U5802 (N_5802,N_5752,N_5799);
and U5803 (N_5803,N_5703,N_5672);
nand U5804 (N_5804,N_5781,N_5667);
nor U5805 (N_5805,N_5604,N_5603);
and U5806 (N_5806,N_5660,N_5640);
nand U5807 (N_5807,N_5771,N_5748);
nand U5808 (N_5808,N_5773,N_5779);
nand U5809 (N_5809,N_5689,N_5627);
or U5810 (N_5810,N_5705,N_5649);
nor U5811 (N_5811,N_5796,N_5696);
or U5812 (N_5812,N_5683,N_5634);
nand U5813 (N_5813,N_5723,N_5795);
or U5814 (N_5814,N_5717,N_5756);
or U5815 (N_5815,N_5636,N_5739);
nand U5816 (N_5816,N_5670,N_5777);
or U5817 (N_5817,N_5747,N_5616);
or U5818 (N_5818,N_5642,N_5663);
nor U5819 (N_5819,N_5624,N_5704);
or U5820 (N_5820,N_5721,N_5630);
or U5821 (N_5821,N_5785,N_5661);
and U5822 (N_5822,N_5633,N_5715);
and U5823 (N_5823,N_5784,N_5653);
nor U5824 (N_5824,N_5780,N_5726);
and U5825 (N_5825,N_5629,N_5716);
xor U5826 (N_5826,N_5608,N_5639);
nor U5827 (N_5827,N_5632,N_5625);
and U5828 (N_5828,N_5798,N_5607);
and U5829 (N_5829,N_5774,N_5646);
and U5830 (N_5830,N_5789,N_5681);
and U5831 (N_5831,N_5678,N_5623);
nand U5832 (N_5832,N_5645,N_5601);
and U5833 (N_5833,N_5791,N_5644);
or U5834 (N_5834,N_5764,N_5686);
and U5835 (N_5835,N_5635,N_5677);
xor U5836 (N_5836,N_5734,N_5758);
and U5837 (N_5837,N_5658,N_5767);
nand U5838 (N_5838,N_5622,N_5743);
and U5839 (N_5839,N_5745,N_5665);
nand U5840 (N_5840,N_5759,N_5637);
or U5841 (N_5841,N_5769,N_5790);
and U5842 (N_5842,N_5760,N_5643);
nand U5843 (N_5843,N_5617,N_5657);
nand U5844 (N_5844,N_5669,N_5620);
nor U5845 (N_5845,N_5659,N_5738);
and U5846 (N_5846,N_5714,N_5631);
nand U5847 (N_5847,N_5770,N_5782);
and U5848 (N_5848,N_5776,N_5668);
and U5849 (N_5849,N_5761,N_5641);
or U5850 (N_5850,N_5730,N_5638);
xnor U5851 (N_5851,N_5797,N_5648);
and U5852 (N_5852,N_5722,N_5609);
and U5853 (N_5853,N_5732,N_5755);
nand U5854 (N_5854,N_5753,N_5697);
nand U5855 (N_5855,N_5712,N_5619);
and U5856 (N_5856,N_5676,N_5706);
and U5857 (N_5857,N_5731,N_5729);
or U5858 (N_5858,N_5662,N_5765);
and U5859 (N_5859,N_5615,N_5700);
and U5860 (N_5860,N_5741,N_5713);
xor U5861 (N_5861,N_5693,N_5724);
or U5862 (N_5862,N_5702,N_5736);
nor U5863 (N_5863,N_5763,N_5610);
nand U5864 (N_5864,N_5684,N_5611);
or U5865 (N_5865,N_5679,N_5709);
nand U5866 (N_5866,N_5650,N_5671);
nand U5867 (N_5867,N_5666,N_5710);
nand U5868 (N_5868,N_5778,N_5602);
or U5869 (N_5869,N_5673,N_5751);
or U5870 (N_5870,N_5691,N_5606);
or U5871 (N_5871,N_5651,N_5699);
nor U5872 (N_5872,N_5727,N_5694);
or U5873 (N_5873,N_5656,N_5718);
nor U5874 (N_5874,N_5737,N_5746);
nor U5875 (N_5875,N_5744,N_5628);
or U5876 (N_5876,N_5626,N_5618);
xor U5877 (N_5877,N_5701,N_5768);
nand U5878 (N_5878,N_5707,N_5742);
nor U5879 (N_5879,N_5621,N_5687);
nand U5880 (N_5880,N_5708,N_5613);
or U5881 (N_5881,N_5698,N_5775);
nand U5882 (N_5882,N_5690,N_5612);
xnor U5883 (N_5883,N_5740,N_5605);
nor U5884 (N_5884,N_5793,N_5762);
or U5885 (N_5885,N_5725,N_5786);
nand U5886 (N_5886,N_5647,N_5682);
nand U5887 (N_5887,N_5749,N_5600);
or U5888 (N_5888,N_5685,N_5794);
or U5889 (N_5889,N_5792,N_5720);
nand U5890 (N_5890,N_5711,N_5675);
nor U5891 (N_5891,N_5654,N_5783);
nor U5892 (N_5892,N_5695,N_5688);
nand U5893 (N_5893,N_5766,N_5719);
nor U5894 (N_5894,N_5728,N_5664);
or U5895 (N_5895,N_5655,N_5680);
nor U5896 (N_5896,N_5733,N_5757);
or U5897 (N_5897,N_5787,N_5750);
nor U5898 (N_5898,N_5614,N_5692);
and U5899 (N_5899,N_5772,N_5674);
xor U5900 (N_5900,N_5679,N_5604);
nor U5901 (N_5901,N_5635,N_5769);
and U5902 (N_5902,N_5604,N_5711);
or U5903 (N_5903,N_5769,N_5699);
and U5904 (N_5904,N_5695,N_5795);
nand U5905 (N_5905,N_5790,N_5674);
nand U5906 (N_5906,N_5677,N_5755);
nand U5907 (N_5907,N_5770,N_5660);
nand U5908 (N_5908,N_5789,N_5675);
nand U5909 (N_5909,N_5621,N_5628);
or U5910 (N_5910,N_5773,N_5669);
and U5911 (N_5911,N_5689,N_5740);
nor U5912 (N_5912,N_5662,N_5793);
or U5913 (N_5913,N_5733,N_5604);
nor U5914 (N_5914,N_5714,N_5747);
and U5915 (N_5915,N_5687,N_5661);
and U5916 (N_5916,N_5699,N_5788);
and U5917 (N_5917,N_5690,N_5770);
nand U5918 (N_5918,N_5739,N_5780);
nor U5919 (N_5919,N_5713,N_5682);
nor U5920 (N_5920,N_5740,N_5719);
xor U5921 (N_5921,N_5778,N_5695);
or U5922 (N_5922,N_5780,N_5644);
nor U5923 (N_5923,N_5708,N_5713);
and U5924 (N_5924,N_5637,N_5795);
or U5925 (N_5925,N_5671,N_5700);
or U5926 (N_5926,N_5771,N_5676);
nor U5927 (N_5927,N_5602,N_5727);
nand U5928 (N_5928,N_5630,N_5760);
nor U5929 (N_5929,N_5705,N_5713);
or U5930 (N_5930,N_5751,N_5771);
nor U5931 (N_5931,N_5758,N_5668);
or U5932 (N_5932,N_5734,N_5683);
or U5933 (N_5933,N_5780,N_5686);
nor U5934 (N_5934,N_5672,N_5766);
nand U5935 (N_5935,N_5784,N_5709);
and U5936 (N_5936,N_5725,N_5633);
or U5937 (N_5937,N_5730,N_5712);
xnor U5938 (N_5938,N_5727,N_5774);
or U5939 (N_5939,N_5728,N_5639);
or U5940 (N_5940,N_5705,N_5765);
and U5941 (N_5941,N_5626,N_5728);
or U5942 (N_5942,N_5641,N_5654);
nor U5943 (N_5943,N_5784,N_5762);
and U5944 (N_5944,N_5699,N_5691);
and U5945 (N_5945,N_5722,N_5675);
nor U5946 (N_5946,N_5773,N_5770);
nand U5947 (N_5947,N_5697,N_5746);
nand U5948 (N_5948,N_5677,N_5604);
or U5949 (N_5949,N_5671,N_5751);
nor U5950 (N_5950,N_5753,N_5649);
nand U5951 (N_5951,N_5728,N_5652);
xor U5952 (N_5952,N_5717,N_5615);
or U5953 (N_5953,N_5677,N_5664);
and U5954 (N_5954,N_5604,N_5789);
and U5955 (N_5955,N_5612,N_5660);
nor U5956 (N_5956,N_5687,N_5770);
or U5957 (N_5957,N_5618,N_5724);
nor U5958 (N_5958,N_5647,N_5796);
nor U5959 (N_5959,N_5749,N_5735);
or U5960 (N_5960,N_5686,N_5738);
nor U5961 (N_5961,N_5712,N_5682);
nor U5962 (N_5962,N_5765,N_5699);
and U5963 (N_5963,N_5768,N_5697);
nor U5964 (N_5964,N_5742,N_5658);
nor U5965 (N_5965,N_5646,N_5672);
nor U5966 (N_5966,N_5789,N_5704);
and U5967 (N_5967,N_5663,N_5636);
or U5968 (N_5968,N_5614,N_5606);
and U5969 (N_5969,N_5676,N_5674);
or U5970 (N_5970,N_5604,N_5619);
nor U5971 (N_5971,N_5615,N_5626);
and U5972 (N_5972,N_5631,N_5602);
nor U5973 (N_5973,N_5781,N_5727);
nor U5974 (N_5974,N_5657,N_5631);
nor U5975 (N_5975,N_5643,N_5757);
and U5976 (N_5976,N_5675,N_5733);
and U5977 (N_5977,N_5787,N_5666);
nor U5978 (N_5978,N_5684,N_5709);
and U5979 (N_5979,N_5799,N_5688);
nand U5980 (N_5980,N_5673,N_5726);
and U5981 (N_5981,N_5738,N_5732);
nand U5982 (N_5982,N_5661,N_5739);
nand U5983 (N_5983,N_5689,N_5785);
nand U5984 (N_5984,N_5744,N_5728);
nor U5985 (N_5985,N_5754,N_5629);
or U5986 (N_5986,N_5605,N_5792);
and U5987 (N_5987,N_5730,N_5603);
nor U5988 (N_5988,N_5664,N_5791);
nor U5989 (N_5989,N_5709,N_5761);
and U5990 (N_5990,N_5764,N_5782);
nor U5991 (N_5991,N_5624,N_5674);
nor U5992 (N_5992,N_5746,N_5618);
and U5993 (N_5993,N_5676,N_5736);
nand U5994 (N_5994,N_5625,N_5659);
or U5995 (N_5995,N_5733,N_5735);
and U5996 (N_5996,N_5602,N_5609);
nand U5997 (N_5997,N_5713,N_5731);
nor U5998 (N_5998,N_5627,N_5697);
and U5999 (N_5999,N_5686,N_5633);
xor U6000 (N_6000,N_5841,N_5892);
and U6001 (N_6001,N_5809,N_5969);
nand U6002 (N_6002,N_5940,N_5998);
nand U6003 (N_6003,N_5949,N_5850);
nand U6004 (N_6004,N_5803,N_5980);
nor U6005 (N_6005,N_5877,N_5893);
and U6006 (N_6006,N_5905,N_5963);
or U6007 (N_6007,N_5900,N_5874);
and U6008 (N_6008,N_5887,N_5921);
nand U6009 (N_6009,N_5978,N_5835);
nor U6010 (N_6010,N_5907,N_5943);
nand U6011 (N_6011,N_5848,N_5955);
and U6012 (N_6012,N_5976,N_5995);
xor U6013 (N_6013,N_5936,N_5912);
and U6014 (N_6014,N_5983,N_5933);
nand U6015 (N_6015,N_5960,N_5984);
and U6016 (N_6016,N_5961,N_5831);
nor U6017 (N_6017,N_5934,N_5979);
xor U6018 (N_6018,N_5842,N_5922);
xnor U6019 (N_6019,N_5811,N_5950);
or U6020 (N_6020,N_5975,N_5826);
or U6021 (N_6021,N_5879,N_5832);
or U6022 (N_6022,N_5991,N_5968);
nand U6023 (N_6023,N_5947,N_5918);
nor U6024 (N_6024,N_5930,N_5830);
and U6025 (N_6025,N_5856,N_5913);
nand U6026 (N_6026,N_5958,N_5816);
nor U6027 (N_6027,N_5972,N_5990);
nand U6028 (N_6028,N_5822,N_5992);
or U6029 (N_6029,N_5906,N_5876);
xnor U6030 (N_6030,N_5970,N_5878);
and U6031 (N_6031,N_5813,N_5847);
and U6032 (N_6032,N_5891,N_5890);
and U6033 (N_6033,N_5820,N_5895);
nand U6034 (N_6034,N_5896,N_5852);
nand U6035 (N_6035,N_5897,N_5810);
and U6036 (N_6036,N_5806,N_5966);
or U6037 (N_6037,N_5805,N_5914);
or U6038 (N_6038,N_5932,N_5957);
nor U6039 (N_6039,N_5861,N_5928);
nand U6040 (N_6040,N_5911,N_5908);
and U6041 (N_6041,N_5935,N_5868);
or U6042 (N_6042,N_5821,N_5920);
nor U6043 (N_6043,N_5817,N_5903);
and U6044 (N_6044,N_5828,N_5871);
nand U6045 (N_6045,N_5882,N_5825);
and U6046 (N_6046,N_5977,N_5858);
nand U6047 (N_6047,N_5942,N_5941);
nor U6048 (N_6048,N_5834,N_5946);
nor U6049 (N_6049,N_5938,N_5862);
nand U6050 (N_6050,N_5989,N_5939);
nor U6051 (N_6051,N_5829,N_5974);
and U6052 (N_6052,N_5999,N_5899);
nand U6053 (N_6053,N_5881,N_5837);
nor U6054 (N_6054,N_5857,N_5833);
nand U6055 (N_6055,N_5927,N_5915);
nand U6056 (N_6056,N_5802,N_5937);
and U6057 (N_6057,N_5888,N_5853);
nor U6058 (N_6058,N_5843,N_5849);
nor U6059 (N_6059,N_5844,N_5889);
nor U6060 (N_6060,N_5959,N_5859);
nand U6061 (N_6061,N_5909,N_5931);
and U6062 (N_6062,N_5839,N_5872);
or U6063 (N_6063,N_5902,N_5836);
xor U6064 (N_6064,N_5886,N_5807);
or U6065 (N_6065,N_5867,N_5883);
nor U6066 (N_6066,N_5840,N_5910);
nor U6067 (N_6067,N_5917,N_5824);
nand U6068 (N_6068,N_5964,N_5814);
nand U6069 (N_6069,N_5956,N_5827);
nor U6070 (N_6070,N_5925,N_5924);
and U6071 (N_6071,N_5919,N_5894);
and U6072 (N_6072,N_5885,N_5866);
xor U6073 (N_6073,N_5846,N_5948);
nor U6074 (N_6074,N_5962,N_5863);
xnor U6075 (N_6075,N_5996,N_5845);
nand U6076 (N_6076,N_5997,N_5873);
and U6077 (N_6077,N_5981,N_5804);
or U6078 (N_6078,N_5954,N_5994);
xor U6079 (N_6079,N_5982,N_5951);
and U6080 (N_6080,N_5965,N_5986);
and U6081 (N_6081,N_5812,N_5971);
nor U6082 (N_6082,N_5985,N_5869);
nand U6083 (N_6083,N_5860,N_5884);
nor U6084 (N_6084,N_5923,N_5875);
nand U6085 (N_6085,N_5864,N_5800);
nand U6086 (N_6086,N_5987,N_5808);
or U6087 (N_6087,N_5953,N_5898);
and U6088 (N_6088,N_5993,N_5944);
xnor U6089 (N_6089,N_5855,N_5865);
nand U6090 (N_6090,N_5926,N_5818);
and U6091 (N_6091,N_5945,N_5952);
nand U6092 (N_6092,N_5929,N_5870);
nand U6093 (N_6093,N_5967,N_5988);
or U6094 (N_6094,N_5904,N_5880);
nand U6095 (N_6095,N_5801,N_5854);
xor U6096 (N_6096,N_5815,N_5819);
xnor U6097 (N_6097,N_5823,N_5838);
and U6098 (N_6098,N_5973,N_5851);
nor U6099 (N_6099,N_5916,N_5901);
nand U6100 (N_6100,N_5987,N_5803);
or U6101 (N_6101,N_5847,N_5922);
or U6102 (N_6102,N_5931,N_5906);
or U6103 (N_6103,N_5998,N_5955);
xnor U6104 (N_6104,N_5843,N_5974);
and U6105 (N_6105,N_5954,N_5813);
or U6106 (N_6106,N_5829,N_5943);
xnor U6107 (N_6107,N_5929,N_5957);
and U6108 (N_6108,N_5937,N_5825);
xnor U6109 (N_6109,N_5835,N_5919);
or U6110 (N_6110,N_5936,N_5856);
and U6111 (N_6111,N_5938,N_5883);
nor U6112 (N_6112,N_5909,N_5884);
nand U6113 (N_6113,N_5875,N_5990);
or U6114 (N_6114,N_5958,N_5933);
nor U6115 (N_6115,N_5981,N_5900);
nand U6116 (N_6116,N_5882,N_5807);
or U6117 (N_6117,N_5913,N_5930);
and U6118 (N_6118,N_5970,N_5831);
nor U6119 (N_6119,N_5849,N_5930);
nand U6120 (N_6120,N_5968,N_5800);
nor U6121 (N_6121,N_5919,N_5883);
xnor U6122 (N_6122,N_5982,N_5977);
nand U6123 (N_6123,N_5935,N_5865);
nor U6124 (N_6124,N_5967,N_5800);
nor U6125 (N_6125,N_5821,N_5892);
nor U6126 (N_6126,N_5868,N_5878);
or U6127 (N_6127,N_5801,N_5828);
nor U6128 (N_6128,N_5896,N_5940);
nand U6129 (N_6129,N_5880,N_5811);
or U6130 (N_6130,N_5804,N_5951);
nand U6131 (N_6131,N_5951,N_5996);
and U6132 (N_6132,N_5945,N_5980);
nand U6133 (N_6133,N_5867,N_5888);
xor U6134 (N_6134,N_5952,N_5957);
and U6135 (N_6135,N_5849,N_5863);
and U6136 (N_6136,N_5846,N_5981);
nor U6137 (N_6137,N_5869,N_5970);
nand U6138 (N_6138,N_5879,N_5913);
or U6139 (N_6139,N_5946,N_5816);
nand U6140 (N_6140,N_5973,N_5823);
nand U6141 (N_6141,N_5893,N_5947);
and U6142 (N_6142,N_5840,N_5800);
nand U6143 (N_6143,N_5971,N_5937);
nor U6144 (N_6144,N_5960,N_5952);
nand U6145 (N_6145,N_5999,N_5918);
nor U6146 (N_6146,N_5821,N_5876);
and U6147 (N_6147,N_5893,N_5895);
nand U6148 (N_6148,N_5904,N_5823);
nor U6149 (N_6149,N_5922,N_5919);
and U6150 (N_6150,N_5972,N_5998);
nand U6151 (N_6151,N_5914,N_5892);
or U6152 (N_6152,N_5874,N_5933);
nand U6153 (N_6153,N_5984,N_5900);
or U6154 (N_6154,N_5918,N_5870);
nor U6155 (N_6155,N_5905,N_5860);
or U6156 (N_6156,N_5987,N_5831);
nand U6157 (N_6157,N_5862,N_5886);
and U6158 (N_6158,N_5932,N_5982);
nand U6159 (N_6159,N_5994,N_5987);
xnor U6160 (N_6160,N_5936,N_5922);
and U6161 (N_6161,N_5884,N_5991);
and U6162 (N_6162,N_5834,N_5979);
or U6163 (N_6163,N_5941,N_5905);
nand U6164 (N_6164,N_5902,N_5883);
nor U6165 (N_6165,N_5874,N_5899);
nor U6166 (N_6166,N_5965,N_5817);
or U6167 (N_6167,N_5855,N_5928);
nor U6168 (N_6168,N_5871,N_5835);
or U6169 (N_6169,N_5903,N_5845);
or U6170 (N_6170,N_5980,N_5860);
or U6171 (N_6171,N_5853,N_5845);
or U6172 (N_6172,N_5823,N_5808);
nor U6173 (N_6173,N_5875,N_5945);
and U6174 (N_6174,N_5814,N_5816);
nor U6175 (N_6175,N_5865,N_5873);
nor U6176 (N_6176,N_5994,N_5809);
or U6177 (N_6177,N_5979,N_5919);
nor U6178 (N_6178,N_5849,N_5888);
nand U6179 (N_6179,N_5924,N_5812);
nand U6180 (N_6180,N_5875,N_5978);
xnor U6181 (N_6181,N_5843,N_5932);
nand U6182 (N_6182,N_5885,N_5925);
and U6183 (N_6183,N_5814,N_5972);
nand U6184 (N_6184,N_5803,N_5861);
or U6185 (N_6185,N_5887,N_5977);
and U6186 (N_6186,N_5949,N_5950);
or U6187 (N_6187,N_5944,N_5860);
and U6188 (N_6188,N_5836,N_5974);
xor U6189 (N_6189,N_5935,N_5820);
and U6190 (N_6190,N_5859,N_5908);
nand U6191 (N_6191,N_5874,N_5905);
or U6192 (N_6192,N_5906,N_5835);
or U6193 (N_6193,N_5915,N_5866);
or U6194 (N_6194,N_5972,N_5975);
and U6195 (N_6195,N_5815,N_5996);
nor U6196 (N_6196,N_5944,N_5919);
and U6197 (N_6197,N_5989,N_5971);
nand U6198 (N_6198,N_5949,N_5975);
nor U6199 (N_6199,N_5820,N_5864);
xor U6200 (N_6200,N_6118,N_6186);
and U6201 (N_6201,N_6166,N_6062);
nor U6202 (N_6202,N_6057,N_6059);
and U6203 (N_6203,N_6172,N_6018);
or U6204 (N_6204,N_6171,N_6194);
nand U6205 (N_6205,N_6000,N_6162);
and U6206 (N_6206,N_6135,N_6070);
nor U6207 (N_6207,N_6167,N_6098);
or U6208 (N_6208,N_6155,N_6144);
or U6209 (N_6209,N_6159,N_6093);
and U6210 (N_6210,N_6082,N_6060);
nand U6211 (N_6211,N_6084,N_6045);
or U6212 (N_6212,N_6113,N_6073);
or U6213 (N_6213,N_6077,N_6019);
and U6214 (N_6214,N_6078,N_6177);
nand U6215 (N_6215,N_6139,N_6039);
and U6216 (N_6216,N_6013,N_6153);
and U6217 (N_6217,N_6140,N_6001);
and U6218 (N_6218,N_6033,N_6106);
nand U6219 (N_6219,N_6141,N_6188);
xor U6220 (N_6220,N_6023,N_6131);
nand U6221 (N_6221,N_6164,N_6046);
nor U6222 (N_6222,N_6008,N_6165);
nor U6223 (N_6223,N_6168,N_6096);
xor U6224 (N_6224,N_6092,N_6130);
and U6225 (N_6225,N_6121,N_6069);
nor U6226 (N_6226,N_6192,N_6199);
xor U6227 (N_6227,N_6031,N_6072);
nand U6228 (N_6228,N_6015,N_6197);
or U6229 (N_6229,N_6095,N_6119);
nand U6230 (N_6230,N_6079,N_6161);
or U6231 (N_6231,N_6043,N_6040);
and U6232 (N_6232,N_6006,N_6016);
and U6233 (N_6233,N_6169,N_6117);
and U6234 (N_6234,N_6116,N_6002);
xnor U6235 (N_6235,N_6150,N_6103);
or U6236 (N_6236,N_6076,N_6053);
nor U6237 (N_6237,N_6085,N_6120);
nor U6238 (N_6238,N_6124,N_6099);
and U6239 (N_6239,N_6065,N_6128);
and U6240 (N_6240,N_6028,N_6145);
nand U6241 (N_6241,N_6003,N_6133);
or U6242 (N_6242,N_6127,N_6012);
nand U6243 (N_6243,N_6071,N_6142);
xor U6244 (N_6244,N_6190,N_6149);
nand U6245 (N_6245,N_6104,N_6022);
and U6246 (N_6246,N_6129,N_6112);
xor U6247 (N_6247,N_6173,N_6042);
or U6248 (N_6248,N_6151,N_6058);
nand U6249 (N_6249,N_6152,N_6146);
or U6250 (N_6250,N_6089,N_6067);
and U6251 (N_6251,N_6086,N_6163);
nor U6252 (N_6252,N_6183,N_6061);
nor U6253 (N_6253,N_6035,N_6179);
nand U6254 (N_6254,N_6102,N_6195);
xnor U6255 (N_6255,N_6185,N_6111);
or U6256 (N_6256,N_6105,N_6100);
and U6257 (N_6257,N_6122,N_6068);
nor U6258 (N_6258,N_6191,N_6196);
xnor U6259 (N_6259,N_6110,N_6181);
and U6260 (N_6260,N_6075,N_6048);
nand U6261 (N_6261,N_6176,N_6126);
and U6262 (N_6262,N_6081,N_6025);
nand U6263 (N_6263,N_6198,N_6087);
or U6264 (N_6264,N_6037,N_6101);
nand U6265 (N_6265,N_6017,N_6034);
nand U6266 (N_6266,N_6026,N_6094);
xnor U6267 (N_6267,N_6114,N_6007);
nand U6268 (N_6268,N_6154,N_6125);
nor U6269 (N_6269,N_6055,N_6049);
nor U6270 (N_6270,N_6050,N_6011);
or U6271 (N_6271,N_6004,N_6041);
nand U6272 (N_6272,N_6066,N_6009);
nand U6273 (N_6273,N_6088,N_6052);
and U6274 (N_6274,N_6132,N_6063);
or U6275 (N_6275,N_6021,N_6108);
nor U6276 (N_6276,N_6074,N_6036);
nand U6277 (N_6277,N_6156,N_6030);
xnor U6278 (N_6278,N_6032,N_6047);
and U6279 (N_6279,N_6148,N_6157);
nor U6280 (N_6280,N_6029,N_6138);
nand U6281 (N_6281,N_6115,N_6184);
nor U6282 (N_6282,N_6158,N_6056);
nor U6283 (N_6283,N_6189,N_6178);
xor U6284 (N_6284,N_6097,N_6147);
nor U6285 (N_6285,N_6182,N_6143);
and U6286 (N_6286,N_6090,N_6170);
nor U6287 (N_6287,N_6080,N_6123);
xnor U6288 (N_6288,N_6187,N_6109);
or U6289 (N_6289,N_6083,N_6027);
nor U6290 (N_6290,N_6064,N_6136);
and U6291 (N_6291,N_6010,N_6014);
nand U6292 (N_6292,N_6175,N_6134);
nor U6293 (N_6293,N_6107,N_6020);
nor U6294 (N_6294,N_6180,N_6005);
nor U6295 (N_6295,N_6044,N_6051);
nand U6296 (N_6296,N_6091,N_6024);
or U6297 (N_6297,N_6174,N_6054);
xor U6298 (N_6298,N_6160,N_6038);
xor U6299 (N_6299,N_6193,N_6137);
nand U6300 (N_6300,N_6014,N_6144);
xnor U6301 (N_6301,N_6157,N_6078);
or U6302 (N_6302,N_6100,N_6135);
or U6303 (N_6303,N_6004,N_6156);
xnor U6304 (N_6304,N_6137,N_6122);
nor U6305 (N_6305,N_6034,N_6113);
nand U6306 (N_6306,N_6027,N_6010);
nor U6307 (N_6307,N_6014,N_6174);
nand U6308 (N_6308,N_6141,N_6176);
nand U6309 (N_6309,N_6108,N_6189);
or U6310 (N_6310,N_6191,N_6162);
nor U6311 (N_6311,N_6004,N_6187);
nor U6312 (N_6312,N_6062,N_6007);
or U6313 (N_6313,N_6143,N_6029);
and U6314 (N_6314,N_6081,N_6160);
or U6315 (N_6315,N_6188,N_6001);
xnor U6316 (N_6316,N_6033,N_6074);
or U6317 (N_6317,N_6009,N_6159);
and U6318 (N_6318,N_6040,N_6092);
xor U6319 (N_6319,N_6125,N_6081);
nor U6320 (N_6320,N_6025,N_6165);
and U6321 (N_6321,N_6088,N_6082);
nand U6322 (N_6322,N_6173,N_6010);
nor U6323 (N_6323,N_6107,N_6169);
or U6324 (N_6324,N_6123,N_6173);
xor U6325 (N_6325,N_6036,N_6185);
nor U6326 (N_6326,N_6099,N_6182);
nand U6327 (N_6327,N_6065,N_6119);
nand U6328 (N_6328,N_6058,N_6012);
and U6329 (N_6329,N_6107,N_6186);
nand U6330 (N_6330,N_6139,N_6057);
xnor U6331 (N_6331,N_6082,N_6025);
nor U6332 (N_6332,N_6135,N_6196);
or U6333 (N_6333,N_6182,N_6076);
nand U6334 (N_6334,N_6083,N_6132);
and U6335 (N_6335,N_6033,N_6063);
or U6336 (N_6336,N_6022,N_6162);
xnor U6337 (N_6337,N_6016,N_6174);
nand U6338 (N_6338,N_6050,N_6071);
and U6339 (N_6339,N_6055,N_6026);
nor U6340 (N_6340,N_6194,N_6107);
and U6341 (N_6341,N_6016,N_6172);
or U6342 (N_6342,N_6132,N_6058);
or U6343 (N_6343,N_6057,N_6199);
and U6344 (N_6344,N_6190,N_6026);
nor U6345 (N_6345,N_6010,N_6158);
and U6346 (N_6346,N_6154,N_6138);
nor U6347 (N_6347,N_6184,N_6025);
and U6348 (N_6348,N_6128,N_6081);
and U6349 (N_6349,N_6063,N_6176);
nand U6350 (N_6350,N_6162,N_6128);
nor U6351 (N_6351,N_6002,N_6087);
or U6352 (N_6352,N_6034,N_6135);
nand U6353 (N_6353,N_6070,N_6095);
xor U6354 (N_6354,N_6124,N_6127);
nor U6355 (N_6355,N_6104,N_6023);
nor U6356 (N_6356,N_6001,N_6044);
nand U6357 (N_6357,N_6003,N_6053);
and U6358 (N_6358,N_6144,N_6142);
nand U6359 (N_6359,N_6172,N_6189);
nand U6360 (N_6360,N_6039,N_6126);
xnor U6361 (N_6361,N_6097,N_6068);
nand U6362 (N_6362,N_6122,N_6072);
nand U6363 (N_6363,N_6184,N_6172);
or U6364 (N_6364,N_6030,N_6109);
or U6365 (N_6365,N_6022,N_6149);
nand U6366 (N_6366,N_6035,N_6091);
nor U6367 (N_6367,N_6059,N_6055);
nor U6368 (N_6368,N_6054,N_6105);
or U6369 (N_6369,N_6185,N_6137);
nor U6370 (N_6370,N_6102,N_6080);
xnor U6371 (N_6371,N_6186,N_6094);
and U6372 (N_6372,N_6017,N_6199);
nor U6373 (N_6373,N_6081,N_6018);
nor U6374 (N_6374,N_6095,N_6040);
nor U6375 (N_6375,N_6128,N_6014);
nand U6376 (N_6376,N_6025,N_6090);
nor U6377 (N_6377,N_6069,N_6026);
nand U6378 (N_6378,N_6097,N_6064);
or U6379 (N_6379,N_6079,N_6104);
nor U6380 (N_6380,N_6191,N_6165);
nand U6381 (N_6381,N_6127,N_6080);
or U6382 (N_6382,N_6119,N_6029);
xnor U6383 (N_6383,N_6030,N_6117);
nor U6384 (N_6384,N_6048,N_6000);
nand U6385 (N_6385,N_6001,N_6161);
and U6386 (N_6386,N_6055,N_6101);
nor U6387 (N_6387,N_6066,N_6071);
nor U6388 (N_6388,N_6011,N_6078);
and U6389 (N_6389,N_6195,N_6049);
and U6390 (N_6390,N_6122,N_6035);
and U6391 (N_6391,N_6111,N_6090);
or U6392 (N_6392,N_6183,N_6101);
nor U6393 (N_6393,N_6081,N_6107);
and U6394 (N_6394,N_6009,N_6079);
and U6395 (N_6395,N_6015,N_6094);
nand U6396 (N_6396,N_6111,N_6192);
or U6397 (N_6397,N_6167,N_6140);
or U6398 (N_6398,N_6171,N_6059);
and U6399 (N_6399,N_6165,N_6159);
nor U6400 (N_6400,N_6207,N_6381);
nor U6401 (N_6401,N_6351,N_6296);
nand U6402 (N_6402,N_6334,N_6350);
and U6403 (N_6403,N_6211,N_6367);
nand U6404 (N_6404,N_6203,N_6247);
and U6405 (N_6405,N_6225,N_6290);
nor U6406 (N_6406,N_6213,N_6226);
nor U6407 (N_6407,N_6231,N_6310);
or U6408 (N_6408,N_6342,N_6284);
nor U6409 (N_6409,N_6388,N_6240);
nand U6410 (N_6410,N_6356,N_6341);
or U6411 (N_6411,N_6304,N_6220);
or U6412 (N_6412,N_6382,N_6317);
or U6413 (N_6413,N_6372,N_6201);
or U6414 (N_6414,N_6306,N_6359);
and U6415 (N_6415,N_6233,N_6303);
nand U6416 (N_6416,N_6320,N_6365);
nand U6417 (N_6417,N_6390,N_6238);
and U6418 (N_6418,N_6232,N_6222);
or U6419 (N_6419,N_6325,N_6254);
nor U6420 (N_6420,N_6312,N_6274);
or U6421 (N_6421,N_6364,N_6329);
nand U6422 (N_6422,N_6386,N_6266);
nand U6423 (N_6423,N_6383,N_6307);
xor U6424 (N_6424,N_6387,N_6309);
nand U6425 (N_6425,N_6328,N_6347);
or U6426 (N_6426,N_6379,N_6260);
nand U6427 (N_6427,N_6227,N_6346);
nand U6428 (N_6428,N_6316,N_6217);
or U6429 (N_6429,N_6242,N_6302);
and U6430 (N_6430,N_6327,N_6218);
or U6431 (N_6431,N_6270,N_6314);
nor U6432 (N_6432,N_6333,N_6300);
xor U6433 (N_6433,N_6361,N_6273);
or U6434 (N_6434,N_6249,N_6397);
or U6435 (N_6435,N_6208,N_6332);
and U6436 (N_6436,N_6338,N_6239);
nor U6437 (N_6437,N_6323,N_6398);
nand U6438 (N_6438,N_6371,N_6344);
or U6439 (N_6439,N_6308,N_6354);
nor U6440 (N_6440,N_6336,N_6214);
and U6441 (N_6441,N_6230,N_6264);
xor U6442 (N_6442,N_6395,N_6392);
or U6443 (N_6443,N_6283,N_6288);
nand U6444 (N_6444,N_6374,N_6298);
and U6445 (N_6445,N_6250,N_6315);
and U6446 (N_6446,N_6268,N_6362);
nand U6447 (N_6447,N_6202,N_6276);
and U6448 (N_6448,N_6272,N_6256);
or U6449 (N_6449,N_6293,N_6349);
and U6450 (N_6450,N_6205,N_6215);
xnor U6451 (N_6451,N_6339,N_6368);
or U6452 (N_6452,N_6209,N_6355);
nor U6453 (N_6453,N_6271,N_6258);
nor U6454 (N_6454,N_6311,N_6263);
nand U6455 (N_6455,N_6235,N_6357);
or U6456 (N_6456,N_6275,N_6352);
and U6457 (N_6457,N_6282,N_6399);
nor U6458 (N_6458,N_6391,N_6353);
nand U6459 (N_6459,N_6384,N_6378);
nor U6460 (N_6460,N_6219,N_6331);
nor U6461 (N_6461,N_6262,N_6380);
or U6462 (N_6462,N_6370,N_6321);
nor U6463 (N_6463,N_6301,N_6322);
xor U6464 (N_6464,N_6210,N_6394);
and U6465 (N_6465,N_6393,N_6377);
and U6466 (N_6466,N_6345,N_6376);
and U6467 (N_6467,N_6241,N_6281);
and U6468 (N_6468,N_6252,N_6236);
nor U6469 (N_6469,N_6337,N_6343);
nand U6470 (N_6470,N_6292,N_6277);
or U6471 (N_6471,N_6295,N_6212);
nand U6472 (N_6472,N_6363,N_6385);
or U6473 (N_6473,N_6253,N_6335);
xor U6474 (N_6474,N_6305,N_6265);
or U6475 (N_6475,N_6286,N_6245);
nand U6476 (N_6476,N_6279,N_6259);
nand U6477 (N_6477,N_6267,N_6285);
nor U6478 (N_6478,N_6200,N_6291);
and U6479 (N_6479,N_6237,N_6216);
or U6480 (N_6480,N_6330,N_6299);
or U6481 (N_6481,N_6278,N_6229);
xnor U6482 (N_6482,N_6221,N_6369);
nor U6483 (N_6483,N_6251,N_6396);
or U6484 (N_6484,N_6280,N_6324);
and U6485 (N_6485,N_6248,N_6389);
or U6486 (N_6486,N_6246,N_6366);
nand U6487 (N_6487,N_6326,N_6319);
xnor U6488 (N_6488,N_6228,N_6269);
nor U6489 (N_6489,N_6223,N_6257);
nor U6490 (N_6490,N_6224,N_6287);
nor U6491 (N_6491,N_6318,N_6289);
nor U6492 (N_6492,N_6360,N_6255);
nor U6493 (N_6493,N_6297,N_6244);
or U6494 (N_6494,N_6261,N_6234);
and U6495 (N_6495,N_6348,N_6358);
and U6496 (N_6496,N_6373,N_6340);
nand U6497 (N_6497,N_6313,N_6204);
or U6498 (N_6498,N_6294,N_6375);
nand U6499 (N_6499,N_6206,N_6243);
or U6500 (N_6500,N_6345,N_6343);
and U6501 (N_6501,N_6345,N_6222);
and U6502 (N_6502,N_6268,N_6297);
nor U6503 (N_6503,N_6365,N_6231);
and U6504 (N_6504,N_6356,N_6266);
nor U6505 (N_6505,N_6321,N_6368);
xor U6506 (N_6506,N_6356,N_6379);
nor U6507 (N_6507,N_6209,N_6368);
nand U6508 (N_6508,N_6307,N_6305);
or U6509 (N_6509,N_6373,N_6386);
or U6510 (N_6510,N_6209,N_6215);
nor U6511 (N_6511,N_6275,N_6319);
or U6512 (N_6512,N_6327,N_6355);
or U6513 (N_6513,N_6322,N_6283);
and U6514 (N_6514,N_6313,N_6373);
xor U6515 (N_6515,N_6308,N_6219);
nor U6516 (N_6516,N_6367,N_6274);
nand U6517 (N_6517,N_6303,N_6250);
and U6518 (N_6518,N_6258,N_6228);
nand U6519 (N_6519,N_6294,N_6318);
xnor U6520 (N_6520,N_6385,N_6312);
xor U6521 (N_6521,N_6358,N_6225);
nand U6522 (N_6522,N_6274,N_6303);
or U6523 (N_6523,N_6239,N_6380);
and U6524 (N_6524,N_6298,N_6276);
nor U6525 (N_6525,N_6383,N_6243);
nand U6526 (N_6526,N_6275,N_6336);
nor U6527 (N_6527,N_6387,N_6366);
and U6528 (N_6528,N_6201,N_6232);
nand U6529 (N_6529,N_6259,N_6218);
nand U6530 (N_6530,N_6333,N_6244);
nor U6531 (N_6531,N_6268,N_6339);
nand U6532 (N_6532,N_6365,N_6371);
nand U6533 (N_6533,N_6349,N_6372);
nand U6534 (N_6534,N_6284,N_6277);
nand U6535 (N_6535,N_6263,N_6281);
and U6536 (N_6536,N_6307,N_6263);
nand U6537 (N_6537,N_6380,N_6264);
and U6538 (N_6538,N_6214,N_6281);
or U6539 (N_6539,N_6346,N_6339);
nor U6540 (N_6540,N_6227,N_6270);
or U6541 (N_6541,N_6365,N_6322);
nor U6542 (N_6542,N_6251,N_6233);
nor U6543 (N_6543,N_6300,N_6388);
nor U6544 (N_6544,N_6228,N_6312);
nor U6545 (N_6545,N_6278,N_6276);
nand U6546 (N_6546,N_6228,N_6208);
and U6547 (N_6547,N_6202,N_6215);
or U6548 (N_6548,N_6397,N_6339);
or U6549 (N_6549,N_6365,N_6288);
nor U6550 (N_6550,N_6330,N_6305);
and U6551 (N_6551,N_6392,N_6256);
nor U6552 (N_6552,N_6224,N_6265);
nand U6553 (N_6553,N_6318,N_6271);
and U6554 (N_6554,N_6368,N_6267);
nand U6555 (N_6555,N_6383,N_6283);
xor U6556 (N_6556,N_6310,N_6236);
nand U6557 (N_6557,N_6313,N_6322);
and U6558 (N_6558,N_6238,N_6370);
nor U6559 (N_6559,N_6353,N_6387);
nor U6560 (N_6560,N_6268,N_6260);
nand U6561 (N_6561,N_6358,N_6260);
nand U6562 (N_6562,N_6346,N_6213);
and U6563 (N_6563,N_6223,N_6212);
xor U6564 (N_6564,N_6385,N_6296);
nand U6565 (N_6565,N_6365,N_6235);
and U6566 (N_6566,N_6256,N_6262);
and U6567 (N_6567,N_6232,N_6376);
xnor U6568 (N_6568,N_6238,N_6271);
nand U6569 (N_6569,N_6297,N_6374);
and U6570 (N_6570,N_6370,N_6352);
nor U6571 (N_6571,N_6256,N_6234);
nor U6572 (N_6572,N_6336,N_6341);
nand U6573 (N_6573,N_6357,N_6208);
and U6574 (N_6574,N_6204,N_6301);
and U6575 (N_6575,N_6224,N_6321);
nor U6576 (N_6576,N_6221,N_6390);
xor U6577 (N_6577,N_6318,N_6214);
xor U6578 (N_6578,N_6356,N_6255);
or U6579 (N_6579,N_6213,N_6352);
nor U6580 (N_6580,N_6275,N_6288);
nand U6581 (N_6581,N_6210,N_6334);
or U6582 (N_6582,N_6373,N_6210);
nor U6583 (N_6583,N_6227,N_6364);
or U6584 (N_6584,N_6393,N_6252);
or U6585 (N_6585,N_6343,N_6229);
or U6586 (N_6586,N_6335,N_6342);
nor U6587 (N_6587,N_6252,N_6226);
nor U6588 (N_6588,N_6254,N_6382);
nor U6589 (N_6589,N_6259,N_6210);
nor U6590 (N_6590,N_6276,N_6270);
or U6591 (N_6591,N_6390,N_6376);
nor U6592 (N_6592,N_6231,N_6383);
nand U6593 (N_6593,N_6329,N_6304);
nor U6594 (N_6594,N_6258,N_6314);
nor U6595 (N_6595,N_6342,N_6399);
nand U6596 (N_6596,N_6351,N_6298);
xor U6597 (N_6597,N_6354,N_6234);
nand U6598 (N_6598,N_6336,N_6265);
or U6599 (N_6599,N_6228,N_6398);
nor U6600 (N_6600,N_6505,N_6520);
and U6601 (N_6601,N_6416,N_6445);
nor U6602 (N_6602,N_6461,N_6471);
or U6603 (N_6603,N_6495,N_6443);
nand U6604 (N_6604,N_6563,N_6430);
nand U6605 (N_6605,N_6433,N_6540);
or U6606 (N_6606,N_6590,N_6537);
and U6607 (N_6607,N_6467,N_6525);
and U6608 (N_6608,N_6411,N_6489);
or U6609 (N_6609,N_6418,N_6577);
nand U6610 (N_6610,N_6484,N_6476);
and U6611 (N_6611,N_6557,N_6569);
and U6612 (N_6612,N_6474,N_6510);
and U6613 (N_6613,N_6522,N_6579);
nor U6614 (N_6614,N_6555,N_6570);
or U6615 (N_6615,N_6500,N_6400);
and U6616 (N_6616,N_6425,N_6597);
or U6617 (N_6617,N_6437,N_6539);
and U6618 (N_6618,N_6465,N_6409);
and U6619 (N_6619,N_6492,N_6571);
and U6620 (N_6620,N_6415,N_6533);
xor U6621 (N_6621,N_6454,N_6482);
or U6622 (N_6622,N_6512,N_6527);
nor U6623 (N_6623,N_6462,N_6450);
nor U6624 (N_6624,N_6548,N_6503);
nor U6625 (N_6625,N_6536,N_6594);
nand U6626 (N_6626,N_6405,N_6432);
and U6627 (N_6627,N_6480,N_6598);
nor U6628 (N_6628,N_6568,N_6434);
and U6629 (N_6629,N_6456,N_6567);
nor U6630 (N_6630,N_6517,N_6499);
or U6631 (N_6631,N_6421,N_6424);
nand U6632 (N_6632,N_6573,N_6401);
nand U6633 (N_6633,N_6488,N_6459);
and U6634 (N_6634,N_6513,N_6455);
nand U6635 (N_6635,N_6560,N_6408);
and U6636 (N_6636,N_6559,N_6477);
nand U6637 (N_6637,N_6506,N_6578);
nor U6638 (N_6638,N_6549,N_6588);
and U6639 (N_6639,N_6413,N_6523);
or U6640 (N_6640,N_6486,N_6496);
nand U6641 (N_6641,N_6550,N_6420);
and U6642 (N_6642,N_6426,N_6404);
or U6643 (N_6643,N_6453,N_6448);
nand U6644 (N_6644,N_6419,N_6532);
nor U6645 (N_6645,N_6584,N_6435);
or U6646 (N_6646,N_6410,N_6516);
nand U6647 (N_6647,N_6468,N_6436);
nor U6648 (N_6648,N_6572,N_6552);
and U6649 (N_6649,N_6494,N_6591);
nor U6650 (N_6650,N_6429,N_6514);
or U6651 (N_6651,N_6478,N_6534);
and U6652 (N_6652,N_6442,N_6530);
and U6653 (N_6653,N_6509,N_6464);
nor U6654 (N_6654,N_6491,N_6451);
nand U6655 (N_6655,N_6439,N_6406);
nor U6656 (N_6656,N_6566,N_6490);
nand U6657 (N_6657,N_6466,N_6551);
and U6658 (N_6658,N_6561,N_6447);
nor U6659 (N_6659,N_6581,N_6515);
and U6660 (N_6660,N_6528,N_6402);
nand U6661 (N_6661,N_6423,N_6595);
or U6662 (N_6662,N_6504,N_6586);
nand U6663 (N_6663,N_6449,N_6583);
nor U6664 (N_6664,N_6556,N_6526);
or U6665 (N_6665,N_6498,N_6481);
xnor U6666 (N_6666,N_6538,N_6440);
nand U6667 (N_6667,N_6599,N_6529);
nor U6668 (N_6668,N_6587,N_6483);
nor U6669 (N_6669,N_6502,N_6427);
nor U6670 (N_6670,N_6441,N_6546);
nand U6671 (N_6671,N_6545,N_6507);
nor U6672 (N_6672,N_6508,N_6589);
or U6673 (N_6673,N_6497,N_6547);
xnor U6674 (N_6674,N_6511,N_6414);
or U6675 (N_6675,N_6558,N_6457);
nor U6676 (N_6676,N_6501,N_6565);
xnor U6677 (N_6677,N_6458,N_6428);
or U6678 (N_6678,N_6438,N_6576);
nand U6679 (N_6679,N_6479,N_6554);
and U6680 (N_6680,N_6582,N_6485);
and U6681 (N_6681,N_6519,N_6472);
xor U6682 (N_6682,N_6562,N_6596);
nor U6683 (N_6683,N_6593,N_6544);
nor U6684 (N_6684,N_6407,N_6553);
nand U6685 (N_6685,N_6487,N_6444);
nand U6686 (N_6686,N_6475,N_6524);
and U6687 (N_6687,N_6493,N_6422);
and U6688 (N_6688,N_6535,N_6564);
or U6689 (N_6689,N_6575,N_6518);
nor U6690 (N_6690,N_6412,N_6469);
nand U6691 (N_6691,N_6417,N_6542);
and U6692 (N_6692,N_6531,N_6473);
and U6693 (N_6693,N_6580,N_6452);
or U6694 (N_6694,N_6431,N_6543);
nor U6695 (N_6695,N_6470,N_6460);
xor U6696 (N_6696,N_6403,N_6574);
nor U6697 (N_6697,N_6463,N_6585);
or U6698 (N_6698,N_6541,N_6592);
xnor U6699 (N_6699,N_6446,N_6521);
nor U6700 (N_6700,N_6428,N_6555);
nor U6701 (N_6701,N_6454,N_6548);
nor U6702 (N_6702,N_6468,N_6513);
and U6703 (N_6703,N_6417,N_6547);
and U6704 (N_6704,N_6475,N_6546);
nand U6705 (N_6705,N_6576,N_6541);
xor U6706 (N_6706,N_6501,N_6481);
and U6707 (N_6707,N_6503,N_6464);
nor U6708 (N_6708,N_6537,N_6549);
nand U6709 (N_6709,N_6531,N_6406);
or U6710 (N_6710,N_6537,N_6403);
nand U6711 (N_6711,N_6439,N_6533);
xor U6712 (N_6712,N_6533,N_6536);
or U6713 (N_6713,N_6571,N_6550);
and U6714 (N_6714,N_6437,N_6491);
nor U6715 (N_6715,N_6509,N_6479);
or U6716 (N_6716,N_6541,N_6451);
and U6717 (N_6717,N_6478,N_6481);
or U6718 (N_6718,N_6489,N_6527);
or U6719 (N_6719,N_6503,N_6557);
and U6720 (N_6720,N_6426,N_6443);
nand U6721 (N_6721,N_6594,N_6466);
nand U6722 (N_6722,N_6546,N_6522);
or U6723 (N_6723,N_6406,N_6515);
nand U6724 (N_6724,N_6418,N_6492);
or U6725 (N_6725,N_6420,N_6548);
nand U6726 (N_6726,N_6581,N_6501);
xor U6727 (N_6727,N_6413,N_6562);
nand U6728 (N_6728,N_6555,N_6458);
and U6729 (N_6729,N_6451,N_6577);
and U6730 (N_6730,N_6411,N_6479);
nand U6731 (N_6731,N_6465,N_6467);
or U6732 (N_6732,N_6564,N_6516);
and U6733 (N_6733,N_6492,N_6528);
nand U6734 (N_6734,N_6494,N_6480);
and U6735 (N_6735,N_6477,N_6524);
and U6736 (N_6736,N_6516,N_6505);
xor U6737 (N_6737,N_6516,N_6404);
xor U6738 (N_6738,N_6583,N_6402);
or U6739 (N_6739,N_6403,N_6414);
nand U6740 (N_6740,N_6594,N_6412);
xor U6741 (N_6741,N_6490,N_6463);
nor U6742 (N_6742,N_6459,N_6476);
nand U6743 (N_6743,N_6511,N_6432);
xnor U6744 (N_6744,N_6460,N_6414);
nor U6745 (N_6745,N_6472,N_6414);
or U6746 (N_6746,N_6599,N_6511);
nor U6747 (N_6747,N_6424,N_6535);
xnor U6748 (N_6748,N_6466,N_6450);
xnor U6749 (N_6749,N_6533,N_6442);
nor U6750 (N_6750,N_6538,N_6592);
or U6751 (N_6751,N_6583,N_6589);
xnor U6752 (N_6752,N_6584,N_6467);
nor U6753 (N_6753,N_6551,N_6494);
and U6754 (N_6754,N_6468,N_6472);
or U6755 (N_6755,N_6500,N_6582);
and U6756 (N_6756,N_6448,N_6530);
nor U6757 (N_6757,N_6406,N_6475);
or U6758 (N_6758,N_6592,N_6447);
nand U6759 (N_6759,N_6574,N_6595);
nand U6760 (N_6760,N_6548,N_6577);
nor U6761 (N_6761,N_6571,N_6430);
nor U6762 (N_6762,N_6556,N_6521);
or U6763 (N_6763,N_6569,N_6471);
nand U6764 (N_6764,N_6449,N_6466);
or U6765 (N_6765,N_6486,N_6564);
or U6766 (N_6766,N_6568,N_6445);
and U6767 (N_6767,N_6415,N_6410);
and U6768 (N_6768,N_6476,N_6576);
nor U6769 (N_6769,N_6459,N_6553);
and U6770 (N_6770,N_6489,N_6416);
nor U6771 (N_6771,N_6554,N_6576);
nand U6772 (N_6772,N_6504,N_6518);
or U6773 (N_6773,N_6582,N_6497);
nand U6774 (N_6774,N_6518,N_6435);
or U6775 (N_6775,N_6446,N_6537);
nor U6776 (N_6776,N_6465,N_6511);
or U6777 (N_6777,N_6468,N_6593);
nor U6778 (N_6778,N_6555,N_6553);
xnor U6779 (N_6779,N_6484,N_6430);
or U6780 (N_6780,N_6517,N_6501);
nand U6781 (N_6781,N_6496,N_6559);
or U6782 (N_6782,N_6427,N_6549);
nand U6783 (N_6783,N_6466,N_6575);
xor U6784 (N_6784,N_6593,N_6570);
nand U6785 (N_6785,N_6454,N_6528);
xnor U6786 (N_6786,N_6520,N_6461);
and U6787 (N_6787,N_6583,N_6502);
or U6788 (N_6788,N_6530,N_6491);
nor U6789 (N_6789,N_6514,N_6576);
nor U6790 (N_6790,N_6411,N_6501);
nor U6791 (N_6791,N_6513,N_6590);
and U6792 (N_6792,N_6450,N_6428);
nand U6793 (N_6793,N_6566,N_6433);
or U6794 (N_6794,N_6462,N_6569);
or U6795 (N_6795,N_6422,N_6525);
nand U6796 (N_6796,N_6510,N_6483);
or U6797 (N_6797,N_6568,N_6577);
nor U6798 (N_6798,N_6468,N_6522);
nor U6799 (N_6799,N_6499,N_6527);
xor U6800 (N_6800,N_6757,N_6618);
or U6801 (N_6801,N_6731,N_6630);
nand U6802 (N_6802,N_6662,N_6667);
nand U6803 (N_6803,N_6775,N_6623);
or U6804 (N_6804,N_6716,N_6733);
nand U6805 (N_6805,N_6639,N_6713);
or U6806 (N_6806,N_6682,N_6719);
and U6807 (N_6807,N_6675,N_6688);
or U6808 (N_6808,N_6786,N_6656);
nand U6809 (N_6809,N_6681,N_6680);
nor U6810 (N_6810,N_6619,N_6717);
nor U6811 (N_6811,N_6777,N_6749);
nand U6812 (N_6812,N_6787,N_6760);
and U6813 (N_6813,N_6774,N_6730);
nand U6814 (N_6814,N_6726,N_6694);
xnor U6815 (N_6815,N_6615,N_6782);
and U6816 (N_6816,N_6651,N_6746);
and U6817 (N_6817,N_6699,N_6710);
nor U6818 (N_6818,N_6744,N_6785);
or U6819 (N_6819,N_6748,N_6658);
or U6820 (N_6820,N_6764,N_6634);
nand U6821 (N_6821,N_6752,N_6758);
nand U6822 (N_6822,N_6720,N_6799);
and U6823 (N_6823,N_6763,N_6700);
and U6824 (N_6824,N_6628,N_6795);
nor U6825 (N_6825,N_6741,N_6684);
nor U6826 (N_6826,N_6709,N_6756);
nor U6827 (N_6827,N_6685,N_6707);
or U6828 (N_6828,N_6725,N_6626);
nand U6829 (N_6829,N_6621,N_6704);
or U6830 (N_6830,N_6672,N_6732);
and U6831 (N_6831,N_6687,N_6692);
or U6832 (N_6832,N_6691,N_6724);
nand U6833 (N_6833,N_6759,N_6705);
nand U6834 (N_6834,N_6772,N_6792);
nor U6835 (N_6835,N_6788,N_6701);
xnor U6836 (N_6836,N_6797,N_6722);
nor U6837 (N_6837,N_6766,N_6604);
nand U6838 (N_6838,N_6611,N_6755);
or U6839 (N_6839,N_6646,N_6649);
nand U6840 (N_6840,N_6796,N_6650);
or U6841 (N_6841,N_6671,N_6762);
and U6842 (N_6842,N_6613,N_6737);
or U6843 (N_6843,N_6683,N_6603);
and U6844 (N_6844,N_6696,N_6614);
or U6845 (N_6845,N_6714,N_6769);
xnor U6846 (N_6846,N_6712,N_6703);
nand U6847 (N_6847,N_6711,N_6776);
nand U6848 (N_6848,N_6745,N_6622);
nand U6849 (N_6849,N_6729,N_6693);
nand U6850 (N_6850,N_6686,N_6679);
or U6851 (N_6851,N_6754,N_6616);
nand U6852 (N_6852,N_6770,N_6697);
nor U6853 (N_6853,N_6750,N_6609);
xor U6854 (N_6854,N_6631,N_6783);
or U6855 (N_6855,N_6640,N_6659);
nor U6856 (N_6856,N_6647,N_6641);
or U6857 (N_6857,N_6663,N_6718);
nand U6858 (N_6858,N_6723,N_6765);
or U6859 (N_6859,N_6602,N_6654);
nand U6860 (N_6860,N_6689,N_6624);
nand U6861 (N_6861,N_6668,N_6753);
nand U6862 (N_6862,N_6698,N_6644);
and U6863 (N_6863,N_6665,N_6791);
and U6864 (N_6864,N_6768,N_6735);
or U6865 (N_6865,N_6798,N_6678);
and U6866 (N_6866,N_6767,N_6661);
nor U6867 (N_6867,N_6600,N_6620);
nor U6868 (N_6868,N_6612,N_6653);
and U6869 (N_6869,N_6690,N_6642);
and U6870 (N_6870,N_6625,N_6666);
nand U6871 (N_6871,N_6738,N_6761);
or U6872 (N_6872,N_6633,N_6778);
nor U6873 (N_6873,N_6677,N_6664);
or U6874 (N_6874,N_6739,N_6648);
or U6875 (N_6875,N_6632,N_6734);
xor U6876 (N_6876,N_6617,N_6608);
xor U6877 (N_6877,N_6715,N_6706);
nand U6878 (N_6878,N_6660,N_6784);
nand U6879 (N_6879,N_6652,N_6674);
or U6880 (N_6880,N_6789,N_6607);
and U6881 (N_6881,N_6742,N_6610);
or U6882 (N_6882,N_6751,N_6779);
and U6883 (N_6883,N_6601,N_6629);
and U6884 (N_6884,N_6605,N_6669);
and U6885 (N_6885,N_6708,N_6773);
nand U6886 (N_6886,N_6636,N_6670);
and U6887 (N_6887,N_6771,N_6747);
nor U6888 (N_6888,N_6676,N_6794);
xnor U6889 (N_6889,N_6702,N_6637);
or U6890 (N_6890,N_6728,N_6780);
and U6891 (N_6891,N_6635,N_6727);
nor U6892 (N_6892,N_6790,N_6645);
or U6893 (N_6893,N_6638,N_6655);
nand U6894 (N_6894,N_6743,N_6736);
xnor U6895 (N_6895,N_6657,N_6673);
and U6896 (N_6896,N_6627,N_6793);
and U6897 (N_6897,N_6606,N_6781);
nor U6898 (N_6898,N_6740,N_6643);
nand U6899 (N_6899,N_6695,N_6721);
or U6900 (N_6900,N_6639,N_6688);
and U6901 (N_6901,N_6664,N_6611);
nand U6902 (N_6902,N_6695,N_6799);
or U6903 (N_6903,N_6727,N_6715);
xnor U6904 (N_6904,N_6759,N_6628);
or U6905 (N_6905,N_6692,N_6683);
nor U6906 (N_6906,N_6741,N_6746);
xor U6907 (N_6907,N_6678,N_6784);
and U6908 (N_6908,N_6771,N_6764);
nand U6909 (N_6909,N_6660,N_6674);
or U6910 (N_6910,N_6726,N_6727);
nor U6911 (N_6911,N_6704,N_6695);
nand U6912 (N_6912,N_6775,N_6641);
nor U6913 (N_6913,N_6687,N_6627);
nand U6914 (N_6914,N_6799,N_6775);
nand U6915 (N_6915,N_6787,N_6697);
nor U6916 (N_6916,N_6652,N_6796);
and U6917 (N_6917,N_6636,N_6681);
nor U6918 (N_6918,N_6718,N_6648);
nor U6919 (N_6919,N_6609,N_6650);
xnor U6920 (N_6920,N_6671,N_6626);
and U6921 (N_6921,N_6755,N_6733);
xor U6922 (N_6922,N_6706,N_6729);
and U6923 (N_6923,N_6788,N_6747);
nor U6924 (N_6924,N_6674,N_6612);
nor U6925 (N_6925,N_6679,N_6749);
or U6926 (N_6926,N_6733,N_6760);
or U6927 (N_6927,N_6604,N_6793);
nor U6928 (N_6928,N_6600,N_6756);
nand U6929 (N_6929,N_6667,N_6689);
or U6930 (N_6930,N_6648,N_6687);
and U6931 (N_6931,N_6637,N_6753);
or U6932 (N_6932,N_6751,N_6612);
nor U6933 (N_6933,N_6793,N_6748);
nor U6934 (N_6934,N_6668,N_6620);
nand U6935 (N_6935,N_6607,N_6678);
or U6936 (N_6936,N_6627,N_6730);
nor U6937 (N_6937,N_6684,N_6657);
or U6938 (N_6938,N_6724,N_6769);
nand U6939 (N_6939,N_6776,N_6610);
or U6940 (N_6940,N_6630,N_6783);
or U6941 (N_6941,N_6601,N_6709);
nor U6942 (N_6942,N_6657,N_6665);
nor U6943 (N_6943,N_6729,N_6659);
nand U6944 (N_6944,N_6751,N_6657);
xor U6945 (N_6945,N_6726,N_6662);
nand U6946 (N_6946,N_6787,N_6781);
or U6947 (N_6947,N_6604,N_6693);
and U6948 (N_6948,N_6644,N_6681);
nand U6949 (N_6949,N_6746,N_6788);
nor U6950 (N_6950,N_6716,N_6670);
or U6951 (N_6951,N_6648,N_6665);
or U6952 (N_6952,N_6777,N_6785);
and U6953 (N_6953,N_6734,N_6600);
nor U6954 (N_6954,N_6735,N_6707);
nand U6955 (N_6955,N_6620,N_6643);
xnor U6956 (N_6956,N_6698,N_6621);
nand U6957 (N_6957,N_6760,N_6694);
nand U6958 (N_6958,N_6643,N_6710);
and U6959 (N_6959,N_6608,N_6755);
nor U6960 (N_6960,N_6694,N_6772);
or U6961 (N_6961,N_6699,N_6687);
nor U6962 (N_6962,N_6760,N_6695);
nor U6963 (N_6963,N_6749,N_6625);
and U6964 (N_6964,N_6622,N_6693);
or U6965 (N_6965,N_6630,N_6680);
nor U6966 (N_6966,N_6737,N_6775);
and U6967 (N_6967,N_6661,N_6792);
nand U6968 (N_6968,N_6730,N_6623);
nand U6969 (N_6969,N_6794,N_6738);
or U6970 (N_6970,N_6697,N_6680);
nor U6971 (N_6971,N_6749,N_6758);
nand U6972 (N_6972,N_6743,N_6650);
nand U6973 (N_6973,N_6738,N_6661);
nor U6974 (N_6974,N_6615,N_6600);
nand U6975 (N_6975,N_6602,N_6771);
xor U6976 (N_6976,N_6794,N_6725);
nor U6977 (N_6977,N_6623,N_6628);
xnor U6978 (N_6978,N_6762,N_6763);
or U6979 (N_6979,N_6649,N_6700);
nor U6980 (N_6980,N_6622,N_6643);
xnor U6981 (N_6981,N_6706,N_6638);
and U6982 (N_6982,N_6791,N_6708);
and U6983 (N_6983,N_6752,N_6607);
nor U6984 (N_6984,N_6635,N_6749);
nor U6985 (N_6985,N_6770,N_6616);
nand U6986 (N_6986,N_6783,N_6693);
xnor U6987 (N_6987,N_6639,N_6747);
or U6988 (N_6988,N_6684,N_6786);
or U6989 (N_6989,N_6733,N_6717);
and U6990 (N_6990,N_6707,N_6633);
or U6991 (N_6991,N_6777,N_6746);
nand U6992 (N_6992,N_6794,N_6718);
or U6993 (N_6993,N_6679,N_6681);
nor U6994 (N_6994,N_6767,N_6778);
and U6995 (N_6995,N_6689,N_6686);
or U6996 (N_6996,N_6621,N_6645);
nand U6997 (N_6997,N_6782,N_6635);
nor U6998 (N_6998,N_6759,N_6728);
nand U6999 (N_6999,N_6609,N_6794);
nand U7000 (N_7000,N_6903,N_6910);
and U7001 (N_7001,N_6886,N_6883);
or U7002 (N_7002,N_6934,N_6956);
nand U7003 (N_7003,N_6999,N_6982);
or U7004 (N_7004,N_6844,N_6894);
nor U7005 (N_7005,N_6897,N_6817);
nor U7006 (N_7006,N_6935,N_6841);
or U7007 (N_7007,N_6834,N_6987);
and U7008 (N_7008,N_6809,N_6976);
nand U7009 (N_7009,N_6922,N_6898);
and U7010 (N_7010,N_6973,N_6947);
or U7011 (N_7011,N_6953,N_6891);
or U7012 (N_7012,N_6871,N_6905);
nor U7013 (N_7013,N_6948,N_6870);
xnor U7014 (N_7014,N_6901,N_6983);
nor U7015 (N_7015,N_6994,N_6885);
and U7016 (N_7016,N_6992,N_6881);
and U7017 (N_7017,N_6907,N_6825);
nand U7018 (N_7018,N_6951,N_6920);
or U7019 (N_7019,N_6832,N_6971);
nor U7020 (N_7020,N_6872,N_6944);
nor U7021 (N_7021,N_6830,N_6968);
nand U7022 (N_7022,N_6923,N_6991);
or U7023 (N_7023,N_6807,N_6842);
or U7024 (N_7024,N_6854,N_6926);
nor U7025 (N_7025,N_6873,N_6952);
and U7026 (N_7026,N_6833,N_6985);
nand U7027 (N_7027,N_6917,N_6853);
nor U7028 (N_7028,N_6965,N_6902);
nor U7029 (N_7029,N_6890,N_6859);
or U7030 (N_7030,N_6846,N_6851);
xor U7031 (N_7031,N_6823,N_6984);
nand U7032 (N_7032,N_6880,N_6961);
or U7033 (N_7033,N_6889,N_6840);
nand U7034 (N_7034,N_6915,N_6927);
or U7035 (N_7035,N_6929,N_6812);
nand U7036 (N_7036,N_6869,N_6946);
and U7037 (N_7037,N_6866,N_6845);
nor U7038 (N_7038,N_6852,N_6925);
xnor U7039 (N_7039,N_6964,N_6822);
or U7040 (N_7040,N_6867,N_6954);
and U7041 (N_7041,N_6950,N_6814);
or U7042 (N_7042,N_6932,N_6824);
nand U7043 (N_7043,N_6997,N_6818);
nand U7044 (N_7044,N_6801,N_6820);
or U7045 (N_7045,N_6969,N_6865);
nand U7046 (N_7046,N_6868,N_6943);
or U7047 (N_7047,N_6970,N_6989);
nor U7048 (N_7048,N_6908,N_6916);
nand U7049 (N_7049,N_6937,N_6849);
nand U7050 (N_7050,N_6936,N_6863);
or U7051 (N_7051,N_6836,N_6924);
nand U7052 (N_7052,N_6888,N_6913);
nor U7053 (N_7053,N_6835,N_6979);
or U7054 (N_7054,N_6877,N_6959);
or U7055 (N_7055,N_6843,N_6899);
nand U7056 (N_7056,N_6806,N_6831);
xnor U7057 (N_7057,N_6904,N_6933);
or U7058 (N_7058,N_6914,N_6819);
nand U7059 (N_7059,N_6860,N_6805);
nand U7060 (N_7060,N_6998,N_6939);
nand U7061 (N_7061,N_6942,N_6804);
nor U7062 (N_7062,N_6856,N_6847);
nor U7063 (N_7063,N_6990,N_6988);
nand U7064 (N_7064,N_6957,N_6827);
xnor U7065 (N_7065,N_6815,N_6975);
xor U7066 (N_7066,N_6900,N_6887);
nor U7067 (N_7067,N_6803,N_6878);
or U7068 (N_7068,N_6955,N_6921);
nand U7069 (N_7069,N_6940,N_6978);
or U7070 (N_7070,N_6839,N_6972);
and U7071 (N_7071,N_6967,N_6893);
or U7072 (N_7072,N_6816,N_6855);
xor U7073 (N_7073,N_6945,N_6996);
nor U7074 (N_7074,N_6864,N_6938);
or U7075 (N_7075,N_6962,N_6980);
xnor U7076 (N_7076,N_6837,N_6918);
nor U7077 (N_7077,N_6829,N_6960);
or U7078 (N_7078,N_6949,N_6857);
or U7079 (N_7079,N_6874,N_6862);
nand U7080 (N_7080,N_6958,N_6966);
nor U7081 (N_7081,N_6906,N_6993);
or U7082 (N_7082,N_6882,N_6802);
nor U7083 (N_7083,N_6912,N_6981);
nand U7084 (N_7084,N_6808,N_6974);
and U7085 (N_7085,N_6963,N_6931);
nand U7086 (N_7086,N_6892,N_6919);
and U7087 (N_7087,N_6811,N_6875);
or U7088 (N_7088,N_6821,N_6828);
and U7089 (N_7089,N_6858,N_6848);
and U7090 (N_7090,N_6800,N_6861);
nand U7091 (N_7091,N_6986,N_6879);
nor U7092 (N_7092,N_6941,N_6895);
nor U7093 (N_7093,N_6911,N_6838);
nor U7094 (N_7094,N_6977,N_6813);
nor U7095 (N_7095,N_6876,N_6909);
and U7096 (N_7096,N_6810,N_6930);
or U7097 (N_7097,N_6850,N_6884);
nor U7098 (N_7098,N_6826,N_6995);
or U7099 (N_7099,N_6928,N_6896);
or U7100 (N_7100,N_6927,N_6878);
nand U7101 (N_7101,N_6997,N_6955);
and U7102 (N_7102,N_6887,N_6910);
or U7103 (N_7103,N_6919,N_6971);
xnor U7104 (N_7104,N_6853,N_6900);
nor U7105 (N_7105,N_6963,N_6893);
nor U7106 (N_7106,N_6981,N_6881);
nand U7107 (N_7107,N_6925,N_6814);
nand U7108 (N_7108,N_6804,N_6833);
nor U7109 (N_7109,N_6872,N_6817);
and U7110 (N_7110,N_6982,N_6919);
nor U7111 (N_7111,N_6904,N_6896);
and U7112 (N_7112,N_6943,N_6808);
nor U7113 (N_7113,N_6924,N_6821);
xnor U7114 (N_7114,N_6920,N_6894);
nand U7115 (N_7115,N_6844,N_6889);
nor U7116 (N_7116,N_6912,N_6815);
xor U7117 (N_7117,N_6805,N_6950);
and U7118 (N_7118,N_6976,N_6897);
nand U7119 (N_7119,N_6889,N_6919);
or U7120 (N_7120,N_6875,N_6835);
xor U7121 (N_7121,N_6959,N_6933);
and U7122 (N_7122,N_6856,N_6941);
nand U7123 (N_7123,N_6925,N_6886);
or U7124 (N_7124,N_6820,N_6846);
nor U7125 (N_7125,N_6802,N_6934);
xor U7126 (N_7126,N_6992,N_6912);
nor U7127 (N_7127,N_6832,N_6997);
nand U7128 (N_7128,N_6989,N_6836);
nor U7129 (N_7129,N_6862,N_6886);
nand U7130 (N_7130,N_6897,N_6994);
nor U7131 (N_7131,N_6827,N_6927);
and U7132 (N_7132,N_6823,N_6807);
or U7133 (N_7133,N_6951,N_6845);
and U7134 (N_7134,N_6868,N_6908);
nand U7135 (N_7135,N_6940,N_6801);
nor U7136 (N_7136,N_6852,N_6886);
nand U7137 (N_7137,N_6979,N_6964);
and U7138 (N_7138,N_6856,N_6878);
nor U7139 (N_7139,N_6845,N_6831);
nand U7140 (N_7140,N_6989,N_6849);
or U7141 (N_7141,N_6858,N_6862);
nor U7142 (N_7142,N_6838,N_6893);
and U7143 (N_7143,N_6973,N_6817);
or U7144 (N_7144,N_6950,N_6966);
and U7145 (N_7145,N_6851,N_6829);
or U7146 (N_7146,N_6936,N_6970);
nor U7147 (N_7147,N_6900,N_6945);
xnor U7148 (N_7148,N_6919,N_6834);
nor U7149 (N_7149,N_6963,N_6846);
nor U7150 (N_7150,N_6916,N_6913);
and U7151 (N_7151,N_6900,N_6805);
nand U7152 (N_7152,N_6907,N_6964);
and U7153 (N_7153,N_6835,N_6874);
and U7154 (N_7154,N_6827,N_6907);
and U7155 (N_7155,N_6907,N_6983);
and U7156 (N_7156,N_6858,N_6929);
and U7157 (N_7157,N_6925,N_6915);
nand U7158 (N_7158,N_6965,N_6820);
and U7159 (N_7159,N_6930,N_6908);
and U7160 (N_7160,N_6871,N_6931);
or U7161 (N_7161,N_6974,N_6894);
and U7162 (N_7162,N_6853,N_6818);
and U7163 (N_7163,N_6827,N_6851);
or U7164 (N_7164,N_6963,N_6803);
and U7165 (N_7165,N_6944,N_6810);
nand U7166 (N_7166,N_6830,N_6867);
or U7167 (N_7167,N_6970,N_6946);
or U7168 (N_7168,N_6806,N_6912);
nor U7169 (N_7169,N_6848,N_6988);
and U7170 (N_7170,N_6917,N_6943);
nor U7171 (N_7171,N_6899,N_6818);
or U7172 (N_7172,N_6886,N_6980);
xor U7173 (N_7173,N_6869,N_6903);
xnor U7174 (N_7174,N_6807,N_6857);
and U7175 (N_7175,N_6931,N_6908);
and U7176 (N_7176,N_6931,N_6950);
nand U7177 (N_7177,N_6952,N_6852);
nand U7178 (N_7178,N_6851,N_6891);
nor U7179 (N_7179,N_6966,N_6955);
or U7180 (N_7180,N_6951,N_6882);
nand U7181 (N_7181,N_6998,N_6892);
and U7182 (N_7182,N_6909,N_6905);
or U7183 (N_7183,N_6810,N_6877);
and U7184 (N_7184,N_6995,N_6851);
nor U7185 (N_7185,N_6847,N_6859);
nand U7186 (N_7186,N_6957,N_6839);
and U7187 (N_7187,N_6895,N_6857);
xnor U7188 (N_7188,N_6866,N_6959);
or U7189 (N_7189,N_6922,N_6827);
or U7190 (N_7190,N_6906,N_6844);
nand U7191 (N_7191,N_6860,N_6980);
and U7192 (N_7192,N_6878,N_6867);
and U7193 (N_7193,N_6923,N_6965);
nand U7194 (N_7194,N_6883,N_6859);
or U7195 (N_7195,N_6830,N_6947);
nand U7196 (N_7196,N_6905,N_6934);
xnor U7197 (N_7197,N_6960,N_6821);
and U7198 (N_7198,N_6893,N_6965);
nor U7199 (N_7199,N_6834,N_6827);
and U7200 (N_7200,N_7039,N_7099);
nand U7201 (N_7201,N_7050,N_7041);
nor U7202 (N_7202,N_7168,N_7080);
and U7203 (N_7203,N_7104,N_7137);
or U7204 (N_7204,N_7071,N_7062);
or U7205 (N_7205,N_7173,N_7154);
nor U7206 (N_7206,N_7183,N_7136);
and U7207 (N_7207,N_7112,N_7105);
and U7208 (N_7208,N_7189,N_7063);
xnor U7209 (N_7209,N_7198,N_7002);
and U7210 (N_7210,N_7019,N_7166);
nand U7211 (N_7211,N_7140,N_7188);
nand U7212 (N_7212,N_7171,N_7124);
and U7213 (N_7213,N_7159,N_7064);
nand U7214 (N_7214,N_7174,N_7008);
and U7215 (N_7215,N_7021,N_7123);
nor U7216 (N_7216,N_7161,N_7184);
nand U7217 (N_7217,N_7084,N_7135);
and U7218 (N_7218,N_7058,N_7165);
xnor U7219 (N_7219,N_7133,N_7069);
or U7220 (N_7220,N_7065,N_7079);
xor U7221 (N_7221,N_7155,N_7082);
nor U7222 (N_7222,N_7077,N_7072);
and U7223 (N_7223,N_7013,N_7005);
and U7224 (N_7224,N_7197,N_7196);
and U7225 (N_7225,N_7017,N_7193);
nand U7226 (N_7226,N_7126,N_7035);
nor U7227 (N_7227,N_7111,N_7045);
xnor U7228 (N_7228,N_7033,N_7040);
and U7229 (N_7229,N_7195,N_7102);
or U7230 (N_7230,N_7032,N_7175);
nand U7231 (N_7231,N_7185,N_7070);
nor U7232 (N_7232,N_7059,N_7088);
and U7233 (N_7233,N_7152,N_7034);
nand U7234 (N_7234,N_7110,N_7142);
xor U7235 (N_7235,N_7143,N_7087);
xor U7236 (N_7236,N_7003,N_7076);
nor U7237 (N_7237,N_7162,N_7117);
and U7238 (N_7238,N_7148,N_7127);
and U7239 (N_7239,N_7116,N_7144);
xnor U7240 (N_7240,N_7078,N_7053);
nand U7241 (N_7241,N_7038,N_7122);
nand U7242 (N_7242,N_7108,N_7051);
xor U7243 (N_7243,N_7007,N_7100);
nor U7244 (N_7244,N_7141,N_7001);
nor U7245 (N_7245,N_7181,N_7028);
or U7246 (N_7246,N_7075,N_7057);
or U7247 (N_7247,N_7056,N_7150);
xnor U7248 (N_7248,N_7132,N_7109);
and U7249 (N_7249,N_7129,N_7119);
nand U7250 (N_7250,N_7043,N_7097);
nand U7251 (N_7251,N_7199,N_7048);
and U7252 (N_7252,N_7020,N_7192);
nor U7253 (N_7253,N_7085,N_7176);
nor U7254 (N_7254,N_7115,N_7047);
and U7255 (N_7255,N_7016,N_7068);
or U7256 (N_7256,N_7054,N_7010);
nand U7257 (N_7257,N_7031,N_7096);
nand U7258 (N_7258,N_7178,N_7151);
nor U7259 (N_7259,N_7012,N_7046);
nand U7260 (N_7260,N_7000,N_7029);
nor U7261 (N_7261,N_7139,N_7042);
nor U7262 (N_7262,N_7023,N_7149);
nor U7263 (N_7263,N_7163,N_7146);
nand U7264 (N_7264,N_7004,N_7044);
nand U7265 (N_7265,N_7066,N_7106);
or U7266 (N_7266,N_7191,N_7052);
xnor U7267 (N_7267,N_7093,N_7113);
xor U7268 (N_7268,N_7026,N_7103);
nand U7269 (N_7269,N_7067,N_7153);
or U7270 (N_7270,N_7055,N_7081);
nand U7271 (N_7271,N_7011,N_7130);
nand U7272 (N_7272,N_7134,N_7179);
or U7273 (N_7273,N_7091,N_7015);
or U7274 (N_7274,N_7180,N_7121);
and U7275 (N_7275,N_7095,N_7169);
and U7276 (N_7276,N_7086,N_7018);
nor U7277 (N_7277,N_7118,N_7092);
or U7278 (N_7278,N_7160,N_7025);
nand U7279 (N_7279,N_7061,N_7138);
and U7280 (N_7280,N_7172,N_7120);
and U7281 (N_7281,N_7145,N_7157);
nand U7282 (N_7282,N_7101,N_7125);
nand U7283 (N_7283,N_7037,N_7030);
and U7284 (N_7284,N_7107,N_7190);
nor U7285 (N_7285,N_7170,N_7158);
xnor U7286 (N_7286,N_7114,N_7186);
or U7287 (N_7287,N_7036,N_7131);
xor U7288 (N_7288,N_7027,N_7194);
or U7289 (N_7289,N_7182,N_7156);
and U7290 (N_7290,N_7089,N_7177);
and U7291 (N_7291,N_7164,N_7022);
or U7292 (N_7292,N_7009,N_7098);
or U7293 (N_7293,N_7090,N_7060);
or U7294 (N_7294,N_7128,N_7167);
xnor U7295 (N_7295,N_7074,N_7049);
or U7296 (N_7296,N_7147,N_7006);
nand U7297 (N_7297,N_7024,N_7014);
and U7298 (N_7298,N_7187,N_7073);
and U7299 (N_7299,N_7083,N_7094);
or U7300 (N_7300,N_7124,N_7170);
or U7301 (N_7301,N_7194,N_7145);
xor U7302 (N_7302,N_7115,N_7096);
and U7303 (N_7303,N_7107,N_7069);
or U7304 (N_7304,N_7170,N_7155);
or U7305 (N_7305,N_7126,N_7002);
nor U7306 (N_7306,N_7034,N_7070);
nor U7307 (N_7307,N_7196,N_7165);
nor U7308 (N_7308,N_7133,N_7181);
nor U7309 (N_7309,N_7194,N_7193);
nand U7310 (N_7310,N_7043,N_7199);
or U7311 (N_7311,N_7099,N_7158);
nand U7312 (N_7312,N_7186,N_7154);
or U7313 (N_7313,N_7026,N_7174);
and U7314 (N_7314,N_7130,N_7197);
or U7315 (N_7315,N_7192,N_7029);
and U7316 (N_7316,N_7130,N_7147);
and U7317 (N_7317,N_7006,N_7165);
nand U7318 (N_7318,N_7155,N_7135);
or U7319 (N_7319,N_7065,N_7082);
and U7320 (N_7320,N_7131,N_7181);
nand U7321 (N_7321,N_7032,N_7054);
nor U7322 (N_7322,N_7047,N_7033);
nor U7323 (N_7323,N_7055,N_7126);
and U7324 (N_7324,N_7013,N_7012);
xor U7325 (N_7325,N_7086,N_7182);
xnor U7326 (N_7326,N_7108,N_7085);
nor U7327 (N_7327,N_7052,N_7082);
nor U7328 (N_7328,N_7120,N_7013);
or U7329 (N_7329,N_7018,N_7058);
xnor U7330 (N_7330,N_7019,N_7043);
xor U7331 (N_7331,N_7089,N_7134);
xnor U7332 (N_7332,N_7175,N_7064);
nor U7333 (N_7333,N_7091,N_7150);
xnor U7334 (N_7334,N_7040,N_7044);
and U7335 (N_7335,N_7192,N_7006);
and U7336 (N_7336,N_7186,N_7032);
nor U7337 (N_7337,N_7082,N_7159);
nand U7338 (N_7338,N_7194,N_7191);
or U7339 (N_7339,N_7023,N_7108);
and U7340 (N_7340,N_7115,N_7182);
nand U7341 (N_7341,N_7033,N_7012);
nor U7342 (N_7342,N_7126,N_7104);
nor U7343 (N_7343,N_7070,N_7063);
and U7344 (N_7344,N_7105,N_7171);
and U7345 (N_7345,N_7186,N_7001);
nand U7346 (N_7346,N_7106,N_7199);
and U7347 (N_7347,N_7083,N_7080);
or U7348 (N_7348,N_7027,N_7000);
nand U7349 (N_7349,N_7096,N_7125);
and U7350 (N_7350,N_7165,N_7007);
and U7351 (N_7351,N_7148,N_7034);
nor U7352 (N_7352,N_7039,N_7078);
nor U7353 (N_7353,N_7181,N_7117);
nand U7354 (N_7354,N_7177,N_7112);
xnor U7355 (N_7355,N_7093,N_7162);
and U7356 (N_7356,N_7099,N_7066);
or U7357 (N_7357,N_7018,N_7168);
nor U7358 (N_7358,N_7121,N_7194);
or U7359 (N_7359,N_7159,N_7011);
nor U7360 (N_7360,N_7003,N_7116);
and U7361 (N_7361,N_7153,N_7085);
or U7362 (N_7362,N_7002,N_7032);
or U7363 (N_7363,N_7067,N_7151);
or U7364 (N_7364,N_7053,N_7007);
and U7365 (N_7365,N_7115,N_7093);
or U7366 (N_7366,N_7093,N_7154);
or U7367 (N_7367,N_7017,N_7114);
xnor U7368 (N_7368,N_7042,N_7101);
nand U7369 (N_7369,N_7044,N_7160);
or U7370 (N_7370,N_7188,N_7020);
and U7371 (N_7371,N_7174,N_7132);
or U7372 (N_7372,N_7129,N_7052);
xnor U7373 (N_7373,N_7195,N_7070);
or U7374 (N_7374,N_7064,N_7018);
xnor U7375 (N_7375,N_7140,N_7105);
xnor U7376 (N_7376,N_7178,N_7060);
or U7377 (N_7377,N_7103,N_7105);
nor U7378 (N_7378,N_7185,N_7157);
and U7379 (N_7379,N_7053,N_7065);
nor U7380 (N_7380,N_7013,N_7043);
nor U7381 (N_7381,N_7033,N_7128);
xnor U7382 (N_7382,N_7169,N_7092);
nor U7383 (N_7383,N_7049,N_7001);
nand U7384 (N_7384,N_7186,N_7195);
nand U7385 (N_7385,N_7175,N_7136);
nor U7386 (N_7386,N_7066,N_7034);
or U7387 (N_7387,N_7027,N_7099);
nor U7388 (N_7388,N_7186,N_7113);
nand U7389 (N_7389,N_7029,N_7083);
and U7390 (N_7390,N_7167,N_7161);
nand U7391 (N_7391,N_7097,N_7044);
xor U7392 (N_7392,N_7121,N_7009);
nor U7393 (N_7393,N_7115,N_7169);
nor U7394 (N_7394,N_7176,N_7020);
nor U7395 (N_7395,N_7193,N_7027);
nor U7396 (N_7396,N_7111,N_7041);
nand U7397 (N_7397,N_7163,N_7016);
and U7398 (N_7398,N_7075,N_7012);
or U7399 (N_7399,N_7072,N_7099);
nand U7400 (N_7400,N_7311,N_7352);
nor U7401 (N_7401,N_7222,N_7378);
nand U7402 (N_7402,N_7323,N_7347);
or U7403 (N_7403,N_7253,N_7343);
and U7404 (N_7404,N_7289,N_7217);
nor U7405 (N_7405,N_7228,N_7300);
nand U7406 (N_7406,N_7208,N_7361);
nor U7407 (N_7407,N_7335,N_7234);
and U7408 (N_7408,N_7390,N_7342);
or U7409 (N_7409,N_7237,N_7202);
and U7410 (N_7410,N_7367,N_7374);
nor U7411 (N_7411,N_7230,N_7272);
or U7412 (N_7412,N_7357,N_7287);
or U7413 (N_7413,N_7284,N_7246);
or U7414 (N_7414,N_7364,N_7298);
nand U7415 (N_7415,N_7281,N_7394);
and U7416 (N_7416,N_7391,N_7212);
nor U7417 (N_7417,N_7250,N_7306);
and U7418 (N_7418,N_7243,N_7326);
nor U7419 (N_7419,N_7249,N_7375);
nand U7420 (N_7420,N_7227,N_7322);
or U7421 (N_7421,N_7276,N_7240);
and U7422 (N_7422,N_7207,N_7239);
nand U7423 (N_7423,N_7201,N_7291);
nand U7424 (N_7424,N_7381,N_7305);
nand U7425 (N_7425,N_7385,N_7331);
or U7426 (N_7426,N_7204,N_7302);
and U7427 (N_7427,N_7319,N_7387);
nor U7428 (N_7428,N_7315,N_7282);
xnor U7429 (N_7429,N_7362,N_7244);
or U7430 (N_7430,N_7236,N_7330);
and U7431 (N_7431,N_7274,N_7370);
nor U7432 (N_7432,N_7273,N_7225);
nor U7433 (N_7433,N_7332,N_7206);
nand U7434 (N_7434,N_7268,N_7238);
and U7435 (N_7435,N_7368,N_7383);
nor U7436 (N_7436,N_7256,N_7221);
nand U7437 (N_7437,N_7382,N_7345);
nor U7438 (N_7438,N_7211,N_7355);
nor U7439 (N_7439,N_7363,N_7340);
or U7440 (N_7440,N_7336,N_7371);
and U7441 (N_7441,N_7266,N_7214);
nor U7442 (N_7442,N_7393,N_7231);
or U7443 (N_7443,N_7325,N_7349);
nand U7444 (N_7444,N_7351,N_7205);
and U7445 (N_7445,N_7280,N_7252);
and U7446 (N_7446,N_7318,N_7337);
and U7447 (N_7447,N_7279,N_7218);
nand U7448 (N_7448,N_7223,N_7308);
and U7449 (N_7449,N_7307,N_7210);
nor U7450 (N_7450,N_7369,N_7278);
and U7451 (N_7451,N_7219,N_7270);
and U7452 (N_7452,N_7312,N_7296);
and U7453 (N_7453,N_7262,N_7327);
and U7454 (N_7454,N_7313,N_7377);
xor U7455 (N_7455,N_7215,N_7386);
and U7456 (N_7456,N_7299,N_7290);
nand U7457 (N_7457,N_7293,N_7294);
or U7458 (N_7458,N_7372,N_7285);
xor U7459 (N_7459,N_7261,N_7286);
nand U7460 (N_7460,N_7288,N_7258);
or U7461 (N_7461,N_7283,N_7264);
nand U7462 (N_7462,N_7257,N_7310);
and U7463 (N_7463,N_7247,N_7398);
nor U7464 (N_7464,N_7229,N_7324);
and U7465 (N_7465,N_7346,N_7316);
xor U7466 (N_7466,N_7353,N_7203);
or U7467 (N_7467,N_7209,N_7328);
and U7468 (N_7468,N_7303,N_7348);
xor U7469 (N_7469,N_7267,N_7226);
or U7470 (N_7470,N_7373,N_7317);
nor U7471 (N_7471,N_7366,N_7338);
nand U7472 (N_7472,N_7339,N_7224);
or U7473 (N_7473,N_7301,N_7251);
nor U7474 (N_7474,N_7333,N_7356);
nor U7475 (N_7475,N_7396,N_7245);
nand U7476 (N_7476,N_7309,N_7265);
nor U7477 (N_7477,N_7376,N_7392);
and U7478 (N_7478,N_7379,N_7232);
nand U7479 (N_7479,N_7216,N_7213);
and U7480 (N_7480,N_7277,N_7220);
xor U7481 (N_7481,N_7388,N_7397);
or U7482 (N_7482,N_7314,N_7359);
or U7483 (N_7483,N_7384,N_7304);
xnor U7484 (N_7484,N_7395,N_7235);
or U7485 (N_7485,N_7329,N_7358);
xnor U7486 (N_7486,N_7233,N_7271);
and U7487 (N_7487,N_7297,N_7295);
nand U7488 (N_7488,N_7344,N_7320);
or U7489 (N_7489,N_7248,N_7399);
or U7490 (N_7490,N_7360,N_7350);
or U7491 (N_7491,N_7259,N_7254);
nand U7492 (N_7492,N_7200,N_7275);
nand U7493 (N_7493,N_7241,N_7260);
or U7494 (N_7494,N_7269,N_7365);
and U7495 (N_7495,N_7380,N_7389);
nand U7496 (N_7496,N_7242,N_7334);
or U7497 (N_7497,N_7341,N_7263);
or U7498 (N_7498,N_7292,N_7255);
nand U7499 (N_7499,N_7354,N_7321);
and U7500 (N_7500,N_7211,N_7206);
and U7501 (N_7501,N_7223,N_7378);
or U7502 (N_7502,N_7381,N_7295);
nor U7503 (N_7503,N_7366,N_7312);
nor U7504 (N_7504,N_7378,N_7339);
nor U7505 (N_7505,N_7340,N_7217);
nand U7506 (N_7506,N_7236,N_7362);
or U7507 (N_7507,N_7368,N_7278);
nor U7508 (N_7508,N_7332,N_7262);
nor U7509 (N_7509,N_7312,N_7284);
nor U7510 (N_7510,N_7219,N_7232);
and U7511 (N_7511,N_7280,N_7393);
nand U7512 (N_7512,N_7238,N_7243);
and U7513 (N_7513,N_7265,N_7357);
nand U7514 (N_7514,N_7283,N_7398);
or U7515 (N_7515,N_7397,N_7362);
and U7516 (N_7516,N_7303,N_7235);
and U7517 (N_7517,N_7338,N_7313);
or U7518 (N_7518,N_7226,N_7364);
xnor U7519 (N_7519,N_7253,N_7304);
or U7520 (N_7520,N_7295,N_7268);
nor U7521 (N_7521,N_7331,N_7375);
or U7522 (N_7522,N_7247,N_7267);
or U7523 (N_7523,N_7335,N_7319);
and U7524 (N_7524,N_7206,N_7380);
and U7525 (N_7525,N_7311,N_7340);
nor U7526 (N_7526,N_7241,N_7259);
and U7527 (N_7527,N_7372,N_7248);
nand U7528 (N_7528,N_7233,N_7250);
xnor U7529 (N_7529,N_7279,N_7243);
or U7530 (N_7530,N_7204,N_7234);
or U7531 (N_7531,N_7343,N_7379);
nand U7532 (N_7532,N_7306,N_7375);
xor U7533 (N_7533,N_7399,N_7257);
nor U7534 (N_7534,N_7351,N_7261);
and U7535 (N_7535,N_7224,N_7387);
or U7536 (N_7536,N_7312,N_7287);
and U7537 (N_7537,N_7259,N_7396);
and U7538 (N_7538,N_7383,N_7372);
and U7539 (N_7539,N_7256,N_7236);
nor U7540 (N_7540,N_7233,N_7321);
nor U7541 (N_7541,N_7394,N_7375);
xnor U7542 (N_7542,N_7228,N_7338);
and U7543 (N_7543,N_7354,N_7377);
and U7544 (N_7544,N_7320,N_7309);
nand U7545 (N_7545,N_7209,N_7244);
and U7546 (N_7546,N_7398,N_7319);
nand U7547 (N_7547,N_7322,N_7205);
nand U7548 (N_7548,N_7383,N_7381);
nor U7549 (N_7549,N_7339,N_7370);
nand U7550 (N_7550,N_7209,N_7384);
and U7551 (N_7551,N_7311,N_7312);
nor U7552 (N_7552,N_7330,N_7256);
nor U7553 (N_7553,N_7303,N_7298);
nor U7554 (N_7554,N_7349,N_7355);
nor U7555 (N_7555,N_7265,N_7379);
or U7556 (N_7556,N_7372,N_7317);
or U7557 (N_7557,N_7388,N_7228);
and U7558 (N_7558,N_7361,N_7231);
and U7559 (N_7559,N_7345,N_7338);
nand U7560 (N_7560,N_7232,N_7278);
and U7561 (N_7561,N_7237,N_7243);
nand U7562 (N_7562,N_7219,N_7298);
nor U7563 (N_7563,N_7384,N_7303);
nand U7564 (N_7564,N_7394,N_7338);
nor U7565 (N_7565,N_7254,N_7332);
xnor U7566 (N_7566,N_7298,N_7315);
nand U7567 (N_7567,N_7381,N_7320);
nor U7568 (N_7568,N_7265,N_7361);
nand U7569 (N_7569,N_7309,N_7230);
and U7570 (N_7570,N_7309,N_7324);
nand U7571 (N_7571,N_7210,N_7359);
nor U7572 (N_7572,N_7217,N_7387);
or U7573 (N_7573,N_7217,N_7366);
nand U7574 (N_7574,N_7269,N_7354);
or U7575 (N_7575,N_7348,N_7239);
nand U7576 (N_7576,N_7312,N_7352);
or U7577 (N_7577,N_7390,N_7204);
nor U7578 (N_7578,N_7280,N_7354);
and U7579 (N_7579,N_7279,N_7213);
nor U7580 (N_7580,N_7302,N_7228);
or U7581 (N_7581,N_7276,N_7381);
or U7582 (N_7582,N_7239,N_7211);
nor U7583 (N_7583,N_7339,N_7318);
and U7584 (N_7584,N_7327,N_7215);
nand U7585 (N_7585,N_7249,N_7293);
or U7586 (N_7586,N_7214,N_7236);
nor U7587 (N_7587,N_7377,N_7351);
nor U7588 (N_7588,N_7293,N_7218);
nand U7589 (N_7589,N_7331,N_7277);
xnor U7590 (N_7590,N_7294,N_7259);
or U7591 (N_7591,N_7399,N_7266);
xnor U7592 (N_7592,N_7320,N_7354);
and U7593 (N_7593,N_7249,N_7357);
nand U7594 (N_7594,N_7342,N_7349);
or U7595 (N_7595,N_7340,N_7222);
nor U7596 (N_7596,N_7257,N_7248);
and U7597 (N_7597,N_7376,N_7319);
nand U7598 (N_7598,N_7264,N_7359);
and U7599 (N_7599,N_7266,N_7235);
nand U7600 (N_7600,N_7491,N_7417);
or U7601 (N_7601,N_7535,N_7516);
or U7602 (N_7602,N_7507,N_7482);
or U7603 (N_7603,N_7408,N_7499);
or U7604 (N_7604,N_7532,N_7496);
and U7605 (N_7605,N_7477,N_7416);
nor U7606 (N_7606,N_7591,N_7407);
or U7607 (N_7607,N_7471,N_7510);
and U7608 (N_7608,N_7534,N_7530);
nor U7609 (N_7609,N_7572,N_7587);
nor U7610 (N_7610,N_7564,N_7444);
nor U7611 (N_7611,N_7409,N_7431);
and U7612 (N_7612,N_7460,N_7522);
and U7613 (N_7613,N_7415,N_7552);
nand U7614 (N_7614,N_7536,N_7548);
nand U7615 (N_7615,N_7590,N_7437);
nor U7616 (N_7616,N_7423,N_7419);
or U7617 (N_7617,N_7553,N_7571);
nand U7618 (N_7618,N_7412,N_7595);
nor U7619 (N_7619,N_7574,N_7438);
nand U7620 (N_7620,N_7489,N_7449);
or U7621 (N_7621,N_7483,N_7425);
and U7622 (N_7622,N_7546,N_7511);
xnor U7623 (N_7623,N_7525,N_7433);
and U7624 (N_7624,N_7578,N_7569);
or U7625 (N_7625,N_7582,N_7476);
and U7626 (N_7626,N_7478,N_7599);
nor U7627 (N_7627,N_7426,N_7420);
and U7628 (N_7628,N_7579,N_7461);
and U7629 (N_7629,N_7442,N_7586);
nand U7630 (N_7630,N_7446,N_7422);
and U7631 (N_7631,N_7594,N_7492);
nand U7632 (N_7632,N_7459,N_7480);
nor U7633 (N_7633,N_7580,N_7429);
and U7634 (N_7634,N_7593,N_7598);
nand U7635 (N_7635,N_7528,N_7573);
xor U7636 (N_7636,N_7404,N_7568);
nor U7637 (N_7637,N_7421,N_7521);
or U7638 (N_7638,N_7577,N_7531);
nand U7639 (N_7639,N_7443,N_7466);
or U7640 (N_7640,N_7497,N_7515);
nand U7641 (N_7641,N_7440,N_7427);
nand U7642 (N_7642,N_7547,N_7456);
nand U7643 (N_7643,N_7462,N_7524);
nor U7644 (N_7644,N_7540,N_7469);
nand U7645 (N_7645,N_7596,N_7495);
nor U7646 (N_7646,N_7555,N_7479);
and U7647 (N_7647,N_7463,N_7502);
nor U7648 (N_7648,N_7558,N_7490);
or U7649 (N_7649,N_7411,N_7434);
nor U7650 (N_7650,N_7567,N_7498);
xor U7651 (N_7651,N_7418,N_7472);
nand U7652 (N_7652,N_7550,N_7509);
nand U7653 (N_7653,N_7470,N_7545);
nor U7654 (N_7654,N_7454,N_7430);
xnor U7655 (N_7655,N_7445,N_7556);
nand U7656 (N_7656,N_7468,N_7533);
and U7657 (N_7657,N_7520,N_7441);
nor U7658 (N_7658,N_7453,N_7537);
or U7659 (N_7659,N_7543,N_7424);
nor U7660 (N_7660,N_7538,N_7506);
or U7661 (N_7661,N_7589,N_7455);
or U7662 (N_7662,N_7542,N_7505);
nand U7663 (N_7663,N_7436,N_7405);
nand U7664 (N_7664,N_7467,N_7485);
and U7665 (N_7665,N_7583,N_7557);
or U7666 (N_7666,N_7501,N_7475);
xor U7667 (N_7667,N_7403,N_7435);
or U7668 (N_7668,N_7512,N_7519);
nand U7669 (N_7669,N_7481,N_7488);
and U7670 (N_7670,N_7585,N_7554);
nor U7671 (N_7671,N_7562,N_7432);
and U7672 (N_7672,N_7575,N_7513);
nor U7673 (N_7673,N_7500,N_7563);
or U7674 (N_7674,N_7518,N_7400);
xor U7675 (N_7675,N_7551,N_7504);
xor U7676 (N_7676,N_7451,N_7570);
xnor U7677 (N_7677,N_7526,N_7517);
nor U7678 (N_7678,N_7549,N_7401);
and U7679 (N_7679,N_7588,N_7487);
nand U7680 (N_7680,N_7565,N_7452);
and U7681 (N_7681,N_7402,N_7561);
or U7682 (N_7682,N_7597,N_7406);
nor U7683 (N_7683,N_7503,N_7474);
nand U7684 (N_7684,N_7539,N_7450);
nor U7685 (N_7685,N_7523,N_7428);
nor U7686 (N_7686,N_7457,N_7448);
nand U7687 (N_7687,N_7414,N_7581);
nand U7688 (N_7688,N_7566,N_7576);
or U7689 (N_7689,N_7413,N_7486);
xnor U7690 (N_7690,N_7410,N_7560);
nand U7691 (N_7691,N_7584,N_7458);
xor U7692 (N_7692,N_7541,N_7439);
nor U7693 (N_7693,N_7494,N_7465);
nor U7694 (N_7694,N_7544,N_7514);
nor U7695 (N_7695,N_7493,N_7508);
or U7696 (N_7696,N_7559,N_7464);
nor U7697 (N_7697,N_7592,N_7527);
and U7698 (N_7698,N_7529,N_7484);
nor U7699 (N_7699,N_7473,N_7447);
nand U7700 (N_7700,N_7571,N_7541);
and U7701 (N_7701,N_7583,N_7478);
and U7702 (N_7702,N_7538,N_7499);
xnor U7703 (N_7703,N_7516,N_7439);
or U7704 (N_7704,N_7420,N_7549);
nand U7705 (N_7705,N_7403,N_7468);
and U7706 (N_7706,N_7477,N_7546);
nor U7707 (N_7707,N_7471,N_7560);
or U7708 (N_7708,N_7596,N_7401);
xnor U7709 (N_7709,N_7589,N_7463);
or U7710 (N_7710,N_7569,N_7494);
nor U7711 (N_7711,N_7405,N_7525);
nor U7712 (N_7712,N_7537,N_7477);
or U7713 (N_7713,N_7475,N_7571);
nand U7714 (N_7714,N_7427,N_7581);
and U7715 (N_7715,N_7561,N_7464);
and U7716 (N_7716,N_7551,N_7430);
nand U7717 (N_7717,N_7404,N_7423);
or U7718 (N_7718,N_7459,N_7451);
or U7719 (N_7719,N_7484,N_7480);
nor U7720 (N_7720,N_7418,N_7434);
nor U7721 (N_7721,N_7425,N_7417);
nand U7722 (N_7722,N_7550,N_7438);
and U7723 (N_7723,N_7467,N_7446);
or U7724 (N_7724,N_7439,N_7492);
nand U7725 (N_7725,N_7460,N_7566);
or U7726 (N_7726,N_7408,N_7532);
nand U7727 (N_7727,N_7493,N_7448);
or U7728 (N_7728,N_7559,N_7588);
and U7729 (N_7729,N_7588,N_7581);
nand U7730 (N_7730,N_7550,N_7421);
nand U7731 (N_7731,N_7577,N_7579);
nand U7732 (N_7732,N_7433,N_7421);
nor U7733 (N_7733,N_7467,N_7576);
and U7734 (N_7734,N_7434,N_7429);
or U7735 (N_7735,N_7584,N_7429);
nand U7736 (N_7736,N_7590,N_7430);
nor U7737 (N_7737,N_7531,N_7466);
nor U7738 (N_7738,N_7540,N_7410);
nand U7739 (N_7739,N_7492,N_7479);
nor U7740 (N_7740,N_7569,N_7472);
nand U7741 (N_7741,N_7594,N_7476);
nor U7742 (N_7742,N_7498,N_7565);
nand U7743 (N_7743,N_7444,N_7400);
and U7744 (N_7744,N_7443,N_7405);
or U7745 (N_7745,N_7565,N_7592);
and U7746 (N_7746,N_7459,N_7516);
and U7747 (N_7747,N_7567,N_7464);
nand U7748 (N_7748,N_7402,N_7599);
and U7749 (N_7749,N_7555,N_7403);
xnor U7750 (N_7750,N_7550,N_7485);
nor U7751 (N_7751,N_7542,N_7507);
xor U7752 (N_7752,N_7460,N_7532);
or U7753 (N_7753,N_7570,N_7430);
nor U7754 (N_7754,N_7523,N_7488);
xnor U7755 (N_7755,N_7532,N_7577);
nor U7756 (N_7756,N_7527,N_7505);
nor U7757 (N_7757,N_7473,N_7538);
nand U7758 (N_7758,N_7478,N_7514);
and U7759 (N_7759,N_7500,N_7531);
xnor U7760 (N_7760,N_7526,N_7515);
and U7761 (N_7761,N_7598,N_7525);
or U7762 (N_7762,N_7416,N_7491);
or U7763 (N_7763,N_7405,N_7481);
and U7764 (N_7764,N_7586,N_7439);
or U7765 (N_7765,N_7447,N_7565);
nand U7766 (N_7766,N_7409,N_7483);
nand U7767 (N_7767,N_7447,N_7480);
nor U7768 (N_7768,N_7512,N_7423);
and U7769 (N_7769,N_7448,N_7573);
or U7770 (N_7770,N_7458,N_7405);
nor U7771 (N_7771,N_7566,N_7578);
and U7772 (N_7772,N_7504,N_7407);
nor U7773 (N_7773,N_7479,N_7589);
and U7774 (N_7774,N_7407,N_7455);
nand U7775 (N_7775,N_7481,N_7445);
and U7776 (N_7776,N_7437,N_7430);
nand U7777 (N_7777,N_7488,N_7557);
nand U7778 (N_7778,N_7555,N_7581);
nand U7779 (N_7779,N_7467,N_7529);
nand U7780 (N_7780,N_7447,N_7577);
and U7781 (N_7781,N_7403,N_7574);
and U7782 (N_7782,N_7478,N_7579);
nor U7783 (N_7783,N_7570,N_7404);
or U7784 (N_7784,N_7528,N_7561);
nor U7785 (N_7785,N_7578,N_7542);
or U7786 (N_7786,N_7472,N_7470);
and U7787 (N_7787,N_7570,N_7418);
or U7788 (N_7788,N_7476,N_7529);
and U7789 (N_7789,N_7558,N_7492);
nand U7790 (N_7790,N_7418,N_7432);
nand U7791 (N_7791,N_7536,N_7490);
nand U7792 (N_7792,N_7488,N_7474);
nor U7793 (N_7793,N_7529,N_7434);
or U7794 (N_7794,N_7596,N_7567);
or U7795 (N_7795,N_7503,N_7576);
xor U7796 (N_7796,N_7587,N_7534);
nor U7797 (N_7797,N_7495,N_7430);
nand U7798 (N_7798,N_7477,N_7583);
and U7799 (N_7799,N_7481,N_7587);
nor U7800 (N_7800,N_7631,N_7738);
or U7801 (N_7801,N_7726,N_7785);
nand U7802 (N_7802,N_7696,N_7725);
and U7803 (N_7803,N_7727,N_7660);
or U7804 (N_7804,N_7734,N_7645);
and U7805 (N_7805,N_7736,N_7789);
or U7806 (N_7806,N_7667,N_7761);
nor U7807 (N_7807,N_7677,N_7757);
or U7808 (N_7808,N_7614,N_7796);
or U7809 (N_7809,N_7740,N_7708);
and U7810 (N_7810,N_7753,N_7712);
nor U7811 (N_7811,N_7601,N_7648);
nor U7812 (N_7812,N_7747,N_7735);
and U7813 (N_7813,N_7793,N_7767);
or U7814 (N_7814,N_7602,N_7625);
nand U7815 (N_7815,N_7675,N_7633);
or U7816 (N_7816,N_7632,N_7629);
nor U7817 (N_7817,N_7728,N_7687);
nor U7818 (N_7818,N_7713,N_7788);
nand U7819 (N_7819,N_7673,N_7746);
nand U7820 (N_7820,N_7719,N_7697);
and U7821 (N_7821,N_7775,N_7754);
nor U7822 (N_7822,N_7654,N_7661);
nor U7823 (N_7823,N_7665,N_7776);
nand U7824 (N_7824,N_7662,N_7755);
nand U7825 (N_7825,N_7618,N_7639);
and U7826 (N_7826,N_7682,N_7756);
xnor U7827 (N_7827,N_7739,N_7603);
and U7828 (N_7828,N_7615,N_7798);
nor U7829 (N_7829,N_7792,N_7650);
and U7830 (N_7830,N_7640,N_7758);
and U7831 (N_7831,N_7764,N_7616);
or U7832 (N_7832,N_7600,N_7611);
or U7833 (N_7833,N_7759,N_7745);
xnor U7834 (N_7834,N_7765,N_7636);
nand U7835 (N_7835,N_7679,N_7670);
and U7836 (N_7836,N_7676,N_7609);
or U7837 (N_7837,N_7794,N_7684);
and U7838 (N_7838,N_7718,N_7612);
nand U7839 (N_7839,N_7643,N_7686);
nand U7840 (N_7840,N_7628,N_7622);
nor U7841 (N_7841,N_7651,N_7674);
nor U7842 (N_7842,N_7790,N_7781);
xnor U7843 (N_7843,N_7724,N_7710);
and U7844 (N_7844,N_7627,N_7637);
nor U7845 (N_7845,N_7689,N_7613);
and U7846 (N_7846,N_7700,N_7610);
nand U7847 (N_7847,N_7642,N_7774);
and U7848 (N_7848,N_7644,N_7678);
and U7849 (N_7849,N_7683,N_7690);
and U7850 (N_7850,N_7604,N_7751);
nor U7851 (N_7851,N_7709,N_7723);
and U7852 (N_7852,N_7659,N_7799);
xor U7853 (N_7853,N_7702,N_7634);
or U7854 (N_7854,N_7707,N_7742);
nand U7855 (N_7855,N_7763,N_7646);
and U7856 (N_7856,N_7624,N_7655);
or U7857 (N_7857,N_7783,N_7626);
or U7858 (N_7858,N_7685,N_7649);
nand U7859 (N_7859,N_7704,N_7772);
and U7860 (N_7860,N_7779,N_7656);
xnor U7861 (N_7861,N_7787,N_7671);
xor U7862 (N_7862,N_7717,N_7630);
nor U7863 (N_7863,N_7750,N_7743);
nor U7864 (N_7864,N_7608,N_7784);
nor U7865 (N_7865,N_7606,N_7623);
nor U7866 (N_7866,N_7762,N_7770);
nand U7867 (N_7867,N_7777,N_7732);
nand U7868 (N_7868,N_7795,N_7769);
nor U7869 (N_7869,N_7692,N_7744);
and U7870 (N_7870,N_7619,N_7635);
or U7871 (N_7871,N_7731,N_7714);
nor U7872 (N_7872,N_7720,N_7658);
or U7873 (N_7873,N_7669,N_7711);
nor U7874 (N_7874,N_7733,N_7730);
or U7875 (N_7875,N_7647,N_7703);
xnor U7876 (N_7876,N_7771,N_7638);
or U7877 (N_7877,N_7672,N_7782);
and U7878 (N_7878,N_7653,N_7791);
or U7879 (N_7879,N_7699,N_7701);
and U7880 (N_7880,N_7780,N_7688);
nor U7881 (N_7881,N_7748,N_7716);
and U7882 (N_7882,N_7786,N_7749);
or U7883 (N_7883,N_7668,N_7705);
nor U7884 (N_7884,N_7681,N_7657);
and U7885 (N_7885,N_7760,N_7715);
or U7886 (N_7886,N_7693,N_7617);
and U7887 (N_7887,N_7605,N_7694);
and U7888 (N_7888,N_7621,N_7691);
nand U7889 (N_7889,N_7620,N_7680);
nor U7890 (N_7890,N_7773,N_7752);
and U7891 (N_7891,N_7641,N_7698);
nand U7892 (N_7892,N_7797,N_7778);
nor U7893 (N_7893,N_7695,N_7721);
nand U7894 (N_7894,N_7722,N_7729);
and U7895 (N_7895,N_7766,N_7768);
and U7896 (N_7896,N_7664,N_7666);
nand U7897 (N_7897,N_7706,N_7663);
or U7898 (N_7898,N_7607,N_7741);
nor U7899 (N_7899,N_7737,N_7652);
or U7900 (N_7900,N_7797,N_7603);
nor U7901 (N_7901,N_7769,N_7618);
nor U7902 (N_7902,N_7638,N_7608);
nor U7903 (N_7903,N_7694,N_7674);
nor U7904 (N_7904,N_7668,N_7617);
and U7905 (N_7905,N_7644,N_7634);
xor U7906 (N_7906,N_7743,N_7670);
xor U7907 (N_7907,N_7796,N_7625);
nand U7908 (N_7908,N_7677,N_7717);
and U7909 (N_7909,N_7700,N_7614);
and U7910 (N_7910,N_7601,N_7791);
nor U7911 (N_7911,N_7770,N_7600);
nor U7912 (N_7912,N_7747,N_7682);
nor U7913 (N_7913,N_7709,N_7657);
and U7914 (N_7914,N_7634,N_7739);
or U7915 (N_7915,N_7786,N_7628);
and U7916 (N_7916,N_7732,N_7617);
or U7917 (N_7917,N_7642,N_7672);
or U7918 (N_7918,N_7756,N_7794);
nor U7919 (N_7919,N_7703,N_7628);
or U7920 (N_7920,N_7623,N_7680);
or U7921 (N_7921,N_7756,N_7745);
and U7922 (N_7922,N_7680,N_7671);
nand U7923 (N_7923,N_7694,N_7757);
or U7924 (N_7924,N_7799,N_7634);
nand U7925 (N_7925,N_7601,N_7715);
or U7926 (N_7926,N_7709,N_7600);
nand U7927 (N_7927,N_7671,N_7664);
nor U7928 (N_7928,N_7620,N_7774);
and U7929 (N_7929,N_7797,N_7751);
nand U7930 (N_7930,N_7786,N_7753);
and U7931 (N_7931,N_7626,N_7704);
nand U7932 (N_7932,N_7652,N_7747);
xnor U7933 (N_7933,N_7689,N_7675);
xnor U7934 (N_7934,N_7697,N_7691);
and U7935 (N_7935,N_7600,N_7701);
nand U7936 (N_7936,N_7716,N_7799);
nor U7937 (N_7937,N_7743,N_7739);
nor U7938 (N_7938,N_7708,N_7629);
and U7939 (N_7939,N_7774,N_7672);
nor U7940 (N_7940,N_7779,N_7706);
xor U7941 (N_7941,N_7683,N_7783);
xor U7942 (N_7942,N_7604,N_7712);
and U7943 (N_7943,N_7658,N_7772);
nor U7944 (N_7944,N_7711,N_7639);
or U7945 (N_7945,N_7612,N_7762);
or U7946 (N_7946,N_7744,N_7742);
and U7947 (N_7947,N_7671,N_7741);
or U7948 (N_7948,N_7782,N_7748);
and U7949 (N_7949,N_7685,N_7624);
and U7950 (N_7950,N_7606,N_7776);
and U7951 (N_7951,N_7648,N_7627);
and U7952 (N_7952,N_7745,N_7640);
nor U7953 (N_7953,N_7698,N_7770);
nor U7954 (N_7954,N_7783,N_7771);
nor U7955 (N_7955,N_7698,N_7645);
nor U7956 (N_7956,N_7754,N_7683);
and U7957 (N_7957,N_7766,N_7634);
nand U7958 (N_7958,N_7630,N_7618);
or U7959 (N_7959,N_7794,N_7662);
nand U7960 (N_7960,N_7779,N_7727);
or U7961 (N_7961,N_7796,N_7635);
nand U7962 (N_7962,N_7755,N_7792);
and U7963 (N_7963,N_7619,N_7730);
nand U7964 (N_7964,N_7661,N_7706);
nand U7965 (N_7965,N_7749,N_7604);
nor U7966 (N_7966,N_7612,N_7630);
nand U7967 (N_7967,N_7629,N_7759);
nand U7968 (N_7968,N_7695,N_7740);
or U7969 (N_7969,N_7633,N_7660);
nand U7970 (N_7970,N_7714,N_7694);
and U7971 (N_7971,N_7734,N_7638);
and U7972 (N_7972,N_7682,N_7788);
or U7973 (N_7973,N_7761,N_7729);
and U7974 (N_7974,N_7677,N_7739);
or U7975 (N_7975,N_7785,N_7715);
nand U7976 (N_7976,N_7766,N_7674);
xnor U7977 (N_7977,N_7653,N_7760);
nor U7978 (N_7978,N_7699,N_7641);
nor U7979 (N_7979,N_7759,N_7706);
or U7980 (N_7980,N_7798,N_7796);
nand U7981 (N_7981,N_7729,N_7733);
nor U7982 (N_7982,N_7628,N_7774);
nor U7983 (N_7983,N_7703,N_7675);
nand U7984 (N_7984,N_7622,N_7730);
nand U7985 (N_7985,N_7754,N_7623);
nor U7986 (N_7986,N_7645,N_7610);
xnor U7987 (N_7987,N_7765,N_7677);
nor U7988 (N_7988,N_7679,N_7680);
nand U7989 (N_7989,N_7631,N_7790);
xnor U7990 (N_7990,N_7776,N_7767);
and U7991 (N_7991,N_7617,N_7623);
xor U7992 (N_7992,N_7711,N_7748);
or U7993 (N_7993,N_7771,N_7677);
nand U7994 (N_7994,N_7603,N_7646);
nand U7995 (N_7995,N_7731,N_7631);
nand U7996 (N_7996,N_7779,N_7766);
and U7997 (N_7997,N_7604,N_7630);
and U7998 (N_7998,N_7649,N_7755);
nand U7999 (N_7999,N_7728,N_7600);
or U8000 (N_8000,N_7983,N_7876);
or U8001 (N_8001,N_7841,N_7850);
nor U8002 (N_8002,N_7879,N_7913);
and U8003 (N_8003,N_7940,N_7887);
xnor U8004 (N_8004,N_7809,N_7821);
or U8005 (N_8005,N_7910,N_7816);
or U8006 (N_8006,N_7902,N_7814);
or U8007 (N_8007,N_7939,N_7999);
xor U8008 (N_8008,N_7803,N_7901);
nand U8009 (N_8009,N_7925,N_7843);
xor U8010 (N_8010,N_7893,N_7853);
and U8011 (N_8011,N_7963,N_7981);
nor U8012 (N_8012,N_7811,N_7996);
or U8013 (N_8013,N_7878,N_7896);
nor U8014 (N_8014,N_7865,N_7951);
xnor U8015 (N_8015,N_7802,N_7840);
nand U8016 (N_8016,N_7829,N_7903);
nor U8017 (N_8017,N_7921,N_7942);
nor U8018 (N_8018,N_7884,N_7997);
or U8019 (N_8019,N_7849,N_7958);
nand U8020 (N_8020,N_7881,N_7904);
nor U8021 (N_8021,N_7916,N_7860);
nor U8022 (N_8022,N_7808,N_7810);
or U8023 (N_8023,N_7883,N_7987);
nand U8024 (N_8024,N_7858,N_7974);
or U8025 (N_8025,N_7842,N_7936);
or U8026 (N_8026,N_7817,N_7854);
and U8027 (N_8027,N_7895,N_7872);
nand U8028 (N_8028,N_7859,N_7880);
xnor U8029 (N_8029,N_7863,N_7973);
xor U8030 (N_8030,N_7915,N_7823);
nor U8031 (N_8031,N_7846,N_7833);
nand U8032 (N_8032,N_7815,N_7870);
nor U8033 (N_8033,N_7929,N_7948);
nor U8034 (N_8034,N_7914,N_7969);
nor U8035 (N_8035,N_7978,N_7831);
xnor U8036 (N_8036,N_7839,N_7819);
xnor U8037 (N_8037,N_7947,N_7826);
nor U8038 (N_8038,N_7877,N_7970);
and U8039 (N_8039,N_7824,N_7888);
nor U8040 (N_8040,N_7907,N_7874);
nor U8041 (N_8041,N_7861,N_7834);
nand U8042 (N_8042,N_7968,N_7998);
or U8043 (N_8043,N_7922,N_7830);
and U8044 (N_8044,N_7965,N_7852);
and U8045 (N_8045,N_7889,N_7971);
nand U8046 (N_8046,N_7952,N_7835);
nor U8047 (N_8047,N_7945,N_7825);
or U8048 (N_8048,N_7933,N_7966);
or U8049 (N_8049,N_7924,N_7801);
nand U8050 (N_8050,N_7986,N_7920);
nand U8051 (N_8051,N_7812,N_7931);
or U8052 (N_8052,N_7905,N_7950);
and U8053 (N_8053,N_7908,N_7982);
and U8054 (N_8054,N_7937,N_7934);
nand U8055 (N_8055,N_7857,N_7953);
or U8056 (N_8056,N_7882,N_7837);
or U8057 (N_8057,N_7984,N_7873);
nor U8058 (N_8058,N_7898,N_7805);
and U8059 (N_8059,N_7906,N_7890);
nand U8060 (N_8060,N_7899,N_7979);
nand U8061 (N_8061,N_7868,N_7862);
and U8062 (N_8062,N_7961,N_7990);
nand U8063 (N_8063,N_7957,N_7894);
and U8064 (N_8064,N_7891,N_7962);
or U8065 (N_8065,N_7946,N_7995);
nor U8066 (N_8066,N_7992,N_7960);
nor U8067 (N_8067,N_7855,N_7935);
nand U8068 (N_8068,N_7827,N_7991);
and U8069 (N_8069,N_7836,N_7919);
and U8070 (N_8070,N_7828,N_7926);
or U8071 (N_8071,N_7869,N_7806);
xor U8072 (N_8072,N_7975,N_7800);
and U8073 (N_8073,N_7930,N_7844);
and U8074 (N_8074,N_7911,N_7980);
nor U8075 (N_8075,N_7993,N_7923);
and U8076 (N_8076,N_7832,N_7856);
nor U8077 (N_8077,N_7917,N_7985);
or U8078 (N_8078,N_7964,N_7954);
or U8079 (N_8079,N_7818,N_7956);
or U8080 (N_8080,N_7813,N_7820);
nor U8081 (N_8081,N_7897,N_7967);
and U8082 (N_8082,N_7928,N_7955);
and U8083 (N_8083,N_7909,N_7912);
xor U8084 (N_8084,N_7848,N_7838);
nor U8085 (N_8085,N_7847,N_7900);
or U8086 (N_8086,N_7972,N_7867);
and U8087 (N_8087,N_7851,N_7977);
nor U8088 (N_8088,N_7864,N_7949);
nor U8089 (N_8089,N_7944,N_7871);
or U8090 (N_8090,N_7804,N_7875);
and U8091 (N_8091,N_7932,N_7918);
or U8092 (N_8092,N_7845,N_7866);
nand U8093 (N_8093,N_7927,N_7807);
nand U8094 (N_8094,N_7994,N_7976);
and U8095 (N_8095,N_7988,N_7885);
xnor U8096 (N_8096,N_7989,N_7886);
or U8097 (N_8097,N_7943,N_7938);
and U8098 (N_8098,N_7959,N_7892);
nor U8099 (N_8099,N_7822,N_7941);
xor U8100 (N_8100,N_7808,N_7905);
nor U8101 (N_8101,N_7963,N_7900);
or U8102 (N_8102,N_7976,N_7800);
xor U8103 (N_8103,N_7835,N_7897);
nor U8104 (N_8104,N_7927,N_7931);
nor U8105 (N_8105,N_7832,N_7838);
xnor U8106 (N_8106,N_7893,N_7813);
or U8107 (N_8107,N_7811,N_7889);
or U8108 (N_8108,N_7934,N_7912);
nand U8109 (N_8109,N_7837,N_7832);
and U8110 (N_8110,N_7887,N_7879);
nor U8111 (N_8111,N_7986,N_7971);
nor U8112 (N_8112,N_7861,N_7918);
nand U8113 (N_8113,N_7874,N_7888);
xor U8114 (N_8114,N_7889,N_7836);
and U8115 (N_8115,N_7805,N_7902);
nor U8116 (N_8116,N_7946,N_7844);
xnor U8117 (N_8117,N_7853,N_7972);
nor U8118 (N_8118,N_7977,N_7850);
xor U8119 (N_8119,N_7906,N_7937);
nor U8120 (N_8120,N_7895,N_7855);
and U8121 (N_8121,N_7901,N_7844);
nor U8122 (N_8122,N_7845,N_7973);
nand U8123 (N_8123,N_7872,N_7991);
and U8124 (N_8124,N_7950,N_7819);
or U8125 (N_8125,N_7866,N_7888);
nor U8126 (N_8126,N_7890,N_7807);
or U8127 (N_8127,N_7921,N_7833);
nand U8128 (N_8128,N_7882,N_7998);
and U8129 (N_8129,N_7937,N_7995);
and U8130 (N_8130,N_7975,N_7899);
and U8131 (N_8131,N_7917,N_7949);
and U8132 (N_8132,N_7842,N_7943);
nand U8133 (N_8133,N_7961,N_7831);
and U8134 (N_8134,N_7996,N_7942);
and U8135 (N_8135,N_7903,N_7801);
nand U8136 (N_8136,N_7993,N_7802);
and U8137 (N_8137,N_7817,N_7883);
nor U8138 (N_8138,N_7908,N_7838);
nand U8139 (N_8139,N_7819,N_7876);
or U8140 (N_8140,N_7957,N_7951);
or U8141 (N_8141,N_7886,N_7952);
nand U8142 (N_8142,N_7907,N_7900);
nand U8143 (N_8143,N_7966,N_7960);
nor U8144 (N_8144,N_7841,N_7826);
nor U8145 (N_8145,N_7885,N_7915);
nand U8146 (N_8146,N_7951,N_7805);
and U8147 (N_8147,N_7872,N_7896);
xor U8148 (N_8148,N_7916,N_7948);
nand U8149 (N_8149,N_7901,N_7991);
nor U8150 (N_8150,N_7804,N_7851);
and U8151 (N_8151,N_7984,N_7885);
xnor U8152 (N_8152,N_7805,N_7946);
nor U8153 (N_8153,N_7916,N_7968);
and U8154 (N_8154,N_7850,N_7827);
nor U8155 (N_8155,N_7910,N_7949);
xor U8156 (N_8156,N_7995,N_7919);
nand U8157 (N_8157,N_7998,N_7865);
nand U8158 (N_8158,N_7870,N_7959);
and U8159 (N_8159,N_7976,N_7867);
nand U8160 (N_8160,N_7889,N_7835);
or U8161 (N_8161,N_7849,N_7860);
nand U8162 (N_8162,N_7959,N_7823);
nand U8163 (N_8163,N_7988,N_7890);
nand U8164 (N_8164,N_7875,N_7837);
and U8165 (N_8165,N_7851,N_7865);
and U8166 (N_8166,N_7868,N_7913);
nand U8167 (N_8167,N_7878,N_7845);
nand U8168 (N_8168,N_7918,N_7951);
nor U8169 (N_8169,N_7839,N_7811);
and U8170 (N_8170,N_7856,N_7855);
xor U8171 (N_8171,N_7924,N_7803);
or U8172 (N_8172,N_7880,N_7816);
nor U8173 (N_8173,N_7852,N_7873);
or U8174 (N_8174,N_7844,N_7980);
or U8175 (N_8175,N_7974,N_7959);
or U8176 (N_8176,N_7905,N_7910);
nand U8177 (N_8177,N_7955,N_7896);
xnor U8178 (N_8178,N_7996,N_7974);
nor U8179 (N_8179,N_7802,N_7933);
nand U8180 (N_8180,N_7832,N_7983);
nor U8181 (N_8181,N_7863,N_7889);
xor U8182 (N_8182,N_7953,N_7961);
nor U8183 (N_8183,N_7957,N_7851);
xnor U8184 (N_8184,N_7946,N_7918);
xnor U8185 (N_8185,N_7922,N_7998);
nand U8186 (N_8186,N_7860,N_7957);
or U8187 (N_8187,N_7833,N_7950);
nand U8188 (N_8188,N_7935,N_7857);
nand U8189 (N_8189,N_7974,N_7904);
nor U8190 (N_8190,N_7833,N_7899);
nand U8191 (N_8191,N_7809,N_7882);
nand U8192 (N_8192,N_7868,N_7904);
or U8193 (N_8193,N_7852,N_7835);
or U8194 (N_8194,N_7800,N_7874);
and U8195 (N_8195,N_7921,N_7893);
nor U8196 (N_8196,N_7854,N_7872);
and U8197 (N_8197,N_7959,N_7990);
and U8198 (N_8198,N_7832,N_7829);
and U8199 (N_8199,N_7949,N_7837);
nor U8200 (N_8200,N_8134,N_8010);
and U8201 (N_8201,N_8084,N_8067);
and U8202 (N_8202,N_8099,N_8153);
and U8203 (N_8203,N_8094,N_8112);
or U8204 (N_8204,N_8035,N_8012);
xnor U8205 (N_8205,N_8038,N_8002);
or U8206 (N_8206,N_8106,N_8144);
and U8207 (N_8207,N_8042,N_8048);
nor U8208 (N_8208,N_8162,N_8051);
nor U8209 (N_8209,N_8169,N_8107);
nor U8210 (N_8210,N_8079,N_8114);
nand U8211 (N_8211,N_8104,N_8196);
xor U8212 (N_8212,N_8088,N_8136);
nor U8213 (N_8213,N_8192,N_8052);
nor U8214 (N_8214,N_8062,N_8183);
and U8215 (N_8215,N_8009,N_8050);
or U8216 (N_8216,N_8022,N_8131);
xor U8217 (N_8217,N_8003,N_8014);
nand U8218 (N_8218,N_8057,N_8015);
nor U8219 (N_8219,N_8118,N_8055);
or U8220 (N_8220,N_8066,N_8054);
and U8221 (N_8221,N_8071,N_8121);
and U8222 (N_8222,N_8115,N_8164);
xor U8223 (N_8223,N_8081,N_8069);
nand U8224 (N_8224,N_8182,N_8140);
and U8225 (N_8225,N_8168,N_8004);
or U8226 (N_8226,N_8105,N_8065);
nor U8227 (N_8227,N_8155,N_8158);
nor U8228 (N_8228,N_8124,N_8018);
or U8229 (N_8229,N_8195,N_8150);
nor U8230 (N_8230,N_8117,N_8008);
or U8231 (N_8231,N_8126,N_8111);
nor U8232 (N_8232,N_8093,N_8023);
and U8233 (N_8233,N_8078,N_8113);
or U8234 (N_8234,N_8119,N_8013);
or U8235 (N_8235,N_8040,N_8125);
xnor U8236 (N_8236,N_8146,N_8019);
nand U8237 (N_8237,N_8076,N_8047);
nand U8238 (N_8238,N_8020,N_8075);
nand U8239 (N_8239,N_8089,N_8096);
or U8240 (N_8240,N_8177,N_8072);
nor U8241 (N_8241,N_8049,N_8141);
nor U8242 (N_8242,N_8039,N_8030);
and U8243 (N_8243,N_8036,N_8056);
xnor U8244 (N_8244,N_8142,N_8170);
or U8245 (N_8245,N_8191,N_8083);
and U8246 (N_8246,N_8184,N_8095);
and U8247 (N_8247,N_8100,N_8011);
xnor U8248 (N_8248,N_8154,N_8180);
or U8249 (N_8249,N_8133,N_8090);
nand U8250 (N_8250,N_8034,N_8176);
nor U8251 (N_8251,N_8102,N_8198);
or U8252 (N_8252,N_8122,N_8138);
nand U8253 (N_8253,N_8046,N_8033);
nor U8254 (N_8254,N_8027,N_8001);
nor U8255 (N_8255,N_8109,N_8197);
nor U8256 (N_8256,N_8061,N_8092);
and U8257 (N_8257,N_8173,N_8186);
xnor U8258 (N_8258,N_8108,N_8159);
or U8259 (N_8259,N_8181,N_8139);
or U8260 (N_8260,N_8151,N_8044);
nor U8261 (N_8261,N_8080,N_8145);
nor U8262 (N_8262,N_8127,N_8156);
nor U8263 (N_8263,N_8070,N_8058);
xor U8264 (N_8264,N_8185,N_8161);
nor U8265 (N_8265,N_8123,N_8152);
or U8266 (N_8266,N_8160,N_8025);
nor U8267 (N_8267,N_8194,N_8116);
nand U8268 (N_8268,N_8187,N_8086);
nor U8269 (N_8269,N_8000,N_8016);
or U8270 (N_8270,N_8068,N_8073);
and U8271 (N_8271,N_8179,N_8091);
nand U8272 (N_8272,N_8037,N_8166);
and U8273 (N_8273,N_8026,N_8110);
and U8274 (N_8274,N_8163,N_8147);
nor U8275 (N_8275,N_8053,N_8193);
nand U8276 (N_8276,N_8097,N_8077);
nand U8277 (N_8277,N_8006,N_8157);
and U8278 (N_8278,N_8064,N_8074);
xor U8279 (N_8279,N_8021,N_8043);
or U8280 (N_8280,N_8172,N_8059);
nand U8281 (N_8281,N_8101,N_8199);
xor U8282 (N_8282,N_8024,N_8028);
nand U8283 (N_8283,N_8128,N_8032);
nor U8284 (N_8284,N_8031,N_8130);
or U8285 (N_8285,N_8045,N_8135);
nor U8286 (N_8286,N_8174,N_8017);
and U8287 (N_8287,N_8132,N_8063);
or U8288 (N_8288,N_8149,N_8120);
and U8289 (N_8289,N_8143,N_8129);
nor U8290 (N_8290,N_8029,N_8007);
nand U8291 (N_8291,N_8060,N_8148);
nor U8292 (N_8292,N_8085,N_8082);
xnor U8293 (N_8293,N_8189,N_8098);
nor U8294 (N_8294,N_8188,N_8041);
and U8295 (N_8295,N_8087,N_8103);
xnor U8296 (N_8296,N_8178,N_8165);
or U8297 (N_8297,N_8175,N_8167);
or U8298 (N_8298,N_8137,N_8190);
nand U8299 (N_8299,N_8005,N_8171);
nand U8300 (N_8300,N_8127,N_8148);
and U8301 (N_8301,N_8070,N_8146);
and U8302 (N_8302,N_8117,N_8192);
nand U8303 (N_8303,N_8028,N_8161);
or U8304 (N_8304,N_8037,N_8112);
or U8305 (N_8305,N_8133,N_8189);
or U8306 (N_8306,N_8149,N_8003);
or U8307 (N_8307,N_8171,N_8123);
and U8308 (N_8308,N_8141,N_8104);
nand U8309 (N_8309,N_8029,N_8183);
nor U8310 (N_8310,N_8037,N_8120);
and U8311 (N_8311,N_8012,N_8100);
nor U8312 (N_8312,N_8036,N_8160);
and U8313 (N_8313,N_8081,N_8115);
and U8314 (N_8314,N_8001,N_8008);
nor U8315 (N_8315,N_8143,N_8034);
nor U8316 (N_8316,N_8050,N_8078);
and U8317 (N_8317,N_8000,N_8187);
xor U8318 (N_8318,N_8077,N_8062);
and U8319 (N_8319,N_8193,N_8130);
xor U8320 (N_8320,N_8055,N_8112);
nand U8321 (N_8321,N_8077,N_8195);
nand U8322 (N_8322,N_8146,N_8121);
and U8323 (N_8323,N_8167,N_8080);
nor U8324 (N_8324,N_8101,N_8111);
or U8325 (N_8325,N_8056,N_8032);
or U8326 (N_8326,N_8064,N_8117);
nand U8327 (N_8327,N_8079,N_8130);
nor U8328 (N_8328,N_8000,N_8161);
nor U8329 (N_8329,N_8166,N_8143);
nand U8330 (N_8330,N_8191,N_8117);
nand U8331 (N_8331,N_8105,N_8097);
xnor U8332 (N_8332,N_8016,N_8109);
nor U8333 (N_8333,N_8084,N_8013);
or U8334 (N_8334,N_8161,N_8119);
and U8335 (N_8335,N_8093,N_8092);
or U8336 (N_8336,N_8177,N_8174);
nor U8337 (N_8337,N_8157,N_8175);
nor U8338 (N_8338,N_8082,N_8197);
nor U8339 (N_8339,N_8095,N_8134);
or U8340 (N_8340,N_8115,N_8021);
nand U8341 (N_8341,N_8021,N_8000);
or U8342 (N_8342,N_8025,N_8034);
nand U8343 (N_8343,N_8077,N_8032);
nand U8344 (N_8344,N_8164,N_8002);
and U8345 (N_8345,N_8036,N_8167);
xnor U8346 (N_8346,N_8192,N_8118);
nor U8347 (N_8347,N_8068,N_8176);
nor U8348 (N_8348,N_8030,N_8071);
nor U8349 (N_8349,N_8111,N_8038);
and U8350 (N_8350,N_8147,N_8096);
nand U8351 (N_8351,N_8087,N_8164);
nor U8352 (N_8352,N_8183,N_8054);
nor U8353 (N_8353,N_8090,N_8196);
and U8354 (N_8354,N_8081,N_8097);
and U8355 (N_8355,N_8144,N_8184);
or U8356 (N_8356,N_8075,N_8132);
xor U8357 (N_8357,N_8162,N_8145);
and U8358 (N_8358,N_8114,N_8166);
nand U8359 (N_8359,N_8043,N_8038);
nor U8360 (N_8360,N_8069,N_8140);
nand U8361 (N_8361,N_8178,N_8041);
or U8362 (N_8362,N_8051,N_8068);
nor U8363 (N_8363,N_8031,N_8170);
nand U8364 (N_8364,N_8007,N_8024);
or U8365 (N_8365,N_8024,N_8053);
or U8366 (N_8366,N_8162,N_8104);
or U8367 (N_8367,N_8173,N_8028);
nand U8368 (N_8368,N_8006,N_8038);
nand U8369 (N_8369,N_8142,N_8055);
and U8370 (N_8370,N_8193,N_8017);
or U8371 (N_8371,N_8073,N_8064);
nor U8372 (N_8372,N_8091,N_8182);
xor U8373 (N_8373,N_8190,N_8058);
or U8374 (N_8374,N_8089,N_8041);
nor U8375 (N_8375,N_8047,N_8193);
or U8376 (N_8376,N_8013,N_8191);
nand U8377 (N_8377,N_8034,N_8192);
nor U8378 (N_8378,N_8022,N_8093);
nand U8379 (N_8379,N_8077,N_8173);
xnor U8380 (N_8380,N_8142,N_8085);
nand U8381 (N_8381,N_8059,N_8043);
nand U8382 (N_8382,N_8157,N_8058);
nor U8383 (N_8383,N_8182,N_8108);
or U8384 (N_8384,N_8161,N_8089);
and U8385 (N_8385,N_8188,N_8015);
and U8386 (N_8386,N_8140,N_8051);
or U8387 (N_8387,N_8072,N_8153);
nand U8388 (N_8388,N_8065,N_8066);
nor U8389 (N_8389,N_8070,N_8015);
nor U8390 (N_8390,N_8007,N_8068);
nand U8391 (N_8391,N_8021,N_8096);
and U8392 (N_8392,N_8138,N_8127);
or U8393 (N_8393,N_8094,N_8190);
and U8394 (N_8394,N_8124,N_8148);
nand U8395 (N_8395,N_8143,N_8139);
or U8396 (N_8396,N_8178,N_8059);
and U8397 (N_8397,N_8174,N_8193);
nand U8398 (N_8398,N_8164,N_8066);
or U8399 (N_8399,N_8102,N_8040);
nand U8400 (N_8400,N_8316,N_8380);
nand U8401 (N_8401,N_8272,N_8233);
and U8402 (N_8402,N_8269,N_8254);
xor U8403 (N_8403,N_8318,N_8291);
nor U8404 (N_8404,N_8245,N_8236);
nor U8405 (N_8405,N_8350,N_8284);
nor U8406 (N_8406,N_8265,N_8220);
or U8407 (N_8407,N_8268,N_8280);
nand U8408 (N_8408,N_8369,N_8386);
and U8409 (N_8409,N_8256,N_8359);
nand U8410 (N_8410,N_8261,N_8240);
and U8411 (N_8411,N_8375,N_8344);
and U8412 (N_8412,N_8297,N_8204);
nand U8413 (N_8413,N_8320,N_8317);
and U8414 (N_8414,N_8276,N_8208);
nor U8415 (N_8415,N_8215,N_8299);
xnor U8416 (N_8416,N_8331,N_8293);
or U8417 (N_8417,N_8311,N_8294);
nor U8418 (N_8418,N_8388,N_8252);
or U8419 (N_8419,N_8363,N_8378);
or U8420 (N_8420,N_8301,N_8259);
or U8421 (N_8421,N_8289,N_8360);
and U8422 (N_8422,N_8211,N_8243);
or U8423 (N_8423,N_8342,N_8367);
and U8424 (N_8424,N_8321,N_8308);
nor U8425 (N_8425,N_8307,N_8341);
nand U8426 (N_8426,N_8336,N_8214);
or U8427 (N_8427,N_8387,N_8389);
xor U8428 (N_8428,N_8257,N_8205);
or U8429 (N_8429,N_8264,N_8353);
nand U8430 (N_8430,N_8234,N_8343);
or U8431 (N_8431,N_8248,N_8267);
and U8432 (N_8432,N_8271,N_8393);
nand U8433 (N_8433,N_8273,N_8290);
or U8434 (N_8434,N_8221,N_8326);
or U8435 (N_8435,N_8298,N_8282);
nand U8436 (N_8436,N_8228,N_8315);
nand U8437 (N_8437,N_8223,N_8305);
and U8438 (N_8438,N_8266,N_8366);
or U8439 (N_8439,N_8255,N_8399);
nand U8440 (N_8440,N_8382,N_8246);
nor U8441 (N_8441,N_8242,N_8296);
xor U8442 (N_8442,N_8351,N_8355);
nand U8443 (N_8443,N_8306,N_8209);
and U8444 (N_8444,N_8300,N_8322);
xnor U8445 (N_8445,N_8227,N_8262);
or U8446 (N_8446,N_8295,N_8314);
nand U8447 (N_8447,N_8260,N_8338);
nor U8448 (N_8448,N_8225,N_8325);
and U8449 (N_8449,N_8332,N_8330);
xnor U8450 (N_8450,N_8258,N_8231);
or U8451 (N_8451,N_8218,N_8312);
nor U8452 (N_8452,N_8287,N_8337);
nor U8453 (N_8453,N_8224,N_8244);
and U8454 (N_8454,N_8206,N_8212);
nor U8455 (N_8455,N_8201,N_8286);
nand U8456 (N_8456,N_8381,N_8313);
or U8457 (N_8457,N_8251,N_8373);
xor U8458 (N_8458,N_8370,N_8334);
and U8459 (N_8459,N_8395,N_8340);
and U8460 (N_8460,N_8232,N_8222);
and U8461 (N_8461,N_8207,N_8278);
nand U8462 (N_8462,N_8239,N_8213);
or U8463 (N_8463,N_8217,N_8292);
and U8464 (N_8464,N_8249,N_8302);
and U8465 (N_8465,N_8376,N_8358);
xnor U8466 (N_8466,N_8391,N_8202);
nor U8467 (N_8467,N_8394,N_8200);
xor U8468 (N_8468,N_8319,N_8390);
nand U8469 (N_8469,N_8235,N_8247);
nand U8470 (N_8470,N_8281,N_8396);
nor U8471 (N_8471,N_8323,N_8229);
and U8472 (N_8472,N_8203,N_8329);
nand U8473 (N_8473,N_8398,N_8333);
or U8474 (N_8474,N_8230,N_8374);
nor U8475 (N_8475,N_8279,N_8377);
and U8476 (N_8476,N_8339,N_8361);
nand U8477 (N_8477,N_8241,N_8238);
nor U8478 (N_8478,N_8304,N_8237);
and U8479 (N_8479,N_8349,N_8285);
nor U8480 (N_8480,N_8270,N_8365);
and U8481 (N_8481,N_8354,N_8356);
nand U8482 (N_8482,N_8385,N_8364);
nor U8483 (N_8483,N_8216,N_8328);
or U8484 (N_8484,N_8277,N_8379);
and U8485 (N_8485,N_8324,N_8253);
nor U8486 (N_8486,N_8309,N_8383);
or U8487 (N_8487,N_8303,N_8275);
or U8488 (N_8488,N_8346,N_8348);
nand U8489 (N_8489,N_8327,N_8352);
nor U8490 (N_8490,N_8335,N_8357);
or U8491 (N_8491,N_8397,N_8310);
nor U8492 (N_8492,N_8372,N_8283);
nand U8493 (N_8493,N_8226,N_8219);
nor U8494 (N_8494,N_8263,N_8368);
and U8495 (N_8495,N_8347,N_8392);
xnor U8496 (N_8496,N_8371,N_8362);
nor U8497 (N_8497,N_8210,N_8288);
or U8498 (N_8498,N_8250,N_8274);
and U8499 (N_8499,N_8345,N_8384);
nand U8500 (N_8500,N_8329,N_8395);
and U8501 (N_8501,N_8383,N_8289);
nor U8502 (N_8502,N_8285,N_8301);
nand U8503 (N_8503,N_8312,N_8389);
and U8504 (N_8504,N_8370,N_8355);
and U8505 (N_8505,N_8294,N_8223);
and U8506 (N_8506,N_8282,N_8311);
nand U8507 (N_8507,N_8377,N_8393);
nand U8508 (N_8508,N_8330,N_8274);
nand U8509 (N_8509,N_8289,N_8359);
or U8510 (N_8510,N_8264,N_8363);
or U8511 (N_8511,N_8385,N_8387);
xor U8512 (N_8512,N_8295,N_8241);
xnor U8513 (N_8513,N_8283,N_8276);
nand U8514 (N_8514,N_8279,N_8222);
or U8515 (N_8515,N_8242,N_8342);
or U8516 (N_8516,N_8253,N_8354);
and U8517 (N_8517,N_8224,N_8260);
nor U8518 (N_8518,N_8212,N_8308);
nor U8519 (N_8519,N_8301,N_8204);
and U8520 (N_8520,N_8353,N_8274);
or U8521 (N_8521,N_8239,N_8303);
nand U8522 (N_8522,N_8310,N_8314);
nand U8523 (N_8523,N_8260,N_8340);
nand U8524 (N_8524,N_8249,N_8355);
nor U8525 (N_8525,N_8316,N_8253);
nand U8526 (N_8526,N_8330,N_8381);
nand U8527 (N_8527,N_8274,N_8203);
or U8528 (N_8528,N_8338,N_8268);
xnor U8529 (N_8529,N_8334,N_8342);
xor U8530 (N_8530,N_8392,N_8363);
nand U8531 (N_8531,N_8260,N_8308);
and U8532 (N_8532,N_8354,N_8210);
and U8533 (N_8533,N_8202,N_8246);
nor U8534 (N_8534,N_8377,N_8240);
nand U8535 (N_8535,N_8276,N_8328);
xor U8536 (N_8536,N_8356,N_8243);
and U8537 (N_8537,N_8369,N_8252);
nor U8538 (N_8538,N_8319,N_8374);
nand U8539 (N_8539,N_8242,N_8306);
nor U8540 (N_8540,N_8223,N_8302);
or U8541 (N_8541,N_8320,N_8362);
xnor U8542 (N_8542,N_8397,N_8268);
nor U8543 (N_8543,N_8321,N_8326);
nor U8544 (N_8544,N_8347,N_8272);
nand U8545 (N_8545,N_8329,N_8398);
xnor U8546 (N_8546,N_8291,N_8310);
or U8547 (N_8547,N_8250,N_8261);
xnor U8548 (N_8548,N_8210,N_8314);
or U8549 (N_8549,N_8218,N_8341);
xnor U8550 (N_8550,N_8386,N_8238);
nand U8551 (N_8551,N_8362,N_8395);
nand U8552 (N_8552,N_8396,N_8383);
and U8553 (N_8553,N_8341,N_8258);
xor U8554 (N_8554,N_8237,N_8396);
and U8555 (N_8555,N_8297,N_8306);
or U8556 (N_8556,N_8208,N_8299);
or U8557 (N_8557,N_8367,N_8338);
nor U8558 (N_8558,N_8271,N_8295);
nand U8559 (N_8559,N_8283,N_8330);
or U8560 (N_8560,N_8289,N_8313);
xor U8561 (N_8561,N_8217,N_8307);
xor U8562 (N_8562,N_8333,N_8223);
nor U8563 (N_8563,N_8360,N_8231);
and U8564 (N_8564,N_8377,N_8392);
nand U8565 (N_8565,N_8280,N_8250);
or U8566 (N_8566,N_8299,N_8283);
xnor U8567 (N_8567,N_8224,N_8319);
nand U8568 (N_8568,N_8358,N_8216);
nor U8569 (N_8569,N_8357,N_8328);
nand U8570 (N_8570,N_8275,N_8299);
nor U8571 (N_8571,N_8219,N_8327);
and U8572 (N_8572,N_8385,N_8321);
and U8573 (N_8573,N_8241,N_8232);
nor U8574 (N_8574,N_8286,N_8344);
nor U8575 (N_8575,N_8206,N_8307);
xnor U8576 (N_8576,N_8321,N_8271);
and U8577 (N_8577,N_8320,N_8215);
nand U8578 (N_8578,N_8243,N_8234);
nand U8579 (N_8579,N_8245,N_8201);
nor U8580 (N_8580,N_8208,N_8355);
or U8581 (N_8581,N_8323,N_8258);
xnor U8582 (N_8582,N_8380,N_8322);
nand U8583 (N_8583,N_8269,N_8362);
xor U8584 (N_8584,N_8334,N_8329);
nor U8585 (N_8585,N_8312,N_8383);
or U8586 (N_8586,N_8234,N_8276);
nand U8587 (N_8587,N_8267,N_8258);
and U8588 (N_8588,N_8344,N_8296);
xor U8589 (N_8589,N_8205,N_8396);
or U8590 (N_8590,N_8238,N_8399);
and U8591 (N_8591,N_8234,N_8372);
nand U8592 (N_8592,N_8297,N_8354);
xnor U8593 (N_8593,N_8226,N_8279);
or U8594 (N_8594,N_8224,N_8262);
and U8595 (N_8595,N_8302,N_8352);
and U8596 (N_8596,N_8258,N_8342);
and U8597 (N_8597,N_8369,N_8316);
or U8598 (N_8598,N_8333,N_8208);
xor U8599 (N_8599,N_8224,N_8277);
nand U8600 (N_8600,N_8568,N_8567);
nor U8601 (N_8601,N_8493,N_8468);
and U8602 (N_8602,N_8471,N_8502);
or U8603 (N_8603,N_8559,N_8403);
nor U8604 (N_8604,N_8505,N_8456);
and U8605 (N_8605,N_8474,N_8506);
xor U8606 (N_8606,N_8418,N_8545);
nor U8607 (N_8607,N_8484,N_8566);
and U8608 (N_8608,N_8569,N_8525);
nor U8609 (N_8609,N_8512,N_8571);
or U8610 (N_8610,N_8446,N_8428);
and U8611 (N_8611,N_8576,N_8497);
nand U8612 (N_8612,N_8508,N_8549);
nor U8613 (N_8613,N_8521,N_8432);
and U8614 (N_8614,N_8444,N_8530);
and U8615 (N_8615,N_8542,N_8458);
nand U8616 (N_8616,N_8533,N_8591);
nor U8617 (N_8617,N_8452,N_8597);
nand U8618 (N_8618,N_8478,N_8408);
or U8619 (N_8619,N_8539,N_8570);
nand U8620 (N_8620,N_8555,N_8472);
and U8621 (N_8621,N_8504,N_8548);
nand U8622 (N_8622,N_8494,N_8435);
or U8623 (N_8623,N_8424,N_8422);
or U8624 (N_8624,N_8550,N_8466);
or U8625 (N_8625,N_8415,N_8528);
nand U8626 (N_8626,N_8414,N_8420);
nor U8627 (N_8627,N_8487,N_8522);
xor U8628 (N_8628,N_8437,N_8585);
nor U8629 (N_8629,N_8595,N_8433);
and U8630 (N_8630,N_8573,N_8515);
nand U8631 (N_8631,N_8543,N_8479);
nor U8632 (N_8632,N_8495,N_8455);
xnor U8633 (N_8633,N_8412,N_8473);
and U8634 (N_8634,N_8519,N_8580);
nor U8635 (N_8635,N_8590,N_8514);
nor U8636 (N_8636,N_8501,N_8589);
nor U8637 (N_8637,N_8407,N_8593);
xnor U8638 (N_8638,N_8463,N_8450);
and U8639 (N_8639,N_8477,N_8532);
or U8640 (N_8640,N_8465,N_8535);
or U8641 (N_8641,N_8454,N_8413);
and U8642 (N_8642,N_8560,N_8448);
and U8643 (N_8643,N_8547,N_8459);
nor U8644 (N_8644,N_8475,N_8400);
nand U8645 (N_8645,N_8574,N_8561);
nand U8646 (N_8646,N_8578,N_8598);
or U8647 (N_8647,N_8486,N_8411);
or U8648 (N_8648,N_8469,N_8482);
or U8649 (N_8649,N_8503,N_8592);
or U8650 (N_8650,N_8402,N_8527);
or U8651 (N_8651,N_8404,N_8488);
or U8652 (N_8652,N_8431,N_8565);
nand U8653 (N_8653,N_8575,N_8430);
and U8654 (N_8654,N_8409,N_8577);
nand U8655 (N_8655,N_8546,N_8480);
nor U8656 (N_8656,N_8507,N_8537);
and U8657 (N_8657,N_8558,N_8596);
nand U8658 (N_8658,N_8481,N_8554);
nand U8659 (N_8659,N_8594,N_8538);
or U8660 (N_8660,N_8429,N_8496);
or U8661 (N_8661,N_8540,N_8416);
or U8662 (N_8662,N_8586,N_8564);
xor U8663 (N_8663,N_8457,N_8464);
or U8664 (N_8664,N_8417,N_8572);
and U8665 (N_8665,N_8441,N_8584);
or U8666 (N_8666,N_8524,N_8534);
nand U8667 (N_8667,N_8490,N_8520);
nor U8668 (N_8668,N_8401,N_8438);
and U8669 (N_8669,N_8439,N_8557);
nor U8670 (N_8670,N_8579,N_8553);
xor U8671 (N_8671,N_8491,N_8447);
or U8672 (N_8672,N_8442,N_8536);
nor U8673 (N_8673,N_8423,N_8552);
and U8674 (N_8674,N_8498,N_8562);
or U8675 (N_8675,N_8517,N_8510);
or U8676 (N_8676,N_8513,N_8460);
or U8677 (N_8677,N_8563,N_8531);
nor U8678 (N_8678,N_8489,N_8467);
and U8679 (N_8679,N_8427,N_8421);
nor U8680 (N_8680,N_8445,N_8581);
nand U8681 (N_8681,N_8518,N_8476);
and U8682 (N_8682,N_8434,N_8509);
and U8683 (N_8683,N_8544,N_8406);
nor U8684 (N_8684,N_8523,N_8588);
nor U8685 (N_8685,N_8440,N_8419);
or U8686 (N_8686,N_8583,N_8499);
or U8687 (N_8687,N_8426,N_8410);
nor U8688 (N_8688,N_8470,N_8551);
or U8689 (N_8689,N_8462,N_8587);
nand U8690 (N_8690,N_8599,N_8526);
and U8691 (N_8691,N_8541,N_8516);
nor U8692 (N_8692,N_8461,N_8483);
and U8693 (N_8693,N_8443,N_8449);
nand U8694 (N_8694,N_8436,N_8492);
or U8695 (N_8695,N_8485,N_8405);
nor U8696 (N_8696,N_8451,N_8529);
and U8697 (N_8697,N_8425,N_8453);
nor U8698 (N_8698,N_8582,N_8500);
nor U8699 (N_8699,N_8556,N_8511);
and U8700 (N_8700,N_8431,N_8409);
nor U8701 (N_8701,N_8592,N_8406);
nor U8702 (N_8702,N_8499,N_8541);
nor U8703 (N_8703,N_8411,N_8432);
nand U8704 (N_8704,N_8553,N_8436);
nor U8705 (N_8705,N_8499,N_8497);
and U8706 (N_8706,N_8411,N_8531);
xor U8707 (N_8707,N_8592,N_8467);
xor U8708 (N_8708,N_8498,N_8526);
nor U8709 (N_8709,N_8483,N_8403);
xnor U8710 (N_8710,N_8465,N_8585);
and U8711 (N_8711,N_8475,N_8562);
nand U8712 (N_8712,N_8405,N_8473);
or U8713 (N_8713,N_8598,N_8478);
and U8714 (N_8714,N_8523,N_8562);
nor U8715 (N_8715,N_8560,N_8401);
nand U8716 (N_8716,N_8450,N_8542);
or U8717 (N_8717,N_8584,N_8461);
and U8718 (N_8718,N_8434,N_8482);
nand U8719 (N_8719,N_8525,N_8556);
and U8720 (N_8720,N_8411,N_8584);
and U8721 (N_8721,N_8550,N_8558);
nor U8722 (N_8722,N_8460,N_8436);
and U8723 (N_8723,N_8567,N_8581);
and U8724 (N_8724,N_8458,N_8510);
and U8725 (N_8725,N_8465,N_8592);
and U8726 (N_8726,N_8450,N_8408);
xor U8727 (N_8727,N_8594,N_8506);
nand U8728 (N_8728,N_8420,N_8405);
nor U8729 (N_8729,N_8438,N_8489);
and U8730 (N_8730,N_8487,N_8536);
nor U8731 (N_8731,N_8513,N_8465);
nand U8732 (N_8732,N_8585,N_8466);
or U8733 (N_8733,N_8409,N_8422);
nand U8734 (N_8734,N_8412,N_8560);
or U8735 (N_8735,N_8427,N_8414);
or U8736 (N_8736,N_8533,N_8596);
or U8737 (N_8737,N_8567,N_8542);
nand U8738 (N_8738,N_8494,N_8404);
nor U8739 (N_8739,N_8403,N_8455);
and U8740 (N_8740,N_8550,N_8421);
xnor U8741 (N_8741,N_8559,N_8469);
or U8742 (N_8742,N_8496,N_8493);
xnor U8743 (N_8743,N_8410,N_8580);
nand U8744 (N_8744,N_8477,N_8571);
and U8745 (N_8745,N_8429,N_8570);
xnor U8746 (N_8746,N_8539,N_8555);
and U8747 (N_8747,N_8422,N_8505);
nand U8748 (N_8748,N_8562,N_8567);
or U8749 (N_8749,N_8578,N_8420);
nand U8750 (N_8750,N_8516,N_8487);
and U8751 (N_8751,N_8584,N_8529);
nor U8752 (N_8752,N_8408,N_8466);
nand U8753 (N_8753,N_8415,N_8428);
xor U8754 (N_8754,N_8504,N_8552);
nor U8755 (N_8755,N_8574,N_8497);
or U8756 (N_8756,N_8537,N_8588);
and U8757 (N_8757,N_8520,N_8555);
nor U8758 (N_8758,N_8486,N_8503);
or U8759 (N_8759,N_8446,N_8534);
nor U8760 (N_8760,N_8472,N_8501);
nor U8761 (N_8761,N_8402,N_8488);
nand U8762 (N_8762,N_8443,N_8482);
nor U8763 (N_8763,N_8495,N_8570);
nand U8764 (N_8764,N_8450,N_8582);
and U8765 (N_8765,N_8442,N_8481);
and U8766 (N_8766,N_8469,N_8455);
nand U8767 (N_8767,N_8414,N_8446);
nand U8768 (N_8768,N_8536,N_8521);
or U8769 (N_8769,N_8427,N_8534);
nor U8770 (N_8770,N_8419,N_8541);
nor U8771 (N_8771,N_8438,N_8575);
or U8772 (N_8772,N_8497,N_8598);
or U8773 (N_8773,N_8428,N_8548);
xnor U8774 (N_8774,N_8514,N_8555);
nand U8775 (N_8775,N_8454,N_8405);
nand U8776 (N_8776,N_8566,N_8509);
or U8777 (N_8777,N_8566,N_8545);
xor U8778 (N_8778,N_8574,N_8449);
or U8779 (N_8779,N_8523,N_8547);
xor U8780 (N_8780,N_8467,N_8431);
or U8781 (N_8781,N_8540,N_8489);
nor U8782 (N_8782,N_8448,N_8535);
and U8783 (N_8783,N_8442,N_8448);
or U8784 (N_8784,N_8509,N_8569);
and U8785 (N_8785,N_8546,N_8505);
or U8786 (N_8786,N_8589,N_8557);
and U8787 (N_8787,N_8458,N_8561);
or U8788 (N_8788,N_8506,N_8409);
nand U8789 (N_8789,N_8401,N_8520);
and U8790 (N_8790,N_8577,N_8460);
nand U8791 (N_8791,N_8474,N_8593);
or U8792 (N_8792,N_8416,N_8402);
or U8793 (N_8793,N_8432,N_8523);
xor U8794 (N_8794,N_8464,N_8564);
nor U8795 (N_8795,N_8512,N_8515);
nor U8796 (N_8796,N_8411,N_8419);
nand U8797 (N_8797,N_8457,N_8505);
and U8798 (N_8798,N_8587,N_8576);
and U8799 (N_8799,N_8441,N_8496);
nand U8800 (N_8800,N_8709,N_8666);
nand U8801 (N_8801,N_8639,N_8627);
nor U8802 (N_8802,N_8608,N_8729);
nor U8803 (N_8803,N_8669,N_8740);
or U8804 (N_8804,N_8797,N_8605);
or U8805 (N_8805,N_8705,N_8690);
nor U8806 (N_8806,N_8628,N_8730);
nand U8807 (N_8807,N_8675,N_8771);
nor U8808 (N_8808,N_8699,N_8642);
nor U8809 (N_8809,N_8693,N_8781);
nor U8810 (N_8810,N_8659,N_8621);
xnor U8811 (N_8811,N_8710,N_8791);
or U8812 (N_8812,N_8794,N_8623);
xnor U8813 (N_8813,N_8603,N_8650);
and U8814 (N_8814,N_8719,N_8789);
nand U8815 (N_8815,N_8757,N_8681);
nand U8816 (N_8816,N_8640,N_8651);
nor U8817 (N_8817,N_8672,N_8793);
nor U8818 (N_8818,N_8697,N_8796);
and U8819 (N_8819,N_8717,N_8629);
nor U8820 (N_8820,N_8636,N_8773);
or U8821 (N_8821,N_8616,N_8617);
nand U8822 (N_8822,N_8638,N_8695);
or U8823 (N_8823,N_8725,N_8723);
nor U8824 (N_8824,N_8658,N_8714);
or U8825 (N_8825,N_8698,N_8702);
nand U8826 (N_8826,N_8708,N_8611);
nand U8827 (N_8827,N_8600,N_8780);
xnor U8828 (N_8828,N_8786,N_8612);
nand U8829 (N_8829,N_8674,N_8645);
or U8830 (N_8830,N_8715,N_8700);
and U8831 (N_8831,N_8704,N_8798);
or U8832 (N_8832,N_8678,N_8742);
or U8833 (N_8833,N_8722,N_8785);
and U8834 (N_8834,N_8767,N_8686);
nand U8835 (N_8835,N_8754,N_8706);
xnor U8836 (N_8836,N_8653,N_8787);
xnor U8837 (N_8837,N_8790,N_8676);
or U8838 (N_8838,N_8620,N_8689);
xor U8839 (N_8839,N_8683,N_8788);
or U8840 (N_8840,N_8724,N_8738);
nand U8841 (N_8841,N_8602,N_8718);
xnor U8842 (N_8842,N_8663,N_8726);
and U8843 (N_8843,N_8743,N_8774);
xor U8844 (N_8844,N_8641,N_8684);
or U8845 (N_8845,N_8769,N_8735);
or U8846 (N_8846,N_8631,N_8778);
nor U8847 (N_8847,N_8667,N_8759);
nand U8848 (N_8848,N_8652,N_8604);
nor U8849 (N_8849,N_8707,N_8626);
nor U8850 (N_8850,N_8606,N_8739);
nand U8851 (N_8851,N_8758,N_8688);
or U8852 (N_8852,N_8670,N_8745);
nor U8853 (N_8853,N_8712,N_8637);
nor U8854 (N_8854,N_8749,N_8762);
nor U8855 (N_8855,N_8687,N_8727);
or U8856 (N_8856,N_8614,N_8654);
and U8857 (N_8857,N_8664,N_8682);
nor U8858 (N_8858,N_8673,N_8782);
nand U8859 (N_8859,N_8633,N_8662);
and U8860 (N_8860,N_8752,N_8732);
or U8861 (N_8861,N_8711,N_8635);
xnor U8862 (N_8862,N_8799,N_8747);
or U8863 (N_8863,N_8647,N_8756);
nor U8864 (N_8864,N_8755,N_8613);
xor U8865 (N_8865,N_8618,N_8748);
and U8866 (N_8866,N_8792,N_8691);
nor U8867 (N_8867,N_8660,N_8713);
nand U8868 (N_8868,N_8696,N_8655);
and U8869 (N_8869,N_8685,N_8741);
nor U8870 (N_8870,N_8644,N_8734);
or U8871 (N_8871,N_8753,N_8619);
and U8872 (N_8872,N_8783,N_8760);
nand U8873 (N_8873,N_8779,N_8736);
or U8874 (N_8874,N_8648,N_8607);
and U8875 (N_8875,N_8677,N_8643);
or U8876 (N_8876,N_8737,N_8656);
or U8877 (N_8877,N_8601,N_8770);
or U8878 (N_8878,N_8775,N_8622);
nor U8879 (N_8879,N_8610,N_8646);
or U8880 (N_8880,N_8657,N_8777);
nand U8881 (N_8881,N_8615,N_8632);
nor U8882 (N_8882,N_8721,N_8703);
nand U8883 (N_8883,N_8744,N_8761);
or U8884 (N_8884,N_8763,N_8720);
nor U8885 (N_8885,N_8728,N_8750);
or U8886 (N_8886,N_8766,N_8679);
nand U8887 (N_8887,N_8694,N_8701);
and U8888 (N_8888,N_8764,N_8716);
nor U8889 (N_8889,N_8733,N_8692);
or U8890 (N_8890,N_8772,N_8731);
xnor U8891 (N_8891,N_8671,N_8668);
nor U8892 (N_8892,N_8765,N_8624);
xnor U8893 (N_8893,N_8630,N_8625);
nand U8894 (N_8894,N_8609,N_8751);
nand U8895 (N_8895,N_8649,N_8776);
xnor U8896 (N_8896,N_8795,N_8768);
nand U8897 (N_8897,N_8746,N_8784);
nor U8898 (N_8898,N_8665,N_8634);
and U8899 (N_8899,N_8661,N_8680);
nor U8900 (N_8900,N_8627,N_8778);
nand U8901 (N_8901,N_8783,N_8614);
or U8902 (N_8902,N_8607,N_8650);
or U8903 (N_8903,N_8611,N_8771);
xor U8904 (N_8904,N_8648,N_8610);
nand U8905 (N_8905,N_8677,N_8710);
and U8906 (N_8906,N_8757,N_8748);
xnor U8907 (N_8907,N_8787,N_8699);
nor U8908 (N_8908,N_8659,N_8745);
or U8909 (N_8909,N_8782,N_8703);
or U8910 (N_8910,N_8739,N_8720);
or U8911 (N_8911,N_8710,N_8753);
nor U8912 (N_8912,N_8798,N_8635);
nand U8913 (N_8913,N_8656,N_8775);
or U8914 (N_8914,N_8660,N_8618);
nand U8915 (N_8915,N_8791,N_8718);
xnor U8916 (N_8916,N_8673,N_8718);
and U8917 (N_8917,N_8722,N_8721);
and U8918 (N_8918,N_8718,N_8720);
nor U8919 (N_8919,N_8788,N_8695);
nand U8920 (N_8920,N_8632,N_8751);
nor U8921 (N_8921,N_8672,N_8710);
or U8922 (N_8922,N_8682,N_8755);
nand U8923 (N_8923,N_8737,N_8776);
or U8924 (N_8924,N_8775,N_8619);
and U8925 (N_8925,N_8772,N_8666);
and U8926 (N_8926,N_8661,N_8605);
nor U8927 (N_8927,N_8676,N_8660);
nand U8928 (N_8928,N_8781,N_8677);
xnor U8929 (N_8929,N_8752,N_8727);
nand U8930 (N_8930,N_8623,N_8744);
or U8931 (N_8931,N_8716,N_8622);
and U8932 (N_8932,N_8798,N_8685);
nor U8933 (N_8933,N_8622,N_8670);
nor U8934 (N_8934,N_8798,N_8698);
and U8935 (N_8935,N_8791,N_8782);
and U8936 (N_8936,N_8771,N_8739);
nand U8937 (N_8937,N_8724,N_8731);
nor U8938 (N_8938,N_8608,N_8738);
and U8939 (N_8939,N_8612,N_8721);
or U8940 (N_8940,N_8751,N_8752);
and U8941 (N_8941,N_8772,N_8685);
or U8942 (N_8942,N_8709,N_8731);
nor U8943 (N_8943,N_8684,N_8662);
nand U8944 (N_8944,N_8631,N_8747);
nor U8945 (N_8945,N_8670,N_8709);
nand U8946 (N_8946,N_8619,N_8693);
and U8947 (N_8947,N_8731,N_8780);
or U8948 (N_8948,N_8623,N_8650);
nand U8949 (N_8949,N_8742,N_8664);
nor U8950 (N_8950,N_8774,N_8736);
and U8951 (N_8951,N_8622,N_8665);
xor U8952 (N_8952,N_8625,N_8725);
and U8953 (N_8953,N_8716,N_8674);
and U8954 (N_8954,N_8653,N_8625);
nor U8955 (N_8955,N_8655,N_8635);
or U8956 (N_8956,N_8643,N_8608);
xor U8957 (N_8957,N_8754,N_8797);
nand U8958 (N_8958,N_8660,N_8701);
nor U8959 (N_8959,N_8611,N_8651);
and U8960 (N_8960,N_8672,N_8792);
and U8961 (N_8961,N_8749,N_8746);
nor U8962 (N_8962,N_8737,N_8765);
nand U8963 (N_8963,N_8768,N_8789);
nand U8964 (N_8964,N_8738,N_8660);
and U8965 (N_8965,N_8765,N_8645);
and U8966 (N_8966,N_8780,N_8678);
nor U8967 (N_8967,N_8642,N_8619);
nor U8968 (N_8968,N_8751,N_8634);
and U8969 (N_8969,N_8652,N_8793);
nand U8970 (N_8970,N_8668,N_8615);
or U8971 (N_8971,N_8608,N_8764);
nand U8972 (N_8972,N_8601,N_8690);
nor U8973 (N_8973,N_8756,N_8752);
nor U8974 (N_8974,N_8641,N_8603);
or U8975 (N_8975,N_8617,N_8777);
nand U8976 (N_8976,N_8719,N_8672);
and U8977 (N_8977,N_8682,N_8719);
nand U8978 (N_8978,N_8677,N_8684);
nor U8979 (N_8979,N_8695,N_8613);
and U8980 (N_8980,N_8626,N_8630);
and U8981 (N_8981,N_8712,N_8693);
and U8982 (N_8982,N_8731,N_8675);
nor U8983 (N_8983,N_8657,N_8619);
and U8984 (N_8984,N_8628,N_8767);
or U8985 (N_8985,N_8753,N_8617);
nand U8986 (N_8986,N_8638,N_8655);
nand U8987 (N_8987,N_8625,N_8705);
nor U8988 (N_8988,N_8739,N_8765);
nor U8989 (N_8989,N_8630,N_8719);
or U8990 (N_8990,N_8779,N_8613);
xor U8991 (N_8991,N_8777,N_8788);
nor U8992 (N_8992,N_8790,N_8671);
nor U8993 (N_8993,N_8653,N_8790);
and U8994 (N_8994,N_8708,N_8702);
or U8995 (N_8995,N_8701,N_8684);
or U8996 (N_8996,N_8604,N_8735);
or U8997 (N_8997,N_8779,N_8644);
nor U8998 (N_8998,N_8799,N_8620);
nor U8999 (N_8999,N_8681,N_8677);
xor U9000 (N_9000,N_8971,N_8910);
nand U9001 (N_9001,N_8802,N_8830);
nor U9002 (N_9002,N_8805,N_8997);
and U9003 (N_9003,N_8930,N_8804);
nand U9004 (N_9004,N_8969,N_8922);
and U9005 (N_9005,N_8906,N_8845);
nand U9006 (N_9006,N_8945,N_8836);
nand U9007 (N_9007,N_8839,N_8868);
nand U9008 (N_9008,N_8957,N_8838);
nor U9009 (N_9009,N_8870,N_8886);
nor U9010 (N_9010,N_8872,N_8982);
nand U9011 (N_9011,N_8889,N_8819);
xor U9012 (N_9012,N_8935,N_8824);
nor U9013 (N_9013,N_8967,N_8818);
and U9014 (N_9014,N_8869,N_8899);
nand U9015 (N_9015,N_8865,N_8895);
nand U9016 (N_9016,N_8850,N_8987);
nand U9017 (N_9017,N_8811,N_8807);
and U9018 (N_9018,N_8923,N_8810);
nor U9019 (N_9019,N_8941,N_8874);
xor U9020 (N_9020,N_8988,N_8852);
and U9021 (N_9021,N_8927,N_8984);
or U9022 (N_9022,N_8973,N_8835);
nand U9023 (N_9023,N_8859,N_8902);
and U9024 (N_9024,N_8905,N_8933);
nand U9025 (N_9025,N_8834,N_8879);
or U9026 (N_9026,N_8904,N_8826);
xnor U9027 (N_9027,N_8908,N_8887);
nand U9028 (N_9028,N_8977,N_8832);
or U9029 (N_9029,N_8968,N_8803);
or U9030 (N_9030,N_8900,N_8955);
or U9031 (N_9031,N_8934,N_8885);
nor U9032 (N_9032,N_8847,N_8837);
nand U9033 (N_9033,N_8990,N_8989);
nor U9034 (N_9034,N_8858,N_8944);
nand U9035 (N_9035,N_8999,N_8862);
or U9036 (N_9036,N_8952,N_8806);
nor U9037 (N_9037,N_8809,N_8943);
nor U9038 (N_9038,N_8942,N_8820);
nor U9039 (N_9039,N_8972,N_8864);
nand U9040 (N_9040,N_8829,N_8841);
and U9041 (N_9041,N_8938,N_8926);
nand U9042 (N_9042,N_8947,N_8882);
or U9043 (N_9043,N_8893,N_8915);
nand U9044 (N_9044,N_8974,N_8961);
nand U9045 (N_9045,N_8929,N_8827);
and U9046 (N_9046,N_8979,N_8817);
nand U9047 (N_9047,N_8843,N_8815);
nor U9048 (N_9048,N_8833,N_8928);
xnor U9049 (N_9049,N_8995,N_8860);
or U9050 (N_9050,N_8821,N_8975);
nand U9051 (N_9051,N_8993,N_8966);
or U9052 (N_9052,N_8956,N_8800);
nor U9053 (N_9053,N_8994,N_8960);
nand U9054 (N_9054,N_8855,N_8891);
nand U9055 (N_9055,N_8996,N_8985);
and U9056 (N_9056,N_8937,N_8917);
or U9057 (N_9057,N_8953,N_8925);
nor U9058 (N_9058,N_8911,N_8921);
and U9059 (N_9059,N_8901,N_8876);
or U9060 (N_9060,N_8931,N_8914);
or U9061 (N_9061,N_8848,N_8894);
nor U9062 (N_9062,N_8962,N_8881);
and U9063 (N_9063,N_8981,N_8814);
and U9064 (N_9064,N_8842,N_8965);
nor U9065 (N_9065,N_8863,N_8907);
nand U9066 (N_9066,N_8861,N_8828);
and U9067 (N_9067,N_8880,N_8808);
xnor U9068 (N_9068,N_8875,N_8812);
nor U9069 (N_9069,N_8849,N_8897);
and U9070 (N_9070,N_8939,N_8948);
and U9071 (N_9071,N_8949,N_8853);
xor U9072 (N_9072,N_8963,N_8919);
nand U9073 (N_9073,N_8958,N_8884);
nand U9074 (N_9074,N_8983,N_8976);
nor U9075 (N_9075,N_8946,N_8970);
or U9076 (N_9076,N_8898,N_8823);
nand U9077 (N_9077,N_8959,N_8871);
nand U9078 (N_9078,N_8998,N_8825);
and U9079 (N_9079,N_8890,N_8896);
and U9080 (N_9080,N_8950,N_8840);
or U9081 (N_9081,N_8844,N_8932);
nand U9082 (N_9082,N_8918,N_8888);
xor U9083 (N_9083,N_8936,N_8992);
nand U9084 (N_9084,N_8846,N_8940);
or U9085 (N_9085,N_8856,N_8857);
nand U9086 (N_9086,N_8991,N_8916);
nor U9087 (N_9087,N_8831,N_8912);
and U9088 (N_9088,N_8903,N_8980);
nor U9089 (N_9089,N_8801,N_8867);
and U9090 (N_9090,N_8951,N_8854);
and U9091 (N_9091,N_8873,N_8964);
or U9092 (N_9092,N_8913,N_8822);
or U9093 (N_9093,N_8986,N_8924);
and U9094 (N_9094,N_8954,N_8892);
or U9095 (N_9095,N_8878,N_8920);
or U9096 (N_9096,N_8816,N_8978);
nand U9097 (N_9097,N_8851,N_8813);
nand U9098 (N_9098,N_8877,N_8866);
nand U9099 (N_9099,N_8883,N_8909);
xnor U9100 (N_9100,N_8883,N_8881);
nor U9101 (N_9101,N_8975,N_8883);
xor U9102 (N_9102,N_8920,N_8899);
xnor U9103 (N_9103,N_8910,N_8874);
or U9104 (N_9104,N_8928,N_8849);
nand U9105 (N_9105,N_8982,N_8995);
or U9106 (N_9106,N_8888,N_8967);
or U9107 (N_9107,N_8820,N_8933);
nand U9108 (N_9108,N_8831,N_8981);
nand U9109 (N_9109,N_8896,N_8934);
or U9110 (N_9110,N_8804,N_8884);
nand U9111 (N_9111,N_8976,N_8859);
nor U9112 (N_9112,N_8997,N_8884);
and U9113 (N_9113,N_8958,N_8877);
xor U9114 (N_9114,N_8850,N_8824);
nand U9115 (N_9115,N_8945,N_8924);
nor U9116 (N_9116,N_8980,N_8843);
nand U9117 (N_9117,N_8951,N_8808);
and U9118 (N_9118,N_8999,N_8845);
xnor U9119 (N_9119,N_8818,N_8835);
xnor U9120 (N_9120,N_8959,N_8985);
and U9121 (N_9121,N_8906,N_8880);
and U9122 (N_9122,N_8936,N_8821);
or U9123 (N_9123,N_8864,N_8932);
or U9124 (N_9124,N_8931,N_8858);
nand U9125 (N_9125,N_8998,N_8958);
nor U9126 (N_9126,N_8925,N_8923);
xor U9127 (N_9127,N_8999,N_8842);
xnor U9128 (N_9128,N_8860,N_8928);
nor U9129 (N_9129,N_8940,N_8804);
xor U9130 (N_9130,N_8932,N_8876);
and U9131 (N_9131,N_8832,N_8910);
nor U9132 (N_9132,N_8868,N_8892);
and U9133 (N_9133,N_8858,N_8860);
or U9134 (N_9134,N_8832,N_8971);
and U9135 (N_9135,N_8941,N_8974);
or U9136 (N_9136,N_8948,N_8938);
nand U9137 (N_9137,N_8998,N_8929);
nand U9138 (N_9138,N_8956,N_8871);
or U9139 (N_9139,N_8988,N_8954);
or U9140 (N_9140,N_8856,N_8982);
xor U9141 (N_9141,N_8989,N_8817);
or U9142 (N_9142,N_8810,N_8867);
and U9143 (N_9143,N_8894,N_8870);
and U9144 (N_9144,N_8856,N_8996);
and U9145 (N_9145,N_8938,N_8995);
and U9146 (N_9146,N_8840,N_8841);
or U9147 (N_9147,N_8832,N_8954);
and U9148 (N_9148,N_8874,N_8983);
or U9149 (N_9149,N_8858,N_8976);
and U9150 (N_9150,N_8905,N_8953);
nor U9151 (N_9151,N_8931,N_8843);
nand U9152 (N_9152,N_8827,N_8933);
nand U9153 (N_9153,N_8856,N_8893);
nand U9154 (N_9154,N_8810,N_8881);
and U9155 (N_9155,N_8974,N_8984);
nand U9156 (N_9156,N_8853,N_8882);
and U9157 (N_9157,N_8916,N_8923);
nor U9158 (N_9158,N_8928,N_8812);
and U9159 (N_9159,N_8911,N_8909);
or U9160 (N_9160,N_8883,N_8934);
and U9161 (N_9161,N_8819,N_8848);
nand U9162 (N_9162,N_8992,N_8938);
nor U9163 (N_9163,N_8847,N_8967);
nor U9164 (N_9164,N_8969,N_8828);
nand U9165 (N_9165,N_8966,N_8824);
nor U9166 (N_9166,N_8840,N_8906);
nor U9167 (N_9167,N_8986,N_8856);
or U9168 (N_9168,N_8919,N_8802);
and U9169 (N_9169,N_8936,N_8906);
nand U9170 (N_9170,N_8870,N_8914);
and U9171 (N_9171,N_8846,N_8804);
nor U9172 (N_9172,N_8872,N_8952);
xnor U9173 (N_9173,N_8897,N_8937);
or U9174 (N_9174,N_8900,N_8972);
and U9175 (N_9175,N_8827,N_8810);
nor U9176 (N_9176,N_8924,N_8928);
nor U9177 (N_9177,N_8993,N_8865);
nand U9178 (N_9178,N_8981,N_8821);
xnor U9179 (N_9179,N_8801,N_8934);
xnor U9180 (N_9180,N_8851,N_8914);
nand U9181 (N_9181,N_8884,N_8861);
or U9182 (N_9182,N_8913,N_8984);
nand U9183 (N_9183,N_8930,N_8855);
nor U9184 (N_9184,N_8873,N_8990);
nand U9185 (N_9185,N_8870,N_8912);
xnor U9186 (N_9186,N_8865,N_8899);
and U9187 (N_9187,N_8817,N_8939);
or U9188 (N_9188,N_8898,N_8902);
and U9189 (N_9189,N_8957,N_8897);
and U9190 (N_9190,N_8937,N_8832);
and U9191 (N_9191,N_8970,N_8968);
or U9192 (N_9192,N_8983,N_8826);
and U9193 (N_9193,N_8856,N_8934);
and U9194 (N_9194,N_8929,N_8943);
nand U9195 (N_9195,N_8800,N_8867);
nand U9196 (N_9196,N_8930,N_8957);
nand U9197 (N_9197,N_8978,N_8944);
and U9198 (N_9198,N_8966,N_8915);
and U9199 (N_9199,N_8860,N_8958);
or U9200 (N_9200,N_9081,N_9017);
nor U9201 (N_9201,N_9164,N_9026);
nand U9202 (N_9202,N_9188,N_9048);
nor U9203 (N_9203,N_9120,N_9143);
nor U9204 (N_9204,N_9049,N_9159);
nand U9205 (N_9205,N_9144,N_9077);
or U9206 (N_9206,N_9044,N_9157);
xor U9207 (N_9207,N_9066,N_9057);
nor U9208 (N_9208,N_9027,N_9196);
and U9209 (N_9209,N_9094,N_9113);
and U9210 (N_9210,N_9021,N_9198);
nor U9211 (N_9211,N_9147,N_9142);
or U9212 (N_9212,N_9080,N_9005);
or U9213 (N_9213,N_9031,N_9091);
and U9214 (N_9214,N_9001,N_9110);
or U9215 (N_9215,N_9176,N_9166);
nand U9216 (N_9216,N_9141,N_9010);
nor U9217 (N_9217,N_9009,N_9174);
nor U9218 (N_9218,N_9007,N_9030);
or U9219 (N_9219,N_9053,N_9107);
and U9220 (N_9220,N_9029,N_9032);
xnor U9221 (N_9221,N_9090,N_9151);
nor U9222 (N_9222,N_9126,N_9040);
or U9223 (N_9223,N_9050,N_9084);
nor U9224 (N_9224,N_9088,N_9075);
and U9225 (N_9225,N_9108,N_9193);
nor U9226 (N_9226,N_9002,N_9122);
nor U9227 (N_9227,N_9069,N_9158);
xnor U9228 (N_9228,N_9043,N_9004);
nor U9229 (N_9229,N_9095,N_9192);
and U9230 (N_9230,N_9112,N_9024);
nor U9231 (N_9231,N_9145,N_9167);
nor U9232 (N_9232,N_9102,N_9013);
and U9233 (N_9233,N_9056,N_9067);
nor U9234 (N_9234,N_9117,N_9187);
and U9235 (N_9235,N_9082,N_9123);
xnor U9236 (N_9236,N_9037,N_9152);
nor U9237 (N_9237,N_9129,N_9014);
and U9238 (N_9238,N_9153,N_9041);
nand U9239 (N_9239,N_9137,N_9184);
nor U9240 (N_9240,N_9058,N_9181);
or U9241 (N_9241,N_9051,N_9054);
nand U9242 (N_9242,N_9008,N_9149);
nand U9243 (N_9243,N_9180,N_9020);
nor U9244 (N_9244,N_9185,N_9097);
nor U9245 (N_9245,N_9130,N_9134);
nand U9246 (N_9246,N_9092,N_9072);
and U9247 (N_9247,N_9033,N_9006);
and U9248 (N_9248,N_9045,N_9019);
nor U9249 (N_9249,N_9173,N_9111);
nand U9250 (N_9250,N_9118,N_9087);
nand U9251 (N_9251,N_9105,N_9086);
nor U9252 (N_9252,N_9083,N_9100);
or U9253 (N_9253,N_9131,N_9018);
xnor U9254 (N_9254,N_9068,N_9012);
and U9255 (N_9255,N_9076,N_9127);
xnor U9256 (N_9256,N_9034,N_9154);
nor U9257 (N_9257,N_9064,N_9177);
nor U9258 (N_9258,N_9098,N_9052);
or U9259 (N_9259,N_9168,N_9150);
or U9260 (N_9260,N_9060,N_9119);
and U9261 (N_9261,N_9047,N_9035);
nor U9262 (N_9262,N_9073,N_9070);
nand U9263 (N_9263,N_9194,N_9063);
or U9264 (N_9264,N_9179,N_9025);
nor U9265 (N_9265,N_9162,N_9115);
nor U9266 (N_9266,N_9042,N_9161);
nor U9267 (N_9267,N_9078,N_9011);
or U9268 (N_9268,N_9038,N_9124);
or U9269 (N_9269,N_9135,N_9079);
nand U9270 (N_9270,N_9195,N_9023);
and U9271 (N_9271,N_9046,N_9140);
xor U9272 (N_9272,N_9104,N_9055);
nand U9273 (N_9273,N_9171,N_9106);
nor U9274 (N_9274,N_9085,N_9015);
and U9275 (N_9275,N_9103,N_9132);
nor U9276 (N_9276,N_9116,N_9114);
nand U9277 (N_9277,N_9125,N_9199);
or U9278 (N_9278,N_9071,N_9101);
nor U9279 (N_9279,N_9190,N_9039);
and U9280 (N_9280,N_9036,N_9128);
or U9281 (N_9281,N_9061,N_9028);
nor U9282 (N_9282,N_9093,N_9136);
nor U9283 (N_9283,N_9191,N_9109);
nand U9284 (N_9284,N_9089,N_9186);
and U9285 (N_9285,N_9156,N_9139);
or U9286 (N_9286,N_9155,N_9163);
nor U9287 (N_9287,N_9074,N_9133);
nand U9288 (N_9288,N_9096,N_9059);
or U9289 (N_9289,N_9000,N_9121);
nand U9290 (N_9290,N_9197,N_9178);
nor U9291 (N_9291,N_9003,N_9099);
and U9292 (N_9292,N_9189,N_9165);
and U9293 (N_9293,N_9138,N_9182);
and U9294 (N_9294,N_9169,N_9172);
nand U9295 (N_9295,N_9183,N_9022);
and U9296 (N_9296,N_9062,N_9148);
or U9297 (N_9297,N_9170,N_9175);
or U9298 (N_9298,N_9160,N_9016);
and U9299 (N_9299,N_9065,N_9146);
and U9300 (N_9300,N_9087,N_9091);
nand U9301 (N_9301,N_9067,N_9004);
and U9302 (N_9302,N_9113,N_9118);
xnor U9303 (N_9303,N_9143,N_9184);
and U9304 (N_9304,N_9054,N_9007);
and U9305 (N_9305,N_9125,N_9096);
nand U9306 (N_9306,N_9119,N_9181);
nor U9307 (N_9307,N_9043,N_9107);
and U9308 (N_9308,N_9076,N_9082);
nand U9309 (N_9309,N_9057,N_9134);
nor U9310 (N_9310,N_9103,N_9042);
and U9311 (N_9311,N_9071,N_9080);
or U9312 (N_9312,N_9183,N_9054);
nor U9313 (N_9313,N_9117,N_9190);
xnor U9314 (N_9314,N_9094,N_9017);
nand U9315 (N_9315,N_9116,N_9021);
nor U9316 (N_9316,N_9069,N_9141);
xnor U9317 (N_9317,N_9148,N_9141);
nor U9318 (N_9318,N_9035,N_9176);
xnor U9319 (N_9319,N_9072,N_9014);
or U9320 (N_9320,N_9100,N_9004);
nand U9321 (N_9321,N_9071,N_9092);
xnor U9322 (N_9322,N_9006,N_9169);
and U9323 (N_9323,N_9040,N_9162);
xor U9324 (N_9324,N_9079,N_9063);
nand U9325 (N_9325,N_9169,N_9113);
and U9326 (N_9326,N_9170,N_9191);
nor U9327 (N_9327,N_9169,N_9174);
nand U9328 (N_9328,N_9193,N_9196);
or U9329 (N_9329,N_9165,N_9008);
and U9330 (N_9330,N_9141,N_9007);
nor U9331 (N_9331,N_9183,N_9165);
nor U9332 (N_9332,N_9153,N_9199);
or U9333 (N_9333,N_9106,N_9137);
nand U9334 (N_9334,N_9036,N_9122);
and U9335 (N_9335,N_9057,N_9176);
nand U9336 (N_9336,N_9124,N_9011);
xor U9337 (N_9337,N_9159,N_9093);
nor U9338 (N_9338,N_9108,N_9175);
or U9339 (N_9339,N_9042,N_9061);
nor U9340 (N_9340,N_9056,N_9057);
or U9341 (N_9341,N_9166,N_9054);
and U9342 (N_9342,N_9008,N_9181);
nor U9343 (N_9343,N_9110,N_9000);
and U9344 (N_9344,N_9022,N_9135);
and U9345 (N_9345,N_9117,N_9087);
nand U9346 (N_9346,N_9167,N_9034);
nand U9347 (N_9347,N_9073,N_9194);
or U9348 (N_9348,N_9152,N_9052);
and U9349 (N_9349,N_9122,N_9059);
or U9350 (N_9350,N_9079,N_9085);
and U9351 (N_9351,N_9072,N_9038);
or U9352 (N_9352,N_9109,N_9086);
or U9353 (N_9353,N_9057,N_9084);
nand U9354 (N_9354,N_9061,N_9179);
nor U9355 (N_9355,N_9191,N_9198);
nor U9356 (N_9356,N_9153,N_9104);
and U9357 (N_9357,N_9023,N_9118);
and U9358 (N_9358,N_9049,N_9111);
and U9359 (N_9359,N_9019,N_9174);
and U9360 (N_9360,N_9005,N_9186);
xnor U9361 (N_9361,N_9044,N_9166);
or U9362 (N_9362,N_9017,N_9012);
and U9363 (N_9363,N_9006,N_9148);
xor U9364 (N_9364,N_9153,N_9176);
or U9365 (N_9365,N_9086,N_9146);
and U9366 (N_9366,N_9175,N_9121);
nand U9367 (N_9367,N_9117,N_9098);
and U9368 (N_9368,N_9149,N_9003);
and U9369 (N_9369,N_9018,N_9034);
or U9370 (N_9370,N_9136,N_9004);
or U9371 (N_9371,N_9188,N_9108);
nor U9372 (N_9372,N_9034,N_9193);
or U9373 (N_9373,N_9122,N_9034);
or U9374 (N_9374,N_9015,N_9188);
nand U9375 (N_9375,N_9052,N_9037);
nor U9376 (N_9376,N_9119,N_9073);
and U9377 (N_9377,N_9014,N_9069);
and U9378 (N_9378,N_9027,N_9173);
nand U9379 (N_9379,N_9033,N_9119);
and U9380 (N_9380,N_9067,N_9177);
nand U9381 (N_9381,N_9070,N_9130);
and U9382 (N_9382,N_9033,N_9039);
nor U9383 (N_9383,N_9133,N_9138);
xnor U9384 (N_9384,N_9076,N_9113);
xor U9385 (N_9385,N_9106,N_9145);
or U9386 (N_9386,N_9017,N_9023);
xor U9387 (N_9387,N_9018,N_9045);
nor U9388 (N_9388,N_9093,N_9023);
and U9389 (N_9389,N_9052,N_9187);
and U9390 (N_9390,N_9002,N_9047);
nor U9391 (N_9391,N_9098,N_9196);
nand U9392 (N_9392,N_9112,N_9175);
nor U9393 (N_9393,N_9135,N_9044);
nor U9394 (N_9394,N_9077,N_9023);
or U9395 (N_9395,N_9004,N_9148);
or U9396 (N_9396,N_9007,N_9147);
xor U9397 (N_9397,N_9084,N_9169);
or U9398 (N_9398,N_9153,N_9017);
nor U9399 (N_9399,N_9192,N_9178);
nand U9400 (N_9400,N_9385,N_9344);
nand U9401 (N_9401,N_9267,N_9346);
and U9402 (N_9402,N_9308,N_9348);
and U9403 (N_9403,N_9256,N_9350);
nor U9404 (N_9404,N_9314,N_9264);
nand U9405 (N_9405,N_9363,N_9380);
nor U9406 (N_9406,N_9337,N_9202);
or U9407 (N_9407,N_9396,N_9250);
or U9408 (N_9408,N_9229,N_9210);
nand U9409 (N_9409,N_9276,N_9281);
xnor U9410 (N_9410,N_9374,N_9340);
nand U9411 (N_9411,N_9355,N_9395);
and U9412 (N_9412,N_9296,N_9326);
nand U9413 (N_9413,N_9241,N_9384);
or U9414 (N_9414,N_9323,N_9317);
xor U9415 (N_9415,N_9213,N_9211);
nor U9416 (N_9416,N_9322,N_9273);
or U9417 (N_9417,N_9358,N_9299);
nor U9418 (N_9418,N_9312,N_9215);
nor U9419 (N_9419,N_9290,N_9260);
nand U9420 (N_9420,N_9230,N_9310);
nand U9421 (N_9421,N_9291,N_9367);
and U9422 (N_9422,N_9225,N_9368);
xnor U9423 (N_9423,N_9237,N_9399);
and U9424 (N_9424,N_9372,N_9223);
and U9425 (N_9425,N_9268,N_9284);
nand U9426 (N_9426,N_9239,N_9304);
and U9427 (N_9427,N_9366,N_9219);
nand U9428 (N_9428,N_9297,N_9245);
nor U9429 (N_9429,N_9379,N_9342);
or U9430 (N_9430,N_9364,N_9218);
nand U9431 (N_9431,N_9324,N_9371);
or U9432 (N_9432,N_9391,N_9394);
or U9433 (N_9433,N_9294,N_9327);
and U9434 (N_9434,N_9339,N_9243);
nand U9435 (N_9435,N_9228,N_9397);
or U9436 (N_9436,N_9365,N_9234);
nor U9437 (N_9437,N_9361,N_9388);
xor U9438 (N_9438,N_9277,N_9201);
nor U9439 (N_9439,N_9336,N_9266);
or U9440 (N_9440,N_9376,N_9295);
or U9441 (N_9441,N_9206,N_9207);
xor U9442 (N_9442,N_9216,N_9224);
nor U9443 (N_9443,N_9261,N_9381);
nor U9444 (N_9444,N_9231,N_9360);
and U9445 (N_9445,N_9343,N_9349);
nand U9446 (N_9446,N_9265,N_9298);
nor U9447 (N_9447,N_9378,N_9254);
or U9448 (N_9448,N_9209,N_9272);
and U9449 (N_9449,N_9249,N_9354);
nand U9450 (N_9450,N_9329,N_9393);
nor U9451 (N_9451,N_9301,N_9259);
nand U9452 (N_9452,N_9278,N_9258);
or U9453 (N_9453,N_9247,N_9271);
nand U9454 (N_9454,N_9370,N_9244);
xnor U9455 (N_9455,N_9377,N_9341);
nand U9456 (N_9456,N_9214,N_9300);
and U9457 (N_9457,N_9220,N_9282);
xor U9458 (N_9458,N_9316,N_9319);
nor U9459 (N_9459,N_9383,N_9270);
or U9460 (N_9460,N_9352,N_9217);
or U9461 (N_9461,N_9307,N_9351);
or U9462 (N_9462,N_9212,N_9382);
nor U9463 (N_9463,N_9200,N_9233);
nor U9464 (N_9464,N_9204,N_9335);
nand U9465 (N_9465,N_9232,N_9288);
nor U9466 (N_9466,N_9373,N_9328);
xnor U9467 (N_9467,N_9309,N_9362);
nand U9468 (N_9468,N_9305,N_9255);
or U9469 (N_9469,N_9353,N_9280);
or U9470 (N_9470,N_9246,N_9285);
or U9471 (N_9471,N_9257,N_9248);
or U9472 (N_9472,N_9386,N_9331);
and U9473 (N_9473,N_9292,N_9347);
nor U9474 (N_9474,N_9293,N_9251);
nand U9475 (N_9475,N_9325,N_9375);
xor U9476 (N_9476,N_9390,N_9315);
nor U9477 (N_9477,N_9226,N_9238);
nor U9478 (N_9478,N_9221,N_9369);
nand U9479 (N_9479,N_9227,N_9289);
and U9480 (N_9480,N_9392,N_9313);
xor U9481 (N_9481,N_9240,N_9302);
or U9482 (N_9482,N_9274,N_9303);
nand U9483 (N_9483,N_9275,N_9252);
nand U9484 (N_9484,N_9203,N_9332);
nor U9485 (N_9485,N_9287,N_9286);
or U9486 (N_9486,N_9262,N_9345);
nor U9487 (N_9487,N_9205,N_9389);
or U9488 (N_9488,N_9208,N_9253);
and U9489 (N_9489,N_9235,N_9236);
and U9490 (N_9490,N_9222,N_9359);
or U9491 (N_9491,N_9356,N_9357);
nand U9492 (N_9492,N_9263,N_9320);
nor U9493 (N_9493,N_9306,N_9330);
nand U9494 (N_9494,N_9321,N_9311);
xor U9495 (N_9495,N_9338,N_9269);
nand U9496 (N_9496,N_9318,N_9398);
and U9497 (N_9497,N_9334,N_9242);
xor U9498 (N_9498,N_9387,N_9279);
nor U9499 (N_9499,N_9283,N_9333);
and U9500 (N_9500,N_9301,N_9225);
xor U9501 (N_9501,N_9302,N_9275);
and U9502 (N_9502,N_9242,N_9393);
and U9503 (N_9503,N_9245,N_9399);
and U9504 (N_9504,N_9397,N_9296);
nand U9505 (N_9505,N_9300,N_9324);
nand U9506 (N_9506,N_9255,N_9278);
xor U9507 (N_9507,N_9277,N_9302);
or U9508 (N_9508,N_9241,N_9361);
nor U9509 (N_9509,N_9344,N_9207);
nand U9510 (N_9510,N_9326,N_9351);
or U9511 (N_9511,N_9202,N_9336);
nand U9512 (N_9512,N_9245,N_9327);
nor U9513 (N_9513,N_9352,N_9333);
and U9514 (N_9514,N_9202,N_9264);
nor U9515 (N_9515,N_9226,N_9272);
and U9516 (N_9516,N_9327,N_9222);
or U9517 (N_9517,N_9292,N_9341);
or U9518 (N_9518,N_9373,N_9340);
or U9519 (N_9519,N_9355,N_9302);
nor U9520 (N_9520,N_9221,N_9356);
or U9521 (N_9521,N_9229,N_9230);
xnor U9522 (N_9522,N_9379,N_9271);
or U9523 (N_9523,N_9219,N_9303);
and U9524 (N_9524,N_9367,N_9339);
xor U9525 (N_9525,N_9206,N_9286);
nand U9526 (N_9526,N_9365,N_9392);
nor U9527 (N_9527,N_9356,N_9327);
nand U9528 (N_9528,N_9368,N_9350);
nand U9529 (N_9529,N_9232,N_9234);
nand U9530 (N_9530,N_9252,N_9342);
or U9531 (N_9531,N_9387,N_9234);
nor U9532 (N_9532,N_9303,N_9384);
nor U9533 (N_9533,N_9275,N_9265);
nor U9534 (N_9534,N_9363,N_9377);
and U9535 (N_9535,N_9320,N_9272);
and U9536 (N_9536,N_9292,N_9288);
nor U9537 (N_9537,N_9304,N_9390);
xor U9538 (N_9538,N_9275,N_9208);
nor U9539 (N_9539,N_9382,N_9237);
xnor U9540 (N_9540,N_9307,N_9242);
nor U9541 (N_9541,N_9253,N_9359);
xnor U9542 (N_9542,N_9307,N_9359);
and U9543 (N_9543,N_9333,N_9266);
nand U9544 (N_9544,N_9289,N_9381);
or U9545 (N_9545,N_9274,N_9377);
or U9546 (N_9546,N_9331,N_9244);
nand U9547 (N_9547,N_9211,N_9278);
xor U9548 (N_9548,N_9223,N_9332);
nor U9549 (N_9549,N_9287,N_9201);
nand U9550 (N_9550,N_9326,N_9290);
and U9551 (N_9551,N_9304,N_9312);
or U9552 (N_9552,N_9297,N_9350);
or U9553 (N_9553,N_9334,N_9282);
xor U9554 (N_9554,N_9251,N_9305);
and U9555 (N_9555,N_9331,N_9316);
or U9556 (N_9556,N_9300,N_9243);
nand U9557 (N_9557,N_9308,N_9366);
nor U9558 (N_9558,N_9336,N_9330);
nand U9559 (N_9559,N_9237,N_9209);
or U9560 (N_9560,N_9362,N_9350);
xnor U9561 (N_9561,N_9246,N_9264);
xnor U9562 (N_9562,N_9384,N_9211);
nor U9563 (N_9563,N_9253,N_9357);
or U9564 (N_9564,N_9382,N_9296);
nor U9565 (N_9565,N_9250,N_9350);
nor U9566 (N_9566,N_9217,N_9309);
or U9567 (N_9567,N_9332,N_9275);
nand U9568 (N_9568,N_9263,N_9348);
or U9569 (N_9569,N_9236,N_9251);
or U9570 (N_9570,N_9341,N_9295);
and U9571 (N_9571,N_9258,N_9368);
nor U9572 (N_9572,N_9325,N_9215);
and U9573 (N_9573,N_9370,N_9226);
nor U9574 (N_9574,N_9316,N_9271);
nand U9575 (N_9575,N_9353,N_9372);
nor U9576 (N_9576,N_9389,N_9361);
nor U9577 (N_9577,N_9240,N_9207);
and U9578 (N_9578,N_9235,N_9211);
xnor U9579 (N_9579,N_9228,N_9364);
and U9580 (N_9580,N_9370,N_9345);
nor U9581 (N_9581,N_9330,N_9284);
nor U9582 (N_9582,N_9293,N_9381);
nor U9583 (N_9583,N_9348,N_9273);
and U9584 (N_9584,N_9218,N_9347);
and U9585 (N_9585,N_9240,N_9307);
nor U9586 (N_9586,N_9386,N_9362);
and U9587 (N_9587,N_9306,N_9305);
and U9588 (N_9588,N_9366,N_9305);
or U9589 (N_9589,N_9312,N_9285);
nand U9590 (N_9590,N_9291,N_9395);
or U9591 (N_9591,N_9342,N_9357);
nand U9592 (N_9592,N_9243,N_9209);
nand U9593 (N_9593,N_9360,N_9372);
and U9594 (N_9594,N_9286,N_9315);
nand U9595 (N_9595,N_9397,N_9251);
nand U9596 (N_9596,N_9264,N_9388);
nor U9597 (N_9597,N_9391,N_9223);
xor U9598 (N_9598,N_9233,N_9257);
nor U9599 (N_9599,N_9200,N_9302);
and U9600 (N_9600,N_9494,N_9515);
nor U9601 (N_9601,N_9434,N_9512);
or U9602 (N_9602,N_9590,N_9440);
nor U9603 (N_9603,N_9539,N_9407);
nor U9604 (N_9604,N_9546,N_9487);
or U9605 (N_9605,N_9429,N_9540);
nor U9606 (N_9606,N_9475,N_9542);
or U9607 (N_9607,N_9545,N_9597);
nor U9608 (N_9608,N_9502,N_9519);
nor U9609 (N_9609,N_9451,N_9506);
nand U9610 (N_9610,N_9406,N_9568);
xor U9611 (N_9611,N_9521,N_9589);
nor U9612 (N_9612,N_9446,N_9403);
nand U9613 (N_9613,N_9586,N_9432);
nand U9614 (N_9614,N_9437,N_9495);
and U9615 (N_9615,N_9458,N_9573);
and U9616 (N_9616,N_9491,N_9579);
nor U9617 (N_9617,N_9464,N_9584);
xor U9618 (N_9618,N_9524,N_9538);
nand U9619 (N_9619,N_9427,N_9501);
and U9620 (N_9620,N_9505,N_9588);
nand U9621 (N_9621,N_9415,N_9566);
nand U9622 (N_9622,N_9490,N_9469);
nor U9623 (N_9623,N_9441,N_9422);
xnor U9624 (N_9624,N_9599,N_9531);
or U9625 (N_9625,N_9553,N_9509);
nand U9626 (N_9626,N_9503,N_9517);
nor U9627 (N_9627,N_9444,N_9547);
nor U9628 (N_9628,N_9536,N_9510);
or U9629 (N_9629,N_9466,N_9592);
or U9630 (N_9630,N_9452,N_9420);
and U9631 (N_9631,N_9497,N_9535);
and U9632 (N_9632,N_9496,N_9480);
xor U9633 (N_9633,N_9523,N_9468);
nand U9634 (N_9634,N_9543,N_9555);
and U9635 (N_9635,N_9526,N_9433);
or U9636 (N_9636,N_9426,N_9504);
nand U9637 (N_9637,N_9520,N_9447);
xnor U9638 (N_9638,N_9569,N_9511);
nand U9639 (N_9639,N_9402,N_9529);
and U9640 (N_9640,N_9565,N_9443);
nor U9641 (N_9641,N_9486,N_9435);
nand U9642 (N_9642,N_9476,N_9500);
and U9643 (N_9643,N_9591,N_9474);
nand U9644 (N_9644,N_9561,N_9533);
and U9645 (N_9645,N_9544,N_9598);
nor U9646 (N_9646,N_9488,N_9405);
or U9647 (N_9647,N_9404,N_9562);
nand U9648 (N_9648,N_9493,N_9513);
xor U9649 (N_9649,N_9408,N_9551);
and U9650 (N_9650,N_9552,N_9449);
nor U9651 (N_9651,N_9414,N_9525);
or U9652 (N_9652,N_9456,N_9518);
xnor U9653 (N_9653,N_9499,N_9549);
or U9654 (N_9654,N_9582,N_9438);
nand U9655 (N_9655,N_9537,N_9465);
or U9656 (N_9656,N_9459,N_9571);
xnor U9657 (N_9657,N_9574,N_9467);
nor U9658 (N_9658,N_9460,N_9522);
nand U9659 (N_9659,N_9445,N_9558);
or U9660 (N_9660,N_9548,N_9481);
or U9661 (N_9661,N_9471,N_9457);
or U9662 (N_9662,N_9484,N_9419);
nand U9663 (N_9663,N_9416,N_9430);
or U9664 (N_9664,N_9470,N_9479);
and U9665 (N_9665,N_9514,N_9516);
nor U9666 (N_9666,N_9563,N_9489);
nand U9667 (N_9667,N_9477,N_9485);
nor U9668 (N_9668,N_9483,N_9428);
and U9669 (N_9669,N_9560,N_9556);
nand U9670 (N_9670,N_9559,N_9448);
or U9671 (N_9671,N_9530,N_9575);
and U9672 (N_9672,N_9436,N_9594);
nor U9673 (N_9673,N_9508,N_9424);
nor U9674 (N_9674,N_9528,N_9410);
or U9675 (N_9675,N_9567,N_9431);
and U9676 (N_9676,N_9576,N_9541);
nor U9677 (N_9677,N_9409,N_9564);
and U9678 (N_9678,N_9412,N_9507);
or U9679 (N_9679,N_9577,N_9595);
xnor U9680 (N_9680,N_9411,N_9570);
and U9681 (N_9681,N_9482,N_9442);
nor U9682 (N_9682,N_9425,N_9421);
nor U9683 (N_9683,N_9473,N_9401);
nor U9684 (N_9684,N_9461,N_9596);
or U9685 (N_9685,N_9532,N_9572);
or U9686 (N_9686,N_9413,N_9554);
and U9687 (N_9687,N_9534,N_9455);
nand U9688 (N_9688,N_9581,N_9557);
and U9689 (N_9689,N_9439,N_9593);
nor U9690 (N_9690,N_9587,N_9453);
nand U9691 (N_9691,N_9418,N_9585);
or U9692 (N_9692,N_9498,N_9423);
nand U9693 (N_9693,N_9450,N_9463);
nand U9694 (N_9694,N_9578,N_9492);
nand U9695 (N_9695,N_9472,N_9527);
and U9696 (N_9696,N_9462,N_9583);
or U9697 (N_9697,N_9400,N_9454);
or U9698 (N_9698,N_9478,N_9580);
nand U9699 (N_9699,N_9550,N_9417);
or U9700 (N_9700,N_9500,N_9560);
xor U9701 (N_9701,N_9476,N_9454);
nand U9702 (N_9702,N_9441,N_9504);
or U9703 (N_9703,N_9593,N_9402);
nor U9704 (N_9704,N_9599,N_9497);
and U9705 (N_9705,N_9439,N_9471);
nor U9706 (N_9706,N_9471,N_9480);
xor U9707 (N_9707,N_9443,N_9559);
and U9708 (N_9708,N_9536,N_9534);
nand U9709 (N_9709,N_9560,N_9415);
nor U9710 (N_9710,N_9460,N_9468);
or U9711 (N_9711,N_9504,N_9516);
nand U9712 (N_9712,N_9573,N_9525);
nor U9713 (N_9713,N_9419,N_9426);
nand U9714 (N_9714,N_9590,N_9443);
nor U9715 (N_9715,N_9561,N_9579);
or U9716 (N_9716,N_9430,N_9532);
nand U9717 (N_9717,N_9412,N_9502);
nand U9718 (N_9718,N_9448,N_9566);
nor U9719 (N_9719,N_9582,N_9462);
nand U9720 (N_9720,N_9502,N_9596);
and U9721 (N_9721,N_9410,N_9599);
and U9722 (N_9722,N_9594,N_9430);
or U9723 (N_9723,N_9542,N_9485);
nand U9724 (N_9724,N_9589,N_9518);
and U9725 (N_9725,N_9421,N_9511);
and U9726 (N_9726,N_9517,N_9511);
nor U9727 (N_9727,N_9501,N_9452);
xnor U9728 (N_9728,N_9555,N_9447);
nor U9729 (N_9729,N_9448,N_9402);
or U9730 (N_9730,N_9511,N_9578);
nor U9731 (N_9731,N_9425,N_9548);
nor U9732 (N_9732,N_9495,N_9481);
and U9733 (N_9733,N_9470,N_9516);
nor U9734 (N_9734,N_9547,N_9503);
or U9735 (N_9735,N_9480,N_9560);
or U9736 (N_9736,N_9558,N_9514);
nor U9737 (N_9737,N_9410,N_9448);
nand U9738 (N_9738,N_9554,N_9464);
nor U9739 (N_9739,N_9418,N_9416);
or U9740 (N_9740,N_9414,N_9446);
nand U9741 (N_9741,N_9412,N_9403);
or U9742 (N_9742,N_9438,N_9463);
nand U9743 (N_9743,N_9496,N_9424);
xnor U9744 (N_9744,N_9508,N_9549);
nand U9745 (N_9745,N_9401,N_9412);
nor U9746 (N_9746,N_9520,N_9406);
nor U9747 (N_9747,N_9531,N_9486);
nand U9748 (N_9748,N_9451,N_9459);
nor U9749 (N_9749,N_9423,N_9480);
or U9750 (N_9750,N_9593,N_9523);
nor U9751 (N_9751,N_9500,N_9526);
or U9752 (N_9752,N_9504,N_9436);
nor U9753 (N_9753,N_9565,N_9505);
or U9754 (N_9754,N_9559,N_9564);
xor U9755 (N_9755,N_9599,N_9500);
nor U9756 (N_9756,N_9499,N_9472);
and U9757 (N_9757,N_9546,N_9503);
and U9758 (N_9758,N_9460,N_9487);
nand U9759 (N_9759,N_9528,N_9484);
or U9760 (N_9760,N_9442,N_9530);
or U9761 (N_9761,N_9550,N_9408);
and U9762 (N_9762,N_9429,N_9532);
and U9763 (N_9763,N_9442,N_9457);
nor U9764 (N_9764,N_9492,N_9595);
or U9765 (N_9765,N_9591,N_9437);
nor U9766 (N_9766,N_9549,N_9550);
nor U9767 (N_9767,N_9427,N_9475);
and U9768 (N_9768,N_9509,N_9561);
xnor U9769 (N_9769,N_9466,N_9465);
nor U9770 (N_9770,N_9448,N_9501);
nand U9771 (N_9771,N_9481,N_9556);
nand U9772 (N_9772,N_9589,N_9581);
or U9773 (N_9773,N_9479,N_9446);
nand U9774 (N_9774,N_9429,N_9517);
xnor U9775 (N_9775,N_9416,N_9591);
nand U9776 (N_9776,N_9422,N_9462);
and U9777 (N_9777,N_9414,N_9596);
xor U9778 (N_9778,N_9432,N_9562);
nor U9779 (N_9779,N_9482,N_9472);
or U9780 (N_9780,N_9562,N_9566);
and U9781 (N_9781,N_9556,N_9407);
nor U9782 (N_9782,N_9543,N_9441);
and U9783 (N_9783,N_9575,N_9561);
or U9784 (N_9784,N_9441,N_9583);
or U9785 (N_9785,N_9414,N_9504);
or U9786 (N_9786,N_9408,N_9570);
nand U9787 (N_9787,N_9439,N_9546);
and U9788 (N_9788,N_9442,N_9518);
or U9789 (N_9789,N_9569,N_9449);
nand U9790 (N_9790,N_9544,N_9570);
nand U9791 (N_9791,N_9560,N_9566);
and U9792 (N_9792,N_9585,N_9456);
nand U9793 (N_9793,N_9499,N_9531);
nor U9794 (N_9794,N_9505,N_9589);
xor U9795 (N_9795,N_9435,N_9532);
nor U9796 (N_9796,N_9575,N_9404);
nor U9797 (N_9797,N_9425,N_9555);
and U9798 (N_9798,N_9474,N_9593);
and U9799 (N_9799,N_9585,N_9522);
nand U9800 (N_9800,N_9629,N_9703);
xor U9801 (N_9801,N_9739,N_9698);
nand U9802 (N_9802,N_9697,N_9656);
nand U9803 (N_9803,N_9652,N_9760);
xnor U9804 (N_9804,N_9686,N_9687);
nor U9805 (N_9805,N_9708,N_9669);
or U9806 (N_9806,N_9617,N_9770);
or U9807 (N_9807,N_9619,N_9728);
or U9808 (N_9808,N_9663,N_9717);
or U9809 (N_9809,N_9632,N_9718);
nor U9810 (N_9810,N_9790,N_9620);
or U9811 (N_9811,N_9778,N_9658);
or U9812 (N_9812,N_9692,N_9768);
or U9813 (N_9813,N_9779,N_9773);
and U9814 (N_9814,N_9646,N_9751);
and U9815 (N_9815,N_9732,N_9650);
nor U9816 (N_9816,N_9794,N_9747);
xor U9817 (N_9817,N_9631,N_9613);
and U9818 (N_9818,N_9608,N_9782);
or U9819 (N_9819,N_9735,N_9769);
nand U9820 (N_9820,N_9705,N_9796);
nor U9821 (N_9821,N_9731,N_9603);
xnor U9822 (N_9822,N_9682,N_9737);
nand U9823 (N_9823,N_9727,N_9738);
or U9824 (N_9824,N_9721,N_9635);
or U9825 (N_9825,N_9621,N_9733);
or U9826 (N_9826,N_9634,N_9657);
or U9827 (N_9827,N_9762,N_9606);
nand U9828 (N_9828,N_9798,N_9676);
and U9829 (N_9829,N_9765,N_9683);
and U9830 (N_9830,N_9622,N_9624);
or U9831 (N_9831,N_9653,N_9761);
or U9832 (N_9832,N_9645,N_9766);
nor U9833 (N_9833,N_9699,N_9701);
nor U9834 (N_9834,N_9616,N_9660);
or U9835 (N_9835,N_9786,N_9771);
nor U9836 (N_9836,N_9605,N_9655);
and U9837 (N_9837,N_9710,N_9795);
xnor U9838 (N_9838,N_9691,N_9665);
xor U9839 (N_9839,N_9763,N_9681);
xnor U9840 (N_9840,N_9659,N_9675);
and U9841 (N_9841,N_9723,N_9730);
nand U9842 (N_9842,N_9636,N_9651);
and U9843 (N_9843,N_9623,N_9767);
and U9844 (N_9844,N_9758,N_9734);
xor U9845 (N_9845,N_9744,N_9772);
and U9846 (N_9846,N_9673,N_9670);
nand U9847 (N_9847,N_9604,N_9618);
nand U9848 (N_9848,N_9639,N_9764);
xor U9849 (N_9849,N_9776,N_9746);
or U9850 (N_9850,N_9693,N_9700);
and U9851 (N_9851,N_9695,N_9724);
nor U9852 (N_9852,N_9680,N_9647);
nor U9853 (N_9853,N_9668,N_9677);
nand U9854 (N_9854,N_9713,N_9788);
nand U9855 (N_9855,N_9661,N_9679);
nor U9856 (N_9856,N_9748,N_9667);
nor U9857 (N_9857,N_9637,N_9614);
xnor U9858 (N_9858,N_9704,N_9783);
and U9859 (N_9859,N_9757,N_9789);
or U9860 (N_9860,N_9642,N_9745);
or U9861 (N_9861,N_9654,N_9644);
and U9862 (N_9862,N_9671,N_9684);
nand U9863 (N_9863,N_9602,N_9662);
or U9864 (N_9864,N_9752,N_9706);
nand U9865 (N_9865,N_9689,N_9611);
or U9866 (N_9866,N_9781,N_9702);
or U9867 (N_9867,N_9774,N_9600);
and U9868 (N_9868,N_9780,N_9715);
and U9869 (N_9869,N_9685,N_9719);
nor U9870 (N_9870,N_9625,N_9643);
and U9871 (N_9871,N_9750,N_9787);
nand U9872 (N_9872,N_9609,N_9775);
or U9873 (N_9873,N_9799,N_9690);
and U9874 (N_9874,N_9694,N_9729);
nand U9875 (N_9875,N_9714,N_9688);
or U9876 (N_9876,N_9696,N_9664);
nor U9877 (N_9877,N_9607,N_9601);
nand U9878 (N_9878,N_9736,N_9612);
or U9879 (N_9879,N_9797,N_9638);
xnor U9880 (N_9880,N_9626,N_9674);
and U9881 (N_9881,N_9672,N_9630);
xor U9882 (N_9882,N_9720,N_9793);
nor U9883 (N_9883,N_9707,N_9755);
and U9884 (N_9884,N_9726,N_9742);
and U9885 (N_9885,N_9615,N_9756);
or U9886 (N_9886,N_9784,N_9716);
xor U9887 (N_9887,N_9759,N_9633);
and U9888 (N_9888,N_9666,N_9648);
nor U9889 (N_9889,N_9722,N_9649);
nor U9890 (N_9890,N_9792,N_9678);
nor U9891 (N_9891,N_9628,N_9743);
and U9892 (N_9892,N_9740,N_9711);
and U9893 (N_9893,N_9709,N_9753);
or U9894 (N_9894,N_9610,N_9791);
or U9895 (N_9895,N_9741,N_9640);
and U9896 (N_9896,N_9725,N_9754);
or U9897 (N_9897,N_9749,N_9785);
nand U9898 (N_9898,N_9627,N_9777);
nor U9899 (N_9899,N_9712,N_9641);
nor U9900 (N_9900,N_9734,N_9665);
and U9901 (N_9901,N_9606,N_9691);
nor U9902 (N_9902,N_9727,N_9777);
nand U9903 (N_9903,N_9600,N_9729);
nor U9904 (N_9904,N_9602,N_9624);
nand U9905 (N_9905,N_9768,N_9729);
and U9906 (N_9906,N_9705,N_9620);
xnor U9907 (N_9907,N_9632,N_9731);
nand U9908 (N_9908,N_9645,N_9688);
xor U9909 (N_9909,N_9730,N_9654);
nand U9910 (N_9910,N_9776,N_9744);
nor U9911 (N_9911,N_9724,N_9743);
and U9912 (N_9912,N_9758,N_9774);
and U9913 (N_9913,N_9743,N_9792);
and U9914 (N_9914,N_9681,N_9740);
and U9915 (N_9915,N_9727,N_9634);
or U9916 (N_9916,N_9783,N_9754);
nand U9917 (N_9917,N_9703,N_9610);
and U9918 (N_9918,N_9664,N_9679);
nor U9919 (N_9919,N_9731,N_9665);
or U9920 (N_9920,N_9740,N_9789);
and U9921 (N_9921,N_9747,N_9770);
nand U9922 (N_9922,N_9660,N_9649);
or U9923 (N_9923,N_9714,N_9654);
nor U9924 (N_9924,N_9617,N_9663);
and U9925 (N_9925,N_9790,N_9727);
or U9926 (N_9926,N_9614,N_9663);
nand U9927 (N_9927,N_9675,N_9733);
and U9928 (N_9928,N_9748,N_9708);
and U9929 (N_9929,N_9706,N_9601);
or U9930 (N_9930,N_9783,N_9639);
or U9931 (N_9931,N_9602,N_9674);
nor U9932 (N_9932,N_9705,N_9649);
nand U9933 (N_9933,N_9649,N_9726);
nand U9934 (N_9934,N_9734,N_9705);
or U9935 (N_9935,N_9753,N_9623);
or U9936 (N_9936,N_9764,N_9727);
and U9937 (N_9937,N_9684,N_9645);
nor U9938 (N_9938,N_9621,N_9783);
nand U9939 (N_9939,N_9749,N_9684);
and U9940 (N_9940,N_9691,N_9647);
nor U9941 (N_9941,N_9696,N_9610);
or U9942 (N_9942,N_9624,N_9770);
nand U9943 (N_9943,N_9682,N_9752);
nor U9944 (N_9944,N_9784,N_9758);
nor U9945 (N_9945,N_9672,N_9729);
and U9946 (N_9946,N_9749,N_9759);
nand U9947 (N_9947,N_9684,N_9652);
and U9948 (N_9948,N_9798,N_9623);
xor U9949 (N_9949,N_9780,N_9603);
or U9950 (N_9950,N_9733,N_9681);
xnor U9951 (N_9951,N_9772,N_9780);
and U9952 (N_9952,N_9664,N_9759);
nand U9953 (N_9953,N_9612,N_9709);
nand U9954 (N_9954,N_9750,N_9709);
xnor U9955 (N_9955,N_9713,N_9778);
nand U9956 (N_9956,N_9659,N_9669);
and U9957 (N_9957,N_9673,N_9724);
and U9958 (N_9958,N_9707,N_9740);
xnor U9959 (N_9959,N_9691,N_9728);
or U9960 (N_9960,N_9655,N_9716);
nor U9961 (N_9961,N_9686,N_9759);
xor U9962 (N_9962,N_9674,N_9667);
and U9963 (N_9963,N_9749,N_9656);
xnor U9964 (N_9964,N_9636,N_9630);
and U9965 (N_9965,N_9781,N_9629);
nor U9966 (N_9966,N_9707,N_9663);
nand U9967 (N_9967,N_9799,N_9662);
and U9968 (N_9968,N_9612,N_9644);
nand U9969 (N_9969,N_9714,N_9798);
nand U9970 (N_9970,N_9695,N_9660);
or U9971 (N_9971,N_9767,N_9676);
xnor U9972 (N_9972,N_9639,N_9636);
nand U9973 (N_9973,N_9774,N_9748);
and U9974 (N_9974,N_9650,N_9634);
nand U9975 (N_9975,N_9675,N_9756);
or U9976 (N_9976,N_9657,N_9601);
or U9977 (N_9977,N_9675,N_9697);
and U9978 (N_9978,N_9667,N_9647);
nand U9979 (N_9979,N_9668,N_9756);
nor U9980 (N_9980,N_9600,N_9614);
or U9981 (N_9981,N_9774,N_9622);
nand U9982 (N_9982,N_9653,N_9661);
nor U9983 (N_9983,N_9621,N_9705);
and U9984 (N_9984,N_9730,N_9627);
nor U9985 (N_9985,N_9732,N_9742);
nor U9986 (N_9986,N_9767,N_9748);
nand U9987 (N_9987,N_9650,N_9627);
and U9988 (N_9988,N_9603,N_9666);
nor U9989 (N_9989,N_9614,N_9736);
nor U9990 (N_9990,N_9702,N_9618);
or U9991 (N_9991,N_9696,N_9676);
or U9992 (N_9992,N_9648,N_9657);
or U9993 (N_9993,N_9683,N_9729);
nor U9994 (N_9994,N_9777,N_9735);
nor U9995 (N_9995,N_9707,N_9607);
or U9996 (N_9996,N_9676,N_9632);
nor U9997 (N_9997,N_9623,N_9615);
and U9998 (N_9998,N_9785,N_9798);
nor U9999 (N_9999,N_9652,N_9799);
nor UO_0 (O_0,N_9812,N_9922);
or UO_1 (O_1,N_9873,N_9968);
or UO_2 (O_2,N_9829,N_9889);
and UO_3 (O_3,N_9839,N_9808);
xnor UO_4 (O_4,N_9852,N_9927);
and UO_5 (O_5,N_9934,N_9910);
or UO_6 (O_6,N_9870,N_9987);
nand UO_7 (O_7,N_9996,N_9912);
and UO_8 (O_8,N_9826,N_9882);
nand UO_9 (O_9,N_9865,N_9957);
or UO_10 (O_10,N_9926,N_9817);
nor UO_11 (O_11,N_9810,N_9943);
and UO_12 (O_12,N_9891,N_9902);
or UO_13 (O_13,N_9911,N_9898);
xnor UO_14 (O_14,N_9960,N_9851);
nand UO_15 (O_15,N_9919,N_9853);
and UO_16 (O_16,N_9948,N_9903);
and UO_17 (O_17,N_9917,N_9894);
nand UO_18 (O_18,N_9918,N_9930);
nor UO_19 (O_19,N_9962,N_9884);
or UO_20 (O_20,N_9907,N_9887);
or UO_21 (O_21,N_9834,N_9809);
and UO_22 (O_22,N_9935,N_9897);
nand UO_23 (O_23,N_9967,N_9814);
xnor UO_24 (O_24,N_9835,N_9857);
or UO_25 (O_25,N_9893,N_9939);
and UO_26 (O_26,N_9854,N_9877);
and UO_27 (O_27,N_9971,N_9966);
nand UO_28 (O_28,N_9913,N_9980);
xor UO_29 (O_29,N_9856,N_9855);
nor UO_30 (O_30,N_9961,N_9828);
xor UO_31 (O_31,N_9822,N_9925);
or UO_32 (O_32,N_9909,N_9931);
nand UO_33 (O_33,N_9941,N_9946);
and UO_34 (O_34,N_9832,N_9995);
nand UO_35 (O_35,N_9921,N_9886);
or UO_36 (O_36,N_9973,N_9986);
and UO_37 (O_37,N_9849,N_9938);
xor UO_38 (O_38,N_9819,N_9970);
xnor UO_39 (O_39,N_9837,N_9950);
and UO_40 (O_40,N_9976,N_9982);
and UO_41 (O_41,N_9899,N_9876);
and UO_42 (O_42,N_9949,N_9900);
nand UO_43 (O_43,N_9878,N_9871);
nand UO_44 (O_44,N_9969,N_9896);
nor UO_45 (O_45,N_9860,N_9975);
and UO_46 (O_46,N_9963,N_9844);
or UO_47 (O_47,N_9827,N_9929);
and UO_48 (O_48,N_9908,N_9874);
nand UO_49 (O_49,N_9841,N_9823);
xnor UO_50 (O_50,N_9895,N_9953);
and UO_51 (O_51,N_9985,N_9915);
xor UO_52 (O_52,N_9940,N_9981);
and UO_53 (O_53,N_9848,N_9952);
and UO_54 (O_54,N_9991,N_9999);
xnor UO_55 (O_55,N_9859,N_9956);
nand UO_56 (O_56,N_9824,N_9862);
xor UO_57 (O_57,N_9888,N_9958);
and UO_58 (O_58,N_9892,N_9993);
and UO_59 (O_59,N_9923,N_9833);
and UO_60 (O_60,N_9869,N_9944);
or UO_61 (O_61,N_9932,N_9811);
nand UO_62 (O_62,N_9974,N_9924);
and UO_63 (O_63,N_9984,N_9845);
nor UO_64 (O_64,N_9866,N_9988);
nand UO_65 (O_65,N_9965,N_9977);
or UO_66 (O_66,N_9813,N_9864);
nand UO_67 (O_67,N_9990,N_9881);
and UO_68 (O_68,N_9997,N_9951);
and UO_69 (O_69,N_9803,N_9994);
xnor UO_70 (O_70,N_9979,N_9901);
nand UO_71 (O_71,N_9890,N_9840);
and UO_72 (O_72,N_9847,N_9955);
and UO_73 (O_73,N_9879,N_9861);
and UO_74 (O_74,N_9830,N_9964);
xnor UO_75 (O_75,N_9972,N_9906);
xor UO_76 (O_76,N_9933,N_9858);
and UO_77 (O_77,N_9836,N_9850);
or UO_78 (O_78,N_9916,N_9800);
or UO_79 (O_79,N_9942,N_9816);
nand UO_80 (O_80,N_9937,N_9992);
or UO_81 (O_81,N_9863,N_9945);
or UO_82 (O_82,N_9831,N_9914);
nor UO_83 (O_83,N_9820,N_9920);
nand UO_84 (O_84,N_9998,N_9875);
nand UO_85 (O_85,N_9880,N_9885);
nor UO_86 (O_86,N_9807,N_9821);
and UO_87 (O_87,N_9883,N_9806);
or UO_88 (O_88,N_9928,N_9818);
nand UO_89 (O_89,N_9815,N_9825);
and UO_90 (O_90,N_9867,N_9904);
nand UO_91 (O_91,N_9802,N_9801);
nand UO_92 (O_92,N_9989,N_9978);
nor UO_93 (O_93,N_9805,N_9983);
or UO_94 (O_94,N_9843,N_9872);
or UO_95 (O_95,N_9842,N_9905);
or UO_96 (O_96,N_9838,N_9959);
nor UO_97 (O_97,N_9936,N_9804);
nor UO_98 (O_98,N_9846,N_9954);
or UO_99 (O_99,N_9868,N_9947);
xnor UO_100 (O_100,N_9896,N_9867);
nand UO_101 (O_101,N_9988,N_9800);
xor UO_102 (O_102,N_9984,N_9927);
and UO_103 (O_103,N_9889,N_9887);
nor UO_104 (O_104,N_9862,N_9926);
or UO_105 (O_105,N_9906,N_9981);
or UO_106 (O_106,N_9821,N_9947);
and UO_107 (O_107,N_9908,N_9916);
nor UO_108 (O_108,N_9983,N_9885);
xor UO_109 (O_109,N_9932,N_9959);
or UO_110 (O_110,N_9954,N_9997);
or UO_111 (O_111,N_9921,N_9971);
nand UO_112 (O_112,N_9940,N_9846);
and UO_113 (O_113,N_9917,N_9803);
nand UO_114 (O_114,N_9981,N_9975);
and UO_115 (O_115,N_9809,N_9885);
nor UO_116 (O_116,N_9925,N_9976);
nand UO_117 (O_117,N_9912,N_9891);
and UO_118 (O_118,N_9992,N_9886);
or UO_119 (O_119,N_9960,N_9940);
nand UO_120 (O_120,N_9838,N_9875);
or UO_121 (O_121,N_9952,N_9913);
or UO_122 (O_122,N_9968,N_9854);
and UO_123 (O_123,N_9810,N_9981);
nand UO_124 (O_124,N_9890,N_9850);
nor UO_125 (O_125,N_9936,N_9809);
xor UO_126 (O_126,N_9980,N_9819);
or UO_127 (O_127,N_9979,N_9870);
nand UO_128 (O_128,N_9958,N_9968);
or UO_129 (O_129,N_9828,N_9910);
and UO_130 (O_130,N_9916,N_9825);
or UO_131 (O_131,N_9857,N_9920);
or UO_132 (O_132,N_9823,N_9908);
or UO_133 (O_133,N_9883,N_9926);
nand UO_134 (O_134,N_9844,N_9854);
or UO_135 (O_135,N_9869,N_9960);
or UO_136 (O_136,N_9952,N_9991);
or UO_137 (O_137,N_9914,N_9895);
nor UO_138 (O_138,N_9868,N_9869);
or UO_139 (O_139,N_9814,N_9961);
xnor UO_140 (O_140,N_9972,N_9934);
and UO_141 (O_141,N_9975,N_9820);
nor UO_142 (O_142,N_9812,N_9843);
nor UO_143 (O_143,N_9829,N_9878);
nor UO_144 (O_144,N_9811,N_9933);
xor UO_145 (O_145,N_9832,N_9847);
or UO_146 (O_146,N_9975,N_9986);
or UO_147 (O_147,N_9819,N_9850);
nor UO_148 (O_148,N_9956,N_9935);
and UO_149 (O_149,N_9966,N_9978);
nand UO_150 (O_150,N_9947,N_9946);
or UO_151 (O_151,N_9987,N_9815);
or UO_152 (O_152,N_9971,N_9897);
nand UO_153 (O_153,N_9848,N_9931);
nor UO_154 (O_154,N_9823,N_9837);
nand UO_155 (O_155,N_9960,N_9855);
nand UO_156 (O_156,N_9868,N_9907);
and UO_157 (O_157,N_9832,N_9991);
or UO_158 (O_158,N_9906,N_9975);
nor UO_159 (O_159,N_9850,N_9840);
nand UO_160 (O_160,N_9822,N_9999);
or UO_161 (O_161,N_9916,N_9811);
xnor UO_162 (O_162,N_9810,N_9842);
nor UO_163 (O_163,N_9957,N_9892);
nand UO_164 (O_164,N_9932,N_9990);
or UO_165 (O_165,N_9868,N_9873);
nor UO_166 (O_166,N_9938,N_9911);
xnor UO_167 (O_167,N_9878,N_9992);
nor UO_168 (O_168,N_9927,N_9898);
or UO_169 (O_169,N_9980,N_9941);
nand UO_170 (O_170,N_9977,N_9824);
or UO_171 (O_171,N_9963,N_9878);
nor UO_172 (O_172,N_9909,N_9981);
and UO_173 (O_173,N_9855,N_9904);
nand UO_174 (O_174,N_9806,N_9881);
nand UO_175 (O_175,N_9974,N_9955);
nor UO_176 (O_176,N_9937,N_9978);
nor UO_177 (O_177,N_9993,N_9938);
nand UO_178 (O_178,N_9872,N_9842);
nor UO_179 (O_179,N_9815,N_9947);
xnor UO_180 (O_180,N_9919,N_9868);
and UO_181 (O_181,N_9871,N_9849);
nor UO_182 (O_182,N_9996,N_9872);
and UO_183 (O_183,N_9841,N_9890);
and UO_184 (O_184,N_9911,N_9994);
and UO_185 (O_185,N_9874,N_9858);
nor UO_186 (O_186,N_9959,N_9937);
nand UO_187 (O_187,N_9836,N_9861);
and UO_188 (O_188,N_9836,N_9893);
xor UO_189 (O_189,N_9992,N_9973);
nor UO_190 (O_190,N_9882,N_9966);
and UO_191 (O_191,N_9949,N_9954);
xor UO_192 (O_192,N_9978,N_9963);
and UO_193 (O_193,N_9923,N_9997);
or UO_194 (O_194,N_9970,N_9893);
or UO_195 (O_195,N_9855,N_9892);
or UO_196 (O_196,N_9811,N_9891);
or UO_197 (O_197,N_9914,N_9986);
nand UO_198 (O_198,N_9882,N_9912);
or UO_199 (O_199,N_9824,N_9910);
or UO_200 (O_200,N_9934,N_9926);
nor UO_201 (O_201,N_9848,N_9979);
or UO_202 (O_202,N_9939,N_9977);
or UO_203 (O_203,N_9995,N_9930);
nand UO_204 (O_204,N_9832,N_9861);
nor UO_205 (O_205,N_9926,N_9815);
or UO_206 (O_206,N_9991,N_9903);
nor UO_207 (O_207,N_9916,N_9827);
nand UO_208 (O_208,N_9948,N_9839);
or UO_209 (O_209,N_9819,N_9841);
nand UO_210 (O_210,N_9972,N_9835);
and UO_211 (O_211,N_9867,N_9946);
nand UO_212 (O_212,N_9872,N_9965);
and UO_213 (O_213,N_9858,N_9862);
and UO_214 (O_214,N_9906,N_9947);
xnor UO_215 (O_215,N_9802,N_9835);
and UO_216 (O_216,N_9888,N_9869);
and UO_217 (O_217,N_9924,N_9869);
nand UO_218 (O_218,N_9983,N_9882);
and UO_219 (O_219,N_9958,N_9896);
nor UO_220 (O_220,N_9837,N_9996);
or UO_221 (O_221,N_9989,N_9854);
nor UO_222 (O_222,N_9830,N_9932);
nor UO_223 (O_223,N_9886,N_9922);
or UO_224 (O_224,N_9842,N_9803);
nor UO_225 (O_225,N_9861,N_9969);
nand UO_226 (O_226,N_9922,N_9996);
and UO_227 (O_227,N_9982,N_9898);
xor UO_228 (O_228,N_9870,N_9994);
nor UO_229 (O_229,N_9863,N_9852);
nor UO_230 (O_230,N_9803,N_9992);
nand UO_231 (O_231,N_9982,N_9826);
and UO_232 (O_232,N_9828,N_9857);
and UO_233 (O_233,N_9887,N_9995);
nor UO_234 (O_234,N_9940,N_9970);
or UO_235 (O_235,N_9959,N_9835);
nand UO_236 (O_236,N_9861,N_9945);
nand UO_237 (O_237,N_9882,N_9907);
nor UO_238 (O_238,N_9950,N_9964);
or UO_239 (O_239,N_9858,N_9979);
nand UO_240 (O_240,N_9821,N_9802);
nor UO_241 (O_241,N_9821,N_9966);
or UO_242 (O_242,N_9863,N_9959);
or UO_243 (O_243,N_9902,N_9865);
xnor UO_244 (O_244,N_9940,N_9973);
or UO_245 (O_245,N_9911,N_9941);
nand UO_246 (O_246,N_9932,N_9861);
nand UO_247 (O_247,N_9909,N_9938);
nor UO_248 (O_248,N_9835,N_9821);
xnor UO_249 (O_249,N_9826,N_9991);
nand UO_250 (O_250,N_9970,N_9832);
nor UO_251 (O_251,N_9882,N_9913);
xnor UO_252 (O_252,N_9942,N_9838);
nand UO_253 (O_253,N_9934,N_9859);
xor UO_254 (O_254,N_9905,N_9945);
or UO_255 (O_255,N_9827,N_9931);
nor UO_256 (O_256,N_9911,N_9880);
nor UO_257 (O_257,N_9934,N_9873);
nand UO_258 (O_258,N_9879,N_9874);
or UO_259 (O_259,N_9826,N_9971);
or UO_260 (O_260,N_9894,N_9984);
nand UO_261 (O_261,N_9960,N_9854);
nor UO_262 (O_262,N_9977,N_9851);
or UO_263 (O_263,N_9853,N_9997);
nor UO_264 (O_264,N_9916,N_9968);
xnor UO_265 (O_265,N_9830,N_9840);
nand UO_266 (O_266,N_9876,N_9846);
nand UO_267 (O_267,N_9995,N_9843);
nand UO_268 (O_268,N_9918,N_9837);
or UO_269 (O_269,N_9984,N_9855);
nand UO_270 (O_270,N_9968,N_9875);
and UO_271 (O_271,N_9991,N_9956);
and UO_272 (O_272,N_9818,N_9945);
or UO_273 (O_273,N_9991,N_9852);
nor UO_274 (O_274,N_9904,N_9836);
nor UO_275 (O_275,N_9829,N_9912);
and UO_276 (O_276,N_9848,N_9853);
and UO_277 (O_277,N_9877,N_9985);
nor UO_278 (O_278,N_9821,N_9994);
and UO_279 (O_279,N_9996,N_9967);
or UO_280 (O_280,N_9976,N_9800);
nand UO_281 (O_281,N_9987,N_9869);
nand UO_282 (O_282,N_9995,N_9943);
nand UO_283 (O_283,N_9839,N_9997);
and UO_284 (O_284,N_9966,N_9917);
and UO_285 (O_285,N_9988,N_9994);
xnor UO_286 (O_286,N_9997,N_9914);
nand UO_287 (O_287,N_9832,N_9806);
and UO_288 (O_288,N_9854,N_9905);
nand UO_289 (O_289,N_9943,N_9920);
or UO_290 (O_290,N_9913,N_9870);
nor UO_291 (O_291,N_9958,N_9813);
or UO_292 (O_292,N_9800,N_9939);
nor UO_293 (O_293,N_9982,N_9970);
and UO_294 (O_294,N_9935,N_9835);
nand UO_295 (O_295,N_9846,N_9982);
nand UO_296 (O_296,N_9996,N_9905);
or UO_297 (O_297,N_9914,N_9951);
and UO_298 (O_298,N_9902,N_9860);
nand UO_299 (O_299,N_9937,N_9989);
nand UO_300 (O_300,N_9996,N_9986);
nor UO_301 (O_301,N_9867,N_9954);
and UO_302 (O_302,N_9847,N_9808);
nor UO_303 (O_303,N_9996,N_9881);
xnor UO_304 (O_304,N_9819,N_9942);
nor UO_305 (O_305,N_9882,N_9937);
nand UO_306 (O_306,N_9949,N_9892);
nand UO_307 (O_307,N_9860,N_9965);
nand UO_308 (O_308,N_9918,N_9968);
nand UO_309 (O_309,N_9827,N_9912);
nand UO_310 (O_310,N_9953,N_9963);
nand UO_311 (O_311,N_9842,N_9823);
or UO_312 (O_312,N_9949,N_9849);
or UO_313 (O_313,N_9888,N_9993);
nand UO_314 (O_314,N_9832,N_9945);
nand UO_315 (O_315,N_9995,N_9853);
nand UO_316 (O_316,N_9817,N_9868);
or UO_317 (O_317,N_9837,N_9844);
nor UO_318 (O_318,N_9827,N_9881);
or UO_319 (O_319,N_9825,N_9888);
or UO_320 (O_320,N_9978,N_9988);
or UO_321 (O_321,N_9847,N_9944);
and UO_322 (O_322,N_9964,N_9954);
and UO_323 (O_323,N_9972,N_9942);
nor UO_324 (O_324,N_9801,N_9853);
or UO_325 (O_325,N_9962,N_9814);
or UO_326 (O_326,N_9834,N_9848);
nor UO_327 (O_327,N_9928,N_9845);
or UO_328 (O_328,N_9933,N_9990);
and UO_329 (O_329,N_9927,N_9933);
nand UO_330 (O_330,N_9983,N_9900);
nor UO_331 (O_331,N_9804,N_9818);
and UO_332 (O_332,N_9881,N_9850);
or UO_333 (O_333,N_9956,N_9800);
and UO_334 (O_334,N_9981,N_9862);
nor UO_335 (O_335,N_9924,N_9859);
nor UO_336 (O_336,N_9808,N_9866);
and UO_337 (O_337,N_9849,N_9922);
and UO_338 (O_338,N_9995,N_9813);
or UO_339 (O_339,N_9816,N_9992);
or UO_340 (O_340,N_9957,N_9855);
and UO_341 (O_341,N_9820,N_9836);
xnor UO_342 (O_342,N_9822,N_9869);
or UO_343 (O_343,N_9845,N_9966);
nand UO_344 (O_344,N_9902,N_9959);
nor UO_345 (O_345,N_9838,N_9876);
nor UO_346 (O_346,N_9961,N_9886);
or UO_347 (O_347,N_9967,N_9822);
xnor UO_348 (O_348,N_9954,N_9955);
nor UO_349 (O_349,N_9900,N_9991);
nor UO_350 (O_350,N_9847,N_9905);
or UO_351 (O_351,N_9822,N_9922);
nand UO_352 (O_352,N_9924,N_9995);
xnor UO_353 (O_353,N_9948,N_9957);
and UO_354 (O_354,N_9898,N_9875);
nor UO_355 (O_355,N_9954,N_9971);
and UO_356 (O_356,N_9879,N_9870);
nor UO_357 (O_357,N_9989,N_9964);
and UO_358 (O_358,N_9962,N_9873);
nor UO_359 (O_359,N_9829,N_9916);
nand UO_360 (O_360,N_9839,N_9943);
or UO_361 (O_361,N_9920,N_9813);
nor UO_362 (O_362,N_9967,N_9827);
nand UO_363 (O_363,N_9809,N_9858);
nand UO_364 (O_364,N_9872,N_9947);
nor UO_365 (O_365,N_9875,N_9848);
or UO_366 (O_366,N_9867,N_9840);
nand UO_367 (O_367,N_9996,N_9983);
and UO_368 (O_368,N_9974,N_9885);
and UO_369 (O_369,N_9826,N_9842);
nand UO_370 (O_370,N_9848,N_9928);
nand UO_371 (O_371,N_9913,N_9874);
nor UO_372 (O_372,N_9836,N_9854);
and UO_373 (O_373,N_9918,N_9982);
nor UO_374 (O_374,N_9994,N_9884);
or UO_375 (O_375,N_9826,N_9817);
nand UO_376 (O_376,N_9929,N_9999);
nand UO_377 (O_377,N_9841,N_9936);
and UO_378 (O_378,N_9819,N_9851);
and UO_379 (O_379,N_9885,N_9984);
or UO_380 (O_380,N_9870,N_9924);
or UO_381 (O_381,N_9918,N_9945);
and UO_382 (O_382,N_9803,N_9860);
nor UO_383 (O_383,N_9984,N_9870);
and UO_384 (O_384,N_9984,N_9940);
or UO_385 (O_385,N_9986,N_9807);
nand UO_386 (O_386,N_9967,N_9823);
or UO_387 (O_387,N_9880,N_9977);
and UO_388 (O_388,N_9891,N_9843);
or UO_389 (O_389,N_9977,N_9894);
and UO_390 (O_390,N_9866,N_9998);
nand UO_391 (O_391,N_9845,N_9925);
or UO_392 (O_392,N_9898,N_9818);
nor UO_393 (O_393,N_9816,N_9953);
nor UO_394 (O_394,N_9950,N_9971);
nand UO_395 (O_395,N_9868,N_9950);
xnor UO_396 (O_396,N_9842,N_9865);
nor UO_397 (O_397,N_9866,N_9966);
nor UO_398 (O_398,N_9893,N_9851);
xnor UO_399 (O_399,N_9844,N_9804);
nor UO_400 (O_400,N_9997,N_9872);
and UO_401 (O_401,N_9946,N_9887);
nor UO_402 (O_402,N_9858,N_9989);
or UO_403 (O_403,N_9817,N_9974);
and UO_404 (O_404,N_9971,N_9882);
and UO_405 (O_405,N_9903,N_9860);
nand UO_406 (O_406,N_9882,N_9901);
nand UO_407 (O_407,N_9894,N_9871);
nor UO_408 (O_408,N_9862,N_9976);
xor UO_409 (O_409,N_9969,N_9935);
and UO_410 (O_410,N_9818,N_9849);
or UO_411 (O_411,N_9901,N_9827);
nand UO_412 (O_412,N_9811,N_9853);
xnor UO_413 (O_413,N_9894,N_9870);
and UO_414 (O_414,N_9914,N_9924);
nor UO_415 (O_415,N_9908,N_9994);
nand UO_416 (O_416,N_9936,N_9874);
xor UO_417 (O_417,N_9858,N_9849);
or UO_418 (O_418,N_9865,N_9821);
or UO_419 (O_419,N_9961,N_9933);
xor UO_420 (O_420,N_9890,N_9976);
or UO_421 (O_421,N_9904,N_9925);
or UO_422 (O_422,N_9918,N_9840);
nand UO_423 (O_423,N_9977,N_9909);
and UO_424 (O_424,N_9881,N_9927);
or UO_425 (O_425,N_9973,N_9930);
xnor UO_426 (O_426,N_9832,N_9899);
or UO_427 (O_427,N_9807,N_9877);
and UO_428 (O_428,N_9851,N_9815);
xor UO_429 (O_429,N_9989,N_9800);
xnor UO_430 (O_430,N_9983,N_9852);
nand UO_431 (O_431,N_9890,N_9896);
and UO_432 (O_432,N_9886,N_9998);
nor UO_433 (O_433,N_9964,N_9962);
or UO_434 (O_434,N_9883,N_9853);
nand UO_435 (O_435,N_9861,N_9997);
and UO_436 (O_436,N_9937,N_9848);
or UO_437 (O_437,N_9817,N_9911);
or UO_438 (O_438,N_9985,N_9816);
and UO_439 (O_439,N_9830,N_9949);
nor UO_440 (O_440,N_9925,N_9874);
nand UO_441 (O_441,N_9975,N_9939);
nand UO_442 (O_442,N_9865,N_9891);
or UO_443 (O_443,N_9940,N_9911);
and UO_444 (O_444,N_9861,N_9831);
nor UO_445 (O_445,N_9992,N_9954);
nand UO_446 (O_446,N_9905,N_9874);
nor UO_447 (O_447,N_9855,N_9911);
nor UO_448 (O_448,N_9866,N_9980);
or UO_449 (O_449,N_9961,N_9875);
nor UO_450 (O_450,N_9863,N_9949);
and UO_451 (O_451,N_9837,N_9847);
nand UO_452 (O_452,N_9995,N_9925);
nor UO_453 (O_453,N_9837,N_9941);
nor UO_454 (O_454,N_9918,N_9912);
and UO_455 (O_455,N_9871,N_9898);
xnor UO_456 (O_456,N_9834,N_9907);
nor UO_457 (O_457,N_9811,N_9832);
nor UO_458 (O_458,N_9901,N_9852);
or UO_459 (O_459,N_9895,N_9863);
or UO_460 (O_460,N_9936,N_9885);
and UO_461 (O_461,N_9878,N_9815);
nor UO_462 (O_462,N_9928,N_9802);
and UO_463 (O_463,N_9957,N_9859);
nand UO_464 (O_464,N_9854,N_9907);
and UO_465 (O_465,N_9953,N_9822);
nor UO_466 (O_466,N_9886,N_9933);
or UO_467 (O_467,N_9854,N_9967);
nor UO_468 (O_468,N_9937,N_9836);
or UO_469 (O_469,N_9842,N_9890);
or UO_470 (O_470,N_9912,N_9974);
and UO_471 (O_471,N_9875,N_9834);
nand UO_472 (O_472,N_9816,N_9964);
and UO_473 (O_473,N_9988,N_9814);
nor UO_474 (O_474,N_9961,N_9824);
nor UO_475 (O_475,N_9960,N_9868);
and UO_476 (O_476,N_9982,N_9860);
or UO_477 (O_477,N_9947,N_9938);
and UO_478 (O_478,N_9959,N_9967);
xor UO_479 (O_479,N_9820,N_9821);
nor UO_480 (O_480,N_9948,N_9906);
nand UO_481 (O_481,N_9839,N_9823);
or UO_482 (O_482,N_9935,N_9928);
nor UO_483 (O_483,N_9893,N_9823);
nor UO_484 (O_484,N_9856,N_9926);
nor UO_485 (O_485,N_9890,N_9969);
and UO_486 (O_486,N_9924,N_9887);
or UO_487 (O_487,N_9815,N_9842);
nor UO_488 (O_488,N_9818,N_9900);
nor UO_489 (O_489,N_9961,N_9815);
and UO_490 (O_490,N_9925,N_9921);
nand UO_491 (O_491,N_9878,N_9854);
nand UO_492 (O_492,N_9880,N_9998);
and UO_493 (O_493,N_9926,N_9965);
and UO_494 (O_494,N_9978,N_9896);
or UO_495 (O_495,N_9922,N_9863);
or UO_496 (O_496,N_9837,N_9960);
or UO_497 (O_497,N_9892,N_9836);
nand UO_498 (O_498,N_9975,N_9902);
or UO_499 (O_499,N_9847,N_9844);
nand UO_500 (O_500,N_9883,N_9832);
and UO_501 (O_501,N_9879,N_9927);
and UO_502 (O_502,N_9916,N_9978);
nor UO_503 (O_503,N_9974,N_9954);
nand UO_504 (O_504,N_9850,N_9886);
nand UO_505 (O_505,N_9917,N_9898);
nand UO_506 (O_506,N_9829,N_9806);
or UO_507 (O_507,N_9809,N_9937);
or UO_508 (O_508,N_9977,N_9944);
nor UO_509 (O_509,N_9903,N_9953);
and UO_510 (O_510,N_9938,N_9810);
and UO_511 (O_511,N_9808,N_9976);
nand UO_512 (O_512,N_9866,N_9975);
and UO_513 (O_513,N_9847,N_9913);
nand UO_514 (O_514,N_9932,N_9890);
and UO_515 (O_515,N_9814,N_9861);
or UO_516 (O_516,N_9897,N_9915);
or UO_517 (O_517,N_9918,N_9940);
or UO_518 (O_518,N_9987,N_9831);
xor UO_519 (O_519,N_9983,N_9981);
nand UO_520 (O_520,N_9993,N_9857);
nand UO_521 (O_521,N_9867,N_9865);
or UO_522 (O_522,N_9831,N_9807);
or UO_523 (O_523,N_9853,N_9834);
nor UO_524 (O_524,N_9930,N_9949);
and UO_525 (O_525,N_9856,N_9873);
and UO_526 (O_526,N_9819,N_9880);
or UO_527 (O_527,N_9846,N_9943);
or UO_528 (O_528,N_9947,N_9831);
nor UO_529 (O_529,N_9882,N_9952);
xor UO_530 (O_530,N_9868,N_9976);
or UO_531 (O_531,N_9945,N_9868);
or UO_532 (O_532,N_9996,N_9902);
and UO_533 (O_533,N_9920,N_9814);
nand UO_534 (O_534,N_9817,N_9844);
and UO_535 (O_535,N_9968,N_9984);
nor UO_536 (O_536,N_9920,N_9907);
xnor UO_537 (O_537,N_9962,N_9917);
and UO_538 (O_538,N_9878,N_9998);
or UO_539 (O_539,N_9903,N_9817);
nand UO_540 (O_540,N_9839,N_9820);
and UO_541 (O_541,N_9978,N_9826);
and UO_542 (O_542,N_9847,N_9962);
nand UO_543 (O_543,N_9828,N_9992);
nor UO_544 (O_544,N_9829,N_9856);
nor UO_545 (O_545,N_9807,N_9834);
xor UO_546 (O_546,N_9962,N_9963);
nand UO_547 (O_547,N_9853,N_9993);
or UO_548 (O_548,N_9807,N_9810);
and UO_549 (O_549,N_9888,N_9901);
nor UO_550 (O_550,N_9896,N_9834);
nand UO_551 (O_551,N_9932,N_9817);
nor UO_552 (O_552,N_9929,N_9997);
xnor UO_553 (O_553,N_9892,N_9887);
nand UO_554 (O_554,N_9982,N_9917);
nor UO_555 (O_555,N_9832,N_9859);
nor UO_556 (O_556,N_9849,N_9814);
and UO_557 (O_557,N_9854,N_9923);
and UO_558 (O_558,N_9884,N_9925);
nor UO_559 (O_559,N_9944,N_9931);
or UO_560 (O_560,N_9804,N_9999);
and UO_561 (O_561,N_9914,N_9855);
and UO_562 (O_562,N_9938,N_9915);
or UO_563 (O_563,N_9999,N_9865);
nand UO_564 (O_564,N_9954,N_9879);
and UO_565 (O_565,N_9835,N_9946);
and UO_566 (O_566,N_9928,N_9875);
and UO_567 (O_567,N_9909,N_9855);
and UO_568 (O_568,N_9929,N_9903);
nor UO_569 (O_569,N_9802,N_9829);
nor UO_570 (O_570,N_9980,N_9915);
or UO_571 (O_571,N_9824,N_9938);
and UO_572 (O_572,N_9825,N_9968);
xnor UO_573 (O_573,N_9975,N_9995);
or UO_574 (O_574,N_9921,N_9894);
or UO_575 (O_575,N_9887,N_9830);
nor UO_576 (O_576,N_9925,N_9819);
and UO_577 (O_577,N_9889,N_9872);
or UO_578 (O_578,N_9912,N_9973);
nor UO_579 (O_579,N_9880,N_9901);
or UO_580 (O_580,N_9866,N_9836);
or UO_581 (O_581,N_9943,N_9958);
and UO_582 (O_582,N_9943,N_9951);
nand UO_583 (O_583,N_9931,N_9870);
nor UO_584 (O_584,N_9829,N_9847);
nand UO_585 (O_585,N_9998,N_9847);
nand UO_586 (O_586,N_9948,N_9833);
nor UO_587 (O_587,N_9853,N_9935);
and UO_588 (O_588,N_9860,N_9923);
xnor UO_589 (O_589,N_9889,N_9992);
nor UO_590 (O_590,N_9859,N_9951);
nand UO_591 (O_591,N_9864,N_9870);
nand UO_592 (O_592,N_9833,N_9930);
nor UO_593 (O_593,N_9824,N_9801);
nand UO_594 (O_594,N_9858,N_9864);
or UO_595 (O_595,N_9877,N_9953);
nor UO_596 (O_596,N_9911,N_9836);
or UO_597 (O_597,N_9850,N_9949);
nor UO_598 (O_598,N_9833,N_9813);
nand UO_599 (O_599,N_9813,N_9840);
nor UO_600 (O_600,N_9994,N_9868);
or UO_601 (O_601,N_9955,N_9959);
and UO_602 (O_602,N_9886,N_9839);
nand UO_603 (O_603,N_9999,N_9885);
or UO_604 (O_604,N_9911,N_9944);
xnor UO_605 (O_605,N_9929,N_9821);
or UO_606 (O_606,N_9815,N_9936);
nor UO_607 (O_607,N_9826,N_9968);
nand UO_608 (O_608,N_9891,N_9859);
xnor UO_609 (O_609,N_9806,N_9981);
nand UO_610 (O_610,N_9949,N_9847);
nor UO_611 (O_611,N_9971,N_9810);
nand UO_612 (O_612,N_9958,N_9863);
or UO_613 (O_613,N_9955,N_9969);
or UO_614 (O_614,N_9992,N_9991);
nand UO_615 (O_615,N_9892,N_9943);
or UO_616 (O_616,N_9990,N_9818);
or UO_617 (O_617,N_9898,N_9856);
and UO_618 (O_618,N_9950,N_9925);
xor UO_619 (O_619,N_9995,N_9983);
nor UO_620 (O_620,N_9829,N_9932);
or UO_621 (O_621,N_9998,N_9863);
nand UO_622 (O_622,N_9813,N_9861);
or UO_623 (O_623,N_9888,N_9819);
or UO_624 (O_624,N_9807,N_9912);
nor UO_625 (O_625,N_9988,N_9975);
nor UO_626 (O_626,N_9859,N_9840);
or UO_627 (O_627,N_9850,N_9897);
xnor UO_628 (O_628,N_9842,N_9928);
nand UO_629 (O_629,N_9914,N_9835);
nor UO_630 (O_630,N_9993,N_9828);
nand UO_631 (O_631,N_9941,N_9904);
or UO_632 (O_632,N_9991,N_9982);
or UO_633 (O_633,N_9982,N_9861);
xnor UO_634 (O_634,N_9887,N_9934);
nand UO_635 (O_635,N_9915,N_9979);
nand UO_636 (O_636,N_9847,N_9901);
and UO_637 (O_637,N_9853,N_9829);
or UO_638 (O_638,N_9912,N_9888);
and UO_639 (O_639,N_9919,N_9943);
nand UO_640 (O_640,N_9947,N_9844);
and UO_641 (O_641,N_9836,N_9949);
and UO_642 (O_642,N_9928,N_9830);
xnor UO_643 (O_643,N_9923,N_9992);
nor UO_644 (O_644,N_9918,N_9838);
nand UO_645 (O_645,N_9845,N_9895);
or UO_646 (O_646,N_9939,N_9867);
and UO_647 (O_647,N_9943,N_9842);
and UO_648 (O_648,N_9957,N_9873);
or UO_649 (O_649,N_9866,N_9859);
nor UO_650 (O_650,N_9939,N_9824);
nand UO_651 (O_651,N_9981,N_9844);
and UO_652 (O_652,N_9804,N_9813);
nand UO_653 (O_653,N_9818,N_9878);
or UO_654 (O_654,N_9861,N_9938);
nor UO_655 (O_655,N_9957,N_9856);
or UO_656 (O_656,N_9939,N_9927);
or UO_657 (O_657,N_9860,N_9846);
and UO_658 (O_658,N_9998,N_9977);
or UO_659 (O_659,N_9933,N_9829);
or UO_660 (O_660,N_9993,N_9943);
nand UO_661 (O_661,N_9807,N_9817);
xor UO_662 (O_662,N_9806,N_9867);
nand UO_663 (O_663,N_9840,N_9968);
and UO_664 (O_664,N_9966,N_9905);
xor UO_665 (O_665,N_9995,N_9940);
nor UO_666 (O_666,N_9953,N_9811);
nor UO_667 (O_667,N_9831,N_9997);
nor UO_668 (O_668,N_9934,N_9948);
nor UO_669 (O_669,N_9927,N_9924);
nor UO_670 (O_670,N_9865,N_9974);
nand UO_671 (O_671,N_9967,N_9904);
nand UO_672 (O_672,N_9992,N_9860);
or UO_673 (O_673,N_9995,N_9984);
xnor UO_674 (O_674,N_9875,N_9809);
nand UO_675 (O_675,N_9885,N_9945);
and UO_676 (O_676,N_9859,N_9998);
nand UO_677 (O_677,N_9890,N_9860);
or UO_678 (O_678,N_9896,N_9998);
and UO_679 (O_679,N_9838,N_9960);
nand UO_680 (O_680,N_9845,N_9976);
or UO_681 (O_681,N_9868,N_9918);
nor UO_682 (O_682,N_9966,N_9869);
and UO_683 (O_683,N_9970,N_9978);
nand UO_684 (O_684,N_9936,N_9888);
and UO_685 (O_685,N_9816,N_9966);
nand UO_686 (O_686,N_9880,N_9960);
nor UO_687 (O_687,N_9818,N_9867);
nor UO_688 (O_688,N_9854,N_9930);
nor UO_689 (O_689,N_9942,N_9960);
nor UO_690 (O_690,N_9841,N_9921);
xnor UO_691 (O_691,N_9840,N_9901);
nor UO_692 (O_692,N_9922,N_9834);
and UO_693 (O_693,N_9808,N_9891);
and UO_694 (O_694,N_9807,N_9954);
nand UO_695 (O_695,N_9866,N_9882);
xnor UO_696 (O_696,N_9826,N_9923);
or UO_697 (O_697,N_9936,N_9947);
nor UO_698 (O_698,N_9979,N_9996);
xnor UO_699 (O_699,N_9932,N_9894);
nor UO_700 (O_700,N_9886,N_9944);
and UO_701 (O_701,N_9897,N_9954);
and UO_702 (O_702,N_9966,N_9999);
or UO_703 (O_703,N_9937,N_9879);
nor UO_704 (O_704,N_9894,N_9918);
or UO_705 (O_705,N_9839,N_9884);
nor UO_706 (O_706,N_9856,N_9811);
and UO_707 (O_707,N_9919,N_9852);
or UO_708 (O_708,N_9802,N_9937);
nor UO_709 (O_709,N_9899,N_9978);
and UO_710 (O_710,N_9879,N_9903);
nor UO_711 (O_711,N_9975,N_9803);
xnor UO_712 (O_712,N_9822,N_9841);
nand UO_713 (O_713,N_9867,N_9967);
and UO_714 (O_714,N_9878,N_9866);
or UO_715 (O_715,N_9898,N_9907);
or UO_716 (O_716,N_9908,N_9946);
nand UO_717 (O_717,N_9981,N_9821);
nand UO_718 (O_718,N_9889,N_9812);
nor UO_719 (O_719,N_9897,N_9942);
nand UO_720 (O_720,N_9935,N_9900);
nand UO_721 (O_721,N_9907,N_9852);
nand UO_722 (O_722,N_9954,N_9874);
nor UO_723 (O_723,N_9950,N_9877);
nor UO_724 (O_724,N_9932,N_9804);
xnor UO_725 (O_725,N_9932,N_9855);
or UO_726 (O_726,N_9940,N_9915);
and UO_727 (O_727,N_9946,N_9982);
or UO_728 (O_728,N_9959,N_9823);
nand UO_729 (O_729,N_9971,N_9855);
nand UO_730 (O_730,N_9876,N_9930);
nor UO_731 (O_731,N_9923,N_9831);
and UO_732 (O_732,N_9993,N_9991);
or UO_733 (O_733,N_9801,N_9997);
or UO_734 (O_734,N_9907,N_9869);
nor UO_735 (O_735,N_9820,N_9898);
or UO_736 (O_736,N_9979,N_9837);
and UO_737 (O_737,N_9825,N_9976);
or UO_738 (O_738,N_9977,N_9821);
nor UO_739 (O_739,N_9905,N_9938);
or UO_740 (O_740,N_9903,N_9913);
nor UO_741 (O_741,N_9845,N_9906);
xnor UO_742 (O_742,N_9892,N_9921);
or UO_743 (O_743,N_9962,N_9856);
and UO_744 (O_744,N_9827,N_9961);
nor UO_745 (O_745,N_9815,N_9844);
and UO_746 (O_746,N_9857,N_9816);
xnor UO_747 (O_747,N_9966,N_9841);
nand UO_748 (O_748,N_9805,N_9965);
or UO_749 (O_749,N_9912,N_9892);
or UO_750 (O_750,N_9979,N_9818);
nand UO_751 (O_751,N_9896,N_9891);
and UO_752 (O_752,N_9946,N_9911);
nor UO_753 (O_753,N_9907,N_9896);
or UO_754 (O_754,N_9918,N_9928);
and UO_755 (O_755,N_9892,N_9978);
nand UO_756 (O_756,N_9982,N_9887);
or UO_757 (O_757,N_9997,N_9826);
nand UO_758 (O_758,N_9959,N_9883);
nand UO_759 (O_759,N_9935,N_9948);
and UO_760 (O_760,N_9977,N_9904);
and UO_761 (O_761,N_9968,N_9829);
and UO_762 (O_762,N_9956,N_9964);
nand UO_763 (O_763,N_9817,N_9927);
xor UO_764 (O_764,N_9873,N_9877);
xor UO_765 (O_765,N_9922,N_9902);
and UO_766 (O_766,N_9945,N_9901);
nor UO_767 (O_767,N_9990,N_9866);
nor UO_768 (O_768,N_9949,N_9815);
nand UO_769 (O_769,N_9979,N_9973);
and UO_770 (O_770,N_9980,N_9970);
or UO_771 (O_771,N_9989,N_9948);
or UO_772 (O_772,N_9997,N_9917);
nand UO_773 (O_773,N_9870,N_9926);
and UO_774 (O_774,N_9947,N_9993);
nand UO_775 (O_775,N_9921,N_9913);
nor UO_776 (O_776,N_9851,N_9850);
and UO_777 (O_777,N_9844,N_9929);
and UO_778 (O_778,N_9896,N_9881);
or UO_779 (O_779,N_9918,N_9915);
nand UO_780 (O_780,N_9833,N_9890);
nor UO_781 (O_781,N_9976,N_9949);
xor UO_782 (O_782,N_9929,N_9993);
and UO_783 (O_783,N_9813,N_9870);
nor UO_784 (O_784,N_9909,N_9829);
and UO_785 (O_785,N_9930,N_9994);
nor UO_786 (O_786,N_9953,N_9827);
or UO_787 (O_787,N_9880,N_9873);
xnor UO_788 (O_788,N_9968,N_9888);
and UO_789 (O_789,N_9931,N_9960);
nand UO_790 (O_790,N_9834,N_9827);
or UO_791 (O_791,N_9997,N_9903);
nand UO_792 (O_792,N_9962,N_9838);
nand UO_793 (O_793,N_9882,N_9885);
and UO_794 (O_794,N_9888,N_9949);
nand UO_795 (O_795,N_9887,N_9917);
nand UO_796 (O_796,N_9811,N_9917);
nand UO_797 (O_797,N_9965,N_9909);
nor UO_798 (O_798,N_9918,N_9820);
and UO_799 (O_799,N_9869,N_9829);
or UO_800 (O_800,N_9901,N_9898);
nand UO_801 (O_801,N_9829,N_9976);
and UO_802 (O_802,N_9926,N_9852);
nand UO_803 (O_803,N_9907,N_9843);
xor UO_804 (O_804,N_9990,N_9940);
or UO_805 (O_805,N_9828,N_9839);
nor UO_806 (O_806,N_9926,N_9804);
nor UO_807 (O_807,N_9814,N_9942);
nor UO_808 (O_808,N_9960,N_9800);
nand UO_809 (O_809,N_9817,N_9876);
or UO_810 (O_810,N_9987,N_9985);
and UO_811 (O_811,N_9902,N_9855);
nor UO_812 (O_812,N_9929,N_9911);
nor UO_813 (O_813,N_9879,N_9972);
and UO_814 (O_814,N_9951,N_9925);
xor UO_815 (O_815,N_9884,N_9882);
or UO_816 (O_816,N_9904,N_9884);
or UO_817 (O_817,N_9963,N_9982);
or UO_818 (O_818,N_9967,N_9906);
xnor UO_819 (O_819,N_9913,N_9901);
nor UO_820 (O_820,N_9950,N_9805);
nor UO_821 (O_821,N_9813,N_9936);
nor UO_822 (O_822,N_9925,N_9978);
and UO_823 (O_823,N_9833,N_9994);
nor UO_824 (O_824,N_9998,N_9971);
nor UO_825 (O_825,N_9826,N_9962);
nand UO_826 (O_826,N_9807,N_9908);
or UO_827 (O_827,N_9861,N_9869);
xor UO_828 (O_828,N_9945,N_9864);
or UO_829 (O_829,N_9835,N_9824);
nor UO_830 (O_830,N_9905,N_9903);
xor UO_831 (O_831,N_9961,N_9860);
or UO_832 (O_832,N_9825,N_9810);
nand UO_833 (O_833,N_9910,N_9924);
xor UO_834 (O_834,N_9815,N_9916);
and UO_835 (O_835,N_9821,N_9809);
or UO_836 (O_836,N_9823,N_9849);
xor UO_837 (O_837,N_9881,N_9942);
or UO_838 (O_838,N_9925,N_9888);
or UO_839 (O_839,N_9913,N_9919);
or UO_840 (O_840,N_9850,N_9906);
and UO_841 (O_841,N_9802,N_9874);
nand UO_842 (O_842,N_9990,N_9844);
nand UO_843 (O_843,N_9983,N_9974);
nand UO_844 (O_844,N_9873,N_9824);
and UO_845 (O_845,N_9880,N_9968);
nor UO_846 (O_846,N_9839,N_9995);
nor UO_847 (O_847,N_9913,N_9801);
nand UO_848 (O_848,N_9937,N_9914);
or UO_849 (O_849,N_9919,N_9880);
and UO_850 (O_850,N_9818,N_9861);
xor UO_851 (O_851,N_9875,N_9976);
nor UO_852 (O_852,N_9873,N_9847);
nand UO_853 (O_853,N_9904,N_9937);
and UO_854 (O_854,N_9959,N_9854);
or UO_855 (O_855,N_9999,N_9809);
or UO_856 (O_856,N_9955,N_9929);
nor UO_857 (O_857,N_9854,N_9982);
or UO_858 (O_858,N_9801,N_9954);
nor UO_859 (O_859,N_9865,N_9855);
and UO_860 (O_860,N_9855,N_9868);
nand UO_861 (O_861,N_9834,N_9805);
nor UO_862 (O_862,N_9877,N_9912);
and UO_863 (O_863,N_9918,N_9863);
or UO_864 (O_864,N_9944,N_9936);
nand UO_865 (O_865,N_9999,N_9987);
nor UO_866 (O_866,N_9891,N_9987);
nor UO_867 (O_867,N_9922,N_9970);
or UO_868 (O_868,N_9836,N_9938);
nor UO_869 (O_869,N_9959,N_9919);
or UO_870 (O_870,N_9915,N_9914);
or UO_871 (O_871,N_9846,N_9820);
xor UO_872 (O_872,N_9979,N_9930);
and UO_873 (O_873,N_9928,N_9872);
nor UO_874 (O_874,N_9913,N_9959);
xnor UO_875 (O_875,N_9983,N_9919);
and UO_876 (O_876,N_9976,N_9970);
nand UO_877 (O_877,N_9800,N_9972);
and UO_878 (O_878,N_9811,N_9977);
nor UO_879 (O_879,N_9953,N_9931);
xnor UO_880 (O_880,N_9891,N_9853);
and UO_881 (O_881,N_9819,N_9859);
and UO_882 (O_882,N_9835,N_9828);
nand UO_883 (O_883,N_9877,N_9994);
nor UO_884 (O_884,N_9951,N_9844);
nor UO_885 (O_885,N_9919,N_9953);
nor UO_886 (O_886,N_9816,N_9859);
and UO_887 (O_887,N_9892,N_9944);
nand UO_888 (O_888,N_9992,N_9870);
nand UO_889 (O_889,N_9882,N_9978);
nand UO_890 (O_890,N_9839,N_9893);
or UO_891 (O_891,N_9976,N_9953);
nand UO_892 (O_892,N_9993,N_9935);
or UO_893 (O_893,N_9982,N_9912);
nor UO_894 (O_894,N_9876,N_9923);
xnor UO_895 (O_895,N_9974,N_9899);
nor UO_896 (O_896,N_9814,N_9813);
nor UO_897 (O_897,N_9999,N_9956);
or UO_898 (O_898,N_9956,N_9813);
or UO_899 (O_899,N_9857,N_9959);
nor UO_900 (O_900,N_9860,N_9883);
nand UO_901 (O_901,N_9888,N_9833);
or UO_902 (O_902,N_9995,N_9859);
nor UO_903 (O_903,N_9923,N_9889);
nor UO_904 (O_904,N_9881,N_9980);
or UO_905 (O_905,N_9923,N_9801);
or UO_906 (O_906,N_9996,N_9882);
nor UO_907 (O_907,N_9829,N_9961);
nor UO_908 (O_908,N_9838,N_9912);
nand UO_909 (O_909,N_9985,N_9993);
or UO_910 (O_910,N_9934,N_9816);
and UO_911 (O_911,N_9882,N_9934);
or UO_912 (O_912,N_9892,N_9951);
or UO_913 (O_913,N_9817,N_9962);
nand UO_914 (O_914,N_9855,N_9873);
nand UO_915 (O_915,N_9952,N_9893);
nor UO_916 (O_916,N_9892,N_9965);
nand UO_917 (O_917,N_9933,N_9917);
or UO_918 (O_918,N_9983,N_9827);
and UO_919 (O_919,N_9906,N_9882);
and UO_920 (O_920,N_9896,N_9862);
and UO_921 (O_921,N_9880,N_9844);
nand UO_922 (O_922,N_9806,N_9890);
nor UO_923 (O_923,N_9894,N_9998);
nor UO_924 (O_924,N_9887,N_9825);
or UO_925 (O_925,N_9978,N_9903);
nor UO_926 (O_926,N_9956,N_9897);
and UO_927 (O_927,N_9950,N_9878);
xnor UO_928 (O_928,N_9859,N_9960);
and UO_929 (O_929,N_9802,N_9960);
nand UO_930 (O_930,N_9828,N_9998);
and UO_931 (O_931,N_9814,N_9936);
and UO_932 (O_932,N_9954,N_9816);
nand UO_933 (O_933,N_9803,N_9879);
and UO_934 (O_934,N_9927,N_9994);
nor UO_935 (O_935,N_9848,N_9961);
or UO_936 (O_936,N_9928,N_9940);
xnor UO_937 (O_937,N_9834,N_9874);
xnor UO_938 (O_938,N_9821,N_9852);
nor UO_939 (O_939,N_9999,N_9815);
and UO_940 (O_940,N_9999,N_9801);
or UO_941 (O_941,N_9820,N_9961);
or UO_942 (O_942,N_9800,N_9892);
nand UO_943 (O_943,N_9880,N_9827);
and UO_944 (O_944,N_9998,N_9929);
and UO_945 (O_945,N_9857,N_9960);
or UO_946 (O_946,N_9806,N_9986);
nand UO_947 (O_947,N_9969,N_9984);
nand UO_948 (O_948,N_9985,N_9846);
and UO_949 (O_949,N_9844,N_9952);
and UO_950 (O_950,N_9901,N_9917);
and UO_951 (O_951,N_9967,N_9980);
or UO_952 (O_952,N_9801,N_9993);
nand UO_953 (O_953,N_9887,N_9999);
nand UO_954 (O_954,N_9876,N_9858);
nand UO_955 (O_955,N_9981,N_9953);
nor UO_956 (O_956,N_9824,N_9816);
nand UO_957 (O_957,N_9965,N_9981);
nor UO_958 (O_958,N_9906,N_9939);
nand UO_959 (O_959,N_9958,N_9970);
nand UO_960 (O_960,N_9933,N_9867);
nand UO_961 (O_961,N_9916,N_9813);
and UO_962 (O_962,N_9955,N_9813);
nand UO_963 (O_963,N_9968,N_9998);
nand UO_964 (O_964,N_9961,N_9972);
nand UO_965 (O_965,N_9804,N_9939);
nand UO_966 (O_966,N_9953,N_9961);
and UO_967 (O_967,N_9843,N_9838);
and UO_968 (O_968,N_9873,N_9944);
nand UO_969 (O_969,N_9951,N_9893);
xor UO_970 (O_970,N_9983,N_9815);
and UO_971 (O_971,N_9859,N_9839);
or UO_972 (O_972,N_9847,N_9856);
nor UO_973 (O_973,N_9916,N_9932);
and UO_974 (O_974,N_9816,N_9881);
xor UO_975 (O_975,N_9884,N_9892);
xor UO_976 (O_976,N_9827,N_9945);
xnor UO_977 (O_977,N_9887,N_9850);
and UO_978 (O_978,N_9805,N_9954);
xor UO_979 (O_979,N_9849,N_9848);
nand UO_980 (O_980,N_9989,N_9851);
nand UO_981 (O_981,N_9820,N_9803);
nor UO_982 (O_982,N_9816,N_9988);
nand UO_983 (O_983,N_9834,N_9935);
or UO_984 (O_984,N_9849,N_9988);
nor UO_985 (O_985,N_9811,N_9879);
nor UO_986 (O_986,N_9966,N_9873);
nand UO_987 (O_987,N_9988,N_9870);
nor UO_988 (O_988,N_9825,N_9841);
and UO_989 (O_989,N_9824,N_9865);
and UO_990 (O_990,N_9914,N_9994);
xnor UO_991 (O_991,N_9992,N_9817);
xnor UO_992 (O_992,N_9887,N_9904);
and UO_993 (O_993,N_9970,N_9897);
and UO_994 (O_994,N_9974,N_9832);
and UO_995 (O_995,N_9974,N_9868);
nor UO_996 (O_996,N_9949,N_9935);
nor UO_997 (O_997,N_9931,N_9829);
or UO_998 (O_998,N_9812,N_9903);
and UO_999 (O_999,N_9997,N_9806);
and UO_1000 (O_1000,N_9898,N_9959);
nor UO_1001 (O_1001,N_9885,N_9881);
nor UO_1002 (O_1002,N_9899,N_9993);
nor UO_1003 (O_1003,N_9853,N_9892);
and UO_1004 (O_1004,N_9846,N_9840);
and UO_1005 (O_1005,N_9928,N_9924);
xor UO_1006 (O_1006,N_9877,N_9812);
nor UO_1007 (O_1007,N_9977,N_9937);
nand UO_1008 (O_1008,N_9981,N_9864);
and UO_1009 (O_1009,N_9985,N_9828);
nand UO_1010 (O_1010,N_9902,N_9871);
nor UO_1011 (O_1011,N_9897,N_9939);
or UO_1012 (O_1012,N_9928,N_9899);
xnor UO_1013 (O_1013,N_9825,N_9907);
nor UO_1014 (O_1014,N_9810,N_9811);
nand UO_1015 (O_1015,N_9928,N_9846);
or UO_1016 (O_1016,N_9875,N_9916);
or UO_1017 (O_1017,N_9964,N_9975);
or UO_1018 (O_1018,N_9995,N_9936);
nand UO_1019 (O_1019,N_9999,N_9820);
nand UO_1020 (O_1020,N_9817,N_9964);
nor UO_1021 (O_1021,N_9857,N_9921);
and UO_1022 (O_1022,N_9888,N_9947);
and UO_1023 (O_1023,N_9911,N_9816);
and UO_1024 (O_1024,N_9831,N_9863);
xnor UO_1025 (O_1025,N_9978,N_9808);
nor UO_1026 (O_1026,N_9926,N_9887);
nand UO_1027 (O_1027,N_9915,N_9854);
nor UO_1028 (O_1028,N_9971,N_9928);
nor UO_1029 (O_1029,N_9918,N_9919);
and UO_1030 (O_1030,N_9898,N_9916);
nand UO_1031 (O_1031,N_9892,N_9804);
or UO_1032 (O_1032,N_9960,N_9973);
and UO_1033 (O_1033,N_9835,N_9984);
nand UO_1034 (O_1034,N_9906,N_9953);
nand UO_1035 (O_1035,N_9872,N_9841);
nor UO_1036 (O_1036,N_9984,N_9979);
nor UO_1037 (O_1037,N_9924,N_9929);
nor UO_1038 (O_1038,N_9802,N_9966);
and UO_1039 (O_1039,N_9815,N_9974);
nor UO_1040 (O_1040,N_9952,N_9809);
and UO_1041 (O_1041,N_9842,N_9862);
or UO_1042 (O_1042,N_9924,N_9840);
nand UO_1043 (O_1043,N_9960,N_9824);
nor UO_1044 (O_1044,N_9945,N_9964);
nor UO_1045 (O_1045,N_9861,N_9864);
nor UO_1046 (O_1046,N_9951,N_9986);
nor UO_1047 (O_1047,N_9875,N_9974);
nand UO_1048 (O_1048,N_9890,N_9882);
nand UO_1049 (O_1049,N_9899,N_9844);
nand UO_1050 (O_1050,N_9803,N_9862);
nor UO_1051 (O_1051,N_9828,N_9988);
or UO_1052 (O_1052,N_9926,N_9812);
and UO_1053 (O_1053,N_9967,N_9857);
or UO_1054 (O_1054,N_9966,N_9959);
or UO_1055 (O_1055,N_9953,N_9883);
and UO_1056 (O_1056,N_9971,N_9967);
nand UO_1057 (O_1057,N_9859,N_9968);
nand UO_1058 (O_1058,N_9843,N_9841);
and UO_1059 (O_1059,N_9969,N_9889);
and UO_1060 (O_1060,N_9856,N_9967);
and UO_1061 (O_1061,N_9994,N_9918);
and UO_1062 (O_1062,N_9992,N_9969);
and UO_1063 (O_1063,N_9982,N_9848);
and UO_1064 (O_1064,N_9908,N_9934);
and UO_1065 (O_1065,N_9853,N_9946);
and UO_1066 (O_1066,N_9954,N_9812);
and UO_1067 (O_1067,N_9891,N_9988);
or UO_1068 (O_1068,N_9907,N_9965);
nand UO_1069 (O_1069,N_9875,N_9890);
nor UO_1070 (O_1070,N_9898,N_9994);
xor UO_1071 (O_1071,N_9955,N_9892);
or UO_1072 (O_1072,N_9983,N_9941);
or UO_1073 (O_1073,N_9959,N_9956);
nor UO_1074 (O_1074,N_9877,N_9938);
nand UO_1075 (O_1075,N_9919,N_9844);
or UO_1076 (O_1076,N_9838,N_9801);
or UO_1077 (O_1077,N_9983,N_9903);
nor UO_1078 (O_1078,N_9836,N_9833);
nand UO_1079 (O_1079,N_9850,N_9963);
and UO_1080 (O_1080,N_9893,N_9905);
xnor UO_1081 (O_1081,N_9966,N_9992);
or UO_1082 (O_1082,N_9924,N_9802);
and UO_1083 (O_1083,N_9860,N_9931);
or UO_1084 (O_1084,N_9922,N_9939);
or UO_1085 (O_1085,N_9854,N_9976);
and UO_1086 (O_1086,N_9999,N_9989);
xor UO_1087 (O_1087,N_9912,N_9966);
nand UO_1088 (O_1088,N_9816,N_9962);
nor UO_1089 (O_1089,N_9914,N_9868);
xnor UO_1090 (O_1090,N_9899,N_9802);
and UO_1091 (O_1091,N_9899,N_9890);
or UO_1092 (O_1092,N_9800,N_9822);
or UO_1093 (O_1093,N_9867,N_9917);
xnor UO_1094 (O_1094,N_9967,N_9993);
and UO_1095 (O_1095,N_9852,N_9825);
nor UO_1096 (O_1096,N_9890,N_9855);
nand UO_1097 (O_1097,N_9845,N_9988);
or UO_1098 (O_1098,N_9893,N_9903);
or UO_1099 (O_1099,N_9925,N_9841);
nand UO_1100 (O_1100,N_9828,N_9861);
or UO_1101 (O_1101,N_9965,N_9863);
nand UO_1102 (O_1102,N_9801,N_9888);
or UO_1103 (O_1103,N_9983,N_9969);
or UO_1104 (O_1104,N_9953,N_9950);
nor UO_1105 (O_1105,N_9928,N_9987);
or UO_1106 (O_1106,N_9948,N_9842);
or UO_1107 (O_1107,N_9979,N_9815);
nor UO_1108 (O_1108,N_9908,N_9800);
nand UO_1109 (O_1109,N_9827,N_9956);
xor UO_1110 (O_1110,N_9877,N_9933);
or UO_1111 (O_1111,N_9974,N_9959);
or UO_1112 (O_1112,N_9923,N_9810);
and UO_1113 (O_1113,N_9889,N_9988);
xor UO_1114 (O_1114,N_9849,N_9841);
or UO_1115 (O_1115,N_9930,N_9923);
nand UO_1116 (O_1116,N_9818,N_9833);
nand UO_1117 (O_1117,N_9892,N_9835);
or UO_1118 (O_1118,N_9953,N_9851);
nand UO_1119 (O_1119,N_9830,N_9958);
or UO_1120 (O_1120,N_9939,N_9811);
nor UO_1121 (O_1121,N_9845,N_9944);
nor UO_1122 (O_1122,N_9940,N_9883);
and UO_1123 (O_1123,N_9824,N_9857);
nor UO_1124 (O_1124,N_9894,N_9933);
or UO_1125 (O_1125,N_9903,N_9895);
and UO_1126 (O_1126,N_9994,N_9975);
nand UO_1127 (O_1127,N_9832,N_9809);
nor UO_1128 (O_1128,N_9934,N_9858);
nor UO_1129 (O_1129,N_9854,N_9879);
and UO_1130 (O_1130,N_9923,N_9857);
nor UO_1131 (O_1131,N_9954,N_9860);
or UO_1132 (O_1132,N_9859,N_9836);
or UO_1133 (O_1133,N_9952,N_9909);
and UO_1134 (O_1134,N_9969,N_9904);
nor UO_1135 (O_1135,N_9952,N_9919);
nor UO_1136 (O_1136,N_9917,N_9903);
nor UO_1137 (O_1137,N_9933,N_9975);
and UO_1138 (O_1138,N_9966,N_9988);
and UO_1139 (O_1139,N_9958,N_9966);
nand UO_1140 (O_1140,N_9997,N_9879);
and UO_1141 (O_1141,N_9818,N_9967);
or UO_1142 (O_1142,N_9878,N_9995);
or UO_1143 (O_1143,N_9967,N_9949);
or UO_1144 (O_1144,N_9813,N_9878);
or UO_1145 (O_1145,N_9901,N_9998);
nand UO_1146 (O_1146,N_9959,N_9978);
nand UO_1147 (O_1147,N_9842,N_9844);
or UO_1148 (O_1148,N_9995,N_9999);
and UO_1149 (O_1149,N_9893,N_9965);
nand UO_1150 (O_1150,N_9935,N_9822);
or UO_1151 (O_1151,N_9872,N_9852);
nor UO_1152 (O_1152,N_9809,N_9906);
and UO_1153 (O_1153,N_9864,N_9936);
or UO_1154 (O_1154,N_9983,N_9838);
and UO_1155 (O_1155,N_9855,N_9974);
xnor UO_1156 (O_1156,N_9982,N_9868);
nor UO_1157 (O_1157,N_9860,N_9827);
nand UO_1158 (O_1158,N_9827,N_9972);
nor UO_1159 (O_1159,N_9891,N_9936);
nand UO_1160 (O_1160,N_9889,N_9830);
and UO_1161 (O_1161,N_9909,N_9877);
nand UO_1162 (O_1162,N_9935,N_9846);
or UO_1163 (O_1163,N_9863,N_9983);
nand UO_1164 (O_1164,N_9851,N_9825);
nand UO_1165 (O_1165,N_9930,N_9801);
xor UO_1166 (O_1166,N_9946,N_9880);
xnor UO_1167 (O_1167,N_9919,N_9925);
or UO_1168 (O_1168,N_9874,N_9800);
nand UO_1169 (O_1169,N_9831,N_9806);
nor UO_1170 (O_1170,N_9885,N_9830);
or UO_1171 (O_1171,N_9940,N_9887);
and UO_1172 (O_1172,N_9936,N_9952);
nand UO_1173 (O_1173,N_9976,N_9992);
nor UO_1174 (O_1174,N_9909,N_9985);
nand UO_1175 (O_1175,N_9834,N_9920);
nor UO_1176 (O_1176,N_9942,N_9922);
nand UO_1177 (O_1177,N_9883,N_9840);
nor UO_1178 (O_1178,N_9806,N_9873);
nor UO_1179 (O_1179,N_9862,N_9947);
xnor UO_1180 (O_1180,N_9989,N_9904);
or UO_1181 (O_1181,N_9948,N_9884);
nor UO_1182 (O_1182,N_9929,N_9896);
nand UO_1183 (O_1183,N_9829,N_9843);
and UO_1184 (O_1184,N_9917,N_9990);
xnor UO_1185 (O_1185,N_9934,N_9823);
or UO_1186 (O_1186,N_9927,N_9841);
or UO_1187 (O_1187,N_9983,N_9803);
or UO_1188 (O_1188,N_9896,N_9993);
nand UO_1189 (O_1189,N_9925,N_9807);
nand UO_1190 (O_1190,N_9923,N_9832);
nor UO_1191 (O_1191,N_9811,N_9860);
and UO_1192 (O_1192,N_9911,N_9850);
nand UO_1193 (O_1193,N_9806,N_9951);
and UO_1194 (O_1194,N_9837,N_9955);
xor UO_1195 (O_1195,N_9858,N_9942);
or UO_1196 (O_1196,N_9848,N_9951);
or UO_1197 (O_1197,N_9871,N_9814);
nand UO_1198 (O_1198,N_9941,N_9825);
and UO_1199 (O_1199,N_9966,N_9921);
nor UO_1200 (O_1200,N_9879,N_9816);
or UO_1201 (O_1201,N_9867,N_9894);
or UO_1202 (O_1202,N_9872,N_9968);
and UO_1203 (O_1203,N_9855,N_9916);
nor UO_1204 (O_1204,N_9997,N_9859);
nor UO_1205 (O_1205,N_9929,N_9838);
and UO_1206 (O_1206,N_9844,N_9816);
and UO_1207 (O_1207,N_9919,N_9817);
or UO_1208 (O_1208,N_9849,N_9863);
and UO_1209 (O_1209,N_9988,N_9873);
nor UO_1210 (O_1210,N_9970,N_9805);
or UO_1211 (O_1211,N_9943,N_9885);
nand UO_1212 (O_1212,N_9803,N_9937);
nand UO_1213 (O_1213,N_9844,N_9814);
or UO_1214 (O_1214,N_9804,N_9973);
or UO_1215 (O_1215,N_9852,N_9903);
nor UO_1216 (O_1216,N_9900,N_9932);
nand UO_1217 (O_1217,N_9836,N_9987);
nand UO_1218 (O_1218,N_9837,N_9989);
or UO_1219 (O_1219,N_9812,N_9980);
and UO_1220 (O_1220,N_9921,N_9973);
nor UO_1221 (O_1221,N_9818,N_9851);
nand UO_1222 (O_1222,N_9971,N_9873);
nand UO_1223 (O_1223,N_9975,N_9873);
and UO_1224 (O_1224,N_9941,N_9886);
and UO_1225 (O_1225,N_9937,N_9806);
nor UO_1226 (O_1226,N_9853,N_9970);
xnor UO_1227 (O_1227,N_9898,N_9866);
nor UO_1228 (O_1228,N_9989,N_9839);
or UO_1229 (O_1229,N_9858,N_9983);
or UO_1230 (O_1230,N_9971,N_9815);
nor UO_1231 (O_1231,N_9820,N_9893);
and UO_1232 (O_1232,N_9918,N_9914);
or UO_1233 (O_1233,N_9818,N_9835);
nor UO_1234 (O_1234,N_9868,N_9966);
nand UO_1235 (O_1235,N_9868,N_9944);
nor UO_1236 (O_1236,N_9982,N_9929);
or UO_1237 (O_1237,N_9891,N_9942);
or UO_1238 (O_1238,N_9927,N_9937);
and UO_1239 (O_1239,N_9946,N_9838);
and UO_1240 (O_1240,N_9986,N_9814);
nand UO_1241 (O_1241,N_9886,N_9841);
nor UO_1242 (O_1242,N_9870,N_9963);
or UO_1243 (O_1243,N_9939,N_9945);
nand UO_1244 (O_1244,N_9830,N_9929);
nor UO_1245 (O_1245,N_9968,N_9816);
and UO_1246 (O_1246,N_9923,N_9928);
nor UO_1247 (O_1247,N_9858,N_9879);
nand UO_1248 (O_1248,N_9940,N_9916);
nor UO_1249 (O_1249,N_9992,N_9809);
or UO_1250 (O_1250,N_9837,N_9885);
or UO_1251 (O_1251,N_9843,N_9892);
or UO_1252 (O_1252,N_9971,N_9984);
or UO_1253 (O_1253,N_9933,N_9812);
xnor UO_1254 (O_1254,N_9840,N_9805);
or UO_1255 (O_1255,N_9829,N_9990);
nor UO_1256 (O_1256,N_9887,N_9912);
nand UO_1257 (O_1257,N_9851,N_9884);
and UO_1258 (O_1258,N_9905,N_9870);
nand UO_1259 (O_1259,N_9864,N_9872);
nor UO_1260 (O_1260,N_9917,N_9920);
and UO_1261 (O_1261,N_9841,N_9924);
and UO_1262 (O_1262,N_9932,N_9935);
and UO_1263 (O_1263,N_9962,N_9850);
and UO_1264 (O_1264,N_9875,N_9933);
xnor UO_1265 (O_1265,N_9848,N_9809);
nand UO_1266 (O_1266,N_9980,N_9998);
nor UO_1267 (O_1267,N_9850,N_9826);
nand UO_1268 (O_1268,N_9887,N_9936);
or UO_1269 (O_1269,N_9914,N_9887);
and UO_1270 (O_1270,N_9881,N_9993);
or UO_1271 (O_1271,N_9897,N_9880);
nor UO_1272 (O_1272,N_9858,N_9951);
nand UO_1273 (O_1273,N_9939,N_9879);
or UO_1274 (O_1274,N_9876,N_9895);
nand UO_1275 (O_1275,N_9977,N_9910);
xnor UO_1276 (O_1276,N_9857,N_9831);
or UO_1277 (O_1277,N_9874,N_9871);
xor UO_1278 (O_1278,N_9840,N_9976);
nor UO_1279 (O_1279,N_9961,N_9900);
and UO_1280 (O_1280,N_9918,N_9988);
or UO_1281 (O_1281,N_9928,N_9869);
or UO_1282 (O_1282,N_9870,N_9965);
or UO_1283 (O_1283,N_9852,N_9814);
nand UO_1284 (O_1284,N_9948,N_9821);
or UO_1285 (O_1285,N_9887,N_9994);
nor UO_1286 (O_1286,N_9822,N_9942);
nor UO_1287 (O_1287,N_9901,N_9976);
nor UO_1288 (O_1288,N_9902,N_9842);
nand UO_1289 (O_1289,N_9806,N_9809);
nor UO_1290 (O_1290,N_9843,N_9906);
and UO_1291 (O_1291,N_9979,N_9893);
nand UO_1292 (O_1292,N_9986,N_9847);
and UO_1293 (O_1293,N_9933,N_9825);
and UO_1294 (O_1294,N_9985,N_9917);
or UO_1295 (O_1295,N_9884,N_9875);
or UO_1296 (O_1296,N_9905,N_9881);
nand UO_1297 (O_1297,N_9820,N_9956);
nand UO_1298 (O_1298,N_9824,N_9887);
and UO_1299 (O_1299,N_9958,N_9942);
nor UO_1300 (O_1300,N_9898,N_9997);
and UO_1301 (O_1301,N_9899,N_9999);
and UO_1302 (O_1302,N_9974,N_9902);
and UO_1303 (O_1303,N_9823,N_9864);
and UO_1304 (O_1304,N_9966,N_9861);
nor UO_1305 (O_1305,N_9863,N_9987);
or UO_1306 (O_1306,N_9917,N_9928);
nand UO_1307 (O_1307,N_9814,N_9845);
nand UO_1308 (O_1308,N_9953,N_9809);
or UO_1309 (O_1309,N_9938,N_9874);
and UO_1310 (O_1310,N_9918,N_9974);
nand UO_1311 (O_1311,N_9996,N_9857);
nor UO_1312 (O_1312,N_9922,N_9967);
or UO_1313 (O_1313,N_9866,N_9832);
nand UO_1314 (O_1314,N_9813,N_9883);
nand UO_1315 (O_1315,N_9888,N_9805);
nand UO_1316 (O_1316,N_9927,N_9847);
or UO_1317 (O_1317,N_9805,N_9955);
and UO_1318 (O_1318,N_9970,N_9812);
nor UO_1319 (O_1319,N_9815,N_9992);
and UO_1320 (O_1320,N_9959,N_9976);
nand UO_1321 (O_1321,N_9931,N_9906);
nand UO_1322 (O_1322,N_9835,N_9947);
nand UO_1323 (O_1323,N_9984,N_9961);
or UO_1324 (O_1324,N_9800,N_9911);
nor UO_1325 (O_1325,N_9812,N_9925);
nor UO_1326 (O_1326,N_9941,N_9894);
nor UO_1327 (O_1327,N_9828,N_9974);
nor UO_1328 (O_1328,N_9884,N_9826);
or UO_1329 (O_1329,N_9999,N_9851);
xor UO_1330 (O_1330,N_9938,N_9902);
or UO_1331 (O_1331,N_9821,N_9877);
nand UO_1332 (O_1332,N_9806,N_9987);
nor UO_1333 (O_1333,N_9926,N_9859);
and UO_1334 (O_1334,N_9943,N_9873);
and UO_1335 (O_1335,N_9893,N_9909);
or UO_1336 (O_1336,N_9945,N_9809);
xor UO_1337 (O_1337,N_9898,N_9868);
nor UO_1338 (O_1338,N_9933,N_9881);
or UO_1339 (O_1339,N_9877,N_9974);
or UO_1340 (O_1340,N_9811,N_9804);
or UO_1341 (O_1341,N_9896,N_9863);
nand UO_1342 (O_1342,N_9979,N_9924);
nand UO_1343 (O_1343,N_9886,N_9925);
nor UO_1344 (O_1344,N_9925,N_9803);
xnor UO_1345 (O_1345,N_9976,N_9966);
nand UO_1346 (O_1346,N_9908,N_9931);
nor UO_1347 (O_1347,N_9855,N_9869);
and UO_1348 (O_1348,N_9833,N_9892);
or UO_1349 (O_1349,N_9965,N_9970);
nor UO_1350 (O_1350,N_9838,N_9901);
or UO_1351 (O_1351,N_9934,N_9907);
and UO_1352 (O_1352,N_9976,N_9978);
nor UO_1353 (O_1353,N_9917,N_9992);
xnor UO_1354 (O_1354,N_9829,N_9813);
nor UO_1355 (O_1355,N_9895,N_9924);
or UO_1356 (O_1356,N_9946,N_9844);
and UO_1357 (O_1357,N_9934,N_9855);
and UO_1358 (O_1358,N_9856,N_9901);
and UO_1359 (O_1359,N_9918,N_9938);
nand UO_1360 (O_1360,N_9964,N_9947);
nor UO_1361 (O_1361,N_9810,N_9822);
nor UO_1362 (O_1362,N_9965,N_9815);
or UO_1363 (O_1363,N_9877,N_9973);
or UO_1364 (O_1364,N_9891,N_9828);
or UO_1365 (O_1365,N_9914,N_9913);
or UO_1366 (O_1366,N_9963,N_9864);
nor UO_1367 (O_1367,N_9857,N_9887);
or UO_1368 (O_1368,N_9839,N_9971);
nand UO_1369 (O_1369,N_9807,N_9833);
or UO_1370 (O_1370,N_9943,N_9833);
and UO_1371 (O_1371,N_9863,N_9985);
and UO_1372 (O_1372,N_9970,N_9830);
nand UO_1373 (O_1373,N_9887,N_9915);
or UO_1374 (O_1374,N_9908,N_9987);
or UO_1375 (O_1375,N_9970,N_9840);
nand UO_1376 (O_1376,N_9912,N_9947);
and UO_1377 (O_1377,N_9852,N_9961);
and UO_1378 (O_1378,N_9926,N_9805);
and UO_1379 (O_1379,N_9957,N_9814);
nand UO_1380 (O_1380,N_9821,N_9892);
and UO_1381 (O_1381,N_9825,N_9918);
xnor UO_1382 (O_1382,N_9922,N_9803);
xnor UO_1383 (O_1383,N_9800,N_9843);
nor UO_1384 (O_1384,N_9976,N_9963);
nand UO_1385 (O_1385,N_9927,N_9973);
nor UO_1386 (O_1386,N_9816,N_9901);
and UO_1387 (O_1387,N_9812,N_9913);
nand UO_1388 (O_1388,N_9944,N_9990);
or UO_1389 (O_1389,N_9963,N_9896);
nor UO_1390 (O_1390,N_9997,N_9855);
and UO_1391 (O_1391,N_9861,N_9833);
nand UO_1392 (O_1392,N_9939,N_9813);
xnor UO_1393 (O_1393,N_9904,N_9938);
nand UO_1394 (O_1394,N_9978,N_9927);
nor UO_1395 (O_1395,N_9959,N_9895);
nor UO_1396 (O_1396,N_9901,N_9956);
or UO_1397 (O_1397,N_9920,N_9987);
nand UO_1398 (O_1398,N_9942,N_9827);
nor UO_1399 (O_1399,N_9921,N_9906);
and UO_1400 (O_1400,N_9805,N_9809);
nand UO_1401 (O_1401,N_9917,N_9934);
or UO_1402 (O_1402,N_9947,N_9927);
or UO_1403 (O_1403,N_9981,N_9875);
or UO_1404 (O_1404,N_9996,N_9885);
and UO_1405 (O_1405,N_9933,N_9871);
nand UO_1406 (O_1406,N_9941,N_9908);
and UO_1407 (O_1407,N_9805,N_9947);
nor UO_1408 (O_1408,N_9991,N_9989);
or UO_1409 (O_1409,N_9985,N_9931);
nand UO_1410 (O_1410,N_9835,N_9913);
xor UO_1411 (O_1411,N_9844,N_9922);
nor UO_1412 (O_1412,N_9822,N_9837);
and UO_1413 (O_1413,N_9981,N_9971);
and UO_1414 (O_1414,N_9898,N_9846);
nand UO_1415 (O_1415,N_9927,N_9819);
and UO_1416 (O_1416,N_9931,N_9895);
or UO_1417 (O_1417,N_9965,N_9897);
and UO_1418 (O_1418,N_9898,N_9933);
xor UO_1419 (O_1419,N_9854,N_9974);
and UO_1420 (O_1420,N_9958,N_9857);
nand UO_1421 (O_1421,N_9819,N_9969);
or UO_1422 (O_1422,N_9867,N_9956);
nor UO_1423 (O_1423,N_9903,N_9938);
nand UO_1424 (O_1424,N_9818,N_9845);
nand UO_1425 (O_1425,N_9854,N_9965);
nor UO_1426 (O_1426,N_9936,N_9920);
nor UO_1427 (O_1427,N_9934,N_9849);
xor UO_1428 (O_1428,N_9923,N_9805);
or UO_1429 (O_1429,N_9919,N_9838);
and UO_1430 (O_1430,N_9975,N_9947);
nor UO_1431 (O_1431,N_9990,N_9849);
and UO_1432 (O_1432,N_9936,N_9960);
and UO_1433 (O_1433,N_9808,N_9989);
nor UO_1434 (O_1434,N_9903,N_9877);
or UO_1435 (O_1435,N_9980,N_9968);
and UO_1436 (O_1436,N_9952,N_9884);
nor UO_1437 (O_1437,N_9987,N_9952);
nand UO_1438 (O_1438,N_9980,N_9981);
nand UO_1439 (O_1439,N_9898,N_9958);
nand UO_1440 (O_1440,N_9894,N_9981);
nor UO_1441 (O_1441,N_9855,N_9872);
xnor UO_1442 (O_1442,N_9929,N_9983);
and UO_1443 (O_1443,N_9916,N_9995);
nand UO_1444 (O_1444,N_9804,N_9929);
nor UO_1445 (O_1445,N_9813,N_9879);
or UO_1446 (O_1446,N_9961,N_9915);
or UO_1447 (O_1447,N_9978,N_9922);
and UO_1448 (O_1448,N_9978,N_9967);
nor UO_1449 (O_1449,N_9865,N_9976);
nand UO_1450 (O_1450,N_9936,N_9974);
and UO_1451 (O_1451,N_9888,N_9961);
or UO_1452 (O_1452,N_9938,N_9820);
or UO_1453 (O_1453,N_9922,N_9927);
nand UO_1454 (O_1454,N_9856,N_9807);
nor UO_1455 (O_1455,N_9807,N_9804);
nor UO_1456 (O_1456,N_9936,N_9965);
and UO_1457 (O_1457,N_9938,N_9895);
nor UO_1458 (O_1458,N_9876,N_9926);
nor UO_1459 (O_1459,N_9816,N_9839);
or UO_1460 (O_1460,N_9809,N_9981);
xnor UO_1461 (O_1461,N_9933,N_9810);
nor UO_1462 (O_1462,N_9814,N_9946);
or UO_1463 (O_1463,N_9853,N_9934);
nand UO_1464 (O_1464,N_9824,N_9837);
and UO_1465 (O_1465,N_9977,N_9879);
xnor UO_1466 (O_1466,N_9833,N_9922);
and UO_1467 (O_1467,N_9919,N_9821);
nor UO_1468 (O_1468,N_9912,N_9907);
xor UO_1469 (O_1469,N_9876,N_9937);
and UO_1470 (O_1470,N_9949,N_9972);
and UO_1471 (O_1471,N_9968,N_9928);
or UO_1472 (O_1472,N_9821,N_9867);
xnor UO_1473 (O_1473,N_9814,N_9904);
nand UO_1474 (O_1474,N_9950,N_9839);
nand UO_1475 (O_1475,N_9819,N_9989);
nor UO_1476 (O_1476,N_9923,N_9800);
or UO_1477 (O_1477,N_9855,N_9962);
nor UO_1478 (O_1478,N_9890,N_9995);
or UO_1479 (O_1479,N_9893,N_9870);
or UO_1480 (O_1480,N_9984,N_9925);
nor UO_1481 (O_1481,N_9968,N_9938);
or UO_1482 (O_1482,N_9990,N_9860);
nand UO_1483 (O_1483,N_9991,N_9949);
nand UO_1484 (O_1484,N_9837,N_9865);
and UO_1485 (O_1485,N_9988,N_9910);
or UO_1486 (O_1486,N_9967,N_9929);
nor UO_1487 (O_1487,N_9992,N_9872);
and UO_1488 (O_1488,N_9845,N_9977);
xnor UO_1489 (O_1489,N_9966,N_9945);
nand UO_1490 (O_1490,N_9999,N_9842);
or UO_1491 (O_1491,N_9880,N_9852);
nor UO_1492 (O_1492,N_9941,N_9976);
nand UO_1493 (O_1493,N_9896,N_9947);
or UO_1494 (O_1494,N_9973,N_9974);
nand UO_1495 (O_1495,N_9856,N_9991);
or UO_1496 (O_1496,N_9831,N_9991);
nor UO_1497 (O_1497,N_9993,N_9844);
nand UO_1498 (O_1498,N_9818,N_9961);
xnor UO_1499 (O_1499,N_9987,N_9878);
endmodule