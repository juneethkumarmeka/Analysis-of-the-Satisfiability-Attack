module basic_500_3000_500_30_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_68,In_342);
and U1 (N_1,In_229,In_368);
nand U2 (N_2,In_121,In_177);
and U3 (N_3,In_258,In_377);
nand U4 (N_4,In_154,In_433);
and U5 (N_5,In_458,In_244);
nor U6 (N_6,In_348,In_33);
or U7 (N_7,In_274,In_242);
nor U8 (N_8,In_98,In_115);
or U9 (N_9,In_145,In_210);
nor U10 (N_10,In_496,In_487);
nand U11 (N_11,In_40,In_142);
nor U12 (N_12,In_259,In_223);
and U13 (N_13,In_466,In_343);
or U14 (N_14,In_42,In_125);
nand U15 (N_15,In_491,In_234);
or U16 (N_16,In_139,In_389);
nand U17 (N_17,In_287,In_416);
nor U18 (N_18,In_448,In_134);
nand U19 (N_19,In_245,In_489);
nor U20 (N_20,In_320,In_69);
nor U21 (N_21,In_216,In_335);
nand U22 (N_22,In_122,In_429);
and U23 (N_23,In_301,In_249);
and U24 (N_24,In_441,In_0);
and U25 (N_25,In_374,In_332);
or U26 (N_26,In_240,In_372);
or U27 (N_27,In_472,In_225);
and U28 (N_28,In_326,In_251);
nor U29 (N_29,In_17,In_435);
nand U30 (N_30,In_172,In_285);
nor U31 (N_31,In_41,In_200);
nor U32 (N_32,In_175,In_19);
nor U33 (N_33,In_45,In_366);
nor U34 (N_34,In_463,In_347);
or U35 (N_35,In_462,In_10);
or U36 (N_36,In_213,In_163);
or U37 (N_37,In_336,In_203);
and U38 (N_38,In_208,In_334);
nor U39 (N_39,In_392,In_298);
nor U40 (N_40,In_432,In_35);
nand U41 (N_41,In_202,In_191);
or U42 (N_42,In_243,In_188);
nand U43 (N_43,In_246,In_302);
and U44 (N_44,In_367,In_194);
nor U45 (N_45,In_230,In_488);
nand U46 (N_46,In_384,In_97);
and U47 (N_47,In_470,In_476);
nor U48 (N_48,In_206,In_63);
nor U49 (N_49,In_211,In_27);
or U50 (N_50,In_140,In_165);
or U51 (N_51,In_212,In_410);
nor U52 (N_52,In_80,In_456);
nand U53 (N_53,In_411,In_397);
nor U54 (N_54,In_486,In_179);
and U55 (N_55,In_157,In_196);
and U56 (N_56,In_484,In_102);
nor U57 (N_57,In_32,In_21);
nand U58 (N_58,In_481,In_468);
or U59 (N_59,In_493,In_113);
and U60 (N_60,In_127,In_350);
nor U61 (N_61,In_215,In_281);
and U62 (N_62,In_262,In_232);
nand U63 (N_63,In_47,In_296);
xor U64 (N_64,In_152,In_446);
nor U65 (N_65,In_1,In_44);
and U66 (N_66,In_166,In_183);
and U67 (N_67,In_478,In_461);
nor U68 (N_68,In_290,In_239);
nand U69 (N_69,In_14,In_138);
nand U70 (N_70,In_352,In_109);
nor U71 (N_71,In_137,In_319);
nor U72 (N_72,In_357,In_293);
nand U73 (N_73,In_222,In_445);
xor U74 (N_74,In_57,In_220);
and U75 (N_75,In_112,In_387);
nand U76 (N_76,In_497,In_146);
or U77 (N_77,In_317,In_271);
nor U78 (N_78,In_116,In_226);
and U79 (N_79,In_20,In_252);
nand U80 (N_80,In_195,In_304);
nand U81 (N_81,In_54,In_419);
or U82 (N_82,In_457,In_403);
nor U83 (N_83,In_214,In_64);
or U84 (N_84,In_120,In_380);
nand U85 (N_85,In_451,In_393);
or U86 (N_86,In_438,In_104);
nor U87 (N_87,In_442,In_60);
or U88 (N_88,In_75,In_406);
nand U89 (N_89,In_117,In_371);
and U90 (N_90,In_375,In_305);
or U91 (N_91,In_114,In_74);
or U92 (N_92,In_404,In_82);
nand U93 (N_93,In_201,In_159);
and U94 (N_94,In_358,In_382);
or U95 (N_95,In_286,In_428);
or U96 (N_96,In_464,In_53);
xnor U97 (N_97,In_363,In_189);
xor U98 (N_98,In_50,In_492);
nor U99 (N_99,In_217,In_198);
nand U100 (N_100,In_36,In_339);
nor U101 (N_101,In_383,In_409);
nand U102 (N_102,In_401,N_42);
nor U103 (N_103,N_11,In_241);
nand U104 (N_104,In_313,In_48);
nand U105 (N_105,In_153,In_71);
and U106 (N_106,In_67,N_56);
or U107 (N_107,In_454,In_221);
nor U108 (N_108,In_431,In_61);
nand U109 (N_109,N_94,In_303);
nor U110 (N_110,N_84,In_427);
nor U111 (N_111,In_280,In_425);
and U112 (N_112,In_181,In_379);
or U113 (N_113,In_93,N_86);
nand U114 (N_114,In_37,In_362);
nand U115 (N_115,In_38,N_16);
nand U116 (N_116,N_10,In_133);
nand U117 (N_117,In_130,In_260);
and U118 (N_118,In_386,N_0);
nor U119 (N_119,In_43,In_297);
nand U120 (N_120,In_325,N_51);
nand U121 (N_121,N_70,In_345);
nand U122 (N_122,In_76,N_23);
xor U123 (N_123,In_340,N_64);
and U124 (N_124,In_250,N_58);
and U125 (N_125,In_88,In_308);
nor U126 (N_126,N_98,In_311);
and U127 (N_127,In_227,In_381);
nor U128 (N_128,N_17,In_209);
nand U129 (N_129,In_439,In_118);
or U130 (N_130,In_277,In_312);
and U131 (N_131,N_14,In_465);
nand U132 (N_132,In_30,In_228);
and U133 (N_133,In_423,In_24);
and U134 (N_134,In_49,In_89);
and U135 (N_135,In_388,N_97);
or U136 (N_136,In_34,N_40);
nor U137 (N_137,In_158,In_59);
and U138 (N_138,In_25,In_365);
nand U139 (N_139,In_498,N_39);
nand U140 (N_140,In_219,N_43);
nor U141 (N_141,In_204,In_180);
nor U142 (N_142,In_72,In_52);
or U143 (N_143,N_92,In_405);
nand U144 (N_144,In_176,In_96);
and U145 (N_145,In_449,In_376);
or U146 (N_146,In_4,In_328);
or U147 (N_147,In_337,In_309);
nor U148 (N_148,In_205,In_103);
nand U149 (N_149,In_276,In_450);
nand U150 (N_150,N_83,N_29);
nand U151 (N_151,In_331,N_19);
or U152 (N_152,N_82,In_105);
nor U153 (N_153,In_197,In_90);
and U154 (N_154,N_95,In_174);
and U155 (N_155,In_394,In_207);
and U156 (N_156,In_467,In_126);
xnor U157 (N_157,N_15,N_72);
and U158 (N_158,In_391,N_7);
nand U159 (N_159,In_257,In_12);
nor U160 (N_160,In_9,N_13);
nand U161 (N_161,In_94,In_400);
or U162 (N_162,In_355,N_45);
nand U163 (N_163,In_485,N_91);
nor U164 (N_164,In_344,In_224);
and U165 (N_165,In_135,N_34);
or U166 (N_166,In_272,In_417);
and U167 (N_167,In_407,In_370);
nand U168 (N_168,In_263,In_95);
and U169 (N_169,In_360,N_93);
or U170 (N_170,In_495,In_474);
nand U171 (N_171,N_85,In_70);
and U172 (N_172,In_422,In_73);
and U173 (N_173,N_5,N_31);
nand U174 (N_174,In_300,In_396);
nand U175 (N_175,In_13,In_81);
or U176 (N_176,In_101,In_291);
nand U177 (N_177,In_143,In_131);
or U178 (N_178,In_6,In_385);
and U179 (N_179,N_90,In_412);
nor U180 (N_180,In_231,N_55);
or U181 (N_181,In_255,In_106);
nand U182 (N_182,In_256,N_21);
nor U183 (N_183,In_141,N_52);
nor U184 (N_184,In_238,In_306);
nand U185 (N_185,In_494,In_475);
or U186 (N_186,N_18,N_36);
and U187 (N_187,In_346,In_329);
nor U188 (N_188,In_269,N_33);
and U189 (N_189,In_264,In_235);
xnor U190 (N_190,In_268,In_233);
nand U191 (N_191,In_15,In_150);
nand U192 (N_192,N_61,N_89);
nor U193 (N_193,In_499,In_430);
and U194 (N_194,N_26,In_399);
nor U195 (N_195,In_23,In_237);
and U196 (N_196,In_185,In_295);
nand U197 (N_197,In_26,In_341);
or U198 (N_198,In_84,N_41);
nor U199 (N_199,In_408,N_4);
nor U200 (N_200,N_54,N_119);
and U201 (N_201,In_164,N_178);
or U202 (N_202,In_420,N_194);
or U203 (N_203,In_155,In_167);
nor U204 (N_204,In_86,N_32);
or U205 (N_205,N_116,N_109);
xnor U206 (N_206,N_197,N_101);
nand U207 (N_207,N_102,N_187);
or U208 (N_208,N_117,In_161);
or U209 (N_209,N_38,In_193);
or U210 (N_210,N_155,N_183);
or U211 (N_211,N_190,N_134);
or U212 (N_212,N_9,In_190);
nand U213 (N_213,In_349,N_171);
or U214 (N_214,N_126,In_436);
and U215 (N_215,N_73,In_292);
nand U216 (N_216,N_140,In_354);
and U217 (N_217,In_87,N_112);
and U218 (N_218,In_483,In_390);
nand U219 (N_219,In_279,In_353);
or U220 (N_220,In_247,In_92);
or U221 (N_221,In_55,In_16);
or U222 (N_222,N_199,In_3);
or U223 (N_223,N_141,N_96);
nand U224 (N_224,In_147,N_142);
nor U225 (N_225,In_413,In_266);
nand U226 (N_226,N_123,N_154);
nor U227 (N_227,In_182,In_192);
and U228 (N_228,In_278,N_57);
nand U229 (N_229,In_471,In_482);
xor U230 (N_230,In_170,In_2);
nor U231 (N_231,N_20,In_169);
nand U232 (N_232,N_2,In_310);
or U233 (N_233,In_254,N_146);
nor U234 (N_234,N_69,In_22);
or U235 (N_235,In_168,In_330);
and U236 (N_236,In_111,N_156);
nand U237 (N_237,N_120,In_378);
and U238 (N_238,In_148,In_58);
nor U239 (N_239,N_193,N_145);
nor U240 (N_240,N_107,N_113);
nand U241 (N_241,N_147,N_65);
or U242 (N_242,N_138,N_122);
and U243 (N_243,N_165,N_106);
nand U244 (N_244,In_267,In_288);
nand U245 (N_245,N_164,In_66);
nand U246 (N_246,In_453,In_373);
nor U247 (N_247,In_119,N_63);
nand U248 (N_248,N_37,N_53);
or U249 (N_249,In_294,N_182);
or U250 (N_250,In_83,In_369);
and U251 (N_251,In_187,N_127);
nand U252 (N_252,N_172,In_424);
nand U253 (N_253,N_128,In_39);
nor U254 (N_254,N_79,In_395);
nand U255 (N_255,N_77,In_473);
nor U256 (N_256,In_173,In_356);
and U257 (N_257,In_108,In_56);
or U258 (N_258,N_151,N_175);
or U259 (N_259,In_469,N_196);
or U260 (N_260,N_169,In_459);
nor U261 (N_261,In_99,N_103);
or U262 (N_262,N_46,In_46);
nor U263 (N_263,N_62,In_129);
xnor U264 (N_264,N_135,N_35);
nor U265 (N_265,N_44,In_8);
or U266 (N_266,N_179,N_1);
nand U267 (N_267,N_144,N_27);
and U268 (N_268,In_426,In_316);
nand U269 (N_269,N_191,In_398);
nor U270 (N_270,N_80,In_414);
or U271 (N_271,In_289,In_107);
nand U272 (N_272,In_444,N_105);
nand U273 (N_273,N_6,N_137);
nor U274 (N_274,In_136,N_192);
nor U275 (N_275,N_71,N_150);
and U276 (N_276,N_115,N_99);
nor U277 (N_277,In_65,N_78);
nand U278 (N_278,In_5,In_443);
nor U279 (N_279,N_131,In_479);
or U280 (N_280,N_49,In_315);
or U281 (N_281,In_434,N_153);
nor U282 (N_282,N_124,N_139);
or U283 (N_283,In_11,N_67);
or U284 (N_284,In_447,N_157);
and U285 (N_285,In_490,N_184);
or U286 (N_286,N_185,In_151);
nand U287 (N_287,N_110,N_162);
and U288 (N_288,In_477,N_176);
nor U289 (N_289,N_166,N_152);
and U290 (N_290,In_18,In_124);
nor U291 (N_291,N_114,In_314);
or U292 (N_292,In_452,In_364);
nand U293 (N_293,N_177,N_76);
or U294 (N_294,N_163,N_75);
and U295 (N_295,In_440,In_359);
or U296 (N_296,In_265,N_186);
or U297 (N_297,N_30,In_110);
nand U298 (N_298,N_148,In_123);
nand U299 (N_299,In_283,In_144);
or U300 (N_300,N_195,N_292);
nor U301 (N_301,In_51,In_275);
nor U302 (N_302,N_48,N_130);
nor U303 (N_303,In_418,In_437);
or U304 (N_304,N_180,N_261);
nand U305 (N_305,N_188,N_104);
nand U306 (N_306,In_324,N_244);
nand U307 (N_307,N_291,N_158);
nor U308 (N_308,In_78,In_29);
nor U309 (N_309,N_216,In_162);
xnor U310 (N_310,N_287,N_210);
or U311 (N_311,In_62,N_241);
nor U312 (N_312,In_184,N_219);
nor U313 (N_313,N_236,N_253);
nand U314 (N_314,In_455,N_222);
or U315 (N_315,In_333,In_178);
nand U316 (N_316,In_323,N_280);
nor U317 (N_317,N_267,N_239);
nor U318 (N_318,N_270,In_460);
nor U319 (N_319,In_31,N_259);
or U320 (N_320,N_202,N_294);
and U321 (N_321,N_59,N_235);
and U322 (N_322,N_231,N_159);
and U323 (N_323,N_225,N_240);
and U324 (N_324,N_232,N_257);
and U325 (N_325,N_262,In_149);
and U326 (N_326,In_132,N_269);
or U327 (N_327,N_220,N_246);
nor U328 (N_328,N_8,N_170);
and U329 (N_329,N_295,N_136);
and U330 (N_330,N_296,N_254);
or U331 (N_331,N_25,N_255);
or U332 (N_332,N_22,N_268);
nor U333 (N_333,N_108,N_214);
and U334 (N_334,In_160,N_242);
nor U335 (N_335,In_351,N_266);
and U336 (N_336,N_208,In_236);
or U337 (N_337,N_251,N_181);
or U338 (N_338,N_260,N_207);
nand U339 (N_339,N_200,In_361);
nor U340 (N_340,N_263,N_160);
or U341 (N_341,N_3,In_218);
nor U342 (N_342,N_252,N_60);
or U343 (N_343,N_284,N_283);
and U344 (N_344,N_226,In_322);
and U345 (N_345,N_189,N_47);
nand U346 (N_346,N_74,In_270);
or U347 (N_347,N_87,N_204);
nor U348 (N_348,N_198,N_211);
and U349 (N_349,In_28,N_230);
nand U350 (N_350,N_227,N_223);
nand U351 (N_351,N_174,In_282);
or U352 (N_352,N_274,In_307);
nand U353 (N_353,N_133,N_272);
and U354 (N_354,N_233,N_281);
and U355 (N_355,N_173,In_253);
nand U356 (N_356,In_273,In_415);
and U357 (N_357,N_247,N_276);
nor U358 (N_358,In_261,In_171);
or U359 (N_359,N_203,N_68);
or U360 (N_360,N_149,N_118);
nand U361 (N_361,N_111,In_402);
nand U362 (N_362,N_249,N_217);
or U363 (N_363,N_161,N_24);
nand U364 (N_364,N_279,N_221);
and U365 (N_365,In_156,N_243);
or U366 (N_366,N_278,In_321);
and U367 (N_367,N_237,In_91);
xor U368 (N_368,N_121,N_206);
or U369 (N_369,N_81,N_12);
or U370 (N_370,N_224,N_212);
nand U371 (N_371,N_28,In_318);
or U372 (N_372,N_264,N_298);
or U373 (N_373,N_290,In_7);
or U374 (N_374,N_100,In_299);
and U375 (N_375,N_209,In_480);
nand U376 (N_376,N_228,In_327);
nand U377 (N_377,In_284,N_229);
and U378 (N_378,N_258,In_77);
and U379 (N_379,N_277,In_128);
and U380 (N_380,N_289,In_100);
and U381 (N_381,N_66,N_299);
or U382 (N_382,N_88,N_168);
nor U383 (N_383,N_286,N_271);
or U384 (N_384,In_248,N_256);
and U385 (N_385,N_129,N_265);
xnor U386 (N_386,N_132,N_205);
nand U387 (N_387,In_79,N_245);
and U388 (N_388,N_250,In_421);
or U389 (N_389,N_215,N_125);
nor U390 (N_390,N_293,N_167);
or U391 (N_391,N_275,N_285);
nand U392 (N_392,N_248,N_201);
or U393 (N_393,N_288,N_297);
or U394 (N_394,N_234,N_218);
and U395 (N_395,In_186,N_50);
and U396 (N_396,In_199,N_143);
and U397 (N_397,In_338,N_213);
and U398 (N_398,In_85,N_273);
or U399 (N_399,N_238,N_282);
or U400 (N_400,N_378,N_388);
nand U401 (N_401,N_382,N_399);
or U402 (N_402,N_352,N_335);
or U403 (N_403,N_369,N_317);
nor U404 (N_404,N_384,N_365);
and U405 (N_405,N_398,N_303);
and U406 (N_406,N_306,N_336);
or U407 (N_407,N_389,N_372);
nand U408 (N_408,N_391,N_387);
or U409 (N_409,N_377,N_311);
nand U410 (N_410,N_357,N_380);
nor U411 (N_411,N_326,N_361);
and U412 (N_412,N_337,N_310);
and U413 (N_413,N_343,N_325);
nand U414 (N_414,N_355,N_308);
and U415 (N_415,N_373,N_386);
and U416 (N_416,N_359,N_395);
and U417 (N_417,N_323,N_312);
and U418 (N_418,N_360,N_397);
and U419 (N_419,N_385,N_338);
or U420 (N_420,N_362,N_364);
or U421 (N_421,N_342,N_307);
nand U422 (N_422,N_327,N_328);
xor U423 (N_423,N_370,N_374);
nand U424 (N_424,N_381,N_315);
or U425 (N_425,N_390,N_316);
nor U426 (N_426,N_319,N_375);
and U427 (N_427,N_353,N_333);
nand U428 (N_428,N_366,N_383);
nand U429 (N_429,N_349,N_330);
or U430 (N_430,N_301,N_332);
nor U431 (N_431,N_367,N_329);
nand U432 (N_432,N_347,N_339);
nand U433 (N_433,N_321,N_322);
or U434 (N_434,N_345,N_302);
and U435 (N_435,N_348,N_376);
nand U436 (N_436,N_392,N_371);
and U437 (N_437,N_320,N_351);
nand U438 (N_438,N_305,N_313);
and U439 (N_439,N_340,N_300);
nor U440 (N_440,N_309,N_368);
nor U441 (N_441,N_346,N_356);
and U442 (N_442,N_354,N_396);
or U443 (N_443,N_394,N_341);
or U444 (N_444,N_379,N_350);
nor U445 (N_445,N_393,N_318);
xor U446 (N_446,N_304,N_314);
nand U447 (N_447,N_344,N_363);
xnor U448 (N_448,N_324,N_358);
nand U449 (N_449,N_334,N_331);
or U450 (N_450,N_312,N_390);
and U451 (N_451,N_326,N_393);
and U452 (N_452,N_381,N_332);
xor U453 (N_453,N_399,N_335);
and U454 (N_454,N_301,N_312);
or U455 (N_455,N_368,N_306);
nor U456 (N_456,N_385,N_359);
nand U457 (N_457,N_396,N_346);
nand U458 (N_458,N_330,N_395);
and U459 (N_459,N_340,N_383);
and U460 (N_460,N_395,N_305);
or U461 (N_461,N_320,N_312);
and U462 (N_462,N_376,N_395);
nor U463 (N_463,N_336,N_316);
or U464 (N_464,N_393,N_377);
nor U465 (N_465,N_333,N_330);
or U466 (N_466,N_369,N_352);
or U467 (N_467,N_357,N_373);
and U468 (N_468,N_382,N_397);
or U469 (N_469,N_304,N_319);
or U470 (N_470,N_356,N_318);
nand U471 (N_471,N_392,N_314);
or U472 (N_472,N_387,N_350);
nor U473 (N_473,N_342,N_321);
nand U474 (N_474,N_379,N_398);
nand U475 (N_475,N_363,N_339);
and U476 (N_476,N_308,N_325);
nor U477 (N_477,N_300,N_364);
nand U478 (N_478,N_355,N_362);
and U479 (N_479,N_363,N_347);
nand U480 (N_480,N_381,N_394);
nand U481 (N_481,N_336,N_362);
or U482 (N_482,N_340,N_334);
nand U483 (N_483,N_376,N_342);
or U484 (N_484,N_390,N_388);
nand U485 (N_485,N_321,N_398);
and U486 (N_486,N_388,N_377);
xor U487 (N_487,N_306,N_318);
nand U488 (N_488,N_374,N_381);
nor U489 (N_489,N_386,N_309);
nand U490 (N_490,N_368,N_316);
nor U491 (N_491,N_314,N_326);
nand U492 (N_492,N_371,N_301);
nand U493 (N_493,N_304,N_321);
and U494 (N_494,N_316,N_377);
nand U495 (N_495,N_327,N_329);
or U496 (N_496,N_302,N_335);
and U497 (N_497,N_353,N_384);
nor U498 (N_498,N_333,N_377);
xor U499 (N_499,N_340,N_355);
nor U500 (N_500,N_456,N_494);
nor U501 (N_501,N_458,N_482);
xor U502 (N_502,N_438,N_448);
and U503 (N_503,N_406,N_404);
and U504 (N_504,N_410,N_434);
nor U505 (N_505,N_450,N_496);
and U506 (N_506,N_408,N_469);
and U507 (N_507,N_433,N_427);
and U508 (N_508,N_431,N_444);
nand U509 (N_509,N_471,N_480);
nand U510 (N_510,N_467,N_409);
nand U511 (N_511,N_403,N_483);
nand U512 (N_512,N_489,N_417);
or U513 (N_513,N_420,N_412);
nor U514 (N_514,N_475,N_439);
and U515 (N_515,N_415,N_421);
nand U516 (N_516,N_457,N_424);
or U517 (N_517,N_414,N_432);
or U518 (N_518,N_495,N_487);
and U519 (N_519,N_479,N_472);
and U520 (N_520,N_402,N_484);
nor U521 (N_521,N_446,N_419);
or U522 (N_522,N_468,N_430);
nor U523 (N_523,N_499,N_443);
nand U524 (N_524,N_455,N_413);
nor U525 (N_525,N_493,N_465);
or U526 (N_526,N_400,N_490);
nand U527 (N_527,N_411,N_474);
or U528 (N_528,N_473,N_442);
nor U529 (N_529,N_426,N_454);
or U530 (N_530,N_436,N_435);
and U531 (N_531,N_491,N_441);
or U532 (N_532,N_477,N_425);
nand U533 (N_533,N_449,N_451);
nand U534 (N_534,N_422,N_488);
or U535 (N_535,N_447,N_498);
or U536 (N_536,N_429,N_407);
or U537 (N_537,N_492,N_486);
nand U538 (N_538,N_428,N_440);
and U539 (N_539,N_485,N_401);
nand U540 (N_540,N_481,N_466);
and U541 (N_541,N_418,N_459);
nand U542 (N_542,N_423,N_497);
nor U543 (N_543,N_462,N_445);
and U544 (N_544,N_461,N_463);
nand U545 (N_545,N_405,N_437);
or U546 (N_546,N_478,N_464);
nand U547 (N_547,N_460,N_416);
and U548 (N_548,N_452,N_476);
and U549 (N_549,N_453,N_470);
or U550 (N_550,N_453,N_463);
and U551 (N_551,N_489,N_423);
and U552 (N_552,N_464,N_410);
or U553 (N_553,N_442,N_423);
or U554 (N_554,N_450,N_457);
or U555 (N_555,N_453,N_487);
and U556 (N_556,N_499,N_488);
nand U557 (N_557,N_498,N_463);
or U558 (N_558,N_455,N_462);
and U559 (N_559,N_467,N_490);
xnor U560 (N_560,N_486,N_457);
nand U561 (N_561,N_414,N_479);
nor U562 (N_562,N_400,N_463);
or U563 (N_563,N_440,N_470);
nor U564 (N_564,N_438,N_440);
nand U565 (N_565,N_417,N_494);
nand U566 (N_566,N_491,N_429);
nor U567 (N_567,N_409,N_440);
and U568 (N_568,N_453,N_456);
nand U569 (N_569,N_438,N_436);
and U570 (N_570,N_467,N_427);
nand U571 (N_571,N_473,N_460);
nand U572 (N_572,N_477,N_426);
or U573 (N_573,N_475,N_420);
nand U574 (N_574,N_450,N_475);
or U575 (N_575,N_405,N_413);
nand U576 (N_576,N_473,N_428);
or U577 (N_577,N_448,N_481);
and U578 (N_578,N_417,N_444);
nor U579 (N_579,N_408,N_463);
xnor U580 (N_580,N_458,N_497);
nor U581 (N_581,N_463,N_478);
nand U582 (N_582,N_499,N_414);
nor U583 (N_583,N_431,N_441);
or U584 (N_584,N_419,N_492);
and U585 (N_585,N_481,N_424);
or U586 (N_586,N_451,N_456);
or U587 (N_587,N_425,N_413);
and U588 (N_588,N_415,N_403);
and U589 (N_589,N_401,N_452);
nor U590 (N_590,N_460,N_406);
or U591 (N_591,N_400,N_418);
nor U592 (N_592,N_492,N_463);
nor U593 (N_593,N_486,N_490);
nand U594 (N_594,N_483,N_430);
nand U595 (N_595,N_416,N_493);
nor U596 (N_596,N_403,N_451);
and U597 (N_597,N_470,N_498);
nand U598 (N_598,N_450,N_455);
and U599 (N_599,N_463,N_462);
xor U600 (N_600,N_540,N_511);
nor U601 (N_601,N_523,N_584);
and U602 (N_602,N_588,N_533);
and U603 (N_603,N_549,N_504);
or U604 (N_604,N_508,N_590);
or U605 (N_605,N_531,N_514);
and U606 (N_606,N_550,N_597);
or U607 (N_607,N_576,N_532);
nor U608 (N_608,N_548,N_541);
xnor U609 (N_609,N_587,N_507);
or U610 (N_610,N_552,N_566);
and U611 (N_611,N_595,N_559);
or U612 (N_612,N_562,N_589);
nor U613 (N_613,N_527,N_594);
and U614 (N_614,N_585,N_555);
nor U615 (N_615,N_554,N_505);
and U616 (N_616,N_557,N_503);
xor U617 (N_617,N_517,N_596);
and U618 (N_618,N_581,N_565);
nand U619 (N_619,N_520,N_564);
nand U620 (N_620,N_519,N_500);
nor U621 (N_621,N_545,N_510);
nand U622 (N_622,N_506,N_582);
or U623 (N_623,N_586,N_556);
and U624 (N_624,N_573,N_524);
nand U625 (N_625,N_522,N_512);
nand U626 (N_626,N_572,N_551);
or U627 (N_627,N_537,N_538);
or U628 (N_628,N_558,N_567);
and U629 (N_629,N_547,N_546);
and U630 (N_630,N_578,N_521);
nor U631 (N_631,N_529,N_561);
nor U632 (N_632,N_502,N_569);
and U633 (N_633,N_530,N_568);
or U634 (N_634,N_518,N_583);
or U635 (N_635,N_515,N_509);
and U636 (N_636,N_574,N_528);
and U637 (N_637,N_571,N_539);
nor U638 (N_638,N_591,N_575);
nor U639 (N_639,N_560,N_593);
nor U640 (N_640,N_501,N_577);
nand U641 (N_641,N_579,N_526);
or U642 (N_642,N_570,N_553);
nor U643 (N_643,N_516,N_535);
or U644 (N_644,N_563,N_536);
and U645 (N_645,N_542,N_513);
xnor U646 (N_646,N_580,N_598);
and U647 (N_647,N_599,N_592);
nand U648 (N_648,N_534,N_525);
nor U649 (N_649,N_543,N_544);
and U650 (N_650,N_597,N_507);
nand U651 (N_651,N_585,N_578);
nor U652 (N_652,N_579,N_580);
nor U653 (N_653,N_540,N_599);
or U654 (N_654,N_519,N_597);
nor U655 (N_655,N_521,N_564);
and U656 (N_656,N_508,N_583);
nor U657 (N_657,N_596,N_511);
or U658 (N_658,N_551,N_502);
and U659 (N_659,N_575,N_523);
and U660 (N_660,N_560,N_564);
nor U661 (N_661,N_570,N_587);
xor U662 (N_662,N_582,N_540);
xnor U663 (N_663,N_564,N_537);
and U664 (N_664,N_595,N_586);
and U665 (N_665,N_591,N_531);
or U666 (N_666,N_587,N_590);
nor U667 (N_667,N_599,N_552);
or U668 (N_668,N_502,N_572);
nor U669 (N_669,N_513,N_592);
or U670 (N_670,N_516,N_597);
and U671 (N_671,N_525,N_503);
and U672 (N_672,N_507,N_511);
or U673 (N_673,N_551,N_553);
and U674 (N_674,N_598,N_549);
or U675 (N_675,N_515,N_518);
and U676 (N_676,N_540,N_530);
nor U677 (N_677,N_563,N_520);
nor U678 (N_678,N_599,N_541);
nand U679 (N_679,N_599,N_570);
or U680 (N_680,N_578,N_556);
nand U681 (N_681,N_589,N_590);
nand U682 (N_682,N_576,N_594);
nand U683 (N_683,N_562,N_533);
or U684 (N_684,N_566,N_579);
nand U685 (N_685,N_554,N_555);
or U686 (N_686,N_566,N_530);
nand U687 (N_687,N_577,N_514);
or U688 (N_688,N_512,N_565);
or U689 (N_689,N_528,N_542);
nand U690 (N_690,N_527,N_534);
or U691 (N_691,N_543,N_567);
nand U692 (N_692,N_529,N_549);
or U693 (N_693,N_599,N_525);
nand U694 (N_694,N_555,N_518);
and U695 (N_695,N_510,N_517);
nor U696 (N_696,N_549,N_541);
xnor U697 (N_697,N_533,N_555);
and U698 (N_698,N_569,N_579);
and U699 (N_699,N_519,N_510);
or U700 (N_700,N_680,N_636);
nand U701 (N_701,N_621,N_661);
nor U702 (N_702,N_681,N_672);
xnor U703 (N_703,N_625,N_610);
nor U704 (N_704,N_626,N_637);
nand U705 (N_705,N_691,N_644);
or U706 (N_706,N_601,N_673);
nand U707 (N_707,N_614,N_646);
nand U708 (N_708,N_613,N_675);
nor U709 (N_709,N_645,N_632);
and U710 (N_710,N_652,N_663);
and U711 (N_711,N_648,N_690);
and U712 (N_712,N_699,N_677);
nand U713 (N_713,N_602,N_650);
nor U714 (N_714,N_694,N_612);
xor U715 (N_715,N_620,N_693);
and U716 (N_716,N_654,N_696);
or U717 (N_717,N_639,N_684);
nor U718 (N_718,N_617,N_624);
nand U719 (N_719,N_660,N_605);
nand U720 (N_720,N_678,N_679);
nand U721 (N_721,N_668,N_649);
and U722 (N_722,N_689,N_697);
or U723 (N_723,N_669,N_615);
nor U724 (N_724,N_657,N_695);
nor U725 (N_725,N_640,N_603);
or U726 (N_726,N_609,N_662);
and U727 (N_727,N_651,N_653);
or U728 (N_728,N_688,N_630);
nor U729 (N_729,N_667,N_698);
nor U730 (N_730,N_635,N_634);
nor U731 (N_731,N_611,N_642);
nand U732 (N_732,N_606,N_631);
nand U733 (N_733,N_608,N_607);
and U734 (N_734,N_685,N_616);
and U735 (N_735,N_666,N_658);
and U736 (N_736,N_627,N_676);
or U737 (N_737,N_618,N_665);
xnor U738 (N_738,N_687,N_623);
and U739 (N_739,N_692,N_643);
and U740 (N_740,N_671,N_674);
or U741 (N_741,N_628,N_638);
nand U742 (N_742,N_619,N_604);
nand U743 (N_743,N_683,N_655);
nand U744 (N_744,N_670,N_656);
xnor U745 (N_745,N_641,N_633);
nor U746 (N_746,N_682,N_686);
or U747 (N_747,N_629,N_659);
or U748 (N_748,N_664,N_600);
nor U749 (N_749,N_622,N_647);
and U750 (N_750,N_680,N_656);
or U751 (N_751,N_623,N_673);
or U752 (N_752,N_685,N_680);
or U753 (N_753,N_669,N_644);
nor U754 (N_754,N_618,N_697);
or U755 (N_755,N_603,N_682);
or U756 (N_756,N_653,N_604);
nor U757 (N_757,N_685,N_651);
nand U758 (N_758,N_680,N_678);
nand U759 (N_759,N_646,N_627);
and U760 (N_760,N_665,N_622);
nor U761 (N_761,N_624,N_686);
and U762 (N_762,N_655,N_628);
nand U763 (N_763,N_683,N_613);
nand U764 (N_764,N_686,N_617);
and U765 (N_765,N_635,N_676);
or U766 (N_766,N_638,N_699);
nor U767 (N_767,N_612,N_647);
or U768 (N_768,N_617,N_691);
xor U769 (N_769,N_627,N_631);
xnor U770 (N_770,N_605,N_673);
nand U771 (N_771,N_641,N_689);
nor U772 (N_772,N_647,N_645);
or U773 (N_773,N_612,N_686);
nor U774 (N_774,N_636,N_600);
or U775 (N_775,N_623,N_643);
xnor U776 (N_776,N_629,N_645);
xnor U777 (N_777,N_606,N_603);
or U778 (N_778,N_602,N_640);
nand U779 (N_779,N_631,N_695);
or U780 (N_780,N_622,N_624);
nor U781 (N_781,N_657,N_631);
nand U782 (N_782,N_629,N_600);
or U783 (N_783,N_616,N_643);
xnor U784 (N_784,N_677,N_653);
nand U785 (N_785,N_690,N_605);
or U786 (N_786,N_656,N_645);
nand U787 (N_787,N_679,N_656);
or U788 (N_788,N_665,N_608);
nor U789 (N_789,N_637,N_612);
xor U790 (N_790,N_638,N_624);
and U791 (N_791,N_651,N_640);
or U792 (N_792,N_669,N_631);
and U793 (N_793,N_666,N_677);
nor U794 (N_794,N_664,N_697);
nand U795 (N_795,N_608,N_678);
nand U796 (N_796,N_685,N_600);
and U797 (N_797,N_637,N_634);
nand U798 (N_798,N_683,N_698);
or U799 (N_799,N_680,N_643);
nand U800 (N_800,N_737,N_762);
nor U801 (N_801,N_756,N_703);
nor U802 (N_802,N_715,N_724);
nand U803 (N_803,N_729,N_789);
nand U804 (N_804,N_781,N_702);
xnor U805 (N_805,N_746,N_772);
nor U806 (N_806,N_782,N_766);
nand U807 (N_807,N_739,N_757);
xor U808 (N_808,N_767,N_710);
and U809 (N_809,N_707,N_753);
xor U810 (N_810,N_741,N_765);
nor U811 (N_811,N_764,N_768);
nor U812 (N_812,N_714,N_706);
nand U813 (N_813,N_731,N_754);
or U814 (N_814,N_773,N_790);
nand U815 (N_815,N_722,N_749);
nand U816 (N_816,N_745,N_717);
and U817 (N_817,N_760,N_777);
and U818 (N_818,N_733,N_784);
or U819 (N_819,N_711,N_793);
nor U820 (N_820,N_778,N_796);
nor U821 (N_821,N_743,N_770);
and U822 (N_822,N_709,N_740);
nor U823 (N_823,N_788,N_736);
nor U824 (N_824,N_771,N_774);
nand U825 (N_825,N_759,N_751);
or U826 (N_826,N_723,N_704);
nand U827 (N_827,N_748,N_783);
nand U828 (N_828,N_797,N_799);
nor U829 (N_829,N_727,N_728);
or U830 (N_830,N_730,N_763);
or U831 (N_831,N_791,N_752);
and U832 (N_832,N_734,N_755);
xnor U833 (N_833,N_735,N_761);
or U834 (N_834,N_794,N_776);
and U835 (N_835,N_795,N_726);
or U836 (N_836,N_747,N_738);
nand U837 (N_837,N_725,N_792);
or U838 (N_838,N_742,N_713);
or U839 (N_839,N_779,N_750);
xnor U840 (N_840,N_700,N_732);
or U841 (N_841,N_775,N_708);
and U842 (N_842,N_787,N_719);
nor U843 (N_843,N_798,N_769);
and U844 (N_844,N_780,N_716);
nand U845 (N_845,N_701,N_744);
or U846 (N_846,N_721,N_786);
and U847 (N_847,N_758,N_785);
and U848 (N_848,N_712,N_720);
nor U849 (N_849,N_705,N_718);
nand U850 (N_850,N_752,N_710);
and U851 (N_851,N_741,N_796);
nor U852 (N_852,N_761,N_764);
or U853 (N_853,N_712,N_789);
and U854 (N_854,N_754,N_752);
or U855 (N_855,N_720,N_750);
or U856 (N_856,N_712,N_773);
nand U857 (N_857,N_790,N_714);
and U858 (N_858,N_710,N_796);
nand U859 (N_859,N_702,N_734);
nor U860 (N_860,N_740,N_782);
and U861 (N_861,N_797,N_747);
nor U862 (N_862,N_784,N_701);
nor U863 (N_863,N_714,N_727);
xor U864 (N_864,N_722,N_723);
and U865 (N_865,N_727,N_739);
and U866 (N_866,N_739,N_787);
nor U867 (N_867,N_755,N_751);
nand U868 (N_868,N_751,N_770);
and U869 (N_869,N_795,N_701);
nor U870 (N_870,N_755,N_772);
and U871 (N_871,N_792,N_781);
nor U872 (N_872,N_700,N_783);
xor U873 (N_873,N_702,N_717);
xor U874 (N_874,N_766,N_772);
nand U875 (N_875,N_786,N_790);
nor U876 (N_876,N_787,N_770);
nor U877 (N_877,N_737,N_794);
or U878 (N_878,N_730,N_790);
and U879 (N_879,N_704,N_763);
nor U880 (N_880,N_740,N_717);
or U881 (N_881,N_752,N_781);
nand U882 (N_882,N_711,N_709);
nand U883 (N_883,N_779,N_771);
nand U884 (N_884,N_773,N_781);
nor U885 (N_885,N_766,N_776);
nor U886 (N_886,N_731,N_773);
or U887 (N_887,N_773,N_714);
or U888 (N_888,N_720,N_758);
nand U889 (N_889,N_764,N_720);
or U890 (N_890,N_716,N_738);
xor U891 (N_891,N_751,N_762);
nor U892 (N_892,N_764,N_734);
nor U893 (N_893,N_727,N_736);
nor U894 (N_894,N_734,N_729);
nand U895 (N_895,N_753,N_774);
nand U896 (N_896,N_717,N_714);
or U897 (N_897,N_700,N_760);
and U898 (N_898,N_728,N_731);
xor U899 (N_899,N_715,N_755);
and U900 (N_900,N_846,N_855);
nand U901 (N_901,N_889,N_804);
and U902 (N_902,N_813,N_847);
nand U903 (N_903,N_893,N_836);
nand U904 (N_904,N_874,N_803);
xor U905 (N_905,N_818,N_867);
nor U906 (N_906,N_890,N_887);
and U907 (N_907,N_831,N_827);
nor U908 (N_908,N_863,N_800);
and U909 (N_909,N_856,N_861);
nor U910 (N_910,N_883,N_850);
or U911 (N_911,N_802,N_848);
and U912 (N_912,N_885,N_898);
nand U913 (N_913,N_860,N_859);
nand U914 (N_914,N_875,N_814);
and U915 (N_915,N_842,N_844);
and U916 (N_916,N_837,N_816);
and U917 (N_917,N_891,N_880);
or U918 (N_918,N_871,N_857);
nor U919 (N_919,N_862,N_817);
and U920 (N_920,N_878,N_808);
nand U921 (N_921,N_858,N_822);
and U922 (N_922,N_834,N_841);
nand U923 (N_923,N_852,N_838);
nor U924 (N_924,N_812,N_892);
or U925 (N_925,N_882,N_868);
nand U926 (N_926,N_870,N_879);
nand U927 (N_927,N_886,N_897);
nand U928 (N_928,N_821,N_843);
or U929 (N_929,N_811,N_884);
or U930 (N_930,N_853,N_833);
nand U931 (N_931,N_888,N_801);
or U932 (N_932,N_806,N_826);
and U933 (N_933,N_873,N_820);
or U934 (N_934,N_830,N_832);
nand U935 (N_935,N_849,N_807);
or U936 (N_936,N_896,N_809);
or U937 (N_937,N_845,N_851);
nand U938 (N_938,N_824,N_819);
and U939 (N_939,N_839,N_835);
or U940 (N_940,N_881,N_866);
nand U941 (N_941,N_840,N_895);
and U942 (N_942,N_876,N_823);
or U943 (N_943,N_872,N_899);
nand U944 (N_944,N_854,N_825);
or U945 (N_945,N_894,N_815);
nor U946 (N_946,N_869,N_805);
nand U947 (N_947,N_810,N_865);
nand U948 (N_948,N_877,N_828);
nand U949 (N_949,N_864,N_829);
and U950 (N_950,N_871,N_840);
nor U951 (N_951,N_803,N_826);
or U952 (N_952,N_860,N_814);
or U953 (N_953,N_832,N_838);
or U954 (N_954,N_896,N_849);
and U955 (N_955,N_816,N_884);
nand U956 (N_956,N_867,N_875);
or U957 (N_957,N_837,N_854);
and U958 (N_958,N_889,N_827);
nand U959 (N_959,N_812,N_817);
and U960 (N_960,N_829,N_854);
and U961 (N_961,N_803,N_837);
nor U962 (N_962,N_865,N_895);
or U963 (N_963,N_889,N_819);
nand U964 (N_964,N_882,N_856);
nand U965 (N_965,N_895,N_861);
xor U966 (N_966,N_876,N_806);
or U967 (N_967,N_882,N_822);
and U968 (N_968,N_847,N_859);
nor U969 (N_969,N_870,N_876);
and U970 (N_970,N_891,N_857);
nand U971 (N_971,N_885,N_803);
and U972 (N_972,N_862,N_826);
or U973 (N_973,N_833,N_866);
nor U974 (N_974,N_825,N_850);
or U975 (N_975,N_803,N_836);
and U976 (N_976,N_859,N_868);
nand U977 (N_977,N_891,N_809);
and U978 (N_978,N_871,N_898);
and U979 (N_979,N_889,N_801);
and U980 (N_980,N_889,N_814);
or U981 (N_981,N_858,N_839);
or U982 (N_982,N_819,N_860);
and U983 (N_983,N_823,N_873);
nand U984 (N_984,N_851,N_869);
and U985 (N_985,N_848,N_813);
nand U986 (N_986,N_815,N_838);
nand U987 (N_987,N_833,N_837);
or U988 (N_988,N_857,N_845);
nor U989 (N_989,N_891,N_846);
or U990 (N_990,N_868,N_840);
nand U991 (N_991,N_883,N_869);
nor U992 (N_992,N_801,N_831);
or U993 (N_993,N_894,N_829);
or U994 (N_994,N_889,N_893);
nand U995 (N_995,N_884,N_812);
nor U996 (N_996,N_838,N_892);
nand U997 (N_997,N_815,N_830);
nor U998 (N_998,N_849,N_872);
nand U999 (N_999,N_812,N_865);
nor U1000 (N_1000,N_922,N_967);
or U1001 (N_1001,N_935,N_960);
and U1002 (N_1002,N_947,N_995);
or U1003 (N_1003,N_912,N_963);
nand U1004 (N_1004,N_980,N_918);
nor U1005 (N_1005,N_934,N_905);
or U1006 (N_1006,N_965,N_983);
nand U1007 (N_1007,N_933,N_902);
nand U1008 (N_1008,N_944,N_999);
nand U1009 (N_1009,N_919,N_997);
nor U1010 (N_1010,N_906,N_911);
nand U1011 (N_1011,N_953,N_928);
or U1012 (N_1012,N_923,N_982);
and U1013 (N_1013,N_937,N_961);
nand U1014 (N_1014,N_998,N_917);
and U1015 (N_1015,N_925,N_931);
and U1016 (N_1016,N_926,N_952);
or U1017 (N_1017,N_978,N_959);
nor U1018 (N_1018,N_991,N_968);
and U1019 (N_1019,N_913,N_969);
nand U1020 (N_1020,N_941,N_977);
and U1021 (N_1021,N_920,N_939);
nand U1022 (N_1022,N_908,N_985);
or U1023 (N_1023,N_994,N_981);
and U1024 (N_1024,N_976,N_924);
or U1025 (N_1025,N_972,N_930);
nor U1026 (N_1026,N_943,N_990);
and U1027 (N_1027,N_903,N_979);
or U1028 (N_1028,N_916,N_958);
nor U1029 (N_1029,N_927,N_956);
nor U1030 (N_1030,N_989,N_907);
nor U1031 (N_1031,N_954,N_915);
nand U1032 (N_1032,N_932,N_945);
nand U1033 (N_1033,N_955,N_940);
nor U1034 (N_1034,N_929,N_986);
xor U1035 (N_1035,N_942,N_938);
nor U1036 (N_1036,N_975,N_910);
and U1037 (N_1037,N_984,N_946);
and U1038 (N_1038,N_909,N_950);
or U1039 (N_1039,N_949,N_900);
nand U1040 (N_1040,N_974,N_904);
and U1041 (N_1041,N_948,N_971);
nor U1042 (N_1042,N_966,N_957);
xor U1043 (N_1043,N_962,N_936);
nor U1044 (N_1044,N_993,N_992);
and U1045 (N_1045,N_988,N_901);
nor U1046 (N_1046,N_921,N_973);
and U1047 (N_1047,N_951,N_970);
or U1048 (N_1048,N_996,N_964);
nand U1049 (N_1049,N_914,N_987);
or U1050 (N_1050,N_904,N_999);
or U1051 (N_1051,N_942,N_967);
xnor U1052 (N_1052,N_929,N_974);
nand U1053 (N_1053,N_924,N_919);
or U1054 (N_1054,N_964,N_905);
and U1055 (N_1055,N_901,N_944);
nor U1056 (N_1056,N_969,N_989);
nor U1057 (N_1057,N_919,N_977);
nor U1058 (N_1058,N_993,N_985);
and U1059 (N_1059,N_961,N_990);
nand U1060 (N_1060,N_966,N_949);
nand U1061 (N_1061,N_951,N_988);
nor U1062 (N_1062,N_931,N_944);
nor U1063 (N_1063,N_943,N_931);
nor U1064 (N_1064,N_955,N_904);
nand U1065 (N_1065,N_923,N_910);
or U1066 (N_1066,N_945,N_915);
nand U1067 (N_1067,N_982,N_985);
nor U1068 (N_1068,N_933,N_917);
nor U1069 (N_1069,N_996,N_972);
nor U1070 (N_1070,N_939,N_917);
and U1071 (N_1071,N_902,N_999);
nor U1072 (N_1072,N_937,N_989);
or U1073 (N_1073,N_917,N_910);
nand U1074 (N_1074,N_965,N_985);
and U1075 (N_1075,N_915,N_909);
nand U1076 (N_1076,N_928,N_996);
and U1077 (N_1077,N_986,N_956);
or U1078 (N_1078,N_971,N_913);
nor U1079 (N_1079,N_968,N_902);
or U1080 (N_1080,N_942,N_934);
xnor U1081 (N_1081,N_921,N_992);
and U1082 (N_1082,N_938,N_947);
nor U1083 (N_1083,N_942,N_939);
or U1084 (N_1084,N_957,N_986);
nor U1085 (N_1085,N_922,N_973);
and U1086 (N_1086,N_961,N_940);
or U1087 (N_1087,N_959,N_980);
nor U1088 (N_1088,N_994,N_939);
and U1089 (N_1089,N_963,N_961);
and U1090 (N_1090,N_938,N_945);
nor U1091 (N_1091,N_934,N_965);
and U1092 (N_1092,N_926,N_998);
or U1093 (N_1093,N_926,N_957);
and U1094 (N_1094,N_952,N_965);
or U1095 (N_1095,N_941,N_994);
nor U1096 (N_1096,N_977,N_932);
or U1097 (N_1097,N_933,N_984);
nor U1098 (N_1098,N_907,N_932);
and U1099 (N_1099,N_919,N_963);
or U1100 (N_1100,N_1092,N_1012);
nand U1101 (N_1101,N_1095,N_1048);
nor U1102 (N_1102,N_1099,N_1054);
nor U1103 (N_1103,N_1075,N_1055);
and U1104 (N_1104,N_1064,N_1000);
nor U1105 (N_1105,N_1019,N_1010);
nand U1106 (N_1106,N_1018,N_1032);
and U1107 (N_1107,N_1034,N_1052);
and U1108 (N_1108,N_1029,N_1090);
or U1109 (N_1109,N_1063,N_1069);
nor U1110 (N_1110,N_1085,N_1071);
nand U1111 (N_1111,N_1066,N_1093);
or U1112 (N_1112,N_1074,N_1073);
and U1113 (N_1113,N_1087,N_1047);
nor U1114 (N_1114,N_1098,N_1081);
nand U1115 (N_1115,N_1036,N_1078);
nor U1116 (N_1116,N_1091,N_1037);
or U1117 (N_1117,N_1053,N_1041);
or U1118 (N_1118,N_1077,N_1027);
and U1119 (N_1119,N_1050,N_1079);
or U1120 (N_1120,N_1006,N_1039);
nor U1121 (N_1121,N_1057,N_1016);
and U1122 (N_1122,N_1045,N_1030);
or U1123 (N_1123,N_1083,N_1094);
or U1124 (N_1124,N_1026,N_1065);
and U1125 (N_1125,N_1068,N_1003);
and U1126 (N_1126,N_1040,N_1033);
or U1127 (N_1127,N_1096,N_1009);
and U1128 (N_1128,N_1042,N_1014);
nand U1129 (N_1129,N_1004,N_1049);
and U1130 (N_1130,N_1017,N_1025);
nor U1131 (N_1131,N_1015,N_1021);
nor U1132 (N_1132,N_1005,N_1028);
and U1133 (N_1133,N_1061,N_1011);
and U1134 (N_1134,N_1088,N_1082);
nor U1135 (N_1135,N_1001,N_1062);
or U1136 (N_1136,N_1084,N_1024);
nor U1137 (N_1137,N_1072,N_1097);
or U1138 (N_1138,N_1031,N_1023);
or U1139 (N_1139,N_1046,N_1059);
or U1140 (N_1140,N_1020,N_1058);
nand U1141 (N_1141,N_1008,N_1022);
and U1142 (N_1142,N_1007,N_1043);
nor U1143 (N_1143,N_1060,N_1002);
or U1144 (N_1144,N_1070,N_1035);
and U1145 (N_1145,N_1044,N_1089);
or U1146 (N_1146,N_1080,N_1013);
xor U1147 (N_1147,N_1038,N_1056);
nand U1148 (N_1148,N_1067,N_1051);
and U1149 (N_1149,N_1086,N_1076);
nor U1150 (N_1150,N_1037,N_1047);
nand U1151 (N_1151,N_1010,N_1055);
and U1152 (N_1152,N_1034,N_1009);
and U1153 (N_1153,N_1062,N_1003);
nand U1154 (N_1154,N_1016,N_1051);
nand U1155 (N_1155,N_1016,N_1084);
and U1156 (N_1156,N_1094,N_1036);
nor U1157 (N_1157,N_1067,N_1040);
or U1158 (N_1158,N_1020,N_1041);
or U1159 (N_1159,N_1066,N_1041);
and U1160 (N_1160,N_1023,N_1017);
nor U1161 (N_1161,N_1037,N_1076);
nand U1162 (N_1162,N_1057,N_1015);
or U1163 (N_1163,N_1071,N_1033);
or U1164 (N_1164,N_1071,N_1095);
and U1165 (N_1165,N_1058,N_1064);
nand U1166 (N_1166,N_1043,N_1046);
nand U1167 (N_1167,N_1038,N_1086);
nand U1168 (N_1168,N_1094,N_1058);
nand U1169 (N_1169,N_1083,N_1037);
or U1170 (N_1170,N_1073,N_1053);
or U1171 (N_1171,N_1035,N_1062);
nand U1172 (N_1172,N_1078,N_1025);
nand U1173 (N_1173,N_1048,N_1031);
or U1174 (N_1174,N_1094,N_1066);
nor U1175 (N_1175,N_1085,N_1067);
and U1176 (N_1176,N_1012,N_1082);
or U1177 (N_1177,N_1057,N_1068);
and U1178 (N_1178,N_1090,N_1003);
and U1179 (N_1179,N_1016,N_1011);
nand U1180 (N_1180,N_1006,N_1072);
and U1181 (N_1181,N_1021,N_1058);
nand U1182 (N_1182,N_1085,N_1042);
or U1183 (N_1183,N_1014,N_1045);
and U1184 (N_1184,N_1080,N_1041);
nor U1185 (N_1185,N_1088,N_1026);
or U1186 (N_1186,N_1077,N_1063);
or U1187 (N_1187,N_1011,N_1069);
or U1188 (N_1188,N_1065,N_1006);
or U1189 (N_1189,N_1079,N_1083);
or U1190 (N_1190,N_1000,N_1061);
nor U1191 (N_1191,N_1057,N_1095);
or U1192 (N_1192,N_1006,N_1024);
nand U1193 (N_1193,N_1072,N_1068);
and U1194 (N_1194,N_1007,N_1091);
and U1195 (N_1195,N_1016,N_1074);
nand U1196 (N_1196,N_1059,N_1052);
and U1197 (N_1197,N_1053,N_1039);
nor U1198 (N_1198,N_1054,N_1020);
and U1199 (N_1199,N_1018,N_1033);
nand U1200 (N_1200,N_1106,N_1195);
and U1201 (N_1201,N_1168,N_1196);
and U1202 (N_1202,N_1143,N_1148);
and U1203 (N_1203,N_1188,N_1198);
nor U1204 (N_1204,N_1119,N_1181);
and U1205 (N_1205,N_1115,N_1103);
and U1206 (N_1206,N_1153,N_1158);
nand U1207 (N_1207,N_1173,N_1156);
nand U1208 (N_1208,N_1101,N_1199);
xnor U1209 (N_1209,N_1192,N_1138);
nand U1210 (N_1210,N_1147,N_1129);
and U1211 (N_1211,N_1141,N_1110);
and U1212 (N_1212,N_1175,N_1191);
and U1213 (N_1213,N_1111,N_1176);
or U1214 (N_1214,N_1179,N_1165);
and U1215 (N_1215,N_1128,N_1127);
and U1216 (N_1216,N_1124,N_1146);
nand U1217 (N_1217,N_1154,N_1135);
nor U1218 (N_1218,N_1162,N_1190);
xor U1219 (N_1219,N_1140,N_1169);
nand U1220 (N_1220,N_1150,N_1117);
nand U1221 (N_1221,N_1197,N_1108);
nand U1222 (N_1222,N_1113,N_1121);
or U1223 (N_1223,N_1112,N_1102);
nor U1224 (N_1224,N_1180,N_1167);
or U1225 (N_1225,N_1160,N_1159);
or U1226 (N_1226,N_1155,N_1163);
or U1227 (N_1227,N_1157,N_1130);
or U1228 (N_1228,N_1100,N_1122);
nand U1229 (N_1229,N_1125,N_1109);
nand U1230 (N_1230,N_1136,N_1174);
or U1231 (N_1231,N_1151,N_1123);
nand U1232 (N_1232,N_1126,N_1114);
nor U1233 (N_1233,N_1161,N_1120);
or U1234 (N_1234,N_1104,N_1116);
nand U1235 (N_1235,N_1132,N_1134);
nand U1236 (N_1236,N_1145,N_1139);
nand U1237 (N_1237,N_1166,N_1170);
and U1238 (N_1238,N_1186,N_1187);
or U1239 (N_1239,N_1189,N_1164);
or U1240 (N_1240,N_1142,N_1177);
nand U1241 (N_1241,N_1137,N_1182);
and U1242 (N_1242,N_1152,N_1193);
nand U1243 (N_1243,N_1118,N_1171);
and U1244 (N_1244,N_1105,N_1183);
nor U1245 (N_1245,N_1178,N_1185);
and U1246 (N_1246,N_1184,N_1133);
or U1247 (N_1247,N_1107,N_1131);
nand U1248 (N_1248,N_1149,N_1172);
and U1249 (N_1249,N_1194,N_1144);
nand U1250 (N_1250,N_1120,N_1105);
and U1251 (N_1251,N_1197,N_1109);
nor U1252 (N_1252,N_1113,N_1175);
or U1253 (N_1253,N_1185,N_1125);
or U1254 (N_1254,N_1110,N_1147);
nand U1255 (N_1255,N_1159,N_1136);
and U1256 (N_1256,N_1181,N_1137);
nand U1257 (N_1257,N_1187,N_1169);
and U1258 (N_1258,N_1176,N_1157);
nand U1259 (N_1259,N_1176,N_1159);
nand U1260 (N_1260,N_1171,N_1106);
or U1261 (N_1261,N_1107,N_1157);
nand U1262 (N_1262,N_1118,N_1110);
xnor U1263 (N_1263,N_1115,N_1109);
nor U1264 (N_1264,N_1157,N_1127);
nand U1265 (N_1265,N_1150,N_1125);
nor U1266 (N_1266,N_1122,N_1169);
and U1267 (N_1267,N_1168,N_1107);
or U1268 (N_1268,N_1108,N_1184);
nor U1269 (N_1269,N_1198,N_1116);
xor U1270 (N_1270,N_1169,N_1104);
nor U1271 (N_1271,N_1195,N_1103);
or U1272 (N_1272,N_1182,N_1144);
xnor U1273 (N_1273,N_1114,N_1180);
nand U1274 (N_1274,N_1123,N_1121);
nand U1275 (N_1275,N_1140,N_1133);
and U1276 (N_1276,N_1174,N_1121);
nand U1277 (N_1277,N_1191,N_1181);
xnor U1278 (N_1278,N_1161,N_1191);
and U1279 (N_1279,N_1162,N_1191);
nand U1280 (N_1280,N_1187,N_1125);
and U1281 (N_1281,N_1194,N_1175);
or U1282 (N_1282,N_1123,N_1147);
nor U1283 (N_1283,N_1179,N_1122);
nor U1284 (N_1284,N_1148,N_1172);
xor U1285 (N_1285,N_1156,N_1105);
and U1286 (N_1286,N_1165,N_1196);
nand U1287 (N_1287,N_1191,N_1148);
or U1288 (N_1288,N_1175,N_1171);
nor U1289 (N_1289,N_1151,N_1191);
and U1290 (N_1290,N_1172,N_1133);
xor U1291 (N_1291,N_1169,N_1108);
and U1292 (N_1292,N_1145,N_1133);
and U1293 (N_1293,N_1191,N_1159);
and U1294 (N_1294,N_1142,N_1179);
or U1295 (N_1295,N_1130,N_1144);
or U1296 (N_1296,N_1150,N_1172);
and U1297 (N_1297,N_1119,N_1110);
or U1298 (N_1298,N_1140,N_1121);
nand U1299 (N_1299,N_1103,N_1184);
and U1300 (N_1300,N_1230,N_1218);
nand U1301 (N_1301,N_1250,N_1211);
nor U1302 (N_1302,N_1231,N_1276);
or U1303 (N_1303,N_1245,N_1253);
and U1304 (N_1304,N_1240,N_1252);
nand U1305 (N_1305,N_1202,N_1235);
or U1306 (N_1306,N_1279,N_1283);
and U1307 (N_1307,N_1299,N_1241);
or U1308 (N_1308,N_1296,N_1206);
nor U1309 (N_1309,N_1272,N_1200);
and U1310 (N_1310,N_1285,N_1207);
nor U1311 (N_1311,N_1239,N_1219);
nand U1312 (N_1312,N_1214,N_1268);
or U1313 (N_1313,N_1247,N_1261);
nand U1314 (N_1314,N_1216,N_1273);
or U1315 (N_1315,N_1234,N_1286);
or U1316 (N_1316,N_1204,N_1233);
xor U1317 (N_1317,N_1269,N_1280);
and U1318 (N_1318,N_1228,N_1229);
and U1319 (N_1319,N_1238,N_1221);
xor U1320 (N_1320,N_1242,N_1267);
nand U1321 (N_1321,N_1264,N_1265);
or U1322 (N_1322,N_1232,N_1260);
nor U1323 (N_1323,N_1222,N_1224);
xor U1324 (N_1324,N_1237,N_1278);
and U1325 (N_1325,N_1289,N_1256);
or U1326 (N_1326,N_1215,N_1227);
and U1327 (N_1327,N_1275,N_1293);
nand U1328 (N_1328,N_1294,N_1292);
nand U1329 (N_1329,N_1258,N_1217);
nor U1330 (N_1330,N_1208,N_1277);
and U1331 (N_1331,N_1259,N_1281);
or U1332 (N_1332,N_1271,N_1295);
or U1333 (N_1333,N_1251,N_1270);
nor U1334 (N_1334,N_1212,N_1255);
xor U1335 (N_1335,N_1201,N_1284);
nor U1336 (N_1336,N_1288,N_1210);
nor U1337 (N_1337,N_1274,N_1249);
nand U1338 (N_1338,N_1225,N_1297);
or U1339 (N_1339,N_1220,N_1243);
nand U1340 (N_1340,N_1257,N_1246);
nor U1341 (N_1341,N_1244,N_1205);
nand U1342 (N_1342,N_1262,N_1203);
nor U1343 (N_1343,N_1236,N_1254);
nand U1344 (N_1344,N_1287,N_1226);
and U1345 (N_1345,N_1213,N_1223);
or U1346 (N_1346,N_1209,N_1248);
nand U1347 (N_1347,N_1266,N_1263);
nand U1348 (N_1348,N_1282,N_1298);
nor U1349 (N_1349,N_1290,N_1291);
nand U1350 (N_1350,N_1261,N_1276);
and U1351 (N_1351,N_1209,N_1273);
nand U1352 (N_1352,N_1259,N_1289);
xor U1353 (N_1353,N_1216,N_1257);
nor U1354 (N_1354,N_1278,N_1209);
nand U1355 (N_1355,N_1246,N_1295);
nand U1356 (N_1356,N_1272,N_1298);
and U1357 (N_1357,N_1277,N_1273);
nand U1358 (N_1358,N_1266,N_1210);
or U1359 (N_1359,N_1206,N_1295);
nor U1360 (N_1360,N_1234,N_1262);
or U1361 (N_1361,N_1269,N_1279);
or U1362 (N_1362,N_1237,N_1220);
nand U1363 (N_1363,N_1232,N_1296);
nor U1364 (N_1364,N_1208,N_1256);
and U1365 (N_1365,N_1246,N_1217);
or U1366 (N_1366,N_1235,N_1288);
or U1367 (N_1367,N_1211,N_1221);
and U1368 (N_1368,N_1263,N_1233);
nor U1369 (N_1369,N_1259,N_1260);
nand U1370 (N_1370,N_1284,N_1274);
or U1371 (N_1371,N_1200,N_1297);
and U1372 (N_1372,N_1226,N_1297);
nor U1373 (N_1373,N_1245,N_1252);
or U1374 (N_1374,N_1241,N_1248);
or U1375 (N_1375,N_1240,N_1254);
xnor U1376 (N_1376,N_1268,N_1215);
and U1377 (N_1377,N_1273,N_1283);
nor U1378 (N_1378,N_1244,N_1295);
nor U1379 (N_1379,N_1212,N_1209);
or U1380 (N_1380,N_1265,N_1236);
nor U1381 (N_1381,N_1270,N_1290);
or U1382 (N_1382,N_1203,N_1296);
or U1383 (N_1383,N_1202,N_1264);
nor U1384 (N_1384,N_1212,N_1210);
or U1385 (N_1385,N_1228,N_1281);
nand U1386 (N_1386,N_1225,N_1222);
or U1387 (N_1387,N_1205,N_1206);
nor U1388 (N_1388,N_1224,N_1239);
nor U1389 (N_1389,N_1264,N_1269);
and U1390 (N_1390,N_1269,N_1212);
and U1391 (N_1391,N_1278,N_1262);
or U1392 (N_1392,N_1269,N_1260);
or U1393 (N_1393,N_1272,N_1281);
and U1394 (N_1394,N_1282,N_1202);
or U1395 (N_1395,N_1269,N_1281);
nand U1396 (N_1396,N_1213,N_1233);
nor U1397 (N_1397,N_1220,N_1251);
nand U1398 (N_1398,N_1265,N_1203);
nand U1399 (N_1399,N_1288,N_1286);
and U1400 (N_1400,N_1300,N_1372);
nor U1401 (N_1401,N_1312,N_1333);
nand U1402 (N_1402,N_1383,N_1341);
or U1403 (N_1403,N_1330,N_1399);
and U1404 (N_1404,N_1386,N_1348);
or U1405 (N_1405,N_1322,N_1391);
nor U1406 (N_1406,N_1344,N_1393);
nor U1407 (N_1407,N_1352,N_1357);
nor U1408 (N_1408,N_1310,N_1343);
or U1409 (N_1409,N_1331,N_1354);
nor U1410 (N_1410,N_1321,N_1345);
and U1411 (N_1411,N_1377,N_1389);
nand U1412 (N_1412,N_1374,N_1395);
and U1413 (N_1413,N_1396,N_1359);
and U1414 (N_1414,N_1304,N_1375);
and U1415 (N_1415,N_1368,N_1365);
and U1416 (N_1416,N_1337,N_1379);
or U1417 (N_1417,N_1319,N_1392);
and U1418 (N_1418,N_1371,N_1384);
and U1419 (N_1419,N_1323,N_1380);
and U1420 (N_1420,N_1335,N_1353);
or U1421 (N_1421,N_1361,N_1303);
and U1422 (N_1422,N_1315,N_1308);
nand U1423 (N_1423,N_1306,N_1324);
nor U1424 (N_1424,N_1326,N_1356);
nand U1425 (N_1425,N_1362,N_1364);
or U1426 (N_1426,N_1369,N_1340);
nand U1427 (N_1427,N_1376,N_1328);
and U1428 (N_1428,N_1370,N_1334);
and U1429 (N_1429,N_1302,N_1390);
nand U1430 (N_1430,N_1349,N_1373);
or U1431 (N_1431,N_1301,N_1381);
nor U1432 (N_1432,N_1305,N_1336);
or U1433 (N_1433,N_1320,N_1325);
or U1434 (N_1434,N_1355,N_1338);
or U1435 (N_1435,N_1332,N_1318);
and U1436 (N_1436,N_1347,N_1385);
nand U1437 (N_1437,N_1314,N_1397);
and U1438 (N_1438,N_1339,N_1387);
and U1439 (N_1439,N_1398,N_1311);
nor U1440 (N_1440,N_1316,N_1388);
and U1441 (N_1441,N_1329,N_1327);
nand U1442 (N_1442,N_1313,N_1346);
and U1443 (N_1443,N_1309,N_1350);
nor U1444 (N_1444,N_1342,N_1378);
or U1445 (N_1445,N_1382,N_1394);
or U1446 (N_1446,N_1366,N_1358);
and U1447 (N_1447,N_1360,N_1317);
nor U1448 (N_1448,N_1307,N_1363);
nor U1449 (N_1449,N_1351,N_1367);
and U1450 (N_1450,N_1367,N_1363);
nor U1451 (N_1451,N_1316,N_1325);
and U1452 (N_1452,N_1387,N_1332);
or U1453 (N_1453,N_1320,N_1330);
nand U1454 (N_1454,N_1316,N_1301);
or U1455 (N_1455,N_1306,N_1373);
nor U1456 (N_1456,N_1337,N_1303);
and U1457 (N_1457,N_1387,N_1321);
nand U1458 (N_1458,N_1321,N_1384);
and U1459 (N_1459,N_1337,N_1376);
or U1460 (N_1460,N_1386,N_1335);
nand U1461 (N_1461,N_1344,N_1305);
or U1462 (N_1462,N_1321,N_1308);
nand U1463 (N_1463,N_1356,N_1392);
nand U1464 (N_1464,N_1390,N_1369);
nor U1465 (N_1465,N_1325,N_1314);
nor U1466 (N_1466,N_1311,N_1371);
and U1467 (N_1467,N_1325,N_1312);
or U1468 (N_1468,N_1327,N_1335);
and U1469 (N_1469,N_1337,N_1314);
or U1470 (N_1470,N_1339,N_1332);
nor U1471 (N_1471,N_1380,N_1310);
or U1472 (N_1472,N_1379,N_1354);
or U1473 (N_1473,N_1313,N_1369);
nor U1474 (N_1474,N_1346,N_1388);
nor U1475 (N_1475,N_1378,N_1318);
or U1476 (N_1476,N_1341,N_1364);
nor U1477 (N_1477,N_1380,N_1361);
or U1478 (N_1478,N_1319,N_1339);
and U1479 (N_1479,N_1372,N_1349);
or U1480 (N_1480,N_1337,N_1347);
nor U1481 (N_1481,N_1324,N_1309);
and U1482 (N_1482,N_1379,N_1342);
nor U1483 (N_1483,N_1369,N_1333);
and U1484 (N_1484,N_1346,N_1368);
nor U1485 (N_1485,N_1358,N_1302);
xor U1486 (N_1486,N_1322,N_1346);
and U1487 (N_1487,N_1358,N_1342);
or U1488 (N_1488,N_1377,N_1386);
and U1489 (N_1489,N_1344,N_1330);
nor U1490 (N_1490,N_1392,N_1381);
nor U1491 (N_1491,N_1349,N_1391);
nor U1492 (N_1492,N_1368,N_1366);
nor U1493 (N_1493,N_1348,N_1320);
nand U1494 (N_1494,N_1310,N_1324);
or U1495 (N_1495,N_1330,N_1385);
and U1496 (N_1496,N_1389,N_1329);
nor U1497 (N_1497,N_1364,N_1365);
and U1498 (N_1498,N_1312,N_1358);
nand U1499 (N_1499,N_1365,N_1375);
nand U1500 (N_1500,N_1465,N_1451);
nand U1501 (N_1501,N_1446,N_1440);
nand U1502 (N_1502,N_1493,N_1434);
nand U1503 (N_1503,N_1484,N_1403);
or U1504 (N_1504,N_1453,N_1481);
nand U1505 (N_1505,N_1496,N_1487);
or U1506 (N_1506,N_1477,N_1448);
or U1507 (N_1507,N_1490,N_1409);
and U1508 (N_1508,N_1483,N_1498);
xor U1509 (N_1509,N_1444,N_1435);
nand U1510 (N_1510,N_1429,N_1458);
or U1511 (N_1511,N_1442,N_1402);
or U1512 (N_1512,N_1460,N_1405);
nand U1513 (N_1513,N_1426,N_1425);
nand U1514 (N_1514,N_1478,N_1464);
nor U1515 (N_1515,N_1412,N_1470);
nand U1516 (N_1516,N_1488,N_1447);
nor U1517 (N_1517,N_1480,N_1420);
and U1518 (N_1518,N_1492,N_1400);
nor U1519 (N_1519,N_1443,N_1404);
or U1520 (N_1520,N_1457,N_1479);
xnor U1521 (N_1521,N_1494,N_1455);
nor U1522 (N_1522,N_1449,N_1406);
nor U1523 (N_1523,N_1469,N_1411);
nand U1524 (N_1524,N_1463,N_1410);
nand U1525 (N_1525,N_1495,N_1486);
nand U1526 (N_1526,N_1430,N_1456);
and U1527 (N_1527,N_1454,N_1472);
nand U1528 (N_1528,N_1473,N_1467);
nand U1529 (N_1529,N_1474,N_1418);
xnor U1530 (N_1530,N_1427,N_1415);
xnor U1531 (N_1531,N_1401,N_1441);
nand U1532 (N_1532,N_1482,N_1445);
nor U1533 (N_1533,N_1437,N_1439);
nor U1534 (N_1534,N_1428,N_1423);
or U1535 (N_1535,N_1424,N_1462);
nand U1536 (N_1536,N_1452,N_1475);
and U1537 (N_1537,N_1421,N_1497);
nand U1538 (N_1538,N_1407,N_1459);
or U1539 (N_1539,N_1468,N_1413);
nor U1540 (N_1540,N_1466,N_1489);
nand U1541 (N_1541,N_1476,N_1485);
or U1542 (N_1542,N_1432,N_1408);
or U1543 (N_1543,N_1416,N_1414);
nor U1544 (N_1544,N_1491,N_1461);
nor U1545 (N_1545,N_1471,N_1419);
nor U1546 (N_1546,N_1499,N_1417);
nand U1547 (N_1547,N_1431,N_1450);
nor U1548 (N_1548,N_1438,N_1433);
and U1549 (N_1549,N_1422,N_1436);
nor U1550 (N_1550,N_1443,N_1478);
nor U1551 (N_1551,N_1452,N_1411);
nand U1552 (N_1552,N_1458,N_1423);
xnor U1553 (N_1553,N_1445,N_1497);
nor U1554 (N_1554,N_1433,N_1497);
or U1555 (N_1555,N_1414,N_1466);
and U1556 (N_1556,N_1431,N_1417);
nand U1557 (N_1557,N_1472,N_1462);
nand U1558 (N_1558,N_1468,N_1466);
nor U1559 (N_1559,N_1487,N_1472);
nand U1560 (N_1560,N_1455,N_1490);
and U1561 (N_1561,N_1495,N_1425);
nor U1562 (N_1562,N_1416,N_1415);
nand U1563 (N_1563,N_1452,N_1457);
nor U1564 (N_1564,N_1444,N_1460);
nand U1565 (N_1565,N_1452,N_1454);
xnor U1566 (N_1566,N_1492,N_1472);
or U1567 (N_1567,N_1479,N_1464);
xor U1568 (N_1568,N_1434,N_1407);
nor U1569 (N_1569,N_1456,N_1490);
and U1570 (N_1570,N_1438,N_1430);
nor U1571 (N_1571,N_1430,N_1478);
xnor U1572 (N_1572,N_1409,N_1445);
nand U1573 (N_1573,N_1405,N_1451);
nand U1574 (N_1574,N_1446,N_1409);
and U1575 (N_1575,N_1488,N_1408);
and U1576 (N_1576,N_1443,N_1416);
or U1577 (N_1577,N_1461,N_1467);
or U1578 (N_1578,N_1417,N_1440);
and U1579 (N_1579,N_1425,N_1412);
nor U1580 (N_1580,N_1444,N_1432);
nor U1581 (N_1581,N_1411,N_1423);
nor U1582 (N_1582,N_1422,N_1493);
or U1583 (N_1583,N_1420,N_1458);
nor U1584 (N_1584,N_1449,N_1466);
nor U1585 (N_1585,N_1401,N_1439);
and U1586 (N_1586,N_1418,N_1425);
nor U1587 (N_1587,N_1457,N_1480);
nand U1588 (N_1588,N_1451,N_1464);
nor U1589 (N_1589,N_1421,N_1456);
nor U1590 (N_1590,N_1461,N_1495);
and U1591 (N_1591,N_1489,N_1400);
nand U1592 (N_1592,N_1498,N_1427);
and U1593 (N_1593,N_1494,N_1406);
or U1594 (N_1594,N_1457,N_1413);
nor U1595 (N_1595,N_1493,N_1440);
nor U1596 (N_1596,N_1463,N_1481);
and U1597 (N_1597,N_1469,N_1410);
nor U1598 (N_1598,N_1455,N_1422);
and U1599 (N_1599,N_1469,N_1498);
nand U1600 (N_1600,N_1535,N_1572);
nand U1601 (N_1601,N_1500,N_1534);
or U1602 (N_1602,N_1564,N_1553);
nor U1603 (N_1603,N_1516,N_1510);
or U1604 (N_1604,N_1504,N_1532);
xor U1605 (N_1605,N_1547,N_1527);
nor U1606 (N_1606,N_1568,N_1587);
nand U1607 (N_1607,N_1530,N_1543);
nand U1608 (N_1608,N_1573,N_1581);
nor U1609 (N_1609,N_1597,N_1550);
nand U1610 (N_1610,N_1554,N_1537);
nand U1611 (N_1611,N_1552,N_1520);
and U1612 (N_1612,N_1517,N_1565);
and U1613 (N_1613,N_1596,N_1570);
nor U1614 (N_1614,N_1525,N_1590);
or U1615 (N_1615,N_1558,N_1578);
and U1616 (N_1616,N_1509,N_1592);
nand U1617 (N_1617,N_1585,N_1577);
and U1618 (N_1618,N_1508,N_1519);
nor U1619 (N_1619,N_1546,N_1513);
nor U1620 (N_1620,N_1584,N_1561);
nand U1621 (N_1621,N_1599,N_1563);
and U1622 (N_1622,N_1544,N_1515);
or U1623 (N_1623,N_1583,N_1507);
nor U1624 (N_1624,N_1538,N_1523);
and U1625 (N_1625,N_1506,N_1566);
nand U1626 (N_1626,N_1528,N_1594);
and U1627 (N_1627,N_1512,N_1560);
nor U1628 (N_1628,N_1505,N_1571);
nor U1629 (N_1629,N_1501,N_1548);
nand U1630 (N_1630,N_1569,N_1589);
nand U1631 (N_1631,N_1522,N_1531);
and U1632 (N_1632,N_1562,N_1502);
nand U1633 (N_1633,N_1524,N_1511);
and U1634 (N_1634,N_1586,N_1514);
nor U1635 (N_1635,N_1556,N_1557);
or U1636 (N_1636,N_1580,N_1539);
or U1637 (N_1637,N_1576,N_1503);
and U1638 (N_1638,N_1591,N_1521);
nor U1639 (N_1639,N_1588,N_1545);
nand U1640 (N_1640,N_1551,N_1559);
and U1641 (N_1641,N_1526,N_1598);
nand U1642 (N_1642,N_1549,N_1593);
or U1643 (N_1643,N_1555,N_1575);
and U1644 (N_1644,N_1541,N_1533);
or U1645 (N_1645,N_1595,N_1542);
or U1646 (N_1646,N_1567,N_1582);
nand U1647 (N_1647,N_1540,N_1529);
or U1648 (N_1648,N_1574,N_1518);
nand U1649 (N_1649,N_1536,N_1579);
nand U1650 (N_1650,N_1539,N_1543);
or U1651 (N_1651,N_1544,N_1592);
and U1652 (N_1652,N_1599,N_1568);
nand U1653 (N_1653,N_1585,N_1576);
nand U1654 (N_1654,N_1586,N_1545);
nand U1655 (N_1655,N_1524,N_1513);
nor U1656 (N_1656,N_1543,N_1507);
nand U1657 (N_1657,N_1558,N_1520);
or U1658 (N_1658,N_1573,N_1563);
nand U1659 (N_1659,N_1546,N_1594);
nor U1660 (N_1660,N_1554,N_1599);
nor U1661 (N_1661,N_1594,N_1507);
nand U1662 (N_1662,N_1550,N_1547);
and U1663 (N_1663,N_1514,N_1564);
or U1664 (N_1664,N_1536,N_1591);
and U1665 (N_1665,N_1588,N_1527);
nor U1666 (N_1666,N_1580,N_1516);
or U1667 (N_1667,N_1531,N_1581);
xor U1668 (N_1668,N_1538,N_1560);
or U1669 (N_1669,N_1572,N_1544);
or U1670 (N_1670,N_1593,N_1530);
and U1671 (N_1671,N_1526,N_1515);
and U1672 (N_1672,N_1515,N_1509);
nor U1673 (N_1673,N_1508,N_1592);
and U1674 (N_1674,N_1588,N_1569);
nor U1675 (N_1675,N_1591,N_1562);
or U1676 (N_1676,N_1572,N_1592);
nor U1677 (N_1677,N_1558,N_1518);
and U1678 (N_1678,N_1510,N_1595);
nand U1679 (N_1679,N_1504,N_1503);
and U1680 (N_1680,N_1569,N_1502);
nand U1681 (N_1681,N_1579,N_1558);
or U1682 (N_1682,N_1540,N_1537);
nor U1683 (N_1683,N_1569,N_1544);
nor U1684 (N_1684,N_1584,N_1564);
nor U1685 (N_1685,N_1547,N_1572);
or U1686 (N_1686,N_1582,N_1518);
and U1687 (N_1687,N_1518,N_1507);
nand U1688 (N_1688,N_1595,N_1505);
and U1689 (N_1689,N_1589,N_1547);
or U1690 (N_1690,N_1572,N_1567);
and U1691 (N_1691,N_1553,N_1554);
nand U1692 (N_1692,N_1522,N_1535);
nand U1693 (N_1693,N_1584,N_1501);
or U1694 (N_1694,N_1571,N_1520);
xor U1695 (N_1695,N_1540,N_1512);
and U1696 (N_1696,N_1538,N_1541);
nand U1697 (N_1697,N_1577,N_1575);
nand U1698 (N_1698,N_1538,N_1505);
nor U1699 (N_1699,N_1507,N_1595);
and U1700 (N_1700,N_1623,N_1692);
and U1701 (N_1701,N_1610,N_1688);
or U1702 (N_1702,N_1622,N_1613);
nand U1703 (N_1703,N_1638,N_1618);
nor U1704 (N_1704,N_1607,N_1637);
xor U1705 (N_1705,N_1639,N_1633);
and U1706 (N_1706,N_1624,N_1691);
nor U1707 (N_1707,N_1629,N_1602);
or U1708 (N_1708,N_1676,N_1620);
xnor U1709 (N_1709,N_1634,N_1668);
or U1710 (N_1710,N_1601,N_1677);
nor U1711 (N_1711,N_1650,N_1681);
nor U1712 (N_1712,N_1645,N_1615);
and U1713 (N_1713,N_1687,N_1664);
and U1714 (N_1714,N_1671,N_1667);
nor U1715 (N_1715,N_1636,N_1665);
or U1716 (N_1716,N_1680,N_1698);
or U1717 (N_1717,N_1648,N_1619);
or U1718 (N_1718,N_1684,N_1647);
nor U1719 (N_1719,N_1616,N_1657);
or U1720 (N_1720,N_1612,N_1694);
nor U1721 (N_1721,N_1654,N_1682);
and U1722 (N_1722,N_1621,N_1672);
or U1723 (N_1723,N_1693,N_1641);
nor U1724 (N_1724,N_1630,N_1690);
or U1725 (N_1725,N_1656,N_1609);
and U1726 (N_1726,N_1652,N_1663);
nand U1727 (N_1727,N_1697,N_1658);
nand U1728 (N_1728,N_1651,N_1699);
and U1729 (N_1729,N_1640,N_1614);
nand U1730 (N_1730,N_1662,N_1600);
or U1731 (N_1731,N_1649,N_1605);
nand U1732 (N_1732,N_1673,N_1695);
and U1733 (N_1733,N_1683,N_1661);
nand U1734 (N_1734,N_1653,N_1689);
nor U1735 (N_1735,N_1627,N_1679);
nand U1736 (N_1736,N_1655,N_1644);
nor U1737 (N_1737,N_1631,N_1611);
or U1738 (N_1738,N_1660,N_1626);
xor U1739 (N_1739,N_1678,N_1606);
nand U1740 (N_1740,N_1617,N_1685);
or U1741 (N_1741,N_1659,N_1669);
nand U1742 (N_1742,N_1674,N_1643);
or U1743 (N_1743,N_1686,N_1608);
or U1744 (N_1744,N_1642,N_1603);
nand U1745 (N_1745,N_1696,N_1632);
and U1746 (N_1746,N_1666,N_1670);
or U1747 (N_1747,N_1646,N_1628);
or U1748 (N_1748,N_1635,N_1604);
xor U1749 (N_1749,N_1625,N_1675);
nor U1750 (N_1750,N_1637,N_1601);
and U1751 (N_1751,N_1606,N_1673);
nor U1752 (N_1752,N_1696,N_1605);
nor U1753 (N_1753,N_1684,N_1688);
nor U1754 (N_1754,N_1628,N_1603);
or U1755 (N_1755,N_1647,N_1619);
or U1756 (N_1756,N_1676,N_1649);
nand U1757 (N_1757,N_1690,N_1642);
or U1758 (N_1758,N_1662,N_1665);
nor U1759 (N_1759,N_1686,N_1655);
or U1760 (N_1760,N_1648,N_1609);
and U1761 (N_1761,N_1620,N_1698);
nand U1762 (N_1762,N_1640,N_1672);
xor U1763 (N_1763,N_1690,N_1664);
or U1764 (N_1764,N_1677,N_1624);
or U1765 (N_1765,N_1601,N_1626);
or U1766 (N_1766,N_1628,N_1641);
and U1767 (N_1767,N_1646,N_1618);
nand U1768 (N_1768,N_1657,N_1663);
and U1769 (N_1769,N_1639,N_1666);
or U1770 (N_1770,N_1613,N_1696);
nand U1771 (N_1771,N_1695,N_1615);
nor U1772 (N_1772,N_1653,N_1680);
nor U1773 (N_1773,N_1604,N_1668);
xor U1774 (N_1774,N_1641,N_1604);
and U1775 (N_1775,N_1625,N_1678);
or U1776 (N_1776,N_1604,N_1603);
nor U1777 (N_1777,N_1650,N_1666);
or U1778 (N_1778,N_1604,N_1651);
or U1779 (N_1779,N_1664,N_1641);
and U1780 (N_1780,N_1608,N_1610);
nand U1781 (N_1781,N_1608,N_1691);
nand U1782 (N_1782,N_1600,N_1668);
nor U1783 (N_1783,N_1633,N_1623);
nor U1784 (N_1784,N_1602,N_1653);
and U1785 (N_1785,N_1634,N_1659);
or U1786 (N_1786,N_1634,N_1639);
nor U1787 (N_1787,N_1682,N_1658);
xor U1788 (N_1788,N_1649,N_1621);
nand U1789 (N_1789,N_1658,N_1690);
nor U1790 (N_1790,N_1669,N_1645);
nand U1791 (N_1791,N_1689,N_1608);
nand U1792 (N_1792,N_1661,N_1694);
or U1793 (N_1793,N_1685,N_1636);
and U1794 (N_1794,N_1672,N_1693);
or U1795 (N_1795,N_1640,N_1692);
nand U1796 (N_1796,N_1655,N_1678);
xor U1797 (N_1797,N_1656,N_1676);
and U1798 (N_1798,N_1696,N_1681);
or U1799 (N_1799,N_1696,N_1602);
nor U1800 (N_1800,N_1765,N_1740);
nor U1801 (N_1801,N_1726,N_1718);
nand U1802 (N_1802,N_1753,N_1700);
or U1803 (N_1803,N_1711,N_1735);
or U1804 (N_1804,N_1799,N_1792);
nor U1805 (N_1805,N_1703,N_1755);
or U1806 (N_1806,N_1757,N_1778);
or U1807 (N_1807,N_1720,N_1713);
or U1808 (N_1808,N_1791,N_1717);
xnor U1809 (N_1809,N_1721,N_1732);
nor U1810 (N_1810,N_1752,N_1743);
and U1811 (N_1811,N_1716,N_1722);
nand U1812 (N_1812,N_1744,N_1771);
nand U1813 (N_1813,N_1729,N_1706);
or U1814 (N_1814,N_1746,N_1764);
xor U1815 (N_1815,N_1714,N_1793);
and U1816 (N_1816,N_1769,N_1787);
xor U1817 (N_1817,N_1773,N_1772);
nor U1818 (N_1818,N_1761,N_1739);
and U1819 (N_1819,N_1785,N_1727);
nor U1820 (N_1820,N_1798,N_1704);
or U1821 (N_1821,N_1719,N_1725);
nor U1822 (N_1822,N_1745,N_1749);
nor U1823 (N_1823,N_1741,N_1760);
nand U1824 (N_1824,N_1707,N_1774);
nor U1825 (N_1825,N_1750,N_1770);
and U1826 (N_1826,N_1781,N_1758);
nand U1827 (N_1827,N_1784,N_1782);
or U1828 (N_1828,N_1754,N_1797);
nor U1829 (N_1829,N_1783,N_1728);
nand U1830 (N_1830,N_1756,N_1767);
and U1831 (N_1831,N_1724,N_1738);
and U1832 (N_1832,N_1789,N_1747);
nand U1833 (N_1833,N_1790,N_1709);
nor U1834 (N_1834,N_1705,N_1708);
and U1835 (N_1835,N_1780,N_1734);
nand U1836 (N_1836,N_1715,N_1731);
and U1837 (N_1837,N_1701,N_1763);
nand U1838 (N_1838,N_1723,N_1779);
or U1839 (N_1839,N_1710,N_1733);
and U1840 (N_1840,N_1712,N_1788);
or U1841 (N_1841,N_1766,N_1759);
nand U1842 (N_1842,N_1736,N_1777);
or U1843 (N_1843,N_1795,N_1751);
nand U1844 (N_1844,N_1737,N_1796);
or U1845 (N_1845,N_1748,N_1762);
nor U1846 (N_1846,N_1786,N_1768);
nand U1847 (N_1847,N_1730,N_1742);
nand U1848 (N_1848,N_1702,N_1775);
or U1849 (N_1849,N_1794,N_1776);
or U1850 (N_1850,N_1795,N_1719);
and U1851 (N_1851,N_1776,N_1791);
nor U1852 (N_1852,N_1770,N_1751);
and U1853 (N_1853,N_1788,N_1711);
nand U1854 (N_1854,N_1728,N_1702);
and U1855 (N_1855,N_1744,N_1796);
nor U1856 (N_1856,N_1764,N_1728);
xor U1857 (N_1857,N_1746,N_1718);
xnor U1858 (N_1858,N_1782,N_1749);
and U1859 (N_1859,N_1786,N_1755);
nand U1860 (N_1860,N_1738,N_1779);
nand U1861 (N_1861,N_1737,N_1728);
nand U1862 (N_1862,N_1793,N_1709);
nor U1863 (N_1863,N_1745,N_1750);
or U1864 (N_1864,N_1766,N_1731);
nor U1865 (N_1865,N_1748,N_1719);
nor U1866 (N_1866,N_1779,N_1729);
nor U1867 (N_1867,N_1783,N_1725);
nand U1868 (N_1868,N_1723,N_1761);
nor U1869 (N_1869,N_1750,N_1701);
or U1870 (N_1870,N_1752,N_1762);
xnor U1871 (N_1871,N_1782,N_1713);
nor U1872 (N_1872,N_1711,N_1718);
and U1873 (N_1873,N_1767,N_1737);
nand U1874 (N_1874,N_1743,N_1737);
nor U1875 (N_1875,N_1712,N_1703);
and U1876 (N_1876,N_1763,N_1738);
nand U1877 (N_1877,N_1708,N_1740);
nor U1878 (N_1878,N_1793,N_1766);
and U1879 (N_1879,N_1790,N_1719);
nor U1880 (N_1880,N_1789,N_1777);
xnor U1881 (N_1881,N_1720,N_1787);
nand U1882 (N_1882,N_1769,N_1770);
nor U1883 (N_1883,N_1719,N_1718);
or U1884 (N_1884,N_1708,N_1714);
nor U1885 (N_1885,N_1756,N_1712);
nand U1886 (N_1886,N_1716,N_1765);
and U1887 (N_1887,N_1769,N_1724);
nand U1888 (N_1888,N_1731,N_1704);
nor U1889 (N_1889,N_1713,N_1761);
or U1890 (N_1890,N_1790,N_1730);
and U1891 (N_1891,N_1799,N_1729);
nand U1892 (N_1892,N_1719,N_1717);
or U1893 (N_1893,N_1731,N_1756);
and U1894 (N_1894,N_1794,N_1762);
nor U1895 (N_1895,N_1707,N_1758);
nor U1896 (N_1896,N_1734,N_1713);
and U1897 (N_1897,N_1706,N_1784);
nand U1898 (N_1898,N_1714,N_1758);
or U1899 (N_1899,N_1790,N_1715);
or U1900 (N_1900,N_1800,N_1873);
nand U1901 (N_1901,N_1858,N_1886);
or U1902 (N_1902,N_1808,N_1820);
and U1903 (N_1903,N_1894,N_1850);
or U1904 (N_1904,N_1893,N_1888);
and U1905 (N_1905,N_1853,N_1803);
nand U1906 (N_1906,N_1848,N_1824);
and U1907 (N_1907,N_1863,N_1859);
and U1908 (N_1908,N_1841,N_1831);
and U1909 (N_1909,N_1818,N_1851);
nand U1910 (N_1910,N_1891,N_1814);
nand U1911 (N_1911,N_1829,N_1849);
nor U1912 (N_1912,N_1882,N_1826);
nor U1913 (N_1913,N_1867,N_1811);
or U1914 (N_1914,N_1855,N_1857);
or U1915 (N_1915,N_1835,N_1898);
and U1916 (N_1916,N_1843,N_1889);
nand U1917 (N_1917,N_1812,N_1881);
nor U1918 (N_1918,N_1887,N_1842);
nand U1919 (N_1919,N_1844,N_1836);
or U1920 (N_1920,N_1871,N_1883);
nand U1921 (N_1921,N_1813,N_1874);
xnor U1922 (N_1922,N_1884,N_1864);
nor U1923 (N_1923,N_1823,N_1827);
nor U1924 (N_1924,N_1825,N_1838);
xor U1925 (N_1925,N_1876,N_1805);
or U1926 (N_1926,N_1847,N_1892);
nand U1927 (N_1927,N_1895,N_1807);
xor U1928 (N_1928,N_1804,N_1861);
or U1929 (N_1929,N_1899,N_1802);
nor U1930 (N_1930,N_1879,N_1862);
and U1931 (N_1931,N_1837,N_1880);
nand U1932 (N_1932,N_1806,N_1817);
and U1933 (N_1933,N_1845,N_1860);
or U1934 (N_1934,N_1877,N_1821);
or U1935 (N_1935,N_1815,N_1828);
nand U1936 (N_1936,N_1869,N_1822);
nor U1937 (N_1937,N_1868,N_1832);
nand U1938 (N_1938,N_1872,N_1897);
and U1939 (N_1939,N_1865,N_1875);
and U1940 (N_1940,N_1866,N_1856);
nand U1941 (N_1941,N_1809,N_1839);
nor U1942 (N_1942,N_1834,N_1819);
nor U1943 (N_1943,N_1816,N_1833);
or U1944 (N_1944,N_1830,N_1854);
or U1945 (N_1945,N_1890,N_1885);
or U1946 (N_1946,N_1878,N_1810);
nand U1947 (N_1947,N_1852,N_1840);
xor U1948 (N_1948,N_1846,N_1896);
and U1949 (N_1949,N_1870,N_1801);
nand U1950 (N_1950,N_1860,N_1843);
and U1951 (N_1951,N_1847,N_1883);
or U1952 (N_1952,N_1806,N_1800);
nor U1953 (N_1953,N_1856,N_1859);
nor U1954 (N_1954,N_1843,N_1866);
nor U1955 (N_1955,N_1882,N_1871);
and U1956 (N_1956,N_1864,N_1853);
nand U1957 (N_1957,N_1876,N_1842);
nor U1958 (N_1958,N_1862,N_1872);
or U1959 (N_1959,N_1817,N_1852);
nor U1960 (N_1960,N_1888,N_1863);
and U1961 (N_1961,N_1861,N_1809);
nor U1962 (N_1962,N_1866,N_1815);
nor U1963 (N_1963,N_1897,N_1892);
nand U1964 (N_1964,N_1819,N_1865);
and U1965 (N_1965,N_1881,N_1801);
or U1966 (N_1966,N_1814,N_1892);
nor U1967 (N_1967,N_1858,N_1880);
nor U1968 (N_1968,N_1824,N_1895);
or U1969 (N_1969,N_1812,N_1890);
nand U1970 (N_1970,N_1883,N_1874);
nor U1971 (N_1971,N_1879,N_1887);
and U1972 (N_1972,N_1814,N_1821);
or U1973 (N_1973,N_1873,N_1881);
nand U1974 (N_1974,N_1819,N_1848);
or U1975 (N_1975,N_1820,N_1819);
and U1976 (N_1976,N_1825,N_1821);
and U1977 (N_1977,N_1858,N_1881);
and U1978 (N_1978,N_1861,N_1825);
and U1979 (N_1979,N_1896,N_1866);
nand U1980 (N_1980,N_1845,N_1875);
or U1981 (N_1981,N_1827,N_1844);
nand U1982 (N_1982,N_1899,N_1853);
nand U1983 (N_1983,N_1881,N_1854);
or U1984 (N_1984,N_1844,N_1857);
or U1985 (N_1985,N_1884,N_1811);
or U1986 (N_1986,N_1839,N_1893);
nand U1987 (N_1987,N_1883,N_1889);
or U1988 (N_1988,N_1885,N_1847);
or U1989 (N_1989,N_1882,N_1835);
nor U1990 (N_1990,N_1830,N_1897);
nor U1991 (N_1991,N_1841,N_1842);
or U1992 (N_1992,N_1840,N_1809);
nor U1993 (N_1993,N_1835,N_1862);
or U1994 (N_1994,N_1847,N_1836);
nand U1995 (N_1995,N_1896,N_1823);
nor U1996 (N_1996,N_1818,N_1881);
and U1997 (N_1997,N_1847,N_1870);
nand U1998 (N_1998,N_1886,N_1847);
and U1999 (N_1999,N_1851,N_1829);
nand U2000 (N_2000,N_1922,N_1985);
and U2001 (N_2001,N_1949,N_1952);
nor U2002 (N_2002,N_1973,N_1900);
nand U2003 (N_2003,N_1914,N_1953);
or U2004 (N_2004,N_1912,N_1906);
nor U2005 (N_2005,N_1980,N_1966);
nand U2006 (N_2006,N_1988,N_1908);
nand U2007 (N_2007,N_1916,N_1942);
or U2008 (N_2008,N_1928,N_1948);
and U2009 (N_2009,N_1934,N_1929);
nor U2010 (N_2010,N_1998,N_1992);
and U2011 (N_2011,N_1956,N_1958);
and U2012 (N_2012,N_1936,N_1911);
nand U2013 (N_2013,N_1935,N_1984);
and U2014 (N_2014,N_1937,N_1947);
nand U2015 (N_2015,N_1990,N_1991);
nor U2016 (N_2016,N_1976,N_1975);
or U2017 (N_2017,N_1959,N_1963);
and U2018 (N_2018,N_1915,N_1999);
nand U2019 (N_2019,N_1968,N_1967);
nor U2020 (N_2020,N_1931,N_1905);
nor U2021 (N_2021,N_1920,N_1932);
nor U2022 (N_2022,N_1971,N_1978);
nor U2023 (N_2023,N_1977,N_1945);
nand U2024 (N_2024,N_1909,N_1981);
or U2025 (N_2025,N_1944,N_1960);
and U2026 (N_2026,N_1995,N_1965);
nand U2027 (N_2027,N_1940,N_1903);
nor U2028 (N_2028,N_1974,N_1939);
or U2029 (N_2029,N_1902,N_1989);
and U2030 (N_2030,N_1913,N_1983);
and U2031 (N_2031,N_1964,N_1962);
nand U2032 (N_2032,N_1982,N_1950);
nand U2033 (N_2033,N_1970,N_1930);
nor U2034 (N_2034,N_1987,N_1919);
nor U2035 (N_2035,N_1972,N_1925);
nand U2036 (N_2036,N_1933,N_1997);
nor U2037 (N_2037,N_1943,N_1993);
nor U2038 (N_2038,N_1921,N_1955);
nor U2039 (N_2039,N_1996,N_1951);
and U2040 (N_2040,N_1917,N_1904);
or U2041 (N_2041,N_1923,N_1918);
and U2042 (N_2042,N_1994,N_1961);
nand U2043 (N_2043,N_1926,N_1954);
and U2044 (N_2044,N_1901,N_1957);
nor U2045 (N_2045,N_1938,N_1979);
nor U2046 (N_2046,N_1907,N_1910);
or U2047 (N_2047,N_1946,N_1986);
nor U2048 (N_2048,N_1924,N_1941);
or U2049 (N_2049,N_1927,N_1969);
or U2050 (N_2050,N_1955,N_1948);
nor U2051 (N_2051,N_1982,N_1993);
and U2052 (N_2052,N_1971,N_1926);
nand U2053 (N_2053,N_1957,N_1961);
or U2054 (N_2054,N_1918,N_1950);
nor U2055 (N_2055,N_1992,N_1987);
nand U2056 (N_2056,N_1942,N_1905);
and U2057 (N_2057,N_1916,N_1965);
nand U2058 (N_2058,N_1960,N_1953);
and U2059 (N_2059,N_1912,N_1999);
and U2060 (N_2060,N_1961,N_1969);
nor U2061 (N_2061,N_1940,N_1907);
or U2062 (N_2062,N_1926,N_1938);
and U2063 (N_2063,N_1906,N_1928);
and U2064 (N_2064,N_1992,N_1910);
or U2065 (N_2065,N_1953,N_1992);
or U2066 (N_2066,N_1950,N_1965);
nand U2067 (N_2067,N_1935,N_1947);
and U2068 (N_2068,N_1991,N_1933);
nor U2069 (N_2069,N_1978,N_1958);
nand U2070 (N_2070,N_1978,N_1976);
or U2071 (N_2071,N_1996,N_1988);
nand U2072 (N_2072,N_1901,N_1956);
or U2073 (N_2073,N_1948,N_1923);
nand U2074 (N_2074,N_1906,N_1947);
nand U2075 (N_2075,N_1974,N_1918);
and U2076 (N_2076,N_1974,N_1992);
or U2077 (N_2077,N_1959,N_1954);
nor U2078 (N_2078,N_1924,N_1995);
nor U2079 (N_2079,N_1955,N_1902);
nand U2080 (N_2080,N_1960,N_1942);
or U2081 (N_2081,N_1920,N_1962);
or U2082 (N_2082,N_1920,N_1927);
nor U2083 (N_2083,N_1936,N_1962);
and U2084 (N_2084,N_1936,N_1999);
and U2085 (N_2085,N_1983,N_1901);
nor U2086 (N_2086,N_1961,N_1960);
nand U2087 (N_2087,N_1916,N_1985);
and U2088 (N_2088,N_1981,N_1987);
nand U2089 (N_2089,N_1939,N_1969);
nor U2090 (N_2090,N_1956,N_1992);
and U2091 (N_2091,N_1938,N_1912);
nand U2092 (N_2092,N_1983,N_1990);
or U2093 (N_2093,N_1909,N_1989);
and U2094 (N_2094,N_1959,N_1907);
or U2095 (N_2095,N_1995,N_1991);
and U2096 (N_2096,N_1955,N_1928);
nand U2097 (N_2097,N_1948,N_1921);
and U2098 (N_2098,N_1990,N_1917);
nand U2099 (N_2099,N_1985,N_1940);
nor U2100 (N_2100,N_2055,N_2018);
and U2101 (N_2101,N_2046,N_2088);
or U2102 (N_2102,N_2041,N_2062);
nor U2103 (N_2103,N_2039,N_2001);
nand U2104 (N_2104,N_2028,N_2094);
xor U2105 (N_2105,N_2006,N_2075);
nand U2106 (N_2106,N_2054,N_2071);
nand U2107 (N_2107,N_2012,N_2030);
or U2108 (N_2108,N_2096,N_2080);
nor U2109 (N_2109,N_2025,N_2031);
or U2110 (N_2110,N_2020,N_2005);
and U2111 (N_2111,N_2082,N_2023);
and U2112 (N_2112,N_2092,N_2078);
and U2113 (N_2113,N_2087,N_2069);
and U2114 (N_2114,N_2060,N_2059);
nor U2115 (N_2115,N_2061,N_2016);
or U2116 (N_2116,N_2007,N_2033);
nand U2117 (N_2117,N_2019,N_2026);
and U2118 (N_2118,N_2093,N_2050);
nand U2119 (N_2119,N_2065,N_2052);
or U2120 (N_2120,N_2097,N_2017);
nor U2121 (N_2121,N_2064,N_2038);
nor U2122 (N_2122,N_2044,N_2066);
and U2123 (N_2123,N_2009,N_2027);
or U2124 (N_2124,N_2058,N_2013);
nor U2125 (N_2125,N_2004,N_2089);
nand U2126 (N_2126,N_2008,N_2090);
nor U2127 (N_2127,N_2081,N_2049);
and U2128 (N_2128,N_2032,N_2079);
and U2129 (N_2129,N_2015,N_2011);
nand U2130 (N_2130,N_2073,N_2002);
or U2131 (N_2131,N_2095,N_2003);
nor U2132 (N_2132,N_2048,N_2068);
nand U2133 (N_2133,N_2014,N_2034);
nand U2134 (N_2134,N_2042,N_2036);
nand U2135 (N_2135,N_2099,N_2035);
or U2136 (N_2136,N_2076,N_2057);
or U2137 (N_2137,N_2084,N_2083);
or U2138 (N_2138,N_2067,N_2086);
and U2139 (N_2139,N_2063,N_2072);
or U2140 (N_2140,N_2070,N_2037);
or U2141 (N_2141,N_2085,N_2021);
nand U2142 (N_2142,N_2047,N_2040);
nand U2143 (N_2143,N_2045,N_2053);
nand U2144 (N_2144,N_2010,N_2051);
nor U2145 (N_2145,N_2091,N_2074);
xor U2146 (N_2146,N_2077,N_2022);
nand U2147 (N_2147,N_2043,N_2024);
or U2148 (N_2148,N_2098,N_2056);
nor U2149 (N_2149,N_2029,N_2000);
and U2150 (N_2150,N_2008,N_2006);
nand U2151 (N_2151,N_2062,N_2007);
and U2152 (N_2152,N_2082,N_2033);
nand U2153 (N_2153,N_2035,N_2032);
or U2154 (N_2154,N_2002,N_2030);
nand U2155 (N_2155,N_2023,N_2060);
nor U2156 (N_2156,N_2045,N_2093);
nor U2157 (N_2157,N_2083,N_2017);
or U2158 (N_2158,N_2015,N_2056);
or U2159 (N_2159,N_2007,N_2082);
or U2160 (N_2160,N_2054,N_2045);
nand U2161 (N_2161,N_2060,N_2038);
and U2162 (N_2162,N_2000,N_2015);
nand U2163 (N_2163,N_2045,N_2057);
nor U2164 (N_2164,N_2062,N_2019);
and U2165 (N_2165,N_2003,N_2024);
or U2166 (N_2166,N_2013,N_2031);
and U2167 (N_2167,N_2041,N_2092);
or U2168 (N_2168,N_2064,N_2019);
nand U2169 (N_2169,N_2057,N_2067);
nor U2170 (N_2170,N_2096,N_2076);
nor U2171 (N_2171,N_2064,N_2002);
nand U2172 (N_2172,N_2092,N_2021);
and U2173 (N_2173,N_2030,N_2026);
nand U2174 (N_2174,N_2033,N_2060);
or U2175 (N_2175,N_2029,N_2016);
and U2176 (N_2176,N_2092,N_2050);
nand U2177 (N_2177,N_2046,N_2030);
nor U2178 (N_2178,N_2005,N_2050);
or U2179 (N_2179,N_2067,N_2039);
and U2180 (N_2180,N_2088,N_2041);
or U2181 (N_2181,N_2010,N_2076);
nor U2182 (N_2182,N_2033,N_2067);
nor U2183 (N_2183,N_2009,N_2022);
nand U2184 (N_2184,N_2032,N_2072);
or U2185 (N_2185,N_2064,N_2095);
nand U2186 (N_2186,N_2016,N_2079);
nand U2187 (N_2187,N_2051,N_2008);
and U2188 (N_2188,N_2021,N_2093);
or U2189 (N_2189,N_2063,N_2003);
nor U2190 (N_2190,N_2093,N_2035);
xor U2191 (N_2191,N_2034,N_2030);
xor U2192 (N_2192,N_2019,N_2008);
nand U2193 (N_2193,N_2035,N_2062);
nand U2194 (N_2194,N_2057,N_2088);
or U2195 (N_2195,N_2026,N_2004);
and U2196 (N_2196,N_2096,N_2050);
and U2197 (N_2197,N_2025,N_2086);
or U2198 (N_2198,N_2097,N_2072);
nor U2199 (N_2199,N_2045,N_2019);
or U2200 (N_2200,N_2177,N_2172);
nor U2201 (N_2201,N_2145,N_2159);
nor U2202 (N_2202,N_2179,N_2123);
xnor U2203 (N_2203,N_2132,N_2185);
nand U2204 (N_2204,N_2100,N_2106);
nand U2205 (N_2205,N_2197,N_2141);
nand U2206 (N_2206,N_2144,N_2109);
and U2207 (N_2207,N_2157,N_2108);
or U2208 (N_2208,N_2127,N_2174);
or U2209 (N_2209,N_2161,N_2135);
and U2210 (N_2210,N_2122,N_2110);
or U2211 (N_2211,N_2117,N_2175);
or U2212 (N_2212,N_2107,N_2111);
and U2213 (N_2213,N_2136,N_2126);
xor U2214 (N_2214,N_2162,N_2189);
nand U2215 (N_2215,N_2143,N_2102);
and U2216 (N_2216,N_2140,N_2182);
nor U2217 (N_2217,N_2173,N_2104);
and U2218 (N_2218,N_2184,N_2134);
nor U2219 (N_2219,N_2166,N_2116);
and U2220 (N_2220,N_2198,N_2149);
nor U2221 (N_2221,N_2120,N_2180);
or U2222 (N_2222,N_2169,N_2158);
nand U2223 (N_2223,N_2115,N_2130);
and U2224 (N_2224,N_2187,N_2196);
xor U2225 (N_2225,N_2105,N_2155);
and U2226 (N_2226,N_2192,N_2178);
or U2227 (N_2227,N_2131,N_2101);
nor U2228 (N_2228,N_2183,N_2191);
nand U2229 (N_2229,N_2171,N_2112);
or U2230 (N_2230,N_2121,N_2113);
and U2231 (N_2231,N_2193,N_2188);
or U2232 (N_2232,N_2165,N_2103);
and U2233 (N_2233,N_2147,N_2199);
nand U2234 (N_2234,N_2133,N_2148);
nor U2235 (N_2235,N_2160,N_2153);
or U2236 (N_2236,N_2139,N_2167);
or U2237 (N_2237,N_2137,N_2186);
nor U2238 (N_2238,N_2118,N_2164);
nand U2239 (N_2239,N_2194,N_2138);
nor U2240 (N_2240,N_2190,N_2170);
and U2241 (N_2241,N_2150,N_2163);
or U2242 (N_2242,N_2125,N_2146);
and U2243 (N_2243,N_2154,N_2176);
and U2244 (N_2244,N_2181,N_2168);
nand U2245 (N_2245,N_2129,N_2156);
nand U2246 (N_2246,N_2142,N_2114);
xor U2247 (N_2247,N_2128,N_2152);
nor U2248 (N_2248,N_2119,N_2195);
nand U2249 (N_2249,N_2151,N_2124);
or U2250 (N_2250,N_2181,N_2119);
and U2251 (N_2251,N_2157,N_2169);
or U2252 (N_2252,N_2109,N_2164);
and U2253 (N_2253,N_2161,N_2114);
and U2254 (N_2254,N_2101,N_2187);
and U2255 (N_2255,N_2158,N_2143);
or U2256 (N_2256,N_2124,N_2166);
nand U2257 (N_2257,N_2149,N_2163);
nand U2258 (N_2258,N_2106,N_2156);
nand U2259 (N_2259,N_2188,N_2158);
and U2260 (N_2260,N_2187,N_2139);
xnor U2261 (N_2261,N_2176,N_2101);
nor U2262 (N_2262,N_2164,N_2151);
or U2263 (N_2263,N_2165,N_2184);
nor U2264 (N_2264,N_2172,N_2169);
and U2265 (N_2265,N_2123,N_2140);
or U2266 (N_2266,N_2142,N_2138);
and U2267 (N_2267,N_2147,N_2114);
nor U2268 (N_2268,N_2170,N_2140);
and U2269 (N_2269,N_2154,N_2164);
xnor U2270 (N_2270,N_2158,N_2176);
nand U2271 (N_2271,N_2127,N_2171);
and U2272 (N_2272,N_2181,N_2171);
and U2273 (N_2273,N_2160,N_2134);
or U2274 (N_2274,N_2157,N_2183);
nor U2275 (N_2275,N_2196,N_2182);
nand U2276 (N_2276,N_2114,N_2133);
nor U2277 (N_2277,N_2170,N_2182);
and U2278 (N_2278,N_2189,N_2146);
or U2279 (N_2279,N_2102,N_2113);
and U2280 (N_2280,N_2125,N_2192);
nor U2281 (N_2281,N_2182,N_2198);
nor U2282 (N_2282,N_2126,N_2107);
nor U2283 (N_2283,N_2118,N_2192);
nand U2284 (N_2284,N_2197,N_2116);
nor U2285 (N_2285,N_2132,N_2100);
and U2286 (N_2286,N_2183,N_2159);
and U2287 (N_2287,N_2186,N_2113);
nor U2288 (N_2288,N_2147,N_2115);
and U2289 (N_2289,N_2155,N_2188);
xnor U2290 (N_2290,N_2199,N_2145);
or U2291 (N_2291,N_2133,N_2138);
and U2292 (N_2292,N_2144,N_2187);
or U2293 (N_2293,N_2178,N_2179);
or U2294 (N_2294,N_2179,N_2106);
nor U2295 (N_2295,N_2189,N_2164);
nor U2296 (N_2296,N_2136,N_2130);
nand U2297 (N_2297,N_2163,N_2158);
and U2298 (N_2298,N_2113,N_2160);
nor U2299 (N_2299,N_2183,N_2102);
nor U2300 (N_2300,N_2211,N_2241);
xor U2301 (N_2301,N_2275,N_2219);
nand U2302 (N_2302,N_2276,N_2285);
or U2303 (N_2303,N_2260,N_2256);
and U2304 (N_2304,N_2247,N_2265);
and U2305 (N_2305,N_2281,N_2224);
nor U2306 (N_2306,N_2272,N_2287);
nor U2307 (N_2307,N_2289,N_2296);
nand U2308 (N_2308,N_2283,N_2259);
and U2309 (N_2309,N_2203,N_2210);
nor U2310 (N_2310,N_2294,N_2233);
nor U2311 (N_2311,N_2274,N_2288);
nand U2312 (N_2312,N_2269,N_2243);
and U2313 (N_2313,N_2250,N_2229);
and U2314 (N_2314,N_2220,N_2201);
nor U2315 (N_2315,N_2251,N_2235);
or U2316 (N_2316,N_2222,N_2290);
nand U2317 (N_2317,N_2258,N_2298);
and U2318 (N_2318,N_2244,N_2227);
nor U2319 (N_2319,N_2277,N_2264);
or U2320 (N_2320,N_2257,N_2249);
nor U2321 (N_2321,N_2239,N_2279);
xor U2322 (N_2322,N_2252,N_2212);
and U2323 (N_2323,N_2299,N_2207);
or U2324 (N_2324,N_2284,N_2206);
nor U2325 (N_2325,N_2273,N_2291);
nor U2326 (N_2326,N_2217,N_2268);
nand U2327 (N_2327,N_2245,N_2293);
nand U2328 (N_2328,N_2271,N_2204);
and U2329 (N_2329,N_2234,N_2232);
nand U2330 (N_2330,N_2248,N_2202);
and U2331 (N_2331,N_2213,N_2262);
nand U2332 (N_2332,N_2228,N_2218);
nor U2333 (N_2333,N_2237,N_2255);
nand U2334 (N_2334,N_2286,N_2209);
nand U2335 (N_2335,N_2238,N_2214);
nor U2336 (N_2336,N_2297,N_2223);
and U2337 (N_2337,N_2221,N_2280);
and U2338 (N_2338,N_2231,N_2208);
or U2339 (N_2339,N_2236,N_2282);
and U2340 (N_2340,N_2267,N_2242);
or U2341 (N_2341,N_2261,N_2270);
nand U2342 (N_2342,N_2266,N_2205);
and U2343 (N_2343,N_2240,N_2230);
and U2344 (N_2344,N_2200,N_2225);
or U2345 (N_2345,N_2254,N_2292);
or U2346 (N_2346,N_2215,N_2278);
nand U2347 (N_2347,N_2246,N_2226);
or U2348 (N_2348,N_2253,N_2295);
and U2349 (N_2349,N_2216,N_2263);
nor U2350 (N_2350,N_2216,N_2283);
or U2351 (N_2351,N_2298,N_2288);
or U2352 (N_2352,N_2254,N_2256);
and U2353 (N_2353,N_2236,N_2240);
and U2354 (N_2354,N_2288,N_2225);
nand U2355 (N_2355,N_2253,N_2240);
and U2356 (N_2356,N_2273,N_2261);
and U2357 (N_2357,N_2264,N_2251);
nor U2358 (N_2358,N_2275,N_2208);
nand U2359 (N_2359,N_2263,N_2218);
or U2360 (N_2360,N_2204,N_2284);
nand U2361 (N_2361,N_2268,N_2270);
nand U2362 (N_2362,N_2280,N_2204);
nand U2363 (N_2363,N_2228,N_2274);
and U2364 (N_2364,N_2293,N_2216);
nand U2365 (N_2365,N_2237,N_2240);
or U2366 (N_2366,N_2212,N_2208);
or U2367 (N_2367,N_2209,N_2292);
and U2368 (N_2368,N_2206,N_2207);
and U2369 (N_2369,N_2228,N_2249);
nor U2370 (N_2370,N_2284,N_2264);
nor U2371 (N_2371,N_2294,N_2238);
nand U2372 (N_2372,N_2222,N_2242);
nand U2373 (N_2373,N_2234,N_2241);
nor U2374 (N_2374,N_2222,N_2257);
nor U2375 (N_2375,N_2238,N_2259);
and U2376 (N_2376,N_2212,N_2246);
nand U2377 (N_2377,N_2230,N_2287);
and U2378 (N_2378,N_2266,N_2298);
nor U2379 (N_2379,N_2252,N_2210);
nor U2380 (N_2380,N_2230,N_2234);
and U2381 (N_2381,N_2255,N_2294);
nor U2382 (N_2382,N_2201,N_2279);
nand U2383 (N_2383,N_2249,N_2244);
and U2384 (N_2384,N_2251,N_2263);
and U2385 (N_2385,N_2251,N_2207);
nand U2386 (N_2386,N_2293,N_2233);
and U2387 (N_2387,N_2218,N_2276);
and U2388 (N_2388,N_2296,N_2238);
nand U2389 (N_2389,N_2266,N_2227);
and U2390 (N_2390,N_2271,N_2227);
nor U2391 (N_2391,N_2263,N_2259);
or U2392 (N_2392,N_2283,N_2289);
and U2393 (N_2393,N_2218,N_2280);
nor U2394 (N_2394,N_2280,N_2200);
and U2395 (N_2395,N_2213,N_2223);
nor U2396 (N_2396,N_2264,N_2213);
or U2397 (N_2397,N_2231,N_2287);
nand U2398 (N_2398,N_2204,N_2240);
nand U2399 (N_2399,N_2267,N_2236);
or U2400 (N_2400,N_2368,N_2377);
nand U2401 (N_2401,N_2342,N_2348);
nand U2402 (N_2402,N_2350,N_2365);
nand U2403 (N_2403,N_2376,N_2398);
and U2404 (N_2404,N_2354,N_2352);
and U2405 (N_2405,N_2312,N_2341);
nand U2406 (N_2406,N_2375,N_2330);
nand U2407 (N_2407,N_2382,N_2369);
nor U2408 (N_2408,N_2300,N_2310);
or U2409 (N_2409,N_2345,N_2370);
and U2410 (N_2410,N_2309,N_2379);
or U2411 (N_2411,N_2320,N_2332);
nand U2412 (N_2412,N_2339,N_2385);
or U2413 (N_2413,N_2353,N_2367);
nand U2414 (N_2414,N_2351,N_2395);
and U2415 (N_2415,N_2317,N_2337);
nor U2416 (N_2416,N_2380,N_2314);
nor U2417 (N_2417,N_2336,N_2374);
or U2418 (N_2418,N_2321,N_2335);
or U2419 (N_2419,N_2399,N_2307);
nor U2420 (N_2420,N_2366,N_2386);
and U2421 (N_2421,N_2331,N_2347);
nor U2422 (N_2422,N_2378,N_2329);
or U2423 (N_2423,N_2362,N_2396);
and U2424 (N_2424,N_2392,N_2334);
nor U2425 (N_2425,N_2394,N_2303);
or U2426 (N_2426,N_2322,N_2338);
nor U2427 (N_2427,N_2357,N_2349);
nor U2428 (N_2428,N_2390,N_2360);
or U2429 (N_2429,N_2383,N_2356);
nor U2430 (N_2430,N_2304,N_2373);
nor U2431 (N_2431,N_2371,N_2363);
nand U2432 (N_2432,N_2358,N_2308);
and U2433 (N_2433,N_2325,N_2388);
and U2434 (N_2434,N_2319,N_2324);
and U2435 (N_2435,N_2306,N_2311);
nand U2436 (N_2436,N_2346,N_2393);
or U2437 (N_2437,N_2318,N_2387);
and U2438 (N_2438,N_2359,N_2384);
nand U2439 (N_2439,N_2302,N_2361);
or U2440 (N_2440,N_2397,N_2326);
or U2441 (N_2441,N_2323,N_2391);
or U2442 (N_2442,N_2328,N_2315);
and U2443 (N_2443,N_2301,N_2340);
and U2444 (N_2444,N_2327,N_2389);
nor U2445 (N_2445,N_2305,N_2313);
nor U2446 (N_2446,N_2355,N_2364);
nand U2447 (N_2447,N_2381,N_2343);
and U2448 (N_2448,N_2372,N_2316);
and U2449 (N_2449,N_2344,N_2333);
nand U2450 (N_2450,N_2379,N_2343);
nor U2451 (N_2451,N_2387,N_2302);
or U2452 (N_2452,N_2358,N_2363);
nor U2453 (N_2453,N_2397,N_2316);
nor U2454 (N_2454,N_2317,N_2331);
nor U2455 (N_2455,N_2304,N_2364);
nand U2456 (N_2456,N_2397,N_2395);
nand U2457 (N_2457,N_2336,N_2345);
or U2458 (N_2458,N_2308,N_2372);
or U2459 (N_2459,N_2396,N_2316);
or U2460 (N_2460,N_2332,N_2368);
nor U2461 (N_2461,N_2392,N_2300);
or U2462 (N_2462,N_2371,N_2304);
nor U2463 (N_2463,N_2398,N_2305);
or U2464 (N_2464,N_2368,N_2309);
nand U2465 (N_2465,N_2347,N_2377);
nor U2466 (N_2466,N_2361,N_2316);
nand U2467 (N_2467,N_2353,N_2326);
nand U2468 (N_2468,N_2310,N_2374);
nor U2469 (N_2469,N_2360,N_2301);
or U2470 (N_2470,N_2329,N_2364);
nand U2471 (N_2471,N_2376,N_2332);
or U2472 (N_2472,N_2399,N_2377);
nor U2473 (N_2473,N_2371,N_2301);
nand U2474 (N_2474,N_2368,N_2306);
nand U2475 (N_2475,N_2339,N_2381);
and U2476 (N_2476,N_2387,N_2397);
and U2477 (N_2477,N_2354,N_2391);
or U2478 (N_2478,N_2378,N_2398);
or U2479 (N_2479,N_2366,N_2320);
nand U2480 (N_2480,N_2369,N_2334);
or U2481 (N_2481,N_2320,N_2346);
and U2482 (N_2482,N_2340,N_2345);
nand U2483 (N_2483,N_2314,N_2370);
or U2484 (N_2484,N_2327,N_2302);
nor U2485 (N_2485,N_2365,N_2361);
nand U2486 (N_2486,N_2376,N_2354);
or U2487 (N_2487,N_2305,N_2344);
nand U2488 (N_2488,N_2347,N_2329);
or U2489 (N_2489,N_2332,N_2355);
or U2490 (N_2490,N_2386,N_2336);
nand U2491 (N_2491,N_2355,N_2302);
nand U2492 (N_2492,N_2359,N_2302);
or U2493 (N_2493,N_2334,N_2309);
nor U2494 (N_2494,N_2351,N_2310);
and U2495 (N_2495,N_2343,N_2301);
nand U2496 (N_2496,N_2304,N_2306);
nand U2497 (N_2497,N_2301,N_2339);
nor U2498 (N_2498,N_2359,N_2320);
or U2499 (N_2499,N_2385,N_2354);
nor U2500 (N_2500,N_2412,N_2467);
or U2501 (N_2501,N_2468,N_2498);
nor U2502 (N_2502,N_2478,N_2481);
nand U2503 (N_2503,N_2496,N_2410);
or U2504 (N_2504,N_2408,N_2449);
and U2505 (N_2505,N_2402,N_2466);
nand U2506 (N_2506,N_2451,N_2443);
and U2507 (N_2507,N_2420,N_2457);
nor U2508 (N_2508,N_2444,N_2454);
nand U2509 (N_2509,N_2452,N_2414);
or U2510 (N_2510,N_2491,N_2484);
or U2511 (N_2511,N_2483,N_2461);
or U2512 (N_2512,N_2440,N_2470);
or U2513 (N_2513,N_2476,N_2458);
nand U2514 (N_2514,N_2431,N_2447);
nor U2515 (N_2515,N_2475,N_2494);
nand U2516 (N_2516,N_2495,N_2403);
nor U2517 (N_2517,N_2455,N_2469);
or U2518 (N_2518,N_2480,N_2499);
nor U2519 (N_2519,N_2409,N_2479);
nor U2520 (N_2520,N_2464,N_2426);
nor U2521 (N_2521,N_2487,N_2427);
nor U2522 (N_2522,N_2460,N_2419);
nand U2523 (N_2523,N_2430,N_2492);
nand U2524 (N_2524,N_2493,N_2488);
or U2525 (N_2525,N_2445,N_2400);
or U2526 (N_2526,N_2425,N_2432);
nand U2527 (N_2527,N_2456,N_2446);
xor U2528 (N_2528,N_2442,N_2474);
or U2529 (N_2529,N_2441,N_2424);
or U2530 (N_2530,N_2473,N_2407);
and U2531 (N_2531,N_2471,N_2429);
and U2532 (N_2532,N_2435,N_2489);
nand U2533 (N_2533,N_2453,N_2405);
nor U2534 (N_2534,N_2448,N_2404);
or U2535 (N_2535,N_2463,N_2477);
nor U2536 (N_2536,N_2437,N_2415);
or U2537 (N_2537,N_2459,N_2436);
or U2538 (N_2538,N_2428,N_2401);
and U2539 (N_2539,N_2497,N_2462);
nand U2540 (N_2540,N_2485,N_2450);
nand U2541 (N_2541,N_2421,N_2472);
nor U2542 (N_2542,N_2439,N_2417);
nor U2543 (N_2543,N_2438,N_2433);
nand U2544 (N_2544,N_2423,N_2482);
or U2545 (N_2545,N_2465,N_2411);
nor U2546 (N_2546,N_2406,N_2413);
or U2547 (N_2547,N_2486,N_2434);
nor U2548 (N_2548,N_2490,N_2416);
nand U2549 (N_2549,N_2422,N_2418);
or U2550 (N_2550,N_2410,N_2458);
or U2551 (N_2551,N_2423,N_2407);
and U2552 (N_2552,N_2411,N_2468);
nor U2553 (N_2553,N_2418,N_2410);
nand U2554 (N_2554,N_2427,N_2417);
nand U2555 (N_2555,N_2475,N_2451);
nor U2556 (N_2556,N_2433,N_2430);
or U2557 (N_2557,N_2448,N_2469);
xor U2558 (N_2558,N_2457,N_2410);
nand U2559 (N_2559,N_2405,N_2488);
nor U2560 (N_2560,N_2451,N_2457);
nand U2561 (N_2561,N_2468,N_2420);
nand U2562 (N_2562,N_2448,N_2457);
nand U2563 (N_2563,N_2406,N_2461);
and U2564 (N_2564,N_2416,N_2402);
or U2565 (N_2565,N_2414,N_2476);
nand U2566 (N_2566,N_2497,N_2469);
and U2567 (N_2567,N_2471,N_2496);
nor U2568 (N_2568,N_2487,N_2408);
or U2569 (N_2569,N_2419,N_2477);
and U2570 (N_2570,N_2424,N_2438);
or U2571 (N_2571,N_2406,N_2466);
nor U2572 (N_2572,N_2456,N_2451);
nand U2573 (N_2573,N_2490,N_2410);
nand U2574 (N_2574,N_2480,N_2486);
nor U2575 (N_2575,N_2427,N_2430);
nand U2576 (N_2576,N_2433,N_2465);
nor U2577 (N_2577,N_2430,N_2421);
nor U2578 (N_2578,N_2431,N_2451);
nand U2579 (N_2579,N_2487,N_2479);
or U2580 (N_2580,N_2421,N_2481);
or U2581 (N_2581,N_2452,N_2476);
nor U2582 (N_2582,N_2400,N_2401);
nor U2583 (N_2583,N_2490,N_2400);
nand U2584 (N_2584,N_2403,N_2470);
or U2585 (N_2585,N_2463,N_2456);
nand U2586 (N_2586,N_2428,N_2406);
and U2587 (N_2587,N_2465,N_2441);
nor U2588 (N_2588,N_2429,N_2464);
and U2589 (N_2589,N_2409,N_2413);
nor U2590 (N_2590,N_2485,N_2433);
xor U2591 (N_2591,N_2418,N_2463);
and U2592 (N_2592,N_2473,N_2442);
nand U2593 (N_2593,N_2436,N_2441);
or U2594 (N_2594,N_2448,N_2470);
nor U2595 (N_2595,N_2460,N_2475);
nor U2596 (N_2596,N_2477,N_2464);
nand U2597 (N_2597,N_2468,N_2430);
nand U2598 (N_2598,N_2441,N_2444);
or U2599 (N_2599,N_2408,N_2495);
or U2600 (N_2600,N_2508,N_2538);
nand U2601 (N_2601,N_2523,N_2511);
nand U2602 (N_2602,N_2548,N_2554);
or U2603 (N_2603,N_2567,N_2577);
nor U2604 (N_2604,N_2505,N_2564);
or U2605 (N_2605,N_2551,N_2581);
nor U2606 (N_2606,N_2586,N_2574);
and U2607 (N_2607,N_2562,N_2596);
nand U2608 (N_2608,N_2516,N_2582);
or U2609 (N_2609,N_2553,N_2587);
nand U2610 (N_2610,N_2509,N_2506);
xnor U2611 (N_2611,N_2552,N_2583);
nand U2612 (N_2612,N_2537,N_2503);
or U2613 (N_2613,N_2580,N_2534);
or U2614 (N_2614,N_2539,N_2535);
and U2615 (N_2615,N_2558,N_2500);
or U2616 (N_2616,N_2566,N_2502);
or U2617 (N_2617,N_2588,N_2594);
and U2618 (N_2618,N_2561,N_2532);
or U2619 (N_2619,N_2571,N_2540);
nor U2620 (N_2620,N_2578,N_2584);
and U2621 (N_2621,N_2512,N_2514);
and U2622 (N_2622,N_2569,N_2531);
nor U2623 (N_2623,N_2573,N_2542);
nand U2624 (N_2624,N_2533,N_2563);
xor U2625 (N_2625,N_2555,N_2510);
nor U2626 (N_2626,N_2520,N_2579);
xor U2627 (N_2627,N_2526,N_2515);
or U2628 (N_2628,N_2518,N_2559);
nand U2629 (N_2629,N_2591,N_2545);
and U2630 (N_2630,N_2560,N_2543);
nand U2631 (N_2631,N_2522,N_2556);
nand U2632 (N_2632,N_2524,N_2504);
or U2633 (N_2633,N_2549,N_2507);
nand U2634 (N_2634,N_2599,N_2550);
nand U2635 (N_2635,N_2570,N_2589);
nor U2636 (N_2636,N_2530,N_2585);
and U2637 (N_2637,N_2598,N_2525);
nor U2638 (N_2638,N_2519,N_2501);
or U2639 (N_2639,N_2528,N_2536);
or U2640 (N_2640,N_2517,N_2546);
and U2641 (N_2641,N_2597,N_2568);
nand U2642 (N_2642,N_2565,N_2595);
nor U2643 (N_2643,N_2529,N_2541);
nand U2644 (N_2644,N_2544,N_2547);
nand U2645 (N_2645,N_2592,N_2527);
nor U2646 (N_2646,N_2593,N_2576);
and U2647 (N_2647,N_2575,N_2557);
or U2648 (N_2648,N_2590,N_2521);
nor U2649 (N_2649,N_2572,N_2513);
nand U2650 (N_2650,N_2571,N_2531);
and U2651 (N_2651,N_2563,N_2571);
xnor U2652 (N_2652,N_2508,N_2537);
nor U2653 (N_2653,N_2588,N_2506);
nand U2654 (N_2654,N_2502,N_2536);
xor U2655 (N_2655,N_2595,N_2573);
or U2656 (N_2656,N_2563,N_2582);
nand U2657 (N_2657,N_2572,N_2510);
or U2658 (N_2658,N_2599,N_2592);
nand U2659 (N_2659,N_2551,N_2586);
nand U2660 (N_2660,N_2509,N_2569);
or U2661 (N_2661,N_2534,N_2573);
and U2662 (N_2662,N_2587,N_2508);
nand U2663 (N_2663,N_2595,N_2563);
or U2664 (N_2664,N_2582,N_2514);
nand U2665 (N_2665,N_2536,N_2592);
nor U2666 (N_2666,N_2552,N_2502);
and U2667 (N_2667,N_2523,N_2593);
or U2668 (N_2668,N_2529,N_2559);
nand U2669 (N_2669,N_2536,N_2520);
nor U2670 (N_2670,N_2550,N_2578);
nor U2671 (N_2671,N_2537,N_2561);
or U2672 (N_2672,N_2564,N_2593);
nor U2673 (N_2673,N_2569,N_2505);
and U2674 (N_2674,N_2582,N_2594);
nor U2675 (N_2675,N_2529,N_2510);
and U2676 (N_2676,N_2534,N_2589);
xnor U2677 (N_2677,N_2503,N_2546);
nand U2678 (N_2678,N_2556,N_2502);
or U2679 (N_2679,N_2575,N_2505);
nor U2680 (N_2680,N_2537,N_2527);
nand U2681 (N_2681,N_2550,N_2524);
or U2682 (N_2682,N_2540,N_2580);
nand U2683 (N_2683,N_2550,N_2548);
or U2684 (N_2684,N_2500,N_2501);
nor U2685 (N_2685,N_2519,N_2522);
nor U2686 (N_2686,N_2556,N_2500);
nor U2687 (N_2687,N_2584,N_2523);
or U2688 (N_2688,N_2544,N_2527);
nor U2689 (N_2689,N_2585,N_2511);
xor U2690 (N_2690,N_2505,N_2592);
nor U2691 (N_2691,N_2553,N_2513);
xor U2692 (N_2692,N_2519,N_2521);
nand U2693 (N_2693,N_2506,N_2586);
or U2694 (N_2694,N_2575,N_2501);
or U2695 (N_2695,N_2575,N_2526);
and U2696 (N_2696,N_2505,N_2528);
xor U2697 (N_2697,N_2596,N_2520);
and U2698 (N_2698,N_2550,N_2596);
and U2699 (N_2699,N_2500,N_2591);
and U2700 (N_2700,N_2660,N_2688);
nor U2701 (N_2701,N_2613,N_2615);
or U2702 (N_2702,N_2669,N_2639);
and U2703 (N_2703,N_2627,N_2637);
and U2704 (N_2704,N_2699,N_2681);
xnor U2705 (N_2705,N_2640,N_2631);
or U2706 (N_2706,N_2624,N_2674);
nand U2707 (N_2707,N_2695,N_2610);
nand U2708 (N_2708,N_2634,N_2672);
nor U2709 (N_2709,N_2632,N_2612);
nand U2710 (N_2710,N_2665,N_2630);
and U2711 (N_2711,N_2654,N_2697);
and U2712 (N_2712,N_2647,N_2641);
nand U2713 (N_2713,N_2684,N_2680);
nand U2714 (N_2714,N_2633,N_2605);
or U2715 (N_2715,N_2603,N_2608);
xor U2716 (N_2716,N_2609,N_2606);
nand U2717 (N_2717,N_2623,N_2694);
nor U2718 (N_2718,N_2677,N_2618);
and U2719 (N_2719,N_2662,N_2692);
nor U2720 (N_2720,N_2687,N_2679);
or U2721 (N_2721,N_2646,N_2670);
nand U2722 (N_2722,N_2607,N_2621);
or U2723 (N_2723,N_2696,N_2655);
nand U2724 (N_2724,N_2653,N_2622);
and U2725 (N_2725,N_2656,N_2626);
and U2726 (N_2726,N_2651,N_2658);
and U2727 (N_2727,N_2676,N_2635);
nand U2728 (N_2728,N_2685,N_2657);
nor U2729 (N_2729,N_2649,N_2682);
nand U2730 (N_2730,N_2650,N_2645);
and U2731 (N_2731,N_2625,N_2661);
nor U2732 (N_2732,N_2617,N_2601);
or U2733 (N_2733,N_2698,N_2693);
nand U2734 (N_2734,N_2690,N_2604);
or U2735 (N_2735,N_2671,N_2648);
and U2736 (N_2736,N_2666,N_2636);
or U2737 (N_2737,N_2600,N_2619);
and U2738 (N_2738,N_2652,N_2611);
nor U2739 (N_2739,N_2629,N_2659);
or U2740 (N_2740,N_2683,N_2664);
nor U2741 (N_2741,N_2663,N_2675);
and U2742 (N_2742,N_2602,N_2673);
and U2743 (N_2743,N_2620,N_2616);
nor U2744 (N_2744,N_2642,N_2628);
nor U2745 (N_2745,N_2689,N_2678);
nor U2746 (N_2746,N_2644,N_2614);
and U2747 (N_2747,N_2668,N_2638);
nor U2748 (N_2748,N_2667,N_2643);
and U2749 (N_2749,N_2691,N_2686);
nor U2750 (N_2750,N_2690,N_2622);
or U2751 (N_2751,N_2692,N_2666);
nor U2752 (N_2752,N_2600,N_2634);
nor U2753 (N_2753,N_2695,N_2671);
and U2754 (N_2754,N_2678,N_2621);
nand U2755 (N_2755,N_2649,N_2606);
nor U2756 (N_2756,N_2645,N_2648);
nand U2757 (N_2757,N_2636,N_2615);
or U2758 (N_2758,N_2658,N_2647);
nand U2759 (N_2759,N_2684,N_2622);
or U2760 (N_2760,N_2601,N_2655);
and U2761 (N_2761,N_2635,N_2631);
nand U2762 (N_2762,N_2620,N_2606);
and U2763 (N_2763,N_2617,N_2606);
and U2764 (N_2764,N_2674,N_2677);
nor U2765 (N_2765,N_2649,N_2620);
or U2766 (N_2766,N_2620,N_2605);
nor U2767 (N_2767,N_2652,N_2632);
nand U2768 (N_2768,N_2686,N_2606);
nand U2769 (N_2769,N_2631,N_2618);
or U2770 (N_2770,N_2630,N_2632);
or U2771 (N_2771,N_2640,N_2609);
nor U2772 (N_2772,N_2695,N_2651);
nand U2773 (N_2773,N_2603,N_2678);
nand U2774 (N_2774,N_2696,N_2671);
nand U2775 (N_2775,N_2628,N_2654);
or U2776 (N_2776,N_2698,N_2682);
or U2777 (N_2777,N_2636,N_2627);
nand U2778 (N_2778,N_2615,N_2627);
and U2779 (N_2779,N_2640,N_2647);
nand U2780 (N_2780,N_2600,N_2613);
or U2781 (N_2781,N_2669,N_2601);
xnor U2782 (N_2782,N_2626,N_2697);
nand U2783 (N_2783,N_2666,N_2680);
or U2784 (N_2784,N_2640,N_2674);
or U2785 (N_2785,N_2648,N_2649);
nand U2786 (N_2786,N_2662,N_2603);
nor U2787 (N_2787,N_2664,N_2648);
nand U2788 (N_2788,N_2629,N_2678);
nor U2789 (N_2789,N_2664,N_2695);
or U2790 (N_2790,N_2655,N_2677);
nand U2791 (N_2791,N_2671,N_2666);
nand U2792 (N_2792,N_2632,N_2640);
and U2793 (N_2793,N_2683,N_2684);
or U2794 (N_2794,N_2612,N_2670);
nor U2795 (N_2795,N_2618,N_2675);
nor U2796 (N_2796,N_2656,N_2614);
and U2797 (N_2797,N_2632,N_2613);
and U2798 (N_2798,N_2644,N_2613);
nand U2799 (N_2799,N_2657,N_2655);
nor U2800 (N_2800,N_2769,N_2762);
nor U2801 (N_2801,N_2776,N_2714);
or U2802 (N_2802,N_2711,N_2790);
nor U2803 (N_2803,N_2728,N_2716);
nor U2804 (N_2804,N_2747,N_2704);
nor U2805 (N_2805,N_2787,N_2737);
or U2806 (N_2806,N_2763,N_2715);
nand U2807 (N_2807,N_2785,N_2792);
nand U2808 (N_2808,N_2779,N_2721);
nand U2809 (N_2809,N_2734,N_2745);
or U2810 (N_2810,N_2700,N_2774);
and U2811 (N_2811,N_2794,N_2783);
nand U2812 (N_2812,N_2732,N_2718);
or U2813 (N_2813,N_2731,N_2736);
xor U2814 (N_2814,N_2772,N_2723);
nand U2815 (N_2815,N_2740,N_2744);
or U2816 (N_2816,N_2735,N_2764);
and U2817 (N_2817,N_2777,N_2749);
and U2818 (N_2818,N_2786,N_2742);
nor U2819 (N_2819,N_2722,N_2738);
xnor U2820 (N_2820,N_2720,N_2708);
and U2821 (N_2821,N_2754,N_2767);
nor U2822 (N_2822,N_2788,N_2756);
xor U2823 (N_2823,N_2701,N_2705);
or U2824 (N_2824,N_2770,N_2725);
nand U2825 (N_2825,N_2797,N_2778);
xnor U2826 (N_2826,N_2741,N_2739);
and U2827 (N_2827,N_2768,N_2765);
and U2828 (N_2828,N_2771,N_2773);
nand U2829 (N_2829,N_2727,N_2793);
and U2830 (N_2830,N_2724,N_2706);
or U2831 (N_2831,N_2702,N_2746);
nand U2832 (N_2832,N_2748,N_2766);
or U2833 (N_2833,N_2759,N_2795);
nor U2834 (N_2834,N_2789,N_2750);
or U2835 (N_2835,N_2781,N_2757);
nor U2836 (N_2836,N_2707,N_2730);
or U2837 (N_2837,N_2761,N_2775);
or U2838 (N_2838,N_2799,N_2791);
or U2839 (N_2839,N_2726,N_2758);
nand U2840 (N_2840,N_2760,N_2796);
nand U2841 (N_2841,N_2751,N_2717);
nand U2842 (N_2842,N_2712,N_2782);
nor U2843 (N_2843,N_2713,N_2733);
nor U2844 (N_2844,N_2729,N_2709);
and U2845 (N_2845,N_2710,N_2784);
nor U2846 (N_2846,N_2780,N_2703);
nand U2847 (N_2847,N_2719,N_2743);
nand U2848 (N_2848,N_2798,N_2753);
and U2849 (N_2849,N_2752,N_2755);
and U2850 (N_2850,N_2746,N_2733);
or U2851 (N_2851,N_2792,N_2765);
nor U2852 (N_2852,N_2798,N_2732);
nand U2853 (N_2853,N_2720,N_2779);
xor U2854 (N_2854,N_2775,N_2718);
and U2855 (N_2855,N_2741,N_2784);
nand U2856 (N_2856,N_2785,N_2715);
and U2857 (N_2857,N_2792,N_2752);
and U2858 (N_2858,N_2780,N_2791);
nand U2859 (N_2859,N_2797,N_2727);
and U2860 (N_2860,N_2740,N_2784);
nor U2861 (N_2861,N_2761,N_2759);
xor U2862 (N_2862,N_2751,N_2766);
xor U2863 (N_2863,N_2760,N_2743);
and U2864 (N_2864,N_2798,N_2797);
or U2865 (N_2865,N_2796,N_2712);
nand U2866 (N_2866,N_2790,N_2726);
nand U2867 (N_2867,N_2716,N_2747);
nor U2868 (N_2868,N_2710,N_2779);
nor U2869 (N_2869,N_2728,N_2701);
nor U2870 (N_2870,N_2782,N_2796);
nor U2871 (N_2871,N_2745,N_2705);
nor U2872 (N_2872,N_2723,N_2765);
or U2873 (N_2873,N_2741,N_2743);
and U2874 (N_2874,N_2752,N_2729);
or U2875 (N_2875,N_2787,N_2774);
and U2876 (N_2876,N_2717,N_2759);
xor U2877 (N_2877,N_2763,N_2778);
and U2878 (N_2878,N_2763,N_2734);
or U2879 (N_2879,N_2779,N_2775);
nor U2880 (N_2880,N_2732,N_2728);
or U2881 (N_2881,N_2727,N_2730);
and U2882 (N_2882,N_2731,N_2734);
nand U2883 (N_2883,N_2732,N_2715);
nand U2884 (N_2884,N_2756,N_2742);
and U2885 (N_2885,N_2779,N_2713);
nor U2886 (N_2886,N_2766,N_2700);
nor U2887 (N_2887,N_2736,N_2755);
and U2888 (N_2888,N_2773,N_2739);
nor U2889 (N_2889,N_2762,N_2799);
nand U2890 (N_2890,N_2789,N_2738);
nor U2891 (N_2891,N_2776,N_2764);
or U2892 (N_2892,N_2769,N_2784);
nor U2893 (N_2893,N_2772,N_2795);
nor U2894 (N_2894,N_2730,N_2700);
or U2895 (N_2895,N_2768,N_2721);
and U2896 (N_2896,N_2796,N_2769);
and U2897 (N_2897,N_2785,N_2724);
nand U2898 (N_2898,N_2798,N_2771);
and U2899 (N_2899,N_2719,N_2796);
nand U2900 (N_2900,N_2896,N_2885);
nand U2901 (N_2901,N_2859,N_2814);
nor U2902 (N_2902,N_2887,N_2879);
and U2903 (N_2903,N_2881,N_2876);
and U2904 (N_2904,N_2833,N_2869);
and U2905 (N_2905,N_2823,N_2874);
xor U2906 (N_2906,N_2880,N_2839);
or U2907 (N_2907,N_2840,N_2865);
and U2908 (N_2908,N_2849,N_2845);
and U2909 (N_2909,N_2808,N_2861);
or U2910 (N_2910,N_2806,N_2851);
nand U2911 (N_2911,N_2888,N_2801);
and U2912 (N_2912,N_2877,N_2830);
nand U2913 (N_2913,N_2847,N_2807);
xor U2914 (N_2914,N_2875,N_2821);
nor U2915 (N_2915,N_2815,N_2809);
nor U2916 (N_2916,N_2856,N_2802);
or U2917 (N_2917,N_2884,N_2810);
or U2918 (N_2918,N_2812,N_2813);
nor U2919 (N_2919,N_2844,N_2852);
nand U2920 (N_2920,N_2837,N_2853);
xnor U2921 (N_2921,N_2834,N_2832);
nor U2922 (N_2922,N_2886,N_2873);
xor U2923 (N_2923,N_2890,N_2824);
nor U2924 (N_2924,N_2811,N_2829);
nand U2925 (N_2925,N_2848,N_2835);
nor U2926 (N_2926,N_2846,N_2866);
or U2927 (N_2927,N_2838,N_2842);
nor U2928 (N_2928,N_2891,N_2855);
and U2929 (N_2929,N_2892,N_2820);
and U2930 (N_2930,N_2863,N_2867);
nor U2931 (N_2931,N_2858,N_2827);
nor U2932 (N_2932,N_2872,N_2898);
or U2933 (N_2933,N_2831,N_2800);
and U2934 (N_2934,N_2816,N_2857);
nor U2935 (N_2935,N_2878,N_2819);
nor U2936 (N_2936,N_2818,N_2894);
or U2937 (N_2937,N_2862,N_2843);
nor U2938 (N_2938,N_2899,N_2854);
nor U2939 (N_2939,N_2805,N_2870);
nor U2940 (N_2940,N_2883,N_2897);
and U2941 (N_2941,N_2826,N_2803);
or U2942 (N_2942,N_2895,N_2825);
or U2943 (N_2943,N_2822,N_2889);
and U2944 (N_2944,N_2828,N_2882);
nand U2945 (N_2945,N_2817,N_2868);
nand U2946 (N_2946,N_2871,N_2860);
nor U2947 (N_2947,N_2864,N_2841);
nand U2948 (N_2948,N_2804,N_2893);
nand U2949 (N_2949,N_2850,N_2836);
xor U2950 (N_2950,N_2837,N_2881);
and U2951 (N_2951,N_2860,N_2823);
nand U2952 (N_2952,N_2877,N_2849);
nor U2953 (N_2953,N_2880,N_2831);
nor U2954 (N_2954,N_2898,N_2854);
nand U2955 (N_2955,N_2840,N_2842);
or U2956 (N_2956,N_2823,N_2815);
or U2957 (N_2957,N_2812,N_2833);
and U2958 (N_2958,N_2889,N_2809);
or U2959 (N_2959,N_2833,N_2803);
and U2960 (N_2960,N_2833,N_2896);
nor U2961 (N_2961,N_2815,N_2875);
nor U2962 (N_2962,N_2848,N_2880);
nand U2963 (N_2963,N_2842,N_2889);
and U2964 (N_2964,N_2884,N_2813);
and U2965 (N_2965,N_2882,N_2829);
nand U2966 (N_2966,N_2898,N_2850);
nand U2967 (N_2967,N_2851,N_2831);
nand U2968 (N_2968,N_2831,N_2829);
or U2969 (N_2969,N_2886,N_2838);
or U2970 (N_2970,N_2873,N_2891);
xor U2971 (N_2971,N_2863,N_2814);
nor U2972 (N_2972,N_2859,N_2807);
nor U2973 (N_2973,N_2801,N_2821);
xor U2974 (N_2974,N_2883,N_2877);
nand U2975 (N_2975,N_2818,N_2848);
nor U2976 (N_2976,N_2812,N_2808);
and U2977 (N_2977,N_2823,N_2812);
or U2978 (N_2978,N_2890,N_2823);
nand U2979 (N_2979,N_2823,N_2887);
nand U2980 (N_2980,N_2858,N_2873);
xor U2981 (N_2981,N_2832,N_2858);
or U2982 (N_2982,N_2856,N_2843);
nor U2983 (N_2983,N_2892,N_2875);
nor U2984 (N_2984,N_2844,N_2827);
nor U2985 (N_2985,N_2834,N_2871);
nor U2986 (N_2986,N_2820,N_2890);
and U2987 (N_2987,N_2844,N_2873);
nor U2988 (N_2988,N_2812,N_2885);
and U2989 (N_2989,N_2818,N_2889);
and U2990 (N_2990,N_2883,N_2882);
nand U2991 (N_2991,N_2838,N_2885);
nor U2992 (N_2992,N_2813,N_2878);
nor U2993 (N_2993,N_2884,N_2895);
and U2994 (N_2994,N_2868,N_2860);
nand U2995 (N_2995,N_2860,N_2827);
nand U2996 (N_2996,N_2894,N_2825);
or U2997 (N_2997,N_2837,N_2843);
or U2998 (N_2998,N_2895,N_2816);
or U2999 (N_2999,N_2836,N_2860);
and UO_0 (O_0,N_2903,N_2991);
nor UO_1 (O_1,N_2938,N_2916);
or UO_2 (O_2,N_2912,N_2910);
nand UO_3 (O_3,N_2974,N_2981);
nand UO_4 (O_4,N_2967,N_2932);
nor UO_5 (O_5,N_2906,N_2923);
and UO_6 (O_6,N_2951,N_2914);
and UO_7 (O_7,N_2950,N_2953);
nand UO_8 (O_8,N_2986,N_2922);
nand UO_9 (O_9,N_2934,N_2901);
or UO_10 (O_10,N_2965,N_2966);
nand UO_11 (O_11,N_2969,N_2918);
nand UO_12 (O_12,N_2907,N_2957);
nor UO_13 (O_13,N_2982,N_2988);
nor UO_14 (O_14,N_2952,N_2977);
nand UO_15 (O_15,N_2905,N_2954);
nand UO_16 (O_16,N_2931,N_2921);
and UO_17 (O_17,N_2917,N_2930);
and UO_18 (O_18,N_2996,N_2998);
nor UO_19 (O_19,N_2971,N_2978);
nand UO_20 (O_20,N_2999,N_2961);
nand UO_21 (O_21,N_2929,N_2911);
nand UO_22 (O_22,N_2983,N_2924);
and UO_23 (O_23,N_2925,N_2968);
and UO_24 (O_24,N_2979,N_2990);
or UO_25 (O_25,N_2959,N_2956);
nor UO_26 (O_26,N_2993,N_2972);
nand UO_27 (O_27,N_2928,N_2975);
or UO_28 (O_28,N_2985,N_2955);
and UO_29 (O_29,N_2963,N_2970);
nand UO_30 (O_30,N_2927,N_2958);
and UO_31 (O_31,N_2937,N_2936);
and UO_32 (O_32,N_2989,N_2992);
or UO_33 (O_33,N_2941,N_2946);
and UO_34 (O_34,N_2909,N_2915);
nand UO_35 (O_35,N_2976,N_2904);
nand UO_36 (O_36,N_2995,N_2943);
nor UO_37 (O_37,N_2997,N_2949);
nor UO_38 (O_38,N_2944,N_2973);
or UO_39 (O_39,N_2908,N_2902);
and UO_40 (O_40,N_2940,N_2962);
and UO_41 (O_41,N_2964,N_2948);
or UO_42 (O_42,N_2913,N_2980);
or UO_43 (O_43,N_2900,N_2939);
xnor UO_44 (O_44,N_2984,N_2920);
and UO_45 (O_45,N_2945,N_2935);
or UO_46 (O_46,N_2960,N_2926);
nor UO_47 (O_47,N_2942,N_2933);
and UO_48 (O_48,N_2994,N_2947);
nand UO_49 (O_49,N_2919,N_2987);
nor UO_50 (O_50,N_2944,N_2956);
nor UO_51 (O_51,N_2986,N_2933);
nor UO_52 (O_52,N_2922,N_2972);
nand UO_53 (O_53,N_2943,N_2961);
nand UO_54 (O_54,N_2975,N_2964);
nand UO_55 (O_55,N_2927,N_2939);
or UO_56 (O_56,N_2904,N_2988);
nand UO_57 (O_57,N_2995,N_2914);
nor UO_58 (O_58,N_2942,N_2906);
nand UO_59 (O_59,N_2979,N_2982);
nor UO_60 (O_60,N_2950,N_2992);
or UO_61 (O_61,N_2989,N_2985);
or UO_62 (O_62,N_2991,N_2985);
and UO_63 (O_63,N_2911,N_2904);
or UO_64 (O_64,N_2977,N_2940);
or UO_65 (O_65,N_2991,N_2958);
nor UO_66 (O_66,N_2953,N_2931);
nand UO_67 (O_67,N_2978,N_2956);
nor UO_68 (O_68,N_2946,N_2953);
nor UO_69 (O_69,N_2905,N_2969);
or UO_70 (O_70,N_2978,N_2912);
or UO_71 (O_71,N_2921,N_2980);
nand UO_72 (O_72,N_2939,N_2932);
nor UO_73 (O_73,N_2910,N_2932);
and UO_74 (O_74,N_2956,N_2967);
and UO_75 (O_75,N_2984,N_2974);
nor UO_76 (O_76,N_2957,N_2917);
and UO_77 (O_77,N_2964,N_2925);
nand UO_78 (O_78,N_2981,N_2915);
or UO_79 (O_79,N_2994,N_2970);
and UO_80 (O_80,N_2996,N_2979);
nor UO_81 (O_81,N_2929,N_2955);
nand UO_82 (O_82,N_2961,N_2903);
nor UO_83 (O_83,N_2913,N_2925);
or UO_84 (O_84,N_2929,N_2990);
or UO_85 (O_85,N_2967,N_2996);
and UO_86 (O_86,N_2946,N_2951);
nand UO_87 (O_87,N_2992,N_2966);
and UO_88 (O_88,N_2958,N_2942);
nand UO_89 (O_89,N_2946,N_2966);
or UO_90 (O_90,N_2941,N_2928);
or UO_91 (O_91,N_2958,N_2957);
nand UO_92 (O_92,N_2939,N_2907);
nand UO_93 (O_93,N_2952,N_2945);
nor UO_94 (O_94,N_2994,N_2996);
and UO_95 (O_95,N_2998,N_2910);
nor UO_96 (O_96,N_2938,N_2937);
xnor UO_97 (O_97,N_2952,N_2921);
nor UO_98 (O_98,N_2907,N_2963);
and UO_99 (O_99,N_2904,N_2951);
or UO_100 (O_100,N_2991,N_2901);
and UO_101 (O_101,N_2905,N_2943);
and UO_102 (O_102,N_2909,N_2944);
nand UO_103 (O_103,N_2934,N_2914);
nand UO_104 (O_104,N_2989,N_2914);
and UO_105 (O_105,N_2928,N_2920);
nand UO_106 (O_106,N_2992,N_2976);
nand UO_107 (O_107,N_2977,N_2994);
nand UO_108 (O_108,N_2967,N_2901);
or UO_109 (O_109,N_2978,N_2977);
or UO_110 (O_110,N_2940,N_2949);
nor UO_111 (O_111,N_2900,N_2943);
and UO_112 (O_112,N_2973,N_2966);
nand UO_113 (O_113,N_2991,N_2937);
and UO_114 (O_114,N_2937,N_2979);
nor UO_115 (O_115,N_2926,N_2980);
nor UO_116 (O_116,N_2966,N_2980);
nor UO_117 (O_117,N_2969,N_2973);
nand UO_118 (O_118,N_2993,N_2925);
or UO_119 (O_119,N_2969,N_2947);
and UO_120 (O_120,N_2928,N_2915);
and UO_121 (O_121,N_2933,N_2947);
nor UO_122 (O_122,N_2990,N_2977);
and UO_123 (O_123,N_2912,N_2940);
nor UO_124 (O_124,N_2988,N_2943);
nor UO_125 (O_125,N_2999,N_2926);
nor UO_126 (O_126,N_2969,N_2903);
and UO_127 (O_127,N_2980,N_2911);
nand UO_128 (O_128,N_2941,N_2940);
nor UO_129 (O_129,N_2986,N_2910);
nor UO_130 (O_130,N_2973,N_2922);
nor UO_131 (O_131,N_2980,N_2965);
and UO_132 (O_132,N_2902,N_2937);
nor UO_133 (O_133,N_2905,N_2933);
or UO_134 (O_134,N_2939,N_2977);
nand UO_135 (O_135,N_2907,N_2978);
nor UO_136 (O_136,N_2989,N_2978);
or UO_137 (O_137,N_2949,N_2912);
nand UO_138 (O_138,N_2959,N_2979);
nand UO_139 (O_139,N_2903,N_2910);
or UO_140 (O_140,N_2948,N_2914);
or UO_141 (O_141,N_2916,N_2965);
or UO_142 (O_142,N_2938,N_2906);
xnor UO_143 (O_143,N_2908,N_2996);
or UO_144 (O_144,N_2954,N_2998);
nor UO_145 (O_145,N_2951,N_2926);
nand UO_146 (O_146,N_2911,N_2900);
and UO_147 (O_147,N_2906,N_2949);
or UO_148 (O_148,N_2999,N_2907);
nor UO_149 (O_149,N_2994,N_2910);
and UO_150 (O_150,N_2976,N_2958);
and UO_151 (O_151,N_2960,N_2969);
nor UO_152 (O_152,N_2912,N_2914);
and UO_153 (O_153,N_2975,N_2920);
nor UO_154 (O_154,N_2945,N_2913);
nand UO_155 (O_155,N_2998,N_2975);
or UO_156 (O_156,N_2902,N_2909);
nor UO_157 (O_157,N_2901,N_2904);
nand UO_158 (O_158,N_2935,N_2917);
nor UO_159 (O_159,N_2964,N_2941);
nor UO_160 (O_160,N_2986,N_2944);
nor UO_161 (O_161,N_2988,N_2942);
nor UO_162 (O_162,N_2996,N_2923);
nand UO_163 (O_163,N_2988,N_2900);
or UO_164 (O_164,N_2977,N_2965);
or UO_165 (O_165,N_2995,N_2973);
or UO_166 (O_166,N_2999,N_2983);
nor UO_167 (O_167,N_2960,N_2999);
nor UO_168 (O_168,N_2905,N_2906);
and UO_169 (O_169,N_2996,N_2901);
nand UO_170 (O_170,N_2964,N_2960);
nand UO_171 (O_171,N_2924,N_2964);
or UO_172 (O_172,N_2986,N_2968);
or UO_173 (O_173,N_2953,N_2997);
nor UO_174 (O_174,N_2956,N_2941);
nor UO_175 (O_175,N_2912,N_2929);
or UO_176 (O_176,N_2927,N_2916);
and UO_177 (O_177,N_2907,N_2943);
and UO_178 (O_178,N_2906,N_2916);
nor UO_179 (O_179,N_2958,N_2928);
nand UO_180 (O_180,N_2953,N_2907);
nand UO_181 (O_181,N_2913,N_2956);
nor UO_182 (O_182,N_2991,N_2993);
or UO_183 (O_183,N_2917,N_2906);
and UO_184 (O_184,N_2911,N_2935);
and UO_185 (O_185,N_2962,N_2979);
nor UO_186 (O_186,N_2977,N_2999);
and UO_187 (O_187,N_2991,N_2908);
nand UO_188 (O_188,N_2925,N_2916);
nand UO_189 (O_189,N_2930,N_2991);
nand UO_190 (O_190,N_2921,N_2981);
nor UO_191 (O_191,N_2954,N_2935);
and UO_192 (O_192,N_2939,N_2904);
nand UO_193 (O_193,N_2908,N_2926);
or UO_194 (O_194,N_2935,N_2957);
or UO_195 (O_195,N_2908,N_2995);
nand UO_196 (O_196,N_2994,N_2998);
nor UO_197 (O_197,N_2924,N_2987);
and UO_198 (O_198,N_2907,N_2977);
nand UO_199 (O_199,N_2937,N_2960);
or UO_200 (O_200,N_2941,N_2939);
nand UO_201 (O_201,N_2912,N_2969);
and UO_202 (O_202,N_2983,N_2927);
xnor UO_203 (O_203,N_2907,N_2987);
nand UO_204 (O_204,N_2953,N_2967);
or UO_205 (O_205,N_2980,N_2936);
or UO_206 (O_206,N_2952,N_2981);
and UO_207 (O_207,N_2909,N_2985);
or UO_208 (O_208,N_2926,N_2963);
and UO_209 (O_209,N_2930,N_2952);
or UO_210 (O_210,N_2954,N_2980);
nand UO_211 (O_211,N_2975,N_2934);
nand UO_212 (O_212,N_2985,N_2936);
nor UO_213 (O_213,N_2999,N_2947);
nand UO_214 (O_214,N_2905,N_2919);
or UO_215 (O_215,N_2972,N_2958);
xor UO_216 (O_216,N_2970,N_2912);
or UO_217 (O_217,N_2908,N_2907);
or UO_218 (O_218,N_2914,N_2910);
xor UO_219 (O_219,N_2947,N_2975);
nor UO_220 (O_220,N_2962,N_2956);
nand UO_221 (O_221,N_2915,N_2962);
or UO_222 (O_222,N_2996,N_2942);
nor UO_223 (O_223,N_2946,N_2931);
or UO_224 (O_224,N_2964,N_2978);
and UO_225 (O_225,N_2940,N_2974);
and UO_226 (O_226,N_2915,N_2912);
and UO_227 (O_227,N_2923,N_2900);
nand UO_228 (O_228,N_2973,N_2926);
nand UO_229 (O_229,N_2988,N_2902);
and UO_230 (O_230,N_2933,N_2952);
nand UO_231 (O_231,N_2993,N_2970);
nand UO_232 (O_232,N_2904,N_2931);
nand UO_233 (O_233,N_2917,N_2988);
and UO_234 (O_234,N_2992,N_2949);
nor UO_235 (O_235,N_2927,N_2975);
and UO_236 (O_236,N_2957,N_2967);
or UO_237 (O_237,N_2975,N_2944);
nor UO_238 (O_238,N_2996,N_2919);
nor UO_239 (O_239,N_2989,N_2991);
or UO_240 (O_240,N_2954,N_2937);
nor UO_241 (O_241,N_2935,N_2915);
nand UO_242 (O_242,N_2915,N_2951);
nor UO_243 (O_243,N_2992,N_2973);
or UO_244 (O_244,N_2928,N_2901);
nand UO_245 (O_245,N_2918,N_2973);
nor UO_246 (O_246,N_2972,N_2971);
nand UO_247 (O_247,N_2947,N_2944);
or UO_248 (O_248,N_2938,N_2977);
nand UO_249 (O_249,N_2915,N_2910);
or UO_250 (O_250,N_2940,N_2905);
and UO_251 (O_251,N_2920,N_2982);
xnor UO_252 (O_252,N_2937,N_2949);
or UO_253 (O_253,N_2966,N_2972);
nor UO_254 (O_254,N_2952,N_2910);
nand UO_255 (O_255,N_2999,N_2927);
or UO_256 (O_256,N_2921,N_2950);
and UO_257 (O_257,N_2922,N_2952);
or UO_258 (O_258,N_2906,N_2933);
and UO_259 (O_259,N_2977,N_2948);
nor UO_260 (O_260,N_2918,N_2949);
nand UO_261 (O_261,N_2945,N_2973);
and UO_262 (O_262,N_2905,N_2973);
or UO_263 (O_263,N_2904,N_2989);
or UO_264 (O_264,N_2923,N_2955);
nor UO_265 (O_265,N_2924,N_2916);
nor UO_266 (O_266,N_2943,N_2918);
or UO_267 (O_267,N_2969,N_2966);
and UO_268 (O_268,N_2996,N_2970);
nand UO_269 (O_269,N_2910,N_2935);
nor UO_270 (O_270,N_2910,N_2929);
and UO_271 (O_271,N_2921,N_2979);
or UO_272 (O_272,N_2905,N_2925);
nand UO_273 (O_273,N_2908,N_2999);
nand UO_274 (O_274,N_2984,N_2994);
or UO_275 (O_275,N_2979,N_2900);
nand UO_276 (O_276,N_2984,N_2979);
and UO_277 (O_277,N_2932,N_2946);
nand UO_278 (O_278,N_2999,N_2920);
nand UO_279 (O_279,N_2957,N_2937);
or UO_280 (O_280,N_2970,N_2937);
nor UO_281 (O_281,N_2999,N_2911);
nand UO_282 (O_282,N_2958,N_2929);
nor UO_283 (O_283,N_2911,N_2905);
or UO_284 (O_284,N_2923,N_2915);
nor UO_285 (O_285,N_2943,N_2997);
nand UO_286 (O_286,N_2975,N_2950);
nor UO_287 (O_287,N_2938,N_2945);
nand UO_288 (O_288,N_2934,N_2968);
nor UO_289 (O_289,N_2920,N_2964);
or UO_290 (O_290,N_2907,N_2930);
or UO_291 (O_291,N_2915,N_2940);
or UO_292 (O_292,N_2913,N_2976);
xnor UO_293 (O_293,N_2933,N_2935);
nor UO_294 (O_294,N_2907,N_2986);
nor UO_295 (O_295,N_2921,N_2925);
or UO_296 (O_296,N_2960,N_2976);
nor UO_297 (O_297,N_2963,N_2964);
nor UO_298 (O_298,N_2988,N_2973);
nor UO_299 (O_299,N_2984,N_2971);
and UO_300 (O_300,N_2974,N_2957);
or UO_301 (O_301,N_2900,N_2931);
or UO_302 (O_302,N_2945,N_2993);
nand UO_303 (O_303,N_2921,N_2901);
nand UO_304 (O_304,N_2931,N_2975);
nand UO_305 (O_305,N_2906,N_2991);
nor UO_306 (O_306,N_2971,N_2974);
or UO_307 (O_307,N_2980,N_2940);
or UO_308 (O_308,N_2973,N_2900);
or UO_309 (O_309,N_2959,N_2985);
or UO_310 (O_310,N_2915,N_2933);
and UO_311 (O_311,N_2933,N_2972);
nor UO_312 (O_312,N_2963,N_2901);
and UO_313 (O_313,N_2940,N_2978);
or UO_314 (O_314,N_2981,N_2922);
nor UO_315 (O_315,N_2952,N_2937);
or UO_316 (O_316,N_2917,N_2985);
nand UO_317 (O_317,N_2948,N_2902);
nand UO_318 (O_318,N_2997,N_2910);
nor UO_319 (O_319,N_2910,N_2965);
nor UO_320 (O_320,N_2931,N_2933);
nand UO_321 (O_321,N_2979,N_2931);
or UO_322 (O_322,N_2940,N_2989);
nor UO_323 (O_323,N_2954,N_2948);
or UO_324 (O_324,N_2941,N_2942);
nor UO_325 (O_325,N_2939,N_2996);
xor UO_326 (O_326,N_2928,N_2976);
and UO_327 (O_327,N_2947,N_2964);
nand UO_328 (O_328,N_2984,N_2959);
nor UO_329 (O_329,N_2988,N_2990);
or UO_330 (O_330,N_2979,N_2942);
or UO_331 (O_331,N_2970,N_2944);
and UO_332 (O_332,N_2907,N_2985);
xnor UO_333 (O_333,N_2970,N_2904);
or UO_334 (O_334,N_2952,N_2993);
nand UO_335 (O_335,N_2906,N_2948);
or UO_336 (O_336,N_2913,N_2955);
and UO_337 (O_337,N_2969,N_2965);
nor UO_338 (O_338,N_2987,N_2937);
and UO_339 (O_339,N_2935,N_2994);
or UO_340 (O_340,N_2996,N_2963);
and UO_341 (O_341,N_2913,N_2979);
or UO_342 (O_342,N_2941,N_2914);
nor UO_343 (O_343,N_2996,N_2912);
and UO_344 (O_344,N_2922,N_2901);
nand UO_345 (O_345,N_2941,N_2911);
nand UO_346 (O_346,N_2989,N_2935);
nand UO_347 (O_347,N_2986,N_2932);
or UO_348 (O_348,N_2945,N_2983);
nor UO_349 (O_349,N_2971,N_2954);
nor UO_350 (O_350,N_2917,N_2955);
nor UO_351 (O_351,N_2903,N_2994);
or UO_352 (O_352,N_2976,N_2916);
and UO_353 (O_353,N_2919,N_2962);
and UO_354 (O_354,N_2991,N_2977);
nor UO_355 (O_355,N_2905,N_2932);
and UO_356 (O_356,N_2926,N_2987);
nor UO_357 (O_357,N_2986,N_2984);
nor UO_358 (O_358,N_2963,N_2920);
or UO_359 (O_359,N_2930,N_2913);
or UO_360 (O_360,N_2985,N_2903);
nand UO_361 (O_361,N_2929,N_2918);
nand UO_362 (O_362,N_2907,N_2931);
or UO_363 (O_363,N_2925,N_2959);
and UO_364 (O_364,N_2975,N_2904);
nand UO_365 (O_365,N_2992,N_2948);
nor UO_366 (O_366,N_2910,N_2955);
and UO_367 (O_367,N_2914,N_2944);
and UO_368 (O_368,N_2967,N_2978);
or UO_369 (O_369,N_2918,N_2974);
or UO_370 (O_370,N_2900,N_2949);
or UO_371 (O_371,N_2948,N_2913);
or UO_372 (O_372,N_2988,N_2979);
and UO_373 (O_373,N_2960,N_2904);
or UO_374 (O_374,N_2967,N_2921);
nor UO_375 (O_375,N_2930,N_2921);
nor UO_376 (O_376,N_2959,N_2970);
and UO_377 (O_377,N_2980,N_2947);
nand UO_378 (O_378,N_2977,N_2909);
and UO_379 (O_379,N_2948,N_2999);
and UO_380 (O_380,N_2902,N_2997);
nor UO_381 (O_381,N_2945,N_2956);
nand UO_382 (O_382,N_2928,N_2911);
nor UO_383 (O_383,N_2967,N_2964);
or UO_384 (O_384,N_2945,N_2959);
and UO_385 (O_385,N_2973,N_2937);
nor UO_386 (O_386,N_2979,N_2947);
or UO_387 (O_387,N_2940,N_2982);
nor UO_388 (O_388,N_2999,N_2956);
and UO_389 (O_389,N_2961,N_2908);
and UO_390 (O_390,N_2994,N_2936);
or UO_391 (O_391,N_2960,N_2971);
nand UO_392 (O_392,N_2963,N_2942);
or UO_393 (O_393,N_2988,N_2911);
and UO_394 (O_394,N_2935,N_2918);
or UO_395 (O_395,N_2971,N_2938);
and UO_396 (O_396,N_2953,N_2901);
nand UO_397 (O_397,N_2957,N_2945);
nand UO_398 (O_398,N_2915,N_2979);
and UO_399 (O_399,N_2973,N_2934);
or UO_400 (O_400,N_2905,N_2963);
nor UO_401 (O_401,N_2909,N_2935);
nand UO_402 (O_402,N_2953,N_2982);
nand UO_403 (O_403,N_2901,N_2956);
or UO_404 (O_404,N_2906,N_2947);
and UO_405 (O_405,N_2911,N_2987);
nand UO_406 (O_406,N_2908,N_2934);
nor UO_407 (O_407,N_2926,N_2967);
and UO_408 (O_408,N_2960,N_2932);
or UO_409 (O_409,N_2900,N_2901);
or UO_410 (O_410,N_2917,N_2916);
or UO_411 (O_411,N_2986,N_2931);
or UO_412 (O_412,N_2947,N_2985);
or UO_413 (O_413,N_2982,N_2913);
nand UO_414 (O_414,N_2939,N_2958);
nor UO_415 (O_415,N_2989,N_2984);
nor UO_416 (O_416,N_2950,N_2907);
nand UO_417 (O_417,N_2958,N_2982);
nand UO_418 (O_418,N_2927,N_2900);
or UO_419 (O_419,N_2914,N_2965);
or UO_420 (O_420,N_2984,N_2969);
and UO_421 (O_421,N_2955,N_2947);
nand UO_422 (O_422,N_2904,N_2919);
or UO_423 (O_423,N_2923,N_2983);
and UO_424 (O_424,N_2903,N_2913);
and UO_425 (O_425,N_2918,N_2965);
and UO_426 (O_426,N_2998,N_2906);
or UO_427 (O_427,N_2974,N_2972);
and UO_428 (O_428,N_2900,N_2956);
and UO_429 (O_429,N_2913,N_2908);
nand UO_430 (O_430,N_2932,N_2981);
or UO_431 (O_431,N_2936,N_2908);
nand UO_432 (O_432,N_2952,N_2944);
nor UO_433 (O_433,N_2940,N_2953);
or UO_434 (O_434,N_2986,N_2963);
and UO_435 (O_435,N_2978,N_2973);
and UO_436 (O_436,N_2995,N_2929);
nor UO_437 (O_437,N_2986,N_2991);
nor UO_438 (O_438,N_2974,N_2992);
or UO_439 (O_439,N_2976,N_2930);
and UO_440 (O_440,N_2941,N_2910);
and UO_441 (O_441,N_2901,N_2902);
or UO_442 (O_442,N_2978,N_2929);
and UO_443 (O_443,N_2980,N_2984);
nand UO_444 (O_444,N_2906,N_2926);
and UO_445 (O_445,N_2954,N_2946);
or UO_446 (O_446,N_2936,N_2929);
nand UO_447 (O_447,N_2998,N_2985);
and UO_448 (O_448,N_2916,N_2973);
or UO_449 (O_449,N_2965,N_2981);
and UO_450 (O_450,N_2916,N_2956);
nand UO_451 (O_451,N_2931,N_2926);
xnor UO_452 (O_452,N_2939,N_2984);
nand UO_453 (O_453,N_2943,N_2902);
xnor UO_454 (O_454,N_2958,N_2945);
or UO_455 (O_455,N_2978,N_2906);
nand UO_456 (O_456,N_2927,N_2994);
and UO_457 (O_457,N_2969,N_2907);
or UO_458 (O_458,N_2975,N_2970);
and UO_459 (O_459,N_2951,N_2980);
xor UO_460 (O_460,N_2950,N_2985);
nand UO_461 (O_461,N_2967,N_2989);
nor UO_462 (O_462,N_2912,N_2966);
or UO_463 (O_463,N_2978,N_2983);
and UO_464 (O_464,N_2986,N_2926);
nand UO_465 (O_465,N_2953,N_2937);
and UO_466 (O_466,N_2951,N_2953);
and UO_467 (O_467,N_2943,N_2994);
nand UO_468 (O_468,N_2953,N_2996);
and UO_469 (O_469,N_2946,N_2921);
nand UO_470 (O_470,N_2961,N_2958);
nor UO_471 (O_471,N_2946,N_2909);
and UO_472 (O_472,N_2950,N_2973);
nand UO_473 (O_473,N_2987,N_2952);
and UO_474 (O_474,N_2950,N_2974);
xor UO_475 (O_475,N_2908,N_2981);
or UO_476 (O_476,N_2906,N_2921);
nand UO_477 (O_477,N_2978,N_2961);
and UO_478 (O_478,N_2915,N_2917);
nand UO_479 (O_479,N_2947,N_2992);
and UO_480 (O_480,N_2928,N_2973);
nand UO_481 (O_481,N_2917,N_2968);
xor UO_482 (O_482,N_2979,N_2938);
and UO_483 (O_483,N_2987,N_2906);
nor UO_484 (O_484,N_2973,N_2939);
nor UO_485 (O_485,N_2950,N_2909);
nor UO_486 (O_486,N_2945,N_2998);
nand UO_487 (O_487,N_2980,N_2982);
or UO_488 (O_488,N_2966,N_2905);
nand UO_489 (O_489,N_2960,N_2929);
and UO_490 (O_490,N_2944,N_2976);
or UO_491 (O_491,N_2973,N_2902);
and UO_492 (O_492,N_2922,N_2955);
and UO_493 (O_493,N_2916,N_2987);
nor UO_494 (O_494,N_2949,N_2976);
and UO_495 (O_495,N_2967,N_2995);
nor UO_496 (O_496,N_2924,N_2915);
or UO_497 (O_497,N_2902,N_2926);
nand UO_498 (O_498,N_2926,N_2920);
or UO_499 (O_499,N_2975,N_2905);
endmodule