module basic_1000_10000_1500_5_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_638,In_790);
nor U1 (N_1,In_92,In_923);
nor U2 (N_2,In_107,In_264);
xor U3 (N_3,In_838,In_330);
xor U4 (N_4,In_310,In_897);
and U5 (N_5,In_585,In_969);
nand U6 (N_6,In_344,In_710);
xor U7 (N_7,In_993,In_241);
and U8 (N_8,In_527,In_108);
xor U9 (N_9,In_469,In_428);
and U10 (N_10,In_178,In_89);
and U11 (N_11,In_632,In_72);
nand U12 (N_12,In_957,In_326);
nand U13 (N_13,In_780,In_801);
nor U14 (N_14,In_764,In_616);
nor U15 (N_15,In_776,In_270);
or U16 (N_16,In_866,In_892);
nor U17 (N_17,In_890,In_749);
and U18 (N_18,In_146,In_557);
and U19 (N_19,In_454,In_444);
nor U20 (N_20,In_630,In_808);
nor U21 (N_21,In_833,In_767);
nand U22 (N_22,In_839,In_799);
and U23 (N_23,In_576,In_153);
or U24 (N_24,In_949,In_111);
nand U25 (N_25,In_507,In_641);
and U26 (N_26,In_177,In_590);
xor U27 (N_27,In_371,In_735);
nand U28 (N_28,In_132,In_606);
nand U29 (N_29,In_193,In_413);
or U30 (N_30,In_901,In_137);
and U31 (N_31,In_282,In_123);
or U32 (N_32,In_968,In_587);
and U33 (N_33,In_55,In_240);
nor U34 (N_34,In_24,In_640);
or U35 (N_35,In_900,In_143);
nor U36 (N_36,In_588,In_940);
nand U37 (N_37,In_119,In_865);
nand U38 (N_38,In_490,In_386);
nor U39 (N_39,In_813,In_924);
nor U40 (N_40,In_84,In_664);
nor U41 (N_41,In_651,In_579);
or U42 (N_42,In_740,In_872);
xor U43 (N_43,In_459,In_437);
nand U44 (N_44,In_753,In_58);
nand U45 (N_45,In_429,In_921);
or U46 (N_46,In_124,In_403);
xnor U47 (N_47,In_499,In_209);
nand U48 (N_48,In_605,In_16);
and U49 (N_49,In_719,In_198);
or U50 (N_50,In_158,In_537);
xor U51 (N_51,In_811,In_955);
nor U52 (N_52,In_206,In_723);
nand U53 (N_53,In_457,In_635);
or U54 (N_54,In_136,In_360);
and U55 (N_55,In_321,In_674);
nand U56 (N_56,In_443,In_763);
and U57 (N_57,In_681,In_231);
or U58 (N_58,In_959,In_649);
nand U59 (N_59,In_477,In_699);
nand U60 (N_60,In_254,In_170);
and U61 (N_61,In_907,In_703);
and U62 (N_62,In_38,In_165);
xor U63 (N_63,In_19,In_22);
nor U64 (N_64,In_583,In_836);
nor U65 (N_65,In_526,In_73);
or U66 (N_66,In_547,In_757);
and U67 (N_67,In_601,In_953);
xor U68 (N_68,In_243,In_224);
nor U69 (N_69,In_521,In_306);
nand U70 (N_70,In_936,In_75);
nor U71 (N_71,In_709,In_743);
nor U72 (N_72,In_362,In_401);
or U73 (N_73,In_631,In_388);
nand U74 (N_74,In_37,In_602);
nor U75 (N_75,In_244,In_822);
and U76 (N_76,In_36,In_643);
nand U77 (N_77,In_302,In_104);
and U78 (N_78,In_511,In_534);
xor U79 (N_79,In_195,In_835);
nor U80 (N_80,In_440,In_773);
or U81 (N_81,In_922,In_402);
or U82 (N_82,In_524,In_201);
or U83 (N_83,In_106,In_563);
and U84 (N_84,In_468,In_338);
xnor U85 (N_85,In_626,In_329);
or U86 (N_86,In_952,In_97);
or U87 (N_87,In_384,In_196);
or U88 (N_88,In_117,In_725);
nor U89 (N_89,In_250,In_389);
xnor U90 (N_90,In_880,In_164);
or U91 (N_91,In_422,In_934);
nor U92 (N_92,In_560,In_152);
nor U93 (N_93,In_359,In_728);
nor U94 (N_94,In_174,In_120);
or U95 (N_95,In_966,In_891);
nor U96 (N_96,In_289,In_581);
and U97 (N_97,In_971,In_122);
and U98 (N_98,In_214,In_910);
or U99 (N_99,In_286,In_797);
nand U100 (N_100,In_462,In_445);
or U101 (N_101,In_70,In_491);
nor U102 (N_102,In_736,In_40);
nor U103 (N_103,In_693,In_502);
and U104 (N_104,In_669,In_809);
nand U105 (N_105,In_215,In_974);
or U106 (N_106,In_7,In_168);
nor U107 (N_107,In_915,In_567);
xnor U108 (N_108,In_991,In_297);
or U109 (N_109,In_208,In_761);
nor U110 (N_110,In_333,In_251);
or U111 (N_111,In_23,In_395);
nor U112 (N_112,In_568,In_441);
nor U113 (N_113,In_14,In_732);
nand U114 (N_114,In_972,In_139);
and U115 (N_115,In_672,In_39);
nand U116 (N_116,In_603,In_312);
nand U117 (N_117,In_538,In_467);
or U118 (N_118,In_159,In_687);
or U119 (N_119,In_979,In_160);
or U120 (N_120,In_447,In_807);
nor U121 (N_121,In_796,In_508);
and U122 (N_122,In_932,In_671);
xnor U123 (N_123,In_722,In_135);
or U124 (N_124,In_320,In_274);
nor U125 (N_125,In_665,In_791);
nand U126 (N_126,In_582,In_184);
nor U127 (N_127,In_661,In_864);
or U128 (N_128,In_950,In_81);
or U129 (N_129,In_997,In_818);
nor U130 (N_130,In_541,In_842);
and U131 (N_131,In_182,In_339);
nand U132 (N_132,In_309,In_926);
xnor U133 (N_133,In_943,In_420);
nand U134 (N_134,In_110,In_994);
and U135 (N_135,In_252,In_318);
xor U136 (N_136,In_857,In_716);
nor U137 (N_137,In_155,In_20);
nand U138 (N_138,In_460,In_169);
nor U139 (N_139,In_187,In_472);
and U140 (N_140,In_948,In_678);
nand U141 (N_141,In_27,In_845);
nor U142 (N_142,In_919,In_726);
and U143 (N_143,In_628,In_279);
xnor U144 (N_144,In_377,In_43);
and U145 (N_145,In_95,In_962);
nor U146 (N_146,In_225,In_45);
and U147 (N_147,In_506,In_400);
and U148 (N_148,In_700,In_354);
nand U149 (N_149,In_531,In_747);
nand U150 (N_150,In_432,In_180);
or U151 (N_151,In_269,In_268);
and U152 (N_152,In_191,In_109);
or U153 (N_153,In_147,In_930);
or U154 (N_154,In_94,In_397);
nand U155 (N_155,In_562,In_875);
nand U156 (N_156,In_125,In_821);
nor U157 (N_157,In_619,In_730);
or U158 (N_158,In_438,In_272);
and U159 (N_159,In_2,In_101);
or U160 (N_160,In_74,In_478);
and U161 (N_161,In_62,In_66);
xnor U162 (N_162,In_520,In_28);
and U163 (N_163,In_466,In_56);
nand U164 (N_164,In_737,In_226);
nor U165 (N_165,In_817,In_814);
nor U166 (N_166,In_752,In_458);
nor U167 (N_167,In_742,In_658);
and U168 (N_168,In_958,In_599);
xnor U169 (N_169,In_337,In_463);
nand U170 (N_170,In_427,In_803);
and U171 (N_171,In_315,In_416);
nor U172 (N_172,In_181,In_978);
nand U173 (N_173,In_322,In_677);
and U174 (N_174,In_52,In_194);
nand U175 (N_175,In_88,In_116);
nor U176 (N_176,In_188,In_12);
nor U177 (N_177,In_862,In_410);
nor U178 (N_178,In_5,In_867);
nor U179 (N_179,In_798,In_704);
and U180 (N_180,In_713,In_637);
nand U181 (N_181,In_256,In_489);
or U182 (N_182,In_954,In_342);
xnor U183 (N_183,In_343,In_300);
nand U184 (N_184,In_303,In_881);
or U185 (N_185,In_151,In_331);
or U186 (N_186,In_755,In_498);
nor U187 (N_187,In_555,In_235);
nor U188 (N_188,In_262,In_30);
nand U189 (N_189,In_522,In_841);
nand U190 (N_190,In_913,In_986);
nand U191 (N_191,In_358,In_76);
and U192 (N_192,In_3,In_351);
nand U193 (N_193,In_205,In_370);
or U194 (N_194,In_500,In_233);
and U195 (N_195,In_882,In_815);
and U196 (N_196,In_44,In_373);
nor U197 (N_197,In_844,In_566);
and U198 (N_198,In_25,In_707);
xor U199 (N_199,In_142,In_621);
nor U200 (N_200,In_63,In_929);
nand U201 (N_201,In_369,In_247);
and U202 (N_202,In_701,In_481);
nand U203 (N_203,In_324,In_479);
and U204 (N_204,In_611,In_941);
nand U205 (N_205,In_504,In_31);
and U206 (N_206,In_937,In_398);
or U207 (N_207,In_308,In_234);
nor U208 (N_208,In_509,In_899);
xor U209 (N_209,In_189,In_407);
or U210 (N_210,In_470,In_185);
nor U211 (N_211,In_510,In_684);
nor U212 (N_212,In_918,In_210);
xor U213 (N_213,In_266,In_655);
nand U214 (N_214,In_689,In_573);
and U215 (N_215,In_64,In_942);
nand U216 (N_216,In_149,In_781);
nor U217 (N_217,In_532,In_806);
and U218 (N_218,In_731,In_540);
nand U219 (N_219,In_260,In_514);
or U220 (N_220,In_425,In_33);
nand U221 (N_221,In_517,In_673);
and U222 (N_222,In_909,In_65);
xnor U223 (N_223,In_652,In_199);
nand U224 (N_224,In_213,In_102);
and U225 (N_225,In_57,In_624);
xnor U226 (N_226,In_471,In_207);
nand U227 (N_227,In_706,In_975);
and U228 (N_228,In_662,In_718);
and U229 (N_229,In_933,In_375);
or U230 (N_230,In_685,In_381);
and U231 (N_231,In_202,In_529);
and U232 (N_232,In_261,In_748);
and U233 (N_233,In_311,In_211);
nor U234 (N_234,In_883,In_552);
xnor U235 (N_235,In_103,In_734);
or U236 (N_236,In_515,In_777);
xnor U237 (N_237,In_905,In_843);
and U238 (N_238,In_283,In_350);
and U239 (N_239,In_769,In_328);
nand U240 (N_240,In_236,In_253);
and U241 (N_241,In_824,In_645);
and U242 (N_242,In_618,In_32);
and U243 (N_243,In_600,In_17);
nor U244 (N_244,In_727,In_255);
and U245 (N_245,In_288,In_827);
nand U246 (N_246,In_18,In_615);
nand U247 (N_247,In_299,In_387);
and U248 (N_248,In_690,In_622);
and U249 (N_249,In_474,In_648);
nand U250 (N_250,In_497,In_995);
xor U251 (N_251,In_868,In_501);
nand U252 (N_252,In_296,In_816);
nor U253 (N_253,In_965,In_885);
nor U254 (N_254,In_301,In_759);
and U255 (N_255,In_633,In_404);
nand U256 (N_256,In_570,In_130);
nand U257 (N_257,In_414,In_285);
nor U258 (N_258,In_639,In_695);
nand U259 (N_259,In_625,In_702);
nand U260 (N_260,In_694,In_281);
nand U261 (N_261,In_133,In_960);
or U262 (N_262,In_564,In_166);
xor U263 (N_263,In_549,In_391);
and U264 (N_264,In_546,In_48);
or U265 (N_265,In_393,In_190);
nand U266 (N_266,In_484,In_313);
or U267 (N_267,In_424,In_682);
nor U268 (N_268,In_964,In_656);
and U269 (N_269,In_854,In_439);
or U270 (N_270,In_653,In_21);
and U271 (N_271,In_423,In_128);
and U272 (N_272,In_68,In_138);
xor U273 (N_273,In_140,In_295);
xnor U274 (N_274,In_223,In_762);
nor U275 (N_275,In_53,In_348);
and U276 (N_276,In_392,In_212);
xor U277 (N_277,In_411,In_642);
and U278 (N_278,In_528,In_293);
or U279 (N_279,In_984,In_378);
nand U280 (N_280,In_516,In_859);
and U281 (N_281,In_249,In_221);
xnor U282 (N_282,In_591,In_548);
xor U283 (N_283,In_782,In_613);
nand U284 (N_284,In_848,In_873);
and U285 (N_285,In_650,In_519);
nand U286 (N_286,In_448,In_486);
nor U287 (N_287,In_415,In_774);
nand U288 (N_288,In_688,In_172);
xor U289 (N_289,In_981,In_793);
or U290 (N_290,In_746,In_574);
nand U291 (N_291,In_157,In_647);
nand U292 (N_292,In_8,In_4);
and U293 (N_293,In_982,In_766);
and U294 (N_294,In_242,In_456);
or U295 (N_295,In_754,In_9);
or U296 (N_296,In_860,In_850);
xnor U297 (N_297,In_592,In_232);
or U298 (N_298,In_990,In_336);
or U299 (N_299,In_584,In_129);
or U300 (N_300,In_874,In_884);
or U301 (N_301,In_409,In_356);
nand U302 (N_302,In_831,In_134);
nand U303 (N_303,In_973,In_29);
or U304 (N_304,In_488,In_939);
xor U305 (N_305,In_659,In_396);
nor U306 (N_306,In_173,In_715);
xor U307 (N_307,In_779,In_325);
and U308 (N_308,In_697,In_59);
and U309 (N_309,In_545,In_383);
nor U310 (N_310,In_361,In_127);
and U311 (N_311,In_819,In_589);
and U312 (N_312,In_795,In_542);
and U313 (N_313,In_163,In_229);
nor U314 (N_314,In_80,In_904);
or U315 (N_315,In_493,In_593);
and U316 (N_316,In_363,In_598);
nand U317 (N_317,In_851,In_888);
or U318 (N_318,In_192,In_382);
or U319 (N_319,In_787,In_98);
nand U320 (N_320,In_558,In_895);
nand U321 (N_321,In_595,In_399);
nand U322 (N_322,In_523,In_741);
nand U323 (N_323,In_482,In_670);
nand U324 (N_324,In_832,In_784);
and U325 (N_325,In_849,In_556);
or U326 (N_326,In_771,In_0);
nor U327 (N_327,In_544,In_376);
nand U328 (N_328,In_902,In_536);
nand U329 (N_329,In_963,In_724);
or U330 (N_330,In_105,In_436);
or U331 (N_331,In_332,In_219);
or U332 (N_332,In_265,In_518);
nor U333 (N_333,In_533,In_273);
xnor U334 (N_334,In_945,In_374);
or U335 (N_335,In_778,In_406);
and U336 (N_336,In_686,In_316);
and U337 (N_337,In_938,In_464);
nor U338 (N_338,In_898,In_46);
xnor U339 (N_339,In_597,In_176);
and U340 (N_340,In_792,In_451);
and U341 (N_341,In_623,In_35);
nor U342 (N_342,In_218,In_114);
and U343 (N_343,In_291,In_113);
nor U344 (N_344,In_711,In_513);
nor U345 (N_345,In_607,In_596);
and U346 (N_346,In_917,In_237);
or U347 (N_347,In_683,In_666);
nor U348 (N_348,In_434,In_858);
or U349 (N_349,In_503,In_421);
and U350 (N_350,In_970,In_347);
and U351 (N_351,In_203,In_627);
nor U352 (N_352,In_154,In_86);
nand U353 (N_353,In_554,In_996);
nand U354 (N_354,In_314,In_610);
or U355 (N_355,In_987,In_287);
nand U356 (N_356,In_10,In_823);
or U357 (N_357,In_11,In_887);
nand U358 (N_358,In_175,In_530);
or U359 (N_359,In_372,In_720);
nor U360 (N_360,In_450,In_426);
nor U361 (N_361,In_115,In_550);
xnor U362 (N_362,In_227,In_758);
or U363 (N_363,In_41,In_829);
and U364 (N_364,In_961,In_294);
and U365 (N_365,In_644,In_368);
and U366 (N_366,In_634,In_575);
nand U367 (N_367,In_788,In_419);
and U368 (N_368,In_657,In_267);
and U369 (N_369,In_667,In_675);
nor U370 (N_370,In_604,In_162);
nand U371 (N_371,In_569,In_258);
and U372 (N_372,In_465,In_71);
and U373 (N_373,In_271,In_304);
nor U374 (N_374,In_47,In_345);
or U375 (N_375,In_920,In_947);
and U376 (N_376,In_99,In_305);
or U377 (N_377,In_453,In_988);
and U378 (N_378,In_141,In_455);
and U379 (N_379,In_87,In_608);
or U380 (N_380,In_765,In_614);
nand U381 (N_381,In_571,In_77);
and U382 (N_382,In_505,In_341);
or U383 (N_383,In_989,In_834);
or U384 (N_384,In_810,In_983);
or U385 (N_385,In_183,In_535);
or U386 (N_386,In_446,In_380);
and U387 (N_387,In_340,In_435);
nand U388 (N_388,In_161,In_405);
nor U389 (N_389,In_495,In_712);
nand U390 (N_390,In_785,In_93);
nor U391 (N_391,In_121,In_714);
nor U392 (N_392,In_204,In_856);
nor U393 (N_393,In_903,In_914);
and U394 (N_394,In_911,In_442);
nor U395 (N_395,In_525,In_42);
nand U396 (N_396,In_944,In_708);
and U397 (N_397,In_13,In_745);
nor U398 (N_398,In_67,In_935);
nor U399 (N_399,In_257,In_15);
and U400 (N_400,In_837,In_390);
and U401 (N_401,In_629,In_660);
nand U402 (N_402,In_612,In_977);
or U403 (N_403,In_61,In_931);
and U404 (N_404,In_804,In_79);
and U405 (N_405,In_738,In_485);
and U406 (N_406,In_751,In_275);
or U407 (N_407,In_577,In_999);
nor U408 (N_408,In_855,In_772);
xor U409 (N_409,In_770,In_246);
nand U410 (N_410,In_846,In_676);
nor U411 (N_411,In_412,In_729);
xnor U412 (N_412,In_284,In_126);
and U413 (N_413,In_967,In_539);
xnor U414 (N_414,In_366,In_620);
or U415 (N_415,In_50,In_197);
nor U416 (N_416,In_179,In_812);
and U417 (N_417,In_487,In_408);
nand U418 (N_418,In_908,In_876);
and U419 (N_419,In_572,In_636);
nand U420 (N_420,In_654,In_307);
nand U421 (N_421,In_679,In_680);
and U422 (N_422,In_496,In_789);
and U423 (N_423,In_646,In_364);
or U424 (N_424,In_543,In_800);
nand U425 (N_425,In_794,In_317);
nor U426 (N_426,In_663,In_357);
nand U427 (N_427,In_145,In_239);
nor U428 (N_428,In_6,In_385);
nor U429 (N_429,In_112,In_786);
and U430 (N_430,In_167,In_319);
nand U431 (N_431,In_156,In_925);
and U432 (N_432,In_980,In_492);
nor U433 (N_433,In_847,In_449);
nor U434 (N_434,In_717,In_290);
nand U435 (N_435,In_698,In_951);
nor U436 (N_436,In_144,In_476);
or U437 (N_437,In_379,In_82);
nand U438 (N_438,In_580,In_90);
nand U439 (N_439,In_893,In_217);
xor U440 (N_440,In_802,In_561);
or U441 (N_441,In_230,In_768);
nor U442 (N_442,In_228,In_131);
or U443 (N_443,In_259,In_278);
xnor U444 (N_444,In_483,In_705);
nand U445 (N_445,In_353,In_877);
nor U446 (N_446,In_992,In_100);
xnor U447 (N_447,In_334,In_245);
nor U448 (N_448,In_475,In_879);
and U449 (N_449,In_586,In_83);
nand U450 (N_450,In_352,In_889);
nor U451 (N_451,In_394,In_739);
and U452 (N_452,In_826,In_878);
and U453 (N_453,In_494,In_559);
xor U454 (N_454,In_928,In_78);
or U455 (N_455,In_696,In_998);
or U456 (N_456,In_956,In_916);
or U457 (N_457,In_828,In_912);
or U458 (N_458,In_118,In_551);
and U459 (N_459,In_853,In_222);
nand U460 (N_460,In_69,In_346);
or U461 (N_461,In_452,In_171);
nor U462 (N_462,In_461,In_34);
or U463 (N_463,In_756,In_852);
nor U464 (N_464,In_830,In_298);
nand U465 (N_465,In_820,In_276);
and U466 (N_466,In_825,In_335);
nand U467 (N_467,In_418,In_617);
nand U468 (N_468,In_760,In_480);
nor U469 (N_469,In_365,In_238);
nand U470 (N_470,In_871,In_349);
nand U471 (N_471,In_750,In_430);
nand U472 (N_472,In_578,In_248);
and U473 (N_473,In_783,In_553);
and U474 (N_474,In_609,In_692);
nor U475 (N_475,In_60,In_691);
and U476 (N_476,In_148,In_26);
and U477 (N_477,In_869,In_512);
nor U478 (N_478,In_220,In_280);
or U479 (N_479,In_150,In_594);
and U480 (N_480,In_292,In_863);
or U481 (N_481,In_54,In_473);
or U482 (N_482,In_355,In_200);
and U483 (N_483,In_96,In_870);
and U484 (N_484,In_733,In_805);
or U485 (N_485,In_1,In_861);
nor U486 (N_486,In_91,In_367);
nor U487 (N_487,In_277,In_946);
and U488 (N_488,In_976,In_51);
xnor U489 (N_489,In_668,In_49);
or U490 (N_490,In_744,In_323);
nand U491 (N_491,In_327,In_840);
nor U492 (N_492,In_85,In_721);
and U493 (N_493,In_985,In_906);
or U494 (N_494,In_894,In_433);
nand U495 (N_495,In_186,In_896);
nor U496 (N_496,In_927,In_886);
and U497 (N_497,In_775,In_263);
nand U498 (N_498,In_216,In_431);
nand U499 (N_499,In_417,In_565);
or U500 (N_500,In_408,In_448);
and U501 (N_501,In_926,In_345);
nand U502 (N_502,In_657,In_873);
nand U503 (N_503,In_36,In_902);
or U504 (N_504,In_759,In_440);
and U505 (N_505,In_15,In_107);
nor U506 (N_506,In_995,In_9);
nand U507 (N_507,In_769,In_907);
and U508 (N_508,In_991,In_957);
nand U509 (N_509,In_728,In_595);
xor U510 (N_510,In_322,In_258);
nand U511 (N_511,In_76,In_602);
and U512 (N_512,In_735,In_646);
and U513 (N_513,In_658,In_70);
nor U514 (N_514,In_613,In_624);
and U515 (N_515,In_57,In_895);
xor U516 (N_516,In_699,In_738);
or U517 (N_517,In_575,In_479);
nand U518 (N_518,In_409,In_766);
xor U519 (N_519,In_866,In_126);
nor U520 (N_520,In_888,In_152);
nand U521 (N_521,In_365,In_848);
nor U522 (N_522,In_980,In_423);
nand U523 (N_523,In_485,In_184);
nand U524 (N_524,In_969,In_240);
nor U525 (N_525,In_975,In_228);
nor U526 (N_526,In_356,In_464);
or U527 (N_527,In_970,In_950);
and U528 (N_528,In_511,In_846);
nor U529 (N_529,In_244,In_421);
nor U530 (N_530,In_601,In_523);
and U531 (N_531,In_966,In_628);
nor U532 (N_532,In_479,In_310);
and U533 (N_533,In_843,In_259);
or U534 (N_534,In_541,In_28);
or U535 (N_535,In_130,In_778);
xor U536 (N_536,In_86,In_998);
or U537 (N_537,In_167,In_559);
nor U538 (N_538,In_296,In_460);
nand U539 (N_539,In_199,In_467);
nand U540 (N_540,In_77,In_281);
nor U541 (N_541,In_388,In_174);
and U542 (N_542,In_596,In_845);
nor U543 (N_543,In_851,In_479);
nor U544 (N_544,In_437,In_745);
and U545 (N_545,In_746,In_85);
and U546 (N_546,In_476,In_163);
or U547 (N_547,In_87,In_898);
nand U548 (N_548,In_71,In_745);
xor U549 (N_549,In_175,In_267);
nand U550 (N_550,In_700,In_346);
nor U551 (N_551,In_32,In_233);
nand U552 (N_552,In_326,In_43);
xor U553 (N_553,In_900,In_610);
nor U554 (N_554,In_839,In_362);
and U555 (N_555,In_181,In_9);
or U556 (N_556,In_494,In_653);
or U557 (N_557,In_248,In_467);
or U558 (N_558,In_337,In_257);
and U559 (N_559,In_889,In_50);
nor U560 (N_560,In_993,In_803);
and U561 (N_561,In_74,In_911);
and U562 (N_562,In_980,In_789);
nand U563 (N_563,In_837,In_763);
nor U564 (N_564,In_87,In_582);
nor U565 (N_565,In_738,In_172);
or U566 (N_566,In_497,In_676);
or U567 (N_567,In_389,In_345);
nand U568 (N_568,In_245,In_919);
xnor U569 (N_569,In_936,In_767);
and U570 (N_570,In_941,In_375);
xnor U571 (N_571,In_515,In_468);
and U572 (N_572,In_850,In_980);
nor U573 (N_573,In_20,In_881);
xor U574 (N_574,In_535,In_173);
nor U575 (N_575,In_455,In_602);
or U576 (N_576,In_186,In_614);
nor U577 (N_577,In_694,In_732);
nor U578 (N_578,In_453,In_384);
nor U579 (N_579,In_791,In_904);
nand U580 (N_580,In_128,In_212);
and U581 (N_581,In_552,In_721);
nor U582 (N_582,In_586,In_570);
nor U583 (N_583,In_147,In_669);
nor U584 (N_584,In_167,In_278);
or U585 (N_585,In_162,In_141);
nor U586 (N_586,In_680,In_147);
xnor U587 (N_587,In_546,In_878);
xnor U588 (N_588,In_86,In_894);
and U589 (N_589,In_785,In_683);
or U590 (N_590,In_204,In_762);
and U591 (N_591,In_268,In_665);
or U592 (N_592,In_789,In_467);
or U593 (N_593,In_281,In_636);
nor U594 (N_594,In_907,In_460);
and U595 (N_595,In_307,In_614);
nor U596 (N_596,In_327,In_646);
nor U597 (N_597,In_807,In_371);
and U598 (N_598,In_199,In_539);
and U599 (N_599,In_517,In_118);
nand U600 (N_600,In_613,In_500);
or U601 (N_601,In_706,In_256);
or U602 (N_602,In_398,In_289);
nand U603 (N_603,In_883,In_594);
nor U604 (N_604,In_487,In_976);
and U605 (N_605,In_909,In_146);
xnor U606 (N_606,In_711,In_359);
or U607 (N_607,In_256,In_998);
nand U608 (N_608,In_875,In_611);
or U609 (N_609,In_458,In_448);
and U610 (N_610,In_600,In_728);
nand U611 (N_611,In_416,In_875);
nor U612 (N_612,In_624,In_552);
nand U613 (N_613,In_515,In_39);
or U614 (N_614,In_944,In_537);
nand U615 (N_615,In_936,In_389);
nand U616 (N_616,In_355,In_275);
and U617 (N_617,In_944,In_886);
and U618 (N_618,In_306,In_669);
nand U619 (N_619,In_524,In_338);
nor U620 (N_620,In_385,In_261);
or U621 (N_621,In_33,In_67);
nand U622 (N_622,In_319,In_582);
or U623 (N_623,In_623,In_532);
nand U624 (N_624,In_284,In_946);
nand U625 (N_625,In_102,In_165);
nor U626 (N_626,In_56,In_577);
nand U627 (N_627,In_50,In_655);
and U628 (N_628,In_748,In_414);
or U629 (N_629,In_462,In_112);
and U630 (N_630,In_714,In_89);
and U631 (N_631,In_758,In_377);
and U632 (N_632,In_460,In_677);
and U633 (N_633,In_257,In_14);
or U634 (N_634,In_198,In_202);
and U635 (N_635,In_617,In_97);
or U636 (N_636,In_591,In_210);
xnor U637 (N_637,In_503,In_535);
xor U638 (N_638,In_221,In_378);
and U639 (N_639,In_478,In_753);
or U640 (N_640,In_523,In_477);
xnor U641 (N_641,In_531,In_65);
or U642 (N_642,In_360,In_479);
nand U643 (N_643,In_186,In_616);
or U644 (N_644,In_904,In_980);
nand U645 (N_645,In_737,In_285);
nor U646 (N_646,In_821,In_208);
nor U647 (N_647,In_159,In_867);
nor U648 (N_648,In_133,In_213);
or U649 (N_649,In_205,In_347);
or U650 (N_650,In_649,In_611);
nor U651 (N_651,In_469,In_672);
and U652 (N_652,In_228,In_440);
or U653 (N_653,In_706,In_290);
xnor U654 (N_654,In_111,In_677);
or U655 (N_655,In_173,In_378);
nand U656 (N_656,In_302,In_435);
nor U657 (N_657,In_200,In_646);
or U658 (N_658,In_458,In_329);
or U659 (N_659,In_117,In_811);
xor U660 (N_660,In_483,In_485);
nor U661 (N_661,In_656,In_129);
nand U662 (N_662,In_504,In_882);
nor U663 (N_663,In_508,In_89);
or U664 (N_664,In_426,In_343);
xnor U665 (N_665,In_900,In_716);
or U666 (N_666,In_308,In_731);
and U667 (N_667,In_301,In_389);
nand U668 (N_668,In_52,In_738);
nand U669 (N_669,In_249,In_258);
nand U670 (N_670,In_615,In_373);
nand U671 (N_671,In_875,In_193);
xnor U672 (N_672,In_24,In_107);
nor U673 (N_673,In_309,In_631);
or U674 (N_674,In_873,In_380);
nor U675 (N_675,In_869,In_784);
nor U676 (N_676,In_98,In_0);
nand U677 (N_677,In_210,In_529);
or U678 (N_678,In_743,In_658);
or U679 (N_679,In_665,In_369);
nand U680 (N_680,In_128,In_254);
nand U681 (N_681,In_520,In_82);
or U682 (N_682,In_452,In_944);
xnor U683 (N_683,In_447,In_3);
nor U684 (N_684,In_484,In_191);
nor U685 (N_685,In_254,In_754);
and U686 (N_686,In_873,In_878);
xor U687 (N_687,In_884,In_752);
xor U688 (N_688,In_493,In_105);
nor U689 (N_689,In_371,In_601);
or U690 (N_690,In_301,In_390);
nor U691 (N_691,In_8,In_782);
nand U692 (N_692,In_764,In_641);
nor U693 (N_693,In_59,In_572);
nand U694 (N_694,In_299,In_284);
nor U695 (N_695,In_557,In_683);
or U696 (N_696,In_38,In_496);
or U697 (N_697,In_501,In_739);
xor U698 (N_698,In_234,In_328);
and U699 (N_699,In_345,In_290);
and U700 (N_700,In_701,In_974);
nor U701 (N_701,In_705,In_436);
nand U702 (N_702,In_495,In_222);
or U703 (N_703,In_679,In_854);
xor U704 (N_704,In_979,In_468);
nand U705 (N_705,In_825,In_810);
nand U706 (N_706,In_208,In_817);
or U707 (N_707,In_326,In_807);
xnor U708 (N_708,In_346,In_697);
nand U709 (N_709,In_199,In_922);
nor U710 (N_710,In_565,In_559);
nand U711 (N_711,In_219,In_581);
nand U712 (N_712,In_411,In_210);
nor U713 (N_713,In_766,In_386);
or U714 (N_714,In_577,In_443);
nor U715 (N_715,In_854,In_861);
nor U716 (N_716,In_109,In_39);
nand U717 (N_717,In_259,In_434);
xnor U718 (N_718,In_506,In_89);
and U719 (N_719,In_340,In_534);
and U720 (N_720,In_68,In_204);
xor U721 (N_721,In_320,In_888);
nor U722 (N_722,In_738,In_742);
nor U723 (N_723,In_204,In_579);
nor U724 (N_724,In_104,In_664);
nand U725 (N_725,In_126,In_984);
nand U726 (N_726,In_849,In_559);
nor U727 (N_727,In_942,In_472);
xnor U728 (N_728,In_558,In_202);
nand U729 (N_729,In_135,In_281);
nor U730 (N_730,In_660,In_123);
and U731 (N_731,In_139,In_462);
nor U732 (N_732,In_355,In_181);
nor U733 (N_733,In_78,In_240);
or U734 (N_734,In_558,In_280);
and U735 (N_735,In_271,In_224);
nor U736 (N_736,In_524,In_177);
and U737 (N_737,In_670,In_709);
nand U738 (N_738,In_805,In_52);
nand U739 (N_739,In_378,In_611);
xnor U740 (N_740,In_646,In_724);
or U741 (N_741,In_801,In_658);
nor U742 (N_742,In_753,In_829);
nor U743 (N_743,In_270,In_63);
or U744 (N_744,In_767,In_602);
nor U745 (N_745,In_352,In_862);
xnor U746 (N_746,In_306,In_827);
xor U747 (N_747,In_214,In_890);
or U748 (N_748,In_323,In_21);
nor U749 (N_749,In_676,In_65);
nor U750 (N_750,In_812,In_622);
and U751 (N_751,In_106,In_350);
nand U752 (N_752,In_876,In_324);
nor U753 (N_753,In_561,In_851);
and U754 (N_754,In_289,In_45);
nand U755 (N_755,In_874,In_48);
or U756 (N_756,In_467,In_513);
nor U757 (N_757,In_599,In_730);
nor U758 (N_758,In_858,In_669);
nor U759 (N_759,In_630,In_74);
nor U760 (N_760,In_284,In_589);
nand U761 (N_761,In_403,In_263);
nand U762 (N_762,In_797,In_206);
and U763 (N_763,In_6,In_618);
or U764 (N_764,In_964,In_96);
nand U765 (N_765,In_47,In_432);
and U766 (N_766,In_965,In_646);
nand U767 (N_767,In_747,In_925);
and U768 (N_768,In_238,In_625);
nor U769 (N_769,In_394,In_806);
nor U770 (N_770,In_643,In_710);
or U771 (N_771,In_352,In_187);
nand U772 (N_772,In_669,In_822);
or U773 (N_773,In_348,In_518);
and U774 (N_774,In_338,In_85);
nand U775 (N_775,In_53,In_903);
nor U776 (N_776,In_605,In_335);
nand U777 (N_777,In_38,In_263);
nor U778 (N_778,In_97,In_736);
or U779 (N_779,In_200,In_875);
xor U780 (N_780,In_935,In_535);
nor U781 (N_781,In_671,In_475);
and U782 (N_782,In_495,In_64);
nor U783 (N_783,In_724,In_906);
xor U784 (N_784,In_553,In_204);
nand U785 (N_785,In_394,In_43);
and U786 (N_786,In_120,In_44);
nand U787 (N_787,In_802,In_242);
nand U788 (N_788,In_700,In_177);
nand U789 (N_789,In_752,In_897);
and U790 (N_790,In_83,In_561);
nand U791 (N_791,In_615,In_223);
nor U792 (N_792,In_806,In_71);
and U793 (N_793,In_577,In_415);
nand U794 (N_794,In_514,In_372);
and U795 (N_795,In_89,In_411);
nand U796 (N_796,In_848,In_205);
or U797 (N_797,In_49,In_47);
nor U798 (N_798,In_241,In_337);
nand U799 (N_799,In_968,In_129);
or U800 (N_800,In_585,In_538);
nor U801 (N_801,In_333,In_763);
nand U802 (N_802,In_842,In_662);
and U803 (N_803,In_447,In_323);
nand U804 (N_804,In_354,In_384);
or U805 (N_805,In_295,In_984);
xnor U806 (N_806,In_676,In_867);
nor U807 (N_807,In_828,In_955);
and U808 (N_808,In_484,In_891);
nand U809 (N_809,In_564,In_304);
and U810 (N_810,In_638,In_45);
nand U811 (N_811,In_812,In_727);
nand U812 (N_812,In_850,In_164);
nor U813 (N_813,In_316,In_202);
xor U814 (N_814,In_391,In_813);
or U815 (N_815,In_394,In_615);
nand U816 (N_816,In_88,In_475);
and U817 (N_817,In_31,In_309);
xnor U818 (N_818,In_46,In_618);
or U819 (N_819,In_179,In_931);
nor U820 (N_820,In_931,In_903);
or U821 (N_821,In_283,In_722);
nand U822 (N_822,In_668,In_161);
and U823 (N_823,In_576,In_986);
or U824 (N_824,In_305,In_254);
and U825 (N_825,In_3,In_813);
nand U826 (N_826,In_881,In_410);
or U827 (N_827,In_465,In_886);
or U828 (N_828,In_725,In_440);
xor U829 (N_829,In_940,In_889);
nor U830 (N_830,In_848,In_806);
and U831 (N_831,In_208,In_953);
or U832 (N_832,In_266,In_772);
nand U833 (N_833,In_844,In_961);
nor U834 (N_834,In_198,In_998);
or U835 (N_835,In_196,In_805);
or U836 (N_836,In_416,In_800);
and U837 (N_837,In_765,In_13);
xor U838 (N_838,In_13,In_259);
and U839 (N_839,In_108,In_901);
or U840 (N_840,In_817,In_818);
nor U841 (N_841,In_270,In_68);
nand U842 (N_842,In_498,In_262);
and U843 (N_843,In_959,In_138);
nor U844 (N_844,In_747,In_265);
nor U845 (N_845,In_564,In_549);
nand U846 (N_846,In_915,In_44);
nor U847 (N_847,In_157,In_853);
nor U848 (N_848,In_940,In_291);
and U849 (N_849,In_237,In_810);
or U850 (N_850,In_630,In_389);
nand U851 (N_851,In_561,In_229);
or U852 (N_852,In_109,In_739);
or U853 (N_853,In_361,In_128);
or U854 (N_854,In_205,In_726);
or U855 (N_855,In_337,In_88);
xor U856 (N_856,In_870,In_868);
nand U857 (N_857,In_903,In_727);
nand U858 (N_858,In_999,In_793);
and U859 (N_859,In_193,In_805);
nand U860 (N_860,In_360,In_771);
nor U861 (N_861,In_868,In_544);
or U862 (N_862,In_888,In_877);
nand U863 (N_863,In_447,In_387);
or U864 (N_864,In_133,In_228);
and U865 (N_865,In_913,In_538);
nand U866 (N_866,In_55,In_948);
or U867 (N_867,In_434,In_92);
and U868 (N_868,In_1,In_714);
and U869 (N_869,In_194,In_370);
nand U870 (N_870,In_208,In_899);
nand U871 (N_871,In_107,In_297);
nor U872 (N_872,In_782,In_415);
nand U873 (N_873,In_680,In_549);
or U874 (N_874,In_840,In_381);
nor U875 (N_875,In_914,In_172);
nand U876 (N_876,In_749,In_941);
nor U877 (N_877,In_580,In_929);
and U878 (N_878,In_392,In_964);
nor U879 (N_879,In_207,In_34);
nor U880 (N_880,In_704,In_404);
or U881 (N_881,In_946,In_69);
or U882 (N_882,In_52,In_598);
and U883 (N_883,In_904,In_551);
and U884 (N_884,In_767,In_369);
nor U885 (N_885,In_405,In_470);
nand U886 (N_886,In_696,In_29);
and U887 (N_887,In_695,In_352);
nand U888 (N_888,In_30,In_16);
nor U889 (N_889,In_178,In_763);
nand U890 (N_890,In_980,In_793);
xor U891 (N_891,In_411,In_966);
nor U892 (N_892,In_475,In_94);
nor U893 (N_893,In_905,In_464);
nor U894 (N_894,In_480,In_257);
or U895 (N_895,In_823,In_650);
nand U896 (N_896,In_861,In_949);
or U897 (N_897,In_421,In_350);
xnor U898 (N_898,In_463,In_385);
nor U899 (N_899,In_730,In_31);
and U900 (N_900,In_529,In_432);
nor U901 (N_901,In_748,In_204);
xnor U902 (N_902,In_312,In_25);
and U903 (N_903,In_242,In_85);
or U904 (N_904,In_293,In_482);
nand U905 (N_905,In_387,In_143);
nor U906 (N_906,In_859,In_282);
and U907 (N_907,In_457,In_128);
or U908 (N_908,In_237,In_795);
nor U909 (N_909,In_583,In_66);
nor U910 (N_910,In_919,In_246);
nor U911 (N_911,In_429,In_839);
and U912 (N_912,In_553,In_482);
nand U913 (N_913,In_197,In_925);
nor U914 (N_914,In_379,In_301);
and U915 (N_915,In_790,In_635);
nor U916 (N_916,In_527,In_912);
nor U917 (N_917,In_392,In_361);
nand U918 (N_918,In_812,In_923);
or U919 (N_919,In_184,In_229);
nand U920 (N_920,In_776,In_357);
and U921 (N_921,In_542,In_500);
and U922 (N_922,In_434,In_583);
xnor U923 (N_923,In_456,In_286);
nand U924 (N_924,In_439,In_619);
or U925 (N_925,In_568,In_355);
and U926 (N_926,In_267,In_398);
nor U927 (N_927,In_133,In_208);
or U928 (N_928,In_34,In_163);
or U929 (N_929,In_364,In_489);
nand U930 (N_930,In_960,In_11);
and U931 (N_931,In_383,In_514);
and U932 (N_932,In_193,In_736);
and U933 (N_933,In_143,In_903);
or U934 (N_934,In_559,In_823);
nand U935 (N_935,In_543,In_993);
and U936 (N_936,In_137,In_834);
nand U937 (N_937,In_453,In_651);
or U938 (N_938,In_628,In_183);
xor U939 (N_939,In_533,In_166);
and U940 (N_940,In_445,In_325);
nor U941 (N_941,In_606,In_986);
and U942 (N_942,In_900,In_128);
nand U943 (N_943,In_76,In_986);
and U944 (N_944,In_162,In_814);
and U945 (N_945,In_330,In_291);
or U946 (N_946,In_850,In_486);
or U947 (N_947,In_850,In_856);
xor U948 (N_948,In_137,In_548);
and U949 (N_949,In_627,In_917);
nand U950 (N_950,In_898,In_287);
nand U951 (N_951,In_430,In_593);
or U952 (N_952,In_236,In_940);
nor U953 (N_953,In_236,In_883);
nand U954 (N_954,In_706,In_358);
nand U955 (N_955,In_931,In_109);
and U956 (N_956,In_515,In_24);
and U957 (N_957,In_185,In_273);
nand U958 (N_958,In_725,In_577);
nand U959 (N_959,In_131,In_537);
nor U960 (N_960,In_869,In_490);
nor U961 (N_961,In_276,In_554);
nand U962 (N_962,In_467,In_305);
nor U963 (N_963,In_256,In_488);
or U964 (N_964,In_668,In_441);
nor U965 (N_965,In_756,In_737);
and U966 (N_966,In_520,In_205);
xnor U967 (N_967,In_821,In_785);
nand U968 (N_968,In_755,In_968);
nand U969 (N_969,In_245,In_115);
nor U970 (N_970,In_172,In_848);
nand U971 (N_971,In_859,In_441);
nand U972 (N_972,In_913,In_440);
nor U973 (N_973,In_436,In_466);
or U974 (N_974,In_742,In_376);
or U975 (N_975,In_37,In_187);
and U976 (N_976,In_271,In_688);
nand U977 (N_977,In_738,In_219);
or U978 (N_978,In_165,In_174);
nor U979 (N_979,In_104,In_480);
or U980 (N_980,In_434,In_332);
and U981 (N_981,In_730,In_169);
nand U982 (N_982,In_11,In_152);
nand U983 (N_983,In_273,In_43);
or U984 (N_984,In_406,In_806);
or U985 (N_985,In_764,In_451);
and U986 (N_986,In_497,In_886);
nand U987 (N_987,In_893,In_481);
xor U988 (N_988,In_27,In_493);
and U989 (N_989,In_307,In_4);
nand U990 (N_990,In_172,In_284);
xor U991 (N_991,In_289,In_851);
xor U992 (N_992,In_752,In_860);
nand U993 (N_993,In_207,In_844);
nor U994 (N_994,In_30,In_510);
nor U995 (N_995,In_91,In_913);
xor U996 (N_996,In_546,In_575);
nor U997 (N_997,In_112,In_295);
and U998 (N_998,In_29,In_959);
or U999 (N_999,In_992,In_575);
and U1000 (N_1000,In_500,In_717);
nand U1001 (N_1001,In_352,In_666);
nor U1002 (N_1002,In_471,In_608);
or U1003 (N_1003,In_320,In_219);
or U1004 (N_1004,In_330,In_863);
or U1005 (N_1005,In_427,In_549);
nor U1006 (N_1006,In_639,In_700);
nand U1007 (N_1007,In_346,In_837);
nor U1008 (N_1008,In_307,In_935);
nor U1009 (N_1009,In_145,In_564);
nand U1010 (N_1010,In_380,In_640);
xor U1011 (N_1011,In_804,In_228);
or U1012 (N_1012,In_873,In_560);
nor U1013 (N_1013,In_200,In_276);
and U1014 (N_1014,In_29,In_957);
xor U1015 (N_1015,In_474,In_155);
or U1016 (N_1016,In_647,In_795);
nor U1017 (N_1017,In_787,In_198);
and U1018 (N_1018,In_62,In_719);
and U1019 (N_1019,In_570,In_235);
or U1020 (N_1020,In_669,In_153);
or U1021 (N_1021,In_153,In_648);
nor U1022 (N_1022,In_566,In_802);
and U1023 (N_1023,In_366,In_953);
nor U1024 (N_1024,In_106,In_131);
or U1025 (N_1025,In_167,In_997);
and U1026 (N_1026,In_877,In_550);
nand U1027 (N_1027,In_664,In_274);
nand U1028 (N_1028,In_826,In_423);
or U1029 (N_1029,In_346,In_851);
or U1030 (N_1030,In_461,In_272);
and U1031 (N_1031,In_965,In_320);
or U1032 (N_1032,In_732,In_292);
nor U1033 (N_1033,In_660,In_284);
or U1034 (N_1034,In_550,In_771);
nand U1035 (N_1035,In_917,In_4);
or U1036 (N_1036,In_332,In_250);
nor U1037 (N_1037,In_551,In_857);
nor U1038 (N_1038,In_260,In_101);
nor U1039 (N_1039,In_766,In_862);
or U1040 (N_1040,In_150,In_315);
nor U1041 (N_1041,In_503,In_22);
and U1042 (N_1042,In_801,In_465);
nor U1043 (N_1043,In_38,In_273);
xnor U1044 (N_1044,In_285,In_62);
and U1045 (N_1045,In_519,In_263);
nand U1046 (N_1046,In_851,In_526);
or U1047 (N_1047,In_840,In_653);
nor U1048 (N_1048,In_960,In_967);
or U1049 (N_1049,In_26,In_818);
nand U1050 (N_1050,In_561,In_102);
nor U1051 (N_1051,In_180,In_96);
nand U1052 (N_1052,In_72,In_854);
nor U1053 (N_1053,In_620,In_281);
or U1054 (N_1054,In_306,In_282);
or U1055 (N_1055,In_42,In_652);
nand U1056 (N_1056,In_790,In_568);
nor U1057 (N_1057,In_601,In_826);
or U1058 (N_1058,In_943,In_295);
nor U1059 (N_1059,In_660,In_239);
or U1060 (N_1060,In_591,In_770);
or U1061 (N_1061,In_365,In_333);
and U1062 (N_1062,In_595,In_110);
or U1063 (N_1063,In_138,In_117);
nand U1064 (N_1064,In_652,In_644);
and U1065 (N_1065,In_565,In_742);
or U1066 (N_1066,In_701,In_810);
or U1067 (N_1067,In_66,In_745);
nand U1068 (N_1068,In_328,In_194);
and U1069 (N_1069,In_657,In_463);
and U1070 (N_1070,In_290,In_520);
xnor U1071 (N_1071,In_952,In_127);
or U1072 (N_1072,In_592,In_69);
nor U1073 (N_1073,In_442,In_38);
or U1074 (N_1074,In_419,In_54);
nor U1075 (N_1075,In_776,In_647);
nand U1076 (N_1076,In_564,In_615);
and U1077 (N_1077,In_987,In_919);
or U1078 (N_1078,In_582,In_224);
nor U1079 (N_1079,In_487,In_103);
and U1080 (N_1080,In_57,In_365);
nor U1081 (N_1081,In_573,In_759);
nor U1082 (N_1082,In_776,In_196);
or U1083 (N_1083,In_331,In_913);
and U1084 (N_1084,In_898,In_32);
xor U1085 (N_1085,In_120,In_71);
and U1086 (N_1086,In_44,In_287);
nor U1087 (N_1087,In_689,In_754);
xnor U1088 (N_1088,In_892,In_563);
and U1089 (N_1089,In_547,In_153);
and U1090 (N_1090,In_900,In_892);
and U1091 (N_1091,In_347,In_137);
and U1092 (N_1092,In_552,In_775);
nand U1093 (N_1093,In_742,In_486);
nand U1094 (N_1094,In_54,In_118);
nand U1095 (N_1095,In_631,In_598);
nor U1096 (N_1096,In_96,In_164);
and U1097 (N_1097,In_905,In_200);
and U1098 (N_1098,In_197,In_496);
and U1099 (N_1099,In_435,In_714);
nand U1100 (N_1100,In_376,In_885);
nand U1101 (N_1101,In_835,In_135);
or U1102 (N_1102,In_918,In_164);
xnor U1103 (N_1103,In_957,In_548);
or U1104 (N_1104,In_790,In_347);
nor U1105 (N_1105,In_128,In_389);
and U1106 (N_1106,In_933,In_382);
nand U1107 (N_1107,In_857,In_94);
nor U1108 (N_1108,In_212,In_220);
nor U1109 (N_1109,In_936,In_887);
and U1110 (N_1110,In_544,In_94);
or U1111 (N_1111,In_151,In_437);
nand U1112 (N_1112,In_441,In_845);
nand U1113 (N_1113,In_164,In_228);
nor U1114 (N_1114,In_266,In_609);
xor U1115 (N_1115,In_17,In_445);
or U1116 (N_1116,In_968,In_207);
nor U1117 (N_1117,In_534,In_416);
nor U1118 (N_1118,In_894,In_222);
nand U1119 (N_1119,In_129,In_595);
and U1120 (N_1120,In_632,In_400);
xor U1121 (N_1121,In_794,In_329);
nor U1122 (N_1122,In_405,In_297);
or U1123 (N_1123,In_938,In_407);
nor U1124 (N_1124,In_899,In_515);
or U1125 (N_1125,In_231,In_288);
and U1126 (N_1126,In_61,In_545);
nor U1127 (N_1127,In_31,In_966);
and U1128 (N_1128,In_637,In_289);
nor U1129 (N_1129,In_15,In_545);
nand U1130 (N_1130,In_111,In_377);
nor U1131 (N_1131,In_554,In_238);
or U1132 (N_1132,In_758,In_905);
xor U1133 (N_1133,In_555,In_958);
nand U1134 (N_1134,In_125,In_498);
nand U1135 (N_1135,In_564,In_44);
xnor U1136 (N_1136,In_505,In_705);
nand U1137 (N_1137,In_507,In_551);
xnor U1138 (N_1138,In_894,In_49);
and U1139 (N_1139,In_429,In_391);
nor U1140 (N_1140,In_202,In_712);
nand U1141 (N_1141,In_279,In_394);
nor U1142 (N_1142,In_469,In_3);
or U1143 (N_1143,In_313,In_594);
nand U1144 (N_1144,In_670,In_199);
nor U1145 (N_1145,In_975,In_266);
nor U1146 (N_1146,In_699,In_2);
nand U1147 (N_1147,In_348,In_218);
xor U1148 (N_1148,In_560,In_425);
nor U1149 (N_1149,In_354,In_20);
nor U1150 (N_1150,In_408,In_138);
nand U1151 (N_1151,In_64,In_452);
nand U1152 (N_1152,In_419,In_328);
nor U1153 (N_1153,In_340,In_585);
and U1154 (N_1154,In_727,In_800);
and U1155 (N_1155,In_99,In_139);
and U1156 (N_1156,In_884,In_818);
nand U1157 (N_1157,In_294,In_624);
xnor U1158 (N_1158,In_640,In_843);
nor U1159 (N_1159,In_921,In_587);
nand U1160 (N_1160,In_219,In_200);
nand U1161 (N_1161,In_491,In_197);
and U1162 (N_1162,In_804,In_209);
nor U1163 (N_1163,In_994,In_546);
nor U1164 (N_1164,In_477,In_769);
xor U1165 (N_1165,In_628,In_874);
and U1166 (N_1166,In_843,In_714);
nor U1167 (N_1167,In_910,In_319);
or U1168 (N_1168,In_765,In_309);
nor U1169 (N_1169,In_230,In_703);
nor U1170 (N_1170,In_671,In_325);
or U1171 (N_1171,In_142,In_757);
and U1172 (N_1172,In_148,In_611);
and U1173 (N_1173,In_876,In_10);
or U1174 (N_1174,In_949,In_207);
and U1175 (N_1175,In_752,In_945);
or U1176 (N_1176,In_876,In_974);
and U1177 (N_1177,In_173,In_69);
nand U1178 (N_1178,In_623,In_420);
nor U1179 (N_1179,In_624,In_215);
or U1180 (N_1180,In_435,In_407);
or U1181 (N_1181,In_13,In_971);
or U1182 (N_1182,In_309,In_109);
nand U1183 (N_1183,In_93,In_833);
nor U1184 (N_1184,In_418,In_616);
nor U1185 (N_1185,In_20,In_321);
nand U1186 (N_1186,In_851,In_980);
nand U1187 (N_1187,In_802,In_138);
nand U1188 (N_1188,In_84,In_264);
nand U1189 (N_1189,In_712,In_545);
nand U1190 (N_1190,In_600,In_129);
xor U1191 (N_1191,In_113,In_539);
nor U1192 (N_1192,In_567,In_65);
nor U1193 (N_1193,In_501,In_977);
and U1194 (N_1194,In_611,In_56);
nor U1195 (N_1195,In_939,In_119);
and U1196 (N_1196,In_180,In_586);
nor U1197 (N_1197,In_983,In_0);
or U1198 (N_1198,In_408,In_920);
nor U1199 (N_1199,In_42,In_519);
xor U1200 (N_1200,In_264,In_135);
nor U1201 (N_1201,In_349,In_982);
nand U1202 (N_1202,In_141,In_529);
xnor U1203 (N_1203,In_113,In_382);
nor U1204 (N_1204,In_711,In_541);
nor U1205 (N_1205,In_914,In_702);
or U1206 (N_1206,In_397,In_746);
or U1207 (N_1207,In_627,In_186);
nor U1208 (N_1208,In_970,In_560);
or U1209 (N_1209,In_783,In_53);
nor U1210 (N_1210,In_475,In_767);
nand U1211 (N_1211,In_42,In_116);
nor U1212 (N_1212,In_410,In_403);
nand U1213 (N_1213,In_29,In_328);
and U1214 (N_1214,In_740,In_766);
or U1215 (N_1215,In_882,In_125);
and U1216 (N_1216,In_678,In_431);
nor U1217 (N_1217,In_348,In_852);
nand U1218 (N_1218,In_826,In_647);
nand U1219 (N_1219,In_247,In_38);
and U1220 (N_1220,In_931,In_411);
nand U1221 (N_1221,In_763,In_4);
nand U1222 (N_1222,In_716,In_414);
nor U1223 (N_1223,In_404,In_636);
and U1224 (N_1224,In_298,In_950);
nand U1225 (N_1225,In_921,In_504);
or U1226 (N_1226,In_851,In_882);
nand U1227 (N_1227,In_250,In_539);
nand U1228 (N_1228,In_694,In_731);
nor U1229 (N_1229,In_871,In_944);
or U1230 (N_1230,In_770,In_443);
nor U1231 (N_1231,In_223,In_62);
and U1232 (N_1232,In_886,In_1);
nand U1233 (N_1233,In_993,In_952);
or U1234 (N_1234,In_217,In_68);
nor U1235 (N_1235,In_466,In_389);
or U1236 (N_1236,In_518,In_326);
or U1237 (N_1237,In_177,In_426);
and U1238 (N_1238,In_558,In_133);
nand U1239 (N_1239,In_723,In_838);
and U1240 (N_1240,In_854,In_978);
and U1241 (N_1241,In_392,In_664);
nand U1242 (N_1242,In_715,In_483);
or U1243 (N_1243,In_542,In_359);
nor U1244 (N_1244,In_129,In_414);
and U1245 (N_1245,In_872,In_716);
nand U1246 (N_1246,In_997,In_257);
nand U1247 (N_1247,In_42,In_30);
and U1248 (N_1248,In_991,In_837);
and U1249 (N_1249,In_772,In_243);
nand U1250 (N_1250,In_845,In_985);
nand U1251 (N_1251,In_501,In_928);
nand U1252 (N_1252,In_773,In_95);
nor U1253 (N_1253,In_538,In_996);
nand U1254 (N_1254,In_697,In_509);
xnor U1255 (N_1255,In_787,In_331);
nor U1256 (N_1256,In_850,In_981);
nor U1257 (N_1257,In_798,In_173);
or U1258 (N_1258,In_277,In_4);
or U1259 (N_1259,In_647,In_357);
and U1260 (N_1260,In_959,In_259);
nor U1261 (N_1261,In_302,In_571);
nor U1262 (N_1262,In_456,In_250);
or U1263 (N_1263,In_895,In_420);
xor U1264 (N_1264,In_282,In_701);
nor U1265 (N_1265,In_398,In_329);
or U1266 (N_1266,In_971,In_571);
and U1267 (N_1267,In_86,In_474);
nor U1268 (N_1268,In_42,In_901);
nor U1269 (N_1269,In_799,In_383);
or U1270 (N_1270,In_276,In_48);
nand U1271 (N_1271,In_366,In_18);
and U1272 (N_1272,In_336,In_828);
and U1273 (N_1273,In_436,In_952);
nand U1274 (N_1274,In_173,In_616);
or U1275 (N_1275,In_216,In_153);
nor U1276 (N_1276,In_75,In_325);
or U1277 (N_1277,In_175,In_184);
and U1278 (N_1278,In_98,In_395);
nand U1279 (N_1279,In_693,In_931);
xor U1280 (N_1280,In_618,In_588);
and U1281 (N_1281,In_406,In_261);
xnor U1282 (N_1282,In_189,In_531);
nand U1283 (N_1283,In_379,In_28);
nand U1284 (N_1284,In_524,In_708);
nor U1285 (N_1285,In_474,In_728);
or U1286 (N_1286,In_198,In_707);
or U1287 (N_1287,In_791,In_413);
and U1288 (N_1288,In_273,In_658);
nor U1289 (N_1289,In_644,In_34);
nor U1290 (N_1290,In_26,In_790);
xor U1291 (N_1291,In_179,In_845);
nor U1292 (N_1292,In_909,In_620);
xnor U1293 (N_1293,In_993,In_0);
xnor U1294 (N_1294,In_611,In_51);
nor U1295 (N_1295,In_451,In_786);
nor U1296 (N_1296,In_546,In_645);
or U1297 (N_1297,In_316,In_842);
or U1298 (N_1298,In_348,In_457);
xor U1299 (N_1299,In_533,In_447);
nand U1300 (N_1300,In_514,In_519);
and U1301 (N_1301,In_979,In_894);
and U1302 (N_1302,In_879,In_535);
and U1303 (N_1303,In_185,In_133);
nand U1304 (N_1304,In_968,In_30);
and U1305 (N_1305,In_478,In_444);
nor U1306 (N_1306,In_449,In_859);
nand U1307 (N_1307,In_612,In_20);
and U1308 (N_1308,In_246,In_406);
nor U1309 (N_1309,In_37,In_885);
nor U1310 (N_1310,In_647,In_636);
nor U1311 (N_1311,In_864,In_213);
and U1312 (N_1312,In_288,In_573);
or U1313 (N_1313,In_497,In_111);
xor U1314 (N_1314,In_57,In_715);
nand U1315 (N_1315,In_117,In_276);
or U1316 (N_1316,In_985,In_520);
nor U1317 (N_1317,In_301,In_935);
nand U1318 (N_1318,In_621,In_262);
nand U1319 (N_1319,In_745,In_215);
and U1320 (N_1320,In_675,In_27);
nor U1321 (N_1321,In_854,In_1);
nand U1322 (N_1322,In_550,In_933);
nor U1323 (N_1323,In_209,In_114);
nand U1324 (N_1324,In_192,In_444);
or U1325 (N_1325,In_19,In_292);
nand U1326 (N_1326,In_99,In_128);
or U1327 (N_1327,In_63,In_879);
nand U1328 (N_1328,In_987,In_874);
nor U1329 (N_1329,In_532,In_984);
or U1330 (N_1330,In_14,In_6);
nor U1331 (N_1331,In_384,In_112);
or U1332 (N_1332,In_918,In_131);
or U1333 (N_1333,In_500,In_147);
nor U1334 (N_1334,In_538,In_15);
or U1335 (N_1335,In_180,In_142);
and U1336 (N_1336,In_167,In_703);
and U1337 (N_1337,In_24,In_465);
xnor U1338 (N_1338,In_984,In_558);
nor U1339 (N_1339,In_398,In_436);
or U1340 (N_1340,In_784,In_450);
nand U1341 (N_1341,In_471,In_352);
nand U1342 (N_1342,In_60,In_204);
and U1343 (N_1343,In_244,In_273);
and U1344 (N_1344,In_198,In_378);
or U1345 (N_1345,In_230,In_153);
and U1346 (N_1346,In_124,In_940);
nand U1347 (N_1347,In_545,In_664);
and U1348 (N_1348,In_789,In_7);
and U1349 (N_1349,In_918,In_633);
or U1350 (N_1350,In_172,In_996);
and U1351 (N_1351,In_483,In_341);
nand U1352 (N_1352,In_310,In_149);
or U1353 (N_1353,In_870,In_312);
and U1354 (N_1354,In_378,In_635);
nand U1355 (N_1355,In_738,In_666);
and U1356 (N_1356,In_405,In_21);
or U1357 (N_1357,In_161,In_241);
or U1358 (N_1358,In_236,In_665);
or U1359 (N_1359,In_419,In_908);
or U1360 (N_1360,In_818,In_199);
nand U1361 (N_1361,In_49,In_738);
or U1362 (N_1362,In_330,In_788);
nand U1363 (N_1363,In_494,In_937);
nor U1364 (N_1364,In_323,In_966);
nor U1365 (N_1365,In_509,In_723);
or U1366 (N_1366,In_510,In_434);
or U1367 (N_1367,In_740,In_559);
nand U1368 (N_1368,In_895,In_181);
nand U1369 (N_1369,In_691,In_228);
or U1370 (N_1370,In_82,In_175);
nand U1371 (N_1371,In_134,In_863);
xnor U1372 (N_1372,In_289,In_719);
and U1373 (N_1373,In_657,In_201);
xnor U1374 (N_1374,In_561,In_94);
xor U1375 (N_1375,In_475,In_551);
xnor U1376 (N_1376,In_759,In_254);
nor U1377 (N_1377,In_95,In_262);
xor U1378 (N_1378,In_585,In_955);
nor U1379 (N_1379,In_710,In_165);
xnor U1380 (N_1380,In_870,In_383);
nand U1381 (N_1381,In_793,In_501);
nand U1382 (N_1382,In_214,In_291);
nand U1383 (N_1383,In_83,In_20);
or U1384 (N_1384,In_164,In_958);
nand U1385 (N_1385,In_932,In_409);
or U1386 (N_1386,In_214,In_69);
nand U1387 (N_1387,In_392,In_683);
and U1388 (N_1388,In_321,In_189);
nor U1389 (N_1389,In_475,In_561);
xor U1390 (N_1390,In_710,In_261);
nor U1391 (N_1391,In_742,In_794);
nor U1392 (N_1392,In_527,In_657);
and U1393 (N_1393,In_734,In_281);
xnor U1394 (N_1394,In_578,In_646);
and U1395 (N_1395,In_17,In_449);
and U1396 (N_1396,In_805,In_513);
nor U1397 (N_1397,In_170,In_677);
and U1398 (N_1398,In_81,In_428);
nor U1399 (N_1399,In_782,In_237);
and U1400 (N_1400,In_68,In_350);
and U1401 (N_1401,In_850,In_29);
nand U1402 (N_1402,In_152,In_425);
or U1403 (N_1403,In_520,In_128);
nor U1404 (N_1404,In_847,In_823);
and U1405 (N_1405,In_958,In_42);
or U1406 (N_1406,In_708,In_444);
nand U1407 (N_1407,In_651,In_82);
or U1408 (N_1408,In_374,In_513);
or U1409 (N_1409,In_43,In_490);
nand U1410 (N_1410,In_355,In_221);
xor U1411 (N_1411,In_108,In_116);
nor U1412 (N_1412,In_89,In_953);
or U1413 (N_1413,In_769,In_750);
nor U1414 (N_1414,In_771,In_848);
or U1415 (N_1415,In_626,In_10);
or U1416 (N_1416,In_429,In_755);
nand U1417 (N_1417,In_880,In_261);
and U1418 (N_1418,In_286,In_162);
or U1419 (N_1419,In_875,In_346);
nor U1420 (N_1420,In_835,In_960);
nand U1421 (N_1421,In_17,In_479);
nand U1422 (N_1422,In_208,In_150);
or U1423 (N_1423,In_319,In_697);
nand U1424 (N_1424,In_582,In_918);
xor U1425 (N_1425,In_280,In_830);
nand U1426 (N_1426,In_648,In_595);
and U1427 (N_1427,In_138,In_263);
nor U1428 (N_1428,In_230,In_500);
and U1429 (N_1429,In_795,In_343);
and U1430 (N_1430,In_841,In_204);
xnor U1431 (N_1431,In_491,In_506);
and U1432 (N_1432,In_155,In_794);
nand U1433 (N_1433,In_690,In_449);
nand U1434 (N_1434,In_321,In_221);
or U1435 (N_1435,In_582,In_849);
nor U1436 (N_1436,In_874,In_886);
nor U1437 (N_1437,In_16,In_830);
and U1438 (N_1438,In_740,In_913);
or U1439 (N_1439,In_354,In_412);
or U1440 (N_1440,In_199,In_767);
nor U1441 (N_1441,In_520,In_892);
and U1442 (N_1442,In_862,In_218);
and U1443 (N_1443,In_45,In_241);
nand U1444 (N_1444,In_915,In_288);
and U1445 (N_1445,In_689,In_709);
and U1446 (N_1446,In_107,In_299);
nand U1447 (N_1447,In_920,In_768);
nand U1448 (N_1448,In_68,In_802);
or U1449 (N_1449,In_612,In_584);
and U1450 (N_1450,In_968,In_439);
or U1451 (N_1451,In_944,In_160);
nand U1452 (N_1452,In_836,In_662);
nor U1453 (N_1453,In_477,In_668);
and U1454 (N_1454,In_405,In_714);
and U1455 (N_1455,In_46,In_443);
nor U1456 (N_1456,In_737,In_553);
nor U1457 (N_1457,In_159,In_649);
xnor U1458 (N_1458,In_645,In_17);
xor U1459 (N_1459,In_724,In_392);
nor U1460 (N_1460,In_592,In_58);
and U1461 (N_1461,In_146,In_556);
nor U1462 (N_1462,In_693,In_103);
or U1463 (N_1463,In_919,In_441);
nor U1464 (N_1464,In_287,In_952);
and U1465 (N_1465,In_455,In_877);
xnor U1466 (N_1466,In_974,In_589);
and U1467 (N_1467,In_57,In_536);
nand U1468 (N_1468,In_885,In_232);
nand U1469 (N_1469,In_977,In_136);
and U1470 (N_1470,In_196,In_478);
or U1471 (N_1471,In_348,In_573);
and U1472 (N_1472,In_689,In_612);
nor U1473 (N_1473,In_932,In_388);
and U1474 (N_1474,In_73,In_237);
nor U1475 (N_1475,In_907,In_754);
xor U1476 (N_1476,In_72,In_848);
and U1477 (N_1477,In_813,In_360);
or U1478 (N_1478,In_470,In_244);
xnor U1479 (N_1479,In_930,In_493);
and U1480 (N_1480,In_684,In_248);
xor U1481 (N_1481,In_516,In_436);
nand U1482 (N_1482,In_139,In_25);
and U1483 (N_1483,In_417,In_1);
or U1484 (N_1484,In_995,In_382);
or U1485 (N_1485,In_762,In_796);
and U1486 (N_1486,In_768,In_799);
and U1487 (N_1487,In_957,In_70);
nand U1488 (N_1488,In_889,In_135);
nand U1489 (N_1489,In_947,In_315);
nand U1490 (N_1490,In_447,In_922);
and U1491 (N_1491,In_643,In_822);
nand U1492 (N_1492,In_722,In_876);
and U1493 (N_1493,In_594,In_887);
and U1494 (N_1494,In_643,In_516);
nand U1495 (N_1495,In_969,In_354);
nand U1496 (N_1496,In_173,In_858);
nand U1497 (N_1497,In_909,In_214);
and U1498 (N_1498,In_354,In_632);
and U1499 (N_1499,In_383,In_474);
and U1500 (N_1500,In_172,In_839);
xor U1501 (N_1501,In_720,In_965);
nor U1502 (N_1502,In_403,In_407);
nand U1503 (N_1503,In_331,In_849);
nor U1504 (N_1504,In_628,In_208);
xor U1505 (N_1505,In_719,In_656);
or U1506 (N_1506,In_182,In_250);
and U1507 (N_1507,In_212,In_310);
or U1508 (N_1508,In_464,In_217);
and U1509 (N_1509,In_567,In_583);
or U1510 (N_1510,In_106,In_718);
and U1511 (N_1511,In_817,In_409);
nor U1512 (N_1512,In_466,In_928);
or U1513 (N_1513,In_151,In_459);
xnor U1514 (N_1514,In_839,In_780);
nand U1515 (N_1515,In_850,In_481);
or U1516 (N_1516,In_709,In_986);
xor U1517 (N_1517,In_94,In_385);
nand U1518 (N_1518,In_896,In_868);
nor U1519 (N_1519,In_316,In_850);
or U1520 (N_1520,In_186,In_800);
xnor U1521 (N_1521,In_977,In_256);
or U1522 (N_1522,In_903,In_573);
nor U1523 (N_1523,In_964,In_932);
or U1524 (N_1524,In_143,In_700);
or U1525 (N_1525,In_28,In_68);
or U1526 (N_1526,In_84,In_810);
and U1527 (N_1527,In_369,In_875);
nor U1528 (N_1528,In_840,In_689);
and U1529 (N_1529,In_387,In_362);
or U1530 (N_1530,In_117,In_209);
nand U1531 (N_1531,In_435,In_762);
nor U1532 (N_1532,In_182,In_173);
or U1533 (N_1533,In_25,In_459);
xnor U1534 (N_1534,In_595,In_634);
nand U1535 (N_1535,In_841,In_736);
and U1536 (N_1536,In_556,In_158);
or U1537 (N_1537,In_900,In_336);
or U1538 (N_1538,In_702,In_102);
nand U1539 (N_1539,In_62,In_402);
or U1540 (N_1540,In_685,In_8);
and U1541 (N_1541,In_711,In_989);
and U1542 (N_1542,In_976,In_376);
nand U1543 (N_1543,In_277,In_168);
or U1544 (N_1544,In_277,In_597);
nor U1545 (N_1545,In_729,In_287);
nor U1546 (N_1546,In_817,In_304);
nand U1547 (N_1547,In_288,In_927);
or U1548 (N_1548,In_644,In_606);
xor U1549 (N_1549,In_852,In_432);
and U1550 (N_1550,In_383,In_488);
or U1551 (N_1551,In_568,In_699);
nand U1552 (N_1552,In_228,In_484);
and U1553 (N_1553,In_419,In_483);
nand U1554 (N_1554,In_134,In_806);
and U1555 (N_1555,In_711,In_702);
xor U1556 (N_1556,In_810,In_5);
and U1557 (N_1557,In_344,In_944);
or U1558 (N_1558,In_322,In_89);
or U1559 (N_1559,In_536,In_306);
nand U1560 (N_1560,In_735,In_619);
xnor U1561 (N_1561,In_725,In_241);
nor U1562 (N_1562,In_658,In_222);
and U1563 (N_1563,In_281,In_388);
or U1564 (N_1564,In_183,In_255);
and U1565 (N_1565,In_865,In_300);
nor U1566 (N_1566,In_911,In_792);
nand U1567 (N_1567,In_617,In_847);
nand U1568 (N_1568,In_68,In_741);
or U1569 (N_1569,In_789,In_389);
or U1570 (N_1570,In_449,In_801);
nand U1571 (N_1571,In_674,In_611);
nor U1572 (N_1572,In_755,In_3);
or U1573 (N_1573,In_435,In_202);
and U1574 (N_1574,In_321,In_537);
xnor U1575 (N_1575,In_361,In_385);
nor U1576 (N_1576,In_900,In_838);
nor U1577 (N_1577,In_344,In_119);
and U1578 (N_1578,In_483,In_418);
nand U1579 (N_1579,In_102,In_778);
nand U1580 (N_1580,In_894,In_498);
or U1581 (N_1581,In_800,In_690);
xnor U1582 (N_1582,In_619,In_40);
or U1583 (N_1583,In_744,In_874);
nor U1584 (N_1584,In_919,In_870);
and U1585 (N_1585,In_231,In_160);
nand U1586 (N_1586,In_932,In_243);
nand U1587 (N_1587,In_375,In_849);
xor U1588 (N_1588,In_261,In_903);
nand U1589 (N_1589,In_225,In_393);
or U1590 (N_1590,In_398,In_824);
and U1591 (N_1591,In_332,In_992);
or U1592 (N_1592,In_175,In_802);
xnor U1593 (N_1593,In_173,In_579);
and U1594 (N_1594,In_849,In_590);
nand U1595 (N_1595,In_130,In_342);
and U1596 (N_1596,In_935,In_794);
nand U1597 (N_1597,In_596,In_746);
nor U1598 (N_1598,In_249,In_866);
nor U1599 (N_1599,In_525,In_253);
nand U1600 (N_1600,In_342,In_323);
and U1601 (N_1601,In_199,In_580);
nor U1602 (N_1602,In_857,In_98);
or U1603 (N_1603,In_221,In_648);
or U1604 (N_1604,In_494,In_130);
nand U1605 (N_1605,In_704,In_231);
and U1606 (N_1606,In_568,In_67);
and U1607 (N_1607,In_314,In_480);
or U1608 (N_1608,In_135,In_287);
or U1609 (N_1609,In_74,In_736);
and U1610 (N_1610,In_792,In_165);
and U1611 (N_1611,In_257,In_270);
or U1612 (N_1612,In_936,In_647);
or U1613 (N_1613,In_986,In_327);
and U1614 (N_1614,In_814,In_494);
nand U1615 (N_1615,In_377,In_435);
and U1616 (N_1616,In_446,In_25);
and U1617 (N_1617,In_309,In_55);
nor U1618 (N_1618,In_497,In_267);
or U1619 (N_1619,In_331,In_550);
or U1620 (N_1620,In_48,In_747);
nor U1621 (N_1621,In_2,In_546);
nor U1622 (N_1622,In_554,In_603);
and U1623 (N_1623,In_642,In_410);
nor U1624 (N_1624,In_668,In_900);
nor U1625 (N_1625,In_353,In_403);
and U1626 (N_1626,In_127,In_189);
or U1627 (N_1627,In_177,In_793);
nand U1628 (N_1628,In_671,In_269);
nand U1629 (N_1629,In_525,In_566);
or U1630 (N_1630,In_7,In_486);
nand U1631 (N_1631,In_150,In_462);
nand U1632 (N_1632,In_260,In_884);
or U1633 (N_1633,In_688,In_546);
or U1634 (N_1634,In_816,In_88);
or U1635 (N_1635,In_657,In_59);
or U1636 (N_1636,In_777,In_499);
and U1637 (N_1637,In_97,In_308);
or U1638 (N_1638,In_644,In_397);
and U1639 (N_1639,In_940,In_907);
xnor U1640 (N_1640,In_289,In_186);
nor U1641 (N_1641,In_299,In_316);
or U1642 (N_1642,In_875,In_76);
and U1643 (N_1643,In_938,In_681);
or U1644 (N_1644,In_259,In_572);
nand U1645 (N_1645,In_256,In_680);
nand U1646 (N_1646,In_406,In_956);
nand U1647 (N_1647,In_153,In_552);
or U1648 (N_1648,In_444,In_135);
nand U1649 (N_1649,In_491,In_645);
nand U1650 (N_1650,In_864,In_456);
nand U1651 (N_1651,In_56,In_511);
or U1652 (N_1652,In_699,In_203);
nor U1653 (N_1653,In_591,In_7);
nor U1654 (N_1654,In_297,In_403);
nand U1655 (N_1655,In_228,In_740);
or U1656 (N_1656,In_296,In_919);
or U1657 (N_1657,In_595,In_67);
and U1658 (N_1658,In_533,In_433);
nor U1659 (N_1659,In_224,In_34);
nor U1660 (N_1660,In_249,In_559);
nor U1661 (N_1661,In_685,In_624);
nor U1662 (N_1662,In_626,In_863);
nor U1663 (N_1663,In_965,In_64);
nor U1664 (N_1664,In_652,In_261);
nand U1665 (N_1665,In_223,In_421);
or U1666 (N_1666,In_798,In_449);
xor U1667 (N_1667,In_205,In_44);
nor U1668 (N_1668,In_490,In_349);
or U1669 (N_1669,In_659,In_535);
xor U1670 (N_1670,In_984,In_904);
or U1671 (N_1671,In_831,In_265);
or U1672 (N_1672,In_981,In_625);
nor U1673 (N_1673,In_875,In_16);
xor U1674 (N_1674,In_104,In_443);
nand U1675 (N_1675,In_24,In_911);
or U1676 (N_1676,In_85,In_439);
or U1677 (N_1677,In_380,In_59);
and U1678 (N_1678,In_489,In_930);
or U1679 (N_1679,In_766,In_178);
nor U1680 (N_1680,In_407,In_851);
or U1681 (N_1681,In_625,In_177);
xnor U1682 (N_1682,In_936,In_224);
and U1683 (N_1683,In_171,In_435);
nand U1684 (N_1684,In_347,In_346);
and U1685 (N_1685,In_958,In_41);
nor U1686 (N_1686,In_258,In_604);
or U1687 (N_1687,In_192,In_805);
or U1688 (N_1688,In_568,In_274);
and U1689 (N_1689,In_505,In_807);
or U1690 (N_1690,In_358,In_120);
or U1691 (N_1691,In_151,In_521);
or U1692 (N_1692,In_739,In_904);
nand U1693 (N_1693,In_702,In_596);
nor U1694 (N_1694,In_674,In_949);
nor U1695 (N_1695,In_373,In_897);
or U1696 (N_1696,In_996,In_613);
nand U1697 (N_1697,In_2,In_489);
nand U1698 (N_1698,In_1,In_476);
and U1699 (N_1699,In_493,In_68);
and U1700 (N_1700,In_118,In_244);
and U1701 (N_1701,In_903,In_470);
and U1702 (N_1702,In_136,In_319);
nor U1703 (N_1703,In_144,In_836);
and U1704 (N_1704,In_780,In_856);
nor U1705 (N_1705,In_719,In_984);
or U1706 (N_1706,In_629,In_254);
nand U1707 (N_1707,In_132,In_217);
nand U1708 (N_1708,In_474,In_541);
or U1709 (N_1709,In_623,In_658);
and U1710 (N_1710,In_39,In_19);
xor U1711 (N_1711,In_536,In_423);
nand U1712 (N_1712,In_487,In_414);
and U1713 (N_1713,In_546,In_371);
and U1714 (N_1714,In_574,In_153);
and U1715 (N_1715,In_659,In_102);
and U1716 (N_1716,In_823,In_305);
and U1717 (N_1717,In_581,In_601);
nand U1718 (N_1718,In_205,In_490);
nand U1719 (N_1719,In_935,In_942);
nand U1720 (N_1720,In_740,In_348);
or U1721 (N_1721,In_44,In_772);
nand U1722 (N_1722,In_145,In_349);
and U1723 (N_1723,In_858,In_204);
nor U1724 (N_1724,In_600,In_690);
and U1725 (N_1725,In_109,In_52);
xnor U1726 (N_1726,In_923,In_447);
nand U1727 (N_1727,In_221,In_808);
and U1728 (N_1728,In_730,In_905);
nor U1729 (N_1729,In_872,In_512);
nand U1730 (N_1730,In_546,In_969);
nor U1731 (N_1731,In_80,In_136);
nand U1732 (N_1732,In_179,In_565);
or U1733 (N_1733,In_327,In_329);
nor U1734 (N_1734,In_483,In_455);
nand U1735 (N_1735,In_990,In_708);
nor U1736 (N_1736,In_21,In_291);
or U1737 (N_1737,In_247,In_854);
and U1738 (N_1738,In_155,In_228);
nand U1739 (N_1739,In_650,In_382);
xnor U1740 (N_1740,In_728,In_880);
nand U1741 (N_1741,In_547,In_444);
xnor U1742 (N_1742,In_751,In_587);
or U1743 (N_1743,In_588,In_146);
and U1744 (N_1744,In_716,In_730);
xor U1745 (N_1745,In_43,In_457);
nand U1746 (N_1746,In_377,In_446);
nand U1747 (N_1747,In_673,In_879);
and U1748 (N_1748,In_14,In_3);
nand U1749 (N_1749,In_437,In_52);
xnor U1750 (N_1750,In_594,In_492);
nand U1751 (N_1751,In_674,In_420);
nand U1752 (N_1752,In_690,In_837);
and U1753 (N_1753,In_215,In_594);
nor U1754 (N_1754,In_800,In_426);
or U1755 (N_1755,In_330,In_76);
nor U1756 (N_1756,In_3,In_223);
or U1757 (N_1757,In_136,In_463);
and U1758 (N_1758,In_613,In_181);
xnor U1759 (N_1759,In_422,In_618);
nor U1760 (N_1760,In_698,In_22);
and U1761 (N_1761,In_47,In_720);
nor U1762 (N_1762,In_123,In_499);
nand U1763 (N_1763,In_743,In_340);
or U1764 (N_1764,In_155,In_78);
and U1765 (N_1765,In_136,In_73);
or U1766 (N_1766,In_8,In_855);
nand U1767 (N_1767,In_867,In_357);
or U1768 (N_1768,In_469,In_979);
xor U1769 (N_1769,In_272,In_495);
nor U1770 (N_1770,In_130,In_536);
nor U1771 (N_1771,In_684,In_765);
nand U1772 (N_1772,In_907,In_560);
or U1773 (N_1773,In_986,In_216);
nor U1774 (N_1774,In_577,In_152);
nor U1775 (N_1775,In_297,In_470);
and U1776 (N_1776,In_770,In_432);
nor U1777 (N_1777,In_98,In_441);
nand U1778 (N_1778,In_379,In_881);
nand U1779 (N_1779,In_561,In_833);
nor U1780 (N_1780,In_646,In_292);
and U1781 (N_1781,In_933,In_469);
nand U1782 (N_1782,In_395,In_869);
nor U1783 (N_1783,In_76,In_339);
or U1784 (N_1784,In_224,In_119);
nor U1785 (N_1785,In_486,In_761);
or U1786 (N_1786,In_791,In_783);
nor U1787 (N_1787,In_584,In_168);
xnor U1788 (N_1788,In_250,In_658);
or U1789 (N_1789,In_17,In_159);
nor U1790 (N_1790,In_440,In_290);
and U1791 (N_1791,In_149,In_978);
or U1792 (N_1792,In_530,In_696);
or U1793 (N_1793,In_99,In_208);
and U1794 (N_1794,In_88,In_348);
or U1795 (N_1795,In_303,In_254);
or U1796 (N_1796,In_917,In_25);
or U1797 (N_1797,In_289,In_905);
nor U1798 (N_1798,In_947,In_674);
nand U1799 (N_1799,In_133,In_548);
nand U1800 (N_1800,In_926,In_164);
and U1801 (N_1801,In_307,In_537);
nand U1802 (N_1802,In_485,In_426);
nand U1803 (N_1803,In_139,In_811);
nand U1804 (N_1804,In_789,In_335);
or U1805 (N_1805,In_597,In_414);
or U1806 (N_1806,In_39,In_133);
nor U1807 (N_1807,In_500,In_775);
or U1808 (N_1808,In_596,In_768);
nand U1809 (N_1809,In_303,In_109);
nor U1810 (N_1810,In_152,In_215);
nor U1811 (N_1811,In_163,In_262);
or U1812 (N_1812,In_100,In_698);
nand U1813 (N_1813,In_355,In_665);
and U1814 (N_1814,In_597,In_376);
nor U1815 (N_1815,In_975,In_521);
nor U1816 (N_1816,In_609,In_423);
nand U1817 (N_1817,In_382,In_61);
nor U1818 (N_1818,In_386,In_233);
and U1819 (N_1819,In_268,In_337);
or U1820 (N_1820,In_208,In_512);
nand U1821 (N_1821,In_969,In_173);
nand U1822 (N_1822,In_848,In_233);
nor U1823 (N_1823,In_430,In_752);
and U1824 (N_1824,In_710,In_825);
nor U1825 (N_1825,In_711,In_169);
and U1826 (N_1826,In_277,In_571);
or U1827 (N_1827,In_292,In_895);
or U1828 (N_1828,In_139,In_971);
xnor U1829 (N_1829,In_510,In_268);
nor U1830 (N_1830,In_102,In_814);
xnor U1831 (N_1831,In_710,In_514);
nand U1832 (N_1832,In_396,In_550);
and U1833 (N_1833,In_560,In_684);
xnor U1834 (N_1834,In_602,In_196);
or U1835 (N_1835,In_752,In_938);
and U1836 (N_1836,In_636,In_734);
nor U1837 (N_1837,In_112,In_273);
nor U1838 (N_1838,In_587,In_157);
nand U1839 (N_1839,In_453,In_676);
nor U1840 (N_1840,In_61,In_995);
or U1841 (N_1841,In_998,In_984);
xnor U1842 (N_1842,In_222,In_625);
and U1843 (N_1843,In_803,In_67);
or U1844 (N_1844,In_289,In_304);
xnor U1845 (N_1845,In_52,In_195);
nand U1846 (N_1846,In_888,In_362);
and U1847 (N_1847,In_524,In_891);
xor U1848 (N_1848,In_225,In_775);
xor U1849 (N_1849,In_569,In_82);
nor U1850 (N_1850,In_76,In_305);
nor U1851 (N_1851,In_647,In_375);
and U1852 (N_1852,In_8,In_383);
or U1853 (N_1853,In_834,In_453);
nor U1854 (N_1854,In_895,In_357);
xnor U1855 (N_1855,In_882,In_419);
nor U1856 (N_1856,In_921,In_179);
and U1857 (N_1857,In_46,In_703);
nor U1858 (N_1858,In_205,In_513);
nand U1859 (N_1859,In_993,In_635);
and U1860 (N_1860,In_5,In_995);
and U1861 (N_1861,In_876,In_168);
and U1862 (N_1862,In_388,In_377);
nor U1863 (N_1863,In_740,In_649);
xor U1864 (N_1864,In_900,In_688);
nand U1865 (N_1865,In_732,In_828);
nor U1866 (N_1866,In_711,In_310);
or U1867 (N_1867,In_482,In_306);
or U1868 (N_1868,In_117,In_215);
or U1869 (N_1869,In_751,In_25);
nor U1870 (N_1870,In_653,In_16);
nor U1871 (N_1871,In_208,In_559);
or U1872 (N_1872,In_153,In_46);
or U1873 (N_1873,In_270,In_233);
xnor U1874 (N_1874,In_567,In_318);
and U1875 (N_1875,In_29,In_758);
and U1876 (N_1876,In_34,In_234);
and U1877 (N_1877,In_926,In_298);
nand U1878 (N_1878,In_901,In_407);
or U1879 (N_1879,In_499,In_44);
or U1880 (N_1880,In_995,In_526);
and U1881 (N_1881,In_701,In_690);
nor U1882 (N_1882,In_972,In_607);
nor U1883 (N_1883,In_527,In_685);
nand U1884 (N_1884,In_575,In_422);
or U1885 (N_1885,In_89,In_765);
nand U1886 (N_1886,In_584,In_666);
nor U1887 (N_1887,In_922,In_66);
nor U1888 (N_1888,In_191,In_923);
or U1889 (N_1889,In_232,In_226);
and U1890 (N_1890,In_805,In_124);
or U1891 (N_1891,In_156,In_16);
and U1892 (N_1892,In_667,In_609);
xor U1893 (N_1893,In_48,In_528);
nand U1894 (N_1894,In_257,In_950);
nor U1895 (N_1895,In_663,In_393);
nand U1896 (N_1896,In_45,In_160);
nor U1897 (N_1897,In_873,In_355);
nand U1898 (N_1898,In_125,In_260);
and U1899 (N_1899,In_363,In_297);
or U1900 (N_1900,In_179,In_20);
nor U1901 (N_1901,In_144,In_15);
nor U1902 (N_1902,In_797,In_126);
nand U1903 (N_1903,In_252,In_177);
xor U1904 (N_1904,In_329,In_93);
xnor U1905 (N_1905,In_452,In_753);
xnor U1906 (N_1906,In_267,In_41);
nand U1907 (N_1907,In_803,In_126);
nor U1908 (N_1908,In_197,In_181);
nand U1909 (N_1909,In_230,In_231);
nand U1910 (N_1910,In_838,In_391);
nor U1911 (N_1911,In_679,In_92);
or U1912 (N_1912,In_281,In_112);
and U1913 (N_1913,In_585,In_952);
nor U1914 (N_1914,In_626,In_209);
xnor U1915 (N_1915,In_12,In_612);
and U1916 (N_1916,In_676,In_812);
nand U1917 (N_1917,In_927,In_477);
and U1918 (N_1918,In_33,In_277);
xor U1919 (N_1919,In_830,In_116);
and U1920 (N_1920,In_820,In_638);
nor U1921 (N_1921,In_665,In_370);
nor U1922 (N_1922,In_327,In_923);
nand U1923 (N_1923,In_398,In_117);
nand U1924 (N_1924,In_36,In_118);
xor U1925 (N_1925,In_758,In_649);
nor U1926 (N_1926,In_715,In_102);
nor U1927 (N_1927,In_23,In_383);
nand U1928 (N_1928,In_434,In_110);
or U1929 (N_1929,In_537,In_488);
and U1930 (N_1930,In_673,In_981);
and U1931 (N_1931,In_598,In_398);
nand U1932 (N_1932,In_660,In_812);
nor U1933 (N_1933,In_114,In_260);
nand U1934 (N_1934,In_614,In_388);
nor U1935 (N_1935,In_344,In_481);
or U1936 (N_1936,In_878,In_881);
or U1937 (N_1937,In_456,In_598);
nor U1938 (N_1938,In_971,In_698);
or U1939 (N_1939,In_214,In_617);
nor U1940 (N_1940,In_188,In_88);
or U1941 (N_1941,In_1,In_577);
xnor U1942 (N_1942,In_339,In_302);
and U1943 (N_1943,In_195,In_839);
and U1944 (N_1944,In_165,In_127);
nand U1945 (N_1945,In_703,In_536);
or U1946 (N_1946,In_381,In_944);
nor U1947 (N_1947,In_406,In_730);
nor U1948 (N_1948,In_265,In_989);
nor U1949 (N_1949,In_998,In_327);
xnor U1950 (N_1950,In_71,In_908);
nor U1951 (N_1951,In_163,In_52);
nor U1952 (N_1952,In_663,In_948);
or U1953 (N_1953,In_350,In_368);
nor U1954 (N_1954,In_468,In_926);
nand U1955 (N_1955,In_555,In_388);
xor U1956 (N_1956,In_692,In_164);
and U1957 (N_1957,In_668,In_853);
xnor U1958 (N_1958,In_400,In_179);
and U1959 (N_1959,In_944,In_637);
and U1960 (N_1960,In_407,In_130);
nor U1961 (N_1961,In_864,In_112);
xnor U1962 (N_1962,In_941,In_150);
or U1963 (N_1963,In_30,In_870);
nor U1964 (N_1964,In_544,In_381);
xor U1965 (N_1965,In_432,In_150);
nor U1966 (N_1966,In_905,In_292);
and U1967 (N_1967,In_459,In_820);
or U1968 (N_1968,In_387,In_785);
nand U1969 (N_1969,In_61,In_732);
or U1970 (N_1970,In_765,In_241);
xor U1971 (N_1971,In_860,In_458);
nand U1972 (N_1972,In_953,In_104);
and U1973 (N_1973,In_955,In_518);
nand U1974 (N_1974,In_186,In_70);
nand U1975 (N_1975,In_110,In_356);
and U1976 (N_1976,In_271,In_44);
or U1977 (N_1977,In_873,In_421);
and U1978 (N_1978,In_190,In_257);
nand U1979 (N_1979,In_668,In_271);
nor U1980 (N_1980,In_412,In_915);
and U1981 (N_1981,In_973,In_109);
xnor U1982 (N_1982,In_817,In_81);
or U1983 (N_1983,In_123,In_393);
nand U1984 (N_1984,In_397,In_801);
nand U1985 (N_1985,In_71,In_151);
nor U1986 (N_1986,In_333,In_389);
nor U1987 (N_1987,In_913,In_123);
or U1988 (N_1988,In_201,In_180);
nand U1989 (N_1989,In_243,In_340);
nor U1990 (N_1990,In_740,In_927);
and U1991 (N_1991,In_112,In_92);
and U1992 (N_1992,In_792,In_660);
nand U1993 (N_1993,In_902,In_634);
nand U1994 (N_1994,In_66,In_95);
nand U1995 (N_1995,In_287,In_594);
nand U1996 (N_1996,In_142,In_189);
and U1997 (N_1997,In_356,In_438);
or U1998 (N_1998,In_331,In_226);
or U1999 (N_1999,In_213,In_658);
nor U2000 (N_2000,N_1976,N_1395);
nand U2001 (N_2001,N_1329,N_1300);
or U2002 (N_2002,N_424,N_1954);
nor U2003 (N_2003,N_1002,N_307);
and U2004 (N_2004,N_324,N_1853);
or U2005 (N_2005,N_636,N_794);
and U2006 (N_2006,N_360,N_449);
nor U2007 (N_2007,N_1647,N_1104);
or U2008 (N_2008,N_1009,N_1092);
nor U2009 (N_2009,N_1906,N_18);
nor U2010 (N_2010,N_1271,N_1877);
and U2011 (N_2011,N_202,N_1607);
nand U2012 (N_2012,N_291,N_1953);
and U2013 (N_2013,N_1677,N_1416);
nand U2014 (N_2014,N_438,N_1943);
or U2015 (N_2015,N_1094,N_597);
or U2016 (N_2016,N_1926,N_1999);
or U2017 (N_2017,N_1590,N_1553);
and U2018 (N_2018,N_394,N_1156);
or U2019 (N_2019,N_404,N_1628);
xor U2020 (N_2020,N_172,N_669);
or U2021 (N_2021,N_1806,N_119);
or U2022 (N_2022,N_417,N_906);
nor U2023 (N_2023,N_1511,N_405);
xnor U2024 (N_2024,N_414,N_816);
nor U2025 (N_2025,N_1202,N_335);
and U2026 (N_2026,N_317,N_1440);
nor U2027 (N_2027,N_470,N_370);
and U2028 (N_2028,N_1059,N_365);
xnor U2029 (N_2029,N_1579,N_1205);
or U2030 (N_2030,N_1472,N_1606);
nand U2031 (N_2031,N_440,N_259);
nor U2032 (N_2032,N_384,N_252);
nand U2033 (N_2033,N_843,N_1675);
and U2034 (N_2034,N_1324,N_618);
nor U2035 (N_2035,N_1846,N_1214);
nor U2036 (N_2036,N_1354,N_1130);
and U2037 (N_2037,N_631,N_1405);
or U2038 (N_2038,N_61,N_81);
and U2039 (N_2039,N_1198,N_982);
and U2040 (N_2040,N_1701,N_1162);
or U2041 (N_2041,N_277,N_645);
nor U2042 (N_2042,N_1680,N_1077);
nand U2043 (N_2043,N_1805,N_528);
nor U2044 (N_2044,N_443,N_1698);
nor U2045 (N_2045,N_34,N_1688);
or U2046 (N_2046,N_1802,N_1950);
or U2047 (N_2047,N_1133,N_1598);
nand U2048 (N_2048,N_879,N_664);
and U2049 (N_2049,N_1718,N_552);
and U2050 (N_2050,N_500,N_894);
or U2051 (N_2051,N_125,N_1321);
and U2052 (N_2052,N_181,N_1140);
nand U2053 (N_2053,N_817,N_605);
nand U2054 (N_2054,N_1213,N_1549);
and U2055 (N_2055,N_459,N_434);
nand U2056 (N_2056,N_1621,N_355);
nand U2057 (N_2057,N_1111,N_256);
nand U2058 (N_2058,N_1128,N_1801);
and U2059 (N_2059,N_1792,N_1959);
or U2060 (N_2060,N_1945,N_1282);
nand U2061 (N_2061,N_1871,N_1005);
nand U2062 (N_2062,N_680,N_1572);
nand U2063 (N_2063,N_427,N_1931);
or U2064 (N_2064,N_1020,N_677);
and U2065 (N_2065,N_1050,N_1866);
and U2066 (N_2066,N_1061,N_1479);
and U2067 (N_2067,N_1824,N_574);
xnor U2068 (N_2068,N_1788,N_17);
nor U2069 (N_2069,N_850,N_344);
and U2070 (N_2070,N_1990,N_849);
nand U2071 (N_2071,N_1979,N_1619);
or U2072 (N_2072,N_1671,N_863);
and U2073 (N_2073,N_1304,N_1905);
or U2074 (N_2074,N_872,N_798);
or U2075 (N_2075,N_1836,N_1466);
nand U2076 (N_2076,N_1091,N_474);
nand U2077 (N_2077,N_1759,N_1225);
or U2078 (N_2078,N_1316,N_924);
or U2079 (N_2079,N_473,N_38);
or U2080 (N_2080,N_1042,N_1392);
nor U2081 (N_2081,N_829,N_28);
nor U2082 (N_2082,N_1046,N_758);
and U2083 (N_2083,N_547,N_316);
nor U2084 (N_2084,N_1052,N_1192);
or U2085 (N_2085,N_1770,N_1443);
or U2086 (N_2086,N_766,N_604);
and U2087 (N_2087,N_951,N_1276);
nor U2088 (N_2088,N_1022,N_838);
nand U2089 (N_2089,N_1885,N_1404);
nand U2090 (N_2090,N_1844,N_388);
xor U2091 (N_2091,N_1429,N_1894);
and U2092 (N_2092,N_908,N_1177);
or U2093 (N_2093,N_1408,N_841);
xnor U2094 (N_2094,N_1571,N_1922);
nor U2095 (N_2095,N_1068,N_313);
or U2096 (N_2096,N_331,N_925);
nand U2097 (N_2097,N_1123,N_936);
or U2098 (N_2098,N_1311,N_1856);
nand U2099 (N_2099,N_1141,N_1346);
nor U2100 (N_2100,N_88,N_1882);
nand U2101 (N_2101,N_646,N_1188);
and U2102 (N_2102,N_1437,N_379);
nor U2103 (N_2103,N_147,N_840);
and U2104 (N_2104,N_1411,N_897);
and U2105 (N_2105,N_1608,N_251);
nor U2106 (N_2106,N_1576,N_134);
or U2107 (N_2107,N_804,N_1204);
nand U2108 (N_2108,N_1886,N_1758);
nand U2109 (N_2109,N_114,N_1021);
nand U2110 (N_2110,N_1656,N_1626);
and U2111 (N_2111,N_156,N_272);
nand U2112 (N_2112,N_1632,N_511);
nand U2113 (N_2113,N_1870,N_898);
nand U2114 (N_2114,N_382,N_609);
nor U2115 (N_2115,N_284,N_40);
xor U2116 (N_2116,N_42,N_146);
and U2117 (N_2117,N_1266,N_1654);
or U2118 (N_2118,N_989,N_1262);
and U2119 (N_2119,N_654,N_662);
nor U2120 (N_2120,N_1872,N_702);
nor U2121 (N_2121,N_108,N_1107);
nand U2122 (N_2122,N_1224,N_594);
and U2123 (N_2123,N_1791,N_561);
nor U2124 (N_2124,N_1365,N_1461);
nor U2125 (N_2125,N_1536,N_647);
and U2126 (N_2126,N_1138,N_1315);
and U2127 (N_2127,N_705,N_764);
nor U2128 (N_2128,N_1843,N_1566);
nand U2129 (N_2129,N_1968,N_948);
xnor U2130 (N_2130,N_1881,N_682);
or U2131 (N_2131,N_1024,N_615);
xnor U2132 (N_2132,N_32,N_1822);
nand U2133 (N_2133,N_1575,N_1557);
nand U2134 (N_2134,N_550,N_1232);
and U2135 (N_2135,N_448,N_1391);
and U2136 (N_2136,N_1124,N_423);
xnor U2137 (N_2137,N_1089,N_493);
nand U2138 (N_2138,N_1977,N_1384);
or U2139 (N_2139,N_1027,N_701);
and U2140 (N_2140,N_825,N_782);
or U2141 (N_2141,N_929,N_299);
and U2142 (N_2142,N_488,N_189);
xor U2143 (N_2143,N_1119,N_278);
and U2144 (N_2144,N_1927,N_1980);
xor U2145 (N_2145,N_1003,N_1746);
nand U2146 (N_2146,N_868,N_821);
and U2147 (N_2147,N_1431,N_1957);
nand U2148 (N_2148,N_942,N_322);
xnor U2149 (N_2149,N_985,N_120);
xor U2150 (N_2150,N_1339,N_328);
nand U2151 (N_2151,N_45,N_1070);
xor U2152 (N_2152,N_1064,N_1804);
and U2153 (N_2153,N_1149,N_1716);
nor U2154 (N_2154,N_1229,N_191);
xnor U2155 (N_2155,N_1006,N_1246);
nand U2156 (N_2156,N_1817,N_455);
nand U2157 (N_2157,N_625,N_740);
or U2158 (N_2158,N_551,N_1412);
nand U2159 (N_2159,N_602,N_1764);
and U2160 (N_2160,N_1051,N_544);
and U2161 (N_2161,N_707,N_915);
nor U2162 (N_2162,N_1900,N_1397);
or U2163 (N_2163,N_1389,N_1150);
nor U2164 (N_2164,N_1651,N_236);
nor U2165 (N_2165,N_1994,N_1908);
and U2166 (N_2166,N_787,N_1497);
nand U2167 (N_2167,N_1490,N_772);
or U2168 (N_2168,N_1396,N_1445);
nor U2169 (N_2169,N_1215,N_1447);
or U2170 (N_2170,N_52,N_484);
nand U2171 (N_2171,N_506,N_1249);
nand U2172 (N_2172,N_1962,N_1096);
or U2173 (N_2173,N_651,N_1823);
and U2174 (N_2174,N_1142,N_1880);
nand U2175 (N_2175,N_1893,N_973);
nand U2176 (N_2176,N_391,N_1310);
and U2177 (N_2177,N_864,N_1136);
nor U2178 (N_2178,N_1060,N_1206);
or U2179 (N_2179,N_1101,N_472);
xnor U2180 (N_2180,N_714,N_763);
xor U2181 (N_2181,N_161,N_454);
nand U2182 (N_2182,N_1,N_805);
nor U2183 (N_2183,N_856,N_140);
or U2184 (N_2184,N_958,N_652);
xor U2185 (N_2185,N_1784,N_537);
and U2186 (N_2186,N_392,N_212);
nand U2187 (N_2187,N_1648,N_741);
or U2188 (N_2188,N_835,N_318);
nor U2189 (N_2189,N_1196,N_436);
xor U2190 (N_2190,N_409,N_1255);
nand U2191 (N_2191,N_72,N_781);
nor U2192 (N_2192,N_304,N_347);
and U2193 (N_2193,N_1373,N_293);
nor U2194 (N_2194,N_188,N_681);
nand U2195 (N_2195,N_1679,N_1295);
and U2196 (N_2196,N_6,N_1627);
and U2197 (N_2197,N_575,N_1997);
nor U2198 (N_2198,N_1018,N_1505);
nand U2199 (N_2199,N_1251,N_412);
nand U2200 (N_2200,N_1735,N_716);
and U2201 (N_2201,N_730,N_329);
nor U2202 (N_2202,N_1669,N_131);
or U2203 (N_2203,N_1040,N_683);
xnor U2204 (N_2204,N_1121,N_200);
nand U2205 (N_2205,N_503,N_854);
nor U2206 (N_2206,N_1813,N_1201);
nand U2207 (N_2207,N_47,N_803);
or U2208 (N_2208,N_234,N_1768);
nor U2209 (N_2209,N_1819,N_800);
or U2210 (N_2210,N_230,N_11);
xnor U2211 (N_2211,N_1564,N_532);
nor U2212 (N_2212,N_1293,N_938);
or U2213 (N_2213,N_1643,N_797);
and U2214 (N_2214,N_1892,N_1114);
or U2215 (N_2215,N_378,N_877);
nand U2216 (N_2216,N_1936,N_396);
nor U2217 (N_2217,N_1137,N_784);
and U2218 (N_2218,N_1793,N_1666);
xor U2219 (N_2219,N_921,N_214);
and U2220 (N_2220,N_1631,N_599);
or U2221 (N_2221,N_1269,N_495);
or U2222 (N_2222,N_1219,N_576);
or U2223 (N_2223,N_1151,N_1122);
nand U2224 (N_2224,N_1974,N_1973);
nand U2225 (N_2225,N_1868,N_1341);
nor U2226 (N_2226,N_157,N_795);
or U2227 (N_2227,N_1694,N_524);
or U2228 (N_2228,N_1848,N_1320);
or U2229 (N_2229,N_1025,N_1949);
nand U2230 (N_2230,N_1102,N_853);
or U2231 (N_2231,N_1630,N_97);
nand U2232 (N_2232,N_546,N_289);
nor U2233 (N_2233,N_954,N_1812);
and U2234 (N_2234,N_1387,N_295);
and U2235 (N_2235,N_306,N_588);
nand U2236 (N_2236,N_1786,N_1659);
nor U2237 (N_2237,N_1487,N_1363);
xnor U2238 (N_2238,N_567,N_545);
xor U2239 (N_2239,N_1896,N_1076);
and U2240 (N_2240,N_676,N_731);
or U2241 (N_2241,N_1292,N_219);
nor U2242 (N_2242,N_1664,N_762);
and U2243 (N_2243,N_1538,N_1991);
nor U2244 (N_2244,N_240,N_321);
and U2245 (N_2245,N_19,N_279);
nand U2246 (N_2246,N_29,N_1134);
nand U2247 (N_2247,N_628,N_859);
or U2248 (N_2248,N_1542,N_811);
nor U2249 (N_2249,N_1525,N_1634);
and U2250 (N_2250,N_24,N_889);
or U2251 (N_2251,N_606,N_658);
xor U2252 (N_2252,N_1017,N_1482);
or U2253 (N_2253,N_1705,N_1235);
nor U2254 (N_2254,N_1272,N_325);
nand U2255 (N_2255,N_1724,N_198);
nor U2256 (N_2256,N_49,N_1589);
and U2257 (N_2257,N_880,N_1855);
nand U2258 (N_2258,N_261,N_708);
nand U2259 (N_2259,N_1448,N_337);
and U2260 (N_2260,N_1842,N_584);
or U2261 (N_2261,N_96,N_1280);
and U2262 (N_2262,N_1139,N_1955);
nor U2263 (N_2263,N_1738,N_1257);
or U2264 (N_2264,N_80,N_1725);
and U2265 (N_2265,N_142,N_1851);
nand U2266 (N_2266,N_678,N_1222);
nand U2267 (N_2267,N_243,N_640);
and U2268 (N_2268,N_1030,N_1930);
xnor U2269 (N_2269,N_1182,N_266);
nand U2270 (N_2270,N_903,N_182);
or U2271 (N_2271,N_1984,N_287);
and U2272 (N_2272,N_1723,N_100);
and U2273 (N_2273,N_31,N_1921);
and U2274 (N_2274,N_1620,N_1008);
or U2275 (N_2275,N_888,N_608);
nor U2276 (N_2276,N_151,N_920);
xor U2277 (N_2277,N_1432,N_1722);
nor U2278 (N_2278,N_1960,N_184);
or U2279 (N_2279,N_23,N_1147);
or U2280 (N_2280,N_376,N_1670);
nor U2281 (N_2281,N_523,N_1638);
or U2282 (N_2282,N_463,N_861);
and U2283 (N_2283,N_1661,N_1840);
and U2284 (N_2284,N_264,N_559);
nor U2285 (N_2285,N_1709,N_959);
nor U2286 (N_2286,N_1739,N_673);
or U2287 (N_2287,N_381,N_1495);
xnor U2288 (N_2288,N_1889,N_1803);
nor U2289 (N_2289,N_356,N_1464);
nand U2290 (N_2290,N_1504,N_696);
and U2291 (N_2291,N_649,N_916);
nand U2292 (N_2292,N_1517,N_1285);
nand U2293 (N_2293,N_1037,N_1995);
and U2294 (N_2294,N_927,N_59);
or U2295 (N_2295,N_1586,N_112);
xnor U2296 (N_2296,N_1034,N_534);
nor U2297 (N_2297,N_1286,N_536);
nand U2298 (N_2298,N_499,N_565);
or U2299 (N_2299,N_878,N_1938);
xnor U2300 (N_2300,N_441,N_1043);
or U2301 (N_2301,N_456,N_1992);
or U2302 (N_2302,N_380,N_1486);
xnor U2303 (N_2303,N_1820,N_719);
and U2304 (N_2304,N_22,N_826);
or U2305 (N_2305,N_1345,N_1928);
nor U2306 (N_2306,N_1712,N_922);
or U2307 (N_2307,N_896,N_1703);
nand U2308 (N_2308,N_870,N_1736);
and U2309 (N_2309,N_407,N_890);
nand U2310 (N_2310,N_1941,N_1260);
or U2311 (N_2311,N_1583,N_1001);
nor U2312 (N_2312,N_1166,N_519);
and U2313 (N_2313,N_1299,N_1655);
or U2314 (N_2314,N_8,N_312);
nor U2315 (N_2315,N_866,N_1580);
nand U2316 (N_2316,N_1766,N_660);
nand U2317 (N_2317,N_887,N_242);
nor U2318 (N_2318,N_783,N_1312);
nand U2319 (N_2319,N_892,N_1875);
and U2320 (N_2320,N_1985,N_976);
xnor U2321 (N_2321,N_93,N_1132);
xor U2322 (N_2322,N_192,N_15);
and U2323 (N_2323,N_1609,N_290);
and U2324 (N_2324,N_904,N_1438);
nand U2325 (N_2325,N_509,N_1967);
or U2326 (N_2326,N_458,N_148);
xor U2327 (N_2327,N_748,N_471);
nand U2328 (N_2328,N_756,N_209);
nand U2329 (N_2329,N_1406,N_997);
xnor U2330 (N_2330,N_1965,N_1987);
or U2331 (N_2331,N_196,N_1158);
and U2332 (N_2332,N_1217,N_250);
nor U2333 (N_2333,N_1650,N_375);
nor U2334 (N_2334,N_637,N_398);
and U2335 (N_2335,N_1765,N_641);
nor U2336 (N_2336,N_13,N_1665);
nand U2337 (N_2337,N_822,N_1367);
and U2338 (N_2338,N_1263,N_1728);
nor U2339 (N_2339,N_258,N_420);
nand U2340 (N_2340,N_358,N_1131);
nand U2341 (N_2341,N_1568,N_132);
and U2342 (N_2342,N_453,N_1611);
nor U2343 (N_2343,N_1774,N_127);
or U2344 (N_2344,N_1435,N_865);
nor U2345 (N_2345,N_1357,N_1242);
nand U2346 (N_2346,N_170,N_1210);
nor U2347 (N_2347,N_847,N_186);
nor U2348 (N_2348,N_1809,N_178);
xor U2349 (N_2349,N_1072,N_768);
nand U2350 (N_2350,N_1763,N_226);
or U2351 (N_2351,N_1852,N_1913);
nor U2352 (N_2352,N_590,N_1494);
nand U2353 (N_2353,N_1831,N_229);
xor U2354 (N_2354,N_1605,N_773);
and U2355 (N_2355,N_679,N_928);
nor U2356 (N_2356,N_400,N_167);
or U2357 (N_2357,N_1097,N_1704);
nor U2358 (N_2358,N_1358,N_508);
nor U2359 (N_2359,N_43,N_1993);
nor U2360 (N_2360,N_1452,N_1524);
or U2361 (N_2361,N_1773,N_244);
nor U2362 (N_2362,N_207,N_1622);
nor U2363 (N_2363,N_1612,N_642);
and U2364 (N_2364,N_1279,N_109);
or U2365 (N_2365,N_944,N_978);
nor U2366 (N_2366,N_340,N_1693);
nand U2367 (N_2367,N_891,N_227);
and U2368 (N_2368,N_674,N_1436);
and U2369 (N_2369,N_1811,N_268);
nor U2370 (N_2370,N_1625,N_724);
or U2371 (N_2371,N_273,N_1808);
or U2372 (N_2372,N_387,N_468);
or U2373 (N_2373,N_1939,N_369);
and U2374 (N_2374,N_943,N_1932);
nor U2375 (N_2375,N_419,N_1471);
nand U2376 (N_2376,N_1729,N_933);
and U2377 (N_2377,N_1283,N_1468);
and U2378 (N_2378,N_1543,N_1732);
nand U2379 (N_2379,N_1398,N_1726);
xnor U2380 (N_2380,N_1143,N_2);
nor U2381 (N_2381,N_1244,N_962);
and U2382 (N_2382,N_479,N_999);
nor U2383 (N_2383,N_1377,N_839);
nor U2384 (N_2384,N_477,N_1434);
and U2385 (N_2385,N_217,N_64);
or U2386 (N_2386,N_1390,N_504);
nand U2387 (N_2387,N_1423,N_187);
nor U2388 (N_2388,N_812,N_1287);
nor U2389 (N_2389,N_54,N_1569);
xor U2390 (N_2390,N_1252,N_969);
nand U2391 (N_2391,N_1417,N_815);
or U2392 (N_2392,N_1761,N_1193);
nor U2393 (N_2393,N_342,N_1830);
nand U2394 (N_2394,N_981,N_1332);
nand U2395 (N_2395,N_314,N_739);
and U2396 (N_2396,N_1236,N_1319);
nand U2397 (N_2397,N_239,N_1212);
nand U2398 (N_2398,N_1449,N_1530);
or U2399 (N_2399,N_1640,N_1573);
nand U2400 (N_2400,N_1327,N_1845);
nor U2401 (N_2401,N_931,N_1223);
or U2402 (N_2402,N_1488,N_700);
nand U2403 (N_2403,N_778,N_1883);
or U2404 (N_2404,N_1364,N_498);
nor U2405 (N_2405,N_648,N_518);
and U2406 (N_2406,N_1053,N_1270);
and U2407 (N_2407,N_326,N_505);
nand U2408 (N_2408,N_834,N_1424);
or U2409 (N_2409,N_276,N_1646);
or U2410 (N_2410,N_153,N_623);
nand U2411 (N_2411,N_502,N_1103);
or U2412 (N_2412,N_1935,N_308);
nand U2413 (N_2413,N_957,N_1597);
nand U2414 (N_2414,N_949,N_558);
and U2415 (N_2415,N_900,N_1409);
nand U2416 (N_2416,N_1787,N_809);
or U2417 (N_2417,N_1307,N_411);
nor U2418 (N_2418,N_848,N_752);
nand U2419 (N_2419,N_1228,N_1189);
and U2420 (N_2420,N_1190,N_1642);
and U2421 (N_2421,N_712,N_213);
nor U2422 (N_2422,N_672,N_661);
or U2423 (N_2423,N_422,N_1873);
or U2424 (N_2424,N_1918,N_837);
or U2425 (N_2425,N_457,N_1869);
or U2426 (N_2426,N_1847,N_1057);
nand U2427 (N_2427,N_667,N_726);
and U2428 (N_2428,N_934,N_1144);
or U2429 (N_2429,N_338,N_1233);
nor U2430 (N_2430,N_1989,N_123);
or U2431 (N_2431,N_1220,N_1988);
and U2432 (N_2432,N_699,N_1617);
nor U2433 (N_2433,N_1506,N_1983);
or U2434 (N_2434,N_201,N_84);
xnor U2435 (N_2435,N_1273,N_332);
or U2436 (N_2436,N_624,N_1035);
or U2437 (N_2437,N_1187,N_195);
and U2438 (N_2438,N_531,N_1169);
nor U2439 (N_2439,N_1998,N_190);
nand U2440 (N_2440,N_1159,N_1737);
nand U2441 (N_2441,N_445,N_1155);
and U2442 (N_2442,N_1054,N_1231);
or U2443 (N_2443,N_246,N_432);
and U2444 (N_2444,N_53,N_136);
and U2445 (N_2445,N_431,N_452);
nor U2446 (N_2446,N_1668,N_377);
and U2447 (N_2447,N_1972,N_738);
or U2448 (N_2448,N_1065,N_1457);
nand U2449 (N_2449,N_1306,N_1115);
and U2450 (N_2450,N_1278,N_901);
nand U2451 (N_2451,N_155,N_571);
or U2452 (N_2452,N_885,N_1828);
nand U2453 (N_2453,N_1523,N_397);
or U2454 (N_2454,N_610,N_1721);
nor U2455 (N_2455,N_1129,N_1769);
nand U2456 (N_2456,N_543,N_1775);
nor U2457 (N_2457,N_496,N_257);
and U2458 (N_2458,N_361,N_1301);
nor U2459 (N_2459,N_447,N_1550);
nand U2460 (N_2460,N_77,N_1561);
nor U2461 (N_2461,N_248,N_255);
nand U2462 (N_2462,N_115,N_1393);
and U2463 (N_2463,N_851,N_1240);
nor U2464 (N_2464,N_106,N_830);
and U2465 (N_2465,N_1860,N_56);
or U2466 (N_2466,N_1481,N_1760);
nor U2467 (N_2467,N_633,N_1167);
or U2468 (N_2468,N_50,N_1850);
or U2469 (N_2469,N_1499,N_165);
nand U2470 (N_2470,N_1399,N_729);
and U2471 (N_2471,N_621,N_1816);
or U2472 (N_2472,N_749,N_1510);
nor U2473 (N_2473,N_1522,N_1385);
nand U2474 (N_2474,N_1195,N_1917);
nand U2475 (N_2475,N_844,N_698);
or U2476 (N_2476,N_1199,N_1164);
or U2477 (N_2477,N_983,N_1925);
or U2478 (N_2478,N_1857,N_1474);
nand U2479 (N_2479,N_7,N_1541);
nand U2480 (N_2480,N_1653,N_1082);
nand U2481 (N_2481,N_1682,N_1016);
nor U2482 (N_2482,N_385,N_33);
nand U2483 (N_2483,N_1599,N_1975);
nand U2484 (N_2484,N_302,N_1776);
or U2485 (N_2485,N_1191,N_1800);
nand U2486 (N_2486,N_1734,N_1343);
and U2487 (N_2487,N_296,N_1088);
nor U2488 (N_2488,N_223,N_1372);
nor U2489 (N_2489,N_746,N_1378);
nor U2490 (N_2490,N_1298,N_1075);
or U2491 (N_2491,N_952,N_930);
and U2492 (N_2492,N_911,N_94);
nor U2493 (N_2493,N_323,N_1366);
or U2494 (N_2494,N_320,N_267);
nor U2495 (N_2495,N_245,N_171);
nand U2496 (N_2496,N_1827,N_941);
nor U2497 (N_2497,N_1422,N_1551);
nand U2498 (N_2498,N_1208,N_715);
and U2499 (N_2499,N_1982,N_1426);
nand U2500 (N_2500,N_105,N_695);
nor U2501 (N_2501,N_1717,N_912);
or U2502 (N_2502,N_704,N_595);
nor U2503 (N_2503,N_1558,N_1044);
nor U2504 (N_2504,N_1218,N_1326);
and U2505 (N_2505,N_1243,N_393);
and U2506 (N_2506,N_305,N_725);
and U2507 (N_2507,N_970,N_1610);
and U2508 (N_2508,N_937,N_1313);
nor U2509 (N_2509,N_126,N_1731);
nor U2510 (N_2510,N_288,N_1920);
nor U2511 (N_2511,N_1157,N_285);
or U2512 (N_2512,N_280,N_692);
and U2513 (N_2513,N_540,N_1335);
or U2514 (N_2514,N_855,N_910);
nand U2515 (N_2515,N_55,N_1507);
or U2516 (N_2516,N_1261,N_237);
nand U2517 (N_2517,N_1078,N_1601);
nor U2518 (N_2518,N_1618,N_1676);
and U2519 (N_2519,N_600,N_1095);
or U2520 (N_2520,N_294,N_845);
and U2521 (N_2521,N_1083,N_644);
and U2522 (N_2522,N_1349,N_241);
nor U2523 (N_2523,N_1779,N_1032);
nor U2524 (N_2524,N_1200,N_953);
xor U2525 (N_2525,N_1446,N_1689);
nor U2526 (N_2526,N_814,N_1649);
nand U2527 (N_2527,N_566,N_1267);
or U2528 (N_2528,N_1197,N_601);
and U2529 (N_2529,N_150,N_1839);
nand U2530 (N_2530,N_83,N_1433);
nand U2531 (N_2531,N_1713,N_733);
and U2532 (N_2532,N_919,N_1532);
xnor U2533 (N_2533,N_1259,N_286);
nand U2534 (N_2534,N_485,N_582);
and U2535 (N_2535,N_410,N_465);
nor U2536 (N_2536,N_1031,N_1864);
and U2537 (N_2537,N_1480,N_1117);
nand U2538 (N_2538,N_1000,N_1207);
or U2539 (N_2539,N_1832,N_1170);
and U2540 (N_2540,N_1012,N_706);
and U2541 (N_2541,N_852,N_1028);
nor U2542 (N_2542,N_691,N_75);
or U2543 (N_2543,N_104,N_963);
nor U2544 (N_2544,N_1745,N_124);
and U2545 (N_2545,N_1891,N_1547);
or U2546 (N_2546,N_1227,N_1248);
nor U2547 (N_2547,N_1386,N_282);
and U2548 (N_2548,N_556,N_775);
and U2549 (N_2549,N_233,N_476);
or U2550 (N_2550,N_179,N_501);
nand U2551 (N_2551,N_693,N_685);
and U2552 (N_2552,N_330,N_770);
and U2553 (N_2553,N_1498,N_1370);
and U2554 (N_2554,N_204,N_406);
nand U2555 (N_2555,N_359,N_1662);
nor U2556 (N_2556,N_1578,N_907);
xor U2557 (N_2557,N_1264,N_1780);
and U2558 (N_2558,N_1814,N_371);
nor U2559 (N_2559,N_389,N_1374);
nand U2560 (N_2560,N_205,N_1355);
or U2561 (N_2561,N_857,N_1749);
or U2562 (N_2562,N_1347,N_51);
nor U2563 (N_2563,N_996,N_767);
and U2564 (N_2564,N_1552,N_806);
nand U2565 (N_2565,N_1458,N_122);
or U2566 (N_2566,N_1593,N_1318);
nand U2567 (N_2567,N_310,N_833);
and U2568 (N_2568,N_1148,N_668);
nand U2569 (N_2569,N_617,N_16);
nor U2570 (N_2570,N_966,N_1879);
nor U2571 (N_2571,N_1742,N_1838);
nor U2572 (N_2572,N_364,N_1952);
nor U2573 (N_2573,N_1258,N_1833);
and U2574 (N_2574,N_643,N_598);
and U2575 (N_2575,N_158,N_1862);
xor U2576 (N_2576,N_1767,N_629);
and U2577 (N_2577,N_1039,N_1508);
nand U2578 (N_2578,N_1520,N_79);
or U2579 (N_2579,N_569,N_1348);
or U2580 (N_2580,N_1184,N_1041);
nand U2581 (N_2581,N_1407,N_1923);
nand U2582 (N_2582,N_281,N_1544);
nor U2583 (N_2583,N_1577,N_627);
or U2584 (N_2584,N_1069,N_639);
nand U2585 (N_2585,N_1582,N_152);
nor U2586 (N_2586,N_987,N_215);
and U2587 (N_2587,N_352,N_1080);
xnor U2588 (N_2588,N_408,N_1352);
or U2589 (N_2589,N_1265,N_1441);
or U2590 (N_2590,N_1465,N_274);
nand U2591 (N_2591,N_221,N_1777);
and U2592 (N_2592,N_1789,N_1485);
or U2593 (N_2593,N_492,N_228);
and U2594 (N_2594,N_607,N_67);
nor U2595 (N_2595,N_914,N_875);
nand U2596 (N_2596,N_1691,N_428);
nor U2597 (N_2597,N_101,N_1567);
or U2598 (N_2598,N_353,N_1106);
nand U2599 (N_2599,N_975,N_166);
or U2600 (N_2600,N_656,N_1183);
or U2601 (N_2601,N_1719,N_1360);
and U2602 (N_2602,N_1160,N_977);
or U2603 (N_2603,N_58,N_1528);
nand U2604 (N_2604,N_137,N_357);
and U2605 (N_2605,N_1849,N_1337);
or U2606 (N_2606,N_1478,N_1535);
nor U2607 (N_2607,N_1684,N_858);
and U2608 (N_2608,N_1369,N_1708);
nor U2609 (N_2609,N_538,N_703);
nor U2610 (N_2610,N_717,N_1587);
nor U2611 (N_2611,N_961,N_1540);
or U2612 (N_2612,N_1496,N_632);
xnor U2613 (N_2613,N_1451,N_1146);
or U2614 (N_2614,N_1074,N_1116);
or U2615 (N_2615,N_1686,N_521);
xor U2616 (N_2616,N_947,N_298);
nor U2617 (N_2617,N_1476,N_1375);
nor U2618 (N_2618,N_1442,N_659);
xor U2619 (N_2619,N_1048,N_247);
nor U2620 (N_2620,N_450,N_139);
or U2621 (N_2621,N_66,N_1026);
nor U2622 (N_2622,N_655,N_1942);
and U2623 (N_2623,N_254,N_1067);
or U2624 (N_2624,N_950,N_1221);
nand U2625 (N_2625,N_1644,N_1516);
or U2626 (N_2626,N_751,N_1834);
xnor U2627 (N_2627,N_995,N_301);
nor U2628 (N_2628,N_1818,N_222);
and U2629 (N_2629,N_765,N_1081);
nor U2630 (N_2630,N_591,N_899);
xnor U2631 (N_2631,N_1038,N_1956);
nor U2632 (N_2632,N_334,N_596);
and U2633 (N_2633,N_1518,N_886);
and U2634 (N_2634,N_494,N_1477);
nand U2635 (N_2635,N_1029,N_1254);
and U2636 (N_2636,N_742,N_554);
xnor U2637 (N_2637,N_177,N_1047);
or U2638 (N_2638,N_82,N_1376);
and U2639 (N_2639,N_1344,N_1785);
and U2640 (N_2640,N_27,N_1033);
nor U2641 (N_2641,N_1179,N_620);
or U2642 (N_2642,N_354,N_1751);
and U2643 (N_2643,N_1066,N_39);
nor U2644 (N_2644,N_1268,N_1328);
and U2645 (N_2645,N_555,N_3);
and U2646 (N_2646,N_98,N_709);
and U2647 (N_2647,N_786,N_1795);
or U2648 (N_2648,N_1013,N_46);
or U2649 (N_2649,N_1604,N_759);
and U2650 (N_2650,N_1695,N_1602);
xnor U2651 (N_2651,N_734,N_1570);
and U2652 (N_2652,N_1874,N_789);
and U2653 (N_2653,N_721,N_1010);
nand U2654 (N_2654,N_1629,N_128);
nor U2655 (N_2655,N_510,N_1902);
nand U2656 (N_2656,N_1173,N_1624);
nor U2657 (N_2657,N_578,N_1176);
or U2658 (N_2658,N_718,N_535);
and U2659 (N_2659,N_1308,N_1475);
nand U2660 (N_2660,N_372,N_1049);
or U2661 (N_2661,N_1555,N_180);
nand U2662 (N_2662,N_686,N_208);
and U2663 (N_2663,N_827,N_231);
and U2664 (N_2664,N_174,N_429);
nor U2665 (N_2665,N_1019,N_1290);
or U2666 (N_2666,N_143,N_902);
and U2667 (N_2667,N_36,N_1211);
and U2668 (N_2668,N_1460,N_713);
and U2669 (N_2669,N_1165,N_622);
or U2670 (N_2670,N_444,N_95);
and U2671 (N_2671,N_1418,N_1172);
or U2672 (N_2672,N_1623,N_41);
nand U2673 (N_2673,N_203,N_1450);
and U2674 (N_2674,N_1782,N_144);
or U2675 (N_2675,N_73,N_1388);
nor U2676 (N_2676,N_743,N_1519);
or U2677 (N_2677,N_819,N_1401);
or U2678 (N_2678,N_1898,N_1685);
nor U2679 (N_2679,N_583,N_439);
or U2680 (N_2680,N_1175,N_1534);
and U2681 (N_2681,N_832,N_199);
nand U2682 (N_2682,N_1331,N_1294);
nand U2683 (N_2683,N_1382,N_587);
nor U2684 (N_2684,N_1916,N_1752);
nor U2685 (N_2685,N_253,N_489);
nand U2686 (N_2686,N_1645,N_1559);
and U2687 (N_2687,N_194,N_390);
nand U2688 (N_2688,N_30,N_593);
or U2689 (N_2689,N_37,N_761);
or U2690 (N_2690,N_336,N_1512);
or U2691 (N_2691,N_665,N_882);
nand U2692 (N_2692,N_138,N_670);
nand U2693 (N_2693,N_1565,N_283);
nand U2694 (N_2694,N_589,N_1730);
nor U2695 (N_2695,N_1289,N_1161);
or U2696 (N_2696,N_1757,N_1539);
xnor U2697 (N_2697,N_1230,N_309);
nor U2698 (N_2698,N_1297,N_1585);
xnor U2699 (N_2699,N_613,N_614);
nand U2700 (N_2700,N_1772,N_1934);
xnor U2701 (N_2701,N_1109,N_548);
nor U2702 (N_2702,N_568,N_1821);
nand U2703 (N_2703,N_527,N_824);
nor U2704 (N_2704,N_1904,N_619);
nor U2705 (N_2705,N_260,N_1702);
and U2706 (N_2706,N_133,N_998);
and U2707 (N_2707,N_1314,N_168);
or U2708 (N_2708,N_1641,N_1484);
or U2709 (N_2709,N_430,N_1740);
and U2710 (N_2710,N_684,N_1733);
nor U2711 (N_2711,N_1178,N_1798);
nor U2712 (N_2712,N_1673,N_1914);
nor U2713 (N_2713,N_932,N_69);
or U2714 (N_2714,N_141,N_224);
nand U2715 (N_2715,N_1402,N_225);
nor U2716 (N_2716,N_1174,N_481);
and U2717 (N_2717,N_1581,N_657);
or U2718 (N_2718,N_533,N_1216);
nand U2719 (N_2719,N_1678,N_1023);
and U2720 (N_2720,N_480,N_1239);
nor U2721 (N_2721,N_831,N_363);
xor U2722 (N_2722,N_1521,N_514);
and U2723 (N_2723,N_792,N_270);
xnor U2724 (N_2724,N_1556,N_1841);
nor U2725 (N_2725,N_99,N_1720);
or U2726 (N_2726,N_339,N_415);
xor U2727 (N_2727,N_269,N_1897);
nand U2728 (N_2728,N_820,N_560);
nand U2729 (N_2729,N_1444,N_754);
nand U2730 (N_2730,N_1783,N_349);
or U2731 (N_2731,N_413,N_711);
or U2732 (N_2732,N_1087,N_1706);
xor U2733 (N_2733,N_1837,N_1185);
or U2734 (N_2734,N_1924,N_373);
nor U2735 (N_2735,N_1981,N_1303);
and U2736 (N_2736,N_490,N_1062);
nor U2737 (N_2737,N_984,N_1186);
nand U2738 (N_2738,N_1861,N_1501);
nand U2739 (N_2739,N_926,N_1359);
nand U2740 (N_2740,N_416,N_842);
nor U2741 (N_2741,N_1910,N_483);
or U2742 (N_2742,N_1929,N_884);
and U2743 (N_2743,N_175,N_909);
nor U2744 (N_2744,N_65,N_1615);
nand U2745 (N_2745,N_1241,N_163);
and U2746 (N_2746,N_160,N_522);
and U2747 (N_2747,N_635,N_327);
nor U2748 (N_2748,N_1015,N_1529);
xor U2749 (N_2749,N_62,N_791);
nand U2750 (N_2750,N_1500,N_913);
xor U2751 (N_2751,N_968,N_777);
or U2752 (N_2752,N_442,N_249);
nor U2753 (N_2753,N_333,N_1696);
nor U2754 (N_2754,N_1014,N_727);
nand U2755 (N_2755,N_722,N_362);
nor U2756 (N_2756,N_516,N_1108);
nand U2757 (N_2757,N_1493,N_1086);
or U2758 (N_2758,N_1410,N_1697);
or U2759 (N_2759,N_1700,N_1807);
or U2760 (N_2760,N_1381,N_1379);
xnor U2761 (N_2761,N_211,N_585);
xor U2762 (N_2762,N_1888,N_1058);
xnor U2763 (N_2763,N_1755,N_1428);
or U2764 (N_2764,N_116,N_1652);
nor U2765 (N_2765,N_1063,N_1120);
nand U2766 (N_2766,N_1011,N_799);
nor U2767 (N_2767,N_1637,N_808);
nand U2768 (N_2768,N_1907,N_426);
nor U2769 (N_2769,N_1978,N_1361);
xor U2770 (N_2770,N_881,N_1778);
and U2771 (N_2771,N_235,N_1546);
or U2772 (N_2772,N_451,N_1098);
nand U2773 (N_2773,N_580,N_111);
or U2774 (N_2774,N_1325,N_1986);
and U2775 (N_2775,N_745,N_1815);
nand U2776 (N_2776,N_1462,N_1951);
nand U2777 (N_2777,N_1933,N_5);
or U2778 (N_2778,N_1899,N_802);
xnor U2779 (N_2779,N_1351,N_1635);
nand U2780 (N_2780,N_1790,N_1548);
xor U2781 (N_2781,N_1045,N_873);
nor U2782 (N_2782,N_343,N_1284);
xor U2783 (N_2783,N_63,N_1455);
nand U2784 (N_2784,N_303,N_20);
nor U2785 (N_2785,N_1394,N_1658);
nor U2786 (N_2786,N_736,N_586);
and U2787 (N_2787,N_1171,N_1085);
and U2788 (N_2788,N_57,N_630);
and U2789 (N_2789,N_818,N_1383);
xnor U2790 (N_2790,N_1453,N_723);
nand U2791 (N_2791,N_1425,N_539);
nand U2792 (N_2792,N_1560,N_292);
nand U2793 (N_2793,N_1715,N_1594);
and U2794 (N_2794,N_1209,N_232);
nand U2795 (N_2795,N_1469,N_867);
and U2796 (N_2796,N_1247,N_35);
nor U2797 (N_2797,N_271,N_464);
and U2798 (N_2798,N_1826,N_9);
and U2799 (N_2799,N_1463,N_1663);
nand U2800 (N_2800,N_68,N_507);
nor U2801 (N_2801,N_796,N_1591);
nand U2802 (N_2802,N_1274,N_1911);
nor U2803 (N_2803,N_846,N_418);
or U2804 (N_2804,N_1614,N_1071);
or U2805 (N_2805,N_612,N_44);
and U2806 (N_2806,N_1636,N_395);
or U2807 (N_2807,N_836,N_1413);
xnor U2808 (N_2808,N_1825,N_1657);
and U2809 (N_2809,N_1537,N_1887);
nand U2810 (N_2810,N_366,N_421);
nor U2811 (N_2811,N_520,N_433);
nor U2812 (N_2812,N_769,N_570);
and U2813 (N_2813,N_486,N_1090);
nor U2814 (N_2814,N_1439,N_1036);
nand U2815 (N_2815,N_70,N_960);
nand U2816 (N_2816,N_577,N_1305);
or U2817 (N_2817,N_563,N_1683);
and U2818 (N_2818,N_1163,N_460);
and U2819 (N_2819,N_1194,N_118);
nand U2820 (N_2820,N_1747,N_1302);
nor U2821 (N_2821,N_10,N_1256);
and U2822 (N_2822,N_1753,N_0);
nand U2823 (N_2823,N_1592,N_694);
or U2824 (N_2824,N_810,N_103);
or U2825 (N_2825,N_1459,N_579);
and U2826 (N_2826,N_1333,N_1362);
or U2827 (N_2827,N_1711,N_530);
or U2828 (N_2828,N_1687,N_1353);
nand U2829 (N_2829,N_650,N_399);
xnor U2830 (N_2830,N_1859,N_581);
and U2831 (N_2831,N_785,N_1296);
nor U2832 (N_2832,N_1513,N_1168);
nand U2833 (N_2833,N_76,N_48);
nand U2834 (N_2834,N_60,N_1154);
nand U2835 (N_2835,N_974,N_687);
or U2836 (N_2836,N_1963,N_755);
or U2837 (N_2837,N_1181,N_1901);
and U2838 (N_2838,N_1100,N_1356);
nor U2839 (N_2839,N_1858,N_1110);
or U2840 (N_2840,N_801,N_462);
nor U2841 (N_2841,N_1944,N_350);
nor U2842 (N_2842,N_671,N_697);
xor U2843 (N_2843,N_1867,N_262);
nor U2844 (N_2844,N_1470,N_159);
nor U2845 (N_2845,N_1509,N_979);
and U2846 (N_2846,N_346,N_1554);
or U2847 (N_2847,N_1368,N_220);
or U2848 (N_2848,N_525,N_666);
nor U2849 (N_2849,N_25,N_297);
nor U2850 (N_2850,N_1756,N_1180);
nand U2851 (N_2851,N_21,N_1699);
nor U2852 (N_2852,N_1771,N_1961);
nand U2853 (N_2853,N_774,N_780);
and U2854 (N_2854,N_1126,N_149);
or U2855 (N_2855,N_1613,N_92);
xnor U2856 (N_2856,N_1692,N_779);
or U2857 (N_2857,N_517,N_402);
nand U2858 (N_2858,N_1503,N_1084);
nor U2859 (N_2859,N_437,N_1492);
and U2860 (N_2860,N_1562,N_1421);
xor U2861 (N_2861,N_348,N_980);
xnor U2862 (N_2862,N_1969,N_1714);
nand U2863 (N_2863,N_939,N_176);
or U2864 (N_2864,N_1794,N_102);
and U2865 (N_2865,N_690,N_1674);
nor U2866 (N_2866,N_813,N_341);
nor U2867 (N_2867,N_515,N_760);
nand U2868 (N_2868,N_967,N_1113);
nand U2869 (N_2869,N_611,N_1633);
nand U2870 (N_2870,N_541,N_1419);
or U2871 (N_2871,N_757,N_964);
nand U2872 (N_2872,N_1342,N_991);
xnor U2873 (N_2873,N_946,N_871);
and U2874 (N_2874,N_1489,N_1810);
and U2875 (N_2875,N_1741,N_1350);
or U2876 (N_2876,N_1563,N_869);
nand U2877 (N_2877,N_562,N_988);
nor U2878 (N_2878,N_368,N_1754);
and U2879 (N_2879,N_592,N_1380);
xor U2880 (N_2880,N_573,N_497);
or U2881 (N_2881,N_1797,N_1309);
xor U2882 (N_2882,N_1336,N_1152);
nor U2883 (N_2883,N_956,N_572);
nand U2884 (N_2884,N_965,N_1890);
nor U2885 (N_2885,N_874,N_807);
and U2886 (N_2886,N_689,N_1796);
nor U2887 (N_2887,N_737,N_162);
xnor U2888 (N_2888,N_164,N_403);
or U2889 (N_2889,N_1835,N_720);
or U2890 (N_2890,N_1964,N_1415);
or U2891 (N_2891,N_1884,N_1600);
and U2892 (N_2892,N_1291,N_86);
or U2893 (N_2893,N_1946,N_1727);
or U2894 (N_2894,N_1127,N_173);
and U2895 (N_2895,N_1744,N_993);
nor U2896 (N_2896,N_1514,N_529);
nand U2897 (N_2897,N_1596,N_435);
nand U2898 (N_2898,N_557,N_1322);
nand U2899 (N_2899,N_553,N_1533);
nand U2900 (N_2900,N_793,N_1330);
and U2901 (N_2901,N_1903,N_26);
or U2902 (N_2902,N_1234,N_776);
or U2903 (N_2903,N_771,N_1710);
and U2904 (N_2904,N_185,N_1996);
xnor U2905 (N_2905,N_940,N_750);
and U2906 (N_2906,N_1427,N_549);
nor U2907 (N_2907,N_1966,N_345);
nor U2908 (N_2908,N_110,N_1237);
nand U2909 (N_2909,N_383,N_1588);
nand U2910 (N_2910,N_482,N_1245);
or U2911 (N_2911,N_945,N_828);
and U2912 (N_2912,N_401,N_1004);
or U2913 (N_2913,N_1750,N_564);
xor U2914 (N_2914,N_1958,N_1672);
or U2915 (N_2915,N_300,N_917);
and U2916 (N_2916,N_1371,N_107);
nor U2917 (N_2917,N_1403,N_425);
xor U2918 (N_2918,N_1603,N_790);
nand U2919 (N_2919,N_315,N_1919);
or U2920 (N_2920,N_923,N_735);
and U2921 (N_2921,N_1912,N_1574);
nand U2922 (N_2922,N_1948,N_513);
and U2923 (N_2923,N_1105,N_1940);
nor U2924 (N_2924,N_1502,N_1203);
xor U2925 (N_2925,N_1681,N_1527);
and U2926 (N_2926,N_1531,N_1863);
nor U2927 (N_2927,N_895,N_992);
and U2928 (N_2928,N_275,N_1135);
nand U2929 (N_2929,N_1584,N_1454);
and U2930 (N_2930,N_265,N_87);
and U2931 (N_2931,N_918,N_1056);
nor U2932 (N_2932,N_117,N_183);
nand U2933 (N_2933,N_1483,N_634);
or U2934 (N_2934,N_626,N_467);
nor U2935 (N_2935,N_971,N_603);
and U2936 (N_2936,N_972,N_238);
nand U2937 (N_2937,N_1250,N_1829);
and U2938 (N_2938,N_1854,N_130);
or U2939 (N_2939,N_876,N_1660);
and U2940 (N_2940,N_1690,N_216);
nand U2941 (N_2941,N_1895,N_1909);
xor U2942 (N_2942,N_374,N_653);
nand U2943 (N_2943,N_1430,N_675);
or U2944 (N_2944,N_1971,N_1340);
xnor U2945 (N_2945,N_1743,N_78);
and U2946 (N_2946,N_728,N_883);
nor U2947 (N_2947,N_862,N_319);
or U2948 (N_2948,N_475,N_1277);
xnor U2949 (N_2949,N_1125,N_367);
nor U2950 (N_2950,N_1595,N_1145);
or U2951 (N_2951,N_1288,N_90);
nor U2952 (N_2952,N_14,N_1007);
nand U2953 (N_2953,N_4,N_905);
or U2954 (N_2954,N_990,N_1545);
nor U2955 (N_2955,N_145,N_1937);
xnor U2956 (N_2956,N_1079,N_1762);
nor U2957 (N_2957,N_1667,N_1414);
nor U2958 (N_2958,N_12,N_1526);
nand U2959 (N_2959,N_710,N_89);
xor U2960 (N_2960,N_526,N_478);
nor U2961 (N_2961,N_1639,N_1456);
or U2962 (N_2962,N_1093,N_638);
and U2963 (N_2963,N_512,N_747);
nand U2964 (N_2964,N_1947,N_823);
and U2965 (N_2965,N_1799,N_85);
nand U2966 (N_2966,N_466,N_616);
nor U2967 (N_2967,N_1748,N_1153);
nor U2968 (N_2968,N_1238,N_154);
xnor U2969 (N_2969,N_386,N_206);
or U2970 (N_2970,N_218,N_311);
nor U2971 (N_2971,N_1112,N_1275);
nor U2972 (N_2972,N_197,N_788);
and U2973 (N_2973,N_351,N_1515);
nor U2974 (N_2974,N_1400,N_469);
nand U2975 (N_2975,N_1491,N_1420);
xor U2976 (N_2976,N_860,N_487);
nand U2977 (N_2977,N_1338,N_1073);
or U2978 (N_2978,N_1473,N_446);
or U2979 (N_2979,N_1253,N_955);
nand U2980 (N_2980,N_1118,N_113);
or U2981 (N_2981,N_893,N_744);
and U2982 (N_2982,N_732,N_663);
and U2983 (N_2983,N_1616,N_121);
nand U2984 (N_2984,N_91,N_1055);
or U2985 (N_2985,N_1865,N_1099);
or U2986 (N_2986,N_129,N_1781);
or U2987 (N_2987,N_169,N_263);
xor U2988 (N_2988,N_210,N_1317);
xnor U2989 (N_2989,N_1226,N_986);
or U2990 (N_2990,N_1876,N_935);
xnor U2991 (N_2991,N_1334,N_753);
nor U2992 (N_2992,N_1878,N_1467);
and U2993 (N_2993,N_542,N_1323);
nand U2994 (N_2994,N_135,N_1915);
nand U2995 (N_2995,N_461,N_1970);
and U2996 (N_2996,N_71,N_1707);
nand U2997 (N_2997,N_74,N_994);
and U2998 (N_2998,N_193,N_688);
or U2999 (N_2999,N_1281,N_491);
and U3000 (N_3000,N_1731,N_683);
and U3001 (N_3001,N_867,N_699);
nor U3002 (N_3002,N_1159,N_1401);
xor U3003 (N_3003,N_1031,N_383);
xor U3004 (N_3004,N_378,N_848);
or U3005 (N_3005,N_287,N_914);
and U3006 (N_3006,N_1164,N_1487);
nor U3007 (N_3007,N_614,N_95);
nand U3008 (N_3008,N_60,N_1177);
nand U3009 (N_3009,N_118,N_1298);
nor U3010 (N_3010,N_728,N_1423);
nor U3011 (N_3011,N_887,N_830);
nor U3012 (N_3012,N_992,N_1903);
xnor U3013 (N_3013,N_1919,N_1145);
or U3014 (N_3014,N_1408,N_1704);
or U3015 (N_3015,N_450,N_986);
nand U3016 (N_3016,N_1863,N_702);
or U3017 (N_3017,N_1075,N_387);
nand U3018 (N_3018,N_927,N_1769);
nand U3019 (N_3019,N_1475,N_7);
nand U3020 (N_3020,N_1903,N_422);
nand U3021 (N_3021,N_394,N_56);
or U3022 (N_3022,N_1755,N_1820);
or U3023 (N_3023,N_1588,N_495);
nor U3024 (N_3024,N_348,N_124);
or U3025 (N_3025,N_1438,N_1674);
nor U3026 (N_3026,N_1692,N_236);
or U3027 (N_3027,N_1911,N_597);
nand U3028 (N_3028,N_654,N_1285);
or U3029 (N_3029,N_1775,N_95);
nand U3030 (N_3030,N_312,N_911);
and U3031 (N_3031,N_381,N_505);
and U3032 (N_3032,N_662,N_744);
or U3033 (N_3033,N_1555,N_390);
nor U3034 (N_3034,N_1305,N_1353);
nor U3035 (N_3035,N_172,N_1096);
xor U3036 (N_3036,N_189,N_382);
and U3037 (N_3037,N_715,N_318);
nand U3038 (N_3038,N_988,N_1103);
or U3039 (N_3039,N_609,N_694);
and U3040 (N_3040,N_708,N_427);
and U3041 (N_3041,N_1654,N_1947);
and U3042 (N_3042,N_1857,N_461);
nand U3043 (N_3043,N_1767,N_1634);
nand U3044 (N_3044,N_1042,N_1144);
nand U3045 (N_3045,N_362,N_601);
and U3046 (N_3046,N_955,N_206);
and U3047 (N_3047,N_958,N_245);
and U3048 (N_3048,N_1805,N_972);
or U3049 (N_3049,N_1677,N_410);
nor U3050 (N_3050,N_1911,N_650);
nand U3051 (N_3051,N_1219,N_1810);
and U3052 (N_3052,N_910,N_905);
and U3053 (N_3053,N_158,N_1819);
nand U3054 (N_3054,N_1238,N_1952);
nand U3055 (N_3055,N_476,N_1677);
and U3056 (N_3056,N_1703,N_122);
nand U3057 (N_3057,N_1032,N_1113);
nor U3058 (N_3058,N_755,N_1488);
nand U3059 (N_3059,N_189,N_861);
or U3060 (N_3060,N_463,N_1164);
nor U3061 (N_3061,N_1246,N_408);
nand U3062 (N_3062,N_789,N_755);
nand U3063 (N_3063,N_686,N_1564);
nor U3064 (N_3064,N_1809,N_1333);
nor U3065 (N_3065,N_1027,N_365);
nor U3066 (N_3066,N_195,N_725);
nand U3067 (N_3067,N_573,N_1706);
and U3068 (N_3068,N_914,N_828);
or U3069 (N_3069,N_372,N_703);
nor U3070 (N_3070,N_1278,N_1189);
and U3071 (N_3071,N_934,N_194);
nand U3072 (N_3072,N_437,N_146);
nor U3073 (N_3073,N_826,N_1648);
xor U3074 (N_3074,N_1485,N_851);
or U3075 (N_3075,N_1945,N_1719);
and U3076 (N_3076,N_540,N_221);
nor U3077 (N_3077,N_729,N_841);
and U3078 (N_3078,N_726,N_1382);
nand U3079 (N_3079,N_1845,N_233);
nor U3080 (N_3080,N_1044,N_252);
and U3081 (N_3081,N_1404,N_25);
nor U3082 (N_3082,N_1173,N_1082);
nor U3083 (N_3083,N_1235,N_427);
and U3084 (N_3084,N_772,N_517);
or U3085 (N_3085,N_24,N_865);
nor U3086 (N_3086,N_1084,N_631);
nor U3087 (N_3087,N_1258,N_667);
nand U3088 (N_3088,N_1862,N_254);
and U3089 (N_3089,N_1933,N_347);
and U3090 (N_3090,N_762,N_28);
nand U3091 (N_3091,N_751,N_1418);
nand U3092 (N_3092,N_1498,N_1423);
or U3093 (N_3093,N_1655,N_452);
nor U3094 (N_3094,N_1705,N_365);
and U3095 (N_3095,N_1981,N_1197);
nand U3096 (N_3096,N_547,N_338);
nand U3097 (N_3097,N_1624,N_1879);
nand U3098 (N_3098,N_869,N_1297);
or U3099 (N_3099,N_1653,N_1603);
nand U3100 (N_3100,N_908,N_1951);
or U3101 (N_3101,N_652,N_1099);
nand U3102 (N_3102,N_1004,N_1645);
xor U3103 (N_3103,N_810,N_520);
or U3104 (N_3104,N_1668,N_345);
nand U3105 (N_3105,N_935,N_1294);
or U3106 (N_3106,N_1912,N_1691);
nor U3107 (N_3107,N_449,N_1387);
xnor U3108 (N_3108,N_1399,N_1673);
and U3109 (N_3109,N_186,N_502);
nand U3110 (N_3110,N_846,N_1828);
nor U3111 (N_3111,N_1820,N_910);
nor U3112 (N_3112,N_2,N_1745);
or U3113 (N_3113,N_1745,N_717);
xnor U3114 (N_3114,N_1170,N_428);
nand U3115 (N_3115,N_1623,N_1353);
nand U3116 (N_3116,N_1399,N_141);
or U3117 (N_3117,N_10,N_1292);
and U3118 (N_3118,N_267,N_1418);
and U3119 (N_3119,N_960,N_1700);
nand U3120 (N_3120,N_760,N_1584);
nor U3121 (N_3121,N_574,N_403);
and U3122 (N_3122,N_727,N_1495);
xnor U3123 (N_3123,N_716,N_731);
and U3124 (N_3124,N_1389,N_413);
and U3125 (N_3125,N_834,N_1984);
nor U3126 (N_3126,N_103,N_515);
nor U3127 (N_3127,N_1002,N_1293);
or U3128 (N_3128,N_1513,N_962);
and U3129 (N_3129,N_1400,N_628);
or U3130 (N_3130,N_1118,N_1143);
nor U3131 (N_3131,N_1315,N_293);
and U3132 (N_3132,N_1409,N_545);
and U3133 (N_3133,N_495,N_851);
or U3134 (N_3134,N_1255,N_1022);
nor U3135 (N_3135,N_1465,N_1870);
and U3136 (N_3136,N_1016,N_608);
xor U3137 (N_3137,N_104,N_514);
and U3138 (N_3138,N_763,N_1074);
nor U3139 (N_3139,N_1024,N_683);
nor U3140 (N_3140,N_1866,N_312);
and U3141 (N_3141,N_1202,N_1786);
and U3142 (N_3142,N_1361,N_261);
nand U3143 (N_3143,N_1237,N_364);
nand U3144 (N_3144,N_1026,N_350);
xor U3145 (N_3145,N_1349,N_680);
or U3146 (N_3146,N_511,N_1125);
or U3147 (N_3147,N_135,N_264);
nor U3148 (N_3148,N_1402,N_730);
nor U3149 (N_3149,N_1425,N_861);
nand U3150 (N_3150,N_1289,N_1395);
or U3151 (N_3151,N_1087,N_1611);
or U3152 (N_3152,N_1766,N_1588);
nor U3153 (N_3153,N_176,N_1697);
nor U3154 (N_3154,N_1753,N_814);
nor U3155 (N_3155,N_1437,N_1933);
nor U3156 (N_3156,N_1151,N_1825);
nand U3157 (N_3157,N_775,N_1667);
nor U3158 (N_3158,N_597,N_1736);
nor U3159 (N_3159,N_1645,N_1846);
or U3160 (N_3160,N_896,N_218);
nand U3161 (N_3161,N_714,N_1058);
nor U3162 (N_3162,N_443,N_936);
or U3163 (N_3163,N_716,N_1967);
and U3164 (N_3164,N_1510,N_992);
nor U3165 (N_3165,N_1491,N_1776);
or U3166 (N_3166,N_310,N_1053);
nand U3167 (N_3167,N_1339,N_1542);
nor U3168 (N_3168,N_1780,N_1295);
or U3169 (N_3169,N_1337,N_405);
or U3170 (N_3170,N_146,N_269);
and U3171 (N_3171,N_1441,N_567);
xor U3172 (N_3172,N_986,N_843);
nor U3173 (N_3173,N_983,N_1177);
and U3174 (N_3174,N_1727,N_287);
and U3175 (N_3175,N_634,N_576);
nand U3176 (N_3176,N_1650,N_859);
nor U3177 (N_3177,N_793,N_1408);
or U3178 (N_3178,N_1670,N_125);
and U3179 (N_3179,N_1300,N_1030);
nor U3180 (N_3180,N_824,N_256);
xnor U3181 (N_3181,N_228,N_1390);
or U3182 (N_3182,N_1209,N_1399);
or U3183 (N_3183,N_905,N_161);
nand U3184 (N_3184,N_592,N_1602);
or U3185 (N_3185,N_1982,N_1572);
nand U3186 (N_3186,N_1555,N_1801);
and U3187 (N_3187,N_286,N_1571);
nand U3188 (N_3188,N_406,N_1286);
nand U3189 (N_3189,N_64,N_1768);
nand U3190 (N_3190,N_755,N_117);
nand U3191 (N_3191,N_755,N_1076);
and U3192 (N_3192,N_1686,N_15);
nor U3193 (N_3193,N_844,N_478);
xnor U3194 (N_3194,N_1706,N_1965);
nand U3195 (N_3195,N_373,N_477);
and U3196 (N_3196,N_764,N_1533);
or U3197 (N_3197,N_717,N_1866);
and U3198 (N_3198,N_418,N_1307);
or U3199 (N_3199,N_1112,N_1764);
or U3200 (N_3200,N_1873,N_1764);
nor U3201 (N_3201,N_1771,N_627);
nor U3202 (N_3202,N_78,N_1679);
nand U3203 (N_3203,N_1746,N_161);
nor U3204 (N_3204,N_522,N_413);
and U3205 (N_3205,N_187,N_1558);
nor U3206 (N_3206,N_615,N_668);
or U3207 (N_3207,N_159,N_636);
or U3208 (N_3208,N_925,N_1762);
nor U3209 (N_3209,N_1027,N_1266);
and U3210 (N_3210,N_712,N_893);
nand U3211 (N_3211,N_384,N_420);
or U3212 (N_3212,N_452,N_1186);
or U3213 (N_3213,N_1226,N_1470);
nor U3214 (N_3214,N_1063,N_821);
and U3215 (N_3215,N_1714,N_403);
or U3216 (N_3216,N_529,N_702);
nor U3217 (N_3217,N_693,N_80);
xnor U3218 (N_3218,N_319,N_1446);
nand U3219 (N_3219,N_592,N_630);
and U3220 (N_3220,N_374,N_1944);
and U3221 (N_3221,N_625,N_26);
and U3222 (N_3222,N_195,N_497);
and U3223 (N_3223,N_495,N_905);
and U3224 (N_3224,N_1091,N_1218);
nor U3225 (N_3225,N_815,N_1149);
xor U3226 (N_3226,N_1965,N_1094);
nand U3227 (N_3227,N_1908,N_1132);
or U3228 (N_3228,N_460,N_1808);
and U3229 (N_3229,N_1806,N_1329);
nand U3230 (N_3230,N_1603,N_1504);
xor U3231 (N_3231,N_1107,N_556);
or U3232 (N_3232,N_65,N_1643);
nor U3233 (N_3233,N_1837,N_133);
nor U3234 (N_3234,N_26,N_815);
and U3235 (N_3235,N_1080,N_434);
nor U3236 (N_3236,N_40,N_1451);
nor U3237 (N_3237,N_1299,N_484);
and U3238 (N_3238,N_428,N_1693);
or U3239 (N_3239,N_804,N_1618);
nand U3240 (N_3240,N_289,N_922);
nand U3241 (N_3241,N_915,N_605);
nand U3242 (N_3242,N_594,N_1916);
nor U3243 (N_3243,N_101,N_1049);
nand U3244 (N_3244,N_731,N_1202);
and U3245 (N_3245,N_1879,N_23);
nor U3246 (N_3246,N_1413,N_132);
nor U3247 (N_3247,N_1306,N_53);
nor U3248 (N_3248,N_1275,N_1668);
nor U3249 (N_3249,N_1569,N_487);
and U3250 (N_3250,N_1658,N_223);
or U3251 (N_3251,N_259,N_1396);
nor U3252 (N_3252,N_474,N_561);
nor U3253 (N_3253,N_715,N_1135);
nor U3254 (N_3254,N_606,N_114);
nor U3255 (N_3255,N_891,N_769);
or U3256 (N_3256,N_1935,N_1371);
xnor U3257 (N_3257,N_120,N_1244);
xor U3258 (N_3258,N_906,N_130);
or U3259 (N_3259,N_226,N_1503);
nand U3260 (N_3260,N_1071,N_256);
nand U3261 (N_3261,N_767,N_726);
nand U3262 (N_3262,N_1889,N_414);
and U3263 (N_3263,N_1403,N_1752);
nor U3264 (N_3264,N_1792,N_1351);
nand U3265 (N_3265,N_819,N_1220);
or U3266 (N_3266,N_896,N_1048);
nand U3267 (N_3267,N_1446,N_963);
and U3268 (N_3268,N_907,N_450);
xor U3269 (N_3269,N_1144,N_1071);
nand U3270 (N_3270,N_1445,N_1538);
nor U3271 (N_3271,N_348,N_1004);
nor U3272 (N_3272,N_487,N_852);
nand U3273 (N_3273,N_847,N_1780);
or U3274 (N_3274,N_787,N_645);
and U3275 (N_3275,N_1003,N_1751);
nand U3276 (N_3276,N_808,N_1292);
or U3277 (N_3277,N_1942,N_1978);
or U3278 (N_3278,N_485,N_859);
nor U3279 (N_3279,N_863,N_1042);
xnor U3280 (N_3280,N_1526,N_1611);
or U3281 (N_3281,N_684,N_1491);
or U3282 (N_3282,N_1329,N_1701);
nand U3283 (N_3283,N_1731,N_1548);
or U3284 (N_3284,N_1151,N_350);
nor U3285 (N_3285,N_710,N_312);
nand U3286 (N_3286,N_1143,N_375);
or U3287 (N_3287,N_1162,N_1405);
or U3288 (N_3288,N_675,N_165);
nand U3289 (N_3289,N_481,N_7);
nor U3290 (N_3290,N_1709,N_1984);
and U3291 (N_3291,N_1031,N_764);
and U3292 (N_3292,N_1379,N_1394);
xor U3293 (N_3293,N_1833,N_442);
and U3294 (N_3294,N_1403,N_1669);
nor U3295 (N_3295,N_1252,N_225);
and U3296 (N_3296,N_30,N_1840);
or U3297 (N_3297,N_1914,N_564);
nand U3298 (N_3298,N_366,N_318);
xor U3299 (N_3299,N_1364,N_1475);
or U3300 (N_3300,N_1120,N_1177);
or U3301 (N_3301,N_1840,N_1173);
nor U3302 (N_3302,N_1440,N_1223);
nand U3303 (N_3303,N_1268,N_2);
nand U3304 (N_3304,N_1560,N_1261);
and U3305 (N_3305,N_1052,N_78);
nor U3306 (N_3306,N_1043,N_1222);
and U3307 (N_3307,N_973,N_1396);
nand U3308 (N_3308,N_1077,N_1470);
nand U3309 (N_3309,N_1045,N_1831);
or U3310 (N_3310,N_1639,N_1437);
nand U3311 (N_3311,N_1852,N_1926);
nor U3312 (N_3312,N_143,N_1401);
and U3313 (N_3313,N_286,N_681);
and U3314 (N_3314,N_1637,N_603);
nand U3315 (N_3315,N_1857,N_1373);
and U3316 (N_3316,N_1056,N_1565);
nand U3317 (N_3317,N_1251,N_175);
and U3318 (N_3318,N_1848,N_981);
and U3319 (N_3319,N_784,N_394);
or U3320 (N_3320,N_544,N_750);
nor U3321 (N_3321,N_698,N_8);
and U3322 (N_3322,N_554,N_1301);
nand U3323 (N_3323,N_982,N_336);
xnor U3324 (N_3324,N_1129,N_604);
xor U3325 (N_3325,N_1814,N_1955);
nand U3326 (N_3326,N_846,N_235);
or U3327 (N_3327,N_355,N_1816);
nor U3328 (N_3328,N_514,N_1514);
xor U3329 (N_3329,N_223,N_452);
xor U3330 (N_3330,N_1981,N_952);
nor U3331 (N_3331,N_1168,N_844);
and U3332 (N_3332,N_1241,N_645);
nand U3333 (N_3333,N_1354,N_250);
or U3334 (N_3334,N_302,N_1925);
xor U3335 (N_3335,N_1833,N_272);
nor U3336 (N_3336,N_1268,N_1370);
and U3337 (N_3337,N_1210,N_889);
nor U3338 (N_3338,N_1281,N_115);
xor U3339 (N_3339,N_1395,N_30);
and U3340 (N_3340,N_265,N_879);
xnor U3341 (N_3341,N_44,N_1406);
nor U3342 (N_3342,N_1130,N_502);
nand U3343 (N_3343,N_46,N_791);
and U3344 (N_3344,N_398,N_1825);
nor U3345 (N_3345,N_1620,N_1968);
nor U3346 (N_3346,N_1242,N_1719);
and U3347 (N_3347,N_821,N_1319);
nor U3348 (N_3348,N_1102,N_1014);
and U3349 (N_3349,N_817,N_408);
nor U3350 (N_3350,N_1512,N_706);
nor U3351 (N_3351,N_844,N_847);
nor U3352 (N_3352,N_1262,N_674);
and U3353 (N_3353,N_753,N_879);
nor U3354 (N_3354,N_1797,N_1412);
nor U3355 (N_3355,N_1841,N_1427);
nor U3356 (N_3356,N_1789,N_1366);
and U3357 (N_3357,N_184,N_1484);
nand U3358 (N_3358,N_1018,N_1378);
nand U3359 (N_3359,N_1065,N_1423);
nand U3360 (N_3360,N_950,N_1448);
nand U3361 (N_3361,N_1570,N_644);
or U3362 (N_3362,N_1864,N_1247);
nor U3363 (N_3363,N_36,N_1495);
nand U3364 (N_3364,N_1756,N_891);
nor U3365 (N_3365,N_1230,N_71);
or U3366 (N_3366,N_1362,N_1534);
and U3367 (N_3367,N_1717,N_696);
and U3368 (N_3368,N_457,N_1422);
nand U3369 (N_3369,N_1127,N_216);
or U3370 (N_3370,N_362,N_1037);
nand U3371 (N_3371,N_424,N_701);
xnor U3372 (N_3372,N_1103,N_172);
nand U3373 (N_3373,N_895,N_551);
or U3374 (N_3374,N_49,N_592);
or U3375 (N_3375,N_535,N_68);
nor U3376 (N_3376,N_1969,N_484);
nand U3377 (N_3377,N_1465,N_1280);
nand U3378 (N_3378,N_716,N_1184);
nor U3379 (N_3379,N_1199,N_1352);
and U3380 (N_3380,N_1941,N_1845);
nand U3381 (N_3381,N_1189,N_1175);
and U3382 (N_3382,N_1780,N_1592);
nor U3383 (N_3383,N_1310,N_1483);
or U3384 (N_3384,N_89,N_167);
or U3385 (N_3385,N_51,N_1748);
and U3386 (N_3386,N_1118,N_1523);
nand U3387 (N_3387,N_1822,N_629);
nand U3388 (N_3388,N_608,N_323);
nor U3389 (N_3389,N_730,N_539);
nand U3390 (N_3390,N_698,N_247);
nor U3391 (N_3391,N_1081,N_1009);
or U3392 (N_3392,N_1951,N_1449);
and U3393 (N_3393,N_11,N_1344);
nor U3394 (N_3394,N_122,N_1109);
xnor U3395 (N_3395,N_1160,N_1604);
and U3396 (N_3396,N_1955,N_891);
xor U3397 (N_3397,N_887,N_874);
and U3398 (N_3398,N_1524,N_855);
xnor U3399 (N_3399,N_492,N_6);
and U3400 (N_3400,N_266,N_383);
and U3401 (N_3401,N_1628,N_207);
nor U3402 (N_3402,N_1085,N_1938);
and U3403 (N_3403,N_944,N_386);
and U3404 (N_3404,N_393,N_135);
or U3405 (N_3405,N_431,N_1086);
and U3406 (N_3406,N_1463,N_666);
nor U3407 (N_3407,N_79,N_1923);
nand U3408 (N_3408,N_67,N_444);
nor U3409 (N_3409,N_1994,N_372);
nor U3410 (N_3410,N_1686,N_365);
nand U3411 (N_3411,N_841,N_884);
nand U3412 (N_3412,N_369,N_1875);
nand U3413 (N_3413,N_1597,N_327);
or U3414 (N_3414,N_1914,N_1254);
nand U3415 (N_3415,N_1601,N_523);
and U3416 (N_3416,N_1309,N_625);
xor U3417 (N_3417,N_460,N_499);
xor U3418 (N_3418,N_459,N_1652);
or U3419 (N_3419,N_1238,N_1310);
or U3420 (N_3420,N_1505,N_939);
and U3421 (N_3421,N_1348,N_1332);
nor U3422 (N_3422,N_37,N_193);
nor U3423 (N_3423,N_1444,N_952);
xnor U3424 (N_3424,N_484,N_1291);
nor U3425 (N_3425,N_51,N_689);
nor U3426 (N_3426,N_944,N_222);
xnor U3427 (N_3427,N_1263,N_168);
and U3428 (N_3428,N_182,N_678);
nor U3429 (N_3429,N_965,N_245);
or U3430 (N_3430,N_1507,N_1837);
nor U3431 (N_3431,N_616,N_416);
xor U3432 (N_3432,N_1258,N_1806);
or U3433 (N_3433,N_1358,N_1734);
nand U3434 (N_3434,N_1118,N_1622);
nor U3435 (N_3435,N_1805,N_1928);
or U3436 (N_3436,N_1342,N_1977);
and U3437 (N_3437,N_163,N_1375);
and U3438 (N_3438,N_441,N_1744);
and U3439 (N_3439,N_1215,N_707);
and U3440 (N_3440,N_108,N_1029);
nor U3441 (N_3441,N_31,N_299);
or U3442 (N_3442,N_1455,N_74);
or U3443 (N_3443,N_1770,N_1225);
xnor U3444 (N_3444,N_1341,N_1800);
and U3445 (N_3445,N_1163,N_1402);
xor U3446 (N_3446,N_1512,N_473);
nor U3447 (N_3447,N_463,N_1942);
nor U3448 (N_3448,N_86,N_797);
nand U3449 (N_3449,N_1151,N_471);
nor U3450 (N_3450,N_339,N_1410);
or U3451 (N_3451,N_409,N_713);
xnor U3452 (N_3452,N_1976,N_1795);
xor U3453 (N_3453,N_1733,N_902);
xor U3454 (N_3454,N_1128,N_772);
nor U3455 (N_3455,N_1890,N_1035);
nor U3456 (N_3456,N_343,N_118);
xor U3457 (N_3457,N_827,N_39);
nand U3458 (N_3458,N_1748,N_1198);
nor U3459 (N_3459,N_156,N_531);
or U3460 (N_3460,N_159,N_582);
nand U3461 (N_3461,N_409,N_1222);
nand U3462 (N_3462,N_16,N_1870);
nor U3463 (N_3463,N_1634,N_254);
nand U3464 (N_3464,N_1916,N_299);
or U3465 (N_3465,N_1966,N_1055);
and U3466 (N_3466,N_396,N_804);
nand U3467 (N_3467,N_312,N_893);
or U3468 (N_3468,N_476,N_1052);
nand U3469 (N_3469,N_1830,N_127);
nor U3470 (N_3470,N_1398,N_733);
nor U3471 (N_3471,N_1850,N_1827);
or U3472 (N_3472,N_132,N_1282);
and U3473 (N_3473,N_1937,N_301);
nand U3474 (N_3474,N_391,N_810);
nor U3475 (N_3475,N_162,N_803);
nand U3476 (N_3476,N_1945,N_1735);
xor U3477 (N_3477,N_757,N_652);
and U3478 (N_3478,N_1118,N_439);
or U3479 (N_3479,N_1209,N_1959);
and U3480 (N_3480,N_157,N_566);
nand U3481 (N_3481,N_101,N_1759);
nand U3482 (N_3482,N_247,N_171);
nor U3483 (N_3483,N_696,N_1558);
nor U3484 (N_3484,N_1051,N_1285);
nand U3485 (N_3485,N_316,N_19);
or U3486 (N_3486,N_1724,N_1074);
xor U3487 (N_3487,N_865,N_823);
nand U3488 (N_3488,N_230,N_1742);
nor U3489 (N_3489,N_1018,N_1885);
nand U3490 (N_3490,N_1418,N_12);
and U3491 (N_3491,N_20,N_1319);
nand U3492 (N_3492,N_1927,N_1226);
or U3493 (N_3493,N_611,N_857);
and U3494 (N_3494,N_1017,N_101);
or U3495 (N_3495,N_1888,N_1245);
nand U3496 (N_3496,N_1858,N_384);
or U3497 (N_3497,N_824,N_1115);
nand U3498 (N_3498,N_884,N_663);
nor U3499 (N_3499,N_731,N_1022);
nand U3500 (N_3500,N_769,N_477);
and U3501 (N_3501,N_1282,N_1392);
nor U3502 (N_3502,N_1888,N_1039);
and U3503 (N_3503,N_545,N_1816);
nor U3504 (N_3504,N_1642,N_797);
and U3505 (N_3505,N_1436,N_394);
xnor U3506 (N_3506,N_345,N_452);
or U3507 (N_3507,N_240,N_121);
nand U3508 (N_3508,N_297,N_676);
and U3509 (N_3509,N_1649,N_1378);
xor U3510 (N_3510,N_1071,N_1999);
nand U3511 (N_3511,N_1217,N_1957);
and U3512 (N_3512,N_362,N_293);
nor U3513 (N_3513,N_1527,N_1867);
or U3514 (N_3514,N_422,N_1541);
nand U3515 (N_3515,N_942,N_1122);
nor U3516 (N_3516,N_1261,N_432);
and U3517 (N_3517,N_916,N_1042);
or U3518 (N_3518,N_510,N_1876);
and U3519 (N_3519,N_1369,N_1823);
and U3520 (N_3520,N_1304,N_378);
nand U3521 (N_3521,N_683,N_1905);
and U3522 (N_3522,N_1387,N_1614);
xnor U3523 (N_3523,N_1040,N_1456);
nor U3524 (N_3524,N_74,N_1534);
xnor U3525 (N_3525,N_1877,N_1049);
nand U3526 (N_3526,N_471,N_924);
nor U3527 (N_3527,N_773,N_1809);
nand U3528 (N_3528,N_149,N_742);
nor U3529 (N_3529,N_992,N_289);
nand U3530 (N_3530,N_1068,N_802);
and U3531 (N_3531,N_1464,N_856);
nor U3532 (N_3532,N_130,N_1131);
nand U3533 (N_3533,N_717,N_54);
xor U3534 (N_3534,N_1205,N_1508);
and U3535 (N_3535,N_98,N_263);
xor U3536 (N_3536,N_1703,N_1814);
nand U3537 (N_3537,N_982,N_1112);
nand U3538 (N_3538,N_973,N_415);
nand U3539 (N_3539,N_1535,N_313);
and U3540 (N_3540,N_546,N_193);
nor U3541 (N_3541,N_1698,N_462);
nand U3542 (N_3542,N_705,N_873);
and U3543 (N_3543,N_968,N_502);
or U3544 (N_3544,N_77,N_972);
or U3545 (N_3545,N_125,N_506);
nor U3546 (N_3546,N_881,N_21);
xnor U3547 (N_3547,N_1355,N_1164);
and U3548 (N_3548,N_1018,N_623);
nor U3549 (N_3549,N_809,N_288);
and U3550 (N_3550,N_1602,N_211);
and U3551 (N_3551,N_619,N_31);
nor U3552 (N_3552,N_848,N_1604);
nand U3553 (N_3553,N_1563,N_1521);
nand U3554 (N_3554,N_1291,N_556);
and U3555 (N_3555,N_104,N_1338);
nand U3556 (N_3556,N_1920,N_1745);
nand U3557 (N_3557,N_1389,N_638);
nand U3558 (N_3558,N_1674,N_812);
nor U3559 (N_3559,N_1888,N_1798);
nand U3560 (N_3560,N_1819,N_1978);
nand U3561 (N_3561,N_414,N_789);
or U3562 (N_3562,N_808,N_742);
or U3563 (N_3563,N_1366,N_1977);
nand U3564 (N_3564,N_887,N_1043);
xor U3565 (N_3565,N_1446,N_1665);
xor U3566 (N_3566,N_609,N_1482);
and U3567 (N_3567,N_76,N_1665);
and U3568 (N_3568,N_626,N_128);
nand U3569 (N_3569,N_1430,N_314);
and U3570 (N_3570,N_1747,N_348);
or U3571 (N_3571,N_983,N_699);
nor U3572 (N_3572,N_987,N_1124);
nand U3573 (N_3573,N_1562,N_544);
nand U3574 (N_3574,N_1115,N_1722);
xnor U3575 (N_3575,N_752,N_1436);
nor U3576 (N_3576,N_1846,N_1683);
or U3577 (N_3577,N_52,N_1663);
and U3578 (N_3578,N_1305,N_1860);
nand U3579 (N_3579,N_442,N_998);
and U3580 (N_3580,N_1697,N_1187);
nand U3581 (N_3581,N_745,N_874);
nor U3582 (N_3582,N_1279,N_305);
nor U3583 (N_3583,N_1399,N_998);
or U3584 (N_3584,N_1676,N_1235);
or U3585 (N_3585,N_424,N_1334);
nor U3586 (N_3586,N_1769,N_1586);
nand U3587 (N_3587,N_364,N_1422);
xnor U3588 (N_3588,N_102,N_841);
and U3589 (N_3589,N_1103,N_1187);
nor U3590 (N_3590,N_1013,N_458);
or U3591 (N_3591,N_1554,N_448);
and U3592 (N_3592,N_872,N_1524);
or U3593 (N_3593,N_1011,N_1057);
xnor U3594 (N_3594,N_333,N_57);
and U3595 (N_3595,N_340,N_18);
nor U3596 (N_3596,N_676,N_307);
nand U3597 (N_3597,N_1719,N_1499);
nor U3598 (N_3598,N_1036,N_1336);
nand U3599 (N_3599,N_1,N_1542);
nor U3600 (N_3600,N_334,N_747);
nand U3601 (N_3601,N_1631,N_1199);
nand U3602 (N_3602,N_923,N_1825);
nand U3603 (N_3603,N_102,N_1980);
or U3604 (N_3604,N_1017,N_1038);
or U3605 (N_3605,N_0,N_609);
or U3606 (N_3606,N_68,N_1180);
xnor U3607 (N_3607,N_498,N_839);
xor U3608 (N_3608,N_801,N_1748);
or U3609 (N_3609,N_39,N_1075);
and U3610 (N_3610,N_488,N_180);
nand U3611 (N_3611,N_263,N_165);
nand U3612 (N_3612,N_838,N_172);
nor U3613 (N_3613,N_791,N_1867);
nor U3614 (N_3614,N_1265,N_315);
and U3615 (N_3615,N_301,N_111);
and U3616 (N_3616,N_965,N_1760);
nand U3617 (N_3617,N_711,N_474);
nand U3618 (N_3618,N_635,N_1193);
nor U3619 (N_3619,N_674,N_400);
or U3620 (N_3620,N_157,N_461);
and U3621 (N_3621,N_272,N_1432);
xor U3622 (N_3622,N_427,N_1432);
nor U3623 (N_3623,N_1615,N_936);
nand U3624 (N_3624,N_244,N_305);
and U3625 (N_3625,N_749,N_82);
nand U3626 (N_3626,N_734,N_835);
nand U3627 (N_3627,N_1702,N_1834);
or U3628 (N_3628,N_1044,N_288);
nor U3629 (N_3629,N_1179,N_1715);
and U3630 (N_3630,N_1009,N_1369);
xor U3631 (N_3631,N_1995,N_1080);
nor U3632 (N_3632,N_1610,N_1365);
and U3633 (N_3633,N_1808,N_1183);
nand U3634 (N_3634,N_1931,N_1267);
and U3635 (N_3635,N_964,N_128);
nor U3636 (N_3636,N_846,N_943);
nand U3637 (N_3637,N_112,N_1327);
nand U3638 (N_3638,N_756,N_850);
xnor U3639 (N_3639,N_1773,N_327);
or U3640 (N_3640,N_637,N_845);
and U3641 (N_3641,N_1839,N_118);
nand U3642 (N_3642,N_1067,N_161);
or U3643 (N_3643,N_1392,N_1947);
nand U3644 (N_3644,N_895,N_1602);
xor U3645 (N_3645,N_1491,N_996);
nor U3646 (N_3646,N_666,N_950);
and U3647 (N_3647,N_1155,N_989);
nand U3648 (N_3648,N_280,N_1928);
or U3649 (N_3649,N_607,N_1546);
nor U3650 (N_3650,N_1549,N_1404);
nor U3651 (N_3651,N_912,N_813);
or U3652 (N_3652,N_1884,N_555);
or U3653 (N_3653,N_1135,N_1687);
xnor U3654 (N_3654,N_1837,N_1825);
nor U3655 (N_3655,N_384,N_1423);
nand U3656 (N_3656,N_882,N_845);
xnor U3657 (N_3657,N_312,N_63);
nor U3658 (N_3658,N_254,N_1951);
and U3659 (N_3659,N_1157,N_1362);
nor U3660 (N_3660,N_1137,N_1442);
nand U3661 (N_3661,N_289,N_1153);
and U3662 (N_3662,N_1684,N_601);
and U3663 (N_3663,N_582,N_691);
or U3664 (N_3664,N_1034,N_1828);
nand U3665 (N_3665,N_639,N_526);
or U3666 (N_3666,N_1613,N_1369);
or U3667 (N_3667,N_962,N_311);
or U3668 (N_3668,N_441,N_1431);
and U3669 (N_3669,N_642,N_216);
xnor U3670 (N_3670,N_762,N_380);
xor U3671 (N_3671,N_285,N_538);
xnor U3672 (N_3672,N_1388,N_167);
nor U3673 (N_3673,N_1632,N_943);
nand U3674 (N_3674,N_1640,N_967);
and U3675 (N_3675,N_89,N_553);
and U3676 (N_3676,N_1962,N_1674);
and U3677 (N_3677,N_1825,N_1391);
nand U3678 (N_3678,N_142,N_752);
and U3679 (N_3679,N_1310,N_77);
or U3680 (N_3680,N_104,N_1938);
or U3681 (N_3681,N_1839,N_867);
nand U3682 (N_3682,N_1458,N_1522);
nor U3683 (N_3683,N_437,N_518);
nor U3684 (N_3684,N_139,N_1772);
and U3685 (N_3685,N_276,N_1275);
nand U3686 (N_3686,N_1809,N_512);
and U3687 (N_3687,N_27,N_513);
or U3688 (N_3688,N_1067,N_484);
nand U3689 (N_3689,N_1399,N_1462);
nor U3690 (N_3690,N_1978,N_520);
and U3691 (N_3691,N_1604,N_1584);
xnor U3692 (N_3692,N_1821,N_1178);
nor U3693 (N_3693,N_683,N_288);
and U3694 (N_3694,N_1449,N_865);
nand U3695 (N_3695,N_8,N_1899);
nor U3696 (N_3696,N_142,N_1020);
nand U3697 (N_3697,N_91,N_746);
or U3698 (N_3698,N_865,N_818);
and U3699 (N_3699,N_1698,N_1857);
nand U3700 (N_3700,N_180,N_642);
and U3701 (N_3701,N_1388,N_1987);
and U3702 (N_3702,N_497,N_1860);
or U3703 (N_3703,N_508,N_1974);
and U3704 (N_3704,N_71,N_320);
or U3705 (N_3705,N_1945,N_1944);
xnor U3706 (N_3706,N_1851,N_68);
nand U3707 (N_3707,N_1508,N_174);
xor U3708 (N_3708,N_1942,N_428);
xnor U3709 (N_3709,N_1421,N_1393);
and U3710 (N_3710,N_504,N_276);
and U3711 (N_3711,N_1108,N_794);
and U3712 (N_3712,N_1596,N_610);
nor U3713 (N_3713,N_241,N_1954);
or U3714 (N_3714,N_1010,N_710);
nand U3715 (N_3715,N_549,N_646);
or U3716 (N_3716,N_649,N_1593);
nand U3717 (N_3717,N_1736,N_1512);
nand U3718 (N_3718,N_1345,N_196);
and U3719 (N_3719,N_440,N_228);
and U3720 (N_3720,N_1557,N_1087);
or U3721 (N_3721,N_1278,N_1769);
nor U3722 (N_3722,N_913,N_757);
xnor U3723 (N_3723,N_1268,N_214);
xnor U3724 (N_3724,N_1198,N_731);
and U3725 (N_3725,N_1279,N_274);
and U3726 (N_3726,N_240,N_880);
or U3727 (N_3727,N_1369,N_757);
nand U3728 (N_3728,N_520,N_1902);
and U3729 (N_3729,N_1979,N_1951);
or U3730 (N_3730,N_1029,N_1349);
nor U3731 (N_3731,N_821,N_1475);
nand U3732 (N_3732,N_289,N_985);
or U3733 (N_3733,N_1817,N_1723);
xnor U3734 (N_3734,N_1211,N_515);
or U3735 (N_3735,N_1897,N_1552);
nand U3736 (N_3736,N_474,N_1786);
or U3737 (N_3737,N_872,N_1562);
nand U3738 (N_3738,N_512,N_1297);
nand U3739 (N_3739,N_361,N_1518);
and U3740 (N_3740,N_1785,N_925);
xnor U3741 (N_3741,N_474,N_1512);
nor U3742 (N_3742,N_1304,N_1294);
or U3743 (N_3743,N_594,N_660);
and U3744 (N_3744,N_1195,N_1875);
and U3745 (N_3745,N_1811,N_1943);
xor U3746 (N_3746,N_1134,N_842);
and U3747 (N_3747,N_1965,N_620);
and U3748 (N_3748,N_864,N_581);
or U3749 (N_3749,N_630,N_1233);
nor U3750 (N_3750,N_1384,N_1775);
and U3751 (N_3751,N_883,N_520);
or U3752 (N_3752,N_942,N_1037);
and U3753 (N_3753,N_1278,N_244);
or U3754 (N_3754,N_133,N_221);
and U3755 (N_3755,N_443,N_1717);
nor U3756 (N_3756,N_1979,N_1363);
nor U3757 (N_3757,N_1712,N_1733);
and U3758 (N_3758,N_487,N_1299);
nand U3759 (N_3759,N_400,N_1855);
nor U3760 (N_3760,N_1931,N_293);
and U3761 (N_3761,N_787,N_712);
and U3762 (N_3762,N_592,N_1756);
nand U3763 (N_3763,N_1364,N_1984);
or U3764 (N_3764,N_984,N_824);
nor U3765 (N_3765,N_860,N_961);
and U3766 (N_3766,N_100,N_35);
or U3767 (N_3767,N_703,N_1831);
nor U3768 (N_3768,N_1180,N_899);
and U3769 (N_3769,N_167,N_612);
and U3770 (N_3770,N_824,N_298);
nand U3771 (N_3771,N_62,N_1962);
or U3772 (N_3772,N_1758,N_233);
nor U3773 (N_3773,N_52,N_949);
or U3774 (N_3774,N_1693,N_796);
nor U3775 (N_3775,N_319,N_1745);
or U3776 (N_3776,N_1327,N_163);
or U3777 (N_3777,N_703,N_150);
nand U3778 (N_3778,N_12,N_1238);
and U3779 (N_3779,N_1554,N_1185);
nand U3780 (N_3780,N_1302,N_1713);
nand U3781 (N_3781,N_392,N_203);
or U3782 (N_3782,N_1400,N_1146);
nor U3783 (N_3783,N_796,N_768);
and U3784 (N_3784,N_801,N_1905);
nand U3785 (N_3785,N_1917,N_571);
and U3786 (N_3786,N_1361,N_1180);
or U3787 (N_3787,N_1804,N_619);
xor U3788 (N_3788,N_1783,N_568);
and U3789 (N_3789,N_1429,N_52);
or U3790 (N_3790,N_349,N_1521);
nor U3791 (N_3791,N_1767,N_985);
or U3792 (N_3792,N_423,N_359);
nor U3793 (N_3793,N_1188,N_317);
xnor U3794 (N_3794,N_28,N_464);
or U3795 (N_3795,N_1564,N_1667);
nand U3796 (N_3796,N_962,N_1341);
and U3797 (N_3797,N_47,N_1991);
nand U3798 (N_3798,N_1387,N_150);
or U3799 (N_3799,N_799,N_234);
nand U3800 (N_3800,N_726,N_1844);
nand U3801 (N_3801,N_1728,N_1453);
and U3802 (N_3802,N_1210,N_1675);
nand U3803 (N_3803,N_700,N_1770);
or U3804 (N_3804,N_1113,N_1343);
xor U3805 (N_3805,N_408,N_1343);
nor U3806 (N_3806,N_1295,N_441);
nand U3807 (N_3807,N_1351,N_1684);
nor U3808 (N_3808,N_619,N_1832);
nor U3809 (N_3809,N_1893,N_315);
and U3810 (N_3810,N_358,N_178);
xnor U3811 (N_3811,N_1178,N_992);
nor U3812 (N_3812,N_1338,N_1728);
nor U3813 (N_3813,N_581,N_162);
xnor U3814 (N_3814,N_546,N_560);
nor U3815 (N_3815,N_1323,N_1283);
and U3816 (N_3816,N_1801,N_95);
nor U3817 (N_3817,N_1335,N_1100);
nand U3818 (N_3818,N_481,N_1871);
and U3819 (N_3819,N_1502,N_559);
or U3820 (N_3820,N_1975,N_207);
nand U3821 (N_3821,N_1478,N_1620);
or U3822 (N_3822,N_314,N_841);
nand U3823 (N_3823,N_1365,N_244);
and U3824 (N_3824,N_1761,N_391);
nand U3825 (N_3825,N_1613,N_303);
and U3826 (N_3826,N_1437,N_813);
or U3827 (N_3827,N_1461,N_853);
nand U3828 (N_3828,N_322,N_784);
xnor U3829 (N_3829,N_456,N_751);
or U3830 (N_3830,N_5,N_1716);
nand U3831 (N_3831,N_1592,N_1718);
nand U3832 (N_3832,N_569,N_1729);
or U3833 (N_3833,N_1876,N_1819);
or U3834 (N_3834,N_1522,N_1398);
nor U3835 (N_3835,N_1066,N_21);
and U3836 (N_3836,N_1505,N_558);
nand U3837 (N_3837,N_1646,N_584);
nor U3838 (N_3838,N_213,N_729);
nand U3839 (N_3839,N_726,N_1895);
nor U3840 (N_3840,N_897,N_781);
nor U3841 (N_3841,N_174,N_1281);
nand U3842 (N_3842,N_853,N_1782);
and U3843 (N_3843,N_331,N_471);
or U3844 (N_3844,N_1611,N_1439);
and U3845 (N_3845,N_723,N_1504);
nor U3846 (N_3846,N_982,N_609);
and U3847 (N_3847,N_1861,N_985);
nand U3848 (N_3848,N_113,N_1014);
nand U3849 (N_3849,N_1415,N_1609);
or U3850 (N_3850,N_513,N_901);
nor U3851 (N_3851,N_197,N_1369);
xnor U3852 (N_3852,N_832,N_1468);
nor U3853 (N_3853,N_883,N_1703);
nand U3854 (N_3854,N_205,N_475);
or U3855 (N_3855,N_474,N_1806);
xnor U3856 (N_3856,N_1988,N_1715);
and U3857 (N_3857,N_870,N_775);
and U3858 (N_3858,N_1090,N_1554);
nor U3859 (N_3859,N_250,N_1136);
nor U3860 (N_3860,N_1230,N_1917);
nand U3861 (N_3861,N_1354,N_1740);
nand U3862 (N_3862,N_75,N_722);
nand U3863 (N_3863,N_81,N_32);
or U3864 (N_3864,N_201,N_415);
nor U3865 (N_3865,N_1353,N_1859);
and U3866 (N_3866,N_1398,N_763);
nor U3867 (N_3867,N_390,N_724);
and U3868 (N_3868,N_202,N_893);
nor U3869 (N_3869,N_1191,N_959);
and U3870 (N_3870,N_1224,N_1688);
nor U3871 (N_3871,N_322,N_1961);
or U3872 (N_3872,N_689,N_567);
nand U3873 (N_3873,N_979,N_679);
or U3874 (N_3874,N_1035,N_65);
or U3875 (N_3875,N_549,N_466);
xnor U3876 (N_3876,N_1785,N_1509);
nor U3877 (N_3877,N_1821,N_926);
xnor U3878 (N_3878,N_1189,N_313);
nand U3879 (N_3879,N_483,N_2);
or U3880 (N_3880,N_777,N_1238);
nor U3881 (N_3881,N_1637,N_1023);
and U3882 (N_3882,N_1806,N_1058);
nand U3883 (N_3883,N_959,N_427);
or U3884 (N_3884,N_865,N_1834);
or U3885 (N_3885,N_1700,N_343);
and U3886 (N_3886,N_1031,N_926);
and U3887 (N_3887,N_1700,N_688);
or U3888 (N_3888,N_604,N_870);
or U3889 (N_3889,N_14,N_1722);
nand U3890 (N_3890,N_1293,N_1992);
xnor U3891 (N_3891,N_1348,N_1824);
nand U3892 (N_3892,N_1772,N_1751);
and U3893 (N_3893,N_1421,N_1413);
nor U3894 (N_3894,N_550,N_1398);
xnor U3895 (N_3895,N_1781,N_1248);
or U3896 (N_3896,N_1549,N_1044);
and U3897 (N_3897,N_1128,N_1846);
nand U3898 (N_3898,N_1547,N_1043);
nand U3899 (N_3899,N_733,N_125);
or U3900 (N_3900,N_1460,N_54);
or U3901 (N_3901,N_1545,N_1587);
and U3902 (N_3902,N_914,N_249);
nand U3903 (N_3903,N_1576,N_1561);
nand U3904 (N_3904,N_1205,N_1117);
nor U3905 (N_3905,N_137,N_1647);
or U3906 (N_3906,N_1889,N_1825);
or U3907 (N_3907,N_186,N_932);
or U3908 (N_3908,N_806,N_1970);
and U3909 (N_3909,N_1025,N_1879);
nand U3910 (N_3910,N_385,N_1463);
or U3911 (N_3911,N_296,N_247);
and U3912 (N_3912,N_439,N_1792);
nand U3913 (N_3913,N_87,N_1240);
nand U3914 (N_3914,N_819,N_179);
or U3915 (N_3915,N_1096,N_259);
or U3916 (N_3916,N_972,N_186);
xor U3917 (N_3917,N_771,N_1018);
nand U3918 (N_3918,N_1494,N_267);
xnor U3919 (N_3919,N_242,N_1735);
nor U3920 (N_3920,N_1259,N_969);
nor U3921 (N_3921,N_804,N_1217);
and U3922 (N_3922,N_641,N_1956);
and U3923 (N_3923,N_387,N_1936);
or U3924 (N_3924,N_171,N_1224);
nand U3925 (N_3925,N_444,N_1288);
xor U3926 (N_3926,N_799,N_1031);
or U3927 (N_3927,N_1625,N_1768);
nor U3928 (N_3928,N_1159,N_873);
xor U3929 (N_3929,N_1872,N_1126);
and U3930 (N_3930,N_581,N_1205);
and U3931 (N_3931,N_1546,N_1563);
nor U3932 (N_3932,N_1547,N_119);
nor U3933 (N_3933,N_1856,N_1906);
and U3934 (N_3934,N_31,N_385);
nor U3935 (N_3935,N_185,N_237);
nor U3936 (N_3936,N_1375,N_1119);
or U3937 (N_3937,N_1763,N_1585);
nor U3938 (N_3938,N_554,N_291);
or U3939 (N_3939,N_1741,N_1649);
or U3940 (N_3940,N_494,N_1672);
or U3941 (N_3941,N_946,N_101);
and U3942 (N_3942,N_1194,N_1091);
nor U3943 (N_3943,N_1340,N_1273);
nand U3944 (N_3944,N_1681,N_458);
xnor U3945 (N_3945,N_115,N_614);
xor U3946 (N_3946,N_1856,N_784);
and U3947 (N_3947,N_275,N_1910);
and U3948 (N_3948,N_1149,N_209);
nor U3949 (N_3949,N_801,N_1345);
and U3950 (N_3950,N_127,N_190);
or U3951 (N_3951,N_1873,N_365);
xnor U3952 (N_3952,N_1327,N_1067);
and U3953 (N_3953,N_517,N_1851);
or U3954 (N_3954,N_1489,N_1473);
or U3955 (N_3955,N_1027,N_461);
and U3956 (N_3956,N_884,N_1743);
nor U3957 (N_3957,N_754,N_92);
or U3958 (N_3958,N_1716,N_353);
and U3959 (N_3959,N_1635,N_511);
nand U3960 (N_3960,N_593,N_1845);
or U3961 (N_3961,N_1492,N_1914);
nor U3962 (N_3962,N_581,N_318);
or U3963 (N_3963,N_331,N_1251);
or U3964 (N_3964,N_1342,N_1374);
and U3965 (N_3965,N_1271,N_1802);
nand U3966 (N_3966,N_795,N_1168);
or U3967 (N_3967,N_1377,N_526);
or U3968 (N_3968,N_1584,N_1759);
nor U3969 (N_3969,N_84,N_689);
nand U3970 (N_3970,N_633,N_1011);
nand U3971 (N_3971,N_419,N_1733);
and U3972 (N_3972,N_1332,N_29);
nand U3973 (N_3973,N_1678,N_289);
or U3974 (N_3974,N_1729,N_167);
xor U3975 (N_3975,N_370,N_1019);
xnor U3976 (N_3976,N_95,N_1407);
or U3977 (N_3977,N_1165,N_689);
nor U3978 (N_3978,N_815,N_1744);
and U3979 (N_3979,N_918,N_1083);
and U3980 (N_3980,N_1787,N_567);
nor U3981 (N_3981,N_892,N_177);
nor U3982 (N_3982,N_918,N_1085);
or U3983 (N_3983,N_346,N_443);
and U3984 (N_3984,N_524,N_1672);
nor U3985 (N_3985,N_1968,N_1838);
nor U3986 (N_3986,N_1135,N_1636);
nand U3987 (N_3987,N_1028,N_538);
nor U3988 (N_3988,N_775,N_670);
and U3989 (N_3989,N_620,N_1874);
nor U3990 (N_3990,N_581,N_757);
nor U3991 (N_3991,N_1091,N_246);
or U3992 (N_3992,N_1790,N_1352);
nand U3993 (N_3993,N_1306,N_918);
and U3994 (N_3994,N_304,N_1098);
and U3995 (N_3995,N_417,N_1605);
and U3996 (N_3996,N_1087,N_448);
nor U3997 (N_3997,N_1161,N_1112);
or U3998 (N_3998,N_356,N_762);
nor U3999 (N_3999,N_1686,N_1533);
or U4000 (N_4000,N_2680,N_2854);
and U4001 (N_4001,N_2216,N_3919);
nor U4002 (N_4002,N_2954,N_3103);
nand U4003 (N_4003,N_3984,N_2846);
and U4004 (N_4004,N_2898,N_3119);
or U4005 (N_4005,N_3931,N_3894);
xor U4006 (N_4006,N_2416,N_3042);
or U4007 (N_4007,N_2450,N_2805);
nand U4008 (N_4008,N_3829,N_2254);
nand U4009 (N_4009,N_3791,N_3844);
xor U4010 (N_4010,N_2403,N_2966);
or U4011 (N_4011,N_2269,N_2794);
and U4012 (N_4012,N_3780,N_2591);
nor U4013 (N_4013,N_2369,N_2114);
or U4014 (N_4014,N_2701,N_2516);
and U4015 (N_4015,N_2857,N_3084);
nor U4016 (N_4016,N_2359,N_2429);
or U4017 (N_4017,N_3129,N_2070);
nand U4018 (N_4018,N_2776,N_2272);
or U4019 (N_4019,N_3339,N_2512);
or U4020 (N_4020,N_3605,N_2210);
nand U4021 (N_4021,N_2436,N_3724);
nand U4022 (N_4022,N_2159,N_2896);
nor U4023 (N_4023,N_2273,N_2848);
or U4024 (N_4024,N_3632,N_3449);
and U4025 (N_4025,N_2305,N_3257);
nand U4026 (N_4026,N_3874,N_3132);
or U4027 (N_4027,N_3531,N_3029);
nor U4028 (N_4028,N_2021,N_3398);
or U4029 (N_4029,N_3234,N_2354);
nor U4030 (N_4030,N_3429,N_2072);
xnor U4031 (N_4031,N_3364,N_3394);
nand U4032 (N_4032,N_3579,N_3849);
nand U4033 (N_4033,N_2598,N_2692);
and U4034 (N_4034,N_3503,N_3804);
nand U4035 (N_4035,N_3170,N_3157);
nor U4036 (N_4036,N_2376,N_2533);
xnor U4037 (N_4037,N_3896,N_2582);
nor U4038 (N_4038,N_2623,N_3606);
and U4039 (N_4039,N_3920,N_2174);
or U4040 (N_4040,N_3872,N_2517);
xor U4041 (N_4041,N_3341,N_2628);
nor U4042 (N_4042,N_3373,N_3943);
nand U4043 (N_4043,N_3703,N_2382);
xor U4044 (N_4044,N_3087,N_2586);
or U4045 (N_4045,N_3004,N_3773);
and U4046 (N_4046,N_2513,N_2042);
nor U4047 (N_4047,N_2654,N_3682);
and U4048 (N_4048,N_2818,N_2027);
or U4049 (N_4049,N_3971,N_3127);
and U4050 (N_4050,N_2163,N_2478);
xnor U4051 (N_4051,N_2212,N_3291);
xnor U4052 (N_4052,N_3051,N_3768);
or U4053 (N_4053,N_3962,N_2324);
xnor U4054 (N_4054,N_3308,N_3522);
xor U4055 (N_4055,N_2120,N_2464);
nand U4056 (N_4056,N_3450,N_3774);
or U4057 (N_4057,N_2322,N_2064);
and U4058 (N_4058,N_3559,N_3824);
nor U4059 (N_4059,N_3864,N_2521);
nor U4060 (N_4060,N_2566,N_2691);
and U4061 (N_4061,N_2204,N_3360);
nor U4062 (N_4062,N_2226,N_3539);
nand U4063 (N_4063,N_3865,N_3496);
or U4064 (N_4064,N_2507,N_2152);
or U4065 (N_4065,N_3035,N_2677);
nand U4066 (N_4066,N_2798,N_3944);
and U4067 (N_4067,N_2866,N_3616);
and U4068 (N_4068,N_3468,N_3899);
nor U4069 (N_4069,N_3965,N_3996);
nor U4070 (N_4070,N_2388,N_2375);
nor U4071 (N_4071,N_3722,N_3909);
and U4072 (N_4072,N_3715,N_2637);
nand U4073 (N_4073,N_3334,N_2187);
nand U4074 (N_4074,N_3779,N_3858);
nand U4075 (N_4075,N_2585,N_2130);
or U4076 (N_4076,N_3556,N_2283);
nand U4077 (N_4077,N_2752,N_2535);
and U4078 (N_4078,N_3846,N_2518);
nand U4079 (N_4079,N_2017,N_2143);
and U4080 (N_4080,N_3913,N_3174);
nor U4081 (N_4081,N_2786,N_3669);
nand U4082 (N_4082,N_2942,N_3597);
nor U4083 (N_4083,N_2800,N_3305);
or U4084 (N_4084,N_3204,N_2165);
and U4085 (N_4085,N_3240,N_2061);
or U4086 (N_4086,N_3277,N_3440);
nor U4087 (N_4087,N_3419,N_3608);
nor U4088 (N_4088,N_3526,N_3452);
xor U4089 (N_4089,N_3101,N_3749);
or U4090 (N_4090,N_3514,N_3324);
xnor U4091 (N_4091,N_3144,N_3259);
nor U4092 (N_4092,N_3619,N_3941);
nor U4093 (N_4093,N_3842,N_3377);
xnor U4094 (N_4094,N_3106,N_3306);
xnor U4095 (N_4095,N_2648,N_3386);
nor U4096 (N_4096,N_3295,N_2643);
nand U4097 (N_4097,N_3916,N_2964);
nor U4098 (N_4098,N_3908,N_2469);
and U4099 (N_4099,N_3547,N_3243);
or U4100 (N_4100,N_2514,N_2378);
nand U4101 (N_4101,N_2367,N_3983);
nand U4102 (N_4102,N_3262,N_2554);
nor U4103 (N_4103,N_3002,N_3188);
nand U4104 (N_4104,N_3008,N_3302);
or U4105 (N_4105,N_3479,N_2047);
nor U4106 (N_4106,N_2194,N_3426);
or U4107 (N_4107,N_2689,N_3904);
and U4108 (N_4108,N_2844,N_3130);
nor U4109 (N_4109,N_2482,N_2880);
or U4110 (N_4110,N_3043,N_3126);
nor U4111 (N_4111,N_3775,N_3598);
or U4112 (N_4112,N_2013,N_3654);
nor U4113 (N_4113,N_2679,N_3444);
or U4114 (N_4114,N_2780,N_3484);
nor U4115 (N_4115,N_2238,N_2155);
nor U4116 (N_4116,N_3128,N_2922);
xnor U4117 (N_4117,N_2986,N_3124);
nor U4118 (N_4118,N_3843,N_3997);
nand U4119 (N_4119,N_2183,N_2057);
or U4120 (N_4120,N_3544,N_2963);
and U4121 (N_4121,N_2496,N_3210);
nand U4122 (N_4122,N_2756,N_3552);
or U4123 (N_4123,N_2815,N_2162);
and U4124 (N_4124,N_2779,N_2297);
nand U4125 (N_4125,N_3355,N_2601);
and U4126 (N_4126,N_3999,N_2611);
nand U4127 (N_4127,N_2791,N_2649);
nor U4128 (N_4128,N_2332,N_3072);
nor U4129 (N_4129,N_2971,N_3353);
nand U4130 (N_4130,N_3753,N_3873);
or U4131 (N_4131,N_2308,N_3989);
nor U4132 (N_4132,N_3572,N_3211);
nand U4133 (N_4133,N_2783,N_3518);
nor U4134 (N_4134,N_2385,N_3770);
or U4135 (N_4135,N_2852,N_2706);
nor U4136 (N_4136,N_3623,N_2462);
nor U4137 (N_4137,N_3686,N_3528);
or U4138 (N_4138,N_3836,N_3453);
nor U4139 (N_4139,N_2937,N_2240);
xor U4140 (N_4140,N_2171,N_3769);
nand U4141 (N_4141,N_3123,N_3574);
and U4142 (N_4142,N_3033,N_2312);
nand U4143 (N_4143,N_3938,N_3812);
nor U4144 (N_4144,N_2438,N_3995);
and U4145 (N_4145,N_2625,N_3253);
nand U4146 (N_4146,N_3500,N_3629);
nand U4147 (N_4147,N_3886,N_3089);
xor U4148 (N_4148,N_3740,N_3456);
nand U4149 (N_4149,N_2990,N_3617);
nand U4150 (N_4150,N_2956,N_2172);
nor U4151 (N_4151,N_2981,N_3342);
and U4152 (N_4152,N_2446,N_2128);
xor U4153 (N_4153,N_3914,N_2590);
or U4154 (N_4154,N_3557,N_2778);
or U4155 (N_4155,N_3231,N_2492);
nand U4156 (N_4156,N_2144,N_3746);
or U4157 (N_4157,N_2527,N_3918);
nand U4158 (N_4158,N_3609,N_3663);
and U4159 (N_4159,N_3196,N_3809);
or U4160 (N_4160,N_2106,N_3599);
and U4161 (N_4161,N_3146,N_3430);
nor U4162 (N_4162,N_3760,N_3312);
nand U4163 (N_4163,N_2872,N_2141);
or U4164 (N_4164,N_2997,N_3421);
and U4165 (N_4165,N_2111,N_3473);
nor U4166 (N_4166,N_2548,N_2824);
nand U4167 (N_4167,N_3199,N_2301);
xor U4168 (N_4168,N_2614,N_2932);
nand U4169 (N_4169,N_3763,N_3704);
and U4170 (N_4170,N_2959,N_3934);
or U4171 (N_4171,N_2763,N_2698);
and U4172 (N_4172,N_3055,N_3114);
or U4173 (N_4173,N_3534,N_3650);
nor U4174 (N_4174,N_3058,N_2835);
and U4175 (N_4175,N_2870,N_3855);
xor U4176 (N_4176,N_3469,N_3928);
and U4177 (N_4177,N_3154,N_3434);
and U4178 (N_4178,N_3052,N_3645);
nor U4179 (N_4179,N_3165,N_2213);
nand U4180 (N_4180,N_3857,N_2276);
and U4181 (N_4181,N_2020,N_2612);
or U4182 (N_4182,N_2004,N_2653);
nor U4183 (N_4183,N_2743,N_3620);
and U4184 (N_4184,N_3279,N_2443);
or U4185 (N_4185,N_2317,N_2565);
nor U4186 (N_4186,N_3376,N_3541);
nor U4187 (N_4187,N_2769,N_2353);
and U4188 (N_4188,N_3086,N_2840);
nand U4189 (N_4189,N_3054,N_2909);
or U4190 (N_4190,N_3283,N_3074);
nor U4191 (N_4191,N_3671,N_3863);
and U4192 (N_4192,N_2998,N_3251);
nor U4193 (N_4193,N_2864,N_2861);
nor U4194 (N_4194,N_3604,N_2992);
or U4195 (N_4195,N_2231,N_3230);
nand U4196 (N_4196,N_3764,N_2010);
xnor U4197 (N_4197,N_2887,N_2015);
nand U4198 (N_4198,N_3815,N_2747);
nor U4199 (N_4199,N_2250,N_2884);
nor U4200 (N_4200,N_3647,N_2092);
nand U4201 (N_4201,N_2900,N_3796);
and U4202 (N_4202,N_2502,N_3284);
nor U4203 (N_4203,N_2571,N_3177);
nor U4204 (N_4204,N_3725,N_2904);
nand U4205 (N_4205,N_3313,N_3925);
or U4206 (N_4206,N_2982,N_3463);
nor U4207 (N_4207,N_2588,N_3432);
nand U4208 (N_4208,N_3734,N_2040);
xor U4209 (N_4209,N_2775,N_3851);
nand U4210 (N_4210,N_2475,N_2977);
and U4211 (N_4211,N_3411,N_3830);
nor U4212 (N_4212,N_2256,N_3111);
nand U4213 (N_4213,N_3991,N_3571);
nor U4214 (N_4214,N_2728,N_2605);
nand U4215 (N_4215,N_2715,N_3078);
nor U4216 (N_4216,N_2674,N_3751);
and U4217 (N_4217,N_2987,N_3193);
and U4218 (N_4218,N_3238,N_2849);
xnor U4219 (N_4219,N_3733,N_2658);
nand U4220 (N_4220,N_2999,N_3367);
nand U4221 (N_4221,N_3723,N_2316);
and U4222 (N_4222,N_2483,N_2823);
nor U4223 (N_4223,N_3994,N_2967);
nor U4224 (N_4224,N_2820,N_2923);
and U4225 (N_4225,N_3973,N_2827);
and U4226 (N_4226,N_3304,N_3911);
xor U4227 (N_4227,N_2461,N_2871);
or U4228 (N_4228,N_3269,N_2044);
nand U4229 (N_4229,N_3583,N_3612);
xnor U4230 (N_4230,N_2448,N_2893);
nor U4231 (N_4231,N_3718,N_2755);
nand U4232 (N_4232,N_3618,N_2022);
and U4233 (N_4233,N_3201,N_2158);
or U4234 (N_4234,N_2340,N_3362);
nor U4235 (N_4235,N_3881,N_2730);
nor U4236 (N_4236,N_3835,N_2652);
and U4237 (N_4237,N_3792,N_2076);
or U4238 (N_4238,N_3441,N_2676);
nor U4239 (N_4239,N_3820,N_3053);
nand U4240 (N_4240,N_3540,N_2832);
and U4241 (N_4241,N_3121,N_2116);
and U4242 (N_4242,N_3314,N_3626);
or U4243 (N_4243,N_2404,N_3073);
nor U4244 (N_4244,N_2073,N_3800);
nor U4245 (N_4245,N_2321,N_2479);
nand U4246 (N_4246,N_2449,N_2629);
or U4247 (N_4247,N_3900,N_2809);
or U4248 (N_4248,N_3783,N_3589);
nor U4249 (N_4249,N_2828,N_2237);
nand U4250 (N_4250,N_2627,N_2161);
xnor U4251 (N_4251,N_2733,N_2090);
and U4252 (N_4252,N_3678,N_3093);
and U4253 (N_4253,N_3163,N_3443);
nand U4254 (N_4254,N_3197,N_3020);
or U4255 (N_4255,N_2693,N_2694);
or U4256 (N_4256,N_3102,N_3680);
nor U4257 (N_4257,N_3627,N_2039);
or U4258 (N_4258,N_2534,N_3992);
nand U4259 (N_4259,N_2936,N_3600);
nand U4260 (N_4260,N_2968,N_2669);
or U4261 (N_4261,N_3624,N_3927);
and U4262 (N_4262,N_2043,N_3982);
or U4263 (N_4263,N_3532,N_3841);
and U4264 (N_4264,N_2558,N_2442);
or U4265 (N_4265,N_3169,N_2196);
or U4266 (N_4266,N_3412,N_3460);
nor U4267 (N_4267,N_2193,N_2243);
or U4268 (N_4268,N_3859,N_2170);
and U4269 (N_4269,N_3272,N_2935);
xor U4270 (N_4270,N_2729,N_2452);
nand U4271 (N_4271,N_3031,N_3451);
xnor U4272 (N_4272,N_2721,N_3184);
or U4273 (N_4273,N_2642,N_2929);
nand U4274 (N_4274,N_3967,N_2314);
and U4275 (N_4275,N_2300,N_3545);
and U4276 (N_4276,N_3176,N_2683);
or U4277 (N_4277,N_3707,N_2917);
or U4278 (N_4278,N_2067,N_3781);
and U4279 (N_4279,N_2499,N_2651);
nand U4280 (N_4280,N_2224,N_2529);
nand U4281 (N_4281,N_2825,N_3507);
and U4282 (N_4282,N_2408,N_3401);
or U4283 (N_4283,N_3850,N_2184);
nand U4284 (N_4284,N_3290,N_3565);
nand U4285 (N_4285,N_2948,N_3709);
or U4286 (N_4286,N_2875,N_3457);
nand U4287 (N_4287,N_2341,N_3027);
xnor U4288 (N_4288,N_3694,N_3985);
nand U4289 (N_4289,N_2618,N_3611);
nor U4290 (N_4290,N_3375,N_2702);
nor U4291 (N_4291,N_3385,N_2445);
nand U4292 (N_4292,N_2101,N_2320);
and U4293 (N_4293,N_2071,N_2188);
nor U4294 (N_4294,N_3039,N_2028);
or U4295 (N_4295,N_3716,N_2850);
and U4296 (N_4296,N_2168,N_3592);
nand U4297 (N_4297,N_3661,N_3024);
and U4298 (N_4298,N_3838,N_2275);
and U4299 (N_4299,N_2227,N_2953);
nor U4300 (N_4300,N_3228,N_3805);
and U4301 (N_4301,N_3736,N_2038);
nand U4302 (N_4302,N_3428,N_2790);
and U4303 (N_4303,N_3673,N_2933);
and U4304 (N_4304,N_2530,N_2916);
xnor U4305 (N_4305,N_2281,N_3926);
nand U4306 (N_4306,N_3013,N_3461);
nand U4307 (N_4307,N_3071,N_2007);
nand U4308 (N_4308,N_3964,N_2481);
or U4309 (N_4309,N_2773,N_2374);
nor U4310 (N_4310,N_3676,N_3966);
or U4311 (N_4311,N_3391,N_3814);
and U4312 (N_4312,N_3573,N_3383);
or U4313 (N_4313,N_2813,N_2412);
or U4314 (N_4314,N_2716,N_3549);
nand U4315 (N_4315,N_2053,N_2380);
and U4316 (N_4316,N_3282,N_3693);
xnor U4317 (N_4317,N_2665,N_2306);
nor U4318 (N_4318,N_2381,N_3782);
nand U4319 (N_4319,N_2124,N_3372);
nand U4320 (N_4320,N_2687,N_3810);
nand U4321 (N_4321,N_2115,N_3402);
xor U4322 (N_4322,N_2352,N_3333);
or U4323 (N_4323,N_2647,N_2711);
or U4324 (N_4324,N_2700,N_3961);
xor U4325 (N_4325,N_3640,N_2635);
and U4326 (N_4326,N_2265,N_2841);
or U4327 (N_4327,N_2789,N_3798);
xor U4328 (N_4328,N_2459,N_2949);
and U4329 (N_4329,N_2902,N_3637);
or U4330 (N_4330,N_2150,N_3275);
and U4331 (N_4331,N_2863,N_2965);
and U4332 (N_4332,N_2050,N_2091);
or U4333 (N_4333,N_2019,N_2387);
and U4334 (N_4334,N_3254,N_3168);
or U4335 (N_4335,N_3665,N_2899);
or U4336 (N_4336,N_2328,N_2697);
and U4337 (N_4337,N_2012,N_3266);
or U4338 (N_4338,N_3164,N_2418);
nand U4339 (N_4339,N_3097,N_3728);
nor U4340 (N_4340,N_2616,N_3195);
nand U4341 (N_4341,N_3423,N_2860);
xnor U4342 (N_4342,N_3980,N_3465);
xnor U4343 (N_4343,N_2422,N_2803);
or U4344 (N_4344,N_3012,N_3030);
nand U4345 (N_4345,N_3110,N_2808);
and U4346 (N_4346,N_3591,N_2456);
nor U4347 (N_4347,N_3294,N_2768);
or U4348 (N_4348,N_3668,N_2567);
xnor U4349 (N_4349,N_2264,N_2405);
or U4350 (N_4350,N_3041,N_2166);
and U4351 (N_4351,N_3420,N_3424);
and U4352 (N_4352,N_3799,N_3368);
xnor U4353 (N_4353,N_3986,N_3776);
or U4354 (N_4354,N_3656,N_3642);
nor U4355 (N_4355,N_3326,N_2985);
and U4356 (N_4356,N_3511,N_3603);
or U4357 (N_4357,N_2544,N_2097);
nor U4358 (N_4358,N_3777,N_3625);
or U4359 (N_4359,N_2401,N_3521);
or U4360 (N_4360,N_2500,N_2726);
or U4361 (N_4361,N_2239,N_2920);
and U4362 (N_4362,N_3754,N_3179);
and U4363 (N_4363,N_2819,N_3489);
nor U4364 (N_4364,N_2123,N_2371);
xnor U4365 (N_4365,N_3536,N_2303);
nand U4366 (N_4366,N_3771,N_2346);
nand U4367 (N_4367,N_3699,N_2200);
nor U4368 (N_4368,N_2030,N_3570);
xnor U4369 (N_4369,N_3028,N_3389);
xnor U4370 (N_4370,N_2754,N_3587);
xor U4371 (N_4371,N_3194,N_3406);
and U4372 (N_4372,N_2624,N_2862);
xnor U4373 (N_4373,N_3975,N_2682);
nor U4374 (N_4374,N_2621,N_2562);
nor U4375 (N_4375,N_2309,N_3834);
and U4376 (N_4376,N_2704,N_3582);
nand U4377 (N_4377,N_3566,N_2498);
and U4378 (N_4378,N_2178,N_2131);
nor U4379 (N_4379,N_2451,N_3149);
nand U4380 (N_4380,N_3267,N_3327);
nor U4381 (N_4381,N_3517,N_2259);
nor U4382 (N_4382,N_2688,N_3175);
and U4383 (N_4383,N_2228,N_2018);
nor U4384 (N_4384,N_3595,N_3882);
nand U4385 (N_4385,N_2397,N_2447);
nand U4386 (N_4386,N_2415,N_2298);
or U4387 (N_4387,N_3223,N_2058);
nor U4388 (N_4388,N_2262,N_2581);
nor U4389 (N_4389,N_3958,N_2615);
nand U4390 (N_4390,N_3352,N_3268);
nor U4391 (N_4391,N_3328,N_3960);
nand U4392 (N_4392,N_3436,N_2520);
nand U4393 (N_4393,N_3067,N_3447);
xor U4394 (N_4394,N_3229,N_2951);
and U4395 (N_4395,N_3765,N_2632);
or U4396 (N_4396,N_3122,N_3956);
nand U4397 (N_4397,N_2425,N_2838);
or U4398 (N_4398,N_2304,N_2656);
nor U4399 (N_4399,N_2532,N_3150);
nor U4400 (N_4400,N_3712,N_2455);
nand U4401 (N_4401,N_2427,N_2660);
nand U4402 (N_4402,N_3940,N_3091);
nand U4403 (N_4403,N_2191,N_3658);
nor U4404 (N_4404,N_2145,N_3399);
nand U4405 (N_4405,N_2557,N_2709);
and U4406 (N_4406,N_3095,N_3567);
and U4407 (N_4407,N_3879,N_2727);
or U4408 (N_4408,N_3060,N_3166);
or U4409 (N_4409,N_3527,N_2045);
nand U4410 (N_4410,N_3050,N_3875);
nor U4411 (N_4411,N_3246,N_3833);
or U4412 (N_4412,N_2718,N_2433);
nor U4413 (N_4413,N_2181,N_2345);
and U4414 (N_4414,N_2771,N_2630);
nand U4415 (N_4415,N_2753,N_2253);
and U4416 (N_4416,N_2543,N_3331);
and U4417 (N_4417,N_2424,N_3903);
or U4418 (N_4418,N_3017,N_3633);
nand U4419 (N_4419,N_3010,N_3757);
nor U4420 (N_4420,N_2740,N_3329);
and U4421 (N_4421,N_3183,N_3837);
and U4422 (N_4422,N_2041,N_2804);
xor U4423 (N_4423,N_3032,N_2757);
or U4424 (N_4424,N_2258,N_3047);
nand U4425 (N_4425,N_2277,N_3520);
xor U4426 (N_4426,N_3705,N_3794);
xnor U4427 (N_4427,N_3156,N_2016);
or U4428 (N_4428,N_2407,N_2176);
nand U4429 (N_4429,N_3902,N_3801);
or U4430 (N_4430,N_3576,N_2761);
or U4431 (N_4431,N_2552,N_2504);
nor U4432 (N_4432,N_3025,N_3561);
nor U4433 (N_4433,N_2323,N_2218);
and U4434 (N_4434,N_2831,N_3239);
nor U4435 (N_4435,N_3363,N_2025);
and U4436 (N_4436,N_2112,N_3148);
or U4437 (N_4437,N_2559,N_2536);
and U4438 (N_4438,N_3454,N_2703);
or U4439 (N_4439,N_3803,N_3378);
nand U4440 (N_4440,N_3005,N_2147);
nand U4441 (N_4441,N_2506,N_2988);
and U4442 (N_4442,N_2048,N_3232);
nor U4443 (N_4443,N_3727,N_3438);
nor U4444 (N_4444,N_3706,N_3929);
and U4445 (N_4445,N_2160,N_2122);
nand U4446 (N_4446,N_2355,N_3788);
nand U4447 (N_4447,N_2384,N_2357);
nor U4448 (N_4448,N_2881,N_3867);
or U4449 (N_4449,N_2856,N_3319);
and U4450 (N_4450,N_2035,N_2069);
and U4451 (N_4451,N_2006,N_2393);
nand U4452 (N_4452,N_2081,N_2473);
nand U4453 (N_4453,N_2724,N_2329);
nor U4454 (N_4454,N_3993,N_3245);
nor U4455 (N_4455,N_3691,N_3840);
or U4456 (N_4456,N_2569,N_3227);
and U4457 (N_4457,N_2710,N_3252);
nor U4458 (N_4458,N_2389,N_2607);
or U4459 (N_4459,N_3543,N_2468);
xnor U4460 (N_4460,N_2059,N_2105);
and U4461 (N_4461,N_2005,N_3685);
nand U4462 (N_4462,N_2394,N_3936);
or U4463 (N_4463,N_2528,N_3679);
or U4464 (N_4464,N_2503,N_2280);
and U4465 (N_4465,N_3493,N_2372);
or U4466 (N_4466,N_3081,N_3322);
nor U4467 (N_4467,N_2118,N_2961);
and U4468 (N_4468,N_3215,N_2869);
or U4469 (N_4469,N_3159,N_2033);
and U4470 (N_4470,N_3448,N_2600);
and U4471 (N_4471,N_2282,N_2386);
nor U4472 (N_4472,N_3731,N_3737);
and U4473 (N_4473,N_2157,N_2735);
and U4474 (N_4474,N_3066,N_2739);
nor U4475 (N_4475,N_2608,N_2509);
nor U4476 (N_4476,N_2192,N_3970);
nor U4477 (N_4477,N_2540,N_3427);
nor U4478 (N_4478,N_3158,N_2675);
and U4479 (N_4479,N_3495,N_3933);
nor U4480 (N_4480,N_2766,N_2219);
nor U4481 (N_4481,N_2088,N_2913);
and U4482 (N_4482,N_2480,N_2001);
or U4483 (N_4483,N_2731,N_2234);
or U4484 (N_4484,N_2587,N_2930);
and U4485 (N_4485,N_3096,N_2290);
nor U4486 (N_4486,N_2051,N_2926);
nor U4487 (N_4487,N_3040,N_2205);
and U4488 (N_4488,N_2190,N_3242);
and U4489 (N_4489,N_2670,N_2749);
nand U4490 (N_4490,N_3698,N_2351);
and U4491 (N_4491,N_2344,N_2491);
or U4492 (N_4492,N_3924,N_2969);
nand U4493 (N_4493,N_3845,N_3098);
and U4494 (N_4494,N_3652,N_3458);
nand U4495 (N_4495,N_2003,N_3203);
nand U4496 (N_4496,N_2511,N_3046);
or U4497 (N_4497,N_2725,N_3400);
nor U4498 (N_4498,N_3713,N_3387);
or U4499 (N_4499,N_2596,N_2737);
nand U4500 (N_4500,N_2911,N_3720);
nor U4501 (N_4501,N_2400,N_3371);
nand U4502 (N_4502,N_3786,N_3296);
nor U4503 (N_4503,N_2098,N_2945);
xnor U4504 (N_4504,N_3581,N_3289);
or U4505 (N_4505,N_2547,N_2066);
and U4506 (N_4506,N_2722,N_2247);
or U4507 (N_4507,N_3827,N_2132);
nand U4508 (N_4508,N_2661,N_3417);
and U4509 (N_4509,N_3987,N_3653);
or U4510 (N_4510,N_2087,N_2634);
and U4511 (N_4511,N_3807,N_3062);
nor U4512 (N_4512,N_3657,N_3015);
nand U4513 (N_4513,N_3752,N_2620);
nor U4514 (N_4514,N_3813,N_2944);
or U4515 (N_4515,N_2758,N_2759);
and U4516 (N_4516,N_2251,N_3622);
and U4517 (N_4517,N_3346,N_3261);
and U4518 (N_4518,N_3644,N_3088);
or U4519 (N_4519,N_3271,N_3832);
xnor U4520 (N_4520,N_3059,N_2127);
or U4521 (N_4521,N_3405,N_2767);
and U4522 (N_4522,N_3649,N_2242);
and U4523 (N_4523,N_3117,N_2350);
or U4524 (N_4524,N_3335,N_3293);
xnor U4525 (N_4525,N_3743,N_3337);
and U4526 (N_4526,N_2244,N_3191);
or U4527 (N_4527,N_2799,N_3950);
and U4528 (N_4528,N_3988,N_2515);
nand U4529 (N_4529,N_2268,N_3120);
and U4530 (N_4530,N_2667,N_2894);
nor U4531 (N_4531,N_2232,N_2440);
or U4532 (N_4532,N_2858,N_2847);
nand U4533 (N_4533,N_3009,N_2885);
nand U4534 (N_4534,N_2912,N_2542);
nand U4535 (N_4535,N_2851,N_3019);
nand U4536 (N_4536,N_2008,N_2074);
xor U4537 (N_4537,N_2299,N_2545);
and U4538 (N_4538,N_3898,N_3404);
nand U4539 (N_4539,N_3048,N_3351);
and U4540 (N_4540,N_2889,N_2079);
and U4541 (N_4541,N_2198,N_3866);
nor U4542 (N_4542,N_3955,N_2151);
nand U4543 (N_4543,N_3118,N_2905);
nor U4544 (N_4544,N_2390,N_3937);
nor U4545 (N_4545,N_3889,N_3064);
xnor U4546 (N_4546,N_2593,N_2036);
nand U4547 (N_4547,N_3880,N_2622);
or U4548 (N_4548,N_3236,N_3299);
nand U4549 (N_4549,N_2555,N_3381);
or U4550 (N_4550,N_2288,N_3014);
nand U4551 (N_4551,N_2639,N_3710);
nand U4552 (N_4552,N_2444,N_3212);
nand U4553 (N_4553,N_2398,N_2720);
or U4554 (N_4554,N_3614,N_3482);
nand U4555 (N_4555,N_3641,N_3745);
xor U4556 (N_4556,N_3684,N_3505);
xnor U4557 (N_4557,N_2093,N_2741);
nand U4558 (N_4558,N_3806,N_3481);
and U4559 (N_4559,N_2524,N_2221);
or U4560 (N_4560,N_2886,N_3802);
and U4561 (N_4561,N_3689,N_2650);
nand U4562 (N_4562,N_3131,N_2508);
nand U4563 (N_4563,N_2541,N_2373);
and U4564 (N_4564,N_2927,N_3366);
nand U4565 (N_4565,N_3695,N_2531);
and U4566 (N_4566,N_3586,N_3893);
nor U4567 (N_4567,N_3065,N_3946);
nor U4568 (N_4568,N_3761,N_2984);
or U4569 (N_4569,N_2453,N_2426);
xnor U4570 (N_4570,N_2626,N_2082);
or U4571 (N_4571,N_2671,N_2319);
and U4572 (N_4572,N_2736,N_2797);
nand U4573 (N_4573,N_3316,N_2865);
and U4574 (N_4574,N_2261,N_2263);
nor U4575 (N_4575,N_2484,N_2310);
nor U4576 (N_4576,N_3655,N_2583);
xnor U4577 (N_4577,N_3681,N_2023);
xor U4578 (N_4578,N_2829,N_3860);
or U4579 (N_4579,N_3359,N_2845);
or U4580 (N_4580,N_2970,N_3160);
xor U4581 (N_4581,N_2343,N_3852);
nand U4582 (N_4582,N_2362,N_3116);
or U4583 (N_4583,N_3648,N_3410);
nor U4584 (N_4584,N_3082,N_3555);
xnor U4585 (N_4585,N_3719,N_2266);
nor U4586 (N_4586,N_3667,N_2095);
nand U4587 (N_4587,N_3510,N_2089);
nand U4588 (N_4588,N_2203,N_2631);
or U4589 (N_4589,N_3748,N_2295);
or U4590 (N_4590,N_2952,N_2096);
nor U4591 (N_4591,N_2454,N_2663);
and U4592 (N_4592,N_2765,N_3466);
and U4593 (N_4593,N_3153,N_2286);
xnor U4594 (N_4594,N_2026,N_3112);
and U4595 (N_4595,N_2267,N_2817);
and U4596 (N_4596,N_2855,N_3061);
or U4597 (N_4597,N_3906,N_3202);
xnor U4598 (N_4598,N_2644,N_2207);
nor U4599 (N_4599,N_2738,N_3467);
and U4600 (N_4600,N_3049,N_3891);
nand U4601 (N_4601,N_2843,N_3659);
nor U4602 (N_4602,N_3471,N_3501);
and U4603 (N_4603,N_2510,N_3418);
and U4604 (N_4604,N_3172,N_2853);
nor U4605 (N_4605,N_2938,N_2179);
xor U4606 (N_4606,N_3247,N_2560);
nor U4607 (N_4607,N_3077,N_3550);
or U4608 (N_4608,N_2110,N_2934);
nor U4609 (N_4609,N_3811,N_2955);
nor U4610 (N_4610,N_2979,N_3315);
nand U4611 (N_4611,N_3415,N_2714);
xnor U4612 (N_4612,N_3477,N_3949);
nor U4613 (N_4613,N_3739,N_3022);
or U4614 (N_4614,N_2235,N_3332);
xor U4615 (N_4615,N_3189,N_2812);
xnor U4616 (N_4616,N_2338,N_3498);
or U4617 (N_4617,N_2229,N_3286);
nor U4618 (N_4618,N_2167,N_2748);
and U4619 (N_4619,N_2439,N_2678);
nand U4620 (N_4620,N_3963,N_2493);
nand U4621 (N_4621,N_3535,N_2888);
xor U4622 (N_4622,N_3726,N_3590);
nand U4623 (N_4623,N_3330,N_2077);
nand U4624 (N_4624,N_3439,N_3145);
and U4625 (N_4625,N_2795,N_2180);
nor U4626 (N_4626,N_3957,N_3741);
nand U4627 (N_4627,N_2972,N_2209);
nand U4628 (N_4628,N_2821,N_2460);
and U4629 (N_4629,N_2471,N_3285);
or U4630 (N_4630,N_2100,N_2195);
and U4631 (N_4631,N_3396,N_3225);
nand U4632 (N_4632,N_3459,N_3155);
or U4633 (N_4633,N_2148,N_3513);
or U4634 (N_4634,N_3491,N_2140);
nor U4635 (N_4635,N_3478,N_2633);
or U4636 (N_4636,N_2646,N_2573);
and U4637 (N_4637,N_3729,N_2662);
nand U4638 (N_4638,N_2349,N_2943);
nand U4639 (N_4639,N_3990,N_2640);
nor U4640 (N_4640,N_2287,N_2153);
or U4641 (N_4641,N_2417,N_3178);
nor U4642 (N_4642,N_3666,N_2525);
nor U4643 (N_4643,N_3379,N_3133);
or U4644 (N_4644,N_3701,N_3790);
nand U4645 (N_4645,N_3615,N_2490);
nor U4646 (N_4646,N_2062,N_2826);
nand U4647 (N_4647,N_3414,N_2719);
nand U4648 (N_4648,N_3601,N_3023);
nor U4649 (N_4649,N_2556,N_2574);
nand U4650 (N_4650,N_3486,N_2377);
or U4651 (N_4651,N_2084,N_3651);
nor U4652 (N_4652,N_3255,N_3674);
or U4653 (N_4653,N_2024,N_3895);
and U4654 (N_4654,N_3825,N_3374);
nor U4655 (N_4655,N_2293,N_2364);
and U4656 (N_4656,N_2873,N_2202);
nand U4657 (N_4657,N_3206,N_3523);
nor U4658 (N_4658,N_3278,N_3056);
nand U4659 (N_4659,N_2094,N_2011);
or U4660 (N_4660,N_2908,N_2713);
and U4661 (N_4661,N_2419,N_2197);
or U4662 (N_4662,N_2836,N_2336);
or U4663 (N_4663,N_2973,N_3298);
nand U4664 (N_4664,N_3190,N_2278);
xor U4665 (N_4665,N_3356,N_2918);
and U4666 (N_4666,N_2579,N_2796);
or U4667 (N_4667,N_2363,N_2497);
xnor U4668 (N_4668,N_2368,N_2659);
nor U4669 (N_4669,N_2211,N_3136);
nor U4670 (N_4670,N_2996,N_3808);
nor U4671 (N_4671,N_3977,N_2708);
or U4672 (N_4672,N_3789,N_3470);
xor U4673 (N_4673,N_3948,N_2921);
nor U4674 (N_4674,N_2604,N_3369);
or U4675 (N_4675,N_2108,N_3142);
nand U4676 (N_4676,N_2962,N_2037);
nand U4677 (N_4677,N_3735,N_2925);
or U4678 (N_4678,N_2859,N_3584);
or U4679 (N_4679,N_3876,N_3200);
nor U4680 (N_4680,N_2488,N_3358);
and U4681 (N_4681,N_2793,N_3951);
and U4682 (N_4682,N_3750,N_3092);
nor U4683 (N_4683,N_2402,N_3021);
nor U4684 (N_4684,N_3475,N_3099);
nand U4685 (N_4685,N_2135,N_2339);
nand U4686 (N_4686,N_2465,N_3766);
nand U4687 (N_4687,N_3497,N_2810);
and U4688 (N_4688,N_2489,N_3998);
nor U4689 (N_4689,N_3488,N_2522);
xnor U4690 (N_4690,N_2940,N_2572);
and U4691 (N_4691,N_3672,N_2568);
xor U4692 (N_4692,N_3100,N_2891);
nor U4693 (N_4693,N_3696,N_3562);
or U4694 (N_4694,N_2575,N_3797);
nand U4695 (N_4695,N_2107,N_3241);
nand U4696 (N_4696,N_2685,N_3487);
or U4697 (N_4697,N_2208,N_3361);
nor U4698 (N_4698,N_3455,N_3732);
nand U4699 (N_4699,N_2347,N_3533);
and U4700 (N_4700,N_2214,N_3677);
and U4701 (N_4701,N_3472,N_2271);
nand U4702 (N_4702,N_2991,N_2673);
or U4703 (N_4703,N_2878,N_3433);
or U4704 (N_4704,N_3742,N_3393);
or U4705 (N_4705,N_2563,N_2901);
nor U4706 (N_4706,N_2915,N_2201);
nand U4707 (N_4707,N_2126,N_3036);
and U4708 (N_4708,N_3631,N_3321);
or U4709 (N_4709,N_3431,N_2787);
or U4710 (N_4710,N_3636,N_2117);
and U4711 (N_4711,N_2744,N_3888);
nor U4712 (N_4712,N_2764,N_2315);
nand U4713 (N_4713,N_2610,N_3140);
or U4714 (N_4714,N_2248,N_2361);
nand U4715 (N_4715,N_3292,N_3462);
or U4716 (N_4716,N_2657,N_3152);
and U4717 (N_4717,N_2335,N_2217);
or U4718 (N_4718,N_3143,N_2690);
nand U4719 (N_4719,N_3670,N_3884);
nand U4720 (N_4720,N_3000,N_3942);
nand U4721 (N_4721,N_2877,N_3016);
xor U4722 (N_4722,N_2411,N_2113);
or U4723 (N_4723,N_2745,N_3537);
nand U4724 (N_4724,N_3274,N_2584);
xnor U4725 (N_4725,N_3578,N_2874);
xnor U4726 (N_4726,N_2842,N_2762);
and U4727 (N_4727,N_2392,N_3530);
nor U4728 (N_4728,N_3529,N_2619);
nor U4729 (N_4729,N_2421,N_3085);
and U4730 (N_4730,N_2960,N_3182);
or U4731 (N_4731,N_2606,N_3822);
xnor U4732 (N_4732,N_2245,N_3409);
nand U4733 (N_4733,N_2830,N_3675);
or U4734 (N_4734,N_3350,N_3692);
nor U4735 (N_4735,N_2029,N_3070);
and U4736 (N_4736,N_3847,N_3494);
or U4737 (N_4737,N_2599,N_2326);
nand U4738 (N_4738,N_3213,N_3310);
and U4739 (N_4739,N_3890,N_3817);
or U4740 (N_4740,N_2435,N_3554);
and U4741 (N_4741,N_3407,N_3628);
nand U4742 (N_4742,N_3198,N_3209);
and U4743 (N_4743,N_3912,N_3688);
nand U4744 (N_4744,N_2002,N_2539);
nand U4745 (N_4745,N_3422,N_3577);
nand U4746 (N_4746,N_2549,N_3785);
xor U4747 (N_4747,N_3192,N_2342);
and U4748 (N_4748,N_3721,N_3162);
xnor U4749 (N_4749,N_3492,N_3744);
nor U4750 (N_4750,N_2156,N_2487);
and U4751 (N_4751,N_2994,N_2063);
nor U4752 (N_4752,N_2285,N_3826);
nand U4753 (N_4753,N_2358,N_2236);
nor U4754 (N_4754,N_3542,N_3224);
nand U4755 (N_4755,N_3887,N_2538);
and U4756 (N_4756,N_3504,N_3094);
or U4757 (N_4757,N_2307,N_2655);
nor U4758 (N_4758,N_2457,N_2924);
and U4759 (N_4759,N_3580,N_3660);
nand U4760 (N_4760,N_2423,N_3161);
and U4761 (N_4761,N_3256,N_2645);
and U4762 (N_4762,N_2816,N_2519);
xnor U4763 (N_4763,N_3038,N_3248);
nor U4764 (N_4764,N_2958,N_3397);
or U4765 (N_4765,N_2553,N_3506);
or U4766 (N_4766,N_2109,N_3509);
xor U4767 (N_4767,N_2000,N_3755);
nor U4768 (N_4768,N_2760,N_3018);
and U4769 (N_4769,N_2177,N_2723);
nand U4770 (N_4770,N_3167,N_2811);
nand U4771 (N_4771,N_3357,N_3939);
xnor U4772 (N_4772,N_3853,N_2595);
nand U4773 (N_4773,N_2983,N_2995);
or U4774 (N_4774,N_2330,N_3264);
and U4775 (N_4775,N_2366,N_2467);
nor U4776 (N_4776,N_2325,N_3839);
or U4777 (N_4777,N_3907,N_2292);
or U4778 (N_4778,N_3711,N_2215);
or U4779 (N_4779,N_2681,N_3923);
and U4780 (N_4780,N_3502,N_3700);
or U4781 (N_4781,N_2199,N_3395);
or U4782 (N_4782,N_2220,N_2260);
or U4783 (N_4783,N_3344,N_2169);
nand U4784 (N_4784,N_3483,N_2876);
nor U4785 (N_4785,N_3610,N_2494);
or U4786 (N_4786,N_2814,N_2785);
nand U4787 (N_4787,N_3930,N_2428);
and U4788 (N_4788,N_2879,N_2149);
nand U4789 (N_4789,N_3080,N_3795);
and U4790 (N_4790,N_2185,N_3952);
or U4791 (N_4791,N_3607,N_2331);
or U4792 (N_4792,N_3083,N_3425);
nand U4793 (N_4793,N_2406,N_3910);
or U4794 (N_4794,N_3113,N_3784);
nand U4795 (N_4795,N_3287,N_2914);
and U4796 (N_4796,N_2103,N_2233);
and U4797 (N_4797,N_3068,N_2882);
and U4798 (N_4798,N_3125,N_2897);
or U4799 (N_4799,N_3263,N_3878);
nand U4800 (N_4800,N_3515,N_3288);
nand U4801 (N_4801,N_3563,N_2327);
or U4802 (N_4802,N_2136,N_3187);
or U4803 (N_4803,N_3297,N_3336);
nor U4804 (N_4804,N_2822,N_3045);
nor U4805 (N_4805,N_2476,N_3007);
nand U4806 (N_4806,N_3921,N_2638);
and U4807 (N_4807,N_3630,N_3115);
or U4808 (N_4808,N_2495,N_2458);
or U4809 (N_4809,N_3821,N_2078);
nor U4810 (N_4810,N_3664,N_3490);
nand U4811 (N_4811,N_3758,N_3922);
nor U4812 (N_4812,N_3702,N_3001);
nand U4813 (N_4813,N_3181,N_2976);
and U4814 (N_4814,N_2950,N_2255);
nor U4815 (N_4815,N_2980,N_3717);
nand U4816 (N_4816,N_3323,N_2370);
or U4817 (N_4817,N_2684,N_3216);
and U4818 (N_4818,N_3828,N_2225);
or U4819 (N_4819,N_3147,N_3069);
or U4820 (N_4820,N_3476,N_2032);
nand U4821 (N_4821,N_3968,N_2356);
or U4822 (N_4822,N_2989,N_2974);
or U4823 (N_4823,N_2907,N_2410);
or U4824 (N_4824,N_2142,N_3205);
nand U4825 (N_4825,N_3011,N_2919);
nor U4826 (N_4826,N_3485,N_3217);
and U4827 (N_4827,N_2173,N_2892);
nand U4828 (N_4828,N_2434,N_3697);
nand U4829 (N_4829,N_3558,N_2441);
and U4830 (N_4830,N_2732,N_3208);
and U4831 (N_4831,N_3634,N_3347);
and U4832 (N_4832,N_3870,N_3265);
nor U4833 (N_4833,N_2296,N_2121);
and U4834 (N_4834,N_3403,N_3079);
xnor U4835 (N_4835,N_2139,N_3793);
or U4836 (N_4836,N_3138,N_3560);
or U4837 (N_4837,N_3037,N_3105);
nor U4838 (N_4838,N_2699,N_2717);
nand U4839 (N_4839,N_3564,N_3303);
nand U4840 (N_4840,N_3687,N_2931);
xnor U4841 (N_4841,N_3613,N_3273);
nand U4842 (N_4842,N_2686,N_2485);
and U4843 (N_4843,N_3575,N_3551);
or U4844 (N_4844,N_2083,N_2705);
and U4845 (N_4845,N_3508,N_2868);
or U4846 (N_4846,N_2395,N_3974);
xor U4847 (N_4847,N_2270,N_3585);
nor U4848 (N_4848,N_3635,N_3003);
xnor U4849 (N_4849,N_2334,N_2431);
xor U4850 (N_4850,N_2249,N_3141);
nor U4851 (N_4851,N_2978,N_2589);
or U4852 (N_4852,N_2257,N_2031);
nand U4853 (N_4853,N_2046,N_3935);
or U4854 (N_4854,N_2486,N_2284);
xnor U4855 (N_4855,N_3173,N_3787);
nand U4856 (N_4856,N_2668,N_3408);
and U4857 (N_4857,N_2666,N_3683);
and U4858 (N_4858,N_2597,N_2975);
and U4859 (N_4859,N_2437,N_3730);
and U4860 (N_4860,N_3318,N_3818);
and U4861 (N_4861,N_3877,N_2792);
or U4862 (N_4862,N_2085,N_3442);
and U4863 (N_4863,N_2712,N_3104);
nor U4864 (N_4864,N_2279,N_2080);
nor U4865 (N_4865,N_2580,N_2751);
xor U4866 (N_4866,N_3237,N_3222);
nand U4867 (N_4867,N_2561,N_3915);
nand U4868 (N_4868,N_3639,N_2052);
xnor U4869 (N_4869,N_3250,N_3139);
nor U4870 (N_4870,N_3596,N_3524);
xor U4871 (N_4871,N_2505,N_2664);
or U4872 (N_4872,N_3006,N_2839);
or U4873 (N_4873,N_2291,N_2337);
and U4874 (N_4874,N_2641,N_3714);
nor U4875 (N_4875,N_3365,N_2055);
nor U4876 (N_4876,N_3416,N_3819);
nand U4877 (N_4877,N_2223,N_2895);
and U4878 (N_4878,N_3233,N_3854);
or U4879 (N_4879,N_3856,N_3954);
or U4880 (N_4880,N_2383,N_2636);
nand U4881 (N_4881,N_2770,N_3738);
and U4882 (N_4882,N_2501,N_2086);
xnor U4883 (N_4883,N_3107,N_2230);
nor U4884 (N_4884,N_3917,N_2399);
and U4885 (N_4885,N_3309,N_3320);
and U4886 (N_4886,N_3280,N_3643);
nand U4887 (N_4887,N_2154,N_3151);
or U4888 (N_4888,N_3325,N_3349);
and U4889 (N_4889,N_3823,N_3388);
or U4890 (N_4890,N_3848,N_3135);
nor U4891 (N_4891,N_2707,N_3569);
nand U4892 (N_4892,N_2910,N_3602);
xor U4893 (N_4893,N_2466,N_2613);
and U4894 (N_4894,N_3972,N_3075);
nor U4895 (N_4895,N_3762,N_3969);
nor U4896 (N_4896,N_3516,N_3249);
nand U4897 (N_4897,N_2289,N_3553);
nor U4898 (N_4898,N_3311,N_3772);
nor U4899 (N_4899,N_2414,N_2318);
and U4900 (N_4900,N_3959,N_3445);
nor U4901 (N_4901,N_2129,N_2577);
xor U4902 (N_4902,N_3480,N_3076);
nand U4903 (N_4903,N_3435,N_2294);
and U4904 (N_4904,N_3892,N_3382);
xor U4905 (N_4905,N_3662,N_3343);
nand U4906 (N_4906,N_3345,N_3831);
nand U4907 (N_4907,N_2333,N_3090);
nor U4908 (N_4908,N_2594,N_3499);
and U4909 (N_4909,N_2833,N_3338);
or U4910 (N_4910,N_2617,N_2472);
and U4911 (N_4911,N_3464,N_3538);
nand U4912 (N_4912,N_3767,N_2576);
or U4913 (N_4913,N_3953,N_2750);
nand U4914 (N_4914,N_3260,N_2742);
nor U4915 (N_4915,N_2592,N_2890);
nand U4916 (N_4916,N_3869,N_2396);
and U4917 (N_4917,N_2348,N_2138);
and U4918 (N_4918,N_3947,N_2772);
or U4919 (N_4919,N_3932,N_2099);
or U4920 (N_4920,N_2939,N_3219);
nor U4921 (N_4921,N_2807,N_3244);
xnor U4922 (N_4922,N_2946,N_2695);
nand U4923 (N_4923,N_2222,N_3759);
nor U4924 (N_4924,N_3317,N_3026);
or U4925 (N_4925,N_2837,N_3340);
nor U4926 (N_4926,N_2009,N_3380);
nor U4927 (N_4927,N_2182,N_2311);
and U4928 (N_4928,N_3594,N_3897);
nand U4929 (N_4929,N_2034,N_2526);
or U4930 (N_4930,N_2189,N_2175);
nor U4931 (N_4931,N_3185,N_3868);
nand U4932 (N_4932,N_2777,N_2060);
and U4933 (N_4933,N_3588,N_3945);
nand U4934 (N_4934,N_3905,N_2125);
xor U4935 (N_4935,N_3901,N_2578);
and U4936 (N_4936,N_2313,N_2164);
nand U4937 (N_4937,N_2014,N_2365);
and U4938 (N_4938,N_2782,N_2564);
or U4939 (N_4939,N_2146,N_2119);
and U4940 (N_4940,N_2696,N_2413);
and U4941 (N_4941,N_3109,N_2274);
or U4942 (N_4942,N_3370,N_3301);
nor U4943 (N_4943,N_3690,N_3593);
and U4944 (N_4944,N_3621,N_3108);
nand U4945 (N_4945,N_3568,N_3446);
nor U4946 (N_4946,N_3861,N_3307);
nand U4947 (N_4947,N_3978,N_3226);
xnor U4948 (N_4948,N_2379,N_3300);
nand U4949 (N_4949,N_2463,N_2788);
or U4950 (N_4950,N_2903,N_3221);
xor U4951 (N_4951,N_2867,N_2602);
nor U4952 (N_4952,N_3044,N_2802);
or U4953 (N_4953,N_3756,N_3638);
nand U4954 (N_4954,N_2137,N_3384);
nor U4955 (N_4955,N_3034,N_2430);
or U4956 (N_4956,N_3979,N_2941);
or U4957 (N_4957,N_3548,N_3137);
nor U4958 (N_4958,N_2102,N_3390);
or U4959 (N_4959,N_2065,N_2806);
xor U4960 (N_4960,N_3063,N_2834);
nor U4961 (N_4961,N_3778,N_2302);
and U4962 (N_4962,N_3214,N_3816);
nor U4963 (N_4963,N_3057,N_2603);
nor U4964 (N_4964,N_2784,N_3220);
nand U4965 (N_4965,N_3270,N_3862);
or U4966 (N_4966,N_3512,N_2957);
and U4967 (N_4967,N_2801,N_3976);
nand U4968 (N_4968,N_2186,N_2075);
nor U4969 (N_4969,N_3519,N_3474);
nor U4970 (N_4970,N_2993,N_2252);
nor U4971 (N_4971,N_2734,N_2054);
nand U4972 (N_4972,N_3218,N_3258);
nor U4973 (N_4973,N_2928,N_3235);
or U4974 (N_4974,N_3134,N_2241);
nand U4975 (N_4975,N_3747,N_2570);
nor U4976 (N_4976,N_2609,N_3281);
xnor U4977 (N_4977,N_3437,N_2068);
nand U4978 (N_4978,N_2049,N_2550);
nand U4979 (N_4979,N_3171,N_2746);
and U4980 (N_4980,N_2391,N_2774);
nand U4981 (N_4981,N_3207,N_2056);
nor U4982 (N_4982,N_3708,N_3525);
xnor U4983 (N_4983,N_3546,N_2551);
nand U4984 (N_4984,N_2134,N_2420);
and U4985 (N_4985,N_2246,N_2133);
and U4986 (N_4986,N_2546,N_3186);
nand U4987 (N_4987,N_2947,N_2883);
or U4988 (N_4988,N_2470,N_2672);
or U4989 (N_4989,N_2409,N_3885);
or U4990 (N_4990,N_3392,N_3180);
and U4991 (N_4991,N_3276,N_2104);
xor U4992 (N_4992,N_2523,N_3646);
nand U4993 (N_4993,N_2477,N_2432);
nor U4994 (N_4994,N_2474,N_2206);
or U4995 (N_4995,N_3883,N_2781);
nand U4996 (N_4996,N_2906,N_2537);
nand U4997 (N_4997,N_3413,N_3348);
and U4998 (N_4998,N_2360,N_3981);
and U4999 (N_4999,N_3354,N_3871);
and U5000 (N_5000,N_3607,N_3898);
or U5001 (N_5001,N_3698,N_3991);
nor U5002 (N_5002,N_3569,N_3846);
xnor U5003 (N_5003,N_3340,N_2624);
nand U5004 (N_5004,N_3997,N_3050);
and U5005 (N_5005,N_2619,N_3433);
and U5006 (N_5006,N_3377,N_2090);
and U5007 (N_5007,N_2730,N_3723);
or U5008 (N_5008,N_3855,N_2800);
nand U5009 (N_5009,N_2641,N_2877);
or U5010 (N_5010,N_2354,N_2289);
and U5011 (N_5011,N_2062,N_3696);
or U5012 (N_5012,N_3766,N_2474);
or U5013 (N_5013,N_2018,N_3285);
nor U5014 (N_5014,N_2611,N_2985);
nand U5015 (N_5015,N_3987,N_2488);
and U5016 (N_5016,N_3593,N_2765);
nand U5017 (N_5017,N_2676,N_2770);
and U5018 (N_5018,N_2971,N_3586);
or U5019 (N_5019,N_2952,N_3779);
and U5020 (N_5020,N_3767,N_3550);
xor U5021 (N_5021,N_3814,N_3219);
and U5022 (N_5022,N_2037,N_3464);
and U5023 (N_5023,N_2642,N_3069);
nor U5024 (N_5024,N_2696,N_3181);
nand U5025 (N_5025,N_3407,N_2646);
nand U5026 (N_5026,N_2678,N_2298);
nand U5027 (N_5027,N_3277,N_3585);
and U5028 (N_5028,N_3654,N_3428);
nor U5029 (N_5029,N_3733,N_2250);
nor U5030 (N_5030,N_3942,N_2717);
nand U5031 (N_5031,N_3967,N_2915);
and U5032 (N_5032,N_3652,N_3698);
or U5033 (N_5033,N_2685,N_2951);
nor U5034 (N_5034,N_3844,N_2166);
xor U5035 (N_5035,N_3298,N_3567);
nand U5036 (N_5036,N_3609,N_3807);
nor U5037 (N_5037,N_2885,N_2375);
and U5038 (N_5038,N_3651,N_2327);
or U5039 (N_5039,N_3827,N_3459);
and U5040 (N_5040,N_3308,N_2247);
nand U5041 (N_5041,N_2802,N_2136);
and U5042 (N_5042,N_3616,N_3388);
nor U5043 (N_5043,N_2030,N_3973);
nand U5044 (N_5044,N_2231,N_2621);
nand U5045 (N_5045,N_2896,N_3059);
xnor U5046 (N_5046,N_2698,N_3308);
and U5047 (N_5047,N_3680,N_2193);
and U5048 (N_5048,N_3303,N_3440);
nor U5049 (N_5049,N_3285,N_3084);
nand U5050 (N_5050,N_3867,N_2043);
nor U5051 (N_5051,N_2452,N_2403);
and U5052 (N_5052,N_2190,N_2778);
nor U5053 (N_5053,N_3536,N_3022);
or U5054 (N_5054,N_2670,N_2280);
nand U5055 (N_5055,N_2771,N_2891);
xnor U5056 (N_5056,N_3725,N_2238);
or U5057 (N_5057,N_3678,N_2640);
nor U5058 (N_5058,N_3553,N_3619);
nand U5059 (N_5059,N_2176,N_3467);
or U5060 (N_5060,N_3616,N_2882);
xnor U5061 (N_5061,N_2196,N_3579);
nand U5062 (N_5062,N_3070,N_3071);
nor U5063 (N_5063,N_3319,N_3594);
nor U5064 (N_5064,N_3192,N_2579);
nor U5065 (N_5065,N_3857,N_2430);
or U5066 (N_5066,N_3107,N_3628);
nand U5067 (N_5067,N_2840,N_3347);
nand U5068 (N_5068,N_2777,N_2073);
nand U5069 (N_5069,N_2136,N_3447);
nor U5070 (N_5070,N_3937,N_3204);
and U5071 (N_5071,N_2801,N_2743);
xor U5072 (N_5072,N_3701,N_2799);
nor U5073 (N_5073,N_2276,N_2722);
and U5074 (N_5074,N_3157,N_2251);
nor U5075 (N_5075,N_3767,N_3351);
nor U5076 (N_5076,N_3951,N_2388);
and U5077 (N_5077,N_3387,N_3389);
or U5078 (N_5078,N_3334,N_2380);
and U5079 (N_5079,N_3074,N_2216);
nor U5080 (N_5080,N_2604,N_3082);
and U5081 (N_5081,N_3376,N_2987);
xor U5082 (N_5082,N_3456,N_2601);
nand U5083 (N_5083,N_2599,N_3800);
and U5084 (N_5084,N_3329,N_3977);
nor U5085 (N_5085,N_3519,N_2134);
nor U5086 (N_5086,N_2625,N_2802);
nand U5087 (N_5087,N_3099,N_2114);
and U5088 (N_5088,N_2426,N_3994);
nor U5089 (N_5089,N_2015,N_3196);
or U5090 (N_5090,N_2632,N_3671);
nor U5091 (N_5091,N_3620,N_3870);
nand U5092 (N_5092,N_3499,N_2701);
or U5093 (N_5093,N_2110,N_3889);
nand U5094 (N_5094,N_3920,N_2188);
nor U5095 (N_5095,N_2488,N_3660);
and U5096 (N_5096,N_3130,N_2156);
and U5097 (N_5097,N_3766,N_3241);
nor U5098 (N_5098,N_2946,N_2310);
and U5099 (N_5099,N_2110,N_3280);
xnor U5100 (N_5100,N_3149,N_3049);
nor U5101 (N_5101,N_3800,N_3166);
nand U5102 (N_5102,N_3249,N_3628);
xor U5103 (N_5103,N_2509,N_2850);
nor U5104 (N_5104,N_3252,N_3204);
nand U5105 (N_5105,N_2168,N_2772);
nand U5106 (N_5106,N_2211,N_3660);
and U5107 (N_5107,N_3170,N_2293);
nand U5108 (N_5108,N_2751,N_2071);
or U5109 (N_5109,N_3381,N_2481);
xnor U5110 (N_5110,N_3253,N_3683);
nor U5111 (N_5111,N_3539,N_3852);
and U5112 (N_5112,N_2758,N_2713);
and U5113 (N_5113,N_2726,N_3636);
or U5114 (N_5114,N_3666,N_3652);
nor U5115 (N_5115,N_3613,N_3729);
nor U5116 (N_5116,N_2727,N_2991);
nor U5117 (N_5117,N_3814,N_3282);
nand U5118 (N_5118,N_3683,N_3231);
xor U5119 (N_5119,N_3556,N_2676);
nand U5120 (N_5120,N_3551,N_3834);
and U5121 (N_5121,N_3114,N_2955);
nor U5122 (N_5122,N_2999,N_2953);
xnor U5123 (N_5123,N_3374,N_2466);
or U5124 (N_5124,N_3948,N_2715);
or U5125 (N_5125,N_3934,N_3452);
nand U5126 (N_5126,N_2663,N_2629);
nor U5127 (N_5127,N_2842,N_2743);
nor U5128 (N_5128,N_2569,N_3955);
nand U5129 (N_5129,N_2826,N_2128);
nor U5130 (N_5130,N_2263,N_2852);
xnor U5131 (N_5131,N_2949,N_3371);
or U5132 (N_5132,N_3929,N_2324);
and U5133 (N_5133,N_2224,N_2802);
or U5134 (N_5134,N_2391,N_2668);
nand U5135 (N_5135,N_3339,N_2759);
or U5136 (N_5136,N_2582,N_2868);
xnor U5137 (N_5137,N_2222,N_3221);
nand U5138 (N_5138,N_3788,N_3495);
xor U5139 (N_5139,N_2961,N_2192);
nand U5140 (N_5140,N_2222,N_3462);
nand U5141 (N_5141,N_3381,N_2948);
xor U5142 (N_5142,N_2306,N_3874);
nand U5143 (N_5143,N_2832,N_3932);
nand U5144 (N_5144,N_2764,N_3571);
xor U5145 (N_5145,N_3424,N_2871);
nor U5146 (N_5146,N_2121,N_2812);
nand U5147 (N_5147,N_3994,N_2109);
or U5148 (N_5148,N_2028,N_2293);
nand U5149 (N_5149,N_3767,N_3676);
or U5150 (N_5150,N_3571,N_2211);
nand U5151 (N_5151,N_3311,N_3598);
nor U5152 (N_5152,N_2920,N_2627);
and U5153 (N_5153,N_3347,N_2263);
nand U5154 (N_5154,N_2768,N_2205);
and U5155 (N_5155,N_2382,N_2653);
nand U5156 (N_5156,N_2744,N_2489);
nor U5157 (N_5157,N_3581,N_3063);
nand U5158 (N_5158,N_2565,N_3665);
nand U5159 (N_5159,N_2670,N_3963);
nand U5160 (N_5160,N_2773,N_2422);
xor U5161 (N_5161,N_2404,N_2925);
nor U5162 (N_5162,N_3376,N_3357);
nand U5163 (N_5163,N_2845,N_3256);
nor U5164 (N_5164,N_3051,N_3514);
nand U5165 (N_5165,N_2314,N_2910);
or U5166 (N_5166,N_3175,N_3786);
nand U5167 (N_5167,N_2019,N_3862);
nand U5168 (N_5168,N_2105,N_3470);
and U5169 (N_5169,N_3745,N_3983);
nand U5170 (N_5170,N_2747,N_3609);
or U5171 (N_5171,N_3482,N_2260);
and U5172 (N_5172,N_3416,N_2945);
xnor U5173 (N_5173,N_3783,N_2326);
or U5174 (N_5174,N_2429,N_2654);
or U5175 (N_5175,N_3647,N_3285);
nand U5176 (N_5176,N_2654,N_3017);
and U5177 (N_5177,N_2215,N_3553);
or U5178 (N_5178,N_2446,N_3942);
xor U5179 (N_5179,N_3262,N_2056);
and U5180 (N_5180,N_3416,N_3751);
and U5181 (N_5181,N_2722,N_3462);
and U5182 (N_5182,N_3198,N_3804);
or U5183 (N_5183,N_3082,N_2117);
and U5184 (N_5184,N_3399,N_3726);
xor U5185 (N_5185,N_3760,N_2427);
nand U5186 (N_5186,N_3839,N_2750);
nand U5187 (N_5187,N_2385,N_2617);
xor U5188 (N_5188,N_2934,N_3774);
nand U5189 (N_5189,N_2424,N_3221);
nand U5190 (N_5190,N_2207,N_2640);
and U5191 (N_5191,N_3054,N_2880);
nand U5192 (N_5192,N_3570,N_3082);
nor U5193 (N_5193,N_2856,N_2217);
and U5194 (N_5194,N_3698,N_2615);
nor U5195 (N_5195,N_3653,N_3693);
nand U5196 (N_5196,N_3173,N_3328);
nand U5197 (N_5197,N_3836,N_3311);
or U5198 (N_5198,N_2205,N_2119);
or U5199 (N_5199,N_2166,N_2079);
nand U5200 (N_5200,N_2097,N_3544);
xor U5201 (N_5201,N_3649,N_3360);
and U5202 (N_5202,N_2490,N_2162);
nand U5203 (N_5203,N_2155,N_3076);
or U5204 (N_5204,N_3761,N_2009);
nand U5205 (N_5205,N_2694,N_3893);
or U5206 (N_5206,N_2515,N_3055);
nor U5207 (N_5207,N_2373,N_2614);
or U5208 (N_5208,N_2138,N_3616);
nor U5209 (N_5209,N_3130,N_3559);
xnor U5210 (N_5210,N_2565,N_2568);
nor U5211 (N_5211,N_2447,N_2115);
nand U5212 (N_5212,N_2344,N_2346);
and U5213 (N_5213,N_3071,N_3020);
nor U5214 (N_5214,N_3122,N_2906);
or U5215 (N_5215,N_2668,N_2528);
and U5216 (N_5216,N_3564,N_2047);
xor U5217 (N_5217,N_2591,N_2783);
nand U5218 (N_5218,N_3928,N_2703);
nand U5219 (N_5219,N_2989,N_2644);
xnor U5220 (N_5220,N_2071,N_3877);
xor U5221 (N_5221,N_2238,N_3443);
nor U5222 (N_5222,N_2752,N_2349);
nand U5223 (N_5223,N_2352,N_3150);
nand U5224 (N_5224,N_3546,N_2786);
nand U5225 (N_5225,N_2786,N_2774);
and U5226 (N_5226,N_3839,N_2260);
nand U5227 (N_5227,N_2859,N_2280);
and U5228 (N_5228,N_3289,N_3948);
and U5229 (N_5229,N_3864,N_3423);
xnor U5230 (N_5230,N_2050,N_3562);
or U5231 (N_5231,N_3427,N_2693);
nor U5232 (N_5232,N_3700,N_3355);
and U5233 (N_5233,N_3479,N_2014);
or U5234 (N_5234,N_3639,N_3846);
nor U5235 (N_5235,N_2682,N_2229);
and U5236 (N_5236,N_3832,N_3399);
and U5237 (N_5237,N_3288,N_2098);
nand U5238 (N_5238,N_3040,N_3007);
and U5239 (N_5239,N_3415,N_3240);
xnor U5240 (N_5240,N_2287,N_2044);
nand U5241 (N_5241,N_2886,N_3763);
or U5242 (N_5242,N_2638,N_3796);
nor U5243 (N_5243,N_2697,N_3188);
and U5244 (N_5244,N_3641,N_3111);
xnor U5245 (N_5245,N_2673,N_3964);
or U5246 (N_5246,N_3094,N_3643);
nor U5247 (N_5247,N_2431,N_3367);
nor U5248 (N_5248,N_3751,N_2047);
and U5249 (N_5249,N_2791,N_3600);
or U5250 (N_5250,N_2250,N_3348);
or U5251 (N_5251,N_2661,N_3938);
or U5252 (N_5252,N_2637,N_3572);
nor U5253 (N_5253,N_3104,N_3185);
and U5254 (N_5254,N_2950,N_2767);
xor U5255 (N_5255,N_2415,N_3928);
nor U5256 (N_5256,N_3923,N_2658);
and U5257 (N_5257,N_2949,N_3869);
nand U5258 (N_5258,N_2516,N_2943);
nand U5259 (N_5259,N_3119,N_2648);
or U5260 (N_5260,N_2558,N_2515);
or U5261 (N_5261,N_3081,N_3375);
xnor U5262 (N_5262,N_3496,N_3627);
or U5263 (N_5263,N_3826,N_3077);
nor U5264 (N_5264,N_2944,N_2614);
and U5265 (N_5265,N_3834,N_2267);
and U5266 (N_5266,N_3764,N_3706);
xor U5267 (N_5267,N_3216,N_3236);
nand U5268 (N_5268,N_3760,N_3647);
nand U5269 (N_5269,N_3494,N_3953);
nand U5270 (N_5270,N_2762,N_2847);
nor U5271 (N_5271,N_2637,N_2291);
nor U5272 (N_5272,N_3982,N_2714);
or U5273 (N_5273,N_3719,N_2807);
and U5274 (N_5274,N_2825,N_2148);
xnor U5275 (N_5275,N_3362,N_3971);
xor U5276 (N_5276,N_3903,N_3900);
and U5277 (N_5277,N_3006,N_3646);
or U5278 (N_5278,N_3940,N_3347);
nor U5279 (N_5279,N_3045,N_3377);
nand U5280 (N_5280,N_2454,N_2146);
and U5281 (N_5281,N_3174,N_3261);
nor U5282 (N_5282,N_2440,N_3041);
nand U5283 (N_5283,N_3442,N_3314);
nor U5284 (N_5284,N_3183,N_2381);
and U5285 (N_5285,N_3473,N_3133);
nand U5286 (N_5286,N_3415,N_3234);
nor U5287 (N_5287,N_2897,N_3281);
and U5288 (N_5288,N_3458,N_2226);
and U5289 (N_5289,N_2699,N_3544);
or U5290 (N_5290,N_2281,N_3468);
and U5291 (N_5291,N_3180,N_3116);
nor U5292 (N_5292,N_2370,N_2114);
or U5293 (N_5293,N_3060,N_3670);
nor U5294 (N_5294,N_3830,N_3589);
and U5295 (N_5295,N_2344,N_2119);
nor U5296 (N_5296,N_3049,N_2028);
or U5297 (N_5297,N_3651,N_2053);
and U5298 (N_5298,N_2120,N_2921);
and U5299 (N_5299,N_2353,N_3521);
and U5300 (N_5300,N_2870,N_2961);
xnor U5301 (N_5301,N_2146,N_3374);
nand U5302 (N_5302,N_2478,N_2353);
and U5303 (N_5303,N_3720,N_2776);
nor U5304 (N_5304,N_3360,N_2829);
nor U5305 (N_5305,N_2512,N_2507);
and U5306 (N_5306,N_2943,N_2369);
nor U5307 (N_5307,N_3376,N_3633);
xor U5308 (N_5308,N_2241,N_3929);
or U5309 (N_5309,N_3341,N_3696);
nor U5310 (N_5310,N_3391,N_2104);
nor U5311 (N_5311,N_2781,N_2653);
nand U5312 (N_5312,N_2772,N_3854);
or U5313 (N_5313,N_3364,N_3370);
nand U5314 (N_5314,N_2446,N_3478);
nand U5315 (N_5315,N_2546,N_2413);
xor U5316 (N_5316,N_3799,N_3674);
or U5317 (N_5317,N_2891,N_2527);
or U5318 (N_5318,N_3622,N_2827);
or U5319 (N_5319,N_3785,N_2625);
nor U5320 (N_5320,N_2111,N_2308);
nand U5321 (N_5321,N_2388,N_2882);
and U5322 (N_5322,N_3193,N_2095);
and U5323 (N_5323,N_3442,N_3749);
nor U5324 (N_5324,N_3748,N_2076);
and U5325 (N_5325,N_2413,N_3182);
nand U5326 (N_5326,N_2748,N_3771);
and U5327 (N_5327,N_2517,N_2416);
or U5328 (N_5328,N_3613,N_2797);
nor U5329 (N_5329,N_2311,N_3785);
or U5330 (N_5330,N_3381,N_3989);
and U5331 (N_5331,N_2918,N_3549);
or U5332 (N_5332,N_3853,N_2607);
nand U5333 (N_5333,N_3116,N_2826);
and U5334 (N_5334,N_3151,N_2489);
nand U5335 (N_5335,N_2367,N_3836);
and U5336 (N_5336,N_2585,N_2249);
and U5337 (N_5337,N_2527,N_2302);
nand U5338 (N_5338,N_2637,N_2025);
nor U5339 (N_5339,N_2520,N_2157);
nand U5340 (N_5340,N_3465,N_3143);
nor U5341 (N_5341,N_2907,N_3116);
nand U5342 (N_5342,N_3721,N_3201);
nand U5343 (N_5343,N_2651,N_3642);
and U5344 (N_5344,N_2635,N_3028);
or U5345 (N_5345,N_3226,N_3965);
nor U5346 (N_5346,N_3390,N_2670);
or U5347 (N_5347,N_3780,N_2840);
or U5348 (N_5348,N_2292,N_3691);
nand U5349 (N_5349,N_2882,N_2806);
and U5350 (N_5350,N_2044,N_3975);
or U5351 (N_5351,N_3090,N_3513);
nand U5352 (N_5352,N_2843,N_3097);
xor U5353 (N_5353,N_3252,N_2832);
xor U5354 (N_5354,N_3537,N_3635);
nand U5355 (N_5355,N_3670,N_3157);
and U5356 (N_5356,N_3682,N_3929);
nor U5357 (N_5357,N_2952,N_2996);
nand U5358 (N_5358,N_3645,N_2741);
nor U5359 (N_5359,N_3870,N_2274);
nand U5360 (N_5360,N_2625,N_2956);
nand U5361 (N_5361,N_2968,N_3231);
or U5362 (N_5362,N_3960,N_2813);
and U5363 (N_5363,N_2403,N_3373);
nand U5364 (N_5364,N_3507,N_3715);
nor U5365 (N_5365,N_3956,N_2236);
and U5366 (N_5366,N_2252,N_2876);
or U5367 (N_5367,N_3412,N_3527);
and U5368 (N_5368,N_2594,N_3735);
xor U5369 (N_5369,N_2462,N_2589);
xnor U5370 (N_5370,N_3732,N_2218);
or U5371 (N_5371,N_2565,N_3999);
nor U5372 (N_5372,N_2634,N_3084);
nor U5373 (N_5373,N_3596,N_2539);
xnor U5374 (N_5374,N_3742,N_3656);
nand U5375 (N_5375,N_3619,N_3784);
or U5376 (N_5376,N_3502,N_3163);
nor U5377 (N_5377,N_3265,N_2120);
or U5378 (N_5378,N_2334,N_2112);
nand U5379 (N_5379,N_3412,N_2334);
nor U5380 (N_5380,N_3708,N_3638);
or U5381 (N_5381,N_3943,N_2125);
and U5382 (N_5382,N_2673,N_3478);
nand U5383 (N_5383,N_3717,N_3205);
and U5384 (N_5384,N_3934,N_2640);
and U5385 (N_5385,N_2083,N_2449);
nor U5386 (N_5386,N_2563,N_3899);
nor U5387 (N_5387,N_3044,N_3129);
and U5388 (N_5388,N_2147,N_2994);
nand U5389 (N_5389,N_3078,N_2552);
and U5390 (N_5390,N_2982,N_3220);
and U5391 (N_5391,N_3759,N_3963);
nand U5392 (N_5392,N_2996,N_2197);
xnor U5393 (N_5393,N_3961,N_3976);
and U5394 (N_5394,N_3173,N_3155);
or U5395 (N_5395,N_3480,N_3608);
and U5396 (N_5396,N_2966,N_2559);
nor U5397 (N_5397,N_3784,N_2083);
and U5398 (N_5398,N_2779,N_2754);
nand U5399 (N_5399,N_2292,N_2770);
nor U5400 (N_5400,N_2493,N_2105);
or U5401 (N_5401,N_3413,N_2935);
xnor U5402 (N_5402,N_2730,N_3316);
and U5403 (N_5403,N_2514,N_3590);
nor U5404 (N_5404,N_3893,N_3592);
or U5405 (N_5405,N_2273,N_3710);
xnor U5406 (N_5406,N_3588,N_3402);
or U5407 (N_5407,N_2016,N_2050);
xor U5408 (N_5408,N_2887,N_3113);
and U5409 (N_5409,N_2253,N_2963);
or U5410 (N_5410,N_2175,N_2078);
or U5411 (N_5411,N_2526,N_3168);
nand U5412 (N_5412,N_2217,N_2553);
nand U5413 (N_5413,N_3258,N_3336);
nor U5414 (N_5414,N_3407,N_2230);
and U5415 (N_5415,N_2918,N_3505);
and U5416 (N_5416,N_2710,N_3473);
nand U5417 (N_5417,N_3765,N_2619);
or U5418 (N_5418,N_3903,N_2646);
and U5419 (N_5419,N_2368,N_3421);
nand U5420 (N_5420,N_2925,N_2553);
nand U5421 (N_5421,N_2494,N_3157);
and U5422 (N_5422,N_3425,N_3090);
nor U5423 (N_5423,N_2409,N_2589);
nor U5424 (N_5424,N_3794,N_2692);
and U5425 (N_5425,N_3063,N_3629);
nor U5426 (N_5426,N_2097,N_3334);
xor U5427 (N_5427,N_3402,N_3335);
nand U5428 (N_5428,N_3585,N_3806);
or U5429 (N_5429,N_3597,N_2851);
nand U5430 (N_5430,N_3726,N_2949);
nand U5431 (N_5431,N_2595,N_2894);
nand U5432 (N_5432,N_2684,N_2372);
nor U5433 (N_5433,N_3295,N_2380);
and U5434 (N_5434,N_2155,N_2747);
nor U5435 (N_5435,N_2557,N_2584);
and U5436 (N_5436,N_2959,N_2804);
or U5437 (N_5437,N_2567,N_2147);
or U5438 (N_5438,N_3229,N_3210);
nand U5439 (N_5439,N_3102,N_2962);
or U5440 (N_5440,N_3703,N_3033);
nand U5441 (N_5441,N_2695,N_3018);
or U5442 (N_5442,N_2729,N_2994);
nand U5443 (N_5443,N_2515,N_3016);
and U5444 (N_5444,N_2085,N_3701);
nand U5445 (N_5445,N_2071,N_3897);
nor U5446 (N_5446,N_2743,N_3033);
nand U5447 (N_5447,N_3587,N_3860);
nor U5448 (N_5448,N_3572,N_3406);
and U5449 (N_5449,N_3437,N_2409);
nor U5450 (N_5450,N_2976,N_2819);
nand U5451 (N_5451,N_2697,N_2727);
nor U5452 (N_5452,N_2675,N_3048);
xor U5453 (N_5453,N_3463,N_2116);
nand U5454 (N_5454,N_3404,N_2881);
nand U5455 (N_5455,N_2525,N_3849);
nor U5456 (N_5456,N_2301,N_3706);
or U5457 (N_5457,N_2652,N_2628);
nand U5458 (N_5458,N_2065,N_2034);
and U5459 (N_5459,N_3168,N_2808);
nand U5460 (N_5460,N_2487,N_2809);
nand U5461 (N_5461,N_2525,N_2495);
xnor U5462 (N_5462,N_2522,N_2447);
nand U5463 (N_5463,N_3531,N_3149);
nor U5464 (N_5464,N_3362,N_3194);
and U5465 (N_5465,N_2815,N_3219);
nand U5466 (N_5466,N_3588,N_2251);
or U5467 (N_5467,N_2969,N_3757);
nor U5468 (N_5468,N_2914,N_2277);
nor U5469 (N_5469,N_2922,N_2843);
nor U5470 (N_5470,N_3137,N_2092);
or U5471 (N_5471,N_2875,N_2289);
nor U5472 (N_5472,N_3481,N_3539);
nand U5473 (N_5473,N_2152,N_3905);
or U5474 (N_5474,N_2123,N_3788);
nand U5475 (N_5475,N_3700,N_2020);
nor U5476 (N_5476,N_2874,N_2030);
nand U5477 (N_5477,N_2389,N_3123);
xnor U5478 (N_5478,N_2138,N_3986);
and U5479 (N_5479,N_3259,N_3072);
nor U5480 (N_5480,N_2095,N_2270);
nor U5481 (N_5481,N_2499,N_2711);
xor U5482 (N_5482,N_2384,N_2087);
nand U5483 (N_5483,N_2359,N_2756);
nand U5484 (N_5484,N_3403,N_2209);
nand U5485 (N_5485,N_2794,N_2049);
nor U5486 (N_5486,N_3527,N_2052);
nor U5487 (N_5487,N_2875,N_2229);
xor U5488 (N_5488,N_2548,N_3086);
or U5489 (N_5489,N_3095,N_2966);
and U5490 (N_5490,N_3461,N_3059);
nand U5491 (N_5491,N_2208,N_3405);
nand U5492 (N_5492,N_3675,N_2676);
nand U5493 (N_5493,N_2584,N_2549);
or U5494 (N_5494,N_2582,N_2579);
nand U5495 (N_5495,N_3365,N_2813);
nor U5496 (N_5496,N_2366,N_3517);
or U5497 (N_5497,N_2456,N_3944);
and U5498 (N_5498,N_2709,N_2840);
nor U5499 (N_5499,N_2794,N_3538);
nor U5500 (N_5500,N_3844,N_3928);
or U5501 (N_5501,N_2115,N_2937);
or U5502 (N_5502,N_2502,N_3005);
or U5503 (N_5503,N_2463,N_2580);
nand U5504 (N_5504,N_2931,N_3428);
nand U5505 (N_5505,N_2597,N_3011);
and U5506 (N_5506,N_2419,N_2714);
and U5507 (N_5507,N_3577,N_2301);
nor U5508 (N_5508,N_3237,N_3322);
and U5509 (N_5509,N_2030,N_3918);
and U5510 (N_5510,N_2022,N_3931);
nand U5511 (N_5511,N_2544,N_3071);
nor U5512 (N_5512,N_3613,N_3654);
and U5513 (N_5513,N_2511,N_3375);
or U5514 (N_5514,N_3165,N_2047);
xor U5515 (N_5515,N_2900,N_2769);
and U5516 (N_5516,N_3684,N_2561);
nand U5517 (N_5517,N_2528,N_2118);
and U5518 (N_5518,N_2158,N_2761);
nor U5519 (N_5519,N_2086,N_2466);
nand U5520 (N_5520,N_2975,N_2092);
and U5521 (N_5521,N_3739,N_2810);
or U5522 (N_5522,N_2730,N_3735);
nand U5523 (N_5523,N_2248,N_3169);
and U5524 (N_5524,N_3985,N_2608);
and U5525 (N_5525,N_3372,N_3904);
or U5526 (N_5526,N_3826,N_2592);
xnor U5527 (N_5527,N_3101,N_2600);
nor U5528 (N_5528,N_2683,N_2769);
nand U5529 (N_5529,N_2376,N_2087);
nor U5530 (N_5530,N_3913,N_2931);
nor U5531 (N_5531,N_3832,N_2417);
nor U5532 (N_5532,N_3382,N_2903);
nand U5533 (N_5533,N_3584,N_3082);
nand U5534 (N_5534,N_3760,N_2445);
or U5535 (N_5535,N_2718,N_3117);
nand U5536 (N_5536,N_3218,N_2944);
and U5537 (N_5537,N_3015,N_3726);
and U5538 (N_5538,N_3237,N_2296);
xnor U5539 (N_5539,N_2593,N_2993);
or U5540 (N_5540,N_3928,N_3403);
nor U5541 (N_5541,N_2705,N_2279);
nor U5542 (N_5542,N_3004,N_2468);
xnor U5543 (N_5543,N_2301,N_3148);
and U5544 (N_5544,N_2787,N_3956);
and U5545 (N_5545,N_2763,N_3983);
nor U5546 (N_5546,N_2276,N_2208);
nor U5547 (N_5547,N_2106,N_2218);
and U5548 (N_5548,N_3917,N_2217);
and U5549 (N_5549,N_3204,N_3777);
or U5550 (N_5550,N_2564,N_3859);
nor U5551 (N_5551,N_2029,N_2952);
nor U5552 (N_5552,N_2727,N_2966);
nor U5553 (N_5553,N_2639,N_3693);
or U5554 (N_5554,N_2391,N_3212);
nand U5555 (N_5555,N_2824,N_2172);
nor U5556 (N_5556,N_3097,N_3696);
xnor U5557 (N_5557,N_2936,N_3380);
nand U5558 (N_5558,N_2711,N_2954);
nand U5559 (N_5559,N_3817,N_3602);
or U5560 (N_5560,N_3661,N_2343);
nand U5561 (N_5561,N_3029,N_2856);
and U5562 (N_5562,N_2536,N_3860);
nor U5563 (N_5563,N_2385,N_3884);
or U5564 (N_5564,N_3694,N_3616);
or U5565 (N_5565,N_3044,N_3786);
or U5566 (N_5566,N_2789,N_3812);
nand U5567 (N_5567,N_2985,N_3329);
nand U5568 (N_5568,N_3735,N_3725);
nand U5569 (N_5569,N_3646,N_2066);
or U5570 (N_5570,N_3886,N_3334);
nand U5571 (N_5571,N_3825,N_2957);
xor U5572 (N_5572,N_3854,N_3452);
and U5573 (N_5573,N_2297,N_3852);
or U5574 (N_5574,N_3245,N_2722);
or U5575 (N_5575,N_3697,N_3633);
and U5576 (N_5576,N_3684,N_2515);
and U5577 (N_5577,N_2673,N_3091);
and U5578 (N_5578,N_3746,N_2205);
nor U5579 (N_5579,N_2233,N_3379);
and U5580 (N_5580,N_2975,N_3709);
or U5581 (N_5581,N_2539,N_3145);
nor U5582 (N_5582,N_3267,N_3536);
nor U5583 (N_5583,N_2887,N_2201);
and U5584 (N_5584,N_2658,N_2191);
or U5585 (N_5585,N_2504,N_2333);
nor U5586 (N_5586,N_2828,N_2999);
nand U5587 (N_5587,N_2567,N_3739);
nand U5588 (N_5588,N_2585,N_3452);
nand U5589 (N_5589,N_2974,N_3068);
nor U5590 (N_5590,N_2738,N_3130);
nor U5591 (N_5591,N_3887,N_2835);
nor U5592 (N_5592,N_2810,N_3206);
or U5593 (N_5593,N_2528,N_2270);
or U5594 (N_5594,N_3071,N_3133);
nand U5595 (N_5595,N_2089,N_2435);
or U5596 (N_5596,N_3474,N_2161);
nand U5597 (N_5597,N_2133,N_3857);
or U5598 (N_5598,N_3473,N_3730);
and U5599 (N_5599,N_3578,N_2503);
nor U5600 (N_5600,N_3589,N_3610);
nand U5601 (N_5601,N_3419,N_3677);
and U5602 (N_5602,N_3993,N_2695);
nand U5603 (N_5603,N_3770,N_3822);
nor U5604 (N_5604,N_2631,N_3056);
xor U5605 (N_5605,N_2473,N_3032);
or U5606 (N_5606,N_3359,N_2374);
and U5607 (N_5607,N_3865,N_3350);
and U5608 (N_5608,N_2592,N_2161);
nor U5609 (N_5609,N_2729,N_3798);
nor U5610 (N_5610,N_3519,N_2895);
or U5611 (N_5611,N_2895,N_3413);
nand U5612 (N_5612,N_2863,N_3881);
or U5613 (N_5613,N_2752,N_3260);
xor U5614 (N_5614,N_3881,N_2940);
nor U5615 (N_5615,N_3558,N_3294);
xnor U5616 (N_5616,N_2555,N_3437);
or U5617 (N_5617,N_2494,N_3926);
and U5618 (N_5618,N_3534,N_3386);
and U5619 (N_5619,N_2393,N_2009);
nand U5620 (N_5620,N_2766,N_2509);
nand U5621 (N_5621,N_3833,N_3842);
nor U5622 (N_5622,N_3626,N_3399);
nor U5623 (N_5623,N_3935,N_3449);
and U5624 (N_5624,N_2086,N_2697);
nor U5625 (N_5625,N_2023,N_3793);
nand U5626 (N_5626,N_3293,N_2916);
or U5627 (N_5627,N_2035,N_2529);
nor U5628 (N_5628,N_3986,N_2569);
nor U5629 (N_5629,N_2718,N_2371);
and U5630 (N_5630,N_2321,N_2872);
or U5631 (N_5631,N_2052,N_2653);
xor U5632 (N_5632,N_2665,N_2648);
nand U5633 (N_5633,N_3951,N_2632);
nand U5634 (N_5634,N_2047,N_3078);
nor U5635 (N_5635,N_2133,N_3308);
or U5636 (N_5636,N_3256,N_3166);
nand U5637 (N_5637,N_3273,N_3694);
nand U5638 (N_5638,N_2451,N_2145);
nand U5639 (N_5639,N_2184,N_2389);
and U5640 (N_5640,N_3580,N_2378);
nand U5641 (N_5641,N_3384,N_3925);
xor U5642 (N_5642,N_2168,N_3676);
nand U5643 (N_5643,N_3456,N_3632);
nand U5644 (N_5644,N_2567,N_3201);
nand U5645 (N_5645,N_2652,N_3281);
or U5646 (N_5646,N_3712,N_2830);
xnor U5647 (N_5647,N_2795,N_2789);
or U5648 (N_5648,N_3830,N_3053);
or U5649 (N_5649,N_3124,N_2175);
and U5650 (N_5650,N_2510,N_2339);
nand U5651 (N_5651,N_3188,N_3943);
or U5652 (N_5652,N_3074,N_2593);
nor U5653 (N_5653,N_3829,N_3999);
nor U5654 (N_5654,N_2742,N_2862);
nor U5655 (N_5655,N_3210,N_2861);
or U5656 (N_5656,N_2636,N_3706);
nand U5657 (N_5657,N_3888,N_2249);
or U5658 (N_5658,N_3913,N_3436);
nor U5659 (N_5659,N_3209,N_3378);
nor U5660 (N_5660,N_2180,N_2729);
or U5661 (N_5661,N_3715,N_3327);
and U5662 (N_5662,N_3011,N_2810);
or U5663 (N_5663,N_2765,N_3206);
nand U5664 (N_5664,N_2441,N_2311);
nand U5665 (N_5665,N_3785,N_2467);
and U5666 (N_5666,N_2085,N_3292);
nand U5667 (N_5667,N_2044,N_2080);
and U5668 (N_5668,N_2344,N_2838);
nand U5669 (N_5669,N_3351,N_3565);
nor U5670 (N_5670,N_3289,N_2070);
nor U5671 (N_5671,N_2846,N_2993);
or U5672 (N_5672,N_2799,N_2538);
nand U5673 (N_5673,N_2352,N_3789);
or U5674 (N_5674,N_2068,N_2421);
or U5675 (N_5675,N_2613,N_3504);
or U5676 (N_5676,N_2183,N_3479);
and U5677 (N_5677,N_2129,N_2681);
or U5678 (N_5678,N_2750,N_3528);
nor U5679 (N_5679,N_2242,N_3808);
or U5680 (N_5680,N_2717,N_3652);
and U5681 (N_5681,N_3269,N_2145);
or U5682 (N_5682,N_3742,N_2687);
nor U5683 (N_5683,N_2952,N_2664);
and U5684 (N_5684,N_3872,N_2710);
and U5685 (N_5685,N_3596,N_2734);
nand U5686 (N_5686,N_2502,N_2496);
nor U5687 (N_5687,N_2289,N_3052);
or U5688 (N_5688,N_3788,N_2861);
and U5689 (N_5689,N_2325,N_3681);
xnor U5690 (N_5690,N_3461,N_3297);
and U5691 (N_5691,N_2358,N_3538);
or U5692 (N_5692,N_3933,N_2529);
nor U5693 (N_5693,N_3391,N_2172);
nand U5694 (N_5694,N_2429,N_3029);
and U5695 (N_5695,N_2619,N_2899);
nand U5696 (N_5696,N_3271,N_2768);
nor U5697 (N_5697,N_2343,N_3614);
nand U5698 (N_5698,N_2707,N_2288);
nor U5699 (N_5699,N_2379,N_3703);
nand U5700 (N_5700,N_3333,N_2456);
nand U5701 (N_5701,N_2941,N_2569);
nor U5702 (N_5702,N_2538,N_2741);
and U5703 (N_5703,N_3051,N_2476);
nand U5704 (N_5704,N_3800,N_3969);
nand U5705 (N_5705,N_2007,N_2351);
xnor U5706 (N_5706,N_2275,N_3081);
and U5707 (N_5707,N_2905,N_2978);
and U5708 (N_5708,N_3956,N_2963);
nor U5709 (N_5709,N_3894,N_3699);
or U5710 (N_5710,N_2370,N_3617);
or U5711 (N_5711,N_2891,N_3357);
and U5712 (N_5712,N_3052,N_2366);
and U5713 (N_5713,N_3145,N_3751);
or U5714 (N_5714,N_3298,N_3860);
and U5715 (N_5715,N_2508,N_3951);
nor U5716 (N_5716,N_3790,N_2922);
nand U5717 (N_5717,N_3086,N_2695);
nor U5718 (N_5718,N_2044,N_3489);
nand U5719 (N_5719,N_3897,N_3536);
xnor U5720 (N_5720,N_3492,N_2283);
nor U5721 (N_5721,N_3491,N_3206);
nor U5722 (N_5722,N_3573,N_3168);
nand U5723 (N_5723,N_3482,N_3704);
nand U5724 (N_5724,N_3365,N_3190);
or U5725 (N_5725,N_3421,N_3574);
and U5726 (N_5726,N_3026,N_2306);
xor U5727 (N_5727,N_3988,N_2145);
or U5728 (N_5728,N_3079,N_3470);
or U5729 (N_5729,N_2147,N_2338);
nor U5730 (N_5730,N_3958,N_3366);
xnor U5731 (N_5731,N_2510,N_3535);
nor U5732 (N_5732,N_3592,N_3742);
or U5733 (N_5733,N_3534,N_2102);
nand U5734 (N_5734,N_3357,N_3320);
or U5735 (N_5735,N_2980,N_2042);
or U5736 (N_5736,N_2523,N_2761);
and U5737 (N_5737,N_3339,N_2627);
and U5738 (N_5738,N_2497,N_2992);
or U5739 (N_5739,N_2453,N_3032);
and U5740 (N_5740,N_3558,N_2204);
nand U5741 (N_5741,N_3130,N_2225);
nor U5742 (N_5742,N_2453,N_3128);
nor U5743 (N_5743,N_3753,N_3625);
nand U5744 (N_5744,N_3057,N_2199);
and U5745 (N_5745,N_3776,N_3171);
or U5746 (N_5746,N_3172,N_3395);
nor U5747 (N_5747,N_2139,N_2724);
nand U5748 (N_5748,N_2322,N_3816);
and U5749 (N_5749,N_3400,N_3988);
xnor U5750 (N_5750,N_3951,N_2883);
nor U5751 (N_5751,N_2148,N_3474);
xor U5752 (N_5752,N_3113,N_3259);
xor U5753 (N_5753,N_3467,N_3769);
nor U5754 (N_5754,N_2687,N_2745);
nand U5755 (N_5755,N_2259,N_3686);
nor U5756 (N_5756,N_3423,N_3293);
xor U5757 (N_5757,N_3684,N_2907);
or U5758 (N_5758,N_3067,N_2777);
and U5759 (N_5759,N_2824,N_2564);
nand U5760 (N_5760,N_2383,N_2785);
and U5761 (N_5761,N_2696,N_3086);
or U5762 (N_5762,N_2684,N_2266);
nor U5763 (N_5763,N_3837,N_3900);
or U5764 (N_5764,N_2443,N_3084);
xor U5765 (N_5765,N_2881,N_2938);
and U5766 (N_5766,N_3911,N_3941);
or U5767 (N_5767,N_3660,N_3037);
nand U5768 (N_5768,N_3197,N_3368);
nand U5769 (N_5769,N_3332,N_3672);
nand U5770 (N_5770,N_2515,N_3655);
or U5771 (N_5771,N_3054,N_2371);
xnor U5772 (N_5772,N_3837,N_3496);
xor U5773 (N_5773,N_3743,N_3732);
nand U5774 (N_5774,N_3891,N_2546);
or U5775 (N_5775,N_3761,N_3790);
and U5776 (N_5776,N_2938,N_2575);
nand U5777 (N_5777,N_3127,N_3028);
nor U5778 (N_5778,N_2096,N_2906);
and U5779 (N_5779,N_3093,N_2913);
and U5780 (N_5780,N_2878,N_3588);
or U5781 (N_5781,N_3123,N_3538);
or U5782 (N_5782,N_3412,N_2162);
nor U5783 (N_5783,N_2868,N_2908);
nor U5784 (N_5784,N_2880,N_2026);
or U5785 (N_5785,N_2793,N_3833);
nor U5786 (N_5786,N_3990,N_3031);
nand U5787 (N_5787,N_2908,N_3982);
or U5788 (N_5788,N_2411,N_2870);
nor U5789 (N_5789,N_2199,N_3783);
nor U5790 (N_5790,N_2175,N_3996);
and U5791 (N_5791,N_3850,N_2116);
or U5792 (N_5792,N_2061,N_3374);
and U5793 (N_5793,N_3123,N_2900);
or U5794 (N_5794,N_3593,N_2163);
nor U5795 (N_5795,N_2995,N_3258);
nor U5796 (N_5796,N_3350,N_2038);
or U5797 (N_5797,N_3310,N_3894);
and U5798 (N_5798,N_2611,N_3581);
nand U5799 (N_5799,N_3098,N_3046);
nand U5800 (N_5800,N_3849,N_2676);
and U5801 (N_5801,N_3260,N_2764);
nand U5802 (N_5802,N_2340,N_2596);
and U5803 (N_5803,N_2093,N_3799);
nand U5804 (N_5804,N_2391,N_2241);
or U5805 (N_5805,N_2045,N_2846);
and U5806 (N_5806,N_2441,N_3974);
and U5807 (N_5807,N_3256,N_3417);
nand U5808 (N_5808,N_3104,N_2558);
and U5809 (N_5809,N_3734,N_2957);
or U5810 (N_5810,N_3961,N_3805);
or U5811 (N_5811,N_2232,N_3887);
and U5812 (N_5812,N_2387,N_2004);
xnor U5813 (N_5813,N_3192,N_2287);
nor U5814 (N_5814,N_2555,N_2956);
nor U5815 (N_5815,N_2910,N_3477);
nand U5816 (N_5816,N_2710,N_3837);
or U5817 (N_5817,N_3504,N_3138);
or U5818 (N_5818,N_2376,N_2145);
or U5819 (N_5819,N_2836,N_3376);
or U5820 (N_5820,N_2861,N_2624);
nand U5821 (N_5821,N_2281,N_3024);
nand U5822 (N_5822,N_2288,N_3612);
or U5823 (N_5823,N_2887,N_2082);
nor U5824 (N_5824,N_3783,N_2623);
nand U5825 (N_5825,N_3469,N_2480);
or U5826 (N_5826,N_2413,N_2362);
nand U5827 (N_5827,N_2635,N_3244);
and U5828 (N_5828,N_2371,N_3417);
xor U5829 (N_5829,N_3450,N_2448);
nand U5830 (N_5830,N_2276,N_2625);
or U5831 (N_5831,N_2901,N_2778);
nor U5832 (N_5832,N_3803,N_3637);
nand U5833 (N_5833,N_2642,N_2051);
nand U5834 (N_5834,N_3084,N_3488);
xnor U5835 (N_5835,N_2554,N_2378);
or U5836 (N_5836,N_2412,N_2069);
xor U5837 (N_5837,N_3539,N_3760);
nor U5838 (N_5838,N_3839,N_3334);
or U5839 (N_5839,N_3646,N_3009);
or U5840 (N_5840,N_3228,N_3767);
nor U5841 (N_5841,N_3113,N_3496);
or U5842 (N_5842,N_3749,N_3534);
and U5843 (N_5843,N_2516,N_3277);
or U5844 (N_5844,N_3749,N_2744);
or U5845 (N_5845,N_3597,N_3583);
nor U5846 (N_5846,N_3660,N_3056);
nor U5847 (N_5847,N_2344,N_2512);
nor U5848 (N_5848,N_2157,N_2743);
or U5849 (N_5849,N_3985,N_2276);
nor U5850 (N_5850,N_3804,N_2811);
and U5851 (N_5851,N_3097,N_3089);
nor U5852 (N_5852,N_3275,N_2208);
nor U5853 (N_5853,N_3846,N_2487);
nor U5854 (N_5854,N_3991,N_3771);
or U5855 (N_5855,N_3111,N_2974);
and U5856 (N_5856,N_3191,N_2223);
or U5857 (N_5857,N_3286,N_3555);
and U5858 (N_5858,N_3396,N_3951);
nand U5859 (N_5859,N_3889,N_3720);
nor U5860 (N_5860,N_3805,N_2144);
nor U5861 (N_5861,N_2099,N_3580);
nor U5862 (N_5862,N_3606,N_3857);
nand U5863 (N_5863,N_2561,N_2961);
and U5864 (N_5864,N_3866,N_3387);
nand U5865 (N_5865,N_2523,N_2663);
and U5866 (N_5866,N_2478,N_2835);
and U5867 (N_5867,N_2248,N_3906);
nand U5868 (N_5868,N_2058,N_3045);
nor U5869 (N_5869,N_3351,N_3413);
nor U5870 (N_5870,N_2593,N_2479);
and U5871 (N_5871,N_2414,N_3722);
or U5872 (N_5872,N_3421,N_3863);
and U5873 (N_5873,N_2735,N_2907);
nand U5874 (N_5874,N_2130,N_3644);
nand U5875 (N_5875,N_3720,N_3428);
or U5876 (N_5876,N_3501,N_3850);
nand U5877 (N_5877,N_3534,N_3195);
and U5878 (N_5878,N_3388,N_3731);
nor U5879 (N_5879,N_2698,N_3319);
and U5880 (N_5880,N_2302,N_2038);
xnor U5881 (N_5881,N_3171,N_3317);
nand U5882 (N_5882,N_3099,N_3855);
xnor U5883 (N_5883,N_3197,N_2922);
nand U5884 (N_5884,N_3397,N_3733);
or U5885 (N_5885,N_2563,N_3836);
nor U5886 (N_5886,N_2239,N_2699);
nor U5887 (N_5887,N_2257,N_3659);
nand U5888 (N_5888,N_2852,N_2638);
or U5889 (N_5889,N_3409,N_2639);
nand U5890 (N_5890,N_3658,N_2342);
xor U5891 (N_5891,N_2370,N_2363);
nand U5892 (N_5892,N_3034,N_3149);
nand U5893 (N_5893,N_2347,N_3322);
xnor U5894 (N_5894,N_2647,N_3154);
or U5895 (N_5895,N_2899,N_2186);
and U5896 (N_5896,N_2625,N_3543);
or U5897 (N_5897,N_2099,N_3325);
or U5898 (N_5898,N_3951,N_3847);
or U5899 (N_5899,N_2232,N_2030);
nor U5900 (N_5900,N_3388,N_2316);
nor U5901 (N_5901,N_2377,N_2790);
xnor U5902 (N_5902,N_3845,N_3999);
nand U5903 (N_5903,N_3445,N_3301);
nand U5904 (N_5904,N_3601,N_3516);
or U5905 (N_5905,N_2969,N_2126);
xnor U5906 (N_5906,N_3858,N_2117);
or U5907 (N_5907,N_3686,N_3695);
nand U5908 (N_5908,N_3187,N_3341);
or U5909 (N_5909,N_3599,N_2846);
or U5910 (N_5910,N_3114,N_2939);
nand U5911 (N_5911,N_2340,N_2761);
and U5912 (N_5912,N_3724,N_3367);
nor U5913 (N_5913,N_2471,N_3213);
nor U5914 (N_5914,N_2111,N_3513);
or U5915 (N_5915,N_3574,N_3561);
and U5916 (N_5916,N_3257,N_3628);
or U5917 (N_5917,N_2181,N_3283);
nand U5918 (N_5918,N_3239,N_3937);
nand U5919 (N_5919,N_3110,N_3492);
nand U5920 (N_5920,N_2077,N_3710);
and U5921 (N_5921,N_3960,N_3329);
or U5922 (N_5922,N_2576,N_3328);
and U5923 (N_5923,N_3729,N_2157);
or U5924 (N_5924,N_3946,N_3185);
nand U5925 (N_5925,N_3926,N_2714);
nand U5926 (N_5926,N_3582,N_3010);
nand U5927 (N_5927,N_2365,N_2835);
or U5928 (N_5928,N_2303,N_3111);
nor U5929 (N_5929,N_2504,N_3449);
xor U5930 (N_5930,N_2183,N_3789);
or U5931 (N_5931,N_3361,N_3664);
and U5932 (N_5932,N_2533,N_3693);
and U5933 (N_5933,N_3361,N_3327);
nor U5934 (N_5934,N_3545,N_3516);
and U5935 (N_5935,N_2818,N_2662);
xor U5936 (N_5936,N_3931,N_2854);
nand U5937 (N_5937,N_3738,N_2303);
or U5938 (N_5938,N_2776,N_2556);
nand U5939 (N_5939,N_3832,N_2190);
or U5940 (N_5940,N_2109,N_3607);
nand U5941 (N_5941,N_3442,N_2188);
or U5942 (N_5942,N_3676,N_3944);
or U5943 (N_5943,N_2291,N_2868);
nor U5944 (N_5944,N_3494,N_2227);
or U5945 (N_5945,N_2724,N_3026);
or U5946 (N_5946,N_3662,N_2582);
or U5947 (N_5947,N_3307,N_2805);
nand U5948 (N_5948,N_3562,N_2688);
nand U5949 (N_5949,N_3722,N_3675);
nor U5950 (N_5950,N_3707,N_3695);
nand U5951 (N_5951,N_3502,N_3938);
nor U5952 (N_5952,N_2603,N_2997);
or U5953 (N_5953,N_2748,N_3354);
and U5954 (N_5954,N_2000,N_2901);
xnor U5955 (N_5955,N_2056,N_3833);
and U5956 (N_5956,N_3956,N_2619);
or U5957 (N_5957,N_2719,N_3319);
or U5958 (N_5958,N_2014,N_2921);
or U5959 (N_5959,N_3587,N_3416);
and U5960 (N_5960,N_2014,N_3447);
nand U5961 (N_5961,N_3137,N_3765);
nor U5962 (N_5962,N_3253,N_2513);
nand U5963 (N_5963,N_2573,N_3327);
nor U5964 (N_5964,N_2180,N_2382);
nor U5965 (N_5965,N_2417,N_2662);
and U5966 (N_5966,N_3563,N_3157);
nor U5967 (N_5967,N_3724,N_3054);
and U5968 (N_5968,N_3318,N_2743);
nand U5969 (N_5969,N_2475,N_2764);
or U5970 (N_5970,N_2630,N_2647);
nand U5971 (N_5971,N_3820,N_2153);
or U5972 (N_5972,N_3569,N_2731);
nor U5973 (N_5973,N_3223,N_2049);
or U5974 (N_5974,N_2293,N_2523);
or U5975 (N_5975,N_3917,N_3529);
or U5976 (N_5976,N_3464,N_2388);
xnor U5977 (N_5977,N_3025,N_2486);
or U5978 (N_5978,N_3127,N_2018);
and U5979 (N_5979,N_3584,N_2782);
nor U5980 (N_5980,N_2031,N_3982);
nor U5981 (N_5981,N_2392,N_2356);
or U5982 (N_5982,N_3037,N_2716);
nand U5983 (N_5983,N_3417,N_2052);
nor U5984 (N_5984,N_2183,N_2131);
xor U5985 (N_5985,N_3933,N_2206);
or U5986 (N_5986,N_3902,N_2945);
nand U5987 (N_5987,N_3787,N_2628);
nand U5988 (N_5988,N_3703,N_2882);
and U5989 (N_5989,N_2900,N_2627);
and U5990 (N_5990,N_2425,N_2324);
nand U5991 (N_5991,N_3388,N_3704);
and U5992 (N_5992,N_3230,N_3582);
and U5993 (N_5993,N_2071,N_2682);
nand U5994 (N_5994,N_3041,N_2178);
nand U5995 (N_5995,N_3488,N_3990);
nor U5996 (N_5996,N_3923,N_2410);
and U5997 (N_5997,N_2492,N_2337);
and U5998 (N_5998,N_2309,N_3531);
or U5999 (N_5999,N_3271,N_3167);
and U6000 (N_6000,N_4549,N_5332);
xor U6001 (N_6001,N_5528,N_5375);
and U6002 (N_6002,N_4666,N_5762);
or U6003 (N_6003,N_5751,N_5144);
nor U6004 (N_6004,N_5766,N_4216);
or U6005 (N_6005,N_5062,N_4951);
nand U6006 (N_6006,N_4582,N_4046);
nor U6007 (N_6007,N_5094,N_5594);
nand U6008 (N_6008,N_5341,N_5072);
nor U6009 (N_6009,N_5151,N_4130);
nor U6010 (N_6010,N_5630,N_5148);
xor U6011 (N_6011,N_5370,N_5146);
nor U6012 (N_6012,N_5791,N_5291);
and U6013 (N_6013,N_5217,N_4025);
or U6014 (N_6014,N_4357,N_5647);
nor U6015 (N_6015,N_5477,N_5673);
and U6016 (N_6016,N_5920,N_4113);
nand U6017 (N_6017,N_5404,N_5134);
xor U6018 (N_6018,N_4195,N_5018);
nand U6019 (N_6019,N_5118,N_4203);
or U6020 (N_6020,N_5328,N_5206);
or U6021 (N_6021,N_4230,N_5395);
or U6022 (N_6022,N_5973,N_4299);
nor U6023 (N_6023,N_4068,N_4442);
and U6024 (N_6024,N_4161,N_5908);
nand U6025 (N_6025,N_5798,N_4995);
nor U6026 (N_6026,N_5967,N_5150);
nand U6027 (N_6027,N_5759,N_4348);
or U6028 (N_6028,N_4853,N_4172);
and U6029 (N_6029,N_5023,N_4763);
or U6030 (N_6030,N_4278,N_4303);
nand U6031 (N_6031,N_5255,N_5748);
nor U6032 (N_6032,N_4087,N_5447);
nand U6033 (N_6033,N_4286,N_4662);
and U6034 (N_6034,N_5744,N_4351);
nand U6035 (N_6035,N_5989,N_5385);
and U6036 (N_6036,N_5536,N_4788);
xor U6037 (N_6037,N_5911,N_5689);
or U6038 (N_6038,N_5881,N_5698);
nor U6039 (N_6039,N_5520,N_5527);
and U6040 (N_6040,N_4564,N_5548);
and U6041 (N_6041,N_4518,N_5783);
or U6042 (N_6042,N_4345,N_4772);
or U6043 (N_6043,N_4449,N_5020);
and U6044 (N_6044,N_5015,N_4755);
and U6045 (N_6045,N_5164,N_5840);
xor U6046 (N_6046,N_5606,N_5602);
nand U6047 (N_6047,N_4801,N_4370);
nor U6048 (N_6048,N_4577,N_4277);
nand U6049 (N_6049,N_5931,N_5515);
nor U6050 (N_6050,N_5879,N_5032);
nand U6051 (N_6051,N_4349,N_5016);
or U6052 (N_6052,N_5357,N_5670);
nand U6053 (N_6053,N_5243,N_5098);
xor U6054 (N_6054,N_4058,N_5126);
or U6055 (N_6055,N_4287,N_4496);
or U6056 (N_6056,N_5279,N_4857);
xor U6057 (N_6057,N_4960,N_4222);
nand U6058 (N_6058,N_4674,N_4615);
nand U6059 (N_6059,N_4617,N_4503);
and U6060 (N_6060,N_4280,N_5320);
or U6061 (N_6061,N_5232,N_4010);
and U6062 (N_6062,N_4616,N_5066);
and U6063 (N_6063,N_5981,N_5403);
nor U6064 (N_6064,N_4391,N_5999);
nor U6065 (N_6065,N_4234,N_4892);
and U6066 (N_6066,N_4475,N_5728);
xnor U6067 (N_6067,N_5779,N_5005);
or U6068 (N_6068,N_5516,N_4245);
nand U6069 (N_6069,N_4194,N_5982);
nor U6070 (N_6070,N_5607,N_5764);
or U6071 (N_6071,N_4365,N_4780);
or U6072 (N_6072,N_4693,N_5768);
or U6073 (N_6073,N_5180,N_5252);
and U6074 (N_6074,N_4078,N_4974);
or U6075 (N_6075,N_4423,N_5773);
xor U6076 (N_6076,N_4739,N_4556);
and U6077 (N_6077,N_4399,N_4446);
nor U6078 (N_6078,N_5522,N_5771);
nor U6079 (N_6079,N_5414,N_5794);
nor U6080 (N_6080,N_4142,N_4304);
nor U6081 (N_6081,N_5889,N_5551);
and U6082 (N_6082,N_5581,N_4789);
and U6083 (N_6083,N_4288,N_5537);
and U6084 (N_6084,N_4879,N_5081);
nor U6085 (N_6085,N_5137,N_5487);
xnor U6086 (N_6086,N_5242,N_4191);
nand U6087 (N_6087,N_5869,N_5902);
and U6088 (N_6088,N_5208,N_4698);
nor U6089 (N_6089,N_4779,N_5872);
nand U6090 (N_6090,N_5886,N_4192);
nand U6091 (N_6091,N_5884,N_5381);
or U6092 (N_6092,N_4206,N_4353);
nand U6093 (N_6093,N_5914,N_4877);
nor U6094 (N_6094,N_5249,N_4988);
and U6095 (N_6095,N_5742,N_4089);
or U6096 (N_6096,N_5969,N_4590);
nor U6097 (N_6097,N_4724,N_5940);
nor U6098 (N_6098,N_4800,N_5099);
or U6099 (N_6099,N_5874,N_4930);
or U6100 (N_6100,N_4843,N_4606);
nor U6101 (N_6101,N_4175,N_4457);
nand U6102 (N_6102,N_5805,N_4066);
or U6103 (N_6103,N_5984,N_4906);
nand U6104 (N_6104,N_5730,N_5333);
nand U6105 (N_6105,N_4608,N_4229);
xor U6106 (N_6106,N_4821,N_4744);
nor U6107 (N_6107,N_5371,N_5503);
nor U6108 (N_6108,N_5786,N_5177);
and U6109 (N_6109,N_4980,N_5300);
nand U6110 (N_6110,N_5435,N_5642);
or U6111 (N_6111,N_5226,N_5068);
nor U6112 (N_6112,N_4104,N_4659);
and U6113 (N_6113,N_4186,N_5121);
nand U6114 (N_6114,N_5864,N_5039);
nand U6115 (N_6115,N_4088,N_5873);
or U6116 (N_6116,N_4753,N_5233);
nand U6117 (N_6117,N_4181,N_5084);
or U6118 (N_6118,N_4713,N_4574);
nor U6119 (N_6119,N_4211,N_4425);
nand U6120 (N_6120,N_5396,N_4897);
nor U6121 (N_6121,N_4734,N_5464);
nand U6122 (N_6122,N_4591,N_5525);
nand U6123 (N_6123,N_5947,N_4364);
xor U6124 (N_6124,N_4413,N_5212);
nand U6125 (N_6125,N_5076,N_4664);
xnor U6126 (N_6126,N_4411,N_4661);
nor U6127 (N_6127,N_5498,N_5966);
nand U6128 (N_6128,N_5650,N_5221);
and U6129 (N_6129,N_4035,N_5380);
nor U6130 (N_6130,N_4942,N_4377);
and U6131 (N_6131,N_4009,N_4650);
xnor U6132 (N_6132,N_5008,N_4014);
or U6133 (N_6133,N_5053,N_4132);
nor U6134 (N_6134,N_4905,N_5376);
or U6135 (N_6135,N_4311,N_4831);
nand U6136 (N_6136,N_4949,N_4363);
nand U6137 (N_6137,N_5045,N_5885);
nand U6138 (N_6138,N_4008,N_4371);
nand U6139 (N_6139,N_5505,N_5219);
nor U6140 (N_6140,N_4137,N_5882);
nand U6141 (N_6141,N_5955,N_5912);
and U6142 (N_6142,N_5448,N_5968);
xor U6143 (N_6143,N_4251,N_4221);
and U6144 (N_6144,N_4568,N_5796);
nor U6145 (N_6145,N_5059,N_4407);
and U6146 (N_6146,N_4197,N_5750);
nand U6147 (N_6147,N_5553,N_4252);
nand U6148 (N_6148,N_5792,N_5655);
or U6149 (N_6149,N_5245,N_4914);
and U6150 (N_6150,N_4957,N_4307);
or U6151 (N_6151,N_4787,N_4640);
and U6152 (N_6152,N_5535,N_4471);
nor U6153 (N_6153,N_4757,N_5990);
xor U6154 (N_6154,N_4395,N_5962);
nor U6155 (N_6155,N_5286,N_5119);
nand U6156 (N_6156,N_4696,N_4400);
xor U6157 (N_6157,N_4302,N_4096);
nand U6158 (N_6158,N_4219,N_4485);
xnor U6159 (N_6159,N_5697,N_5293);
or U6160 (N_6160,N_5677,N_5679);
nor U6161 (N_6161,N_5163,N_5531);
or U6162 (N_6162,N_5348,N_4810);
or U6163 (N_6163,N_4099,N_5740);
nor U6164 (N_6164,N_5866,N_5408);
and U6165 (N_6165,N_4908,N_5756);
xnor U6166 (N_6166,N_5063,N_5133);
and U6167 (N_6167,N_4547,N_5671);
and U6168 (N_6168,N_4158,N_4467);
nand U6169 (N_6169,N_5721,N_4785);
and U6170 (N_6170,N_4947,N_4510);
nor U6171 (N_6171,N_4835,N_5596);
nand U6172 (N_6172,N_5257,N_4016);
and U6173 (N_6173,N_5574,N_5311);
and U6174 (N_6174,N_5054,N_4599);
nand U6175 (N_6175,N_5316,N_5350);
and U6176 (N_6176,N_4361,N_5430);
or U6177 (N_6177,N_5913,N_4885);
nand U6178 (N_6178,N_4682,N_4913);
nor U6179 (N_6179,N_5563,N_4204);
nor U6180 (N_6180,N_4473,N_5561);
nand U6181 (N_6181,N_4215,N_4898);
nor U6182 (N_6182,N_5135,N_4783);
nand U6183 (N_6183,N_4013,N_4409);
and U6184 (N_6184,N_5024,N_4597);
and U6185 (N_6185,N_4968,N_4404);
xor U6186 (N_6186,N_5562,N_5521);
and U6187 (N_6187,N_5754,N_5711);
nor U6188 (N_6188,N_5860,N_5616);
nor U6189 (N_6189,N_5850,N_5767);
xor U6190 (N_6190,N_4891,N_5268);
nand U6191 (N_6191,N_4490,N_5841);
xnor U6192 (N_6192,N_5317,N_5471);
and U6193 (N_6193,N_5075,N_4105);
nor U6194 (N_6194,N_4474,N_5285);
xor U6195 (N_6195,N_5335,N_4658);
and U6196 (N_6196,N_4808,N_5851);
nand U6197 (N_6197,N_5407,N_5322);
nor U6198 (N_6198,N_5154,N_4502);
or U6199 (N_6199,N_5241,N_4073);
or U6200 (N_6200,N_4188,N_4396);
and U6201 (N_6201,N_5368,N_5567);
nand U6202 (N_6202,N_4356,N_5305);
and U6203 (N_6203,N_5200,N_5389);
nor U6204 (N_6204,N_5443,N_4836);
nand U6205 (N_6205,N_4094,N_5390);
nand U6206 (N_6206,N_4963,N_4289);
nor U6207 (N_6207,N_4943,N_4781);
nand U6208 (N_6208,N_4180,N_5188);
and U6209 (N_6209,N_4902,N_4306);
or U6210 (N_6210,N_4149,N_4634);
or U6211 (N_6211,N_5785,N_5486);
or U6212 (N_6212,N_4402,N_5169);
nor U6213 (N_6213,N_4961,N_5720);
nand U6214 (N_6214,N_4707,N_5096);
nor U6215 (N_6215,N_5472,N_4687);
or U6216 (N_6216,N_5343,N_4032);
and U6217 (N_6217,N_4569,N_4583);
xor U6218 (N_6218,N_4019,N_4776);
nand U6219 (N_6219,N_5559,N_5399);
nor U6220 (N_6220,N_5852,N_5543);
or U6221 (N_6221,N_4486,N_5699);
or U6222 (N_6222,N_5455,N_4579);
and U6223 (N_6223,N_4129,N_4292);
nor U6224 (N_6224,N_5410,N_5131);
nand U6225 (N_6225,N_5079,N_5669);
nor U6226 (N_6226,N_5497,N_4387);
nor U6227 (N_6227,N_5833,N_4163);
xnor U6228 (N_6228,N_5092,N_5731);
and U6229 (N_6229,N_5778,N_4055);
or U6230 (N_6230,N_5945,N_5877);
nor U6231 (N_6231,N_5592,N_5540);
and U6232 (N_6232,N_4170,N_4271);
or U6233 (N_6233,N_5712,N_5411);
nand U6234 (N_6234,N_4895,N_5000);
nor U6235 (N_6235,N_5366,N_4508);
or U6236 (N_6236,N_5113,N_4421);
nand U6237 (N_6237,N_4624,N_5713);
nor U6238 (N_6238,N_5340,N_5351);
and U6239 (N_6239,N_4489,N_4081);
nand U6240 (N_6240,N_4466,N_4765);
or U6241 (N_6241,N_4714,N_5808);
and U6242 (N_6242,N_4354,N_5964);
or U6243 (N_6243,N_5500,N_4838);
or U6244 (N_6244,N_5468,N_4074);
nand U6245 (N_6245,N_4994,N_4944);
and U6246 (N_6246,N_4101,N_5585);
or U6247 (N_6247,N_4575,N_5557);
nand U6248 (N_6248,N_4685,N_5437);
nor U6249 (N_6249,N_5256,N_5619);
or U6250 (N_6250,N_5275,N_4869);
xnor U6251 (N_6251,N_5310,N_5544);
xnor U6252 (N_6252,N_5844,N_4505);
or U6253 (N_6253,N_4177,N_4282);
xor U6254 (N_6254,N_4341,N_5198);
nor U6255 (N_6255,N_4705,N_4342);
or U6256 (N_6256,N_5262,N_4362);
and U6257 (N_6257,N_4632,N_4381);
nor U6258 (N_6258,N_5014,N_5861);
and U6259 (N_6259,N_4822,N_4332);
nor U6260 (N_6260,N_5649,N_5662);
nor U6261 (N_6261,N_5047,N_5265);
or U6262 (N_6262,N_5970,N_4148);
nand U6263 (N_6263,N_5306,N_5122);
or U6264 (N_6264,N_4437,N_4817);
nor U6265 (N_6265,N_5769,N_5052);
xnor U6266 (N_6266,N_4657,N_5895);
nand U6267 (N_6267,N_4500,N_5664);
nand U6268 (N_6268,N_5838,N_4270);
or U6269 (N_6269,N_5462,N_4525);
xor U6270 (N_6270,N_4305,N_5700);
and U6271 (N_6271,N_4325,N_4513);
and U6272 (N_6272,N_4483,N_4903);
and U6273 (N_6273,N_5996,N_5620);
nand U6274 (N_6274,N_5452,N_4213);
or U6275 (N_6275,N_4719,N_4022);
and U6276 (N_6276,N_5813,N_4571);
nor U6277 (N_6277,N_4596,N_4884);
or U6278 (N_6278,N_4570,N_4935);
nand U6279 (N_6279,N_5202,N_5733);
xnor U6280 (N_6280,N_4006,N_4858);
nor U6281 (N_6281,N_5314,N_5761);
xnor U6282 (N_6282,N_5723,N_5070);
nand U6283 (N_6283,N_4764,N_5919);
or U6284 (N_6284,N_5104,N_5901);
and U6285 (N_6285,N_5082,N_5490);
nand U6286 (N_6286,N_4833,N_4840);
nand U6287 (N_6287,N_5871,N_4079);
nand U6288 (N_6288,N_4339,N_4346);
xor U6289 (N_6289,N_4774,N_4359);
and U6290 (N_6290,N_5218,N_4070);
nor U6291 (N_6291,N_4152,N_5278);
nor U6292 (N_6292,N_5201,N_5444);
nor U6293 (N_6293,N_4793,N_4048);
and U6294 (N_6294,N_4390,N_5240);
nand U6295 (N_6295,N_4488,N_5176);
nor U6296 (N_6296,N_4253,N_5203);
and U6297 (N_6297,N_4071,N_5818);
and U6298 (N_6298,N_4126,N_4600);
or U6299 (N_6299,N_5858,N_4217);
nor U6300 (N_6300,N_5821,N_4406);
nor U6301 (N_6301,N_5331,N_5934);
and U6302 (N_6302,N_5654,N_5809);
and U6303 (N_6303,N_4460,N_5405);
nor U6304 (N_6304,N_4504,N_4123);
nor U6305 (N_6305,N_4082,N_4924);
or U6306 (N_6306,N_5010,N_5524);
or U6307 (N_6307,N_5915,N_4536);
or U6308 (N_6308,N_4379,N_4455);
nand U6309 (N_6309,N_5565,N_4737);
nor U6310 (N_6310,N_4829,N_4720);
xor U6311 (N_6311,N_4690,N_4695);
and U6312 (N_6312,N_5264,N_4124);
and U6313 (N_6313,N_4852,N_5356);
nor U6314 (N_6314,N_4040,N_4845);
xor U6315 (N_6315,N_5753,N_4526);
or U6316 (N_6316,N_5211,N_4977);
nor U6317 (N_6317,N_4621,N_4205);
nor U6318 (N_6318,N_4224,N_5186);
nor U6319 (N_6319,N_4804,N_5601);
or U6320 (N_6320,N_4921,N_5246);
nor U6321 (N_6321,N_5458,N_4694);
or U6322 (N_6322,N_4313,N_4760);
nand U6323 (N_6323,N_5037,N_4711);
nor U6324 (N_6324,N_5780,N_4433);
nor U6325 (N_6325,N_5634,N_4340);
or U6326 (N_6326,N_5738,N_4609);
nand U6327 (N_6327,N_5397,N_4702);
nand U6328 (N_6328,N_5077,N_4972);
nand U6329 (N_6329,N_4005,N_5267);
nand U6330 (N_6330,N_4060,N_5022);
or U6331 (N_6331,N_5493,N_4108);
or U6332 (N_6332,N_4168,N_4378);
and U6333 (N_6333,N_4514,N_4915);
or U6334 (N_6334,N_5292,N_5334);
nand U6335 (N_6335,N_4448,N_4594);
and U6336 (N_6336,N_5932,N_4716);
or U6337 (N_6337,N_4939,N_4867);
nand U6338 (N_6338,N_5423,N_5453);
and U6339 (N_6339,N_5632,N_4328);
nand U6340 (N_6340,N_4710,N_4360);
nand U6341 (N_6341,N_5695,N_5238);
and U6342 (N_6342,N_4668,N_4761);
nor U6343 (N_6343,N_4811,N_4777);
nor U6344 (N_6344,N_5853,N_4045);
nand U6345 (N_6345,N_4098,N_5485);
xor U6346 (N_6346,N_5604,N_5299);
or U6347 (N_6347,N_5701,N_4166);
nand U6348 (N_6348,N_4978,N_4532);
nor U6349 (N_6349,N_5875,N_4160);
nor U6350 (N_6350,N_4210,N_4086);
xnor U6351 (N_6351,N_4290,N_5442);
nand U6352 (N_6352,N_4966,N_5019);
nand U6353 (N_6353,N_5504,N_5986);
or U6354 (N_6354,N_5459,N_5237);
xnor U6355 (N_6355,N_4268,N_4117);
nand U6356 (N_6356,N_4746,N_4157);
and U6357 (N_6357,N_5755,N_4647);
nor U6358 (N_6358,N_5213,N_5890);
nor U6359 (N_6359,N_4049,N_4122);
nor U6360 (N_6360,N_5182,N_4015);
nand U6361 (N_6361,N_4626,N_4103);
nand U6362 (N_6362,N_4092,N_4064);
and U6363 (N_6363,N_4805,N_5743);
nand U6364 (N_6364,N_4438,N_4033);
nor U6365 (N_6365,N_4509,N_5752);
nand U6366 (N_6366,N_5646,N_5575);
nand U6367 (N_6367,N_5228,N_5434);
nand U6368 (N_6368,N_4444,N_4434);
nand U6369 (N_6369,N_4775,N_4655);
or U6370 (N_6370,N_5804,N_5749);
nand U6371 (N_6371,N_4227,N_4652);
and U6372 (N_6372,N_5897,N_5958);
and U6373 (N_6373,N_5330,N_4100);
nand U6374 (N_6374,N_4860,N_4826);
nor U6375 (N_6375,N_5765,N_5888);
nor U6376 (N_6376,N_4083,N_4736);
or U6377 (N_6377,N_4771,N_5726);
or U6378 (N_6378,N_5847,N_4233);
and U6379 (N_6379,N_5906,N_4263);
xnor U6380 (N_6380,N_5481,N_4246);
or U6381 (N_6381,N_4000,N_4334);
and U6382 (N_6382,N_4128,N_5400);
nor U6383 (N_6383,N_4431,N_4680);
or U6384 (N_6384,N_5660,N_5367);
and U6385 (N_6385,N_4336,N_5489);
xnor U6386 (N_6386,N_4792,N_5878);
nand U6387 (N_6387,N_4611,N_4709);
or U6388 (N_6388,N_4533,N_4552);
nor U6389 (N_6389,N_5355,N_5980);
nand U6390 (N_6390,N_5529,N_5026);
nor U6391 (N_6391,N_5974,N_5484);
nor U6392 (N_6392,N_4164,N_4796);
and U6393 (N_6393,N_5272,N_4412);
nor U6394 (N_6394,N_5048,N_4589);
xnor U6395 (N_6395,N_4839,N_5976);
xor U6396 (N_6396,N_5261,N_5644);
xnor U6397 (N_6397,N_5067,N_4723);
nor U6398 (N_6398,N_5640,N_5501);
nor U6399 (N_6399,N_5523,N_4844);
nand U6400 (N_6400,N_4894,N_4201);
nand U6401 (N_6401,N_4454,N_5862);
or U6402 (N_6402,N_4459,N_4855);
nand U6403 (N_6403,N_5801,N_5591);
nor U6404 (N_6404,N_4481,N_5009);
nor U6405 (N_6405,N_4135,N_4522);
nor U6406 (N_6406,N_4748,N_4519);
nand U6407 (N_6407,N_4856,N_5588);
and U6408 (N_6408,N_4688,N_5116);
and U6409 (N_6409,N_4144,N_4329);
and U6410 (N_6410,N_5132,N_4971);
nand U6411 (N_6411,N_5635,N_4768);
and U6412 (N_6412,N_5483,N_5933);
and U6413 (N_6413,N_4118,N_5717);
nor U6414 (N_6414,N_5495,N_5419);
nand U6415 (N_6415,N_5454,N_4663);
nor U6416 (N_6416,N_5868,N_5690);
and U6417 (N_6417,N_5883,N_5938);
xnor U6418 (N_6418,N_4063,N_4469);
and U6419 (N_6419,N_4642,N_4029);
nor U6420 (N_6420,N_4382,N_4323);
or U6421 (N_6421,N_4560,N_5952);
and U6422 (N_6422,N_4487,N_5854);
or U6423 (N_6423,N_4740,N_5876);
or U6424 (N_6424,N_4926,N_5281);
and U6425 (N_6425,N_4964,N_5187);
nand U6426 (N_6426,N_5432,N_5149);
nand U6427 (N_6427,N_4706,N_5573);
and U6428 (N_6428,N_5347,N_5600);
or U6429 (N_6429,N_5470,N_5450);
xnor U6430 (N_6430,N_4628,N_4607);
or U6431 (N_6431,N_5109,N_4883);
nand U6432 (N_6432,N_4479,N_4766);
nor U6433 (N_6433,N_4482,N_5001);
or U6434 (N_6434,N_4563,N_5824);
nand U6435 (N_6435,N_4102,N_4044);
nor U6436 (N_6436,N_5044,N_5128);
xor U6437 (N_6437,N_4478,N_5511);
nand U6438 (N_6438,N_4881,N_4633);
or U6439 (N_6439,N_4176,N_4043);
or U6440 (N_6440,N_4531,N_4432);
and U6441 (N_6441,N_5788,N_4672);
or U6442 (N_6442,N_4090,N_4630);
or U6443 (N_6443,N_5849,N_4925);
and U6444 (N_6444,N_4981,N_5645);
or U6445 (N_6445,N_5398,N_5703);
and U6446 (N_6446,N_5239,N_4610);
xor U6447 (N_6447,N_5051,N_5739);
nand U6448 (N_6448,N_4538,N_5142);
nand U6449 (N_6449,N_4795,N_4653);
nor U6450 (N_6450,N_4627,N_4384);
xnor U6451 (N_6451,N_4794,N_5153);
nor U6452 (N_6452,N_4051,N_5280);
and U6453 (N_6453,N_5668,N_5758);
xnor U6454 (N_6454,N_5843,N_5112);
or U6455 (N_6455,N_4612,N_5929);
nor U6456 (N_6456,N_5139,N_5401);
and U6457 (N_6457,N_5820,N_5225);
or U6458 (N_6458,N_4366,N_5492);
nand U6459 (N_6459,N_5339,N_4133);
nand U6460 (N_6460,N_5080,N_5378);
xnor U6461 (N_6461,N_4002,N_4959);
xnor U6462 (N_6462,N_5569,N_4799);
and U6463 (N_6463,N_5629,N_4992);
nor U6464 (N_6464,N_4576,N_5095);
nor U6465 (N_6465,N_4298,N_5383);
xnor U6466 (N_6466,N_5171,N_4871);
and U6467 (N_6467,N_4550,N_4375);
or U6468 (N_6468,N_4383,N_5971);
nor U6469 (N_6469,N_5103,N_4093);
nand U6470 (N_6470,N_4054,N_5597);
and U6471 (N_6471,N_4061,N_4922);
nand U6472 (N_6472,N_4131,N_5174);
and U6473 (N_6473,N_5409,N_4401);
nand U6474 (N_6474,N_5309,N_5181);
nor U6475 (N_6475,N_5922,N_4828);
nor U6476 (N_6476,N_4374,N_4791);
xor U6477 (N_6477,N_5259,N_4430);
xnor U6478 (N_6478,N_4882,N_5956);
and U6479 (N_6479,N_5757,N_5760);
nand U6480 (N_6480,N_5580,N_5294);
and U6481 (N_6481,N_5611,N_4248);
nor U6482 (N_6482,N_4067,N_4372);
nor U6483 (N_6483,N_4984,N_5506);
or U6484 (N_6484,N_4837,N_4851);
and U6485 (N_6485,N_4759,N_5704);
and U6486 (N_6486,N_4279,N_4376);
and U6487 (N_6487,N_4733,N_5360);
nand U6488 (N_6488,N_5961,N_4782);
nand U6489 (N_6489,N_4986,N_5438);
or U6490 (N_6490,N_5512,N_5715);
or U6491 (N_6491,N_4725,N_5110);
and U6492 (N_6492,N_5692,N_4141);
and U6493 (N_6493,N_4675,N_4001);
nor U6494 (N_6494,N_4330,N_4284);
nand U6495 (N_6495,N_5905,N_5071);
or U6496 (N_6496,N_4050,N_4335);
nand U6497 (N_6497,N_5336,N_4445);
nor U6498 (N_6498,N_4187,N_4807);
xor U6499 (N_6499,N_4031,N_4324);
nand U6500 (N_6500,N_4199,N_4727);
xor U6501 (N_6501,N_4752,N_5101);
or U6502 (N_6502,N_5942,N_5165);
and U6503 (N_6503,N_5160,N_4196);
and U6504 (N_6504,N_5572,N_5910);
or U6505 (N_6505,N_4007,N_5276);
nand U6506 (N_6506,N_4708,N_5158);
and U6507 (N_6507,N_4742,N_5994);
nor U6508 (N_6508,N_4169,N_4991);
and U6509 (N_6509,N_4861,N_4692);
xor U6510 (N_6510,N_4834,N_4750);
and U6511 (N_6511,N_4940,N_5582);
and U6512 (N_6512,N_5021,N_5382);
and U6513 (N_6513,N_5936,N_5946);
and U6514 (N_6514,N_5667,N_5993);
nand U6515 (N_6515,N_4173,N_5709);
or U6516 (N_6516,N_4786,N_5013);
and U6517 (N_6517,N_4717,N_5775);
nor U6518 (N_6518,N_5556,N_4472);
and U6519 (N_6519,N_5427,N_5318);
nand U6520 (N_6520,N_5266,N_5948);
xnor U6521 (N_6521,N_5289,N_5325);
and U6522 (N_6522,N_5327,N_5033);
nor U6523 (N_6523,N_5802,N_5125);
or U6524 (N_6524,N_5965,N_4393);
and U6525 (N_6525,N_4084,N_4639);
nand U6526 (N_6526,N_4558,N_5358);
nor U6527 (N_6527,N_5725,N_5896);
and U6528 (N_6528,N_5337,N_5473);
xnor U6529 (N_6529,N_4975,N_5064);
nor U6530 (N_6530,N_4258,N_5954);
nand U6531 (N_6531,N_4427,N_5352);
and U6532 (N_6532,N_5178,N_5819);
and U6533 (N_6533,N_5867,N_4424);
nand U6534 (N_6534,N_5248,N_4876);
nor U6535 (N_6535,N_5078,N_5782);
or U6536 (N_6536,N_4983,N_5735);
nor U6537 (N_6537,N_4405,N_4262);
nand U6538 (N_6538,N_4797,N_4300);
and U6539 (N_6539,N_4156,N_5787);
or U6540 (N_6540,N_5894,N_5959);
or U6541 (N_6541,N_5823,N_4352);
and U6542 (N_6542,N_5183,N_4138);
and U6543 (N_6543,N_5814,N_5927);
nor U6544 (N_6544,N_4017,N_5214);
nor U6545 (N_6545,N_5631,N_5426);
nor U6546 (N_6546,N_5859,N_4480);
nor U6547 (N_6547,N_4110,N_5394);
and U6548 (N_6548,N_5887,N_5034);
or U6549 (N_6549,N_4443,N_4223);
nand U6550 (N_6550,N_4397,N_4119);
nand U6551 (N_6551,N_4095,N_4866);
nand U6552 (N_6552,N_4498,N_4973);
or U6553 (N_6553,N_5857,N_4573);
nand U6554 (N_6554,N_5935,N_5518);
nor U6555 (N_6555,N_5517,N_5393);
nand U6556 (N_6556,N_4237,N_4602);
xor U6557 (N_6557,N_4751,N_4447);
nor U6558 (N_6558,N_4316,N_4967);
and U6559 (N_6559,N_5479,N_4499);
or U6560 (N_6560,N_5329,N_5231);
nor U6561 (N_6561,N_5377,N_5627);
nand U6562 (N_6562,N_5209,N_4107);
nor U6563 (N_6563,N_4976,N_5688);
nor U6564 (N_6564,N_4778,N_5192);
or U6565 (N_6565,N_5475,N_4419);
nand U6566 (N_6566,N_5807,N_5831);
nor U6567 (N_6567,N_4147,N_4641);
nand U6568 (N_6568,N_5577,N_5321);
or U6569 (N_6569,N_4398,N_4150);
or U6570 (N_6570,N_4758,N_5421);
or U6571 (N_6571,N_4996,N_5012);
and U6572 (N_6572,N_5369,N_4605);
xnor U6573 (N_6573,N_5530,N_4111);
nand U6574 (N_6574,N_5324,N_5258);
or U6575 (N_6575,N_4542,N_4465);
and U6576 (N_6576,N_4697,N_5196);
or U6577 (N_6577,N_4979,N_4997);
or U6578 (N_6578,N_4408,N_5166);
nor U6579 (N_6579,N_5770,N_5345);
xor U6580 (N_6580,N_4441,N_4179);
nand U6581 (N_6581,N_4145,N_4998);
nor U6582 (N_6582,N_4901,N_4403);
nand U6583 (N_6583,N_4644,N_4820);
and U6584 (N_6584,N_4272,N_5784);
or U6585 (N_6585,N_5595,N_4729);
nand U6586 (N_6586,N_5584,N_5793);
or U6587 (N_6587,N_4327,N_4458);
nand U6588 (N_6588,N_4613,N_5185);
and U6589 (N_6589,N_4011,N_5161);
nor U6590 (N_6590,N_4830,N_5608);
and U6591 (N_6591,N_5223,N_5917);
or U6592 (N_6592,N_5391,N_5763);
xnor U6593 (N_6593,N_5085,N_4970);
xnor U6594 (N_6594,N_5060,N_5613);
or U6595 (N_6595,N_5848,N_4343);
and U6596 (N_6596,N_4841,N_4721);
or U6597 (N_6597,N_5170,N_5776);
nor U6598 (N_6598,N_4699,N_4301);
or U6599 (N_6599,N_5983,N_5184);
and U6600 (N_6600,N_5041,N_4923);
or U6601 (N_6601,N_4159,N_4517);
nand U6602 (N_6602,N_4167,N_5465);
or U6603 (N_6603,N_4681,N_4076);
and U6604 (N_6604,N_5988,N_5845);
or U6605 (N_6605,N_5615,N_5598);
nor U6606 (N_6606,N_5702,N_5727);
nor U6607 (N_6607,N_5510,N_5552);
and U6608 (N_6608,N_5050,N_4309);
nor U6609 (N_6609,N_5810,N_5365);
xor U6610 (N_6610,N_4769,N_5089);
and U6611 (N_6611,N_4162,N_4056);
and U6612 (N_6612,N_5282,N_4242);
nand U6613 (N_6613,N_5904,N_5666);
and U6614 (N_6614,N_5508,N_4965);
and U6615 (N_6615,N_4394,N_5029);
or U6616 (N_6616,N_4809,N_4470);
and U6617 (N_6617,N_5846,N_4893);
or U6618 (N_6618,N_4917,N_4484);
nand U6619 (N_6619,N_5672,N_5466);
xnor U6620 (N_6620,N_5253,N_5539);
nand U6621 (N_6621,N_4516,N_5446);
or U6622 (N_6622,N_4386,N_4004);
or U6623 (N_6623,N_5195,N_5795);
and U6624 (N_6624,N_4257,N_4493);
nor U6625 (N_6625,N_4601,N_5296);
xor U6626 (N_6626,N_4151,N_5541);
nor U6627 (N_6627,N_5772,N_4651);
xor U6628 (N_6628,N_4027,N_4741);
and U6629 (N_6629,N_4034,N_5621);
and U6630 (N_6630,N_5681,N_4874);
and U6631 (N_6631,N_5056,N_5745);
or U6632 (N_6632,N_5560,N_5127);
and U6633 (N_6633,N_4859,N_4308);
and U6634 (N_6634,N_5460,N_5923);
nor U6635 (N_6635,N_4854,N_5729);
nor U6636 (N_6636,N_4476,N_5921);
or U6637 (N_6637,N_4665,N_5558);
or U6638 (N_6638,N_4320,N_5898);
nor U6639 (N_6639,N_4256,N_4910);
or U6640 (N_6640,N_4297,N_4291);
nand U6641 (N_6641,N_4932,N_4566);
nand U6642 (N_6642,N_4890,N_5207);
nor U6643 (N_6643,N_4109,N_4267);
or U6644 (N_6644,N_5930,N_5046);
and U6645 (N_6645,N_4261,N_5027);
xor U6646 (N_6646,N_5686,N_4784);
nand U6647 (N_6647,N_4812,N_5641);
and U6648 (N_6648,N_5254,N_4847);
and U6649 (N_6649,N_4062,N_4548);
nand U6650 (N_6650,N_4153,N_5985);
xnor U6651 (N_6651,N_5829,N_4461);
nand U6652 (N_6652,N_4945,N_5937);
xnor U6653 (N_6653,N_4134,N_5093);
and U6654 (N_6654,N_5741,N_5514);
and U6655 (N_6655,N_5083,N_5308);
or U6656 (N_6656,N_4738,N_5222);
or U6657 (N_6657,N_5162,N_4020);
xnor U6658 (N_6658,N_4887,N_5599);
or U6659 (N_6659,N_5637,N_4296);
nor U6660 (N_6660,N_4198,N_4728);
nand U6661 (N_6661,N_5230,N_5107);
and U6662 (N_6662,N_5618,N_4429);
and U6663 (N_6663,N_4244,N_4214);
and U6664 (N_6664,N_4190,N_4185);
or U6665 (N_6665,N_4919,N_4580);
or U6666 (N_6666,N_5073,N_5236);
or U6667 (N_6667,N_5361,N_4154);
and U6668 (N_6668,N_4036,N_4207);
or U6669 (N_6669,N_4825,N_4464);
and U6670 (N_6670,N_5880,N_5431);
nor U6671 (N_6671,N_4931,N_4410);
nor U6672 (N_6672,N_5576,N_5179);
and U6673 (N_6673,N_4456,N_5346);
or U6674 (N_6674,N_5412,N_4726);
nor U6675 (N_6675,N_5835,N_4614);
nor U6676 (N_6676,N_4420,N_5892);
nand U6677 (N_6677,N_5141,N_4933);
xor U6678 (N_6678,N_5992,N_5918);
nand U6679 (N_6679,N_5273,N_5747);
or U6680 (N_6680,N_4802,N_5502);
nor U6681 (N_6681,N_5461,N_4112);
xnor U6682 (N_6682,N_4275,N_5799);
nor U6683 (N_6683,N_5718,N_5172);
xnor U6684 (N_6684,N_5156,N_5338);
nor U6685 (N_6685,N_4544,N_4899);
nand U6686 (N_6686,N_5002,N_5656);
nor U6687 (N_6687,N_5433,N_5220);
and U6688 (N_6688,N_4041,N_5304);
xor U6689 (N_6689,N_4731,N_5925);
or U6690 (N_6690,N_5108,N_4028);
or U6691 (N_6691,N_4511,N_5250);
xor U6692 (N_6692,N_4684,N_5418);
and U6693 (N_6693,N_5826,N_4749);
and U6694 (N_6694,N_4264,N_5706);
xor U6695 (N_6695,N_4565,N_4848);
xnor U6696 (N_6696,N_4816,N_5863);
nor U6697 (N_6697,N_5145,N_5190);
and U6698 (N_6698,N_4232,N_4436);
nand U6699 (N_6699,N_5097,N_5714);
or U6700 (N_6700,N_4562,N_4491);
nand U6701 (N_6701,N_4468,N_4896);
nor U6702 (N_6702,N_5665,N_4656);
or U6703 (N_6703,N_4643,N_4247);
nor U6704 (N_6704,N_4072,N_4554);
and U6705 (N_6705,N_4868,N_4527);
xor U6706 (N_6706,N_4178,N_4555);
nand U6707 (N_6707,N_5189,N_4850);
nand U6708 (N_6708,N_5997,N_4136);
nand U6709 (N_6709,N_4355,N_5496);
xor U6710 (N_6710,N_4722,N_4414);
or U6711 (N_6711,N_5696,N_5509);
nor U6712 (N_6712,N_4281,N_5817);
nor U6713 (N_6713,N_5197,N_4226);
xor U6714 (N_6714,N_4417,N_4718);
or U6715 (N_6715,N_5017,N_4620);
and U6716 (N_6716,N_5903,N_5274);
nor U6717 (N_6717,N_5519,N_4603);
nand U6718 (N_6718,N_5724,N_4314);
nand U6719 (N_6719,N_4120,N_4052);
or U6720 (N_6720,N_4637,N_5057);
and U6721 (N_6721,N_5722,N_5251);
nor U6722 (N_6722,N_4018,N_5663);
or U6723 (N_6723,N_5106,N_5534);
xor U6724 (N_6724,N_4551,N_5694);
xnor U6725 (N_6725,N_4545,N_4515);
nor U6726 (N_6726,N_5006,N_5837);
xor U6727 (N_6727,N_5676,N_4106);
xnor U6728 (N_6728,N_5564,N_5031);
nand U6729 (N_6729,N_4561,N_4824);
nor U6730 (N_6730,N_4451,N_4174);
nor U6731 (N_6731,N_4938,N_4712);
nor U6732 (N_6732,N_5583,N_4543);
and U6733 (N_6733,N_4184,N_4115);
xor U6734 (N_6734,N_4059,N_5387);
or U6735 (N_6735,N_4790,N_5812);
nor U6736 (N_6736,N_5855,N_4982);
or U6737 (N_6737,N_5803,N_4598);
and U6738 (N_6738,N_4085,N_5359);
and U6739 (N_6739,N_5977,N_4559);
or U6740 (N_6740,N_5836,N_4704);
nor U6741 (N_6741,N_4380,N_4941);
or U6742 (N_6742,N_4671,N_4814);
nor U6743 (N_6743,N_4806,N_5205);
or U6744 (N_6744,N_5568,N_5307);
or U6745 (N_6745,N_5413,N_5229);
nor U6746 (N_6746,N_4987,N_4862);
nand U6747 (N_6747,N_5891,N_5622);
xor U6748 (N_6748,N_4039,N_4171);
or U6749 (N_6749,N_4023,N_5224);
xnor U6750 (N_6750,N_4732,N_5533);
nand U6751 (N_6751,N_5038,N_5425);
nand U6752 (N_6752,N_4202,N_5661);
nand U6753 (N_6753,N_5953,N_5288);
or U6754 (N_6754,N_5963,N_4849);
and U6755 (N_6755,N_4146,N_5979);
nand U6756 (N_6756,N_4047,N_4530);
or U6757 (N_6757,N_5043,N_4686);
or U6758 (N_6758,N_4638,N_5683);
and U6759 (N_6759,N_5415,N_5480);
or U6760 (N_6760,N_4703,N_4189);
and U6761 (N_6761,N_5087,N_4529);
and U6762 (N_6762,N_4818,N_5284);
and U6763 (N_6763,N_4622,N_5429);
and U6764 (N_6764,N_4798,N_5313);
nand U6765 (N_6765,N_4114,N_5392);
or U6766 (N_6766,N_4541,N_5069);
nand U6767 (N_6767,N_5950,N_4864);
and U6768 (N_6768,N_5025,N_4625);
nand U6769 (N_6769,N_5155,N_4337);
nand U6770 (N_6770,N_5007,N_4368);
nand U6771 (N_6771,N_5379,N_5100);
and U6772 (N_6772,N_4813,N_4586);
nor U6773 (N_6773,N_5123,N_4920);
and U6774 (N_6774,N_5090,N_4962);
and U6775 (N_6775,N_4604,N_5469);
or U6776 (N_6776,N_5102,N_5578);
or U6777 (N_6777,N_4678,N_4946);
and U6778 (N_6778,N_5899,N_4819);
nor U6779 (N_6779,N_4773,N_5800);
nor U6780 (N_6780,N_5830,N_5344);
nand U6781 (N_6781,N_4452,N_5693);
xor U6782 (N_6782,N_5943,N_5372);
or U6783 (N_6783,N_5449,N_4524);
and U6784 (N_6784,N_5175,N_5657);
nand U6785 (N_6785,N_5916,N_5244);
nor U6786 (N_6786,N_5499,N_4770);
nor U6787 (N_6787,N_5839,N_4231);
or U6788 (N_6788,N_5136,N_4026);
nor U6789 (N_6789,N_5682,N_4701);
and U6790 (N_6790,N_4143,N_4388);
or U6791 (N_6791,N_5065,N_4453);
nor U6792 (N_6792,N_4646,N_4347);
or U6793 (N_6793,N_5140,N_5736);
nor U6794 (N_6794,N_5301,N_5825);
and U6795 (N_6795,N_4241,N_4953);
nor U6796 (N_6796,N_5589,N_4635);
nand U6797 (N_6797,N_4936,N_5315);
nor U6798 (N_6798,N_4259,N_5978);
and U6799 (N_6799,N_5260,N_5478);
and U6800 (N_6800,N_5549,N_4827);
nand U6801 (N_6801,N_4911,N_5042);
and U6802 (N_6802,N_5797,N_4075);
and U6803 (N_6803,N_4373,N_5998);
nor U6804 (N_6804,N_4003,N_5651);
or U6805 (N_6805,N_4091,N_5111);
nand U6806 (N_6806,N_5303,N_4540);
and U6807 (N_6807,N_5586,N_4265);
nand U6808 (N_6808,N_4310,N_5734);
or U6809 (N_6809,N_4670,N_4392);
or U6810 (N_6810,N_5710,N_4875);
nand U6811 (N_6811,N_4255,N_5120);
and U6812 (N_6812,N_4948,N_4535);
or U6813 (N_6813,N_4823,N_5374);
and U6814 (N_6814,N_4254,N_5811);
nand U6815 (N_6815,N_5215,N_5168);
nor U6816 (N_6816,N_5463,N_5716);
xor U6817 (N_6817,N_5474,N_4389);
nand U6818 (N_6818,N_4888,N_5388);
or U6819 (N_6819,N_5546,N_5684);
nor U6820 (N_6820,N_4521,N_5789);
nor U6821 (N_6821,N_5147,N_5091);
or U6822 (N_6822,N_5290,N_4956);
and U6823 (N_6823,N_5457,N_5105);
nand U6824 (N_6824,N_4422,N_5658);
or U6825 (N_6825,N_4832,N_4042);
nand U6826 (N_6826,N_4220,N_5626);
and U6827 (N_6827,N_4218,N_5088);
and U6828 (N_6828,N_5124,N_4236);
and U6829 (N_6829,N_5870,N_4065);
nand U6830 (N_6830,N_5491,N_5781);
nand U6831 (N_6831,N_5566,N_4735);
or U6832 (N_6832,N_4250,N_5247);
nand U6833 (N_6833,N_5216,N_4863);
or U6834 (N_6834,N_4523,N_4053);
nand U6835 (N_6835,N_4418,N_4916);
nor U6836 (N_6836,N_5319,N_5086);
nand U6837 (N_6837,N_5822,N_4520);
or U6838 (N_6838,N_4918,N_5944);
nand U6839 (N_6839,N_5028,N_5436);
and U6840 (N_6840,N_5467,N_5828);
nor U6841 (N_6841,N_5924,N_5633);
nor U6842 (N_6842,N_5617,N_4623);
and U6843 (N_6843,N_4546,N_4358);
and U6844 (N_6844,N_4273,N_4440);
nor U6845 (N_6845,N_4238,N_4240);
and U6846 (N_6846,N_4155,N_5652);
and U6847 (N_6847,N_5482,N_5199);
nor U6848 (N_6848,N_4276,N_4283);
xor U6849 (N_6849,N_4969,N_4934);
and U6850 (N_6850,N_4077,N_5542);
nand U6851 (N_6851,N_4269,N_4929);
and U6852 (N_6852,N_4878,N_5298);
or U6853 (N_6853,N_5445,N_5513);
or U6854 (N_6854,N_5707,N_4747);
xnor U6855 (N_6855,N_5055,N_5440);
or U6856 (N_6856,N_5353,N_4618);
nand U6857 (N_6857,N_5774,N_4676);
or U6858 (N_6858,N_4745,N_5705);
nor U6859 (N_6859,N_5349,N_5143);
nand U6860 (N_6860,N_4293,N_4200);
nand U6861 (N_6861,N_5972,N_5625);
xnor U6862 (N_6862,N_4578,N_4249);
or U6863 (N_6863,N_4121,N_4069);
and U6864 (N_6864,N_4333,N_4326);
nand U6865 (N_6865,N_4803,N_5049);
nor U6866 (N_6866,N_5130,N_4462);
and U6867 (N_6867,N_4581,N_5117);
nand U6868 (N_6868,N_5675,N_5708);
nand U6869 (N_6869,N_5571,N_4743);
or U6870 (N_6870,N_4954,N_4955);
nor U6871 (N_6871,N_4900,N_5191);
nand U6872 (N_6872,N_5173,N_5639);
or U6873 (N_6873,N_4294,N_5297);
or U6874 (N_6874,N_5269,N_5806);
nor U6875 (N_6875,N_4243,N_4873);
xor U6876 (N_6876,N_4492,N_5816);
or U6877 (N_6877,N_5507,N_4557);
nor U6878 (N_6878,N_4539,N_5074);
or U6879 (N_6879,N_5777,N_4507);
and U6880 (N_6880,N_5832,N_5732);
nand U6881 (N_6881,N_4239,N_4228);
and U6882 (N_6882,N_5547,N_4912);
or U6883 (N_6883,N_5538,N_4767);
and U6884 (N_6884,N_4585,N_5451);
and U6885 (N_6885,N_5036,N_5987);
or U6886 (N_6886,N_5210,N_5416);
and U6887 (N_6887,N_4322,N_4127);
nor U6888 (N_6888,N_4350,N_4494);
nand U6889 (N_6889,N_5362,N_5193);
and U6890 (N_6890,N_4654,N_4909);
or U6891 (N_6891,N_4846,N_5152);
nand U6892 (N_6892,N_5995,N_4024);
nor U6893 (N_6893,N_4754,N_5687);
and U6894 (N_6894,N_4715,N_4528);
nor U6895 (N_6895,N_4512,N_5949);
nand U6896 (N_6896,N_5234,N_5900);
nand U6897 (N_6897,N_4985,N_5957);
and U6898 (N_6898,N_5636,N_5737);
xnor U6899 (N_6899,N_5928,N_5790);
or U6900 (N_6900,N_4587,N_4631);
nand U6901 (N_6901,N_5550,N_5270);
or U6902 (N_6902,N_5326,N_4030);
and U6903 (N_6903,N_5494,N_4673);
nor U6904 (N_6904,N_5159,N_4588);
nand U6905 (N_6905,N_4435,N_5058);
or U6906 (N_6906,N_5302,N_5865);
nand U6907 (N_6907,N_5428,N_4501);
or U6908 (N_6908,N_5951,N_4534);
nor U6909 (N_6909,N_4592,N_4593);
nor U6910 (N_6910,N_4209,N_4553);
or U6911 (N_6911,N_5610,N_4338);
or U6912 (N_6912,N_5605,N_5815);
or U6913 (N_6913,N_5579,N_5061);
nand U6914 (N_6914,N_4225,N_5194);
xor U6915 (N_6915,N_4038,N_5624);
nor U6916 (N_6916,N_5960,N_4021);
nor U6917 (N_6917,N_4907,N_4677);
and U6918 (N_6918,N_4993,N_5115);
nor U6919 (N_6919,N_4950,N_4385);
xor U6920 (N_6920,N_4756,N_5975);
and U6921 (N_6921,N_4428,N_4870);
nand U6922 (N_6922,N_5417,N_5909);
and U6923 (N_6923,N_5614,N_5354);
xor U6924 (N_6924,N_4312,N_5545);
or U6925 (N_6925,N_4497,N_5295);
nor U6926 (N_6926,N_5277,N_4285);
nand U6927 (N_6927,N_4321,N_4762);
nand U6928 (N_6928,N_5439,N_4165);
or U6929 (N_6929,N_5406,N_5035);
and U6930 (N_6930,N_5678,N_4315);
or U6931 (N_6931,N_5004,N_5235);
nand U6932 (N_6932,N_4319,N_5373);
nor U6933 (N_6933,N_4506,N_4648);
nor U6934 (N_6934,N_4872,N_5363);
nand U6935 (N_6935,N_5287,N_5422);
or U6936 (N_6936,N_4669,N_4415);
and U6937 (N_6937,N_4344,N_5746);
nor U6938 (N_6938,N_4595,N_4012);
or U6939 (N_6939,N_4080,N_4567);
nor U6940 (N_6940,N_4990,N_4235);
and U6941 (N_6941,N_5040,N_4889);
or U6942 (N_6942,N_4266,N_5384);
nand U6943 (N_6943,N_5834,N_4139);
or U6944 (N_6944,N_4952,N_5532);
or U6945 (N_6945,N_5941,N_4928);
nor U6946 (N_6946,N_4367,N_5204);
nand U6947 (N_6947,N_4584,N_5719);
or U6948 (N_6948,N_5991,N_5386);
nand U6949 (N_6949,N_4463,N_5603);
and U6950 (N_6950,N_4660,N_4182);
or U6951 (N_6951,N_5827,N_4537);
nor U6952 (N_6952,N_5227,N_4572);
and U6953 (N_6953,N_5555,N_4886);
and U6954 (N_6954,N_5691,N_5570);
nand U6955 (N_6955,N_5283,N_5685);
or U6956 (N_6956,N_4097,N_5638);
nand U6957 (N_6957,N_4116,N_5939);
or U6958 (N_6958,N_4317,N_4439);
nand U6959 (N_6959,N_4815,N_4937);
nor U6960 (N_6960,N_4667,N_5593);
nand U6961 (N_6961,N_5342,N_4904);
or U6962 (N_6962,N_5488,N_5609);
nor U6963 (N_6963,N_5659,N_4426);
xor U6964 (N_6964,N_5157,N_5653);
or U6965 (N_6965,N_5643,N_5167);
nor U6966 (N_6966,N_4183,N_5114);
nor U6967 (N_6967,N_4331,N_4636);
nand U6968 (N_6968,N_4037,N_5003);
xnor U6969 (N_6969,N_4369,N_4318);
or U6970 (N_6970,N_5856,N_5129);
nor U6971 (N_6971,N_5526,N_5926);
or U6972 (N_6972,N_4477,N_4274);
nor U6973 (N_6973,N_4927,N_5030);
and U6974 (N_6974,N_5680,N_5674);
and U6975 (N_6975,N_4645,N_4683);
nand U6976 (N_6976,N_5263,N_5441);
and U6977 (N_6977,N_5842,N_4260);
or U6978 (N_6978,N_4125,N_4057);
nor U6979 (N_6979,N_4679,N_5420);
nor U6980 (N_6980,N_4416,N_5476);
nand U6981 (N_6981,N_4842,N_5364);
nand U6982 (N_6982,N_5554,N_5587);
or U6983 (N_6983,N_4649,N_4495);
and U6984 (N_6984,N_4140,N_5648);
and U6985 (N_6985,N_4689,N_5623);
or U6986 (N_6986,N_4989,N_5011);
nor U6987 (N_6987,N_5312,N_4999);
and U6988 (N_6988,N_5271,N_4208);
and U6989 (N_6989,N_5612,N_4450);
and U6990 (N_6990,N_5907,N_5590);
and U6991 (N_6991,N_4691,N_4193);
or U6992 (N_6992,N_5323,N_4629);
or U6993 (N_6993,N_4865,N_4700);
nor U6994 (N_6994,N_4295,N_5402);
xnor U6995 (N_6995,N_4212,N_4619);
nor U6996 (N_6996,N_5456,N_5628);
nor U6997 (N_6997,N_5138,N_4958);
nand U6998 (N_6998,N_4880,N_4730);
nand U6999 (N_6999,N_5424,N_5893);
and U7000 (N_7000,N_5126,N_5567);
or U7001 (N_7001,N_5968,N_4962);
xor U7002 (N_7002,N_5080,N_4969);
nand U7003 (N_7003,N_4021,N_5656);
nand U7004 (N_7004,N_5327,N_5884);
nand U7005 (N_7005,N_4931,N_4557);
nand U7006 (N_7006,N_5200,N_4976);
and U7007 (N_7007,N_4907,N_4275);
or U7008 (N_7008,N_5434,N_5061);
nor U7009 (N_7009,N_4166,N_5261);
and U7010 (N_7010,N_5287,N_4605);
nand U7011 (N_7011,N_5614,N_5111);
nand U7012 (N_7012,N_5026,N_5961);
or U7013 (N_7013,N_5857,N_5504);
nor U7014 (N_7014,N_5978,N_4760);
nor U7015 (N_7015,N_5976,N_5320);
or U7016 (N_7016,N_5804,N_4356);
or U7017 (N_7017,N_4602,N_4631);
and U7018 (N_7018,N_4021,N_4642);
xnor U7019 (N_7019,N_5161,N_4699);
or U7020 (N_7020,N_5205,N_5687);
and U7021 (N_7021,N_5551,N_5867);
xnor U7022 (N_7022,N_5365,N_4867);
xnor U7023 (N_7023,N_5965,N_4052);
nand U7024 (N_7024,N_4535,N_5306);
and U7025 (N_7025,N_4064,N_4984);
and U7026 (N_7026,N_4084,N_4778);
and U7027 (N_7027,N_5862,N_5732);
or U7028 (N_7028,N_5533,N_4861);
and U7029 (N_7029,N_4232,N_4851);
nor U7030 (N_7030,N_5728,N_4941);
and U7031 (N_7031,N_5040,N_4731);
or U7032 (N_7032,N_5129,N_5494);
xnor U7033 (N_7033,N_4643,N_5819);
or U7034 (N_7034,N_4517,N_5152);
xor U7035 (N_7035,N_4767,N_4654);
nand U7036 (N_7036,N_4187,N_4204);
or U7037 (N_7037,N_5341,N_4831);
nor U7038 (N_7038,N_4336,N_5223);
nand U7039 (N_7039,N_5957,N_5265);
nand U7040 (N_7040,N_4304,N_4056);
or U7041 (N_7041,N_4831,N_5722);
nand U7042 (N_7042,N_5222,N_5820);
xnor U7043 (N_7043,N_5763,N_5632);
or U7044 (N_7044,N_4276,N_5765);
xor U7045 (N_7045,N_4554,N_5491);
nor U7046 (N_7046,N_4214,N_5247);
nand U7047 (N_7047,N_4340,N_5467);
nand U7048 (N_7048,N_5843,N_5722);
and U7049 (N_7049,N_4721,N_5142);
and U7050 (N_7050,N_4558,N_5161);
or U7051 (N_7051,N_4662,N_4707);
and U7052 (N_7052,N_4633,N_4518);
nor U7053 (N_7053,N_4412,N_4233);
and U7054 (N_7054,N_5363,N_4868);
and U7055 (N_7055,N_4789,N_4393);
nand U7056 (N_7056,N_4354,N_5668);
nor U7057 (N_7057,N_5140,N_5925);
or U7058 (N_7058,N_4008,N_5865);
or U7059 (N_7059,N_5112,N_5218);
nand U7060 (N_7060,N_5365,N_4830);
nor U7061 (N_7061,N_5134,N_5579);
nand U7062 (N_7062,N_5201,N_5494);
xnor U7063 (N_7063,N_4981,N_5942);
and U7064 (N_7064,N_5149,N_4806);
or U7065 (N_7065,N_4302,N_4602);
nor U7066 (N_7066,N_5455,N_5396);
or U7067 (N_7067,N_4188,N_5308);
and U7068 (N_7068,N_5568,N_5325);
and U7069 (N_7069,N_5361,N_5391);
nor U7070 (N_7070,N_4560,N_4444);
nor U7071 (N_7071,N_4568,N_4169);
and U7072 (N_7072,N_4067,N_5629);
or U7073 (N_7073,N_5434,N_4964);
xnor U7074 (N_7074,N_4355,N_5814);
nor U7075 (N_7075,N_4786,N_5212);
or U7076 (N_7076,N_5920,N_5293);
and U7077 (N_7077,N_4652,N_4829);
nor U7078 (N_7078,N_4903,N_4120);
nor U7079 (N_7079,N_5802,N_5301);
and U7080 (N_7080,N_4785,N_4554);
nand U7081 (N_7081,N_4349,N_4544);
nor U7082 (N_7082,N_4714,N_5690);
nor U7083 (N_7083,N_5221,N_5264);
nand U7084 (N_7084,N_5605,N_5000);
or U7085 (N_7085,N_4530,N_4251);
and U7086 (N_7086,N_4093,N_5232);
or U7087 (N_7087,N_5896,N_4318);
nor U7088 (N_7088,N_5098,N_5019);
or U7089 (N_7089,N_5759,N_5356);
nand U7090 (N_7090,N_5901,N_4691);
and U7091 (N_7091,N_5608,N_4922);
and U7092 (N_7092,N_5556,N_5074);
and U7093 (N_7093,N_4025,N_5687);
nor U7094 (N_7094,N_4391,N_4316);
and U7095 (N_7095,N_4457,N_5282);
and U7096 (N_7096,N_5632,N_5955);
nand U7097 (N_7097,N_5236,N_4767);
and U7098 (N_7098,N_4760,N_5524);
and U7099 (N_7099,N_5506,N_4537);
and U7100 (N_7100,N_4247,N_5227);
nand U7101 (N_7101,N_4251,N_5019);
or U7102 (N_7102,N_5617,N_5575);
and U7103 (N_7103,N_5244,N_5441);
nand U7104 (N_7104,N_5865,N_4423);
nand U7105 (N_7105,N_4609,N_4214);
nor U7106 (N_7106,N_5690,N_5131);
nand U7107 (N_7107,N_5809,N_4283);
nor U7108 (N_7108,N_5749,N_5957);
nand U7109 (N_7109,N_4323,N_5879);
nor U7110 (N_7110,N_5998,N_4689);
nand U7111 (N_7111,N_5891,N_4470);
xnor U7112 (N_7112,N_4259,N_4640);
nand U7113 (N_7113,N_4607,N_5996);
and U7114 (N_7114,N_5295,N_4670);
nand U7115 (N_7115,N_4664,N_5561);
or U7116 (N_7116,N_5258,N_4157);
and U7117 (N_7117,N_5907,N_5490);
nor U7118 (N_7118,N_4184,N_4374);
nor U7119 (N_7119,N_5745,N_5562);
xor U7120 (N_7120,N_4998,N_4271);
and U7121 (N_7121,N_4340,N_4804);
nand U7122 (N_7122,N_5299,N_5083);
nand U7123 (N_7123,N_5962,N_4643);
and U7124 (N_7124,N_5580,N_4298);
nor U7125 (N_7125,N_4689,N_5483);
nand U7126 (N_7126,N_5723,N_4211);
nand U7127 (N_7127,N_4001,N_5227);
or U7128 (N_7128,N_5061,N_4333);
nor U7129 (N_7129,N_5855,N_5413);
or U7130 (N_7130,N_4546,N_5756);
nor U7131 (N_7131,N_5382,N_5117);
nand U7132 (N_7132,N_4192,N_5634);
or U7133 (N_7133,N_5374,N_5743);
and U7134 (N_7134,N_4651,N_4168);
or U7135 (N_7135,N_4428,N_5148);
xnor U7136 (N_7136,N_5550,N_4084);
nand U7137 (N_7137,N_5923,N_4183);
nand U7138 (N_7138,N_5924,N_5314);
nand U7139 (N_7139,N_4876,N_5462);
or U7140 (N_7140,N_4975,N_5456);
or U7141 (N_7141,N_5397,N_4260);
nand U7142 (N_7142,N_4445,N_5192);
or U7143 (N_7143,N_4272,N_5549);
nand U7144 (N_7144,N_5436,N_4343);
nand U7145 (N_7145,N_5284,N_4775);
xnor U7146 (N_7146,N_4604,N_5620);
xor U7147 (N_7147,N_5625,N_5739);
and U7148 (N_7148,N_4221,N_4951);
or U7149 (N_7149,N_4340,N_4723);
nand U7150 (N_7150,N_4276,N_5977);
or U7151 (N_7151,N_5611,N_5243);
nand U7152 (N_7152,N_5470,N_5028);
nor U7153 (N_7153,N_4509,N_4153);
and U7154 (N_7154,N_5121,N_5930);
nor U7155 (N_7155,N_5828,N_5108);
xor U7156 (N_7156,N_4649,N_4869);
and U7157 (N_7157,N_4384,N_4577);
nor U7158 (N_7158,N_4870,N_5131);
nand U7159 (N_7159,N_5506,N_4186);
or U7160 (N_7160,N_5150,N_4191);
or U7161 (N_7161,N_5837,N_5954);
and U7162 (N_7162,N_4158,N_5468);
and U7163 (N_7163,N_5102,N_4490);
nand U7164 (N_7164,N_4757,N_5028);
xor U7165 (N_7165,N_5965,N_5238);
and U7166 (N_7166,N_4850,N_5448);
or U7167 (N_7167,N_4533,N_5557);
xor U7168 (N_7168,N_4787,N_5035);
and U7169 (N_7169,N_5698,N_4050);
and U7170 (N_7170,N_5556,N_4889);
xnor U7171 (N_7171,N_4084,N_5058);
nor U7172 (N_7172,N_5216,N_5653);
nor U7173 (N_7173,N_5663,N_4996);
nand U7174 (N_7174,N_5765,N_4780);
xor U7175 (N_7175,N_4581,N_4264);
nor U7176 (N_7176,N_5768,N_5649);
or U7177 (N_7177,N_5426,N_5458);
xnor U7178 (N_7178,N_4227,N_5453);
or U7179 (N_7179,N_5933,N_5455);
xor U7180 (N_7180,N_5320,N_5305);
or U7181 (N_7181,N_5746,N_5446);
and U7182 (N_7182,N_5095,N_5689);
or U7183 (N_7183,N_4756,N_4855);
nand U7184 (N_7184,N_5456,N_5559);
nor U7185 (N_7185,N_4264,N_5289);
nor U7186 (N_7186,N_4337,N_5246);
xor U7187 (N_7187,N_4547,N_5821);
nand U7188 (N_7188,N_5713,N_5670);
nor U7189 (N_7189,N_5110,N_5455);
or U7190 (N_7190,N_5485,N_5055);
and U7191 (N_7191,N_5353,N_5627);
or U7192 (N_7192,N_5485,N_4712);
nand U7193 (N_7193,N_4109,N_4115);
xor U7194 (N_7194,N_4170,N_5431);
nand U7195 (N_7195,N_4706,N_5690);
nand U7196 (N_7196,N_5246,N_5849);
nand U7197 (N_7197,N_5539,N_5019);
nand U7198 (N_7198,N_4724,N_4666);
or U7199 (N_7199,N_4323,N_4757);
nand U7200 (N_7200,N_5025,N_5349);
or U7201 (N_7201,N_4547,N_4139);
or U7202 (N_7202,N_4789,N_5943);
or U7203 (N_7203,N_5881,N_5449);
nor U7204 (N_7204,N_4408,N_4256);
or U7205 (N_7205,N_5100,N_4792);
nor U7206 (N_7206,N_5919,N_4983);
nand U7207 (N_7207,N_4854,N_4766);
nor U7208 (N_7208,N_5671,N_5161);
and U7209 (N_7209,N_4789,N_4449);
or U7210 (N_7210,N_5939,N_5848);
and U7211 (N_7211,N_4298,N_5640);
and U7212 (N_7212,N_4181,N_5656);
or U7213 (N_7213,N_4853,N_4661);
xor U7214 (N_7214,N_4732,N_4276);
and U7215 (N_7215,N_5241,N_5126);
and U7216 (N_7216,N_4141,N_4473);
nand U7217 (N_7217,N_5869,N_5434);
and U7218 (N_7218,N_4563,N_5959);
xor U7219 (N_7219,N_4554,N_4437);
and U7220 (N_7220,N_5077,N_4913);
nand U7221 (N_7221,N_5892,N_4950);
and U7222 (N_7222,N_5927,N_4966);
nand U7223 (N_7223,N_5911,N_4769);
or U7224 (N_7224,N_5322,N_5514);
nor U7225 (N_7225,N_4303,N_5987);
xor U7226 (N_7226,N_5176,N_5556);
or U7227 (N_7227,N_4691,N_5617);
xor U7228 (N_7228,N_5854,N_4838);
nor U7229 (N_7229,N_4912,N_5290);
or U7230 (N_7230,N_5656,N_4281);
and U7231 (N_7231,N_5799,N_4775);
or U7232 (N_7232,N_4469,N_4017);
nand U7233 (N_7233,N_4152,N_5337);
or U7234 (N_7234,N_5052,N_5053);
and U7235 (N_7235,N_4753,N_5202);
nand U7236 (N_7236,N_5379,N_5748);
nand U7237 (N_7237,N_5026,N_5505);
nand U7238 (N_7238,N_4573,N_4859);
nand U7239 (N_7239,N_5874,N_4221);
nor U7240 (N_7240,N_4405,N_4550);
nand U7241 (N_7241,N_4971,N_5700);
xor U7242 (N_7242,N_5397,N_5481);
xor U7243 (N_7243,N_4527,N_4005);
or U7244 (N_7244,N_4582,N_5409);
nand U7245 (N_7245,N_4701,N_5929);
nand U7246 (N_7246,N_5377,N_5114);
nor U7247 (N_7247,N_5224,N_5343);
nand U7248 (N_7248,N_4646,N_5862);
and U7249 (N_7249,N_5436,N_4158);
or U7250 (N_7250,N_5586,N_5847);
and U7251 (N_7251,N_5390,N_4706);
or U7252 (N_7252,N_4101,N_4716);
or U7253 (N_7253,N_5055,N_5988);
xnor U7254 (N_7254,N_5326,N_4883);
nand U7255 (N_7255,N_4561,N_5029);
or U7256 (N_7256,N_5640,N_5475);
nand U7257 (N_7257,N_4024,N_4277);
or U7258 (N_7258,N_5353,N_4819);
nand U7259 (N_7259,N_5357,N_4988);
and U7260 (N_7260,N_4638,N_5174);
and U7261 (N_7261,N_5676,N_4397);
nand U7262 (N_7262,N_5025,N_4569);
xnor U7263 (N_7263,N_4972,N_4471);
and U7264 (N_7264,N_5000,N_4753);
nand U7265 (N_7265,N_5349,N_5718);
and U7266 (N_7266,N_4673,N_5529);
xor U7267 (N_7267,N_4220,N_5912);
nand U7268 (N_7268,N_4483,N_4830);
and U7269 (N_7269,N_4872,N_5776);
or U7270 (N_7270,N_4986,N_4956);
xor U7271 (N_7271,N_5122,N_4593);
nand U7272 (N_7272,N_4271,N_4657);
nand U7273 (N_7273,N_5859,N_4348);
and U7274 (N_7274,N_4124,N_5365);
and U7275 (N_7275,N_5349,N_4639);
nand U7276 (N_7276,N_5836,N_4067);
or U7277 (N_7277,N_5972,N_5045);
nor U7278 (N_7278,N_4855,N_4597);
or U7279 (N_7279,N_5675,N_4891);
nor U7280 (N_7280,N_5872,N_5955);
and U7281 (N_7281,N_4166,N_5830);
nand U7282 (N_7282,N_5783,N_4362);
and U7283 (N_7283,N_4788,N_5282);
nand U7284 (N_7284,N_4974,N_4576);
nand U7285 (N_7285,N_5549,N_4961);
nor U7286 (N_7286,N_4448,N_4831);
nand U7287 (N_7287,N_4105,N_5958);
and U7288 (N_7288,N_5535,N_5434);
and U7289 (N_7289,N_5445,N_5416);
nor U7290 (N_7290,N_4804,N_4438);
nand U7291 (N_7291,N_4799,N_4940);
and U7292 (N_7292,N_4533,N_4591);
nor U7293 (N_7293,N_4184,N_5725);
xnor U7294 (N_7294,N_4373,N_5452);
and U7295 (N_7295,N_5232,N_5083);
and U7296 (N_7296,N_5929,N_4758);
nor U7297 (N_7297,N_4407,N_5211);
nor U7298 (N_7298,N_4311,N_5065);
and U7299 (N_7299,N_5936,N_5906);
nand U7300 (N_7300,N_5031,N_5806);
nor U7301 (N_7301,N_4887,N_5270);
nand U7302 (N_7302,N_4141,N_5493);
nor U7303 (N_7303,N_5113,N_4398);
nor U7304 (N_7304,N_5133,N_4352);
nand U7305 (N_7305,N_5957,N_4844);
and U7306 (N_7306,N_4347,N_5586);
xor U7307 (N_7307,N_4844,N_4917);
nand U7308 (N_7308,N_4918,N_5556);
nor U7309 (N_7309,N_5882,N_4038);
or U7310 (N_7310,N_4495,N_5285);
and U7311 (N_7311,N_4390,N_4788);
and U7312 (N_7312,N_5670,N_5572);
xnor U7313 (N_7313,N_5428,N_4924);
or U7314 (N_7314,N_4087,N_4484);
nand U7315 (N_7315,N_4916,N_5778);
nand U7316 (N_7316,N_5073,N_5592);
and U7317 (N_7317,N_5658,N_4500);
nor U7318 (N_7318,N_4019,N_5035);
nor U7319 (N_7319,N_4099,N_5762);
and U7320 (N_7320,N_5647,N_5461);
nor U7321 (N_7321,N_5300,N_5183);
nor U7322 (N_7322,N_5781,N_5846);
nand U7323 (N_7323,N_4255,N_4696);
nand U7324 (N_7324,N_5949,N_4145);
nor U7325 (N_7325,N_5507,N_5254);
or U7326 (N_7326,N_5061,N_5363);
nor U7327 (N_7327,N_5631,N_5827);
nand U7328 (N_7328,N_4233,N_5390);
or U7329 (N_7329,N_5395,N_5796);
and U7330 (N_7330,N_5891,N_5400);
and U7331 (N_7331,N_4906,N_4668);
nor U7332 (N_7332,N_4907,N_5842);
and U7333 (N_7333,N_4926,N_4596);
and U7334 (N_7334,N_4254,N_5834);
nand U7335 (N_7335,N_5048,N_4124);
and U7336 (N_7336,N_4067,N_5783);
and U7337 (N_7337,N_4767,N_4132);
or U7338 (N_7338,N_4525,N_4991);
or U7339 (N_7339,N_5290,N_5547);
nor U7340 (N_7340,N_4084,N_5342);
and U7341 (N_7341,N_5577,N_4235);
nand U7342 (N_7342,N_4247,N_4011);
or U7343 (N_7343,N_5975,N_5153);
and U7344 (N_7344,N_4957,N_5356);
nor U7345 (N_7345,N_5415,N_5022);
xnor U7346 (N_7346,N_4768,N_4479);
xnor U7347 (N_7347,N_5918,N_5213);
xnor U7348 (N_7348,N_4489,N_4023);
nand U7349 (N_7349,N_5580,N_4885);
nor U7350 (N_7350,N_5346,N_4976);
xnor U7351 (N_7351,N_4224,N_4598);
or U7352 (N_7352,N_5308,N_4317);
and U7353 (N_7353,N_5178,N_4242);
or U7354 (N_7354,N_5859,N_5663);
xor U7355 (N_7355,N_4113,N_4967);
and U7356 (N_7356,N_4488,N_5277);
nand U7357 (N_7357,N_5961,N_4321);
and U7358 (N_7358,N_4071,N_5270);
and U7359 (N_7359,N_4635,N_5080);
nor U7360 (N_7360,N_4801,N_4416);
nand U7361 (N_7361,N_4958,N_4225);
and U7362 (N_7362,N_5824,N_5081);
and U7363 (N_7363,N_4083,N_4209);
nand U7364 (N_7364,N_4574,N_4186);
and U7365 (N_7365,N_5205,N_5615);
and U7366 (N_7366,N_4479,N_4000);
or U7367 (N_7367,N_4367,N_4183);
or U7368 (N_7368,N_4069,N_5593);
and U7369 (N_7369,N_5739,N_5909);
and U7370 (N_7370,N_4937,N_5985);
nor U7371 (N_7371,N_5938,N_5036);
nor U7372 (N_7372,N_4002,N_4413);
and U7373 (N_7373,N_5190,N_5646);
and U7374 (N_7374,N_5014,N_4541);
nand U7375 (N_7375,N_4174,N_5045);
nor U7376 (N_7376,N_4517,N_4539);
xnor U7377 (N_7377,N_4442,N_4105);
nor U7378 (N_7378,N_4282,N_4064);
nand U7379 (N_7379,N_5956,N_4386);
and U7380 (N_7380,N_5918,N_5682);
or U7381 (N_7381,N_5021,N_4188);
and U7382 (N_7382,N_4187,N_4044);
and U7383 (N_7383,N_5353,N_4592);
nor U7384 (N_7384,N_4925,N_5161);
nor U7385 (N_7385,N_4735,N_5885);
or U7386 (N_7386,N_4989,N_4541);
and U7387 (N_7387,N_5121,N_5304);
or U7388 (N_7388,N_4526,N_4560);
and U7389 (N_7389,N_4321,N_4693);
nor U7390 (N_7390,N_5403,N_5544);
nor U7391 (N_7391,N_5713,N_4839);
nand U7392 (N_7392,N_4516,N_4705);
or U7393 (N_7393,N_4579,N_5581);
nor U7394 (N_7394,N_5013,N_4850);
nor U7395 (N_7395,N_4556,N_4539);
nor U7396 (N_7396,N_5445,N_4624);
or U7397 (N_7397,N_4660,N_5071);
or U7398 (N_7398,N_4097,N_5383);
nand U7399 (N_7399,N_5283,N_5689);
nand U7400 (N_7400,N_4630,N_5194);
xor U7401 (N_7401,N_4060,N_4812);
and U7402 (N_7402,N_5562,N_5548);
nand U7403 (N_7403,N_4230,N_4501);
and U7404 (N_7404,N_4462,N_5115);
nand U7405 (N_7405,N_4730,N_4417);
or U7406 (N_7406,N_4749,N_5725);
nor U7407 (N_7407,N_5703,N_4937);
nor U7408 (N_7408,N_4755,N_4883);
or U7409 (N_7409,N_4037,N_5578);
nor U7410 (N_7410,N_5228,N_4741);
or U7411 (N_7411,N_4220,N_4560);
and U7412 (N_7412,N_4876,N_4592);
and U7413 (N_7413,N_5081,N_4444);
or U7414 (N_7414,N_5794,N_4431);
and U7415 (N_7415,N_5117,N_5454);
and U7416 (N_7416,N_4723,N_5594);
or U7417 (N_7417,N_4991,N_5188);
nor U7418 (N_7418,N_4556,N_5748);
nor U7419 (N_7419,N_5451,N_4601);
nor U7420 (N_7420,N_4422,N_4360);
and U7421 (N_7421,N_5216,N_5360);
nand U7422 (N_7422,N_4962,N_5481);
nor U7423 (N_7423,N_5647,N_4457);
nand U7424 (N_7424,N_4249,N_4179);
or U7425 (N_7425,N_4665,N_4856);
nor U7426 (N_7426,N_5627,N_4029);
and U7427 (N_7427,N_5912,N_4175);
nand U7428 (N_7428,N_5644,N_5977);
or U7429 (N_7429,N_5792,N_4730);
and U7430 (N_7430,N_5658,N_4474);
nand U7431 (N_7431,N_5419,N_5272);
nor U7432 (N_7432,N_5535,N_5500);
or U7433 (N_7433,N_4150,N_4498);
xnor U7434 (N_7434,N_5123,N_4268);
nand U7435 (N_7435,N_5902,N_5880);
or U7436 (N_7436,N_4598,N_5930);
nand U7437 (N_7437,N_5675,N_5402);
nor U7438 (N_7438,N_4302,N_4790);
or U7439 (N_7439,N_4844,N_5919);
and U7440 (N_7440,N_5767,N_4335);
xor U7441 (N_7441,N_5571,N_4771);
nor U7442 (N_7442,N_4472,N_4917);
xnor U7443 (N_7443,N_4983,N_4271);
and U7444 (N_7444,N_4916,N_5454);
or U7445 (N_7445,N_4059,N_5551);
nand U7446 (N_7446,N_4734,N_4406);
and U7447 (N_7447,N_4312,N_4600);
and U7448 (N_7448,N_5455,N_4085);
nand U7449 (N_7449,N_5719,N_4945);
or U7450 (N_7450,N_4601,N_4118);
and U7451 (N_7451,N_5270,N_4741);
or U7452 (N_7452,N_5568,N_5925);
or U7453 (N_7453,N_5383,N_4386);
xor U7454 (N_7454,N_5199,N_4232);
nand U7455 (N_7455,N_4790,N_5769);
nor U7456 (N_7456,N_4418,N_5187);
and U7457 (N_7457,N_5759,N_5758);
or U7458 (N_7458,N_5180,N_5037);
and U7459 (N_7459,N_4409,N_4994);
nand U7460 (N_7460,N_4035,N_4659);
xnor U7461 (N_7461,N_4916,N_5647);
and U7462 (N_7462,N_4948,N_5823);
xnor U7463 (N_7463,N_4394,N_4221);
nand U7464 (N_7464,N_5251,N_5125);
nor U7465 (N_7465,N_5962,N_5982);
xnor U7466 (N_7466,N_4132,N_5180);
nand U7467 (N_7467,N_4115,N_4190);
or U7468 (N_7468,N_4179,N_5062);
xnor U7469 (N_7469,N_4665,N_5056);
or U7470 (N_7470,N_4963,N_5358);
xnor U7471 (N_7471,N_4002,N_4948);
nor U7472 (N_7472,N_5169,N_5536);
nand U7473 (N_7473,N_4460,N_5520);
and U7474 (N_7474,N_5431,N_4434);
nor U7475 (N_7475,N_4834,N_5161);
or U7476 (N_7476,N_5043,N_4427);
nand U7477 (N_7477,N_5977,N_4192);
and U7478 (N_7478,N_4924,N_4744);
nand U7479 (N_7479,N_5073,N_5325);
xor U7480 (N_7480,N_4700,N_5168);
or U7481 (N_7481,N_4498,N_5617);
nand U7482 (N_7482,N_4988,N_5218);
or U7483 (N_7483,N_4470,N_4955);
nor U7484 (N_7484,N_4352,N_4793);
nor U7485 (N_7485,N_4324,N_5945);
xor U7486 (N_7486,N_5734,N_4316);
or U7487 (N_7487,N_4102,N_5304);
xnor U7488 (N_7488,N_4557,N_4189);
and U7489 (N_7489,N_4502,N_5899);
nand U7490 (N_7490,N_5804,N_4882);
nor U7491 (N_7491,N_4253,N_5068);
or U7492 (N_7492,N_5608,N_4313);
nand U7493 (N_7493,N_4544,N_4624);
xnor U7494 (N_7494,N_5085,N_5355);
and U7495 (N_7495,N_4086,N_5972);
and U7496 (N_7496,N_4816,N_5528);
nand U7497 (N_7497,N_4173,N_4564);
nor U7498 (N_7498,N_4319,N_5239);
or U7499 (N_7499,N_4905,N_5413);
nand U7500 (N_7500,N_5414,N_5117);
nor U7501 (N_7501,N_4829,N_4709);
nand U7502 (N_7502,N_5812,N_4390);
or U7503 (N_7503,N_4529,N_5513);
nand U7504 (N_7504,N_4262,N_5489);
nor U7505 (N_7505,N_4339,N_4142);
nand U7506 (N_7506,N_5649,N_5338);
xor U7507 (N_7507,N_4279,N_5181);
xnor U7508 (N_7508,N_4360,N_4684);
nor U7509 (N_7509,N_4402,N_4034);
nand U7510 (N_7510,N_5914,N_5041);
nand U7511 (N_7511,N_4861,N_5712);
nor U7512 (N_7512,N_4636,N_5945);
or U7513 (N_7513,N_5505,N_5503);
and U7514 (N_7514,N_5050,N_5392);
or U7515 (N_7515,N_5428,N_5723);
nor U7516 (N_7516,N_5048,N_4664);
nor U7517 (N_7517,N_5551,N_5422);
xor U7518 (N_7518,N_5026,N_5815);
nor U7519 (N_7519,N_5205,N_4063);
or U7520 (N_7520,N_5566,N_5924);
nand U7521 (N_7521,N_4160,N_4741);
nand U7522 (N_7522,N_4850,N_4770);
or U7523 (N_7523,N_4017,N_4121);
and U7524 (N_7524,N_4776,N_4361);
and U7525 (N_7525,N_5180,N_5142);
nor U7526 (N_7526,N_5691,N_5044);
nand U7527 (N_7527,N_5049,N_4460);
nand U7528 (N_7528,N_5757,N_4609);
and U7529 (N_7529,N_5653,N_4595);
xnor U7530 (N_7530,N_5694,N_5577);
and U7531 (N_7531,N_5038,N_5141);
or U7532 (N_7532,N_5439,N_5663);
nand U7533 (N_7533,N_5263,N_4547);
and U7534 (N_7534,N_5389,N_5500);
nor U7535 (N_7535,N_4728,N_4683);
nand U7536 (N_7536,N_4306,N_4988);
or U7537 (N_7537,N_5274,N_4532);
or U7538 (N_7538,N_5906,N_5148);
nor U7539 (N_7539,N_4083,N_5889);
nor U7540 (N_7540,N_4732,N_5577);
or U7541 (N_7541,N_4913,N_4143);
nand U7542 (N_7542,N_5319,N_5212);
xnor U7543 (N_7543,N_4434,N_5928);
and U7544 (N_7544,N_5032,N_4743);
or U7545 (N_7545,N_5647,N_5733);
and U7546 (N_7546,N_4536,N_4104);
nand U7547 (N_7547,N_4612,N_4175);
and U7548 (N_7548,N_5012,N_4804);
or U7549 (N_7549,N_4058,N_5348);
xnor U7550 (N_7550,N_4708,N_4111);
nor U7551 (N_7551,N_5881,N_5448);
and U7552 (N_7552,N_5056,N_4798);
nor U7553 (N_7553,N_4431,N_4185);
or U7554 (N_7554,N_5975,N_5013);
or U7555 (N_7555,N_4341,N_4318);
and U7556 (N_7556,N_5926,N_5850);
nand U7557 (N_7557,N_5827,N_5527);
nand U7558 (N_7558,N_5018,N_4827);
nand U7559 (N_7559,N_5614,N_4845);
nor U7560 (N_7560,N_5696,N_5859);
and U7561 (N_7561,N_5348,N_4867);
nand U7562 (N_7562,N_5565,N_5594);
nor U7563 (N_7563,N_4291,N_4156);
nand U7564 (N_7564,N_5755,N_5893);
or U7565 (N_7565,N_4911,N_4197);
nor U7566 (N_7566,N_5192,N_4458);
or U7567 (N_7567,N_5887,N_5053);
and U7568 (N_7568,N_4497,N_4671);
nor U7569 (N_7569,N_5477,N_5948);
nand U7570 (N_7570,N_5979,N_5820);
or U7571 (N_7571,N_4694,N_4354);
and U7572 (N_7572,N_4370,N_4854);
and U7573 (N_7573,N_5100,N_4386);
nand U7574 (N_7574,N_5055,N_4589);
and U7575 (N_7575,N_5519,N_4955);
or U7576 (N_7576,N_4055,N_4496);
and U7577 (N_7577,N_5812,N_5816);
or U7578 (N_7578,N_5763,N_5127);
or U7579 (N_7579,N_4586,N_4195);
or U7580 (N_7580,N_4200,N_5282);
or U7581 (N_7581,N_5930,N_5586);
and U7582 (N_7582,N_4213,N_4174);
nand U7583 (N_7583,N_5922,N_4074);
xnor U7584 (N_7584,N_4623,N_4421);
or U7585 (N_7585,N_4213,N_4674);
nor U7586 (N_7586,N_4798,N_4473);
nor U7587 (N_7587,N_5188,N_4016);
nor U7588 (N_7588,N_4865,N_5009);
and U7589 (N_7589,N_5669,N_5363);
nand U7590 (N_7590,N_4244,N_4430);
nor U7591 (N_7591,N_4662,N_5542);
xnor U7592 (N_7592,N_5356,N_4635);
or U7593 (N_7593,N_5474,N_4513);
or U7594 (N_7594,N_4333,N_4048);
or U7595 (N_7595,N_5627,N_5366);
and U7596 (N_7596,N_4824,N_4940);
nand U7597 (N_7597,N_4356,N_4075);
xnor U7598 (N_7598,N_5023,N_5971);
nand U7599 (N_7599,N_5771,N_4123);
and U7600 (N_7600,N_4967,N_5522);
and U7601 (N_7601,N_4223,N_4278);
and U7602 (N_7602,N_4036,N_4179);
nor U7603 (N_7603,N_4586,N_4795);
nand U7604 (N_7604,N_5690,N_4357);
xor U7605 (N_7605,N_4393,N_5260);
nand U7606 (N_7606,N_5552,N_4201);
nor U7607 (N_7607,N_4408,N_5640);
and U7608 (N_7608,N_5545,N_4344);
nor U7609 (N_7609,N_5938,N_4675);
nor U7610 (N_7610,N_4557,N_4672);
and U7611 (N_7611,N_5619,N_4396);
and U7612 (N_7612,N_4042,N_4246);
or U7613 (N_7613,N_4782,N_4795);
xnor U7614 (N_7614,N_4757,N_5365);
or U7615 (N_7615,N_4109,N_4260);
or U7616 (N_7616,N_4468,N_4278);
or U7617 (N_7617,N_4596,N_5734);
nand U7618 (N_7618,N_4340,N_5470);
nor U7619 (N_7619,N_4373,N_5030);
or U7620 (N_7620,N_4022,N_5206);
nand U7621 (N_7621,N_5020,N_4545);
nand U7622 (N_7622,N_5476,N_4901);
nor U7623 (N_7623,N_4008,N_4324);
nand U7624 (N_7624,N_4865,N_4752);
or U7625 (N_7625,N_5905,N_5899);
and U7626 (N_7626,N_4278,N_5503);
nor U7627 (N_7627,N_4025,N_4465);
nand U7628 (N_7628,N_4511,N_5780);
nand U7629 (N_7629,N_5419,N_4763);
xor U7630 (N_7630,N_5305,N_5399);
nor U7631 (N_7631,N_4850,N_4035);
and U7632 (N_7632,N_4749,N_5092);
xor U7633 (N_7633,N_4327,N_5294);
or U7634 (N_7634,N_5856,N_4760);
nand U7635 (N_7635,N_4745,N_4392);
nor U7636 (N_7636,N_4937,N_5211);
nor U7637 (N_7637,N_4778,N_5718);
or U7638 (N_7638,N_5646,N_4194);
or U7639 (N_7639,N_5181,N_5891);
or U7640 (N_7640,N_5430,N_5171);
nor U7641 (N_7641,N_5208,N_5065);
and U7642 (N_7642,N_4525,N_5838);
and U7643 (N_7643,N_4500,N_4363);
or U7644 (N_7644,N_4403,N_5845);
nor U7645 (N_7645,N_5621,N_4119);
and U7646 (N_7646,N_4371,N_5945);
or U7647 (N_7647,N_5651,N_5837);
nand U7648 (N_7648,N_4923,N_4016);
and U7649 (N_7649,N_4411,N_4055);
xor U7650 (N_7650,N_4100,N_5551);
nand U7651 (N_7651,N_4647,N_5276);
nor U7652 (N_7652,N_4824,N_4681);
and U7653 (N_7653,N_4620,N_5561);
nor U7654 (N_7654,N_4447,N_5217);
nand U7655 (N_7655,N_4147,N_5690);
nor U7656 (N_7656,N_4871,N_5491);
nand U7657 (N_7657,N_4498,N_5302);
and U7658 (N_7658,N_4807,N_4442);
and U7659 (N_7659,N_5237,N_5624);
nand U7660 (N_7660,N_4923,N_5036);
nor U7661 (N_7661,N_4604,N_5584);
and U7662 (N_7662,N_5634,N_5843);
and U7663 (N_7663,N_4422,N_4868);
and U7664 (N_7664,N_4923,N_5851);
or U7665 (N_7665,N_4217,N_4260);
and U7666 (N_7666,N_5287,N_4144);
and U7667 (N_7667,N_4417,N_5092);
nand U7668 (N_7668,N_4356,N_4468);
nand U7669 (N_7669,N_5753,N_4973);
or U7670 (N_7670,N_4026,N_5402);
nand U7671 (N_7671,N_4090,N_5152);
xnor U7672 (N_7672,N_4719,N_4303);
nand U7673 (N_7673,N_4097,N_4859);
or U7674 (N_7674,N_5813,N_4898);
nand U7675 (N_7675,N_5341,N_4903);
or U7676 (N_7676,N_4378,N_5471);
and U7677 (N_7677,N_4084,N_5303);
nor U7678 (N_7678,N_5763,N_5591);
and U7679 (N_7679,N_4880,N_4339);
nand U7680 (N_7680,N_4668,N_5078);
and U7681 (N_7681,N_4330,N_4666);
nor U7682 (N_7682,N_4181,N_4906);
xor U7683 (N_7683,N_4727,N_4308);
or U7684 (N_7684,N_5318,N_4172);
nand U7685 (N_7685,N_5380,N_5771);
or U7686 (N_7686,N_4305,N_4988);
nor U7687 (N_7687,N_5230,N_5564);
or U7688 (N_7688,N_4298,N_5576);
nand U7689 (N_7689,N_5505,N_5120);
and U7690 (N_7690,N_4431,N_4137);
nand U7691 (N_7691,N_4303,N_5864);
nand U7692 (N_7692,N_5337,N_4578);
and U7693 (N_7693,N_4579,N_5426);
nor U7694 (N_7694,N_5684,N_4652);
nand U7695 (N_7695,N_4786,N_4564);
or U7696 (N_7696,N_5754,N_5056);
or U7697 (N_7697,N_4732,N_5757);
xor U7698 (N_7698,N_5773,N_4524);
and U7699 (N_7699,N_4077,N_4530);
nand U7700 (N_7700,N_4500,N_5753);
nand U7701 (N_7701,N_5220,N_5607);
or U7702 (N_7702,N_4143,N_4498);
or U7703 (N_7703,N_4901,N_4859);
or U7704 (N_7704,N_4951,N_4960);
and U7705 (N_7705,N_5885,N_5370);
nor U7706 (N_7706,N_4200,N_5823);
nor U7707 (N_7707,N_4988,N_4143);
nor U7708 (N_7708,N_5084,N_4000);
nor U7709 (N_7709,N_4689,N_4418);
or U7710 (N_7710,N_5256,N_5545);
nand U7711 (N_7711,N_5330,N_5326);
or U7712 (N_7712,N_5234,N_4385);
and U7713 (N_7713,N_5795,N_4017);
nand U7714 (N_7714,N_5617,N_4983);
or U7715 (N_7715,N_4737,N_4105);
and U7716 (N_7716,N_5963,N_4953);
or U7717 (N_7717,N_4692,N_4897);
nand U7718 (N_7718,N_4623,N_4597);
or U7719 (N_7719,N_4027,N_5952);
nand U7720 (N_7720,N_5365,N_5139);
nor U7721 (N_7721,N_5431,N_4884);
and U7722 (N_7722,N_5729,N_5463);
or U7723 (N_7723,N_5673,N_5481);
nor U7724 (N_7724,N_4914,N_4737);
nand U7725 (N_7725,N_5704,N_5859);
or U7726 (N_7726,N_4246,N_5032);
and U7727 (N_7727,N_4417,N_5723);
and U7728 (N_7728,N_5778,N_4642);
and U7729 (N_7729,N_5381,N_5222);
and U7730 (N_7730,N_4943,N_5648);
nor U7731 (N_7731,N_4978,N_4028);
nand U7732 (N_7732,N_4996,N_4397);
nor U7733 (N_7733,N_4953,N_5974);
and U7734 (N_7734,N_5044,N_5344);
nor U7735 (N_7735,N_4447,N_5159);
and U7736 (N_7736,N_5002,N_4193);
and U7737 (N_7737,N_5311,N_4812);
nand U7738 (N_7738,N_5366,N_5962);
or U7739 (N_7739,N_5413,N_4291);
and U7740 (N_7740,N_4768,N_5819);
and U7741 (N_7741,N_5109,N_4009);
nor U7742 (N_7742,N_5283,N_5819);
and U7743 (N_7743,N_5450,N_4562);
or U7744 (N_7744,N_4411,N_5299);
or U7745 (N_7745,N_4452,N_4751);
or U7746 (N_7746,N_4593,N_4118);
and U7747 (N_7747,N_4822,N_4737);
and U7748 (N_7748,N_5352,N_4254);
nor U7749 (N_7749,N_5158,N_5167);
or U7750 (N_7750,N_5648,N_4148);
and U7751 (N_7751,N_4741,N_5861);
or U7752 (N_7752,N_4831,N_5654);
nand U7753 (N_7753,N_4816,N_5216);
nor U7754 (N_7754,N_5425,N_4925);
and U7755 (N_7755,N_5070,N_4899);
nand U7756 (N_7756,N_5603,N_5885);
nand U7757 (N_7757,N_5210,N_4218);
nor U7758 (N_7758,N_5423,N_4317);
nand U7759 (N_7759,N_4692,N_5899);
and U7760 (N_7760,N_5775,N_5114);
and U7761 (N_7761,N_5267,N_4424);
or U7762 (N_7762,N_4248,N_4400);
nand U7763 (N_7763,N_4788,N_4204);
or U7764 (N_7764,N_5755,N_4451);
or U7765 (N_7765,N_5806,N_4186);
nor U7766 (N_7766,N_5419,N_5673);
xnor U7767 (N_7767,N_4602,N_5668);
xnor U7768 (N_7768,N_5564,N_5106);
nor U7769 (N_7769,N_5511,N_5716);
or U7770 (N_7770,N_5917,N_4577);
or U7771 (N_7771,N_5138,N_5126);
or U7772 (N_7772,N_4692,N_4804);
xnor U7773 (N_7773,N_5348,N_5255);
nand U7774 (N_7774,N_5444,N_4590);
and U7775 (N_7775,N_5538,N_5369);
xnor U7776 (N_7776,N_4110,N_5508);
or U7777 (N_7777,N_5474,N_5574);
and U7778 (N_7778,N_4349,N_5530);
nor U7779 (N_7779,N_5363,N_4736);
or U7780 (N_7780,N_4102,N_5613);
xnor U7781 (N_7781,N_4424,N_4849);
xor U7782 (N_7782,N_5285,N_4882);
xor U7783 (N_7783,N_4716,N_5425);
and U7784 (N_7784,N_4323,N_5404);
and U7785 (N_7785,N_5410,N_5571);
and U7786 (N_7786,N_4322,N_4328);
nor U7787 (N_7787,N_4875,N_5485);
nand U7788 (N_7788,N_5930,N_4647);
and U7789 (N_7789,N_5138,N_5630);
nor U7790 (N_7790,N_4506,N_5619);
nor U7791 (N_7791,N_5845,N_4428);
xnor U7792 (N_7792,N_5690,N_5543);
and U7793 (N_7793,N_5326,N_4468);
nand U7794 (N_7794,N_5534,N_4364);
or U7795 (N_7795,N_5807,N_5877);
or U7796 (N_7796,N_4723,N_5583);
nor U7797 (N_7797,N_5818,N_4708);
or U7798 (N_7798,N_4016,N_5991);
nor U7799 (N_7799,N_5953,N_4150);
nand U7800 (N_7800,N_5644,N_4232);
xnor U7801 (N_7801,N_5662,N_5991);
or U7802 (N_7802,N_5041,N_4414);
nor U7803 (N_7803,N_4641,N_4865);
nor U7804 (N_7804,N_4602,N_5119);
or U7805 (N_7805,N_5400,N_4847);
or U7806 (N_7806,N_5542,N_5191);
or U7807 (N_7807,N_5119,N_5761);
and U7808 (N_7808,N_4390,N_4202);
nand U7809 (N_7809,N_5618,N_5908);
and U7810 (N_7810,N_4274,N_4589);
and U7811 (N_7811,N_5015,N_4734);
or U7812 (N_7812,N_4051,N_5980);
and U7813 (N_7813,N_5236,N_4734);
nand U7814 (N_7814,N_4094,N_5151);
or U7815 (N_7815,N_4111,N_4467);
or U7816 (N_7816,N_5205,N_5533);
and U7817 (N_7817,N_5915,N_5708);
nor U7818 (N_7818,N_4878,N_4693);
or U7819 (N_7819,N_4782,N_5328);
nor U7820 (N_7820,N_4590,N_4189);
or U7821 (N_7821,N_4259,N_5681);
nand U7822 (N_7822,N_5525,N_5040);
and U7823 (N_7823,N_4098,N_5308);
nand U7824 (N_7824,N_5330,N_4048);
and U7825 (N_7825,N_4765,N_5252);
nand U7826 (N_7826,N_5103,N_4083);
nor U7827 (N_7827,N_4639,N_4387);
or U7828 (N_7828,N_4433,N_5918);
and U7829 (N_7829,N_5716,N_5971);
nor U7830 (N_7830,N_4122,N_5485);
and U7831 (N_7831,N_5612,N_5527);
nand U7832 (N_7832,N_5756,N_4911);
or U7833 (N_7833,N_4787,N_4147);
nor U7834 (N_7834,N_5688,N_5784);
nor U7835 (N_7835,N_5738,N_4616);
nor U7836 (N_7836,N_5284,N_5210);
nor U7837 (N_7837,N_4014,N_4855);
xnor U7838 (N_7838,N_5236,N_5067);
nand U7839 (N_7839,N_5589,N_5702);
nand U7840 (N_7840,N_4219,N_4087);
and U7841 (N_7841,N_4121,N_4200);
nand U7842 (N_7842,N_5597,N_4009);
nor U7843 (N_7843,N_5364,N_5739);
nand U7844 (N_7844,N_4812,N_5383);
or U7845 (N_7845,N_4146,N_5598);
or U7846 (N_7846,N_4184,N_4231);
nand U7847 (N_7847,N_5386,N_4650);
nor U7848 (N_7848,N_4428,N_5926);
or U7849 (N_7849,N_5473,N_5245);
nor U7850 (N_7850,N_4036,N_5413);
nand U7851 (N_7851,N_4921,N_4912);
nor U7852 (N_7852,N_5050,N_4718);
nand U7853 (N_7853,N_4590,N_4807);
nor U7854 (N_7854,N_4268,N_5192);
or U7855 (N_7855,N_5169,N_4248);
nand U7856 (N_7856,N_4707,N_5053);
and U7857 (N_7857,N_5016,N_5192);
nand U7858 (N_7858,N_4423,N_4696);
nor U7859 (N_7859,N_5802,N_4875);
nand U7860 (N_7860,N_5584,N_5573);
xnor U7861 (N_7861,N_5395,N_5806);
or U7862 (N_7862,N_4829,N_5339);
and U7863 (N_7863,N_5038,N_5016);
or U7864 (N_7864,N_4452,N_5700);
nor U7865 (N_7865,N_5329,N_4585);
nand U7866 (N_7866,N_4905,N_5338);
nor U7867 (N_7867,N_4094,N_4890);
and U7868 (N_7868,N_4361,N_5547);
or U7869 (N_7869,N_5952,N_4574);
nor U7870 (N_7870,N_5291,N_5518);
nor U7871 (N_7871,N_4265,N_5286);
and U7872 (N_7872,N_5743,N_5362);
or U7873 (N_7873,N_5939,N_5169);
or U7874 (N_7874,N_4946,N_4324);
and U7875 (N_7875,N_4004,N_5842);
nor U7876 (N_7876,N_4699,N_5535);
nor U7877 (N_7877,N_5185,N_4257);
and U7878 (N_7878,N_4626,N_5672);
or U7879 (N_7879,N_5982,N_4556);
nand U7880 (N_7880,N_4315,N_4359);
nor U7881 (N_7881,N_4374,N_5181);
and U7882 (N_7882,N_5469,N_5467);
and U7883 (N_7883,N_4765,N_4245);
nand U7884 (N_7884,N_4943,N_4380);
xor U7885 (N_7885,N_5855,N_5284);
nand U7886 (N_7886,N_4524,N_5123);
nand U7887 (N_7887,N_4556,N_5857);
and U7888 (N_7888,N_4429,N_5078);
nor U7889 (N_7889,N_4433,N_5228);
nor U7890 (N_7890,N_4968,N_4882);
or U7891 (N_7891,N_4430,N_5572);
nand U7892 (N_7892,N_5312,N_5221);
nand U7893 (N_7893,N_5445,N_5873);
nor U7894 (N_7894,N_4427,N_5092);
and U7895 (N_7895,N_5277,N_4267);
and U7896 (N_7896,N_5540,N_5148);
or U7897 (N_7897,N_5596,N_5940);
nor U7898 (N_7898,N_4320,N_4414);
and U7899 (N_7899,N_4242,N_4954);
nand U7900 (N_7900,N_4161,N_5748);
xor U7901 (N_7901,N_5871,N_4563);
or U7902 (N_7902,N_4173,N_5795);
or U7903 (N_7903,N_4663,N_4234);
xor U7904 (N_7904,N_4281,N_4576);
and U7905 (N_7905,N_4664,N_4656);
or U7906 (N_7906,N_4873,N_5707);
and U7907 (N_7907,N_5570,N_4029);
xnor U7908 (N_7908,N_4953,N_4027);
or U7909 (N_7909,N_5072,N_4980);
nand U7910 (N_7910,N_4856,N_4192);
or U7911 (N_7911,N_4436,N_4777);
xnor U7912 (N_7912,N_5650,N_4445);
or U7913 (N_7913,N_5500,N_5039);
nand U7914 (N_7914,N_5706,N_4740);
nand U7915 (N_7915,N_4174,N_4284);
and U7916 (N_7916,N_4746,N_5243);
and U7917 (N_7917,N_5279,N_5509);
xnor U7918 (N_7918,N_4256,N_4281);
xnor U7919 (N_7919,N_4361,N_5529);
or U7920 (N_7920,N_4154,N_4450);
nand U7921 (N_7921,N_4583,N_4498);
or U7922 (N_7922,N_4343,N_4246);
or U7923 (N_7923,N_5727,N_4216);
xnor U7924 (N_7924,N_4759,N_4063);
nand U7925 (N_7925,N_4382,N_5915);
and U7926 (N_7926,N_4410,N_4980);
or U7927 (N_7927,N_5497,N_5730);
or U7928 (N_7928,N_4751,N_5809);
nand U7929 (N_7929,N_5438,N_4069);
and U7930 (N_7930,N_4405,N_5978);
or U7931 (N_7931,N_4730,N_5535);
or U7932 (N_7932,N_4560,N_4461);
nand U7933 (N_7933,N_5330,N_5777);
nor U7934 (N_7934,N_5325,N_4780);
nor U7935 (N_7935,N_4413,N_4283);
and U7936 (N_7936,N_4239,N_4347);
nor U7937 (N_7937,N_5092,N_4454);
or U7938 (N_7938,N_5542,N_4160);
nand U7939 (N_7939,N_5004,N_4064);
nand U7940 (N_7940,N_4097,N_5010);
nand U7941 (N_7941,N_5184,N_5606);
nand U7942 (N_7942,N_4709,N_5873);
nand U7943 (N_7943,N_5773,N_4699);
nor U7944 (N_7944,N_5623,N_5205);
or U7945 (N_7945,N_5141,N_4045);
nor U7946 (N_7946,N_4020,N_4285);
nor U7947 (N_7947,N_4487,N_4968);
and U7948 (N_7948,N_4391,N_4830);
nor U7949 (N_7949,N_5916,N_4386);
nand U7950 (N_7950,N_5670,N_4817);
and U7951 (N_7951,N_4367,N_4258);
and U7952 (N_7952,N_4644,N_4555);
or U7953 (N_7953,N_4660,N_4995);
nor U7954 (N_7954,N_5003,N_4409);
and U7955 (N_7955,N_4176,N_4732);
or U7956 (N_7956,N_5325,N_4677);
or U7957 (N_7957,N_4870,N_4831);
or U7958 (N_7958,N_5582,N_4808);
xnor U7959 (N_7959,N_5250,N_5854);
nor U7960 (N_7960,N_4688,N_4987);
and U7961 (N_7961,N_5103,N_5703);
nand U7962 (N_7962,N_5699,N_4180);
nand U7963 (N_7963,N_4612,N_4778);
nor U7964 (N_7964,N_4264,N_5964);
and U7965 (N_7965,N_5620,N_4916);
xnor U7966 (N_7966,N_4381,N_4344);
nand U7967 (N_7967,N_4508,N_5177);
nand U7968 (N_7968,N_4796,N_5885);
nand U7969 (N_7969,N_4902,N_5315);
or U7970 (N_7970,N_5451,N_5616);
nor U7971 (N_7971,N_4276,N_5203);
and U7972 (N_7972,N_4614,N_5057);
nand U7973 (N_7973,N_4209,N_5104);
nand U7974 (N_7974,N_5715,N_5806);
and U7975 (N_7975,N_5673,N_5403);
nand U7976 (N_7976,N_5386,N_4189);
or U7977 (N_7977,N_4246,N_5484);
nand U7978 (N_7978,N_4240,N_5390);
nor U7979 (N_7979,N_4758,N_5498);
xor U7980 (N_7980,N_4917,N_5230);
and U7981 (N_7981,N_4987,N_5089);
and U7982 (N_7982,N_5568,N_5761);
nor U7983 (N_7983,N_5299,N_5482);
nor U7984 (N_7984,N_5067,N_4548);
nor U7985 (N_7985,N_4155,N_4370);
nand U7986 (N_7986,N_5221,N_4430);
or U7987 (N_7987,N_4033,N_4594);
nor U7988 (N_7988,N_4239,N_5467);
or U7989 (N_7989,N_4043,N_5050);
and U7990 (N_7990,N_5913,N_5793);
or U7991 (N_7991,N_4857,N_5783);
nor U7992 (N_7992,N_4506,N_5373);
xnor U7993 (N_7993,N_4586,N_5964);
and U7994 (N_7994,N_5814,N_4360);
nor U7995 (N_7995,N_5459,N_5069);
or U7996 (N_7996,N_5970,N_5202);
nand U7997 (N_7997,N_5975,N_4758);
xnor U7998 (N_7998,N_4348,N_5732);
nand U7999 (N_7999,N_5877,N_5929);
or U8000 (N_8000,N_6396,N_6691);
nor U8001 (N_8001,N_6677,N_6259);
nand U8002 (N_8002,N_7005,N_7630);
xor U8003 (N_8003,N_7912,N_7326);
nor U8004 (N_8004,N_7610,N_7175);
or U8005 (N_8005,N_7628,N_6348);
xnor U8006 (N_8006,N_7584,N_7523);
or U8007 (N_8007,N_6265,N_7657);
and U8008 (N_8008,N_6084,N_6172);
or U8009 (N_8009,N_7289,N_6080);
or U8010 (N_8010,N_7881,N_7679);
nor U8011 (N_8011,N_6254,N_6641);
nand U8012 (N_8012,N_7270,N_7436);
and U8013 (N_8013,N_7901,N_7578);
nand U8014 (N_8014,N_7233,N_7871);
or U8015 (N_8015,N_6483,N_6945);
nand U8016 (N_8016,N_7329,N_7051);
or U8017 (N_8017,N_6815,N_7660);
and U8018 (N_8018,N_6278,N_7538);
or U8019 (N_8019,N_7713,N_7036);
nand U8020 (N_8020,N_7876,N_7279);
and U8021 (N_8021,N_6380,N_6968);
nor U8022 (N_8022,N_7533,N_7104);
and U8023 (N_8023,N_6471,N_7405);
or U8024 (N_8024,N_6406,N_7656);
nand U8025 (N_8025,N_6123,N_7129);
xnor U8026 (N_8026,N_6447,N_7819);
or U8027 (N_8027,N_7797,N_6714);
nand U8028 (N_8028,N_6159,N_6725);
nor U8029 (N_8029,N_6438,N_7247);
and U8030 (N_8030,N_7798,N_7304);
and U8031 (N_8031,N_7984,N_6391);
xor U8032 (N_8032,N_6863,N_7286);
nand U8033 (N_8033,N_6059,N_6279);
nand U8034 (N_8034,N_6314,N_6659);
and U8035 (N_8035,N_6931,N_6713);
xnor U8036 (N_8036,N_7025,N_7413);
nand U8037 (N_8037,N_7559,N_7121);
or U8038 (N_8038,N_7892,N_7761);
and U8039 (N_8039,N_7554,N_6621);
nor U8040 (N_8040,N_6056,N_6051);
and U8041 (N_8041,N_6989,N_6466);
nand U8042 (N_8042,N_6851,N_6501);
nor U8043 (N_8043,N_7226,N_7781);
nor U8044 (N_8044,N_7064,N_7898);
xnor U8045 (N_8045,N_6162,N_6457);
and U8046 (N_8046,N_7222,N_6246);
nor U8047 (N_8047,N_7654,N_6431);
nand U8048 (N_8048,N_7182,N_6075);
and U8049 (N_8049,N_7084,N_6193);
or U8050 (N_8050,N_7626,N_6735);
and U8051 (N_8051,N_7072,N_6412);
or U8052 (N_8052,N_6083,N_7731);
xnor U8053 (N_8053,N_6502,N_6491);
and U8054 (N_8054,N_7812,N_7935);
nand U8055 (N_8055,N_7725,N_6780);
nand U8056 (N_8056,N_6065,N_7522);
nand U8057 (N_8057,N_6010,N_6346);
nand U8058 (N_8058,N_6847,N_7149);
nand U8059 (N_8059,N_7685,N_6373);
and U8060 (N_8060,N_6036,N_6333);
nor U8061 (N_8061,N_7347,N_7108);
and U8062 (N_8062,N_7494,N_6188);
nand U8063 (N_8063,N_6411,N_7774);
or U8064 (N_8064,N_6577,N_7002);
or U8065 (N_8065,N_7934,N_7927);
and U8066 (N_8066,N_6213,N_6181);
or U8067 (N_8067,N_6536,N_6828);
and U8068 (N_8068,N_7560,N_7942);
nand U8069 (N_8069,N_6048,N_7066);
nand U8070 (N_8070,N_7524,N_7189);
nand U8071 (N_8071,N_7441,N_6323);
xor U8072 (N_8072,N_6381,N_6088);
or U8073 (N_8073,N_6636,N_6848);
xor U8074 (N_8074,N_7545,N_6628);
nand U8075 (N_8075,N_6787,N_6681);
xor U8076 (N_8076,N_7874,N_6670);
or U8077 (N_8077,N_7506,N_7128);
xor U8078 (N_8078,N_7343,N_6860);
and U8079 (N_8079,N_7011,N_6873);
or U8080 (N_8080,N_7454,N_6512);
xnor U8081 (N_8081,N_7255,N_7750);
or U8082 (N_8082,N_6124,N_7899);
nor U8083 (N_8083,N_6493,N_6427);
and U8084 (N_8084,N_7396,N_7817);
xor U8085 (N_8085,N_7473,N_7437);
nand U8086 (N_8086,N_7088,N_6710);
nor U8087 (N_8087,N_7359,N_6876);
xor U8088 (N_8088,N_6850,N_7786);
nor U8089 (N_8089,N_7049,N_6097);
and U8090 (N_8090,N_6767,N_7106);
and U8091 (N_8091,N_6557,N_7069);
and U8092 (N_8092,N_7729,N_6095);
nand U8093 (N_8093,N_7944,N_6023);
xor U8094 (N_8094,N_7068,N_6370);
nand U8095 (N_8095,N_7196,N_6376);
nand U8096 (N_8096,N_6114,N_6955);
or U8097 (N_8097,N_7958,N_7278);
or U8098 (N_8098,N_6569,N_7421);
or U8099 (N_8099,N_6631,N_7294);
and U8100 (N_8100,N_7062,N_7264);
and U8101 (N_8101,N_6375,N_7404);
xnor U8102 (N_8102,N_7290,N_6413);
or U8103 (N_8103,N_6961,N_6591);
or U8104 (N_8104,N_6629,N_6035);
or U8105 (N_8105,N_7198,N_6802);
and U8106 (N_8106,N_7316,N_6118);
xnor U8107 (N_8107,N_6086,N_7397);
or U8108 (N_8108,N_7184,N_7586);
nor U8109 (N_8109,N_6490,N_6495);
nor U8110 (N_8110,N_7737,N_7311);
or U8111 (N_8111,N_7361,N_7742);
and U8112 (N_8112,N_7579,N_6775);
nor U8113 (N_8113,N_7868,N_6230);
nor U8114 (N_8114,N_6378,N_6073);
nand U8115 (N_8115,N_6592,N_7360);
nand U8116 (N_8116,N_7331,N_7831);
and U8117 (N_8117,N_6997,N_6357);
xor U8118 (N_8118,N_7859,N_7720);
nand U8119 (N_8119,N_7583,N_7776);
xor U8120 (N_8120,N_7612,N_7996);
nor U8121 (N_8121,N_6737,N_6524);
and U8122 (N_8122,N_7145,N_7034);
and U8123 (N_8123,N_6999,N_6527);
xnor U8124 (N_8124,N_6004,N_7282);
or U8125 (N_8125,N_7305,N_7668);
or U8126 (N_8126,N_7711,N_6607);
and U8127 (N_8127,N_6277,N_7947);
nand U8128 (N_8128,N_6212,N_6907);
or U8129 (N_8129,N_6283,N_6105);
and U8130 (N_8130,N_6757,N_6831);
nor U8131 (N_8131,N_6773,N_6935);
nor U8132 (N_8132,N_7704,N_6587);
or U8133 (N_8133,N_6068,N_7672);
and U8134 (N_8134,N_6470,N_6429);
or U8135 (N_8135,N_7215,N_7123);
nor U8136 (N_8136,N_6801,N_7461);
xnor U8137 (N_8137,N_6559,N_7120);
nor U8138 (N_8138,N_6957,N_6407);
nor U8139 (N_8139,N_6194,N_6546);
nand U8140 (N_8140,N_7219,N_7362);
or U8141 (N_8141,N_6861,N_7318);
nand U8142 (N_8142,N_6783,N_6732);
and U8143 (N_8143,N_7336,N_7867);
xnor U8144 (N_8144,N_7667,N_7611);
xor U8145 (N_8145,N_6899,N_6892);
nor U8146 (N_8146,N_6533,N_7843);
nor U8147 (N_8147,N_7730,N_6488);
nand U8148 (N_8148,N_7161,N_6285);
xnor U8149 (N_8149,N_6603,N_7211);
and U8150 (N_8150,N_6541,N_7171);
and U8151 (N_8151,N_7585,N_7683);
xnor U8152 (N_8152,N_7665,N_7257);
or U8153 (N_8153,N_6077,N_6155);
or U8154 (N_8154,N_6044,N_6358);
xor U8155 (N_8155,N_7450,N_7692);
nor U8156 (N_8156,N_6271,N_7327);
or U8157 (N_8157,N_7261,N_7357);
or U8158 (N_8158,N_7333,N_7537);
nor U8159 (N_8159,N_7113,N_6178);
and U8160 (N_8160,N_6420,N_7020);
nand U8161 (N_8161,N_7855,N_6505);
nand U8162 (N_8162,N_7079,N_7646);
and U8163 (N_8163,N_7220,N_6869);
and U8164 (N_8164,N_6748,N_6685);
xor U8165 (N_8165,N_6476,N_6335);
or U8166 (N_8166,N_7791,N_6582);
and U8167 (N_8167,N_7228,N_7075);
nand U8168 (N_8168,N_6152,N_6025);
nand U8169 (N_8169,N_7181,N_6221);
nand U8170 (N_8170,N_6418,N_7172);
nor U8171 (N_8171,N_6513,N_6539);
nand U8172 (N_8172,N_6324,N_7863);
or U8173 (N_8173,N_6870,N_7875);
and U8174 (N_8174,N_6664,N_7624);
or U8175 (N_8175,N_7705,N_6206);
or U8176 (N_8176,N_6390,N_7785);
nor U8177 (N_8177,N_6006,N_7777);
and U8178 (N_8178,N_6492,N_6844);
nand U8179 (N_8179,N_6454,N_6252);
and U8180 (N_8180,N_6614,N_6131);
nor U8181 (N_8181,N_7503,N_7806);
nand U8182 (N_8182,N_7259,N_7298);
and U8183 (N_8183,N_6126,N_6377);
nand U8184 (N_8184,N_6988,N_7778);
or U8185 (N_8185,N_6715,N_6785);
xnor U8186 (N_8186,N_7370,N_6547);
nor U8187 (N_8187,N_6833,N_6951);
nand U8188 (N_8188,N_6141,N_7904);
xor U8189 (N_8189,N_7802,N_6689);
xnor U8190 (N_8190,N_6933,N_7745);
nor U8191 (N_8191,N_6797,N_7122);
nand U8192 (N_8192,N_6623,N_6901);
xnor U8193 (N_8193,N_6594,N_7280);
or U8194 (N_8194,N_7613,N_6841);
and U8195 (N_8195,N_6584,N_7815);
or U8196 (N_8196,N_6964,N_6300);
nand U8197 (N_8197,N_7689,N_7050);
nor U8198 (N_8198,N_7492,N_6263);
and U8199 (N_8199,N_7428,N_6705);
and U8200 (N_8200,N_6813,N_7296);
xnor U8201 (N_8201,N_7495,N_7015);
xor U8202 (N_8202,N_7440,N_7137);
or U8203 (N_8203,N_7504,N_7388);
and U8204 (N_8204,N_6291,N_6630);
nor U8205 (N_8205,N_7775,N_6186);
nor U8206 (N_8206,N_7771,N_7784);
or U8207 (N_8207,N_7431,N_6102);
and U8208 (N_8208,N_6819,N_7873);
nor U8209 (N_8209,N_7239,N_7426);
and U8210 (N_8210,N_7111,N_6266);
and U8211 (N_8211,N_7835,N_6679);
and U8212 (N_8212,N_7953,N_6460);
and U8213 (N_8213,N_7682,N_6858);
and U8214 (N_8214,N_7839,N_7766);
nor U8215 (N_8215,N_6948,N_6724);
nand U8216 (N_8216,N_7144,N_7923);
nand U8217 (N_8217,N_6115,N_6020);
nor U8218 (N_8218,N_6682,N_7055);
and U8219 (N_8219,N_6824,N_6489);
nor U8220 (N_8220,N_7054,N_7498);
xor U8221 (N_8221,N_6153,N_6716);
nand U8222 (N_8222,N_7168,N_6455);
or U8223 (N_8223,N_6218,N_7012);
xor U8224 (N_8224,N_7564,N_7520);
or U8225 (N_8225,N_7256,N_6345);
nand U8226 (N_8226,N_7199,N_6538);
or U8227 (N_8227,N_7889,N_6920);
nand U8228 (N_8228,N_6777,N_6468);
nor U8229 (N_8229,N_7432,N_6647);
nor U8230 (N_8230,N_6962,N_7833);
nor U8231 (N_8231,N_7794,N_6012);
or U8232 (N_8232,N_7511,N_6168);
xnor U8233 (N_8233,N_6543,N_6560);
and U8234 (N_8234,N_7518,N_7445);
xnor U8235 (N_8235,N_6936,N_6436);
nand U8236 (N_8236,N_7139,N_7866);
nor U8237 (N_8237,N_6262,N_7986);
nand U8238 (N_8238,N_6039,N_7474);
or U8239 (N_8239,N_7519,N_7529);
nand U8240 (N_8240,N_6825,N_6956);
or U8241 (N_8241,N_6895,N_7915);
or U8242 (N_8242,N_6916,N_7017);
nand U8243 (N_8243,N_7676,N_6298);
or U8244 (N_8244,N_6751,N_7752);
and U8245 (N_8245,N_6698,N_7939);
xnor U8246 (N_8246,N_7476,N_7764);
and U8247 (N_8247,N_7805,N_6877);
nor U8248 (N_8248,N_7086,N_7083);
nand U8249 (N_8249,N_6191,N_7770);
nor U8250 (N_8250,N_7548,N_7045);
and U8251 (N_8251,N_7842,N_7526);
nand U8252 (N_8252,N_6474,N_6857);
or U8253 (N_8253,N_7427,N_7936);
nor U8254 (N_8254,N_6275,N_6202);
and U8255 (N_8255,N_6943,N_6127);
xnor U8256 (N_8256,N_7751,N_7345);
or U8257 (N_8257,N_7342,N_7118);
nor U8258 (N_8258,N_6383,N_6359);
nand U8259 (N_8259,N_7383,N_6076);
and U8260 (N_8260,N_7840,N_7291);
or U8261 (N_8261,N_6929,N_7710);
nor U8262 (N_8262,N_7973,N_6052);
and U8263 (N_8263,N_7747,N_6644);
nand U8264 (N_8264,N_7691,N_6906);
nand U8265 (N_8265,N_7739,N_7807);
or U8266 (N_8266,N_7138,N_7152);
nor U8267 (N_8267,N_7834,N_7512);
and U8268 (N_8268,N_7456,N_6885);
xor U8269 (N_8269,N_6952,N_7916);
xor U8270 (N_8270,N_7391,N_6294);
nand U8271 (N_8271,N_7622,N_7081);
and U8272 (N_8272,N_6695,N_6898);
nand U8273 (N_8273,N_7708,N_6836);
nand U8274 (N_8274,N_7767,N_7283);
nand U8275 (N_8275,N_6409,N_7063);
and U8276 (N_8276,N_7772,N_6410);
xnor U8277 (N_8277,N_7913,N_7605);
and U8278 (N_8278,N_6310,N_6722);
and U8279 (N_8279,N_7303,N_7200);
and U8280 (N_8280,N_6910,N_6484);
nor U8281 (N_8281,N_6874,N_7789);
or U8282 (N_8282,N_7489,N_7659);
and U8283 (N_8283,N_7527,N_7664);
and U8284 (N_8284,N_7557,N_7800);
and U8285 (N_8285,N_7410,N_6408);
xnor U8286 (N_8286,N_7674,N_6764);
and U8287 (N_8287,N_6752,N_7816);
nand U8288 (N_8288,N_6750,N_7678);
nand U8289 (N_8289,N_7561,N_6653);
nand U8290 (N_8290,N_6133,N_7880);
nor U8291 (N_8291,N_6026,N_7858);
nand U8292 (N_8292,N_6441,N_6486);
nand U8293 (N_8293,N_6693,N_7192);
nor U8294 (N_8294,N_7556,N_7634);
xnor U8295 (N_8295,N_7135,N_6549);
nand U8296 (N_8296,N_7543,N_6654);
or U8297 (N_8297,N_6031,N_7961);
xnor U8298 (N_8298,N_7910,N_6009);
nor U8299 (N_8299,N_6143,N_6520);
xnor U8300 (N_8300,N_6496,N_7140);
nand U8301 (N_8301,N_6237,N_6465);
nor U8302 (N_8302,N_6424,N_7043);
nor U8303 (N_8303,N_6157,N_7993);
or U8304 (N_8304,N_6482,N_6183);
and U8305 (N_8305,N_7091,N_7848);
nor U8306 (N_8306,N_7484,N_6444);
nor U8307 (N_8307,N_6276,N_6745);
and U8308 (N_8308,N_6747,N_6589);
nor U8309 (N_8309,N_7468,N_7053);
or U8310 (N_8310,N_7022,N_7723);
nor U8311 (N_8311,N_7204,N_6868);
nor U8312 (N_8312,N_6245,N_6326);
nor U8313 (N_8313,N_6992,N_6960);
nor U8314 (N_8314,N_7074,N_7938);
and U8315 (N_8315,N_6061,N_7675);
xnor U8316 (N_8316,N_6463,N_7073);
or U8317 (N_8317,N_6101,N_7216);
or U8318 (N_8318,N_6849,N_7546);
nor U8319 (N_8319,N_7508,N_7534);
and U8320 (N_8320,N_7929,N_6108);
nor U8321 (N_8321,N_6782,N_7857);
xor U8322 (N_8322,N_7600,N_6665);
nor U8323 (N_8323,N_6531,N_7575);
nor U8324 (N_8324,N_7619,N_6028);
nor U8325 (N_8325,N_6690,N_7852);
or U8326 (N_8326,N_6256,N_7918);
xor U8327 (N_8327,N_7999,N_6827);
xor U8328 (N_8328,N_6064,N_6597);
or U8329 (N_8329,N_6887,N_6417);
xnor U8330 (N_8330,N_7635,N_6545);
nand U8331 (N_8331,N_7131,N_6742);
or U8332 (N_8332,N_7272,N_6128);
and U8333 (N_8333,N_6229,N_7349);
or U8334 (N_8334,N_7603,N_6480);
nand U8335 (N_8335,N_6145,N_6288);
or U8336 (N_8336,N_6954,N_7780);
or U8337 (N_8337,N_6485,N_7317);
xor U8338 (N_8338,N_6307,N_6704);
and U8339 (N_8339,N_6744,N_7864);
xor U8340 (N_8340,N_6565,N_6268);
xnor U8341 (N_8341,N_7232,N_6674);
nor U8342 (N_8342,N_7090,N_6700);
nand U8343 (N_8343,N_6405,N_6741);
or U8344 (N_8344,N_6165,N_7760);
xor U8345 (N_8345,N_7744,N_7156);
nand U8346 (N_8346,N_6600,N_7231);
nor U8347 (N_8347,N_6553,N_6625);
nand U8348 (N_8348,N_7860,N_6329);
or U8349 (N_8349,N_7276,N_7218);
nor U8350 (N_8350,N_7130,N_7371);
nand U8351 (N_8351,N_7014,N_6890);
nand U8352 (N_8352,N_6939,N_7308);
nand U8353 (N_8353,N_6219,N_6421);
nand U8354 (N_8354,N_7267,N_6249);
nand U8355 (N_8355,N_6835,N_7110);
or U8356 (N_8356,N_6763,N_7499);
and U8357 (N_8357,N_6184,N_6313);
nand U8358 (N_8358,N_6731,N_6371);
nand U8359 (N_8359,N_7614,N_6122);
nand U8360 (N_8360,N_7067,N_7618);
and U8361 (N_8361,N_7686,N_6590);
nor U8362 (N_8362,N_7416,N_7340);
and U8363 (N_8363,N_6267,N_6286);
nand U8364 (N_8364,N_6069,N_7008);
or U8365 (N_8365,N_7191,N_7878);
and U8366 (N_8366,N_6994,N_6208);
nor U8367 (N_8367,N_6642,N_7712);
or U8368 (N_8368,N_6464,N_6511);
and U8369 (N_8369,N_7818,N_6729);
or U8370 (N_8370,N_6041,N_6216);
and U8371 (N_8371,N_7162,N_7099);
nand U8372 (N_8372,N_7722,N_7392);
nor U8373 (N_8373,N_7366,N_6834);
xnor U8374 (N_8374,N_7909,N_7102);
nor U8375 (N_8375,N_6382,N_7716);
xor U8376 (N_8376,N_7097,N_6074);
or U8377 (N_8377,N_7472,N_6712);
nor U8378 (N_8378,N_6055,N_7453);
nor U8379 (N_8379,N_6595,N_6509);
nand U8380 (N_8380,N_6399,N_7836);
nand U8381 (N_8381,N_6888,N_7030);
or U8382 (N_8382,N_7024,N_7205);
nor U8383 (N_8383,N_6297,N_6678);
xor U8384 (N_8384,N_7606,N_7862);
nand U8385 (N_8385,N_7382,N_7756);
and U8386 (N_8386,N_7568,N_7460);
or U8387 (N_8387,N_7998,N_6342);
or U8388 (N_8388,N_6226,N_6224);
and U8389 (N_8389,N_7699,N_7921);
and U8390 (N_8390,N_6034,N_7502);
xor U8391 (N_8391,N_6397,N_7743);
and U8392 (N_8392,N_7887,N_7885);
nand U8393 (N_8393,N_6503,N_6138);
nand U8394 (N_8394,N_7879,N_7922);
nor U8395 (N_8395,N_6786,N_6005);
nand U8396 (N_8396,N_6135,N_6881);
nand U8397 (N_8397,N_7669,N_7385);
nand U8398 (N_8398,N_7424,N_6561);
nand U8399 (N_8399,N_6120,N_7647);
xnor U8400 (N_8400,N_6507,N_6320);
nand U8401 (N_8401,N_6459,N_7845);
xnor U8402 (N_8402,N_6318,N_7258);
or U8403 (N_8403,N_6332,N_7244);
and U8404 (N_8404,N_6606,N_6537);
or U8405 (N_8405,N_7224,N_6884);
nor U8406 (N_8406,N_6112,N_6555);
and U8407 (N_8407,N_6164,N_6526);
nor U8408 (N_8408,N_6781,N_7027);
nand U8409 (N_8409,N_7642,N_7830);
or U8410 (N_8410,N_6601,N_6803);
nor U8411 (N_8411,N_7967,N_7414);
nand U8412 (N_8412,N_7407,N_6446);
nor U8413 (N_8413,N_7451,N_6015);
and U8414 (N_8414,N_7225,N_7697);
nor U8415 (N_8415,N_6481,N_7443);
xnor U8416 (N_8416,N_7962,N_7604);
and U8417 (N_8417,N_6598,N_6983);
or U8418 (N_8418,N_6820,N_7071);
nor U8419 (N_8419,N_6842,N_6542);
xnor U8420 (N_8420,N_6882,N_6707);
or U8421 (N_8421,N_7530,N_6806);
and U8422 (N_8422,N_6344,N_6915);
or U8423 (N_8423,N_6167,N_7643);
or U8424 (N_8424,N_7299,N_6054);
nand U8425 (N_8425,N_7467,N_6351);
and U8426 (N_8426,N_6635,N_7924);
or U8427 (N_8427,N_6209,N_7582);
or U8428 (N_8428,N_7146,N_7477);
nor U8429 (N_8429,N_7645,N_7844);
nor U8430 (N_8430,N_7240,N_7214);
nand U8431 (N_8431,N_7095,N_6917);
xnor U8432 (N_8432,N_6189,N_7640);
nand U8433 (N_8433,N_7746,N_6779);
nor U8434 (N_8434,N_7134,N_6702);
xnor U8435 (N_8435,N_7653,N_7169);
or U8436 (N_8436,N_6472,N_7908);
and U8437 (N_8437,N_6897,N_7623);
xnor U8438 (N_8438,N_6352,N_6562);
and U8439 (N_8439,N_6672,N_6984);
nor U8440 (N_8440,N_6872,N_6564);
nand U8441 (N_8441,N_7254,N_6137);
xor U8442 (N_8442,N_7930,N_7422);
or U8443 (N_8443,N_7019,N_6241);
or U8444 (N_8444,N_7763,N_7295);
and U8445 (N_8445,N_6839,N_7563);
nand U8446 (N_8446,N_6889,N_6651);
and U8447 (N_8447,N_7884,N_6771);
or U8448 (N_8448,N_6909,N_6829);
or U8449 (N_8449,N_6225,N_6364);
or U8450 (N_8450,N_6032,N_6749);
nand U8451 (N_8451,N_6422,N_6442);
xor U8452 (N_8452,N_7348,N_7985);
nand U8453 (N_8453,N_7190,N_7790);
nor U8454 (N_8454,N_7732,N_7029);
or U8455 (N_8455,N_7734,N_7933);
xor U8456 (N_8456,N_7070,N_7990);
nand U8457 (N_8457,N_6308,N_7509);
or U8458 (N_8458,N_6154,N_7052);
or U8459 (N_8459,N_6053,N_6580);
nor U8460 (N_8460,N_6106,N_7906);
or U8461 (N_8461,N_6919,N_6728);
nor U8462 (N_8462,N_6680,N_7945);
and U8463 (N_8463,N_7963,N_6477);
nand U8464 (N_8464,N_6683,N_6018);
xnor U8465 (N_8465,N_7332,N_6247);
or U8466 (N_8466,N_7116,N_7949);
or U8467 (N_8467,N_6021,N_6979);
nor U8468 (N_8468,N_7142,N_7719);
xnor U8469 (N_8469,N_6667,N_7517);
or U8470 (N_8470,N_6922,N_6067);
nand U8471 (N_8471,N_6768,N_7810);
nand U8472 (N_8472,N_6369,N_6078);
or U8473 (N_8473,N_7952,N_6305);
nor U8474 (N_8474,N_7652,N_7449);
nand U8475 (N_8475,N_7330,N_7714);
and U8476 (N_8476,N_6599,N_6449);
and U8477 (N_8477,N_6941,N_6618);
xor U8478 (N_8478,N_6739,N_6792);
nor U8479 (N_8479,N_6810,N_7609);
and U8480 (N_8480,N_6942,N_7877);
or U8481 (N_8481,N_7319,N_6287);
nor U8482 (N_8482,N_6394,N_6440);
xor U8483 (N_8483,N_7567,N_7919);
nor U8484 (N_8484,N_6826,N_6991);
or U8485 (N_8485,N_7339,N_7003);
nor U8486 (N_8486,N_6251,N_7375);
nand U8487 (N_8487,N_6604,N_7288);
nand U8488 (N_8488,N_7591,N_7576);
nand U8489 (N_8489,N_7539,N_7693);
and U8490 (N_8490,N_6518,N_6261);
nand U8491 (N_8491,N_6087,N_7894);
and U8492 (N_8492,N_6986,N_6762);
nor U8493 (N_8493,N_6990,N_7521);
or U8494 (N_8494,N_6423,N_6985);
nor U8495 (N_8495,N_6720,N_7117);
nor U8496 (N_8496,N_6953,N_6038);
or U8497 (N_8497,N_6796,N_6756);
and U8498 (N_8498,N_7033,N_6462);
nand U8499 (N_8499,N_7379,N_6458);
nand U8500 (N_8500,N_7565,N_6608);
xnor U8501 (N_8501,N_6456,N_7287);
and U8502 (N_8502,N_6214,N_7010);
and U8503 (N_8503,N_6063,N_6914);
or U8504 (N_8504,N_6347,N_7085);
nand U8505 (N_8505,N_7394,N_7320);
and U8506 (N_8506,N_6790,N_7207);
or U8507 (N_8507,N_6788,N_6554);
nor U8508 (N_8508,N_7418,N_7826);
nor U8509 (N_8509,N_7107,N_6938);
nor U8510 (N_8510,N_6203,N_7594);
and U8511 (N_8511,N_6090,N_6924);
nor U8512 (N_8512,N_6726,N_7037);
nand U8513 (N_8513,N_6119,N_7268);
nor U8514 (N_8514,N_6200,N_6932);
nor U8515 (N_8515,N_6879,N_6269);
nand U8516 (N_8516,N_7615,N_6864);
nand U8517 (N_8517,N_7026,N_7170);
nor U8518 (N_8518,N_7788,N_7013);
nand U8519 (N_8519,N_7602,N_6040);
nor U8520 (N_8520,N_7856,N_7592);
and U8521 (N_8521,N_6894,N_7266);
or U8522 (N_8522,N_6637,N_7155);
or U8523 (N_8523,N_7893,N_6156);
xnor U8524 (N_8524,N_7516,N_6544);
nor U8525 (N_8525,N_6207,N_6822);
xnor U8526 (N_8526,N_6981,N_6292);
xnor U8527 (N_8527,N_6891,N_7419);
or U8528 (N_8528,N_7854,N_6809);
nand U8529 (N_8529,N_7570,N_7827);
nand U8530 (N_8530,N_7411,N_7354);
or U8531 (N_8531,N_6150,N_7447);
nor U8532 (N_8532,N_7528,N_6199);
or U8533 (N_8533,N_7248,N_6198);
xor U8534 (N_8534,N_6387,N_7448);
nor U8535 (N_8535,N_7684,N_7060);
and U8536 (N_8536,N_7093,N_6425);
and U8537 (N_8537,N_6719,N_6563);
nor U8538 (N_8538,N_7589,N_6205);
xnor U8539 (N_8539,N_6475,N_6432);
xor U8540 (N_8540,N_7227,N_6619);
nor U8541 (N_8541,N_7183,N_6081);
or U8542 (N_8542,N_7809,N_6911);
or U8543 (N_8543,N_6615,N_6111);
or U8544 (N_8544,N_7234,N_6743);
nor U8545 (N_8545,N_6540,N_7853);
xnor U8546 (N_8546,N_7814,N_6104);
and U8547 (N_8547,N_6570,N_7946);
and U8548 (N_8548,N_7721,N_6071);
and U8549 (N_8549,N_6374,N_6516);
or U8550 (N_8550,N_7203,N_6711);
and U8551 (N_8551,N_7464,N_6772);
or U8552 (N_8552,N_6299,N_6581);
and U8553 (N_8553,N_7163,N_7458);
or U8554 (N_8554,N_7478,N_6129);
nor U8555 (N_8555,N_6646,N_6385);
and U8556 (N_8556,N_7753,N_7353);
nor U8557 (N_8557,N_6350,N_7727);
nor U8558 (N_8558,N_7356,N_7399);
and U8559 (N_8559,N_6576,N_7243);
or U8560 (N_8560,N_6272,N_6239);
nor U8561 (N_8561,N_7823,N_7847);
or U8562 (N_8562,N_7209,N_6166);
nand U8563 (N_8563,N_7542,N_7590);
nand U8564 (N_8564,N_7673,N_7625);
and U8565 (N_8565,N_7496,N_6494);
and U8566 (N_8566,N_6368,N_7651);
and U8567 (N_8567,N_7080,N_7698);
nand U8568 (N_8568,N_7793,N_7197);
nand U8569 (N_8569,N_7799,N_6403);
or U8570 (N_8570,N_6862,N_7112);
xor U8571 (N_8571,N_7896,N_6687);
or U8572 (N_8572,N_7433,N_7549);
or U8573 (N_8573,N_6567,N_6886);
and U8574 (N_8574,N_6072,N_6389);
and U8575 (N_8575,N_6854,N_6479);
nand U8576 (N_8576,N_6430,N_6322);
or U8577 (N_8577,N_7951,N_6934);
nor U8578 (N_8578,N_7820,N_6349);
nand U8579 (N_8579,N_6865,N_6024);
or U8580 (N_8580,N_6640,N_6930);
nor U8581 (N_8581,N_7147,N_6770);
xor U8582 (N_8582,N_6037,N_6656);
nor U8583 (N_8583,N_7369,N_6017);
and U8584 (N_8584,N_7882,N_6812);
and U8585 (N_8585,N_7978,N_7400);
and U8586 (N_8586,N_6660,N_6130);
and U8587 (N_8587,N_6996,N_6317);
nand U8588 (N_8588,N_7059,N_7813);
nor U8589 (N_8589,N_7639,N_6926);
or U8590 (N_8590,N_7373,N_6179);
nand U8591 (N_8591,N_6530,N_7309);
nor U8592 (N_8592,N_7804,N_6624);
or U8593 (N_8593,N_6343,N_7346);
and U8594 (N_8594,N_7595,N_6330);
nand U8595 (N_8595,N_7687,N_6296);
nor U8596 (N_8596,N_7850,N_6085);
xor U8597 (N_8597,N_6525,N_6649);
and U8598 (N_8598,N_7021,N_6033);
nor U8599 (N_8599,N_6232,N_7479);
nand U8600 (N_8600,N_7133,N_6337);
and U8601 (N_8601,N_6650,N_6627);
nor U8602 (N_8602,N_7393,N_7541);
or U8603 (N_8603,N_7486,N_6363);
and U8604 (N_8604,N_7505,N_6671);
or U8605 (N_8605,N_6395,N_7310);
or U8606 (N_8606,N_7825,N_6753);
and U8607 (N_8607,N_6908,N_7832);
and U8608 (N_8608,N_7769,N_7931);
and U8609 (N_8609,N_6875,N_7412);
or U8610 (N_8610,N_6706,N_7483);
xor U8611 (N_8611,N_7338,N_7325);
nor U8612 (N_8612,N_6686,N_7006);
and U8613 (N_8613,N_6113,N_6210);
and U8614 (N_8614,N_7562,N_7420);
nand U8615 (N_8615,N_6791,N_6027);
nand U8616 (N_8616,N_6180,N_6697);
nand U8617 (N_8617,N_7749,N_6117);
or U8618 (N_8618,N_7940,N_6304);
nor U8619 (N_8619,N_7115,N_7970);
and U8620 (N_8620,N_6784,N_6217);
nand U8621 (N_8621,N_6196,N_7395);
nor U8622 (N_8622,N_6966,N_6499);
or U8623 (N_8623,N_6883,N_6974);
nand U8624 (N_8624,N_7439,N_7637);
nor U8625 (N_8625,N_7959,N_6336);
nor U8626 (N_8626,N_6289,N_7096);
and U8627 (N_8627,N_6937,N_7408);
xnor U8628 (N_8628,N_6284,N_7446);
nor U8629 (N_8629,N_7991,N_6675);
nand U8630 (N_8630,N_7888,N_6816);
nor U8631 (N_8631,N_7350,N_7262);
nand U8632 (N_8632,N_7490,N_7700);
nand U8633 (N_8633,N_7981,N_6498);
and U8634 (N_8634,N_7300,N_7992);
and U8635 (N_8635,N_7381,N_6566);
nand U8636 (N_8636,N_6730,N_6699);
nor U8637 (N_8637,N_7551,N_7000);
or U8638 (N_8638,N_6231,N_7292);
nand U8639 (N_8639,N_7206,N_7870);
xor U8640 (N_8640,N_6185,N_7648);
xnor U8641 (N_8641,N_6794,N_7377);
or U8642 (N_8642,N_6799,N_6845);
or U8643 (N_8643,N_7217,N_6174);
xnor U8644 (N_8644,N_6522,N_6558);
nand U8645 (N_8645,N_6846,N_7457);
and U8646 (N_8646,N_6386,N_6727);
nor U8647 (N_8647,N_7903,N_6893);
nand U8648 (N_8648,N_7757,N_7358);
nand U8649 (N_8649,N_6905,N_6439);
and U8650 (N_8650,N_6978,N_6638);
or U8651 (N_8651,N_6852,N_7048);
nand U8652 (N_8652,N_6579,N_7957);
and U8653 (N_8653,N_6173,N_6837);
nand U8654 (N_8654,N_7966,N_6098);
nand U8655 (N_8655,N_6506,N_7555);
nor U8656 (N_8656,N_6633,N_6652);
or U8657 (N_8657,N_6110,N_6568);
or U8658 (N_8658,N_7795,N_7500);
nand U8659 (N_8659,N_7989,N_7928);
or U8660 (N_8660,N_7971,N_6274);
nor U8661 (N_8661,N_6946,N_7596);
and U8662 (N_8662,N_7865,N_6859);
or U8663 (N_8663,N_6645,N_7550);
or U8664 (N_8664,N_7735,N_7143);
nor U8665 (N_8665,N_7758,N_6661);
and U8666 (N_8666,N_7956,N_7726);
nor U8667 (N_8667,N_6632,N_7620);
nand U8668 (N_8668,N_6878,N_6585);
nor U8669 (N_8669,N_6057,N_7482);
nor U8670 (N_8670,N_7368,N_6774);
and U8671 (N_8671,N_7046,N_6519);
nor U8672 (N_8672,N_7434,N_6616);
and U8673 (N_8673,N_7387,N_7238);
and U8674 (N_8674,N_6993,N_7748);
and U8675 (N_8675,N_6551,N_6925);
and U8676 (N_8676,N_7352,N_6717);
nor U8677 (N_8677,N_6149,N_7250);
or U8678 (N_8678,N_7173,N_7195);
xor U8679 (N_8679,N_6900,N_6855);
nand U8680 (N_8680,N_6233,N_6808);
and U8681 (N_8681,N_7883,N_6192);
nor U8682 (N_8682,N_6282,N_6620);
nand U8683 (N_8683,N_6817,N_6746);
nor U8684 (N_8684,N_6655,N_6182);
and U8685 (N_8685,N_7680,N_6918);
or U8686 (N_8686,N_7983,N_6404);
and U8687 (N_8687,N_6461,N_6734);
xnor U8688 (N_8688,N_6045,N_6107);
nand U8689 (N_8689,N_7822,N_7302);
or U8690 (N_8690,N_6912,N_6552);
and U8691 (N_8691,N_6079,N_6610);
and U8692 (N_8692,N_6393,N_6273);
and U8693 (N_8693,N_6548,N_6987);
nor U8694 (N_8694,N_7821,N_6648);
or U8695 (N_8695,N_6612,N_6022);
nor U8696 (N_8696,N_7210,N_6708);
nand U8697 (N_8697,N_6596,N_6478);
and U8698 (N_8698,N_7872,N_7914);
and U8699 (N_8699,N_6319,N_7581);
or U8700 (N_8700,N_7125,N_6089);
xor U8701 (N_8701,N_6703,N_7403);
and U8702 (N_8702,N_6871,N_7641);
or U8703 (N_8703,N_6197,N_7633);
or U8704 (N_8704,N_6356,N_6419);
nand U8705 (N_8705,N_6016,N_7466);
and U8706 (N_8706,N_7475,N_7435);
nand U8707 (N_8707,N_7964,N_6325);
or U8708 (N_8708,N_6611,N_7265);
xor U8709 (N_8709,N_7415,N_6093);
nor U8710 (N_8710,N_6572,N_7886);
or U8711 (N_8711,N_7588,N_7185);
and U8712 (N_8712,N_6965,N_7861);
or U8713 (N_8713,N_6586,N_7186);
or U8714 (N_8714,N_7782,N_7507);
and U8715 (N_8715,N_7754,N_6658);
nor U8716 (N_8716,N_6316,N_7644);
or U8717 (N_8717,N_7313,N_6696);
or U8718 (N_8718,N_7937,N_6721);
nand U8719 (N_8719,N_6977,N_6361);
or U8720 (N_8720,N_6666,N_7608);
xor U8721 (N_8721,N_7406,N_7341);
xor U8722 (N_8722,N_6588,N_6355);
nand U8723 (N_8723,N_6913,N_7925);
or U8724 (N_8724,N_7658,N_6007);
nor U8725 (N_8725,N_7176,N_7792);
and U8726 (N_8726,N_6366,N_7480);
nor U8727 (N_8727,N_7061,N_6215);
or U8728 (N_8728,N_6709,N_6574);
nand U8729 (N_8729,N_7101,N_7573);
xnor U8730 (N_8730,N_6295,N_7773);
and U8731 (N_8731,N_6321,N_7677);
nor U8732 (N_8732,N_6223,N_6529);
nand U8733 (N_8733,N_6433,N_6657);
or U8734 (N_8734,N_6066,N_6136);
or U8735 (N_8735,N_6593,N_6800);
nand U8736 (N_8736,N_7087,N_6451);
xnor U8737 (N_8737,N_7994,N_6243);
or U8738 (N_8738,N_7389,N_7077);
and U8739 (N_8739,N_6975,N_7398);
nand U8740 (N_8740,N_6100,N_7141);
and U8741 (N_8741,N_7230,N_7188);
and U8742 (N_8742,N_7253,N_6050);
nand U8743 (N_8743,N_7334,N_7955);
and U8744 (N_8744,N_7900,N_6453);
and U8745 (N_8745,N_7969,N_7995);
or U8746 (N_8746,N_6523,N_6694);
and U8747 (N_8747,N_6807,N_7089);
nor U8748 (N_8748,N_7100,N_7158);
or U8749 (N_8749,N_6754,N_7976);
or U8750 (N_8750,N_6163,N_7553);
or U8751 (N_8751,N_7525,N_7463);
xnor U8752 (N_8752,N_7801,N_7236);
nand U8753 (N_8753,N_7044,N_6617);
or U8754 (N_8754,N_6014,N_6228);
nand U8755 (N_8755,N_6362,N_7703);
nand U8756 (N_8756,N_7661,N_7977);
and U8757 (N_8757,N_6190,N_7960);
and U8758 (N_8758,N_6970,N_7811);
or U8759 (N_8759,N_7277,N_7082);
or U8760 (N_8760,N_6995,N_6508);
or U8761 (N_8761,N_7577,N_7363);
and U8762 (N_8762,N_7510,N_7208);
nor U8763 (N_8763,N_6534,N_6450);
nand U8764 (N_8764,N_7707,N_6415);
nand U8765 (N_8765,N_6384,N_7367);
nor U8766 (N_8766,N_6392,N_7201);
nor U8767 (N_8767,N_7297,N_7593);
nand U8768 (N_8768,N_6008,N_6605);
nand U8769 (N_8769,N_7324,N_7314);
and U8770 (N_8770,N_7028,N_7696);
or U8771 (N_8771,N_7690,N_6327);
nand U8772 (N_8772,N_6103,N_7481);
nand U8773 (N_8773,N_6856,N_7762);
nand U8774 (N_8774,N_6175,N_7315);
nor U8775 (N_8775,N_6583,N_7374);
nor U8776 (N_8776,N_6398,N_7569);
nand U8777 (N_8777,N_7895,N_6903);
nand U8778 (N_8778,N_6253,N_6639);
xnor U8779 (N_8779,N_6402,N_6270);
or U8780 (N_8780,N_6281,N_7105);
nand U8781 (N_8781,N_6309,N_6904);
xnor U8782 (N_8782,N_6171,N_6235);
and U8783 (N_8783,N_6146,N_7306);
xor U8784 (N_8784,N_7617,N_7897);
nor U8785 (N_8785,N_7180,N_7702);
nor U8786 (N_8786,N_7177,N_6372);
nand U8787 (N_8787,N_6002,N_7485);
and U8788 (N_8788,N_7941,N_6998);
nor U8789 (N_8789,N_7284,N_7787);
xor U8790 (N_8790,N_7718,N_7580);
xnor U8791 (N_8791,N_7321,N_6765);
nor U8792 (N_8792,N_7902,N_7972);
nand U8793 (N_8793,N_6046,N_6980);
xnor U8794 (N_8794,N_7038,N_6921);
or U8795 (N_8795,N_6556,N_6187);
nor U8796 (N_8796,N_6177,N_7322);
or U8797 (N_8797,N_6092,N_6578);
xor U8798 (N_8798,N_6331,N_7148);
nor U8799 (N_8799,N_7597,N_6211);
or U8800 (N_8800,N_6147,N_6521);
nor U8801 (N_8801,N_6838,N_7058);
nand U8802 (N_8802,N_6096,N_6443);
or U8803 (N_8803,N_6532,N_7891);
and U8804 (N_8804,N_7547,N_6250);
xnor U8805 (N_8805,N_7057,N_7571);
nand U8806 (N_8806,N_7251,N_6947);
nor U8807 (N_8807,N_7765,N_6662);
and U8808 (N_8808,N_6766,N_7323);
and U8809 (N_8809,N_6663,N_7452);
or U8810 (N_8810,N_7783,N_6575);
nand U8811 (N_8811,N_7465,N_6244);
and U8812 (N_8812,N_7890,N_6248);
or U8813 (N_8813,N_6867,N_7462);
or U8814 (N_8814,N_7841,N_6452);
and U8815 (N_8815,N_7094,N_7378);
nor U8816 (N_8816,N_7740,N_6733);
and U8817 (N_8817,N_6435,N_7666);
nor U8818 (N_8818,N_6315,N_6795);
and U8819 (N_8819,N_7285,N_6830);
and U8820 (N_8820,N_6866,N_7598);
nand U8821 (N_8821,N_7109,N_7260);
and U8822 (N_8822,N_7047,N_7004);
and U8823 (N_8823,N_7223,N_6535);
nand U8824 (N_8824,N_7738,N_6448);
nand U8825 (N_8825,N_7023,N_7536);
nor U8826 (N_8826,N_7988,N_6227);
nor U8827 (N_8827,N_6142,N_6160);
nor U8828 (N_8828,N_7599,N_6736);
nand U8829 (N_8829,N_6379,N_7166);
xnor U8830 (N_8830,N_6338,N_7566);
and U8831 (N_8831,N_7846,N_6500);
nand U8832 (N_8832,N_6140,N_7252);
nand U8833 (N_8833,N_7979,N_7365);
xor U8834 (N_8834,N_6293,N_6738);
xnor U8835 (N_8835,N_7124,N_6613);
nand U8836 (N_8836,N_7237,N_7429);
nor U8837 (N_8837,N_6959,N_6242);
nand U8838 (N_8838,N_6445,N_7655);
and U8839 (N_8839,N_6969,N_6776);
nor U8840 (N_8840,N_7212,N_7829);
nand U8841 (N_8841,N_6684,N_7627);
and U8842 (N_8842,N_7076,N_6222);
nand U8843 (N_8843,N_7943,N_6944);
nor U8844 (N_8844,N_7213,N_6517);
nand U8845 (N_8845,N_7018,N_7009);
nor U8846 (N_8846,N_6571,N_7715);
nor U8847 (N_8847,N_7355,N_7417);
or U8848 (N_8848,N_7281,N_6125);
or U8849 (N_8849,N_6148,N_6109);
or U8850 (N_8850,N_6414,N_7098);
or U8851 (N_8851,N_7337,N_7975);
and U8852 (N_8852,N_7249,N_6718);
nor U8853 (N_8853,N_7032,N_6609);
or U8854 (N_8854,N_6778,N_7911);
nand U8855 (N_8855,N_6759,N_7344);
or U8856 (N_8856,N_7293,N_6139);
nor U8857 (N_8857,N_6676,N_6514);
or U8858 (N_8858,N_7041,N_6755);
and U8859 (N_8859,N_6688,N_7455);
nor U8860 (N_8860,N_6550,N_7263);
and U8861 (N_8861,N_7092,N_6832);
nor U8862 (N_8862,N_7997,N_6469);
and U8863 (N_8863,N_7241,N_6234);
and U8864 (N_8864,N_7269,N_6515);
xnor U8865 (N_8865,N_7056,N_6758);
or U8866 (N_8866,N_6668,N_6528);
nor U8867 (N_8867,N_7470,N_7160);
xor U8868 (N_8868,N_7167,N_6401);
nand U8869 (N_8869,N_7497,N_7741);
nand U8870 (N_8870,N_6019,N_7701);
nor U8871 (N_8871,N_7174,N_6928);
or U8872 (N_8872,N_6740,N_7671);
nor U8873 (N_8873,N_6573,N_7488);
and U8874 (N_8874,N_7649,N_7491);
nor U8875 (N_8875,N_7307,N_7535);
or U8876 (N_8876,N_7907,N_6328);
nand U8877 (N_8877,N_6302,N_6011);
nand U8878 (N_8878,N_7531,N_6013);
nor U8879 (N_8879,N_7736,N_7136);
nor U8880 (N_8880,N_7621,N_7728);
nor U8881 (N_8881,N_7335,N_7558);
or U8882 (N_8882,N_7165,N_7275);
or U8883 (N_8883,N_7636,N_7631);
and U8884 (N_8884,N_6982,N_6158);
or U8885 (N_8885,N_6264,N_7471);
nand U8886 (N_8886,N_7755,N_6257);
and U8887 (N_8887,N_7235,N_6000);
xnor U8888 (N_8888,N_7103,N_7114);
or U8889 (N_8889,N_6161,N_7917);
or U8890 (N_8890,N_6340,N_7950);
nand U8891 (N_8891,N_6761,N_6510);
and U8892 (N_8892,N_6354,N_6692);
and U8893 (N_8893,N_6967,N_6972);
and U8894 (N_8894,N_7151,N_6003);
nand U8895 (N_8895,N_6927,N_7768);
xnor U8896 (N_8896,N_6201,N_6280);
xnor U8897 (N_8897,N_7242,N_6902);
and U8898 (N_8898,N_7695,N_7065);
and U8899 (N_8899,N_6258,N_7442);
and U8900 (N_8900,N_6950,N_6255);
xor U8901 (N_8901,N_7694,N_6626);
or U8902 (N_8902,N_7587,N_7402);
nand U8903 (N_8903,N_6811,N_7572);
nor U8904 (N_8904,N_6789,N_7948);
or U8905 (N_8905,N_7153,N_6306);
or U8906 (N_8906,N_6220,N_6963);
and U8907 (N_8907,N_6497,N_7187);
nand U8908 (N_8908,N_6334,N_6769);
nand U8909 (N_8909,N_7179,N_7194);
or U8910 (N_8910,N_7031,N_7954);
nor U8911 (N_8911,N_7709,N_6805);
nand U8912 (N_8912,N_7513,N_7040);
nand U8913 (N_8913,N_6301,N_6367);
and U8914 (N_8914,N_7384,N_7968);
nor U8915 (N_8915,N_6170,N_6240);
nand U8916 (N_8916,N_7351,N_6144);
or U8917 (N_8917,N_7796,N_6821);
and U8918 (N_8918,N_6896,N_7607);
and U8919 (N_8919,N_7001,N_7688);
nor U8920 (N_8920,N_7803,N_7601);
nand U8921 (N_8921,N_7828,N_7515);
nor U8922 (N_8922,N_7552,N_7126);
nor U8923 (N_8923,N_6723,N_7401);
nand U8924 (N_8924,N_6030,N_6049);
nand U8925 (N_8925,N_6169,N_7632);
and U8926 (N_8926,N_7042,N_7271);
nor U8927 (N_8927,N_6132,N_7616);
and U8928 (N_8928,N_7982,N_6818);
and U8929 (N_8929,N_7638,N_6793);
nand U8930 (N_8930,N_6094,N_6504);
nand U8931 (N_8931,N_7459,N_6823);
nand U8932 (N_8932,N_7965,N_6043);
and U8933 (N_8933,N_6880,N_6260);
nand U8934 (N_8934,N_6853,N_6070);
and U8935 (N_8935,N_6290,N_7662);
or U8936 (N_8936,N_6643,N_6434);
or U8937 (N_8937,N_7273,N_7980);
or U8938 (N_8938,N_7670,N_6428);
nor U8939 (N_8939,N_6195,N_6365);
or U8940 (N_8940,N_7150,N_6060);
nor U8941 (N_8941,N_6238,N_6047);
and U8942 (N_8942,N_6923,N_6602);
or U8943 (N_8943,N_6236,N_6001);
and U8944 (N_8944,N_6971,N_6437);
or U8945 (N_8945,N_6976,N_7869);
or U8946 (N_8946,N_7849,N_7987);
nor U8947 (N_8947,N_7444,N_6760);
and U8948 (N_8948,N_7932,N_6949);
xnor U8949 (N_8949,N_7328,N_6940);
or U8950 (N_8950,N_7779,N_6062);
nand U8951 (N_8951,N_7127,N_6360);
nand U8952 (N_8952,N_6121,N_7409);
nand U8953 (N_8953,N_7364,N_7487);
xnor U8954 (N_8954,N_6353,N_6843);
nor U8955 (N_8955,N_7717,N_7920);
nand U8956 (N_8956,N_7650,N_6669);
nor U8957 (N_8957,N_6339,N_7724);
or U8958 (N_8958,N_7438,N_7164);
or U8959 (N_8959,N_6303,N_7838);
or U8960 (N_8960,N_7423,N_6058);
and U8961 (N_8961,N_7202,N_7430);
or U8962 (N_8962,N_7178,N_6467);
nand U8963 (N_8963,N_6426,N_6416);
and U8964 (N_8964,N_7926,N_6400);
and U8965 (N_8965,N_7245,N_7544);
nor U8966 (N_8966,N_7193,N_7246);
nand U8967 (N_8967,N_7221,N_7974);
or U8968 (N_8968,N_6091,N_7301);
nand U8969 (N_8969,N_7629,N_7157);
or U8970 (N_8970,N_6134,N_6701);
nor U8971 (N_8971,N_6082,N_7824);
or U8972 (N_8972,N_6029,N_7132);
nor U8973 (N_8973,N_6634,N_7380);
nand U8974 (N_8974,N_6840,N_6151);
or U8975 (N_8975,N_7540,N_6673);
or U8976 (N_8976,N_7501,N_7837);
nand U8977 (N_8977,N_7851,N_6814);
and U8978 (N_8978,N_6311,N_7372);
or U8979 (N_8979,N_6804,N_7007);
and U8980 (N_8980,N_6973,N_7274);
nor U8981 (N_8981,N_7733,N_7493);
nand U8982 (N_8982,N_7681,N_7016);
and U8983 (N_8983,N_7469,N_7119);
nand U8984 (N_8984,N_6042,N_6487);
and U8985 (N_8985,N_7390,N_7663);
and U8986 (N_8986,N_7078,N_6176);
xor U8987 (N_8987,N_7808,N_6116);
nand U8988 (N_8988,N_6388,N_6341);
nand U8989 (N_8989,N_7039,N_6204);
and U8990 (N_8990,N_7425,N_6798);
or U8991 (N_8991,N_7759,N_6099);
or U8992 (N_8992,N_6958,N_7229);
or U8993 (N_8993,N_7574,N_6473);
and U8994 (N_8994,N_7386,N_7159);
nand U8995 (N_8995,N_7376,N_6622);
nand U8996 (N_8996,N_7706,N_7514);
xnor U8997 (N_8997,N_6312,N_7312);
and U8998 (N_8998,N_7532,N_7154);
and U8999 (N_8999,N_7905,N_7035);
nand U9000 (N_9000,N_6181,N_7015);
nand U9001 (N_9001,N_6669,N_6569);
nand U9002 (N_9002,N_6019,N_6916);
nand U9003 (N_9003,N_7724,N_7564);
and U9004 (N_9004,N_7903,N_6172);
and U9005 (N_9005,N_6187,N_7963);
nand U9006 (N_9006,N_6726,N_6772);
xnor U9007 (N_9007,N_7201,N_6661);
xor U9008 (N_9008,N_6800,N_7453);
nor U9009 (N_9009,N_7799,N_7943);
nand U9010 (N_9010,N_7542,N_7191);
nand U9011 (N_9011,N_7773,N_6622);
or U9012 (N_9012,N_7292,N_6808);
or U9013 (N_9013,N_6897,N_7517);
xnor U9014 (N_9014,N_6993,N_6075);
nand U9015 (N_9015,N_7032,N_7837);
and U9016 (N_9016,N_7716,N_7470);
and U9017 (N_9017,N_7709,N_7276);
nor U9018 (N_9018,N_7133,N_7565);
and U9019 (N_9019,N_6059,N_7366);
and U9020 (N_9020,N_6690,N_7648);
xnor U9021 (N_9021,N_6768,N_7909);
and U9022 (N_9022,N_6874,N_6816);
nor U9023 (N_9023,N_6191,N_6566);
and U9024 (N_9024,N_7554,N_6919);
or U9025 (N_9025,N_7065,N_6113);
and U9026 (N_9026,N_6712,N_6771);
nor U9027 (N_9027,N_6585,N_6424);
nor U9028 (N_9028,N_7616,N_7769);
nand U9029 (N_9029,N_7928,N_7838);
or U9030 (N_9030,N_7021,N_6415);
nand U9031 (N_9031,N_7301,N_6630);
and U9032 (N_9032,N_7704,N_6985);
nand U9033 (N_9033,N_7530,N_7559);
nand U9034 (N_9034,N_7673,N_6861);
or U9035 (N_9035,N_7004,N_6682);
nor U9036 (N_9036,N_7579,N_7339);
nor U9037 (N_9037,N_6231,N_6713);
or U9038 (N_9038,N_6040,N_7454);
or U9039 (N_9039,N_6279,N_7007);
nor U9040 (N_9040,N_7300,N_7567);
nand U9041 (N_9041,N_6088,N_7587);
and U9042 (N_9042,N_6227,N_7101);
nor U9043 (N_9043,N_6671,N_6288);
and U9044 (N_9044,N_7547,N_7891);
nand U9045 (N_9045,N_7845,N_7156);
nand U9046 (N_9046,N_6673,N_7374);
nor U9047 (N_9047,N_6389,N_6281);
nand U9048 (N_9048,N_6227,N_7282);
nand U9049 (N_9049,N_6710,N_7236);
nand U9050 (N_9050,N_6990,N_7641);
nor U9051 (N_9051,N_6146,N_7806);
nor U9052 (N_9052,N_6840,N_6724);
and U9053 (N_9053,N_6173,N_7818);
nand U9054 (N_9054,N_6462,N_7442);
nand U9055 (N_9055,N_6998,N_7395);
or U9056 (N_9056,N_6318,N_7030);
or U9057 (N_9057,N_7303,N_6589);
or U9058 (N_9058,N_6252,N_6186);
nand U9059 (N_9059,N_6804,N_7365);
nor U9060 (N_9060,N_7758,N_7247);
and U9061 (N_9061,N_6290,N_7711);
and U9062 (N_9062,N_6951,N_7508);
nand U9063 (N_9063,N_7288,N_6667);
nand U9064 (N_9064,N_6071,N_6963);
and U9065 (N_9065,N_6269,N_7498);
nand U9066 (N_9066,N_7349,N_6782);
or U9067 (N_9067,N_7417,N_6907);
or U9068 (N_9068,N_6822,N_7017);
nand U9069 (N_9069,N_6338,N_6817);
and U9070 (N_9070,N_6972,N_6200);
nand U9071 (N_9071,N_6903,N_7660);
and U9072 (N_9072,N_7913,N_6539);
xor U9073 (N_9073,N_7762,N_6318);
nand U9074 (N_9074,N_6664,N_7835);
or U9075 (N_9075,N_6103,N_6983);
or U9076 (N_9076,N_7321,N_6827);
nor U9077 (N_9077,N_7015,N_7534);
nor U9078 (N_9078,N_6348,N_6456);
nand U9079 (N_9079,N_7451,N_7435);
and U9080 (N_9080,N_6623,N_6781);
nand U9081 (N_9081,N_6822,N_7258);
and U9082 (N_9082,N_6218,N_7062);
or U9083 (N_9083,N_7519,N_6546);
nor U9084 (N_9084,N_6245,N_7483);
nor U9085 (N_9085,N_6736,N_7138);
xor U9086 (N_9086,N_7836,N_7195);
nor U9087 (N_9087,N_6527,N_7859);
nand U9088 (N_9088,N_6096,N_7017);
xnor U9089 (N_9089,N_6050,N_6734);
nor U9090 (N_9090,N_7784,N_6022);
nor U9091 (N_9091,N_6370,N_6951);
and U9092 (N_9092,N_7579,N_7768);
nor U9093 (N_9093,N_6887,N_6223);
nand U9094 (N_9094,N_6624,N_7935);
nand U9095 (N_9095,N_7300,N_6326);
nand U9096 (N_9096,N_7901,N_6139);
and U9097 (N_9097,N_6067,N_7416);
nand U9098 (N_9098,N_7852,N_7544);
or U9099 (N_9099,N_6696,N_7979);
or U9100 (N_9100,N_6110,N_7394);
or U9101 (N_9101,N_6672,N_6065);
nor U9102 (N_9102,N_7184,N_7329);
nor U9103 (N_9103,N_6146,N_7968);
xnor U9104 (N_9104,N_7387,N_7160);
nand U9105 (N_9105,N_7950,N_6262);
and U9106 (N_9106,N_6590,N_6936);
or U9107 (N_9107,N_7479,N_7167);
and U9108 (N_9108,N_6462,N_6915);
nand U9109 (N_9109,N_6568,N_6920);
and U9110 (N_9110,N_6420,N_7001);
and U9111 (N_9111,N_6265,N_7088);
xnor U9112 (N_9112,N_6955,N_7522);
or U9113 (N_9113,N_7449,N_7698);
and U9114 (N_9114,N_7315,N_6881);
nand U9115 (N_9115,N_7054,N_7556);
nand U9116 (N_9116,N_6063,N_6655);
nand U9117 (N_9117,N_6580,N_6936);
nor U9118 (N_9118,N_7980,N_7013);
nor U9119 (N_9119,N_6418,N_6498);
nand U9120 (N_9120,N_7430,N_7024);
nand U9121 (N_9121,N_6328,N_6892);
and U9122 (N_9122,N_6530,N_7906);
xor U9123 (N_9123,N_7511,N_7662);
nor U9124 (N_9124,N_7253,N_7607);
nand U9125 (N_9125,N_7098,N_7547);
or U9126 (N_9126,N_6552,N_7542);
or U9127 (N_9127,N_6893,N_7549);
or U9128 (N_9128,N_6801,N_6931);
nand U9129 (N_9129,N_7215,N_6210);
or U9130 (N_9130,N_6509,N_6692);
and U9131 (N_9131,N_7129,N_6691);
nor U9132 (N_9132,N_7673,N_6726);
and U9133 (N_9133,N_7028,N_6366);
nand U9134 (N_9134,N_6197,N_7757);
nand U9135 (N_9135,N_6828,N_6805);
and U9136 (N_9136,N_7177,N_7134);
or U9137 (N_9137,N_6598,N_6203);
nand U9138 (N_9138,N_6902,N_7018);
and U9139 (N_9139,N_7158,N_6340);
or U9140 (N_9140,N_6092,N_6694);
or U9141 (N_9141,N_7858,N_6673);
nand U9142 (N_9142,N_7661,N_6120);
nand U9143 (N_9143,N_6116,N_6380);
nor U9144 (N_9144,N_6226,N_6644);
and U9145 (N_9145,N_6214,N_6571);
and U9146 (N_9146,N_6896,N_6580);
and U9147 (N_9147,N_7751,N_6317);
or U9148 (N_9148,N_7305,N_7958);
nand U9149 (N_9149,N_7267,N_7145);
nand U9150 (N_9150,N_6397,N_6751);
or U9151 (N_9151,N_6393,N_7559);
xor U9152 (N_9152,N_7353,N_6012);
nand U9153 (N_9153,N_7541,N_6765);
nand U9154 (N_9154,N_6022,N_7287);
or U9155 (N_9155,N_7727,N_6168);
xnor U9156 (N_9156,N_7123,N_7801);
or U9157 (N_9157,N_6131,N_7999);
and U9158 (N_9158,N_6590,N_7328);
xor U9159 (N_9159,N_7846,N_6653);
or U9160 (N_9160,N_6339,N_7068);
or U9161 (N_9161,N_7391,N_7708);
and U9162 (N_9162,N_7316,N_7486);
or U9163 (N_9163,N_6316,N_6484);
or U9164 (N_9164,N_6457,N_7989);
nand U9165 (N_9165,N_6502,N_7319);
nand U9166 (N_9166,N_7578,N_7850);
nand U9167 (N_9167,N_7373,N_6614);
or U9168 (N_9168,N_6942,N_7617);
nand U9169 (N_9169,N_7910,N_6818);
nor U9170 (N_9170,N_6365,N_7416);
or U9171 (N_9171,N_7232,N_6309);
or U9172 (N_9172,N_7271,N_7352);
or U9173 (N_9173,N_6435,N_7400);
nand U9174 (N_9174,N_6202,N_6194);
xor U9175 (N_9175,N_6122,N_6094);
or U9176 (N_9176,N_6703,N_7797);
nor U9177 (N_9177,N_6069,N_7281);
nand U9178 (N_9178,N_7808,N_6052);
nand U9179 (N_9179,N_7503,N_6058);
and U9180 (N_9180,N_7747,N_7748);
and U9181 (N_9181,N_7280,N_6265);
nand U9182 (N_9182,N_6478,N_7059);
or U9183 (N_9183,N_7074,N_7324);
or U9184 (N_9184,N_6620,N_6276);
and U9185 (N_9185,N_6461,N_7169);
or U9186 (N_9186,N_6686,N_7156);
nand U9187 (N_9187,N_6491,N_6806);
and U9188 (N_9188,N_6376,N_7124);
nand U9189 (N_9189,N_6086,N_7760);
nor U9190 (N_9190,N_6001,N_7808);
nor U9191 (N_9191,N_6420,N_6946);
and U9192 (N_9192,N_7119,N_6382);
nor U9193 (N_9193,N_7496,N_7492);
xnor U9194 (N_9194,N_6403,N_7460);
nand U9195 (N_9195,N_6451,N_6597);
nand U9196 (N_9196,N_6546,N_7894);
and U9197 (N_9197,N_7957,N_6724);
nand U9198 (N_9198,N_7239,N_7414);
and U9199 (N_9199,N_7703,N_6537);
xor U9200 (N_9200,N_7574,N_6973);
xnor U9201 (N_9201,N_6834,N_6655);
or U9202 (N_9202,N_6596,N_7198);
nor U9203 (N_9203,N_7243,N_6439);
and U9204 (N_9204,N_7359,N_6243);
and U9205 (N_9205,N_6987,N_6043);
nor U9206 (N_9206,N_7850,N_6371);
nand U9207 (N_9207,N_7963,N_7696);
nor U9208 (N_9208,N_7119,N_7383);
xor U9209 (N_9209,N_6628,N_7634);
and U9210 (N_9210,N_7172,N_7776);
or U9211 (N_9211,N_6082,N_6973);
nand U9212 (N_9212,N_6178,N_7729);
or U9213 (N_9213,N_7577,N_6587);
nand U9214 (N_9214,N_6714,N_6169);
nor U9215 (N_9215,N_7292,N_6377);
xnor U9216 (N_9216,N_6783,N_6650);
or U9217 (N_9217,N_7403,N_7257);
or U9218 (N_9218,N_7663,N_7885);
nor U9219 (N_9219,N_7470,N_7001);
and U9220 (N_9220,N_6625,N_6249);
nand U9221 (N_9221,N_7741,N_7269);
or U9222 (N_9222,N_7246,N_7419);
xnor U9223 (N_9223,N_7392,N_7126);
nor U9224 (N_9224,N_7129,N_6940);
nor U9225 (N_9225,N_7433,N_7320);
nor U9226 (N_9226,N_6484,N_6877);
or U9227 (N_9227,N_6491,N_6173);
or U9228 (N_9228,N_6062,N_7989);
and U9229 (N_9229,N_7573,N_7073);
and U9230 (N_9230,N_6651,N_6141);
nand U9231 (N_9231,N_7900,N_6529);
nand U9232 (N_9232,N_6751,N_7011);
or U9233 (N_9233,N_6458,N_7263);
xor U9234 (N_9234,N_6256,N_7364);
xnor U9235 (N_9235,N_7503,N_7446);
and U9236 (N_9236,N_7667,N_6135);
nand U9237 (N_9237,N_6944,N_7571);
or U9238 (N_9238,N_6967,N_7132);
nor U9239 (N_9239,N_7720,N_6093);
nand U9240 (N_9240,N_7696,N_7588);
xnor U9241 (N_9241,N_6001,N_7541);
nor U9242 (N_9242,N_7378,N_7782);
or U9243 (N_9243,N_7002,N_6033);
and U9244 (N_9244,N_6331,N_7744);
and U9245 (N_9245,N_7083,N_7788);
xnor U9246 (N_9246,N_6186,N_6813);
nand U9247 (N_9247,N_7218,N_7361);
or U9248 (N_9248,N_7288,N_6591);
or U9249 (N_9249,N_6974,N_6845);
or U9250 (N_9250,N_6024,N_7488);
xnor U9251 (N_9251,N_6361,N_7871);
nand U9252 (N_9252,N_7381,N_7402);
nand U9253 (N_9253,N_7857,N_7063);
xor U9254 (N_9254,N_7697,N_7383);
and U9255 (N_9255,N_7060,N_7011);
nor U9256 (N_9256,N_7513,N_6582);
nor U9257 (N_9257,N_7745,N_6884);
or U9258 (N_9258,N_7060,N_6717);
nor U9259 (N_9259,N_7302,N_6013);
or U9260 (N_9260,N_6479,N_7203);
xnor U9261 (N_9261,N_6561,N_7121);
nor U9262 (N_9262,N_7126,N_6110);
xnor U9263 (N_9263,N_6048,N_6871);
nor U9264 (N_9264,N_6570,N_6082);
nand U9265 (N_9265,N_7284,N_6413);
nand U9266 (N_9266,N_6713,N_7581);
nor U9267 (N_9267,N_6413,N_7210);
or U9268 (N_9268,N_6857,N_6498);
or U9269 (N_9269,N_6412,N_7605);
nor U9270 (N_9270,N_7326,N_6593);
xor U9271 (N_9271,N_6987,N_6185);
or U9272 (N_9272,N_7001,N_7328);
nand U9273 (N_9273,N_6426,N_7144);
or U9274 (N_9274,N_6317,N_7063);
and U9275 (N_9275,N_7971,N_6969);
nor U9276 (N_9276,N_6961,N_7731);
nor U9277 (N_9277,N_6758,N_7245);
or U9278 (N_9278,N_6469,N_6489);
nand U9279 (N_9279,N_6266,N_7358);
nor U9280 (N_9280,N_7769,N_7484);
and U9281 (N_9281,N_6503,N_6716);
nor U9282 (N_9282,N_7104,N_7505);
nor U9283 (N_9283,N_7965,N_7263);
or U9284 (N_9284,N_6835,N_7743);
and U9285 (N_9285,N_7801,N_7792);
or U9286 (N_9286,N_7871,N_7603);
and U9287 (N_9287,N_7396,N_7585);
nor U9288 (N_9288,N_6724,N_7948);
nor U9289 (N_9289,N_7166,N_7015);
xnor U9290 (N_9290,N_6987,N_6809);
nor U9291 (N_9291,N_6552,N_6762);
or U9292 (N_9292,N_7675,N_7011);
nand U9293 (N_9293,N_6726,N_6547);
xnor U9294 (N_9294,N_7810,N_6639);
nor U9295 (N_9295,N_7346,N_7056);
nand U9296 (N_9296,N_7428,N_6530);
or U9297 (N_9297,N_6300,N_7056);
and U9298 (N_9298,N_6948,N_6090);
nand U9299 (N_9299,N_7960,N_6218);
nor U9300 (N_9300,N_6426,N_7707);
and U9301 (N_9301,N_6705,N_6752);
and U9302 (N_9302,N_7746,N_6721);
nand U9303 (N_9303,N_7035,N_6737);
or U9304 (N_9304,N_7046,N_6935);
and U9305 (N_9305,N_6308,N_7746);
or U9306 (N_9306,N_6443,N_6459);
nor U9307 (N_9307,N_6666,N_7531);
nor U9308 (N_9308,N_6433,N_6305);
nand U9309 (N_9309,N_6201,N_6974);
nor U9310 (N_9310,N_7588,N_7795);
nor U9311 (N_9311,N_6104,N_7879);
nand U9312 (N_9312,N_6050,N_6800);
nand U9313 (N_9313,N_6905,N_7515);
nand U9314 (N_9314,N_7756,N_6462);
and U9315 (N_9315,N_6823,N_6786);
or U9316 (N_9316,N_6673,N_6994);
or U9317 (N_9317,N_6153,N_7220);
and U9318 (N_9318,N_6702,N_7317);
and U9319 (N_9319,N_7257,N_7906);
xor U9320 (N_9320,N_7093,N_7475);
or U9321 (N_9321,N_6501,N_7436);
or U9322 (N_9322,N_6929,N_6731);
xnor U9323 (N_9323,N_7544,N_7191);
or U9324 (N_9324,N_7348,N_6997);
or U9325 (N_9325,N_7600,N_7586);
or U9326 (N_9326,N_6518,N_6686);
or U9327 (N_9327,N_7900,N_6352);
and U9328 (N_9328,N_7933,N_7532);
or U9329 (N_9329,N_7220,N_6807);
nand U9330 (N_9330,N_7166,N_7151);
xnor U9331 (N_9331,N_7230,N_7088);
nor U9332 (N_9332,N_7977,N_7250);
nor U9333 (N_9333,N_7093,N_7087);
and U9334 (N_9334,N_6466,N_7842);
and U9335 (N_9335,N_7511,N_7167);
nor U9336 (N_9336,N_6875,N_7806);
and U9337 (N_9337,N_7610,N_6408);
and U9338 (N_9338,N_6016,N_7757);
xor U9339 (N_9339,N_6184,N_6463);
or U9340 (N_9340,N_6449,N_6805);
or U9341 (N_9341,N_7650,N_7914);
nand U9342 (N_9342,N_7944,N_7092);
nand U9343 (N_9343,N_6435,N_7311);
xor U9344 (N_9344,N_6974,N_7987);
nand U9345 (N_9345,N_7769,N_7378);
nand U9346 (N_9346,N_7769,N_6592);
nand U9347 (N_9347,N_6238,N_6789);
nor U9348 (N_9348,N_6658,N_7263);
and U9349 (N_9349,N_7446,N_7493);
or U9350 (N_9350,N_7320,N_6151);
nand U9351 (N_9351,N_6819,N_6734);
nor U9352 (N_9352,N_7740,N_7442);
nand U9353 (N_9353,N_7522,N_6748);
or U9354 (N_9354,N_6214,N_7904);
nand U9355 (N_9355,N_7380,N_6765);
and U9356 (N_9356,N_7273,N_7340);
nand U9357 (N_9357,N_7493,N_7767);
or U9358 (N_9358,N_7671,N_7584);
nor U9359 (N_9359,N_6682,N_6447);
xor U9360 (N_9360,N_7201,N_6547);
nor U9361 (N_9361,N_7533,N_6974);
or U9362 (N_9362,N_6653,N_7061);
xor U9363 (N_9363,N_7188,N_7372);
xnor U9364 (N_9364,N_6671,N_7443);
nor U9365 (N_9365,N_6584,N_6812);
and U9366 (N_9366,N_7466,N_6746);
nand U9367 (N_9367,N_7799,N_7995);
nand U9368 (N_9368,N_6693,N_7438);
and U9369 (N_9369,N_7356,N_6504);
nand U9370 (N_9370,N_7865,N_7455);
xnor U9371 (N_9371,N_7223,N_7895);
nand U9372 (N_9372,N_7771,N_6493);
or U9373 (N_9373,N_6079,N_7010);
nand U9374 (N_9374,N_6641,N_6006);
nor U9375 (N_9375,N_7197,N_7551);
or U9376 (N_9376,N_7808,N_7873);
nand U9377 (N_9377,N_6068,N_7881);
nor U9378 (N_9378,N_7027,N_6322);
nand U9379 (N_9379,N_6234,N_6859);
nand U9380 (N_9380,N_7934,N_6787);
and U9381 (N_9381,N_7787,N_6489);
or U9382 (N_9382,N_7902,N_6276);
nand U9383 (N_9383,N_6267,N_6863);
or U9384 (N_9384,N_6079,N_7286);
or U9385 (N_9385,N_6765,N_6896);
nor U9386 (N_9386,N_6176,N_7126);
or U9387 (N_9387,N_7952,N_7759);
nor U9388 (N_9388,N_6525,N_6059);
nand U9389 (N_9389,N_7717,N_6124);
and U9390 (N_9390,N_6392,N_6251);
nand U9391 (N_9391,N_6218,N_7013);
nor U9392 (N_9392,N_7680,N_7715);
or U9393 (N_9393,N_7639,N_7921);
or U9394 (N_9394,N_6668,N_6799);
and U9395 (N_9395,N_7451,N_6608);
nor U9396 (N_9396,N_7174,N_6253);
or U9397 (N_9397,N_7682,N_7976);
nand U9398 (N_9398,N_6811,N_6843);
or U9399 (N_9399,N_6796,N_7898);
nor U9400 (N_9400,N_6253,N_7916);
and U9401 (N_9401,N_7896,N_6422);
xnor U9402 (N_9402,N_7484,N_6977);
and U9403 (N_9403,N_6621,N_7190);
nor U9404 (N_9404,N_7690,N_7784);
nor U9405 (N_9405,N_6505,N_7028);
or U9406 (N_9406,N_7450,N_6564);
xnor U9407 (N_9407,N_7311,N_7406);
nor U9408 (N_9408,N_7838,N_6969);
xnor U9409 (N_9409,N_6517,N_6705);
and U9410 (N_9410,N_7301,N_6460);
or U9411 (N_9411,N_6015,N_6176);
or U9412 (N_9412,N_7295,N_7590);
nor U9413 (N_9413,N_7603,N_7956);
nor U9414 (N_9414,N_6849,N_6437);
xor U9415 (N_9415,N_6439,N_6959);
and U9416 (N_9416,N_6749,N_7158);
and U9417 (N_9417,N_7011,N_7472);
xor U9418 (N_9418,N_7380,N_6172);
nand U9419 (N_9419,N_7274,N_6714);
or U9420 (N_9420,N_7664,N_7936);
nand U9421 (N_9421,N_7814,N_7991);
nand U9422 (N_9422,N_6012,N_6601);
nand U9423 (N_9423,N_7579,N_7522);
or U9424 (N_9424,N_7989,N_7854);
nor U9425 (N_9425,N_7515,N_7023);
or U9426 (N_9426,N_7439,N_6799);
and U9427 (N_9427,N_6864,N_7782);
nand U9428 (N_9428,N_6743,N_6595);
or U9429 (N_9429,N_6012,N_6426);
nand U9430 (N_9430,N_7392,N_7078);
and U9431 (N_9431,N_7060,N_6696);
nor U9432 (N_9432,N_7477,N_7308);
and U9433 (N_9433,N_7207,N_7705);
nand U9434 (N_9434,N_7883,N_7986);
nor U9435 (N_9435,N_7503,N_7764);
or U9436 (N_9436,N_6412,N_6119);
and U9437 (N_9437,N_7163,N_7016);
nand U9438 (N_9438,N_6076,N_6299);
or U9439 (N_9439,N_6084,N_6965);
nor U9440 (N_9440,N_6699,N_6142);
or U9441 (N_9441,N_7645,N_7808);
nor U9442 (N_9442,N_7322,N_6536);
nor U9443 (N_9443,N_6122,N_7017);
nor U9444 (N_9444,N_6388,N_7951);
and U9445 (N_9445,N_6449,N_7399);
xnor U9446 (N_9446,N_7940,N_7727);
and U9447 (N_9447,N_6093,N_7789);
xnor U9448 (N_9448,N_6370,N_6205);
xnor U9449 (N_9449,N_6823,N_6282);
or U9450 (N_9450,N_7121,N_7601);
xor U9451 (N_9451,N_7885,N_7723);
and U9452 (N_9452,N_7944,N_7058);
or U9453 (N_9453,N_7089,N_6764);
xor U9454 (N_9454,N_7480,N_7715);
nand U9455 (N_9455,N_6937,N_6129);
and U9456 (N_9456,N_7603,N_7952);
and U9457 (N_9457,N_6553,N_6377);
nor U9458 (N_9458,N_6984,N_6959);
nor U9459 (N_9459,N_6900,N_7857);
or U9460 (N_9460,N_6728,N_6116);
or U9461 (N_9461,N_7608,N_6954);
xnor U9462 (N_9462,N_6346,N_7318);
and U9463 (N_9463,N_7424,N_6845);
nand U9464 (N_9464,N_6163,N_6266);
nand U9465 (N_9465,N_7266,N_7392);
or U9466 (N_9466,N_6721,N_7074);
and U9467 (N_9467,N_6530,N_6195);
or U9468 (N_9468,N_6183,N_7061);
xnor U9469 (N_9469,N_7810,N_6594);
and U9470 (N_9470,N_7285,N_7809);
nand U9471 (N_9471,N_6616,N_6487);
or U9472 (N_9472,N_7583,N_6907);
nor U9473 (N_9473,N_6135,N_6839);
nor U9474 (N_9474,N_6783,N_6466);
or U9475 (N_9475,N_6716,N_6430);
xnor U9476 (N_9476,N_7567,N_6899);
or U9477 (N_9477,N_6381,N_7652);
or U9478 (N_9478,N_6245,N_6082);
nand U9479 (N_9479,N_7315,N_7381);
xor U9480 (N_9480,N_6547,N_6062);
xor U9481 (N_9481,N_6186,N_6400);
or U9482 (N_9482,N_7192,N_7658);
or U9483 (N_9483,N_7948,N_6232);
or U9484 (N_9484,N_6413,N_7350);
nand U9485 (N_9485,N_6819,N_6709);
nor U9486 (N_9486,N_7831,N_7074);
nand U9487 (N_9487,N_6296,N_7030);
nand U9488 (N_9488,N_6518,N_6671);
and U9489 (N_9489,N_7342,N_7723);
and U9490 (N_9490,N_7918,N_7145);
nand U9491 (N_9491,N_6242,N_6158);
or U9492 (N_9492,N_6356,N_7311);
nand U9493 (N_9493,N_6541,N_7360);
or U9494 (N_9494,N_7358,N_7043);
and U9495 (N_9495,N_6958,N_6016);
or U9496 (N_9496,N_7966,N_7225);
nand U9497 (N_9497,N_7561,N_7447);
nor U9498 (N_9498,N_7136,N_7890);
or U9499 (N_9499,N_7409,N_6701);
nand U9500 (N_9500,N_7409,N_6656);
nor U9501 (N_9501,N_6495,N_6011);
nor U9502 (N_9502,N_6085,N_6008);
nor U9503 (N_9503,N_6076,N_6611);
and U9504 (N_9504,N_6775,N_6236);
nor U9505 (N_9505,N_7782,N_6499);
nor U9506 (N_9506,N_7940,N_7285);
and U9507 (N_9507,N_7948,N_7588);
or U9508 (N_9508,N_6526,N_7463);
nand U9509 (N_9509,N_7067,N_6207);
nor U9510 (N_9510,N_6962,N_7760);
xor U9511 (N_9511,N_6657,N_7043);
or U9512 (N_9512,N_6274,N_6304);
xnor U9513 (N_9513,N_7772,N_7126);
xor U9514 (N_9514,N_6252,N_7053);
xor U9515 (N_9515,N_6920,N_7552);
nand U9516 (N_9516,N_7185,N_6624);
or U9517 (N_9517,N_7028,N_6753);
nor U9518 (N_9518,N_6010,N_7551);
or U9519 (N_9519,N_7405,N_6336);
nor U9520 (N_9520,N_6164,N_7362);
nor U9521 (N_9521,N_6137,N_6978);
nand U9522 (N_9522,N_7909,N_7512);
or U9523 (N_9523,N_6738,N_7560);
and U9524 (N_9524,N_7328,N_7187);
xnor U9525 (N_9525,N_6027,N_7542);
or U9526 (N_9526,N_6092,N_6991);
nor U9527 (N_9527,N_6164,N_6131);
nand U9528 (N_9528,N_6882,N_7417);
or U9529 (N_9529,N_7761,N_7544);
and U9530 (N_9530,N_7564,N_6863);
nand U9531 (N_9531,N_7445,N_6766);
or U9532 (N_9532,N_7733,N_7128);
nand U9533 (N_9533,N_6140,N_6168);
nand U9534 (N_9534,N_7115,N_6767);
and U9535 (N_9535,N_7189,N_6172);
or U9536 (N_9536,N_7737,N_7807);
and U9537 (N_9537,N_6063,N_7861);
xnor U9538 (N_9538,N_7051,N_6906);
and U9539 (N_9539,N_6664,N_7767);
and U9540 (N_9540,N_6505,N_7752);
nor U9541 (N_9541,N_7140,N_6614);
and U9542 (N_9542,N_6269,N_6443);
nor U9543 (N_9543,N_6953,N_7865);
nor U9544 (N_9544,N_6211,N_7793);
xnor U9545 (N_9545,N_6762,N_6840);
nor U9546 (N_9546,N_6999,N_6378);
nand U9547 (N_9547,N_7918,N_6790);
nor U9548 (N_9548,N_7002,N_7542);
nor U9549 (N_9549,N_7373,N_7211);
or U9550 (N_9550,N_7711,N_7340);
nand U9551 (N_9551,N_6721,N_6416);
or U9552 (N_9552,N_7932,N_7853);
xnor U9553 (N_9553,N_6339,N_7140);
nor U9554 (N_9554,N_6232,N_7749);
nand U9555 (N_9555,N_6324,N_6192);
or U9556 (N_9556,N_7137,N_6916);
nor U9557 (N_9557,N_6961,N_7225);
nor U9558 (N_9558,N_6677,N_6453);
nand U9559 (N_9559,N_7633,N_6453);
nor U9560 (N_9560,N_6746,N_7797);
nor U9561 (N_9561,N_6205,N_6109);
nor U9562 (N_9562,N_6372,N_7638);
and U9563 (N_9563,N_6956,N_6900);
nor U9564 (N_9564,N_6910,N_7020);
or U9565 (N_9565,N_6516,N_6953);
nand U9566 (N_9566,N_6256,N_7946);
or U9567 (N_9567,N_6360,N_6544);
nor U9568 (N_9568,N_6443,N_6629);
nor U9569 (N_9569,N_6745,N_7680);
or U9570 (N_9570,N_6192,N_7557);
and U9571 (N_9571,N_6353,N_7318);
nor U9572 (N_9572,N_7693,N_7729);
nand U9573 (N_9573,N_7145,N_7249);
xnor U9574 (N_9574,N_7807,N_6602);
nand U9575 (N_9575,N_6789,N_6076);
and U9576 (N_9576,N_6171,N_6859);
nor U9577 (N_9577,N_6643,N_6085);
and U9578 (N_9578,N_7557,N_7752);
nand U9579 (N_9579,N_7322,N_6837);
and U9580 (N_9580,N_6346,N_7360);
xnor U9581 (N_9581,N_7219,N_7679);
nand U9582 (N_9582,N_7216,N_7439);
and U9583 (N_9583,N_6799,N_7388);
and U9584 (N_9584,N_6351,N_7924);
and U9585 (N_9585,N_7410,N_7045);
and U9586 (N_9586,N_6089,N_7368);
and U9587 (N_9587,N_7052,N_6478);
nand U9588 (N_9588,N_6546,N_7852);
and U9589 (N_9589,N_6468,N_6356);
or U9590 (N_9590,N_6274,N_7393);
and U9591 (N_9591,N_7880,N_6174);
or U9592 (N_9592,N_7545,N_6322);
or U9593 (N_9593,N_6602,N_7565);
nand U9594 (N_9594,N_6295,N_7883);
nand U9595 (N_9595,N_6693,N_7948);
nor U9596 (N_9596,N_6104,N_7278);
nand U9597 (N_9597,N_7880,N_6041);
nor U9598 (N_9598,N_7986,N_6515);
xor U9599 (N_9599,N_6033,N_7551);
nor U9600 (N_9600,N_7507,N_6381);
xor U9601 (N_9601,N_7587,N_7330);
and U9602 (N_9602,N_6884,N_6176);
nand U9603 (N_9603,N_6987,N_7169);
or U9604 (N_9604,N_7046,N_6774);
nand U9605 (N_9605,N_7890,N_7315);
or U9606 (N_9606,N_6155,N_7098);
nand U9607 (N_9607,N_7958,N_6637);
nor U9608 (N_9608,N_7368,N_7895);
and U9609 (N_9609,N_6102,N_7382);
or U9610 (N_9610,N_7296,N_7247);
and U9611 (N_9611,N_7606,N_7252);
xor U9612 (N_9612,N_6722,N_7267);
or U9613 (N_9613,N_7555,N_7580);
nor U9614 (N_9614,N_7896,N_6183);
or U9615 (N_9615,N_6421,N_7542);
and U9616 (N_9616,N_6069,N_7445);
nand U9617 (N_9617,N_6204,N_6317);
and U9618 (N_9618,N_6329,N_6173);
and U9619 (N_9619,N_6205,N_6578);
or U9620 (N_9620,N_7899,N_6800);
xnor U9621 (N_9621,N_7701,N_7586);
or U9622 (N_9622,N_6168,N_6452);
or U9623 (N_9623,N_6726,N_6754);
or U9624 (N_9624,N_6488,N_7951);
nand U9625 (N_9625,N_6641,N_7342);
and U9626 (N_9626,N_7199,N_6460);
nor U9627 (N_9627,N_7180,N_7441);
and U9628 (N_9628,N_7099,N_7738);
and U9629 (N_9629,N_6089,N_6555);
nand U9630 (N_9630,N_6618,N_6206);
or U9631 (N_9631,N_7855,N_7183);
nor U9632 (N_9632,N_7539,N_6463);
and U9633 (N_9633,N_7073,N_6296);
and U9634 (N_9634,N_6688,N_6056);
xor U9635 (N_9635,N_7329,N_7529);
nor U9636 (N_9636,N_6886,N_6094);
and U9637 (N_9637,N_7227,N_7355);
nor U9638 (N_9638,N_6740,N_6536);
or U9639 (N_9639,N_7433,N_6893);
nand U9640 (N_9640,N_7432,N_7810);
nand U9641 (N_9641,N_6109,N_6704);
and U9642 (N_9642,N_7139,N_7593);
or U9643 (N_9643,N_6928,N_6936);
nor U9644 (N_9644,N_6000,N_7658);
nand U9645 (N_9645,N_7364,N_7203);
nor U9646 (N_9646,N_6425,N_7644);
or U9647 (N_9647,N_7439,N_7375);
or U9648 (N_9648,N_7104,N_6830);
or U9649 (N_9649,N_6766,N_6054);
nor U9650 (N_9650,N_6217,N_7110);
or U9651 (N_9651,N_6948,N_7919);
nand U9652 (N_9652,N_6598,N_6432);
nand U9653 (N_9653,N_7750,N_7810);
and U9654 (N_9654,N_7100,N_7063);
xor U9655 (N_9655,N_7570,N_7326);
nor U9656 (N_9656,N_7908,N_7437);
xor U9657 (N_9657,N_7149,N_6462);
or U9658 (N_9658,N_6113,N_6764);
nor U9659 (N_9659,N_6949,N_6194);
nand U9660 (N_9660,N_6009,N_7545);
nor U9661 (N_9661,N_7495,N_7676);
xor U9662 (N_9662,N_7593,N_6243);
or U9663 (N_9663,N_6285,N_6485);
and U9664 (N_9664,N_6297,N_7129);
or U9665 (N_9665,N_7372,N_6455);
and U9666 (N_9666,N_6027,N_7525);
nand U9667 (N_9667,N_6419,N_6679);
nand U9668 (N_9668,N_6513,N_7208);
nor U9669 (N_9669,N_7262,N_7923);
or U9670 (N_9670,N_7328,N_7705);
and U9671 (N_9671,N_6854,N_7639);
and U9672 (N_9672,N_6451,N_7038);
or U9673 (N_9673,N_7384,N_7884);
and U9674 (N_9674,N_7430,N_6088);
or U9675 (N_9675,N_6932,N_6133);
and U9676 (N_9676,N_6366,N_6850);
nand U9677 (N_9677,N_7207,N_7707);
or U9678 (N_9678,N_7759,N_7431);
and U9679 (N_9679,N_7365,N_7432);
nand U9680 (N_9680,N_6030,N_7375);
or U9681 (N_9681,N_6464,N_7869);
and U9682 (N_9682,N_7764,N_7148);
xnor U9683 (N_9683,N_7523,N_6262);
and U9684 (N_9684,N_6301,N_7289);
nor U9685 (N_9685,N_6700,N_7421);
nand U9686 (N_9686,N_6537,N_6324);
and U9687 (N_9687,N_6116,N_7546);
nand U9688 (N_9688,N_7081,N_7932);
xnor U9689 (N_9689,N_7380,N_7934);
or U9690 (N_9690,N_7032,N_7172);
nand U9691 (N_9691,N_7564,N_7848);
xnor U9692 (N_9692,N_6643,N_7091);
and U9693 (N_9693,N_6930,N_7498);
nand U9694 (N_9694,N_6459,N_7499);
or U9695 (N_9695,N_7589,N_7926);
or U9696 (N_9696,N_6948,N_7197);
or U9697 (N_9697,N_6254,N_6361);
or U9698 (N_9698,N_6377,N_7524);
nand U9699 (N_9699,N_7859,N_6285);
nor U9700 (N_9700,N_6588,N_7862);
nand U9701 (N_9701,N_6893,N_7965);
nor U9702 (N_9702,N_6050,N_6321);
nand U9703 (N_9703,N_6077,N_6574);
nor U9704 (N_9704,N_6112,N_6041);
or U9705 (N_9705,N_7512,N_7059);
and U9706 (N_9706,N_6094,N_6706);
nor U9707 (N_9707,N_7421,N_6590);
or U9708 (N_9708,N_6911,N_7793);
nor U9709 (N_9709,N_7035,N_7181);
nor U9710 (N_9710,N_6571,N_6801);
and U9711 (N_9711,N_6710,N_6576);
or U9712 (N_9712,N_6787,N_6372);
and U9713 (N_9713,N_6397,N_6634);
nor U9714 (N_9714,N_7713,N_7303);
or U9715 (N_9715,N_6565,N_7618);
or U9716 (N_9716,N_7268,N_6833);
xor U9717 (N_9717,N_7356,N_7762);
xnor U9718 (N_9718,N_7038,N_7499);
and U9719 (N_9719,N_6190,N_7363);
nor U9720 (N_9720,N_7867,N_7204);
or U9721 (N_9721,N_6089,N_7230);
nand U9722 (N_9722,N_7637,N_6873);
nand U9723 (N_9723,N_6400,N_7369);
and U9724 (N_9724,N_7861,N_7407);
nand U9725 (N_9725,N_6086,N_6725);
nand U9726 (N_9726,N_6791,N_6013);
xnor U9727 (N_9727,N_6511,N_7520);
and U9728 (N_9728,N_6075,N_7760);
or U9729 (N_9729,N_6547,N_6007);
nand U9730 (N_9730,N_7634,N_7414);
or U9731 (N_9731,N_6051,N_7885);
nor U9732 (N_9732,N_6037,N_7303);
or U9733 (N_9733,N_6295,N_7006);
nor U9734 (N_9734,N_6620,N_7376);
and U9735 (N_9735,N_6393,N_7478);
nand U9736 (N_9736,N_6499,N_7550);
nand U9737 (N_9737,N_7648,N_6536);
nor U9738 (N_9738,N_7732,N_7893);
nor U9739 (N_9739,N_7560,N_6019);
or U9740 (N_9740,N_7473,N_7840);
xnor U9741 (N_9741,N_6652,N_6055);
and U9742 (N_9742,N_7378,N_7124);
xor U9743 (N_9743,N_7014,N_6571);
and U9744 (N_9744,N_7737,N_7017);
nand U9745 (N_9745,N_6202,N_7139);
xor U9746 (N_9746,N_6733,N_7718);
or U9747 (N_9747,N_6525,N_6085);
and U9748 (N_9748,N_6230,N_7484);
nand U9749 (N_9749,N_7870,N_6781);
nor U9750 (N_9750,N_6935,N_7263);
and U9751 (N_9751,N_7294,N_6105);
and U9752 (N_9752,N_6374,N_6026);
nor U9753 (N_9753,N_6789,N_7010);
or U9754 (N_9754,N_6203,N_7930);
nand U9755 (N_9755,N_6635,N_6995);
and U9756 (N_9756,N_7315,N_6228);
or U9757 (N_9757,N_7812,N_6760);
or U9758 (N_9758,N_6590,N_7952);
or U9759 (N_9759,N_7858,N_7052);
and U9760 (N_9760,N_7736,N_7946);
xnor U9761 (N_9761,N_7320,N_6268);
nor U9762 (N_9762,N_7369,N_7316);
xnor U9763 (N_9763,N_6686,N_7000);
nor U9764 (N_9764,N_6157,N_7788);
or U9765 (N_9765,N_7638,N_7025);
nor U9766 (N_9766,N_7007,N_6674);
or U9767 (N_9767,N_6623,N_7805);
nor U9768 (N_9768,N_6045,N_6902);
nand U9769 (N_9769,N_7072,N_6122);
and U9770 (N_9770,N_7094,N_6531);
nor U9771 (N_9771,N_6946,N_6800);
nand U9772 (N_9772,N_6141,N_6582);
nand U9773 (N_9773,N_6210,N_6109);
xor U9774 (N_9774,N_6455,N_7375);
and U9775 (N_9775,N_6472,N_7710);
nor U9776 (N_9776,N_7186,N_6247);
xnor U9777 (N_9777,N_7273,N_7790);
nand U9778 (N_9778,N_6197,N_6491);
nor U9779 (N_9779,N_7541,N_7329);
or U9780 (N_9780,N_6292,N_6011);
and U9781 (N_9781,N_6094,N_6997);
and U9782 (N_9782,N_7460,N_6366);
xor U9783 (N_9783,N_6807,N_6272);
or U9784 (N_9784,N_6612,N_7595);
nor U9785 (N_9785,N_7936,N_7671);
and U9786 (N_9786,N_7590,N_6456);
nor U9787 (N_9787,N_6236,N_6996);
nor U9788 (N_9788,N_6037,N_7778);
nor U9789 (N_9789,N_6012,N_6074);
nor U9790 (N_9790,N_7355,N_7687);
nor U9791 (N_9791,N_6576,N_6512);
and U9792 (N_9792,N_6532,N_7663);
or U9793 (N_9793,N_6050,N_7120);
xnor U9794 (N_9794,N_7549,N_6272);
or U9795 (N_9795,N_7995,N_6470);
and U9796 (N_9796,N_6248,N_7554);
and U9797 (N_9797,N_6525,N_7048);
xor U9798 (N_9798,N_7012,N_7343);
or U9799 (N_9799,N_6041,N_6208);
nor U9800 (N_9800,N_7853,N_6598);
xnor U9801 (N_9801,N_7990,N_7315);
nor U9802 (N_9802,N_6587,N_7560);
nand U9803 (N_9803,N_6119,N_6084);
or U9804 (N_9804,N_6845,N_7043);
and U9805 (N_9805,N_7894,N_6470);
and U9806 (N_9806,N_6250,N_6920);
and U9807 (N_9807,N_7413,N_6682);
nor U9808 (N_9808,N_6892,N_6165);
nor U9809 (N_9809,N_6882,N_7400);
xor U9810 (N_9810,N_7313,N_6701);
nor U9811 (N_9811,N_6904,N_7794);
nand U9812 (N_9812,N_6379,N_7047);
and U9813 (N_9813,N_6293,N_6697);
nor U9814 (N_9814,N_7651,N_7003);
nand U9815 (N_9815,N_6819,N_7670);
nor U9816 (N_9816,N_6241,N_7303);
nand U9817 (N_9817,N_7777,N_6869);
and U9818 (N_9818,N_7014,N_7752);
nand U9819 (N_9819,N_6665,N_6796);
or U9820 (N_9820,N_7989,N_7795);
nand U9821 (N_9821,N_7355,N_6405);
nand U9822 (N_9822,N_6619,N_6638);
nor U9823 (N_9823,N_6048,N_6997);
xor U9824 (N_9824,N_7565,N_7640);
xor U9825 (N_9825,N_6135,N_6004);
or U9826 (N_9826,N_7581,N_6386);
or U9827 (N_9827,N_7376,N_7478);
xor U9828 (N_9828,N_6017,N_7245);
nand U9829 (N_9829,N_7546,N_6863);
xnor U9830 (N_9830,N_7876,N_6421);
nand U9831 (N_9831,N_6664,N_7070);
or U9832 (N_9832,N_6807,N_6281);
nor U9833 (N_9833,N_7269,N_6190);
nand U9834 (N_9834,N_7845,N_7120);
nand U9835 (N_9835,N_6500,N_6694);
nor U9836 (N_9836,N_7561,N_7439);
and U9837 (N_9837,N_7409,N_6373);
or U9838 (N_9838,N_7322,N_6295);
nor U9839 (N_9839,N_7930,N_7099);
and U9840 (N_9840,N_7794,N_7903);
nor U9841 (N_9841,N_7733,N_6857);
nand U9842 (N_9842,N_7571,N_6854);
and U9843 (N_9843,N_7895,N_7617);
and U9844 (N_9844,N_6620,N_7858);
nor U9845 (N_9845,N_7706,N_7732);
nor U9846 (N_9846,N_7676,N_6596);
nor U9847 (N_9847,N_6301,N_6740);
nand U9848 (N_9848,N_7398,N_7996);
xor U9849 (N_9849,N_6087,N_6237);
nand U9850 (N_9850,N_6042,N_6324);
nand U9851 (N_9851,N_7696,N_6737);
and U9852 (N_9852,N_7348,N_7314);
or U9853 (N_9853,N_6115,N_6961);
or U9854 (N_9854,N_6622,N_6614);
nand U9855 (N_9855,N_6706,N_7787);
or U9856 (N_9856,N_7343,N_7404);
nand U9857 (N_9857,N_7007,N_6569);
nand U9858 (N_9858,N_6482,N_7554);
xor U9859 (N_9859,N_6414,N_6983);
or U9860 (N_9860,N_7046,N_6501);
nor U9861 (N_9861,N_6350,N_7604);
nor U9862 (N_9862,N_7410,N_6071);
or U9863 (N_9863,N_6965,N_6282);
and U9864 (N_9864,N_7050,N_7653);
nor U9865 (N_9865,N_6103,N_7003);
and U9866 (N_9866,N_6073,N_6084);
or U9867 (N_9867,N_7441,N_6540);
nand U9868 (N_9868,N_7767,N_6998);
and U9869 (N_9869,N_6306,N_6357);
nand U9870 (N_9870,N_7595,N_6163);
or U9871 (N_9871,N_6623,N_7857);
nor U9872 (N_9872,N_7521,N_6594);
xnor U9873 (N_9873,N_6969,N_7331);
nand U9874 (N_9874,N_6276,N_7529);
nor U9875 (N_9875,N_7499,N_6952);
or U9876 (N_9876,N_6748,N_6098);
or U9877 (N_9877,N_7160,N_7362);
or U9878 (N_9878,N_7619,N_6259);
or U9879 (N_9879,N_7667,N_6334);
xor U9880 (N_9880,N_6079,N_7695);
nand U9881 (N_9881,N_6673,N_6873);
and U9882 (N_9882,N_6287,N_6166);
and U9883 (N_9883,N_6731,N_7611);
and U9884 (N_9884,N_6089,N_6681);
and U9885 (N_9885,N_7128,N_6075);
and U9886 (N_9886,N_7720,N_6265);
xnor U9887 (N_9887,N_7867,N_6305);
xnor U9888 (N_9888,N_6571,N_7920);
and U9889 (N_9889,N_6637,N_7186);
and U9890 (N_9890,N_7610,N_7383);
and U9891 (N_9891,N_6143,N_6560);
nand U9892 (N_9892,N_7501,N_7833);
nor U9893 (N_9893,N_6860,N_7173);
nand U9894 (N_9894,N_6339,N_6441);
nor U9895 (N_9895,N_7585,N_7027);
or U9896 (N_9896,N_6762,N_7135);
or U9897 (N_9897,N_7081,N_6739);
or U9898 (N_9898,N_7572,N_6682);
or U9899 (N_9899,N_7870,N_7029);
nand U9900 (N_9900,N_7047,N_6298);
or U9901 (N_9901,N_7654,N_6936);
or U9902 (N_9902,N_7553,N_7461);
or U9903 (N_9903,N_6946,N_6637);
xnor U9904 (N_9904,N_7077,N_6423);
and U9905 (N_9905,N_6448,N_6119);
or U9906 (N_9906,N_6802,N_6809);
nor U9907 (N_9907,N_7995,N_7454);
xor U9908 (N_9908,N_6203,N_6821);
nand U9909 (N_9909,N_7190,N_7280);
or U9910 (N_9910,N_7574,N_7498);
and U9911 (N_9911,N_7080,N_7210);
nor U9912 (N_9912,N_7824,N_6004);
or U9913 (N_9913,N_6981,N_7481);
nor U9914 (N_9914,N_7460,N_6604);
or U9915 (N_9915,N_6733,N_6074);
and U9916 (N_9916,N_7664,N_6204);
nand U9917 (N_9917,N_7720,N_6555);
xor U9918 (N_9918,N_7339,N_6183);
nor U9919 (N_9919,N_7353,N_6719);
nand U9920 (N_9920,N_7721,N_7725);
nand U9921 (N_9921,N_6417,N_7673);
nand U9922 (N_9922,N_7096,N_7324);
and U9923 (N_9923,N_6691,N_7771);
or U9924 (N_9924,N_6442,N_6487);
or U9925 (N_9925,N_6355,N_6459);
or U9926 (N_9926,N_6207,N_6037);
or U9927 (N_9927,N_7968,N_7122);
nand U9928 (N_9928,N_6491,N_6690);
or U9929 (N_9929,N_6625,N_7563);
nand U9930 (N_9930,N_6211,N_6399);
and U9931 (N_9931,N_6271,N_7536);
and U9932 (N_9932,N_7555,N_7842);
nand U9933 (N_9933,N_7189,N_6019);
or U9934 (N_9934,N_7553,N_7314);
nor U9935 (N_9935,N_6897,N_6023);
nor U9936 (N_9936,N_7218,N_6221);
or U9937 (N_9937,N_7049,N_6405);
or U9938 (N_9938,N_6498,N_7619);
and U9939 (N_9939,N_7229,N_7132);
nand U9940 (N_9940,N_7809,N_6929);
and U9941 (N_9941,N_7287,N_7843);
or U9942 (N_9942,N_7825,N_7543);
or U9943 (N_9943,N_7293,N_7079);
nor U9944 (N_9944,N_6396,N_6096);
nand U9945 (N_9945,N_6770,N_6436);
xnor U9946 (N_9946,N_7461,N_6649);
and U9947 (N_9947,N_6097,N_7440);
and U9948 (N_9948,N_7513,N_7586);
nand U9949 (N_9949,N_6993,N_6807);
nand U9950 (N_9950,N_7186,N_6684);
or U9951 (N_9951,N_7430,N_6604);
or U9952 (N_9952,N_6341,N_6239);
or U9953 (N_9953,N_6709,N_6300);
nor U9954 (N_9954,N_6287,N_6561);
xnor U9955 (N_9955,N_7486,N_7763);
or U9956 (N_9956,N_7482,N_7765);
nor U9957 (N_9957,N_6315,N_7862);
nand U9958 (N_9958,N_6017,N_7473);
or U9959 (N_9959,N_7290,N_7467);
and U9960 (N_9960,N_6962,N_7151);
or U9961 (N_9961,N_7312,N_6560);
or U9962 (N_9962,N_6009,N_6642);
or U9963 (N_9963,N_7903,N_6978);
nand U9964 (N_9964,N_6926,N_7046);
or U9965 (N_9965,N_7936,N_7291);
or U9966 (N_9966,N_6519,N_7823);
nand U9967 (N_9967,N_7140,N_7796);
nor U9968 (N_9968,N_6062,N_6327);
nand U9969 (N_9969,N_7731,N_7203);
nor U9970 (N_9970,N_7310,N_7436);
xnor U9971 (N_9971,N_7232,N_6645);
xnor U9972 (N_9972,N_7257,N_7532);
and U9973 (N_9973,N_7068,N_7962);
or U9974 (N_9974,N_7383,N_6311);
nand U9975 (N_9975,N_6717,N_7283);
and U9976 (N_9976,N_7336,N_6385);
nand U9977 (N_9977,N_7980,N_6630);
nand U9978 (N_9978,N_7938,N_7584);
nand U9979 (N_9979,N_6769,N_7909);
nor U9980 (N_9980,N_7564,N_7705);
nand U9981 (N_9981,N_7664,N_6573);
and U9982 (N_9982,N_6191,N_6112);
nor U9983 (N_9983,N_6914,N_7662);
nor U9984 (N_9984,N_6678,N_7135);
xor U9985 (N_9985,N_7978,N_6268);
xnor U9986 (N_9986,N_7115,N_7094);
nand U9987 (N_9987,N_7530,N_6563);
or U9988 (N_9988,N_6601,N_6334);
nand U9989 (N_9989,N_7744,N_7556);
xor U9990 (N_9990,N_6059,N_7624);
nor U9991 (N_9991,N_7431,N_7238);
nand U9992 (N_9992,N_6019,N_6476);
nand U9993 (N_9993,N_6019,N_7615);
and U9994 (N_9994,N_7162,N_6629);
nand U9995 (N_9995,N_7865,N_6870);
xor U9996 (N_9996,N_6441,N_6297);
nor U9997 (N_9997,N_6342,N_6917);
or U9998 (N_9998,N_7141,N_6028);
nand U9999 (N_9999,N_6315,N_6907);
and UO_0 (O_0,N_9447,N_9313);
xnor UO_1 (O_1,N_9312,N_8680);
and UO_2 (O_2,N_8073,N_8663);
nor UO_3 (O_3,N_8607,N_8134);
nand UO_4 (O_4,N_9462,N_8408);
or UO_5 (O_5,N_9124,N_9552);
and UO_6 (O_6,N_9011,N_8285);
or UO_7 (O_7,N_8967,N_9858);
and UO_8 (O_8,N_8448,N_9862);
or UO_9 (O_9,N_8279,N_8438);
and UO_10 (O_10,N_9448,N_8698);
nand UO_11 (O_11,N_8902,N_8582);
or UO_12 (O_12,N_8604,N_8165);
and UO_13 (O_13,N_8989,N_9794);
and UO_14 (O_14,N_8793,N_9138);
nand UO_15 (O_15,N_8571,N_8394);
nor UO_16 (O_16,N_9179,N_9471);
and UO_17 (O_17,N_8093,N_9082);
and UO_18 (O_18,N_8460,N_8447);
or UO_19 (O_19,N_9573,N_8685);
nand UO_20 (O_20,N_8941,N_9362);
nand UO_21 (O_21,N_8878,N_9997);
nand UO_22 (O_22,N_9140,N_8306);
and UO_23 (O_23,N_8572,N_9943);
nand UO_24 (O_24,N_9682,N_9468);
nand UO_25 (O_25,N_8221,N_9162);
nor UO_26 (O_26,N_8665,N_9657);
nand UO_27 (O_27,N_8526,N_8182);
nor UO_28 (O_28,N_8366,N_8021);
and UO_29 (O_29,N_9078,N_9610);
or UO_30 (O_30,N_9868,N_9830);
and UO_31 (O_31,N_8338,N_9044);
nand UO_32 (O_32,N_9301,N_9617);
nand UO_33 (O_33,N_8435,N_9327);
nand UO_34 (O_34,N_8331,N_8273);
and UO_35 (O_35,N_8617,N_8323);
and UO_36 (O_36,N_9959,N_8032);
xnor UO_37 (O_37,N_8493,N_8642);
and UO_38 (O_38,N_9770,N_8430);
nand UO_39 (O_39,N_9832,N_9798);
and UO_40 (O_40,N_9107,N_8076);
and UO_41 (O_41,N_8468,N_9596);
nor UO_42 (O_42,N_8223,N_8368);
nor UO_43 (O_43,N_9772,N_8217);
and UO_44 (O_44,N_9917,N_9667);
nor UO_45 (O_45,N_9771,N_9562);
and UO_46 (O_46,N_9042,N_9805);
nor UO_47 (O_47,N_9615,N_8048);
nor UO_48 (O_48,N_8973,N_8795);
nor UO_49 (O_49,N_9499,N_9844);
nor UO_50 (O_50,N_9278,N_8940);
xor UO_51 (O_51,N_8896,N_9942);
or UO_52 (O_52,N_8277,N_9674);
or UO_53 (O_53,N_9704,N_9463);
and UO_54 (O_54,N_8875,N_8138);
nand UO_55 (O_55,N_9292,N_9732);
nor UO_56 (O_56,N_8118,N_8361);
or UO_57 (O_57,N_9093,N_9636);
or UO_58 (O_58,N_9120,N_9259);
nor UO_59 (O_59,N_9150,N_9035);
nand UO_60 (O_60,N_8755,N_8262);
nand UO_61 (O_61,N_9381,N_9753);
nand UO_62 (O_62,N_8089,N_8891);
and UO_63 (O_63,N_8653,N_9670);
and UO_64 (O_64,N_9420,N_8471);
or UO_65 (O_65,N_9449,N_9650);
xnor UO_66 (O_66,N_9652,N_8066);
nand UO_67 (O_67,N_8488,N_8614);
and UO_68 (O_68,N_9863,N_8025);
nand UO_69 (O_69,N_8857,N_9626);
nand UO_70 (O_70,N_9779,N_9655);
or UO_71 (O_71,N_8806,N_8002);
nor UO_72 (O_72,N_8883,N_8079);
and UO_73 (O_73,N_9401,N_9700);
or UO_74 (O_74,N_9333,N_9752);
and UO_75 (O_75,N_8329,N_9601);
nand UO_76 (O_76,N_9612,N_8905);
and UO_77 (O_77,N_9932,N_8523);
and UO_78 (O_78,N_8742,N_9566);
or UO_79 (O_79,N_9926,N_8100);
or UO_80 (O_80,N_8606,N_8233);
and UO_81 (O_81,N_9684,N_8850);
nor UO_82 (O_82,N_9857,N_8405);
or UO_83 (O_83,N_8543,N_9902);
nor UO_84 (O_84,N_9483,N_8784);
or UO_85 (O_85,N_8881,N_9708);
and UO_86 (O_86,N_9969,N_8590);
and UO_87 (O_87,N_9939,N_8619);
or UO_88 (O_88,N_9835,N_9656);
and UO_89 (O_89,N_9878,N_9742);
and UO_90 (O_90,N_9791,N_9173);
nand UO_91 (O_91,N_8255,N_9256);
nand UO_92 (O_92,N_9909,N_9072);
nor UO_93 (O_93,N_9125,N_9980);
nor UO_94 (O_94,N_9661,N_8777);
and UO_95 (O_95,N_9892,N_9546);
or UO_96 (O_96,N_8832,N_8498);
xor UO_97 (O_97,N_8596,N_8855);
nand UO_98 (O_98,N_8879,N_9087);
nor UO_99 (O_99,N_8968,N_9789);
nor UO_100 (O_100,N_9616,N_9842);
nand UO_101 (O_101,N_9724,N_9649);
xnor UO_102 (O_102,N_8375,N_9332);
xor UO_103 (O_103,N_8414,N_8101);
nand UO_104 (O_104,N_8268,N_9368);
nor UO_105 (O_105,N_9180,N_9963);
or UO_106 (O_106,N_8239,N_9253);
or UO_107 (O_107,N_9537,N_9554);
and UO_108 (O_108,N_9973,N_8669);
and UO_109 (O_109,N_8834,N_9423);
or UO_110 (O_110,N_8031,N_9002);
and UO_111 (O_111,N_8661,N_9726);
xor UO_112 (O_112,N_9681,N_9677);
nor UO_113 (O_113,N_9116,N_8797);
nand UO_114 (O_114,N_8937,N_8278);
nand UO_115 (O_115,N_9970,N_8336);
nand UO_116 (O_116,N_9641,N_8384);
nand UO_117 (O_117,N_8019,N_8043);
nand UO_118 (O_118,N_8232,N_9936);
nand UO_119 (O_119,N_8580,N_9358);
nand UO_120 (O_120,N_8370,N_9506);
or UO_121 (O_121,N_9538,N_9430);
nor UO_122 (O_122,N_8462,N_9767);
xnor UO_123 (O_123,N_8631,N_8094);
and UO_124 (O_124,N_8303,N_8209);
xnor UO_125 (O_125,N_9911,N_9717);
nor UO_126 (O_126,N_8813,N_9203);
or UO_127 (O_127,N_8684,N_9399);
nor UO_128 (O_128,N_9436,N_8948);
and UO_129 (O_129,N_8355,N_8904);
and UO_130 (O_130,N_9136,N_9269);
or UO_131 (O_131,N_8769,N_8579);
and UO_132 (O_132,N_9157,N_9916);
and UO_133 (O_133,N_9875,N_8871);
nor UO_134 (O_134,N_8981,N_8117);
or UO_135 (O_135,N_9397,N_9500);
nor UO_136 (O_136,N_9769,N_9091);
or UO_137 (O_137,N_8102,N_8372);
nor UO_138 (O_138,N_8672,N_9193);
nor UO_139 (O_139,N_8203,N_8315);
nor UO_140 (O_140,N_8718,N_8081);
nand UO_141 (O_141,N_8719,N_8953);
or UO_142 (O_142,N_8198,N_9266);
and UO_143 (O_143,N_8723,N_9597);
or UO_144 (O_144,N_9824,N_8212);
nand UO_145 (O_145,N_8439,N_8354);
nand UO_146 (O_146,N_9073,N_8467);
nor UO_147 (O_147,N_9893,N_8915);
nand UO_148 (O_148,N_8846,N_9188);
or UO_149 (O_149,N_8720,N_9433);
and UO_150 (O_150,N_9485,N_8103);
or UO_151 (O_151,N_9428,N_8078);
and UO_152 (O_152,N_8131,N_9869);
xor UO_153 (O_153,N_8110,N_8147);
xnor UO_154 (O_154,N_8751,N_9274);
nand UO_155 (O_155,N_9599,N_9293);
and UO_156 (O_156,N_8611,N_9030);
nand UO_157 (O_157,N_8133,N_9502);
or UO_158 (O_158,N_8058,N_9317);
or UO_159 (O_159,N_9170,N_8299);
nor UO_160 (O_160,N_8782,N_9472);
and UO_161 (O_161,N_9714,N_9527);
and UO_162 (O_162,N_8838,N_8284);
or UO_163 (O_163,N_9931,N_8847);
and UO_164 (O_164,N_8528,N_9624);
nand UO_165 (O_165,N_8312,N_8229);
or UO_166 (O_166,N_9570,N_9456);
nand UO_167 (O_167,N_9046,N_8411);
and UO_168 (O_168,N_9922,N_8744);
nor UO_169 (O_169,N_8515,N_8256);
and UO_170 (O_170,N_9071,N_8302);
or UO_171 (O_171,N_8030,N_9385);
nor UO_172 (O_172,N_9414,N_8919);
nor UO_173 (O_173,N_8159,N_8119);
nand UO_174 (O_174,N_9990,N_9937);
nor UO_175 (O_175,N_8704,N_9221);
or UO_176 (O_176,N_9623,N_8433);
nor UO_177 (O_177,N_8666,N_9567);
and UO_178 (O_178,N_8282,N_9131);
nor UO_179 (O_179,N_8286,N_9968);
or UO_180 (O_180,N_8912,N_8739);
nor UO_181 (O_181,N_9803,N_9907);
or UO_182 (O_182,N_9081,N_9400);
nand UO_183 (O_183,N_8794,N_9829);
nand UO_184 (O_184,N_8445,N_8396);
nand UO_185 (O_185,N_8870,N_8441);
nor UO_186 (O_186,N_9646,N_9755);
nand UO_187 (O_187,N_9322,N_9512);
nor UO_188 (O_188,N_9240,N_9786);
and UO_189 (O_189,N_9346,N_8156);
or UO_190 (O_190,N_9279,N_9063);
xor UO_191 (O_191,N_8598,N_9629);
nor UO_192 (O_192,N_8020,N_9920);
and UO_193 (O_193,N_8042,N_8003);
nand UO_194 (O_194,N_8272,N_8550);
nand UO_195 (O_195,N_8332,N_8773);
xnor UO_196 (O_196,N_8074,N_9643);
nor UO_197 (O_197,N_9064,N_8860);
nand UO_198 (O_198,N_8911,N_9085);
or UO_199 (O_199,N_9784,N_8722);
nand UO_200 (O_200,N_9880,N_8135);
and UO_201 (O_201,N_8613,N_9508);
and UO_202 (O_202,N_8766,N_9225);
nand UO_203 (O_203,N_9437,N_9678);
nor UO_204 (O_204,N_9209,N_8862);
and UO_205 (O_205,N_8290,N_9737);
or UO_206 (O_206,N_9564,N_8819);
nand UO_207 (O_207,N_8393,N_9895);
nor UO_208 (O_208,N_9024,N_8087);
nor UO_209 (O_209,N_8573,N_8972);
nand UO_210 (O_210,N_8242,N_8296);
nor UO_211 (O_211,N_8533,N_9134);
nand UO_212 (O_212,N_9999,N_8346);
nor UO_213 (O_213,N_8949,N_9187);
nand UO_214 (O_214,N_9101,N_8310);
and UO_215 (O_215,N_9799,N_9768);
nor UO_216 (O_216,N_9204,N_8214);
nand UO_217 (O_217,N_9692,N_8564);
nor UO_218 (O_218,N_9325,N_9979);
and UO_219 (O_219,N_8950,N_8045);
nand UO_220 (O_220,N_9244,N_9183);
nor UO_221 (O_221,N_9631,N_9475);
xnor UO_222 (O_222,N_8178,N_9574);
nand UO_223 (O_223,N_9642,N_9613);
xor UO_224 (O_224,N_8207,N_8213);
and UO_225 (O_225,N_8506,N_9645);
or UO_226 (O_226,N_9001,N_9380);
nand UO_227 (O_227,N_8179,N_9248);
nand UO_228 (O_228,N_8235,N_9533);
and UO_229 (O_229,N_9739,N_9930);
nand UO_230 (O_230,N_9944,N_9580);
nand UO_231 (O_231,N_9861,N_8190);
and UO_232 (O_232,N_8417,N_8099);
and UO_233 (O_233,N_8283,N_8645);
nor UO_234 (O_234,N_8839,N_9996);
nor UO_235 (O_235,N_8222,N_8809);
or UO_236 (O_236,N_8916,N_9812);
or UO_237 (O_237,N_9718,N_9127);
nor UO_238 (O_238,N_9915,N_8535);
or UO_239 (O_239,N_9370,N_8309);
and UO_240 (O_240,N_9320,N_9137);
or UO_241 (O_241,N_9060,N_8443);
and UO_242 (O_242,N_9286,N_9154);
nor UO_243 (O_243,N_8593,N_9347);
nor UO_244 (O_244,N_9254,N_8215);
or UO_245 (O_245,N_9490,N_8798);
or UO_246 (O_246,N_8995,N_8899);
xnor UO_247 (O_247,N_8330,N_9149);
nor UO_248 (O_248,N_8097,N_8216);
or UO_249 (O_249,N_8051,N_8056);
nor UO_250 (O_250,N_9242,N_8261);
nand UO_251 (O_251,N_8345,N_8432);
nor UO_252 (O_252,N_9745,N_9584);
nor UO_253 (O_253,N_8401,N_9727);
nand UO_254 (O_254,N_8900,N_8511);
or UO_255 (O_255,N_8587,N_9429);
or UO_256 (O_256,N_8426,N_9146);
and UO_257 (O_257,N_8141,N_8226);
or UO_258 (O_258,N_8077,N_8630);
and UO_259 (O_259,N_9860,N_8162);
nand UO_260 (O_260,N_8091,N_8544);
and UO_261 (O_261,N_8893,N_8601);
nor UO_262 (O_262,N_9453,N_8028);
nor UO_263 (O_263,N_8369,N_8690);
nand UO_264 (O_264,N_9948,N_9310);
or UO_265 (O_265,N_9166,N_9051);
nor UO_266 (O_266,N_9432,N_9918);
and UO_267 (O_267,N_8926,N_8068);
nand UO_268 (O_268,N_8470,N_8188);
or UO_269 (O_269,N_9142,N_8745);
and UO_270 (O_270,N_8691,N_8276);
nor UO_271 (O_271,N_8970,N_9473);
nand UO_272 (O_272,N_9470,N_8116);
nand UO_273 (O_273,N_9343,N_8907);
or UO_274 (O_274,N_8576,N_8602);
nor UO_275 (O_275,N_9455,N_8933);
nor UO_276 (O_276,N_8339,N_9634);
or UO_277 (O_277,N_9062,N_8145);
or UO_278 (O_278,N_8481,N_8748);
or UO_279 (O_279,N_8854,N_8407);
nand UO_280 (O_280,N_8497,N_9205);
or UO_281 (O_281,N_8489,N_9495);
xnor UO_282 (O_282,N_8906,N_9509);
nand UO_283 (O_283,N_9043,N_9602);
and UO_284 (O_284,N_8787,N_8901);
or UO_285 (O_285,N_8126,N_9820);
nor UO_286 (O_286,N_9439,N_8274);
nand UO_287 (O_287,N_8344,N_8199);
nor UO_288 (O_288,N_8674,N_9938);
and UO_289 (O_289,N_9021,N_8749);
nor UO_290 (O_290,N_8326,N_9498);
and UO_291 (O_291,N_8562,N_8731);
nor UO_292 (O_292,N_8466,N_9738);
xor UO_293 (O_293,N_8792,N_9489);
and UO_294 (O_294,N_9625,N_9689);
nor UO_295 (O_295,N_9339,N_9912);
nand UO_296 (O_296,N_9033,N_9773);
nand UO_297 (O_297,N_9800,N_9129);
and UO_298 (O_298,N_8120,N_9666);
and UO_299 (O_299,N_9776,N_9846);
nand UO_300 (O_300,N_8501,N_8985);
nor UO_301 (O_301,N_9000,N_8741);
nand UO_302 (O_302,N_8541,N_9598);
or UO_303 (O_303,N_9790,N_8542);
nand UO_304 (O_304,N_8649,N_9231);
or UO_305 (O_305,N_8477,N_8636);
nor UO_306 (O_306,N_8801,N_8740);
nand UO_307 (O_307,N_9496,N_9268);
or UO_308 (O_308,N_8422,N_8808);
and UO_309 (O_309,N_9352,N_9925);
nand UO_310 (O_310,N_8772,N_8173);
nor UO_311 (O_311,N_9484,N_8646);
nor UO_312 (O_312,N_9628,N_9549);
nor UO_313 (O_313,N_8584,N_8936);
and UO_314 (O_314,N_9763,N_8965);
or UO_315 (O_315,N_9984,N_8292);
or UO_316 (O_316,N_8993,N_9199);
and UO_317 (O_317,N_9633,N_9705);
or UO_318 (O_318,N_9518,N_9295);
or UO_319 (O_319,N_8708,N_8668);
and UO_320 (O_320,N_9885,N_9560);
or UO_321 (O_321,N_8454,N_9810);
or UO_322 (O_322,N_8880,N_8037);
nand UO_323 (O_323,N_8423,N_9898);
nor UO_324 (O_324,N_9547,N_8457);
nor UO_325 (O_325,N_9321,N_8531);
or UO_326 (O_326,N_9836,N_9006);
or UO_327 (O_327,N_8492,N_9144);
or UO_328 (O_328,N_8856,N_8183);
nor UO_329 (O_329,N_8342,N_9066);
or UO_330 (O_330,N_8828,N_8660);
nor UO_331 (O_331,N_8410,N_8496);
nand UO_332 (O_332,N_8007,N_8565);
nand UO_333 (O_333,N_8238,N_8465);
and UO_334 (O_334,N_9614,N_9565);
xnor UO_335 (O_335,N_9017,N_8267);
and UO_336 (O_336,N_9079,N_8510);
xnor UO_337 (O_337,N_8352,N_9958);
nand UO_338 (O_338,N_9572,N_9735);
and UO_339 (O_339,N_8829,N_8867);
nand UO_340 (O_340,N_9059,N_8169);
nor UO_341 (O_341,N_8865,N_9395);
nor UO_342 (O_342,N_8696,N_8491);
or UO_343 (O_343,N_9593,N_8415);
nor UO_344 (O_344,N_8035,N_8189);
and UO_345 (O_345,N_9294,N_9806);
and UO_346 (O_346,N_9351,N_9505);
nor UO_347 (O_347,N_9644,N_8799);
or UO_348 (O_348,N_9964,N_9581);
nor UO_349 (O_349,N_9444,N_9476);
nor UO_350 (O_350,N_8754,N_9672);
and UO_351 (O_351,N_9741,N_9659);
and UO_352 (O_352,N_8574,N_9874);
nor UO_353 (O_353,N_9298,N_9843);
nand UO_354 (O_354,N_9353,N_8699);
nor UO_355 (O_355,N_8098,N_8929);
nor UO_356 (O_356,N_8052,N_8882);
nor UO_357 (O_357,N_8783,N_8337);
nand UO_358 (O_358,N_9185,N_9442);
nor UO_359 (O_359,N_9838,N_8791);
and UO_360 (O_360,N_8758,N_9540);
or UO_361 (O_361,N_9426,N_8264);
nor UO_362 (O_362,N_9775,N_9622);
xor UO_363 (O_363,N_9637,N_9693);
nor UO_364 (O_364,N_8086,N_8321);
and UO_365 (O_365,N_8513,N_9675);
or UO_366 (O_366,N_9276,N_8265);
nand UO_367 (O_367,N_8577,N_9184);
or UO_368 (O_368,N_8958,N_9034);
nand UO_369 (O_369,N_9220,N_9924);
nand UO_370 (O_370,N_8804,N_9872);
or UO_371 (O_371,N_9323,N_9019);
xnor UO_372 (O_372,N_8026,N_8805);
or UO_373 (O_373,N_8583,N_8537);
nand UO_374 (O_374,N_8317,N_8210);
xnor UO_375 (O_375,N_8934,N_9378);
or UO_376 (O_376,N_8931,N_9685);
or UO_377 (O_377,N_8530,N_8534);
or UO_378 (O_378,N_8248,N_8538);
or UO_379 (O_379,N_9635,N_9976);
or UO_380 (O_380,N_9630,N_8313);
or UO_381 (O_381,N_8942,N_8236);
xor UO_382 (O_382,N_9450,N_9639);
nand UO_383 (O_383,N_9416,N_9045);
nand UO_384 (O_384,N_9284,N_8557);
nor UO_385 (O_385,N_8055,N_8304);
nor UO_386 (O_386,N_9270,N_8129);
nand UO_387 (O_387,N_8288,N_8823);
nand UO_388 (O_388,N_8689,N_8810);
and UO_389 (O_389,N_9403,N_8923);
nand UO_390 (O_390,N_8259,N_9515);
or UO_391 (O_391,N_8503,N_8623);
nor UO_392 (O_392,N_8560,N_9023);
nand UO_393 (O_393,N_9523,N_9954);
nand UO_394 (O_394,N_8177,N_9531);
xnor UO_395 (O_395,N_8171,N_8114);
nand UO_396 (O_396,N_8391,N_8898);
nor UO_397 (O_397,N_9558,N_8966);
or UO_398 (O_398,N_8301,N_8084);
nand UO_399 (O_399,N_9757,N_9519);
or UO_400 (O_400,N_9594,N_9910);
nand UO_401 (O_401,N_8127,N_8340);
or UO_402 (O_402,N_8765,N_8472);
nor UO_403 (O_403,N_9522,N_8049);
or UO_404 (O_404,N_9961,N_9454);
nand UO_405 (O_405,N_9307,N_9854);
or UO_406 (O_406,N_9853,N_8016);
nand UO_407 (O_407,N_9383,N_9516);
or UO_408 (O_408,N_8195,N_8320);
nor UO_409 (O_409,N_8559,N_8736);
or UO_410 (O_410,N_9406,N_8727);
nand UO_411 (O_411,N_9663,N_9725);
nor UO_412 (O_412,N_8886,N_9905);
or UO_413 (O_413,N_9065,N_8759);
or UO_414 (O_414,N_8566,N_8874);
or UO_415 (O_415,N_9796,N_8548);
xnor UO_416 (O_416,N_9966,N_9047);
nand UO_417 (O_417,N_8975,N_9813);
nor UO_418 (O_418,N_8353,N_8701);
nor UO_419 (O_419,N_9354,N_9344);
nor UO_420 (O_420,N_8647,N_8225);
or UO_421 (O_421,N_9673,N_8123);
nand UO_422 (O_422,N_9342,N_8873);
nor UO_423 (O_423,N_9335,N_9543);
and UO_424 (O_424,N_9299,N_8597);
nor UO_425 (O_425,N_8908,N_8640);
or UO_426 (O_426,N_9955,N_9251);
or UO_427 (O_427,N_8293,N_9336);
nand UO_428 (O_428,N_9840,N_8569);
nand UO_429 (O_429,N_9913,N_9049);
or UO_430 (O_430,N_8191,N_9591);
xnor UO_431 (O_431,N_8633,N_9576);
and UO_432 (O_432,N_8756,N_9713);
nand UO_433 (O_433,N_8763,N_9788);
nor UO_434 (O_434,N_9553,N_8122);
and UO_435 (O_435,N_9109,N_8667);
and UO_436 (O_436,N_8108,N_9272);
or UO_437 (O_437,N_8107,N_9367);
and UO_438 (O_438,N_8984,N_9707);
xor UO_439 (O_439,N_9394,N_8512);
or UO_440 (O_440,N_8298,N_8918);
or UO_441 (O_441,N_9418,N_9215);
and UO_442 (O_442,N_8376,N_8767);
xnor UO_443 (O_443,N_9097,N_9056);
nor UO_444 (O_444,N_8271,N_8603);
nor UO_445 (O_445,N_9219,N_8735);
nor UO_446 (O_446,N_8206,N_8047);
nor UO_447 (O_447,N_8943,N_8888);
nand UO_448 (O_448,N_8788,N_8157);
nand UO_449 (O_449,N_9891,N_9621);
xnor UO_450 (O_450,N_9903,N_8452);
xor UO_451 (O_451,N_9477,N_9927);
and UO_452 (O_452,N_8451,N_9291);
or UO_453 (O_453,N_8747,N_9172);
nor UO_454 (O_454,N_9882,N_8446);
nor UO_455 (O_455,N_9052,N_8518);
nand UO_456 (O_456,N_8062,N_8529);
or UO_457 (O_457,N_8017,N_8022);
nand UO_458 (O_458,N_9384,N_9290);
and UO_459 (O_459,N_8517,N_9192);
or UO_460 (O_460,N_9702,N_8692);
and UO_461 (O_461,N_9460,N_8616);
and UO_462 (O_462,N_9398,N_9921);
nand UO_463 (O_463,N_9316,N_8453);
nand UO_464 (O_464,N_8504,N_9126);
nand UO_465 (O_465,N_8914,N_9491);
xor UO_466 (O_466,N_9348,N_9080);
nand UO_467 (O_467,N_9972,N_8487);
and UO_468 (O_468,N_9458,N_8715);
nor UO_469 (O_469,N_8884,N_9112);
and UO_470 (O_470,N_9876,N_8418);
and UO_471 (O_471,N_8673,N_8036);
and UO_472 (O_472,N_9595,N_9532);
nor UO_473 (O_473,N_9809,N_8687);
and UO_474 (O_474,N_8525,N_9671);
and UO_475 (O_475,N_9239,N_8132);
nor UO_476 (O_476,N_9451,N_9711);
or UO_477 (O_477,N_9092,N_9425);
xnor UO_478 (O_478,N_9855,N_9949);
and UO_479 (O_479,N_9361,N_8551);
nand UO_480 (O_480,N_8395,N_9619);
nand UO_481 (O_481,N_8743,N_8686);
and UO_482 (O_482,N_8187,N_8254);
and UO_483 (O_483,N_9828,N_9440);
nor UO_484 (O_484,N_8591,N_8351);
and UO_485 (O_485,N_8644,N_8656);
or UO_486 (O_486,N_9556,N_8851);
nor UO_487 (O_487,N_8090,N_8567);
or UO_488 (O_488,N_8054,N_9664);
nor UO_489 (O_489,N_9265,N_9337);
and UO_490 (O_490,N_9147,N_9094);
nor UO_491 (O_491,N_9994,N_8796);
and UO_492 (O_492,N_9946,N_8681);
or UO_493 (O_493,N_9818,N_9410);
or UO_494 (O_494,N_8046,N_8612);
nand UO_495 (O_495,N_8520,N_9764);
or UO_496 (O_496,N_8027,N_8275);
or UO_497 (O_497,N_8963,N_8335);
nor UO_498 (O_498,N_8664,N_9419);
xnor UO_499 (O_499,N_8170,N_9494);
nand UO_500 (O_500,N_9007,N_8626);
nor UO_501 (O_501,N_9578,N_8291);
nand UO_502 (O_502,N_8897,N_8979);
nand UO_503 (O_503,N_9113,N_9890);
and UO_504 (O_504,N_9196,N_9257);
xnor UO_505 (O_505,N_9234,N_8634);
xor UO_506 (O_506,N_8821,N_9371);
or UO_507 (O_507,N_9366,N_9823);
nand UO_508 (O_508,N_8869,N_9762);
or UO_509 (O_509,N_9245,N_8153);
and UO_510 (O_510,N_9901,N_9900);
xor UO_511 (O_511,N_9716,N_9743);
and UO_512 (O_512,N_9283,N_8982);
xnor UO_513 (O_513,N_9089,N_9856);
or UO_514 (O_514,N_8234,N_8494);
or UO_515 (O_515,N_9983,N_9632);
or UO_516 (O_516,N_8925,N_8539);
or UO_517 (O_517,N_9504,N_9638);
or UO_518 (O_518,N_8954,N_8244);
or UO_519 (O_519,N_9058,N_8409);
or UO_520 (O_520,N_8281,N_8890);
nand UO_521 (O_521,N_8161,N_9226);
nor UO_522 (O_522,N_8155,N_8251);
nand UO_523 (O_523,N_9758,N_9559);
or UO_524 (O_524,N_8001,N_8263);
or UO_525 (O_525,N_8760,N_8628);
xor UO_526 (O_526,N_9161,N_9409);
or UO_527 (O_527,N_9402,N_9445);
and UO_528 (O_528,N_8554,N_8137);
and UO_529 (O_529,N_8381,N_8246);
nand UO_530 (O_530,N_9801,N_8946);
and UO_531 (O_531,N_9237,N_8944);
and UO_532 (O_532,N_9759,N_9376);
xor UO_533 (O_533,N_8677,N_9018);
or UO_534 (O_534,N_9488,N_9514);
and UO_535 (O_535,N_8679,N_8064);
xnor UO_536 (O_536,N_8746,N_9871);
nor UO_537 (O_537,N_9548,N_8627);
and UO_538 (O_538,N_8913,N_8347);
and UO_539 (O_539,N_9686,N_8961);
and UO_540 (O_540,N_8519,N_8311);
and UO_541 (O_541,N_8951,N_9482);
xnor UO_542 (O_542,N_8521,N_8459);
nor UO_543 (O_543,N_9665,N_9139);
nor UO_544 (O_544,N_8753,N_8175);
or UO_545 (O_545,N_9088,N_8781);
or UO_546 (O_546,N_8420,N_8289);
nor UO_547 (O_547,N_8181,N_8670);
or UO_548 (O_548,N_9105,N_9988);
nor UO_549 (O_549,N_8154,N_8478);
nor UO_550 (O_550,N_9302,N_9356);
nor UO_551 (O_551,N_9217,N_8474);
or UO_552 (O_552,N_8243,N_9914);
and UO_553 (O_553,N_9676,N_9151);
or UO_554 (O_554,N_9777,N_8816);
xnor UO_555 (O_555,N_9202,N_8508);
and UO_556 (O_556,N_9501,N_8514);
nand UO_557 (O_557,N_8067,N_9747);
nor UO_558 (O_558,N_9213,N_8280);
nor UO_559 (O_559,N_9068,N_9104);
nor UO_560 (O_560,N_8700,N_9600);
or UO_561 (O_561,N_9841,N_9411);
or UO_562 (O_562,N_8682,N_9363);
nor UO_563 (O_563,N_8359,N_8151);
and UO_564 (O_564,N_9350,N_8622);
and UO_565 (O_565,N_9730,N_9551);
or UO_566 (O_566,N_8714,N_9864);
or UO_567 (O_567,N_8618,N_8499);
or UO_568 (O_568,N_8818,N_8057);
nand UO_569 (O_569,N_9611,N_9870);
nor UO_570 (O_570,N_9555,N_9859);
and UO_571 (O_571,N_8142,N_8938);
nor UO_572 (O_572,N_8683,N_8479);
nand UO_573 (O_573,N_9582,N_8658);
nor UO_574 (O_574,N_9375,N_8992);
xor UO_575 (O_575,N_8877,N_9252);
and UO_576 (O_576,N_8654,N_9783);
nor UO_577 (O_577,N_9492,N_9261);
xor UO_578 (O_578,N_8341,N_8476);
nand UO_579 (O_579,N_8922,N_8662);
nor UO_580 (O_580,N_9474,N_9487);
nor UO_581 (O_581,N_9324,N_9427);
and UO_582 (O_582,N_9744,N_8349);
nand UO_583 (O_583,N_9404,N_8706);
nand UO_584 (O_584,N_9951,N_8357);
or UO_585 (O_585,N_9698,N_8978);
or UO_586 (O_586,N_9372,N_9412);
and UO_587 (O_587,N_9015,N_9176);
and UO_588 (O_588,N_9568,N_9728);
nand UO_589 (O_589,N_8845,N_9503);
and UO_590 (O_590,N_8615,N_8397);
and UO_591 (O_591,N_8428,N_8532);
and UO_592 (O_592,N_9163,N_8437);
nor UO_593 (O_593,N_8034,N_9178);
nand UO_594 (O_594,N_8803,N_8143);
nand UO_595 (O_595,N_9760,N_8778);
xnor UO_596 (O_596,N_8115,N_9379);
nand UO_597 (O_597,N_8012,N_8676);
and UO_598 (O_598,N_8389,N_8581);
and UO_599 (O_599,N_9275,N_9797);
xnor UO_600 (O_600,N_8149,N_8575);
nand UO_601 (O_601,N_9987,N_8322);
nand UO_602 (O_602,N_8711,N_9721);
nand UO_603 (O_603,N_8413,N_8610);
xnor UO_604 (O_604,N_8671,N_9194);
or UO_605 (O_605,N_8833,N_9706);
nand UO_606 (O_606,N_9210,N_8991);
nand UO_607 (O_607,N_9544,N_9941);
nor UO_608 (O_608,N_8996,N_9765);
nand UO_609 (O_609,N_8319,N_9155);
xnor UO_610 (O_610,N_9981,N_9620);
or UO_611 (O_611,N_9719,N_8297);
nand UO_612 (O_612,N_9679,N_8876);
nand UO_613 (O_613,N_8522,N_9238);
nand UO_614 (O_614,N_8750,N_8945);
nor UO_615 (O_615,N_8842,N_9821);
and UO_616 (O_616,N_9029,N_9604);
and UO_617 (O_617,N_8377,N_8358);
nor UO_618 (O_618,N_8294,N_9074);
and UO_619 (O_619,N_9577,N_8400);
nand UO_620 (O_620,N_9422,N_9067);
xor UO_621 (O_621,N_8412,N_9466);
or UO_622 (O_622,N_9746,N_9694);
or UO_623 (O_623,N_8815,N_9834);
or UO_624 (O_624,N_8814,N_8717);
nand UO_625 (O_625,N_8712,N_8713);
or UO_626 (O_626,N_9695,N_9119);
nor UO_627 (O_627,N_8092,N_9446);
and UO_628 (O_628,N_8609,N_8659);
nor UO_629 (O_629,N_9651,N_9881);
nand UO_630 (O_630,N_8121,N_9025);
and UO_631 (O_631,N_8536,N_9683);
nor UO_632 (O_632,N_8629,N_8558);
and UO_633 (O_633,N_9434,N_8125);
and UO_634 (O_634,N_9223,N_8779);
nand UO_635 (O_635,N_9083,N_9647);
and UO_636 (O_636,N_8325,N_8406);
nand UO_637 (O_637,N_9793,N_9609);
and UO_638 (O_638,N_8475,N_9586);
nand UO_639 (O_639,N_8675,N_8148);
nand UO_640 (O_640,N_8392,N_8861);
nand UO_641 (O_641,N_8269,N_9431);
and UO_642 (O_642,N_8257,N_8327);
xor UO_643 (O_643,N_9075,N_8450);
nor UO_644 (O_644,N_9897,N_9208);
and UO_645 (O_645,N_8194,N_9004);
nand UO_646 (O_646,N_9575,N_8252);
nand UO_647 (O_647,N_8463,N_9285);
and UO_648 (O_648,N_9145,N_9703);
nand UO_649 (O_649,N_8053,N_8927);
or UO_650 (O_650,N_8624,N_8378);
nor UO_651 (O_651,N_9304,N_8863);
nand UO_652 (O_652,N_9115,N_8374);
and UO_653 (O_653,N_9699,N_9005);
and UO_654 (O_654,N_8652,N_9096);
nand UO_655 (O_655,N_8356,N_9012);
or UO_656 (O_656,N_8044,N_9040);
nor UO_657 (O_657,N_9883,N_9879);
nor UO_658 (O_658,N_9241,N_9212);
and UO_659 (O_659,N_8549,N_8495);
nand UO_660 (O_660,N_9364,N_8085);
nor UO_661 (O_661,N_8318,N_9103);
nor UO_662 (O_662,N_9550,N_8848);
or UO_663 (O_663,N_9687,N_9528);
or UO_664 (O_664,N_8737,N_9592);
and UO_665 (O_665,N_9696,N_8947);
and UO_666 (O_666,N_9054,N_9169);
nand UO_667 (O_667,N_8160,N_9053);
and UO_668 (O_668,N_9908,N_9391);
nand UO_669 (O_669,N_8348,N_8295);
and UO_670 (O_670,N_9975,N_9027);
or UO_671 (O_671,N_8193,N_9392);
nand UO_672 (O_672,N_8811,N_8071);
or UO_673 (O_673,N_9833,N_8218);
or UO_674 (O_674,N_9608,N_9408);
or UO_675 (O_675,N_8648,N_9816);
or UO_676 (O_676,N_8599,N_9754);
xnor UO_677 (O_677,N_8111,N_8253);
xor UO_678 (O_678,N_9099,N_9731);
nand UO_679 (O_679,N_8910,N_8419);
xnor UO_680 (O_680,N_8008,N_8703);
nor UO_681 (O_681,N_8500,N_9848);
and UO_682 (O_682,N_8657,N_9326);
nor UO_683 (O_683,N_9435,N_8469);
and UO_684 (O_684,N_8775,N_9845);
nand UO_685 (O_685,N_8444,N_9165);
nand UO_686 (O_686,N_8040,N_8545);
nand UO_687 (O_687,N_9282,N_8721);
nor UO_688 (O_688,N_8563,N_8436);
nor UO_689 (O_689,N_8632,N_9357);
xnor UO_690 (O_690,N_8716,N_9814);
nand UO_691 (O_691,N_8018,N_8600);
nand UO_692 (O_692,N_8464,N_9110);
nor UO_693 (O_693,N_8449,N_8786);
or UO_694 (O_694,N_9989,N_9417);
nand UO_695 (O_695,N_9050,N_9766);
or UO_696 (O_696,N_9386,N_8096);
nand UO_697 (O_697,N_8570,N_9839);
and UO_698 (O_698,N_9229,N_9756);
or UO_699 (O_699,N_9026,N_8894);
nor UO_700 (O_700,N_9534,N_8552);
nand UO_701 (O_701,N_8429,N_9355);
nand UO_702 (O_702,N_9952,N_8702);
xor UO_703 (O_703,N_9525,N_9130);
nand UO_704 (O_704,N_8228,N_9303);
and UO_705 (O_705,N_9090,N_8762);
nand UO_706 (O_706,N_9971,N_9175);
nor UO_707 (O_707,N_9709,N_9782);
nor UO_708 (O_708,N_9712,N_9720);
or UO_709 (O_709,N_9894,N_8650);
and UO_710 (O_710,N_9070,N_8732);
or UO_711 (O_711,N_9945,N_8697);
and UO_712 (O_712,N_8000,N_9811);
xnor UO_713 (O_713,N_8885,N_8490);
and UO_714 (O_714,N_9513,N_8130);
and UO_715 (O_715,N_9143,N_9819);
or UO_716 (O_716,N_8987,N_8385);
and UO_717 (O_717,N_9114,N_9481);
or UO_718 (O_718,N_8822,N_8964);
or UO_719 (O_719,N_9232,N_9057);
nor UO_720 (O_720,N_9956,N_8425);
and UO_721 (O_721,N_8362,N_9247);
nor UO_722 (O_722,N_8757,N_8176);
nor UO_723 (O_723,N_9701,N_8015);
or UO_724 (O_724,N_9947,N_9271);
nand UO_725 (O_725,N_9960,N_9349);
nand UO_726 (O_726,N_8924,N_8637);
or UO_727 (O_727,N_9873,N_8050);
xor UO_728 (O_728,N_9396,N_9978);
or UO_729 (O_729,N_9211,N_8859);
nand UO_730 (O_730,N_9561,N_8868);
nand UO_731 (O_731,N_9465,N_8895);
and UO_732 (O_732,N_8903,N_9106);
or UO_733 (O_733,N_8069,N_8080);
or UO_734 (O_734,N_8009,N_9013);
and UO_735 (O_735,N_9545,N_8305);
nand UO_736 (O_736,N_8023,N_9539);
nor UO_737 (O_737,N_9135,N_9201);
nor UO_738 (O_738,N_9148,N_9438);
and UO_739 (O_739,N_9181,N_8163);
and UO_740 (O_740,N_8761,N_9887);
nand UO_741 (O_741,N_8841,N_8620);
and UO_742 (O_742,N_9986,N_9452);
or UO_743 (O_743,N_8780,N_9929);
nand UO_744 (O_744,N_9467,N_8635);
or UO_745 (O_745,N_8258,N_8039);
xor UO_746 (O_746,N_8314,N_8005);
nor UO_747 (O_747,N_8128,N_9214);
nor UO_748 (O_748,N_9831,N_8399);
and UO_749 (O_749,N_8962,N_8969);
nand UO_750 (O_750,N_8245,N_9723);
and UO_751 (O_751,N_8920,N_8561);
and UO_752 (O_752,N_8866,N_9588);
nor UO_753 (O_753,N_9263,N_9524);
xnor UO_754 (O_754,N_8434,N_8776);
or UO_755 (O_755,N_8485,N_8421);
or UO_756 (O_756,N_8858,N_9517);
and UO_757 (O_757,N_9520,N_9998);
or UO_758 (O_758,N_9390,N_9825);
nand UO_759 (O_759,N_8586,N_8307);
or UO_760 (O_760,N_9413,N_8072);
or UO_761 (O_761,N_9098,N_8360);
nand UO_762 (O_762,N_9688,N_9627);
nor UO_763 (O_763,N_9690,N_9479);
xor UO_764 (O_764,N_9486,N_8553);
nor UO_765 (O_765,N_9345,N_9255);
nor UO_766 (O_766,N_9388,N_9359);
or UO_767 (O_767,N_8887,N_9511);
or UO_768 (O_768,N_8174,N_9653);
nor UO_769 (O_769,N_8167,N_9309);
or UO_770 (O_770,N_8260,N_9530);
nor UO_771 (O_771,N_8270,N_9660);
xnor UO_772 (O_772,N_8427,N_8817);
and UO_773 (O_773,N_8844,N_9607);
and UO_774 (O_774,N_8932,N_9153);
nand UO_775 (O_775,N_8424,N_8728);
and UO_776 (O_776,N_8480,N_9262);
or UO_777 (O_777,N_9167,N_9300);
nor UO_778 (O_778,N_9497,N_9847);
nand UO_779 (O_779,N_8524,N_8196);
xor UO_780 (O_780,N_9605,N_9010);
nand UO_781 (O_781,N_8184,N_8373);
or UO_782 (O_782,N_9393,N_9111);
nand UO_783 (O_783,N_8219,N_8186);
nand UO_784 (O_784,N_8038,N_9851);
nor UO_785 (O_785,N_8333,N_9016);
nand UO_786 (O_786,N_8390,N_9076);
or UO_787 (O_787,N_9585,N_8830);
nand UO_788 (O_788,N_9950,N_9227);
nand UO_789 (O_789,N_9529,N_8840);
nand UO_790 (O_790,N_8928,N_8802);
and UO_791 (O_791,N_8789,N_9778);
xor UO_792 (O_792,N_8224,N_8546);
and UO_793 (O_793,N_9311,N_9373);
xor UO_794 (O_794,N_8502,N_9478);
xor UO_795 (O_795,N_8367,N_8166);
and UO_796 (O_796,N_8158,N_8955);
nand UO_797 (O_797,N_9258,N_8308);
nand UO_798 (O_798,N_8825,N_9933);
nor UO_799 (O_799,N_9207,N_8152);
and UO_800 (O_800,N_8729,N_8033);
and UO_801 (O_801,N_9817,N_8364);
nand UO_802 (O_802,N_9850,N_8589);
xnor UO_803 (O_803,N_8440,N_9077);
xor UO_804 (O_804,N_9795,N_9329);
or UO_805 (O_805,N_9541,N_9934);
nor UO_806 (O_806,N_9186,N_9974);
or UO_807 (O_807,N_8379,N_9521);
and UO_808 (O_808,N_9122,N_8638);
or UO_809 (O_809,N_8621,N_9493);
or UO_810 (O_810,N_9906,N_8853);
nand UO_811 (O_811,N_9507,N_9250);
nand UO_812 (O_812,N_8643,N_9957);
or UO_813 (O_813,N_8820,N_9587);
and UO_814 (O_814,N_8921,N_9991);
nor UO_815 (O_815,N_9877,N_8843);
nand UO_816 (O_816,N_8180,N_8835);
nand UO_817 (O_817,N_9128,N_8688);
and UO_818 (O_818,N_9246,N_9039);
nand UO_819 (O_819,N_9164,N_9953);
nand UO_820 (O_820,N_9787,N_9038);
and UO_821 (O_821,N_8726,N_8956);
nor UO_822 (O_822,N_9736,N_9589);
or UO_823 (O_823,N_9280,N_9780);
xnor UO_824 (O_824,N_8249,N_8112);
nand UO_825 (O_825,N_9222,N_8328);
or UO_826 (O_826,N_8768,N_8807);
nor UO_827 (O_827,N_8431,N_9792);
and UO_828 (O_828,N_9100,N_9648);
nand UO_829 (O_829,N_8509,N_8484);
and UO_830 (O_830,N_9123,N_8710);
and UO_831 (O_831,N_9305,N_8365);
nor UO_832 (O_832,N_8930,N_8461);
nor UO_833 (O_833,N_8105,N_9141);
nor UO_834 (O_834,N_8957,N_8486);
or UO_835 (O_835,N_9159,N_9028);
nand UO_836 (O_836,N_8800,N_9338);
or UO_837 (O_837,N_9967,N_8693);
or UO_838 (O_838,N_9748,N_8404);
nor UO_839 (O_839,N_9009,N_8061);
and UO_840 (O_840,N_8482,N_8771);
and UO_841 (O_841,N_9314,N_9377);
nor UO_842 (O_842,N_8568,N_8146);
nor UO_843 (O_843,N_9118,N_9733);
or UO_844 (O_844,N_9867,N_9387);
nand UO_845 (O_845,N_8836,N_8205);
and UO_846 (O_846,N_9160,N_8977);
nor UO_847 (O_847,N_8104,N_8266);
or UO_848 (O_848,N_9297,N_8608);
nand UO_849 (O_849,N_8124,N_9365);
and UO_850 (O_850,N_9031,N_9669);
nand UO_851 (O_851,N_8398,N_9190);
nor UO_852 (O_852,N_8473,N_9569);
nor UO_853 (O_853,N_8507,N_8651);
and UO_854 (O_854,N_9243,N_8812);
nor UO_855 (O_855,N_9224,N_8733);
or UO_856 (O_856,N_8774,N_8088);
or UO_857 (O_857,N_8200,N_8959);
or UO_858 (O_858,N_9415,N_8852);
or UO_859 (O_859,N_8324,N_8029);
nor UO_860 (O_860,N_8363,N_9866);
and UO_861 (O_861,N_8220,N_8872);
xor UO_862 (O_862,N_9328,N_9233);
or UO_863 (O_863,N_9459,N_9340);
nand UO_864 (O_864,N_9405,N_9095);
nor UO_865 (O_865,N_8416,N_8082);
or UO_866 (O_866,N_9084,N_9571);
and UO_867 (O_867,N_9837,N_8555);
or UO_868 (O_868,N_8960,N_9583);
nand UO_869 (O_869,N_9102,N_9715);
nand UO_870 (O_870,N_8316,N_8106);
or UO_871 (O_871,N_9982,N_8041);
nor UO_872 (O_872,N_8140,N_9923);
nor UO_873 (O_873,N_8864,N_9886);
or UO_874 (O_874,N_9264,N_9904);
nor UO_875 (O_875,N_8011,N_9536);
nor UO_876 (O_876,N_8211,N_9680);
nand UO_877 (O_877,N_8988,N_9774);
xor UO_878 (O_878,N_9802,N_8237);
nor UO_879 (O_879,N_8202,N_8540);
or UO_880 (O_880,N_8976,N_9235);
nand UO_881 (O_881,N_9287,N_8730);
nand UO_882 (O_882,N_8343,N_9826);
and UO_883 (O_883,N_8939,N_8300);
nand UO_884 (O_884,N_9055,N_9003);
xnor UO_885 (O_885,N_9198,N_9249);
xor UO_886 (O_886,N_9697,N_9761);
or UO_887 (O_887,N_8192,N_9319);
xor UO_888 (O_888,N_9156,N_9808);
nand UO_889 (O_889,N_9480,N_9133);
nor UO_890 (O_890,N_9751,N_9267);
nor UO_891 (O_891,N_8752,N_9804);
xor UO_892 (O_892,N_8849,N_9785);
or UO_893 (O_893,N_9200,N_8605);
and UO_894 (O_894,N_8588,N_8388);
nor UO_895 (O_895,N_8556,N_9888);
nor UO_896 (O_896,N_9962,N_8382);
and UO_897 (O_897,N_8004,N_8371);
nand UO_898 (O_898,N_9389,N_9985);
or UO_899 (O_899,N_9691,N_8075);
or UO_900 (O_900,N_9036,N_9230);
or UO_901 (O_901,N_9117,N_8442);
and UO_902 (O_902,N_8980,N_9424);
and UO_903 (O_903,N_9899,N_8095);
xor UO_904 (O_904,N_9884,N_8625);
and UO_905 (O_905,N_9288,N_8013);
and UO_906 (O_906,N_8150,N_9443);
nand UO_907 (O_907,N_8707,N_8250);
or UO_908 (O_908,N_9369,N_8402);
and UO_909 (O_909,N_9407,N_9457);
and UO_910 (O_910,N_8952,N_9195);
nor UO_911 (O_911,N_8585,N_8197);
and UO_912 (O_912,N_9993,N_9461);
nand UO_913 (O_913,N_9318,N_8889);
or UO_914 (O_914,N_8695,N_8483);
or UO_915 (O_915,N_9729,N_9158);
or UO_916 (O_916,N_9216,N_9330);
and UO_917 (O_917,N_9331,N_9940);
nand UO_918 (O_918,N_9995,N_9061);
or UO_919 (O_919,N_8705,N_9441);
xor UO_920 (O_920,N_8139,N_8144);
nor UO_921 (O_921,N_9526,N_9469);
or UO_922 (O_922,N_9557,N_9935);
nor UO_923 (O_923,N_8935,N_9281);
nand UO_924 (O_924,N_9020,N_9236);
nor UO_925 (O_925,N_8738,N_9722);
nor UO_926 (O_926,N_8994,N_9822);
or UO_927 (O_927,N_8201,N_9749);
nor UO_928 (O_928,N_8983,N_9108);
or UO_929 (O_929,N_8770,N_8247);
and UO_930 (O_930,N_9654,N_9191);
and UO_931 (O_931,N_8547,N_8831);
nor UO_932 (O_932,N_9041,N_9662);
nand UO_933 (O_933,N_8527,N_9919);
and UO_934 (O_934,N_9260,N_8999);
nand UO_935 (O_935,N_8241,N_9228);
nand UO_936 (O_936,N_9889,N_9014);
nor UO_937 (O_937,N_9606,N_9510);
and UO_938 (O_938,N_9965,N_9132);
xnor UO_939 (O_939,N_8709,N_8113);
and UO_940 (O_940,N_9928,N_9734);
nor UO_941 (O_941,N_8065,N_8724);
nor UO_942 (O_942,N_9710,N_8109);
or UO_943 (O_943,N_8230,N_8998);
and UO_944 (O_944,N_8909,N_9008);
nand UO_945 (O_945,N_9182,N_8006);
and UO_946 (O_946,N_8164,N_8455);
or UO_947 (O_947,N_9296,N_8231);
nand UO_948 (O_948,N_8505,N_9334);
and UO_949 (O_949,N_8971,N_8014);
nand UO_950 (O_950,N_8024,N_8986);
and UO_951 (O_951,N_9896,N_8639);
or UO_952 (O_952,N_8059,N_9069);
and UO_953 (O_953,N_9603,N_9168);
nor UO_954 (O_954,N_8595,N_8764);
nand UO_955 (O_955,N_8641,N_9206);
xor UO_956 (O_956,N_9032,N_8824);
and UO_957 (O_957,N_8594,N_8456);
nor UO_958 (O_958,N_8892,N_9277);
nand UO_959 (O_959,N_9668,N_8083);
nand UO_960 (O_960,N_8403,N_9171);
and UO_961 (O_961,N_9563,N_9542);
nand UO_962 (O_962,N_8678,N_9658);
nand UO_963 (O_963,N_8516,N_9579);
or UO_964 (O_964,N_9421,N_9618);
xnor UO_965 (O_965,N_8694,N_9086);
nor UO_966 (O_966,N_8386,N_9197);
nand UO_967 (O_967,N_8227,N_8350);
or UO_968 (O_968,N_8997,N_9640);
or UO_969 (O_969,N_9590,N_8240);
or UO_970 (O_970,N_8655,N_9022);
nand UO_971 (O_971,N_8785,N_8592);
or UO_972 (O_972,N_9218,N_8380);
nor UO_973 (O_973,N_8917,N_9308);
xor UO_974 (O_974,N_9750,N_8136);
and UO_975 (O_975,N_8010,N_8827);
or UO_976 (O_976,N_9037,N_8070);
or UO_977 (O_977,N_8725,N_8734);
and UO_978 (O_978,N_9535,N_8458);
nand UO_979 (O_979,N_9740,N_8790);
or UO_980 (O_980,N_8383,N_8578);
xnor UO_981 (O_981,N_9807,N_9189);
nand UO_982 (O_982,N_8168,N_9177);
nand UO_983 (O_983,N_9815,N_9152);
nand UO_984 (O_984,N_9382,N_9992);
nor UO_985 (O_985,N_8387,N_8185);
and UO_986 (O_986,N_9174,N_9374);
and UO_987 (O_987,N_8287,N_9852);
nor UO_988 (O_988,N_9306,N_8063);
nor UO_989 (O_989,N_9865,N_8837);
nor UO_990 (O_990,N_9315,N_9781);
nor UO_991 (O_991,N_9360,N_9048);
nand UO_992 (O_992,N_9341,N_9849);
and UO_993 (O_993,N_9289,N_8334);
xnor UO_994 (O_994,N_8208,N_9827);
nand UO_995 (O_995,N_9464,N_8204);
or UO_996 (O_996,N_8990,N_9121);
nand UO_997 (O_997,N_8826,N_8060);
nand UO_998 (O_998,N_9977,N_8974);
nor UO_999 (O_999,N_9273,N_8172);
or UO_1000 (O_1000,N_8578,N_9596);
and UO_1001 (O_1001,N_9285,N_9127);
or UO_1002 (O_1002,N_8700,N_9531);
or UO_1003 (O_1003,N_9575,N_8101);
nand UO_1004 (O_1004,N_9520,N_8300);
nor UO_1005 (O_1005,N_9934,N_8165);
or UO_1006 (O_1006,N_9343,N_8437);
or UO_1007 (O_1007,N_9616,N_8367);
or UO_1008 (O_1008,N_8755,N_8023);
nor UO_1009 (O_1009,N_8036,N_8542);
and UO_1010 (O_1010,N_8558,N_8203);
nand UO_1011 (O_1011,N_8046,N_9655);
nor UO_1012 (O_1012,N_9305,N_8995);
nor UO_1013 (O_1013,N_8701,N_8167);
xor UO_1014 (O_1014,N_8890,N_8461);
or UO_1015 (O_1015,N_8603,N_9243);
nor UO_1016 (O_1016,N_8867,N_8043);
or UO_1017 (O_1017,N_8162,N_9620);
nor UO_1018 (O_1018,N_9430,N_9316);
nor UO_1019 (O_1019,N_9369,N_8797);
and UO_1020 (O_1020,N_8917,N_8647);
or UO_1021 (O_1021,N_9210,N_9769);
or UO_1022 (O_1022,N_9128,N_8824);
and UO_1023 (O_1023,N_8543,N_8075);
xor UO_1024 (O_1024,N_8283,N_8881);
or UO_1025 (O_1025,N_8136,N_8660);
and UO_1026 (O_1026,N_8518,N_9924);
and UO_1027 (O_1027,N_8323,N_8487);
nand UO_1028 (O_1028,N_8138,N_8843);
nor UO_1029 (O_1029,N_9497,N_9915);
and UO_1030 (O_1030,N_8701,N_8942);
nor UO_1031 (O_1031,N_8307,N_9454);
nor UO_1032 (O_1032,N_9428,N_8300);
xnor UO_1033 (O_1033,N_8635,N_9869);
nor UO_1034 (O_1034,N_8712,N_8168);
xor UO_1035 (O_1035,N_9435,N_8103);
nand UO_1036 (O_1036,N_8830,N_8722);
nor UO_1037 (O_1037,N_8767,N_8149);
nor UO_1038 (O_1038,N_9928,N_8181);
or UO_1039 (O_1039,N_9685,N_8060);
and UO_1040 (O_1040,N_9061,N_8885);
xnor UO_1041 (O_1041,N_8956,N_8454);
nand UO_1042 (O_1042,N_8654,N_8458);
and UO_1043 (O_1043,N_9124,N_9340);
and UO_1044 (O_1044,N_8095,N_9673);
and UO_1045 (O_1045,N_9469,N_8051);
nand UO_1046 (O_1046,N_8347,N_8061);
nor UO_1047 (O_1047,N_9142,N_8427);
or UO_1048 (O_1048,N_8343,N_8178);
or UO_1049 (O_1049,N_8443,N_9099);
or UO_1050 (O_1050,N_9431,N_9563);
nand UO_1051 (O_1051,N_8944,N_9918);
and UO_1052 (O_1052,N_9676,N_8532);
and UO_1053 (O_1053,N_8540,N_9136);
or UO_1054 (O_1054,N_9466,N_8243);
nor UO_1055 (O_1055,N_9721,N_8866);
or UO_1056 (O_1056,N_9357,N_9325);
nand UO_1057 (O_1057,N_8849,N_8237);
nand UO_1058 (O_1058,N_8144,N_8318);
nand UO_1059 (O_1059,N_9127,N_8585);
nor UO_1060 (O_1060,N_9454,N_9840);
and UO_1061 (O_1061,N_9786,N_9746);
and UO_1062 (O_1062,N_8251,N_8168);
nor UO_1063 (O_1063,N_8704,N_8938);
nand UO_1064 (O_1064,N_8802,N_9727);
nor UO_1065 (O_1065,N_8541,N_9049);
and UO_1066 (O_1066,N_8701,N_9179);
xor UO_1067 (O_1067,N_8718,N_9426);
or UO_1068 (O_1068,N_8404,N_9791);
and UO_1069 (O_1069,N_9139,N_8255);
xor UO_1070 (O_1070,N_9197,N_8113);
nor UO_1071 (O_1071,N_8386,N_8400);
nor UO_1072 (O_1072,N_8380,N_9826);
nor UO_1073 (O_1073,N_8440,N_9761);
or UO_1074 (O_1074,N_9186,N_8808);
or UO_1075 (O_1075,N_9321,N_8034);
nand UO_1076 (O_1076,N_9509,N_9210);
xnor UO_1077 (O_1077,N_9071,N_8742);
nor UO_1078 (O_1078,N_9063,N_9173);
or UO_1079 (O_1079,N_9541,N_8206);
nor UO_1080 (O_1080,N_9512,N_8177);
nand UO_1081 (O_1081,N_8683,N_9961);
nor UO_1082 (O_1082,N_9004,N_9403);
xnor UO_1083 (O_1083,N_8956,N_9488);
nor UO_1084 (O_1084,N_9838,N_8799);
or UO_1085 (O_1085,N_8074,N_8436);
nand UO_1086 (O_1086,N_9296,N_8235);
nand UO_1087 (O_1087,N_9766,N_8582);
nand UO_1088 (O_1088,N_8624,N_9481);
nor UO_1089 (O_1089,N_9196,N_8909);
and UO_1090 (O_1090,N_9906,N_9295);
and UO_1091 (O_1091,N_9500,N_8976);
and UO_1092 (O_1092,N_9339,N_8761);
nor UO_1093 (O_1093,N_8649,N_8582);
xnor UO_1094 (O_1094,N_9986,N_9918);
xor UO_1095 (O_1095,N_8938,N_9000);
nand UO_1096 (O_1096,N_9577,N_8221);
nor UO_1097 (O_1097,N_9502,N_8092);
xor UO_1098 (O_1098,N_8926,N_9289);
and UO_1099 (O_1099,N_9295,N_8900);
nand UO_1100 (O_1100,N_9245,N_8490);
or UO_1101 (O_1101,N_8237,N_8346);
and UO_1102 (O_1102,N_9319,N_9695);
or UO_1103 (O_1103,N_9320,N_9782);
xnor UO_1104 (O_1104,N_8647,N_8112);
and UO_1105 (O_1105,N_8258,N_9359);
nand UO_1106 (O_1106,N_8917,N_9277);
or UO_1107 (O_1107,N_8312,N_9837);
nor UO_1108 (O_1108,N_9509,N_9881);
nor UO_1109 (O_1109,N_8049,N_9112);
nand UO_1110 (O_1110,N_8527,N_8095);
and UO_1111 (O_1111,N_8079,N_8115);
and UO_1112 (O_1112,N_9222,N_8333);
nand UO_1113 (O_1113,N_9297,N_9677);
nor UO_1114 (O_1114,N_8811,N_8056);
or UO_1115 (O_1115,N_9055,N_9608);
nor UO_1116 (O_1116,N_9260,N_8981);
and UO_1117 (O_1117,N_8871,N_8692);
nand UO_1118 (O_1118,N_8057,N_8328);
nor UO_1119 (O_1119,N_9025,N_9595);
nor UO_1120 (O_1120,N_9129,N_8379);
nand UO_1121 (O_1121,N_8021,N_8754);
nor UO_1122 (O_1122,N_9099,N_8731);
nand UO_1123 (O_1123,N_8144,N_9705);
and UO_1124 (O_1124,N_9532,N_8370);
and UO_1125 (O_1125,N_8831,N_9937);
nor UO_1126 (O_1126,N_9008,N_9999);
nor UO_1127 (O_1127,N_8532,N_8214);
nand UO_1128 (O_1128,N_8796,N_9166);
nand UO_1129 (O_1129,N_8831,N_9983);
and UO_1130 (O_1130,N_8650,N_9475);
nor UO_1131 (O_1131,N_8488,N_9994);
xnor UO_1132 (O_1132,N_8637,N_9458);
nand UO_1133 (O_1133,N_9168,N_8623);
or UO_1134 (O_1134,N_8767,N_9642);
nor UO_1135 (O_1135,N_9470,N_8871);
nor UO_1136 (O_1136,N_8092,N_8455);
xor UO_1137 (O_1137,N_8693,N_9673);
or UO_1138 (O_1138,N_9139,N_9199);
nor UO_1139 (O_1139,N_8004,N_9980);
nand UO_1140 (O_1140,N_9643,N_8994);
or UO_1141 (O_1141,N_9540,N_8135);
or UO_1142 (O_1142,N_9969,N_9708);
nand UO_1143 (O_1143,N_9947,N_8007);
or UO_1144 (O_1144,N_9858,N_8994);
xor UO_1145 (O_1145,N_8258,N_8092);
nand UO_1146 (O_1146,N_9641,N_9844);
and UO_1147 (O_1147,N_9542,N_8567);
or UO_1148 (O_1148,N_8689,N_9293);
nor UO_1149 (O_1149,N_9134,N_8234);
and UO_1150 (O_1150,N_9625,N_9611);
or UO_1151 (O_1151,N_8269,N_9605);
and UO_1152 (O_1152,N_9753,N_9585);
and UO_1153 (O_1153,N_8941,N_8919);
nor UO_1154 (O_1154,N_8691,N_9249);
and UO_1155 (O_1155,N_8647,N_9291);
and UO_1156 (O_1156,N_9430,N_9368);
xnor UO_1157 (O_1157,N_9466,N_9805);
xnor UO_1158 (O_1158,N_9710,N_8939);
or UO_1159 (O_1159,N_9690,N_8857);
and UO_1160 (O_1160,N_8309,N_8092);
nor UO_1161 (O_1161,N_9259,N_9170);
and UO_1162 (O_1162,N_9914,N_9198);
xor UO_1163 (O_1163,N_8243,N_9540);
or UO_1164 (O_1164,N_9329,N_8734);
or UO_1165 (O_1165,N_9659,N_8648);
and UO_1166 (O_1166,N_9325,N_8694);
nor UO_1167 (O_1167,N_8614,N_9537);
and UO_1168 (O_1168,N_9977,N_8055);
and UO_1169 (O_1169,N_8705,N_8471);
or UO_1170 (O_1170,N_9566,N_8720);
or UO_1171 (O_1171,N_9659,N_8864);
nor UO_1172 (O_1172,N_9378,N_9942);
nor UO_1173 (O_1173,N_8196,N_8531);
or UO_1174 (O_1174,N_8540,N_8949);
nand UO_1175 (O_1175,N_8434,N_9701);
nor UO_1176 (O_1176,N_9962,N_9640);
or UO_1177 (O_1177,N_8471,N_8105);
nand UO_1178 (O_1178,N_9330,N_8527);
xnor UO_1179 (O_1179,N_9815,N_8968);
nor UO_1180 (O_1180,N_9909,N_8931);
xnor UO_1181 (O_1181,N_9982,N_9628);
nor UO_1182 (O_1182,N_9698,N_9895);
or UO_1183 (O_1183,N_8412,N_9438);
nand UO_1184 (O_1184,N_8057,N_8909);
or UO_1185 (O_1185,N_9001,N_9269);
nand UO_1186 (O_1186,N_8560,N_9386);
or UO_1187 (O_1187,N_9078,N_9248);
and UO_1188 (O_1188,N_9244,N_8626);
nor UO_1189 (O_1189,N_9188,N_8908);
nand UO_1190 (O_1190,N_8099,N_9896);
nor UO_1191 (O_1191,N_9662,N_9883);
and UO_1192 (O_1192,N_9783,N_8677);
xnor UO_1193 (O_1193,N_9637,N_8867);
or UO_1194 (O_1194,N_8722,N_8871);
nand UO_1195 (O_1195,N_9842,N_8797);
and UO_1196 (O_1196,N_9272,N_8149);
or UO_1197 (O_1197,N_8322,N_9003);
xor UO_1198 (O_1198,N_9931,N_8396);
nand UO_1199 (O_1199,N_9315,N_8530);
or UO_1200 (O_1200,N_9107,N_9064);
nand UO_1201 (O_1201,N_8697,N_9342);
nor UO_1202 (O_1202,N_9357,N_8271);
nor UO_1203 (O_1203,N_8996,N_9896);
xnor UO_1204 (O_1204,N_9837,N_9836);
or UO_1205 (O_1205,N_9241,N_8505);
nor UO_1206 (O_1206,N_8513,N_8411);
xor UO_1207 (O_1207,N_8812,N_8212);
nand UO_1208 (O_1208,N_8831,N_8037);
nor UO_1209 (O_1209,N_9537,N_8670);
and UO_1210 (O_1210,N_8358,N_9157);
nand UO_1211 (O_1211,N_9729,N_9642);
or UO_1212 (O_1212,N_9487,N_8993);
or UO_1213 (O_1213,N_8403,N_8684);
or UO_1214 (O_1214,N_8262,N_9853);
and UO_1215 (O_1215,N_9228,N_8295);
nor UO_1216 (O_1216,N_9703,N_8497);
nand UO_1217 (O_1217,N_8828,N_9000);
nand UO_1218 (O_1218,N_8954,N_9396);
nor UO_1219 (O_1219,N_8149,N_8287);
nand UO_1220 (O_1220,N_8753,N_8711);
and UO_1221 (O_1221,N_9582,N_9905);
or UO_1222 (O_1222,N_8148,N_9949);
and UO_1223 (O_1223,N_8682,N_8975);
xor UO_1224 (O_1224,N_9506,N_8987);
nor UO_1225 (O_1225,N_8562,N_8071);
nor UO_1226 (O_1226,N_9724,N_9016);
nor UO_1227 (O_1227,N_8530,N_8900);
xor UO_1228 (O_1228,N_8319,N_8446);
nor UO_1229 (O_1229,N_8747,N_8231);
and UO_1230 (O_1230,N_8624,N_8537);
or UO_1231 (O_1231,N_8496,N_9640);
or UO_1232 (O_1232,N_8893,N_9172);
and UO_1233 (O_1233,N_9092,N_9373);
nor UO_1234 (O_1234,N_8402,N_9165);
nand UO_1235 (O_1235,N_8195,N_9478);
nand UO_1236 (O_1236,N_9276,N_9127);
nor UO_1237 (O_1237,N_9630,N_9910);
nor UO_1238 (O_1238,N_9309,N_9194);
and UO_1239 (O_1239,N_9739,N_8734);
nand UO_1240 (O_1240,N_8645,N_8891);
and UO_1241 (O_1241,N_8615,N_8071);
nand UO_1242 (O_1242,N_8700,N_9872);
nor UO_1243 (O_1243,N_9206,N_9630);
xor UO_1244 (O_1244,N_8156,N_9193);
or UO_1245 (O_1245,N_9905,N_9280);
nand UO_1246 (O_1246,N_9991,N_9538);
nor UO_1247 (O_1247,N_8954,N_8073);
nor UO_1248 (O_1248,N_9155,N_9635);
and UO_1249 (O_1249,N_8165,N_8922);
or UO_1250 (O_1250,N_8374,N_8111);
nand UO_1251 (O_1251,N_8135,N_9593);
and UO_1252 (O_1252,N_9897,N_8557);
and UO_1253 (O_1253,N_8290,N_9817);
nor UO_1254 (O_1254,N_8793,N_8567);
and UO_1255 (O_1255,N_9926,N_8429);
nor UO_1256 (O_1256,N_9351,N_9576);
nor UO_1257 (O_1257,N_8272,N_9860);
nand UO_1258 (O_1258,N_8249,N_8063);
xor UO_1259 (O_1259,N_8538,N_8672);
nand UO_1260 (O_1260,N_8426,N_8132);
xnor UO_1261 (O_1261,N_9292,N_9221);
nor UO_1262 (O_1262,N_9164,N_8490);
nor UO_1263 (O_1263,N_8613,N_9734);
nand UO_1264 (O_1264,N_9305,N_8277);
or UO_1265 (O_1265,N_9143,N_9103);
or UO_1266 (O_1266,N_9691,N_8719);
nor UO_1267 (O_1267,N_9297,N_8781);
and UO_1268 (O_1268,N_9689,N_9532);
nand UO_1269 (O_1269,N_9284,N_8706);
or UO_1270 (O_1270,N_9417,N_8101);
xnor UO_1271 (O_1271,N_8646,N_8893);
nand UO_1272 (O_1272,N_8743,N_9221);
xor UO_1273 (O_1273,N_8680,N_9093);
and UO_1274 (O_1274,N_9695,N_9341);
and UO_1275 (O_1275,N_9157,N_9580);
nand UO_1276 (O_1276,N_9277,N_8221);
or UO_1277 (O_1277,N_9146,N_9841);
nor UO_1278 (O_1278,N_8072,N_8858);
and UO_1279 (O_1279,N_9253,N_9448);
nor UO_1280 (O_1280,N_9147,N_9075);
or UO_1281 (O_1281,N_8859,N_8448);
nor UO_1282 (O_1282,N_8456,N_8884);
or UO_1283 (O_1283,N_9632,N_9753);
nand UO_1284 (O_1284,N_8152,N_8289);
or UO_1285 (O_1285,N_9622,N_9982);
nor UO_1286 (O_1286,N_8103,N_8868);
xnor UO_1287 (O_1287,N_9108,N_8043);
or UO_1288 (O_1288,N_8984,N_9589);
nor UO_1289 (O_1289,N_8240,N_8335);
and UO_1290 (O_1290,N_8072,N_9205);
and UO_1291 (O_1291,N_9731,N_9089);
nor UO_1292 (O_1292,N_9960,N_9547);
and UO_1293 (O_1293,N_8653,N_8536);
nand UO_1294 (O_1294,N_8505,N_8610);
or UO_1295 (O_1295,N_9267,N_9756);
and UO_1296 (O_1296,N_9957,N_8638);
and UO_1297 (O_1297,N_9712,N_9063);
and UO_1298 (O_1298,N_9469,N_8041);
nand UO_1299 (O_1299,N_8338,N_9832);
nor UO_1300 (O_1300,N_9642,N_8540);
or UO_1301 (O_1301,N_9094,N_9475);
xnor UO_1302 (O_1302,N_8758,N_8184);
or UO_1303 (O_1303,N_8139,N_8808);
or UO_1304 (O_1304,N_9667,N_8624);
and UO_1305 (O_1305,N_8093,N_8455);
and UO_1306 (O_1306,N_9827,N_9225);
xor UO_1307 (O_1307,N_9702,N_8585);
nor UO_1308 (O_1308,N_8134,N_8975);
nand UO_1309 (O_1309,N_9611,N_9395);
nor UO_1310 (O_1310,N_9920,N_8541);
nor UO_1311 (O_1311,N_9093,N_9419);
xor UO_1312 (O_1312,N_9560,N_8798);
or UO_1313 (O_1313,N_9878,N_9556);
xnor UO_1314 (O_1314,N_9008,N_9741);
or UO_1315 (O_1315,N_9997,N_9414);
and UO_1316 (O_1316,N_9933,N_9448);
nand UO_1317 (O_1317,N_9455,N_9033);
nor UO_1318 (O_1318,N_9631,N_8032);
nor UO_1319 (O_1319,N_9029,N_8276);
nor UO_1320 (O_1320,N_8579,N_8068);
or UO_1321 (O_1321,N_8248,N_9787);
or UO_1322 (O_1322,N_9425,N_9390);
nor UO_1323 (O_1323,N_8600,N_9259);
and UO_1324 (O_1324,N_9570,N_8909);
nor UO_1325 (O_1325,N_9896,N_8055);
or UO_1326 (O_1326,N_9794,N_8722);
nor UO_1327 (O_1327,N_8318,N_8129);
nand UO_1328 (O_1328,N_9706,N_8831);
and UO_1329 (O_1329,N_8368,N_8173);
nand UO_1330 (O_1330,N_8938,N_8560);
nand UO_1331 (O_1331,N_9115,N_9485);
nand UO_1332 (O_1332,N_8093,N_9667);
xnor UO_1333 (O_1333,N_9907,N_9212);
nor UO_1334 (O_1334,N_9757,N_8245);
nor UO_1335 (O_1335,N_8602,N_8198);
nand UO_1336 (O_1336,N_9257,N_8847);
nor UO_1337 (O_1337,N_8007,N_8983);
nor UO_1338 (O_1338,N_9149,N_9492);
nor UO_1339 (O_1339,N_9903,N_9932);
or UO_1340 (O_1340,N_8749,N_9844);
nor UO_1341 (O_1341,N_9699,N_9769);
or UO_1342 (O_1342,N_9519,N_8547);
nor UO_1343 (O_1343,N_8974,N_9663);
and UO_1344 (O_1344,N_8827,N_9706);
nand UO_1345 (O_1345,N_9827,N_9306);
nand UO_1346 (O_1346,N_9680,N_8139);
and UO_1347 (O_1347,N_9630,N_9101);
and UO_1348 (O_1348,N_8562,N_9246);
or UO_1349 (O_1349,N_8575,N_9561);
nand UO_1350 (O_1350,N_8917,N_9809);
nor UO_1351 (O_1351,N_9636,N_8186);
xnor UO_1352 (O_1352,N_9337,N_8667);
and UO_1353 (O_1353,N_9231,N_9755);
and UO_1354 (O_1354,N_9821,N_9741);
nor UO_1355 (O_1355,N_9601,N_9840);
and UO_1356 (O_1356,N_8882,N_9177);
or UO_1357 (O_1357,N_8026,N_9664);
and UO_1358 (O_1358,N_8295,N_9122);
nor UO_1359 (O_1359,N_8987,N_8680);
nand UO_1360 (O_1360,N_8195,N_8045);
or UO_1361 (O_1361,N_8147,N_8578);
or UO_1362 (O_1362,N_8143,N_8221);
xor UO_1363 (O_1363,N_8581,N_8010);
nor UO_1364 (O_1364,N_9918,N_9882);
nand UO_1365 (O_1365,N_8259,N_8784);
or UO_1366 (O_1366,N_9152,N_9626);
nor UO_1367 (O_1367,N_9849,N_9913);
and UO_1368 (O_1368,N_8248,N_9160);
or UO_1369 (O_1369,N_8740,N_8686);
or UO_1370 (O_1370,N_9666,N_9109);
or UO_1371 (O_1371,N_9283,N_9404);
nor UO_1372 (O_1372,N_9081,N_9670);
or UO_1373 (O_1373,N_8128,N_9495);
nor UO_1374 (O_1374,N_8344,N_8354);
nor UO_1375 (O_1375,N_8963,N_9598);
or UO_1376 (O_1376,N_8056,N_8626);
nand UO_1377 (O_1377,N_8397,N_9567);
nor UO_1378 (O_1378,N_8591,N_8006);
nor UO_1379 (O_1379,N_8962,N_9749);
and UO_1380 (O_1380,N_9014,N_9058);
nand UO_1381 (O_1381,N_8679,N_9894);
nor UO_1382 (O_1382,N_8044,N_8347);
nand UO_1383 (O_1383,N_9835,N_8855);
nand UO_1384 (O_1384,N_8325,N_9162);
xor UO_1385 (O_1385,N_8974,N_8471);
nor UO_1386 (O_1386,N_9341,N_9113);
or UO_1387 (O_1387,N_9322,N_9044);
and UO_1388 (O_1388,N_8603,N_8491);
xnor UO_1389 (O_1389,N_8352,N_9437);
nor UO_1390 (O_1390,N_8159,N_8537);
nor UO_1391 (O_1391,N_8779,N_9427);
nor UO_1392 (O_1392,N_8127,N_9288);
nand UO_1393 (O_1393,N_8259,N_9913);
and UO_1394 (O_1394,N_8447,N_9835);
and UO_1395 (O_1395,N_9074,N_9269);
nand UO_1396 (O_1396,N_9402,N_8640);
and UO_1397 (O_1397,N_9980,N_9992);
and UO_1398 (O_1398,N_9732,N_9889);
and UO_1399 (O_1399,N_9507,N_8461);
or UO_1400 (O_1400,N_8246,N_9110);
xnor UO_1401 (O_1401,N_9343,N_9021);
and UO_1402 (O_1402,N_8068,N_9967);
xor UO_1403 (O_1403,N_9478,N_9118);
nand UO_1404 (O_1404,N_9721,N_9433);
nor UO_1405 (O_1405,N_9260,N_8909);
and UO_1406 (O_1406,N_9163,N_8647);
or UO_1407 (O_1407,N_9042,N_9402);
xnor UO_1408 (O_1408,N_8136,N_9740);
or UO_1409 (O_1409,N_9672,N_9309);
and UO_1410 (O_1410,N_8152,N_8067);
nor UO_1411 (O_1411,N_8889,N_9900);
xnor UO_1412 (O_1412,N_8162,N_8531);
or UO_1413 (O_1413,N_9079,N_9813);
xor UO_1414 (O_1414,N_8152,N_9632);
or UO_1415 (O_1415,N_9942,N_9557);
xor UO_1416 (O_1416,N_9261,N_9601);
or UO_1417 (O_1417,N_9967,N_8023);
or UO_1418 (O_1418,N_9604,N_9558);
nand UO_1419 (O_1419,N_8167,N_8486);
and UO_1420 (O_1420,N_9745,N_9191);
xor UO_1421 (O_1421,N_9683,N_8253);
or UO_1422 (O_1422,N_9539,N_9516);
or UO_1423 (O_1423,N_8131,N_9830);
or UO_1424 (O_1424,N_9932,N_9558);
or UO_1425 (O_1425,N_9783,N_8037);
nor UO_1426 (O_1426,N_8277,N_9911);
xnor UO_1427 (O_1427,N_8488,N_8414);
nor UO_1428 (O_1428,N_9480,N_8024);
nor UO_1429 (O_1429,N_9843,N_8601);
nand UO_1430 (O_1430,N_9862,N_9181);
nor UO_1431 (O_1431,N_9593,N_8932);
and UO_1432 (O_1432,N_8133,N_8039);
xor UO_1433 (O_1433,N_8669,N_8632);
nand UO_1434 (O_1434,N_9453,N_9417);
nor UO_1435 (O_1435,N_8593,N_9936);
nand UO_1436 (O_1436,N_8158,N_9717);
or UO_1437 (O_1437,N_9125,N_9032);
nand UO_1438 (O_1438,N_9983,N_8627);
nand UO_1439 (O_1439,N_8526,N_9488);
nand UO_1440 (O_1440,N_8653,N_8725);
or UO_1441 (O_1441,N_9476,N_8708);
or UO_1442 (O_1442,N_8269,N_8205);
nand UO_1443 (O_1443,N_9413,N_8684);
xnor UO_1444 (O_1444,N_9368,N_9702);
and UO_1445 (O_1445,N_9953,N_8243);
xnor UO_1446 (O_1446,N_9502,N_8809);
or UO_1447 (O_1447,N_8317,N_9267);
and UO_1448 (O_1448,N_9391,N_8166);
xor UO_1449 (O_1449,N_8458,N_9590);
or UO_1450 (O_1450,N_8713,N_8187);
nor UO_1451 (O_1451,N_8378,N_8517);
nor UO_1452 (O_1452,N_9875,N_9775);
nand UO_1453 (O_1453,N_9217,N_9863);
or UO_1454 (O_1454,N_9682,N_9298);
nand UO_1455 (O_1455,N_9985,N_9002);
nor UO_1456 (O_1456,N_8008,N_9729);
nand UO_1457 (O_1457,N_9400,N_8211);
and UO_1458 (O_1458,N_9824,N_9113);
xor UO_1459 (O_1459,N_8995,N_9106);
nand UO_1460 (O_1460,N_9064,N_9852);
and UO_1461 (O_1461,N_9559,N_9016);
nand UO_1462 (O_1462,N_8359,N_8038);
or UO_1463 (O_1463,N_9819,N_8320);
or UO_1464 (O_1464,N_8935,N_9496);
and UO_1465 (O_1465,N_8694,N_9342);
and UO_1466 (O_1466,N_9452,N_9471);
nand UO_1467 (O_1467,N_9960,N_9543);
xor UO_1468 (O_1468,N_9027,N_8032);
and UO_1469 (O_1469,N_8426,N_9653);
and UO_1470 (O_1470,N_9430,N_8348);
nor UO_1471 (O_1471,N_8738,N_8159);
nand UO_1472 (O_1472,N_8799,N_8528);
nand UO_1473 (O_1473,N_8923,N_9804);
nand UO_1474 (O_1474,N_9957,N_8127);
or UO_1475 (O_1475,N_9842,N_8450);
nor UO_1476 (O_1476,N_9446,N_9692);
and UO_1477 (O_1477,N_8008,N_8779);
nand UO_1478 (O_1478,N_9289,N_9182);
or UO_1479 (O_1479,N_9574,N_9012);
and UO_1480 (O_1480,N_9028,N_8454);
nor UO_1481 (O_1481,N_9555,N_9181);
nand UO_1482 (O_1482,N_9570,N_9792);
or UO_1483 (O_1483,N_8128,N_9812);
or UO_1484 (O_1484,N_9764,N_9587);
nor UO_1485 (O_1485,N_9156,N_8467);
nand UO_1486 (O_1486,N_9996,N_8216);
nand UO_1487 (O_1487,N_9322,N_9285);
and UO_1488 (O_1488,N_9293,N_8746);
nand UO_1489 (O_1489,N_9011,N_9809);
or UO_1490 (O_1490,N_8303,N_9913);
nor UO_1491 (O_1491,N_8206,N_8490);
nand UO_1492 (O_1492,N_8162,N_9523);
and UO_1493 (O_1493,N_8950,N_8913);
or UO_1494 (O_1494,N_9977,N_8221);
nand UO_1495 (O_1495,N_9121,N_9671);
xnor UO_1496 (O_1496,N_8506,N_8915);
or UO_1497 (O_1497,N_8912,N_9913);
and UO_1498 (O_1498,N_8671,N_9808);
nor UO_1499 (O_1499,N_8522,N_9679);
endmodule